module basic_5000_50000_5000_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_147,In_1836);
and U1 (N_1,In_672,In_2509);
nand U2 (N_2,In_1466,In_623);
nand U3 (N_3,In_1801,In_2727);
nor U4 (N_4,In_2313,In_1661);
and U5 (N_5,In_2012,In_4924);
nor U6 (N_6,In_4716,In_4199);
and U7 (N_7,In_2411,In_2144);
xnor U8 (N_8,In_4145,In_395);
nand U9 (N_9,In_4976,In_4484);
nand U10 (N_10,In_517,In_3791);
nand U11 (N_11,In_1142,In_3840);
and U12 (N_12,In_3368,In_896);
or U13 (N_13,In_4703,In_797);
nor U14 (N_14,In_4657,In_1697);
xor U15 (N_15,In_1886,In_1257);
or U16 (N_16,In_4286,In_2353);
nand U17 (N_17,In_67,In_1820);
and U18 (N_18,In_3403,In_3871);
nand U19 (N_19,In_2369,In_2889);
or U20 (N_20,In_2883,In_951);
nor U21 (N_21,In_3991,In_944);
and U22 (N_22,In_2090,In_3646);
and U23 (N_23,In_557,In_2361);
xor U24 (N_24,In_2760,In_1734);
or U25 (N_25,In_1550,In_2895);
nand U26 (N_26,In_680,In_283);
nor U27 (N_27,In_1402,In_2828);
and U28 (N_28,In_3141,In_4784);
nor U29 (N_29,In_749,In_4335);
and U30 (N_30,In_4333,In_3808);
xor U31 (N_31,In_4517,In_4215);
and U32 (N_32,In_4800,In_2673);
or U33 (N_33,In_134,In_4537);
and U34 (N_34,In_800,In_4000);
and U35 (N_35,In_4123,In_465);
nand U36 (N_36,In_1792,In_3425);
nand U37 (N_37,In_3032,In_3708);
nor U38 (N_38,In_622,In_1669);
nand U39 (N_39,In_231,In_3535);
and U40 (N_40,In_3561,In_4229);
nand U41 (N_41,In_563,In_97);
xor U42 (N_42,In_1290,In_2972);
or U43 (N_43,In_1396,In_4995);
nand U44 (N_44,In_1410,In_1101);
or U45 (N_45,In_3742,In_3539);
xor U46 (N_46,In_4167,In_2503);
xor U47 (N_47,In_2933,In_253);
nor U48 (N_48,In_459,In_2851);
and U49 (N_49,In_1742,In_4826);
nor U50 (N_50,In_4701,In_685);
xor U51 (N_51,In_1058,In_4266);
and U52 (N_52,In_19,In_4090);
and U53 (N_53,In_2885,In_3471);
nor U54 (N_54,In_2970,In_3634);
nor U55 (N_55,In_1007,In_2077);
xor U56 (N_56,In_1537,In_3467);
and U57 (N_57,In_3518,In_2608);
and U58 (N_58,In_2706,In_1393);
and U59 (N_59,In_1242,In_4219);
xnor U60 (N_60,In_3302,In_16);
and U61 (N_61,In_3743,In_142);
xor U62 (N_62,In_1804,In_3470);
nor U63 (N_63,In_4283,In_2835);
nand U64 (N_64,In_171,In_3906);
nand U65 (N_65,In_870,In_1429);
nor U66 (N_66,In_1654,In_3855);
nor U67 (N_67,In_2942,In_1508);
or U68 (N_68,In_2722,In_1911);
or U69 (N_69,In_3792,In_977);
or U70 (N_70,In_3321,In_1525);
and U71 (N_71,In_129,In_3845);
and U72 (N_72,In_637,In_2508);
or U73 (N_73,In_4550,In_3714);
and U74 (N_74,In_1602,In_3515);
or U75 (N_75,In_3418,In_2534);
nand U76 (N_76,In_1065,In_2242);
xnor U77 (N_77,In_1825,In_3622);
or U78 (N_78,In_4601,In_2935);
nor U79 (N_79,In_2291,In_3129);
nand U80 (N_80,In_2341,In_3605);
nand U81 (N_81,In_411,In_393);
nand U82 (N_82,In_510,In_1044);
nand U83 (N_83,In_577,In_58);
and U84 (N_84,In_3484,In_1133);
or U85 (N_85,In_3147,In_4241);
and U86 (N_86,In_1965,In_4788);
nor U87 (N_87,In_3200,In_948);
or U88 (N_88,In_3932,In_2670);
and U89 (N_89,In_1373,In_1326);
or U90 (N_90,In_966,In_3199);
nand U91 (N_91,In_2538,In_2060);
xor U92 (N_92,In_3268,In_120);
nor U93 (N_93,In_2629,In_3657);
and U94 (N_94,In_4693,In_3364);
nand U95 (N_95,In_2097,In_1307);
nor U96 (N_96,In_2631,In_519);
xor U97 (N_97,In_4503,In_2698);
xnor U98 (N_98,In_3987,In_3434);
nand U99 (N_99,In_2480,In_1263);
xor U100 (N_100,In_2403,In_1366);
xnor U101 (N_101,In_3435,In_2100);
nand U102 (N_102,In_4098,In_2159);
nor U103 (N_103,In_550,In_2019);
or U104 (N_104,In_2875,In_1013);
xor U105 (N_105,In_354,In_773);
xor U106 (N_106,In_3257,In_4817);
or U107 (N_107,In_2894,In_4099);
and U108 (N_108,In_2607,In_3398);
or U109 (N_109,In_4152,In_3514);
xor U110 (N_110,In_2719,In_382);
nand U111 (N_111,In_2276,In_151);
nand U112 (N_112,In_879,In_2917);
nand U113 (N_113,In_4481,In_953);
nor U114 (N_114,In_2452,In_3087);
nor U115 (N_115,In_4758,In_3395);
xnor U116 (N_116,In_1706,In_3860);
nor U117 (N_117,In_3079,In_1968);
and U118 (N_118,In_2767,In_3633);
and U119 (N_119,In_4709,In_289);
xor U120 (N_120,In_4393,In_4822);
and U121 (N_121,In_514,In_3239);
xnor U122 (N_122,In_2737,In_4223);
nor U123 (N_123,In_38,In_3626);
nand U124 (N_124,In_2869,In_3360);
and U125 (N_125,In_2168,In_1122);
nor U126 (N_126,In_370,In_1980);
xnor U127 (N_127,In_905,In_2213);
nand U128 (N_128,In_2056,In_2667);
nor U129 (N_129,In_4454,In_4058);
or U130 (N_130,In_2375,In_858);
xor U131 (N_131,In_217,In_1251);
or U132 (N_132,In_4607,In_3649);
or U133 (N_133,In_3267,In_3084);
and U134 (N_134,In_644,In_2442);
nand U135 (N_135,In_154,In_3055);
xor U136 (N_136,In_2026,In_4105);
or U137 (N_137,In_2797,In_1030);
nand U138 (N_138,In_2592,In_1931);
and U139 (N_139,In_3061,In_1763);
and U140 (N_140,In_2799,In_4136);
and U141 (N_141,In_578,In_2426);
nand U142 (N_142,In_983,In_36);
nor U143 (N_143,In_326,In_4463);
and U144 (N_144,In_1880,In_2622);
or U145 (N_145,In_1424,In_2418);
or U146 (N_146,In_2841,In_1423);
or U147 (N_147,In_1566,In_551);
or U148 (N_148,In_3009,In_1505);
nand U149 (N_149,In_1492,In_1561);
nor U150 (N_150,In_1805,In_4009);
and U151 (N_151,In_4018,In_1253);
nand U152 (N_152,In_3503,In_320);
nor U153 (N_153,In_1649,In_1309);
and U154 (N_154,In_3441,In_4113);
xnor U155 (N_155,In_2932,In_85);
nand U156 (N_156,In_566,In_4272);
nand U157 (N_157,In_2323,In_346);
nand U158 (N_158,In_2469,In_4328);
and U159 (N_159,In_1962,In_3121);
nor U160 (N_160,In_1448,In_1428);
nor U161 (N_161,In_4727,In_4101);
nand U162 (N_162,In_3986,In_4411);
nor U163 (N_163,In_2890,In_3988);
and U164 (N_164,In_1964,In_4008);
or U165 (N_165,In_2048,In_3002);
nand U166 (N_166,In_544,In_3540);
xor U167 (N_167,In_4653,In_2316);
nand U168 (N_168,In_2396,In_1589);
nand U169 (N_169,In_3495,In_814);
nand U170 (N_170,In_923,In_3075);
nor U171 (N_171,In_4271,In_774);
nand U172 (N_172,In_2888,In_1304);
or U173 (N_173,In_3182,In_4862);
or U174 (N_174,In_3105,In_4978);
and U175 (N_175,In_493,In_929);
and U176 (N_176,In_4831,In_2043);
nand U177 (N_177,In_4336,In_4348);
and U178 (N_178,In_299,In_1540);
and U179 (N_179,In_1231,In_3191);
xor U180 (N_180,In_3137,In_43);
xor U181 (N_181,In_2794,In_281);
nand U182 (N_182,In_3511,In_4143);
nor U183 (N_183,In_3553,In_3946);
nand U184 (N_184,In_2179,In_787);
nand U185 (N_185,In_2416,In_3872);
xor U186 (N_186,In_3071,In_2188);
and U187 (N_187,In_3729,In_4933);
nand U188 (N_188,In_1728,In_634);
nor U189 (N_189,In_4694,In_790);
nand U190 (N_190,In_529,In_1370);
nand U191 (N_191,In_4226,In_3548);
nor U192 (N_192,In_1614,In_389);
nand U193 (N_193,In_3064,In_4710);
xnor U194 (N_194,In_2856,In_1786);
or U195 (N_195,In_18,In_3285);
nor U196 (N_196,In_4796,In_3314);
nand U197 (N_197,In_2867,In_2032);
nor U198 (N_198,In_4093,In_4876);
nand U199 (N_199,In_198,In_3361);
nor U200 (N_200,In_831,In_3139);
and U201 (N_201,In_3751,In_702);
or U202 (N_202,In_1340,In_2123);
xnor U203 (N_203,In_1571,In_1362);
nand U204 (N_204,In_1882,In_1703);
nor U205 (N_205,In_4501,In_3858);
nor U206 (N_206,In_3393,In_2581);
or U207 (N_207,In_2387,In_1765);
or U208 (N_208,In_1311,In_2300);
xor U209 (N_209,In_4474,In_1730);
nand U210 (N_210,In_4061,In_2813);
nor U211 (N_211,In_3215,In_4449);
or U212 (N_212,In_4104,In_973);
nand U213 (N_213,In_2904,In_2674);
nand U214 (N_214,In_3336,In_4031);
nor U215 (N_215,In_1636,In_2107);
xnor U216 (N_216,In_1102,In_4803);
or U217 (N_217,In_3480,In_2065);
nor U218 (N_218,In_4905,In_418);
or U219 (N_219,In_4736,In_2456);
or U220 (N_220,In_4857,In_338);
nor U221 (N_221,In_4786,In_2236);
nor U222 (N_222,In_294,In_1633);
nor U223 (N_223,In_2591,In_829);
or U224 (N_224,In_2712,In_3221);
and U225 (N_225,In_3297,In_1105);
nand U226 (N_226,In_3530,In_4288);
and U227 (N_227,In_3311,In_4611);
and U228 (N_228,In_2891,In_2114);
and U229 (N_229,In_943,In_832);
or U230 (N_230,In_3236,In_4824);
xnor U231 (N_231,In_928,In_4198);
or U232 (N_232,In_4030,In_4749);
and U233 (N_233,In_205,In_282);
nand U234 (N_234,In_705,In_2069);
nor U235 (N_235,In_4951,In_3893);
nand U236 (N_236,In_2818,In_3342);
or U237 (N_237,In_871,In_161);
and U238 (N_238,In_3213,In_2080);
nor U239 (N_239,In_603,In_838);
xnor U240 (N_240,In_2800,In_4497);
xnor U241 (N_241,In_1790,In_4609);
nand U242 (N_242,In_2016,In_2170);
and U243 (N_243,In_2998,In_1539);
or U244 (N_244,In_2253,In_89);
and U245 (N_245,In_3831,In_1045);
nor U246 (N_246,In_887,In_3173);
nor U247 (N_247,In_3572,In_4006);
and U248 (N_248,In_474,In_410);
or U249 (N_249,In_4029,In_1859);
nor U250 (N_250,In_2413,In_850);
nand U251 (N_251,In_3357,In_287);
nand U252 (N_252,In_2965,In_2180);
xnor U253 (N_253,In_606,In_4785);
nor U254 (N_254,In_1659,In_1708);
nor U255 (N_255,In_4878,In_3911);
or U256 (N_256,In_249,In_3809);
nand U257 (N_257,In_2333,In_4274);
and U258 (N_258,In_4513,In_582);
nor U259 (N_259,In_2600,In_4913);
or U260 (N_260,In_3431,In_988);
or U261 (N_261,In_1470,In_1710);
nand U262 (N_262,In_237,In_837);
nor U263 (N_263,In_4419,In_3091);
or U264 (N_264,In_3458,In_1346);
nor U265 (N_265,In_3867,In_4997);
nor U266 (N_266,In_4869,In_2512);
nand U267 (N_267,In_559,In_1764);
xor U268 (N_268,In_1134,In_525);
nand U269 (N_269,In_2284,In_2819);
xor U270 (N_270,In_1951,In_4433);
nand U271 (N_271,In_3177,In_15);
or U272 (N_272,In_2140,In_3619);
nand U273 (N_273,In_2587,In_2146);
and U274 (N_274,In_818,In_4263);
nor U275 (N_275,In_376,In_8);
and U276 (N_276,In_1642,In_1660);
nor U277 (N_277,In_4806,In_2775);
or U278 (N_278,In_1611,In_3167);
nor U279 (N_279,In_4069,In_2269);
and U280 (N_280,In_1475,In_378);
or U281 (N_281,In_271,In_27);
nor U282 (N_282,In_3376,In_3273);
nand U283 (N_283,In_3135,In_4131);
nor U284 (N_284,In_4895,In_4154);
or U285 (N_285,In_4868,In_4702);
and U286 (N_286,In_4354,In_1500);
and U287 (N_287,In_4516,In_1536);
nor U288 (N_288,In_737,In_4776);
xor U289 (N_289,In_4442,In_1834);
xnor U290 (N_290,In_2204,In_4401);
and U291 (N_291,In_1843,In_979);
xnor U292 (N_292,In_3735,In_761);
or U293 (N_293,In_821,In_2964);
and U294 (N_294,In_3026,In_3485);
or U295 (N_295,In_1979,In_3081);
xnor U296 (N_296,In_4511,In_3020);
nor U297 (N_297,In_3278,In_3262);
or U298 (N_298,In_2514,In_1892);
or U299 (N_299,In_427,In_2331);
nor U300 (N_300,In_3916,In_3122);
or U301 (N_301,In_1835,In_4346);
nor U302 (N_302,In_1054,In_2870);
xnor U303 (N_303,In_1680,In_1897);
nor U304 (N_304,In_3781,In_645);
nor U305 (N_305,In_2211,In_1063);
nor U306 (N_306,In_2934,In_3505);
nor U307 (N_307,In_325,In_23);
nand U308 (N_308,In_1782,In_830);
nor U309 (N_309,In_4221,In_941);
nor U310 (N_310,In_4084,In_3195);
nor U311 (N_311,In_4282,In_4841);
nor U312 (N_312,In_1844,In_2913);
and U313 (N_313,In_1993,In_2944);
nand U314 (N_314,In_2381,In_3320);
xnor U315 (N_315,In_1502,In_2435);
nand U316 (N_316,In_788,In_3385);
nor U317 (N_317,In_1573,In_137);
nor U318 (N_318,In_3259,In_189);
nand U319 (N_319,In_4811,In_2268);
nand U320 (N_320,In_1905,In_2379);
xnor U321 (N_321,In_1119,In_4875);
nor U322 (N_322,In_1281,In_1450);
and U323 (N_323,In_3876,In_3538);
and U324 (N_324,In_1890,In_4003);
and U325 (N_325,In_497,In_856);
xor U326 (N_326,In_4999,In_351);
and U327 (N_327,In_4420,In_4952);
nand U328 (N_328,In_4486,In_3717);
nor U329 (N_329,In_4573,In_3152);
xnor U330 (N_330,In_95,In_158);
or U331 (N_331,In_2928,In_3163);
and U332 (N_332,In_2185,In_2303);
or U333 (N_333,In_3698,In_4002);
nor U334 (N_334,In_4279,In_2786);
or U335 (N_335,In_2318,In_3789);
nor U336 (N_336,In_1084,In_236);
and U337 (N_337,In_3638,In_3062);
and U338 (N_338,In_847,In_2617);
nor U339 (N_339,In_1895,In_4043);
or U340 (N_340,In_4208,In_2919);
xor U341 (N_341,In_347,In_1598);
xor U342 (N_342,In_1230,In_3856);
xnor U343 (N_343,In_3018,In_4122);
xnor U344 (N_344,In_1077,In_1438);
or U345 (N_345,In_4415,In_3896);
or U346 (N_346,In_1607,In_4965);
xnor U347 (N_347,In_3914,In_697);
and U348 (N_348,In_3424,In_1998);
nor U349 (N_349,In_2866,In_934);
nand U350 (N_350,In_1451,In_854);
or U351 (N_351,In_4262,In_267);
or U352 (N_352,In_2085,In_1940);
xor U353 (N_353,In_1696,In_4410);
and U354 (N_354,In_2848,In_324);
nor U355 (N_355,In_2768,In_1707);
or U356 (N_356,In_3296,In_460);
xor U357 (N_357,In_3125,In_2504);
nor U358 (N_358,In_2730,In_696);
nor U359 (N_359,In_1535,In_4319);
nand U360 (N_360,In_2422,In_4790);
or U361 (N_361,In_453,In_4494);
or U362 (N_362,In_54,In_1797);
nor U363 (N_363,In_2606,In_4050);
or U364 (N_364,In_3188,In_413);
and U365 (N_365,In_4287,In_540);
nand U366 (N_366,In_107,In_4626);
or U367 (N_367,In_3145,In_2155);
nand U368 (N_368,In_3041,In_3693);
nand U369 (N_369,In_1096,In_2531);
xor U370 (N_370,In_2152,In_3124);
nand U371 (N_371,In_2930,In_3235);
nor U372 (N_372,In_1773,In_1411);
nand U373 (N_373,In_125,In_4576);
and U374 (N_374,In_4931,In_579);
and U375 (N_375,In_846,In_2654);
nor U376 (N_376,In_972,In_3593);
or U377 (N_377,In_3536,In_1595);
nand U378 (N_378,In_914,In_2227);
and U379 (N_379,In_3740,In_3306);
and U380 (N_380,In_4659,In_528);
xor U381 (N_381,In_3596,In_4349);
nor U382 (N_382,In_4480,In_3254);
or U383 (N_383,In_4548,In_2642);
xnor U384 (N_384,In_2363,In_4252);
nor U385 (N_385,In_2311,In_2054);
or U386 (N_386,In_3029,In_1568);
or U387 (N_387,In_1893,In_4887);
nand U388 (N_388,In_3017,In_4555);
nor U389 (N_389,In_1435,In_4707);
nand U390 (N_390,In_946,In_1186);
nand U391 (N_391,In_1196,In_1856);
nand U392 (N_392,In_1594,In_2241);
nor U393 (N_393,In_4673,In_1870);
xnor U394 (N_394,In_1567,In_4042);
or U395 (N_395,In_3687,In_4755);
xnor U396 (N_396,In_1228,In_4178);
nand U397 (N_397,In_2494,In_3701);
or U398 (N_398,In_3624,In_280);
or U399 (N_399,In_1970,In_39);
nand U400 (N_400,In_4744,In_3115);
and U401 (N_401,In_4840,In_756);
xor U402 (N_402,In_648,In_3172);
or U403 (N_403,In_3941,In_1829);
nor U404 (N_404,In_3716,In_1533);
xnor U405 (N_405,In_2506,In_4981);
and U406 (N_406,In_166,In_2424);
nand U407 (N_407,In_3318,In_50);
nand U408 (N_408,In_3885,In_2612);
nand U409 (N_409,In_1275,In_1343);
nand U410 (N_410,In_4129,In_3774);
nand U411 (N_411,In_3734,In_3192);
and U412 (N_412,In_4450,In_511);
nor U413 (N_413,In_2075,In_2182);
xor U414 (N_414,In_2249,In_4763);
and U415 (N_415,In_2939,In_3448);
or U416 (N_416,In_3256,In_4374);
nand U417 (N_417,In_4426,In_1896);
nor U418 (N_418,In_4519,In_4406);
nand U419 (N_419,In_4455,In_1158);
and U420 (N_420,In_580,In_2840);
xnor U421 (N_421,In_422,In_52);
or U422 (N_422,In_2126,In_4205);
nand U423 (N_423,In_4149,In_4545);
and U424 (N_424,In_4212,In_2973);
and U425 (N_425,In_1928,In_2738);
nor U426 (N_426,In_4813,In_4430);
nor U427 (N_427,In_4473,In_3761);
nand U428 (N_428,In_2092,In_3577);
nor U429 (N_429,In_1456,In_621);
nand U430 (N_430,In_1436,In_2036);
and U431 (N_431,In_633,In_2390);
xor U432 (N_432,In_175,In_2920);
and U433 (N_433,In_1552,In_3689);
and U434 (N_434,In_2620,In_4327);
or U435 (N_435,In_3578,In_1264);
nand U436 (N_436,In_954,In_259);
nor U437 (N_437,In_646,In_429);
nand U438 (N_438,In_1916,In_2257);
and U439 (N_439,In_3620,In_288);
nor U440 (N_440,In_1591,In_3479);
and U441 (N_441,In_4565,In_1314);
nor U442 (N_442,In_3848,In_2559);
nand U443 (N_443,In_2334,In_1496);
or U444 (N_444,In_3658,In_467);
or U445 (N_445,In_1222,In_4357);
and U446 (N_446,In_573,In_796);
and U447 (N_447,In_2486,In_4649);
or U448 (N_448,In_679,In_2646);
nor U449 (N_449,In_2164,In_574);
nor U450 (N_450,In_4405,In_218);
xor U451 (N_451,In_342,In_3030);
and U452 (N_452,In_3834,In_415);
and U453 (N_453,In_55,In_3552);
nor U454 (N_454,In_4569,In_2338);
xnor U455 (N_455,In_3008,In_2493);
xnor U456 (N_456,In_3294,In_2199);
and U457 (N_457,In_1061,In_1898);
nor U458 (N_458,In_1506,In_152);
nand U459 (N_459,In_690,In_808);
or U460 (N_460,In_3951,In_1732);
or U461 (N_461,In_3207,In_4360);
and U462 (N_462,In_1503,In_651);
xor U463 (N_463,In_1912,In_1827);
nor U464 (N_464,In_1254,In_2438);
and U465 (N_465,In_4371,In_4834);
nand U466 (N_466,In_848,In_3884);
nand U467 (N_467,In_3563,In_968);
and U468 (N_468,In_2811,In_1983);
xor U469 (N_469,In_4838,In_1043);
xnor U470 (N_470,In_1809,In_2321);
nor U471 (N_471,In_1215,In_4828);
or U472 (N_472,In_3979,In_666);
or U473 (N_473,In_4487,In_4423);
xnor U474 (N_474,In_2298,In_4893);
nor U475 (N_475,In_74,In_1627);
nor U476 (N_476,In_2415,In_1305);
and U477 (N_477,In_4603,In_3021);
or U478 (N_478,In_1592,In_664);
or U479 (N_479,In_1619,In_2791);
nand U480 (N_480,In_629,In_715);
nand U481 (N_481,In_2002,In_286);
xnor U482 (N_482,In_4285,In_233);
nor U483 (N_483,In_4805,In_4139);
and U484 (N_484,In_2425,In_4705);
and U485 (N_485,In_2844,In_4134);
and U486 (N_486,In_4089,In_179);
nor U487 (N_487,In_2771,In_3377);
nand U488 (N_488,In_3274,In_4164);
nor U489 (N_489,In_3901,In_1783);
or U490 (N_490,In_2150,In_3110);
or U491 (N_491,In_2058,In_581);
or U492 (N_492,In_4459,In_2529);
nor U493 (N_493,In_3132,In_4067);
or U494 (N_494,In_2769,In_3089);
nand U495 (N_495,In_3948,In_2167);
and U496 (N_496,In_2033,In_2011);
nand U497 (N_497,In_555,In_261);
and U498 (N_498,In_3963,In_755);
nand U499 (N_499,In_2235,In_3463);
xor U500 (N_500,In_263,In_2874);
nand U501 (N_501,In_1067,In_4369);
nand U502 (N_502,In_1877,In_1048);
xnor U503 (N_503,In_3873,In_2757);
nor U504 (N_504,In_4213,In_319);
and U505 (N_505,In_1579,In_2232);
nand U506 (N_506,In_4258,In_4617);
nand U507 (N_507,In_3654,In_2325);
and U508 (N_508,In_298,In_2393);
nand U509 (N_509,In_4257,In_2658);
and U510 (N_510,In_3183,In_3114);
and U511 (N_511,In_3555,In_2556);
xor U512 (N_512,In_469,In_588);
and U513 (N_513,In_396,In_2838);
xnor U514 (N_514,In_1034,In_674);
nor U515 (N_515,In_40,In_4019);
and U516 (N_516,In_2250,In_1819);
or U517 (N_517,In_182,In_1012);
and U518 (N_518,In_3928,In_1513);
and U519 (N_519,In_3420,In_485);
xnor U520 (N_520,In_1398,In_1079);
or U521 (N_521,In_1319,In_3971);
xnor U522 (N_522,In_2400,In_3526);
nand U523 (N_523,In_103,In_3304);
or U524 (N_524,In_183,In_1555);
nand U525 (N_525,In_883,In_2899);
or U526 (N_526,In_4827,In_1073);
or U527 (N_527,In_616,In_4500);
and U528 (N_528,In_1840,In_1772);
nand U529 (N_529,In_906,In_4842);
nand U530 (N_530,In_1616,In_1179);
nor U531 (N_531,In_2320,In_613);
xor U532 (N_532,In_3205,In_2410);
or U533 (N_533,In_374,In_735);
or U534 (N_534,In_1081,In_1511);
nor U535 (N_535,In_4639,In_245);
nand U536 (N_536,In_2878,In_4294);
nor U537 (N_537,In_1194,In_3949);
or U538 (N_538,In_3892,In_4938);
nand U539 (N_539,In_1368,In_1883);
xor U540 (N_540,In_90,In_4233);
nand U541 (N_541,In_3144,In_3350);
nand U542 (N_542,In_2279,In_1243);
nor U543 (N_543,In_212,In_1872);
nor U544 (N_544,In_3373,In_2383);
or U545 (N_545,In_1651,In_1051);
and U546 (N_546,In_3338,In_4529);
nand U547 (N_547,In_345,In_291);
nor U548 (N_548,In_3639,In_1107);
xnor U549 (N_549,In_902,In_817);
and U550 (N_550,In_4413,In_3090);
and U551 (N_551,In_4446,In_2812);
or U552 (N_552,In_3665,In_3732);
nor U553 (N_553,In_113,In_3117);
and U554 (N_554,In_3814,In_4015);
nand U555 (N_555,In_4435,In_2849);
nand U556 (N_556,In_1881,In_4525);
xor U557 (N_557,In_3753,In_2348);
nor U558 (N_558,In_4175,In_2308);
xor U559 (N_559,In_9,In_2655);
or U560 (N_560,In_4391,In_4969);
nand U561 (N_561,In_3838,In_47);
xor U562 (N_562,In_2062,In_2478);
nor U563 (N_563,In_2831,In_4083);
nor U564 (N_564,In_3721,In_72);
xnor U565 (N_565,In_3568,In_1632);
nor U566 (N_566,In_3462,In_14);
and U567 (N_567,In_1498,In_509);
xnor U568 (N_568,In_3575,In_1794);
nand U569 (N_569,In_3417,In_4290);
nor U570 (N_570,In_869,In_251);
xor U571 (N_571,In_3457,In_2863);
nor U572 (N_572,In_3047,In_4836);
xnor U573 (N_573,In_24,In_3547);
xnor U574 (N_574,In_2611,In_4663);
and U575 (N_575,In_150,In_2575);
nand U576 (N_576,In_2482,In_4124);
xor U577 (N_577,In_4119,In_3541);
xor U578 (N_578,In_3439,In_2368);
nand U579 (N_579,In_4536,In_3123);
and U580 (N_580,In_2850,In_2490);
or U581 (N_581,In_2548,In_1449);
nor U582 (N_582,In_3322,In_730);
nor U583 (N_583,In_4771,In_1260);
xnor U584 (N_584,In_1578,In_1325);
or U585 (N_585,In_2349,In_2703);
xnor U586 (N_586,In_227,In_1355);
nor U587 (N_587,In_4078,In_3673);
xor U588 (N_588,In_1437,In_3460);
or U589 (N_589,In_3497,In_4192);
nor U590 (N_590,In_1586,In_3899);
nor U591 (N_591,In_4665,In_2963);
xor U592 (N_592,In_4608,In_1780);
nor U593 (N_593,In_2560,In_1295);
nand U594 (N_594,In_1433,In_184);
nand U595 (N_595,In_4186,In_388);
xnor U596 (N_596,In_860,In_3094);
nor U597 (N_597,In_2277,In_3204);
or U598 (N_598,In_3961,In_2326);
or U599 (N_599,In_1767,In_489);
nor U600 (N_600,In_2623,In_3113);
xor U601 (N_601,In_1403,In_1);
or U602 (N_602,In_3813,In_3027);
or U603 (N_603,In_3168,In_207);
or U604 (N_604,In_3203,In_1664);
or U605 (N_605,In_4216,In_507);
nand U606 (N_606,In_2082,In_4345);
nor U607 (N_607,In_1570,In_4849);
nand U608 (N_608,In_1686,In_1369);
or U609 (N_609,In_2709,In_3607);
and U610 (N_610,In_1170,In_4970);
or U611 (N_611,In_486,In_3788);
nand U612 (N_612,In_2634,In_2713);
nand U613 (N_613,In_1480,In_1838);
or U614 (N_614,In_1933,In_1672);
xor U615 (N_615,In_1313,In_3883);
nor U616 (N_616,In_4993,In_2163);
or U617 (N_617,In_1676,In_4142);
nand U618 (N_618,In_2013,In_4724);
nand U619 (N_619,In_4530,In_1556);
xnor U620 (N_620,In_3052,In_430);
xor U621 (N_621,In_1903,In_1320);
xnor U622 (N_622,In_296,In_3613);
xor U623 (N_623,In_4355,In_1564);
nor U624 (N_624,In_3022,In_2796);
and U625 (N_625,In_2562,In_2527);
and U626 (N_626,In_1648,In_2772);
nor U627 (N_627,In_4467,In_3891);
nand U628 (N_628,In_3214,In_4927);
nor U629 (N_629,In_4769,In_4443);
nor U630 (N_630,In_2519,In_1816);
and U631 (N_631,In_1737,In_2224);
nor U632 (N_632,In_1489,In_3245);
nand U633 (N_633,In_1738,In_1959);
nor U634 (N_634,In_268,In_4239);
and U635 (N_635,In_3001,In_862);
nor U636 (N_636,In_2817,In_1984);
xnor U637 (N_637,In_1127,In_2409);
nor U638 (N_638,In_3606,In_1291);
nor U639 (N_639,In_1027,In_2597);
nor U640 (N_640,In_1954,In_105);
and U641 (N_641,In_1683,In_4585);
and U642 (N_642,In_4631,In_34);
xnor U643 (N_643,In_3625,In_4498);
or U644 (N_644,In_2975,In_4708);
nand U645 (N_645,In_806,In_2541);
xnor U646 (N_646,In_2647,In_1997);
xor U647 (N_647,In_3817,In_3587);
nand U648 (N_648,In_3266,In_4958);
xnor U649 (N_649,In_4818,In_1799);
nand U650 (N_650,In_4384,In_400);
and U651 (N_651,In_4133,In_3768);
nand U652 (N_652,In_3033,In_1640);
and U653 (N_653,In_4350,In_247);
xnor U654 (N_654,In_855,In_4379);
xor U655 (N_655,In_1289,In_2350);
xor U656 (N_656,In_377,In_533);
nand U657 (N_657,In_3007,In_2023);
nor U658 (N_658,In_1157,In_1606);
nand U659 (N_659,In_3863,In_2266);
nor U660 (N_660,In_2726,In_587);
nand U661 (N_661,In_3136,In_4725);
and U662 (N_662,In_2859,In_4322);
or U663 (N_663,In_4602,In_1025);
or U664 (N_664,In_4889,In_1670);
xnor U665 (N_665,In_295,In_2621);
nand U666 (N_666,In_44,In_4546);
and U667 (N_667,In_2051,In_2347);
nor U668 (N_668,In_119,In_4988);
or U669 (N_669,In_1245,In_1863);
and U670 (N_670,In_22,In_1445);
xor U671 (N_671,In_3551,In_4801);
nand U672 (N_672,In_3579,In_609);
nand U673 (N_673,In_1944,In_1176);
xnor U674 (N_674,In_3058,In_1615);
nor U675 (N_675,In_190,In_35);
nor U676 (N_676,In_2672,In_420);
nand U677 (N_677,In_2448,In_3284);
xor U678 (N_678,In_234,In_976);
and U679 (N_679,In_4808,In_1292);
nand U680 (N_680,In_434,In_3);
and U681 (N_681,In_4852,In_172);
or U682 (N_682,In_3942,In_4921);
nor U683 (N_683,In_4163,In_3252);
xnor U684 (N_684,In_4650,In_3486);
nor U685 (N_685,In_2255,In_3651);
and U686 (N_686,In_2367,In_1971);
or U687 (N_687,In_604,In_3574);
xor U688 (N_688,In_2549,In_3851);
xnor U689 (N_689,In_596,In_1562);
nand U690 (N_690,In_1509,In_4306);
xor U691 (N_691,In_4044,In_1006);
xor U692 (N_692,In_1652,In_1237);
and U693 (N_693,In_1351,In_3394);
nand U694 (N_694,In_1848,In_1705);
and U695 (N_695,In_3787,In_138);
nand U696 (N_696,In_794,In_4116);
nand U697 (N_697,In_1851,In_2927);
nand U698 (N_698,In_1140,In_2830);
nand U699 (N_699,In_2958,In_2789);
nor U700 (N_700,In_2099,In_11);
or U701 (N_701,In_4385,In_691);
nor U702 (N_702,In_3315,In_4111);
or U703 (N_703,In_4676,In_4597);
or U704 (N_704,In_2045,In_2461);
or U705 (N_705,In_1258,In_2217);
nand U706 (N_706,In_1922,In_2414);
and U707 (N_707,In_4033,In_1609);
and U708 (N_708,In_2441,In_4839);
or U709 (N_709,In_4690,In_2025);
xnor U710 (N_710,In_1490,In_3456);
xor U711 (N_711,In_3006,In_594);
nor U712 (N_712,In_68,In_4340);
and U713 (N_713,In_3286,In_1798);
or U714 (N_714,In_1285,In_2892);
and U715 (N_715,In_3158,In_4972);
or U716 (N_716,In_516,In_1294);
xor U717 (N_717,In_4583,In_57);
and U718 (N_718,In_4886,In_2024);
or U719 (N_719,In_3407,In_4132);
xnor U720 (N_720,In_328,In_4815);
or U721 (N_721,In_1138,In_3869);
xnor U722 (N_722,In_1557,In_335);
nor U723 (N_723,In_2487,In_4049);
xnor U724 (N_724,In_1232,In_1286);
or U725 (N_725,In_3422,In_4949);
nand U726 (N_726,In_741,In_3450);
and U727 (N_727,In_3190,In_1748);
and U728 (N_728,In_4483,In_4307);
or U729 (N_729,In_4013,In_3359);
nor U730 (N_730,In_4447,In_1658);
xor U731 (N_731,In_2793,In_4331);
or U732 (N_732,In_1753,In_2267);
or U733 (N_733,In_4194,In_1235);
xnor U734 (N_734,In_155,In_3309);
nand U735 (N_735,In_2485,In_3220);
nor U736 (N_736,In_1832,In_1280);
and U737 (N_737,In_2820,In_1149);
nand U738 (N_738,In_3216,In_1118);
or U739 (N_739,In_4488,In_3637);
xor U740 (N_740,In_202,In_4353);
or U741 (N_741,In_2136,In_4157);
nor U742 (N_742,In_1937,In_1418);
nand U743 (N_743,In_4751,In_1390);
and U744 (N_744,In_1941,In_2281);
and U745 (N_745,In_4961,In_2259);
and U746 (N_746,In_1657,In_2115);
or U747 (N_747,In_4270,In_1775);
and U748 (N_748,In_1349,In_1715);
or U749 (N_749,In_1688,In_1183);
xor U750 (N_750,In_3573,In_4037);
or U751 (N_751,In_4738,In_4863);
nor U752 (N_752,In_3260,In_4882);
xor U753 (N_753,In_2008,In_4679);
nand U754 (N_754,In_2955,In_962);
nor U755 (N_755,In_4193,In_4623);
and U756 (N_756,In_2143,In_2020);
and U757 (N_757,In_1274,In_2953);
or U758 (N_758,In_4173,In_4695);
or U759 (N_759,In_1647,In_3162);
nor U760 (N_760,In_2103,In_228);
nor U761 (N_761,In_1404,In_4733);
xor U762 (N_762,In_1849,In_2868);
or U763 (N_763,In_3782,In_2921);
xnor U764 (N_764,In_723,In_2704);
nand U765 (N_765,In_2806,In_3864);
xnor U766 (N_766,In_1327,In_2364);
xor U767 (N_767,In_2022,In_2651);
xnor U768 (N_768,In_2271,In_4432);
and U769 (N_769,In_4246,In_1910);
xnor U770 (N_770,In_3882,In_936);
xor U771 (N_771,In_45,In_909);
xnor U772 (N_772,In_4217,In_1995);
and U773 (N_773,In_3715,In_3586);
xor U774 (N_774,In_1620,In_2206);
or U775 (N_775,In_4661,In_2433);
and U776 (N_776,In_964,In_823);
nand U777 (N_777,In_2785,In_310);
or U778 (N_778,In_73,In_2044);
nand U779 (N_779,In_704,In_1581);
and U780 (N_780,In_1066,In_3498);
and U781 (N_781,In_4466,In_1784);
and U782 (N_782,In_4196,In_2070);
nand U783 (N_783,In_3647,In_2344);
or U784 (N_784,In_1926,In_3410);
xor U785 (N_785,In_4383,In_404);
and U786 (N_786,In_156,In_3842);
or U787 (N_787,In_1414,In_4745);
nor U788 (N_788,In_1103,In_2710);
nor U789 (N_789,In_3584,In_4475);
and U790 (N_790,In_2699,In_1088);
nand U791 (N_791,In_2488,In_593);
nand U792 (N_792,In_258,In_4866);
or U793 (N_793,In_2650,In_3242);
xor U794 (N_794,In_624,In_1419);
xnor U795 (N_795,In_3962,In_3844);
or U796 (N_796,In_3074,In_3472);
or U797 (N_797,In_121,In_70);
nand U798 (N_798,In_717,In_4176);
nor U799 (N_799,In_31,In_708);
nor U800 (N_800,In_1766,In_4341);
nand U801 (N_801,In_3815,In_4251);
nor U802 (N_802,In_543,In_3543);
xnor U803 (N_803,In_2501,In_352);
xor U804 (N_804,In_3046,In_2040);
and U805 (N_805,In_284,In_4916);
nand U806 (N_806,In_3493,In_4747);
or U807 (N_807,In_2453,In_4259);
and U808 (N_808,In_1454,In_2111);
nand U809 (N_809,In_1634,In_1873);
or U810 (N_810,In_3179,In_4510);
or U811 (N_811,In_3108,In_2815);
and U812 (N_812,In_4641,In_2059);
nand U813 (N_813,In_4458,In_1518);
xnor U814 (N_814,In_3793,In_3012);
and U815 (N_815,In_2265,In_2225);
xnor U816 (N_816,In_3250,In_4461);
nor U817 (N_817,In_2916,In_4871);
or U818 (N_818,In_2550,In_3015);
or U819 (N_819,In_2021,In_3779);
xnor U820 (N_820,In_562,In_2102);
xor U821 (N_821,In_3662,In_2668);
nand U822 (N_822,In_4774,In_2429);
or U823 (N_823,In_764,In_3875);
nor U824 (N_824,In_3825,In_1348);
and U825 (N_825,In_2572,In_269);
nand U826 (N_826,In_2089,In_2676);
nor U827 (N_827,In_759,In_4575);
or U828 (N_828,In_640,In_315);
nor U829 (N_829,In_1850,In_3853);
or U830 (N_830,In_3580,In_512);
nor U831 (N_831,In_1986,In_3667);
or U832 (N_832,In_312,In_3354);
nor U833 (N_833,In_3777,In_1526);
nand U834 (N_834,In_3972,In_1335);
and U835 (N_835,In_499,In_3668);
nand U836 (N_836,In_3968,In_952);
or U837 (N_837,In_475,In_4441);
and U838 (N_838,In_4877,In_2362);
xnor U839 (N_839,In_2173,In_4606);
or U840 (N_840,In_3704,In_2076);
nor U841 (N_841,In_4936,In_340);
or U842 (N_842,In_1206,In_2784);
xor U843 (N_843,In_128,In_1582);
nand U844 (N_844,In_1098,In_3341);
xor U845 (N_845,In_192,In_548);
nand U846 (N_846,In_2352,In_625);
or U847 (N_847,In_3237,In_3756);
or U848 (N_848,In_165,In_4566);
or U849 (N_849,In_1227,In_1412);
xor U850 (N_850,In_1247,In_4932);
or U851 (N_851,In_3727,In_561);
and U852 (N_852,In_3201,In_1646);
nor U853 (N_853,In_482,In_3165);
and U854 (N_854,In_2980,In_130);
or U855 (N_855,In_1392,In_2081);
nor U856 (N_856,In_1769,In_820);
xnor U857 (N_857,In_479,In_3253);
xnor U858 (N_858,In_3386,In_3677);
nand U859 (N_859,In_2565,In_975);
xnor U860 (N_860,In_4362,In_894);
nor U861 (N_861,In_60,In_4558);
and U862 (N_862,In_508,In_3421);
xnor U863 (N_863,In_1548,In_2736);
xor U864 (N_864,In_3180,In_3263);
and U865 (N_865,In_804,In_3644);
and U866 (N_866,In_3003,In_4248);
or U867 (N_867,In_3653,In_1584);
xor U868 (N_868,In_1491,In_1399);
xor U869 (N_869,In_4552,In_1891);
nand U870 (N_870,In_903,In_1643);
and U871 (N_871,In_4637,In_3507);
nor U872 (N_872,In_2648,In_1381);
and U873 (N_873,In_716,In_450);
or U874 (N_874,In_3680,In_3444);
and U875 (N_875,In_2477,In_3519);
or U876 (N_876,In_3955,In_4648);
and U877 (N_877,In_1190,In_678);
or U878 (N_878,In_4390,In_4072);
xnor U879 (N_879,In_1610,In_4210);
and U880 (N_880,In_3910,In_2105);
or U881 (N_881,In_3198,In_709);
xnor U882 (N_882,In_4296,In_4022);
nand U883 (N_883,In_3513,In_1861);
xnor U884 (N_884,In_4077,In_3218);
and U885 (N_885,In_4438,In_4505);
nor U886 (N_886,In_101,In_1100);
or U887 (N_887,In_4055,In_2989);
and U888 (N_888,In_4948,In_472);
or U889 (N_889,In_226,In_1413);
nand U890 (N_890,In_424,In_706);
or U891 (N_891,In_1181,In_3612);
nand U892 (N_892,In_1211,In_4728);
nand U893 (N_893,In_2765,In_4942);
nor U894 (N_894,In_3591,In_2774);
or U895 (N_895,In_4064,In_1405);
and U896 (N_896,In_1388,In_199);
or U897 (N_897,In_661,In_4914);
and U898 (N_898,In_1527,In_4781);
nor U899 (N_899,In_1174,In_4177);
nor U900 (N_900,In_1831,In_2900);
and U901 (N_901,In_1221,In_1871);
xnor U902 (N_902,In_2643,In_4853);
or U903 (N_903,In_83,In_635);
and U904 (N_904,In_701,In_2570);
and U905 (N_905,In_186,In_1724);
or U906 (N_906,In_807,In_597);
xnor U907 (N_907,In_4046,In_117);
and U908 (N_908,In_1342,In_1457);
nand U909 (N_909,In_4074,In_1499);
xor U910 (N_910,In_4521,In_3153);
nand U911 (N_911,In_3329,In_116);
or U912 (N_912,In_456,In_4032);
nand U913 (N_913,In_3148,In_3970);
and U914 (N_914,In_2909,In_3004);
nand U915 (N_915,In_4417,In_502);
or U916 (N_916,In_133,In_4613);
and U917 (N_917,In_1495,In_3978);
and U918 (N_918,In_96,In_4855);
or U919 (N_919,In_4097,In_1789);
nor U920 (N_920,In_3391,In_2564);
nand U921 (N_921,In_3767,In_4540);
xor U922 (N_922,In_1547,In_3836);
and U923 (N_923,In_1461,In_2962);
nor U924 (N_924,In_4571,In_379);
or U925 (N_925,In_4366,In_2296);
xnor U926 (N_926,In_4079,In_1296);
and U927 (N_927,In_2798,In_1416);
nor U928 (N_928,In_4034,In_2346);
nand U929 (N_929,In_1837,In_1553);
xor U930 (N_930,In_4462,In_3980);
nor U931 (N_931,In_3862,In_2761);
and U932 (N_932,In_4973,In_2824);
nor U933 (N_933,In_4376,In_3544);
xor U934 (N_934,In_17,In_3778);
and U935 (N_935,In_380,In_309);
or U936 (N_936,In_2260,In_601);
nand U937 (N_937,In_783,In_2746);
and U938 (N_938,In_1385,In_122);
nor U939 (N_939,In_2360,In_4380);
nand U940 (N_940,In_118,In_3339);
or U941 (N_941,In_86,In_1300);
xor U942 (N_942,In_191,In_401);
nor U943 (N_943,In_4677,In_1205);
or U944 (N_944,In_4630,In_4963);
and U945 (N_945,In_76,In_4535);
or U946 (N_946,In_4795,In_3936);
nand U947 (N_947,In_4892,In_1956);
and U948 (N_948,In_3611,In_3666);
and U949 (N_949,In_2359,In_4670);
xnor U950 (N_950,In_1339,In_3546);
xnor U951 (N_951,In_1015,In_4713);
nand U952 (N_952,In_700,In_3404);
nor U953 (N_953,In_330,In_4378);
or U954 (N_954,In_2366,In_1439);
xor U955 (N_955,In_398,In_4170);
or U956 (N_956,In_4397,In_4373);
nor U957 (N_957,In_3408,In_1569);
xnor U958 (N_958,In_1626,In_994);
or U959 (N_959,In_3566,In_2055);
and U960 (N_960,In_4275,In_992);
or U961 (N_961,In_3025,In_3889);
nor U962 (N_962,In_1685,In_3154);
nand U963 (N_963,In_537,In_792);
xnor U964 (N_964,In_916,In_3174);
and U965 (N_965,In_1758,In_2695);
xnor U966 (N_966,In_1347,In_1189);
nor U967 (N_967,In_1717,In_3344);
nand U968 (N_968,In_3769,In_1583);
nand U969 (N_969,In_4634,In_3275);
and U970 (N_970,In_2795,In_3375);
and U971 (N_971,In_638,In_3053);
xor U972 (N_972,In_1255,In_4940);
nand U973 (N_973,In_2319,In_65);
or U974 (N_974,In_1052,In_4996);
xnor U975 (N_975,In_4491,In_2386);
nand U976 (N_976,In_991,In_1704);
xnor U977 (N_977,In_1108,In_3897);
nor U978 (N_978,In_2419,In_3343);
nor U979 (N_979,In_971,In_417);
and U980 (N_980,In_518,In_4954);
or U981 (N_981,In_285,In_4);
nand U982 (N_982,In_2197,In_3939);
and U983 (N_983,In_4169,In_167);
or U984 (N_984,In_2926,In_1515);
or U985 (N_985,In_4504,In_1018);
nand U986 (N_986,In_1761,In_3509);
or U987 (N_987,In_1455,In_2216);
xnor U988 (N_988,In_4107,In_4719);
xnor U989 (N_989,In_1382,In_1144);
or U990 (N_990,In_3642,In_4945);
nand U991 (N_991,In_1010,In_1698);
nand U992 (N_992,In_1152,In_1441);
xor U993 (N_993,In_3140,In_4645);
xnor U994 (N_994,In_2852,In_1091);
nand U995 (N_995,In_1842,In_584);
nor U996 (N_996,In_2231,In_4236);
nor U997 (N_997,In_4231,In_3524);
or U998 (N_998,In_3307,In_3065);
and U999 (N_999,In_4005,In_3748);
xnor U1000 (N_1000,In_3000,In_1887);
xor U1001 (N_1001,In_3533,In_3770);
nand U1002 (N_1002,In_2568,In_2590);
or U1003 (N_1003,In_359,In_3251);
nand U1004 (N_1004,In_1431,In_4171);
xnor U1005 (N_1005,In_3161,In_149);
nand U1006 (N_1006,In_4605,In_2491);
nor U1007 (N_1007,In_2139,In_2293);
or U1008 (N_1008,In_1746,In_2749);
and U1009 (N_1009,In_3531,In_2861);
or U1010 (N_1010,In_3672,In_4820);
xnor U1011 (N_1011,In_2083,In_3826);
and U1012 (N_1012,In_4759,In_1467);
nor U1013 (N_1013,In_4615,In_699);
and U1014 (N_1014,In_3379,In_784);
and U1015 (N_1015,In_2743,In_653);
and U1016 (N_1016,In_2860,In_2582);
nor U1017 (N_1017,In_2748,In_2814);
and U1018 (N_1018,In_4457,In_4512);
nor U1019 (N_1019,In_3473,In_1747);
and U1020 (N_1020,In_863,In_1130);
or U1021 (N_1021,In_2049,In_4026);
or U1022 (N_1022,In_3670,In_2351);
and U1023 (N_1023,In_1213,In_3760);
or U1024 (N_1024,In_655,In_2678);
xnor U1025 (N_1025,In_201,In_1148);
xor U1026 (N_1026,In_4499,In_2148);
nor U1027 (N_1027,In_2017,In_1344);
and U1028 (N_1028,In_632,In_891);
nand U1029 (N_1029,In_1575,In_3879);
nor U1030 (N_1030,In_2628,In_3909);
nor U1031 (N_1031,In_221,In_2222);
xor U1032 (N_1032,In_3056,In_780);
nor U1033 (N_1033,In_4359,In_2219);
and U1034 (N_1034,In_4843,In_4668);
or U1035 (N_1035,In_2306,In_1803);
xor U1036 (N_1036,In_619,In_2332);
xor U1037 (N_1037,In_4783,In_844);
nand U1038 (N_1038,In_2776,In_865);
nor U1039 (N_1039,In_3710,In_3870);
xnor U1040 (N_1040,In_2178,In_3588);
and U1041 (N_1041,In_160,In_2931);
nor U1042 (N_1042,In_114,In_3895);
xor U1043 (N_1043,In_1656,In_733);
nor U1044 (N_1044,In_2816,In_1318);
or U1045 (N_1045,In_4115,In_3608);
nand U1046 (N_1046,In_4823,In_2946);
and U1047 (N_1047,In_428,In_2585);
nand U1048 (N_1048,In_2558,In_4669);
nand U1049 (N_1049,In_1558,In_2317);
or U1050 (N_1050,In_2372,In_1963);
xnor U1051 (N_1051,In_3525,In_1988);
nor U1052 (N_1052,In_2484,In_3085);
and U1053 (N_1053,In_1365,In_1110);
xor U1054 (N_1054,In_2690,In_3119);
nand U1055 (N_1055,In_3502,In_1358);
or U1056 (N_1056,In_1090,In_2278);
xor U1057 (N_1057,In_2826,In_1721);
and U1058 (N_1058,In_3337,In_4742);
nand U1059 (N_1059,In_2714,In_872);
xor U1060 (N_1060,In_1184,In_1812);
or U1061 (N_1061,In_306,In_3692);
or U1062 (N_1062,In_4662,In_127);
nand U1063 (N_1063,In_2463,In_2971);
nor U1064 (N_1064,In_3324,In_3406);
and U1065 (N_1065,In_2228,In_688);
nor U1066 (N_1066,In_2445,In_4904);
and U1067 (N_1067,In_602,In_3459);
and U1068 (N_1068,In_3880,In_1474);
or U1069 (N_1069,In_4394,In_2427);
xnor U1070 (N_1070,In_1605,In_262);
nand U1071 (N_1071,In_304,In_3346);
xnor U1072 (N_1072,In_3234,In_955);
nand U1073 (N_1073,In_2660,In_4561);
nor U1074 (N_1074,In_3290,In_3947);
nand U1075 (N_1075,In_3797,In_3104);
nor U1076 (N_1076,In_3031,In_2067);
and U1077 (N_1077,In_3282,In_2637);
and U1078 (N_1078,In_4687,In_2880);
or U1079 (N_1079,In_3746,In_2392);
and U1080 (N_1080,In_3131,In_441);
nor U1081 (N_1081,In_2833,In_3291);
nor U1082 (N_1082,In_4844,In_3981);
xnor U1083 (N_1083,In_1479,In_7);
nand U1084 (N_1084,In_1476,In_851);
nor U1085 (N_1085,In_1287,In_2521);
nor U1086 (N_1086,In_1909,In_215);
and U1087 (N_1087,In_360,In_3232);
or U1088 (N_1088,In_4830,In_2843);
nor U1089 (N_1089,In_1723,In_675);
nand U1090 (N_1090,In_3506,In_3630);
nor U1091 (N_1091,In_1925,In_3446);
or U1092 (N_1092,In_940,In_763);
nand U1093 (N_1093,In_3483,In_809);
nand U1094 (N_1094,In_141,In_1002);
nand U1095 (N_1095,In_3024,In_451);
nand U1096 (N_1096,In_3697,In_4472);
nor U1097 (N_1097,In_4468,In_3452);
xnor U1098 (N_1098,In_1864,In_2285);
nor U1099 (N_1099,In_995,In_4633);
or U1100 (N_1100,In_185,In_4203);
or U1101 (N_1101,In_209,In_206);
nor U1102 (N_1102,In_4888,In_2547);
nand U1103 (N_1103,In_4225,In_3868);
nor U1104 (N_1104,In_4460,In_2778);
nand U1105 (N_1105,In_985,In_3202);
nand U1106 (N_1106,In_3592,In_2312);
or U1107 (N_1107,In_1768,In_350);
or U1108 (N_1108,In_3281,In_327);
xor U1109 (N_1109,In_2340,In_2614);
nor U1110 (N_1110,In_3305,In_795);
nor U1111 (N_1111,In_793,In_4625);
nor U1112 (N_1112,In_4983,In_3194);
nand U1113 (N_1113,In_3581,In_3859);
or U1114 (N_1114,In_1427,In_4158);
or U1115 (N_1115,In_3803,In_2264);
xnor U1116 (N_1116,In_1401,In_3819);
or U1117 (N_1117,In_1885,In_3562);
nand U1118 (N_1118,In_4651,In_2995);
nor U1119 (N_1119,In_835,In_729);
or U1120 (N_1120,In_3783,In_1981);
or U1121 (N_1121,In_1852,In_2759);
or U1122 (N_1122,In_1879,In_827);
nor U1123 (N_1123,In_3126,In_3301);
nor U1124 (N_1124,In_4114,In_3636);
nor U1125 (N_1125,In_4756,In_1106);
nand U1126 (N_1126,In_1203,In_2978);
xnor U1127 (N_1127,In_2310,In_1041);
or U1128 (N_1128,In_3877,In_3604);
nor U1129 (N_1129,In_1074,In_3614);
xor U1130 (N_1130,In_779,In_3433);
nor U1131 (N_1131,In_1714,In_4011);
and U1132 (N_1132,In_4873,In_583);
xor U1133 (N_1133,In_4172,In_4207);
xnor U1134 (N_1134,In_3839,In_2243);
nor U1135 (N_1135,In_4159,In_886);
and U1136 (N_1136,In_3241,In_4444);
nor U1137 (N_1137,In_3233,In_4184);
nand U1138 (N_1138,In_630,In_4640);
nand U1139 (N_1139,In_3185,In_3784);
nand U1140 (N_1140,In_4330,In_3904);
nand U1141 (N_1141,In_2711,In_918);
and U1142 (N_1142,In_950,In_4479);
or U1143 (N_1143,In_1733,In_1376);
xor U1144 (N_1144,In_2823,In_4514);
and U1145 (N_1145,In_2208,In_681);
xor U1146 (N_1146,In_423,In_2583);
and U1147 (N_1147,In_2122,In_1510);
nor U1148 (N_1148,In_3718,In_4737);
nor U1149 (N_1149,In_2990,In_2896);
and U1150 (N_1150,In_1514,In_1282);
nand U1151 (N_1151,In_1057,In_3299);
xor U1152 (N_1152,In_3958,In_546);
or U1153 (N_1153,In_1139,In_4833);
or U1154 (N_1154,In_1217,In_4985);
nor U1155 (N_1155,In_4804,In_922);
nor U1156 (N_1156,In_4682,In_2406);
nand U1157 (N_1157,In_2314,In_1225);
nand U1158 (N_1158,In_2196,In_334);
xnor U1159 (N_1159,In_4425,In_1301);
nor U1160 (N_1160,In_462,In_1813);
and U1161 (N_1161,In_4553,In_3683);
and U1162 (N_1162,In_2914,In_1604);
nand U1163 (N_1163,In_907,In_99);
xnor U1164 (N_1164,In_867,In_956);
nor U1165 (N_1165,In_170,In_2468);
and U1166 (N_1166,In_4478,In_1900);
nand U1167 (N_1167,In_4907,In_2223);
nand U1168 (N_1168,In_3726,In_3974);
nand U1169 (N_1169,In_1244,In_455);
and U1170 (N_1170,In_2725,In_738);
xnor U1171 (N_1171,In_4323,In_1126);
nand U1172 (N_1172,In_2035,In_2671);
nor U1173 (N_1173,In_2526,In_2742);
or U1174 (N_1174,In_4883,In_1129);
nand U1175 (N_1175,In_2474,In_3092);
nand U1176 (N_1176,In_2653,In_4789);
nor U1177 (N_1177,In_698,In_136);
and U1178 (N_1178,In_1580,In_4387);
nand U1179 (N_1179,In_4760,In_3138);
xnor U1180 (N_1180,In_4777,In_1407);
nor U1181 (N_1181,In_484,In_126);
xnor U1182 (N_1182,In_3739,In_626);
nand U1183 (N_1183,In_1092,In_3641);
and U1184 (N_1184,In_2872,In_1128);
nor U1185 (N_1185,In_3550,In_2943);
xnor U1186 (N_1186,In_2272,In_3231);
or U1187 (N_1187,In_2098,In_3292);
nor U1188 (N_1188,In_3829,In_926);
or U1189 (N_1189,In_2524,In_3400);
nor U1190 (N_1190,In_3685,In_728);
or U1191 (N_1191,In_4578,In_4386);
or U1192 (N_1192,In_4986,In_48);
nand U1193 (N_1193,In_3388,In_4780);
or U1194 (N_1194,In_3143,In_3051);
nand U1195 (N_1195,In_3943,In_1146);
nand U1196 (N_1196,In_986,In_193);
nor U1197 (N_1197,In_3929,In_828);
or U1198 (N_1198,In_3569,In_727);
and U1199 (N_1199,In_4234,In_4792);
and U1200 (N_1200,In_1028,In_4688);
nand U1201 (N_1201,In_3969,In_2694);
nand U1202 (N_1202,In_240,In_1720);
nand U1203 (N_1203,In_4277,In_3841);
or U1204 (N_1204,In_4934,In_1519);
xor U1205 (N_1205,In_2050,In_2609);
xnor U1206 (N_1206,In_4398,In_2925);
nor U1207 (N_1207,In_2810,In_4232);
nor U1208 (N_1208,In_1497,In_1425);
nand U1209 (N_1209,In_4066,In_3099);
xor U1210 (N_1210,In_1641,In_4301);
nor U1211 (N_1211,In_4848,In_159);
or U1212 (N_1212,In_786,In_2902);
nor U1213 (N_1213,In_3686,In_4994);
xnor U1214 (N_1214,In_2404,In_3931);
and U1215 (N_1215,In_111,In_4920);
or U1216 (N_1216,In_3582,In_4303);
nand U1217 (N_1217,In_2420,In_536);
nor U1218 (N_1218,In_3010,In_1996);
or U1219 (N_1219,In_318,In_477);
and U1220 (N_1220,In_2717,In_4588);
xnor U1221 (N_1221,In_938,In_3413);
nand U1222 (N_1222,In_1432,In_3098);
nor U1223 (N_1223,In_4717,In_4748);
xor U1224 (N_1224,In_2000,In_4361);
or U1225 (N_1225,In_4448,In_612);
nand U1226 (N_1226,In_2610,In_4691);
xor U1227 (N_1227,In_2542,In_3954);
and U1228 (N_1228,In_3935,In_967);
nor U1229 (N_1229,In_1173,In_3528);
and U1230 (N_1230,In_2696,In_387);
nand U1231 (N_1231,In_4746,In_3849);
nand U1232 (N_1232,In_1919,In_4689);
or U1233 (N_1233,In_2741,In_4201);
nor U1234 (N_1234,In_123,In_1175);
and U1235 (N_1235,In_317,In_2322);
nor U1236 (N_1236,In_2947,In_2053);
xor U1237 (N_1237,In_1241,In_693);
and U1238 (N_1238,In_4187,In_4539);
nand U1239 (N_1239,In_4299,In_2605);
nand U1240 (N_1240,In_2184,In_1675);
nor U1241 (N_1241,In_4638,In_4911);
or U1242 (N_1242,In_667,In_2258);
nor U1243 (N_1243,In_1779,In_356);
and U1244 (N_1244,In_4592,In_37);
nor U1245 (N_1245,In_4041,In_2500);
nor U1246 (N_1246,In_4204,In_3994);
nand U1247 (N_1247,In_414,In_888);
or U1248 (N_1248,In_4968,In_1026);
and U1249 (N_1249,In_4741,In_4260);
and U1250 (N_1250,In_3790,In_2700);
nand U1251 (N_1251,In_2263,In_3453);
nor U1252 (N_1252,In_2466,In_3227);
and U1253 (N_1253,In_1123,In_1824);
and U1254 (N_1254,In_2109,In_2911);
nor U1255 (N_1255,In_3371,In_4268);
nor U1256 (N_1256,In_3449,In_26);
nand U1257 (N_1257,In_492,In_4595);
or U1258 (N_1258,In_1689,In_4621);
and U1259 (N_1259,In_1071,In_1534);
nor U1260 (N_1260,In_2959,In_3208);
or U1261 (N_1261,In_965,In_3828);
xor U1262 (N_1262,In_656,In_3374);
nand U1263 (N_1263,In_2431,In_464);
xor U1264 (N_1264,In_1906,In_4218);
and U1265 (N_1265,In_4698,In_4071);
xor U1266 (N_1266,In_657,In_4082);
or U1267 (N_1267,In_1315,In_3086);
or U1268 (N_1268,In_1585,In_4680);
or U1269 (N_1269,In_3679,In_4364);
and U1270 (N_1270,In_1334,In_4683);
and U1271 (N_1271,In_1172,In_3957);
and U1272 (N_1272,In_3246,In_93);
nand U1273 (N_1273,In_4150,In_2619);
xnor U1274 (N_1274,In_2462,In_1991);
nor U1275 (N_1275,In_2827,In_239);
nand U1276 (N_1276,In_1132,In_1277);
or U1277 (N_1277,In_3149,In_1930);
or U1278 (N_1278,In_2664,In_945);
or U1279 (N_1279,In_3801,In_1960);
or U1280 (N_1280,In_3621,In_3684);
nand U1281 (N_1281,In_798,In_532);
nor U1282 (N_1282,In_2809,In_471);
or U1283 (N_1283,In_1718,In_1201);
xnor U1284 (N_1284,In_4428,In_1973);
xnor U1285 (N_1285,In_4108,In_900);
nand U1286 (N_1286,In_3993,In_4518);
xor U1287 (N_1287,In_1395,In_1833);
and U1288 (N_1288,In_1209,In_2087);
xnor U1289 (N_1289,In_3352,In_1324);
or U1290 (N_1290,In_3157,In_1493);
and U1291 (N_1291,In_2189,In_4370);
xor U1292 (N_1292,In_4714,In_3248);
nor U1293 (N_1293,In_997,In_958);
nand U1294 (N_1294,In_1485,In_920);
nand U1295 (N_1295,In_2151,In_4389);
xor U1296 (N_1296,In_2571,In_3039);
nand U1297 (N_1297,In_1857,In_2716);
or U1298 (N_1298,In_3225,In_452);
xor U1299 (N_1299,In_3776,In_1019);
and U1300 (N_1300,In_4445,In_3358);
xor U1301 (N_1301,In_2898,In_595);
nand U1302 (N_1302,In_2074,In_4382);
nor U1303 (N_1303,In_3711,In_1791);
or U1304 (N_1304,In_3918,In_392);
nor U1305 (N_1305,In_375,In_3109);
nand U1306 (N_1306,In_1942,In_3806);
nand U1307 (N_1307,In_293,In_3724);
xor U1308 (N_1308,In_426,In_213);
nand U1309 (N_1309,In_20,In_2465);
and U1310 (N_1310,In_4915,In_1478);
nor U1311 (N_1311,In_2822,In_3076);
nor U1312 (N_1312,In_1185,In_989);
or U1313 (N_1313,In_2302,In_1692);
and U1314 (N_1314,In_3166,In_3706);
xor U1315 (N_1315,In_591,In_1961);
xnor U1316 (N_1316,In_1749,In_2498);
nand U1317 (N_1317,In_1169,In_1350);
nand U1318 (N_1318,In_188,In_568);
and U1319 (N_1319,In_4035,In_3816);
nand U1320 (N_1320,In_826,In_32);
xnor U1321 (N_1321,In_4574,In_3728);
nand U1322 (N_1322,In_3512,In_893);
and U1323 (N_1323,In_2096,In_1663);
and U1324 (N_1324,In_911,In_2038);
nand U1325 (N_1325,In_2238,In_444);
nor U1326 (N_1326,In_2649,In_3917);
and U1327 (N_1327,In_866,In_4109);
and U1328 (N_1328,In_2543,In_4729);
nand U1329 (N_1329,In_3402,In_1363);
and U1330 (N_1330,In_4982,In_3818);
xor U1331 (N_1331,In_3733,In_4264);
xor U1332 (N_1332,In_3671,In_3478);
xor U1333 (N_1333,In_553,In_4739);
and U1334 (N_1334,In_4502,In_4144);
or U1335 (N_1335,In_740,In_503);
or U1336 (N_1336,In_4559,In_4339);
nor U1337 (N_1337,In_3303,In_1483);
or U1338 (N_1338,In_3037,In_4684);
nor U1339 (N_1339,In_1504,In_195);
and U1340 (N_1340,In_4627,In_1631);
nand U1341 (N_1341,In_1577,In_4943);
nor U1342 (N_1342,In_3102,In_2599);
nand U1343 (N_1343,In_300,In_4135);
nor U1344 (N_1344,In_2449,In_2638);
xor U1345 (N_1345,In_1389,In_864);
xnor U1346 (N_1346,In_2015,In_383);
nand U1347 (N_1347,In_921,In_1551);
nand U1348 (N_1348,In_2315,In_4533);
nand U1349 (N_1349,In_3244,In_734);
xor U1350 (N_1350,In_4944,In_2483);
and U1351 (N_1351,In_1337,In_3399);
nor U1352 (N_1352,In_1735,In_2684);
or U1353 (N_1353,In_3752,In_2578);
nor U1354 (N_1354,In_2124,In_1695);
nor U1355 (N_1355,In_3249,In_1888);
nand U1356 (N_1356,In_3944,In_1754);
nor U1357 (N_1357,In_3786,In_4421);
nand U1358 (N_1358,In_337,In_4127);
xor U1359 (N_1359,In_4928,In_4315);
xor U1360 (N_1360,In_109,In_4837);
or U1361 (N_1361,In_1023,In_4750);
nor U1362 (N_1362,In_1855,In_2829);
and U1363 (N_1363,In_3650,In_3999);
nor U1364 (N_1364,In_4766,In_432);
or U1365 (N_1365,In_1017,In_1299);
nor U1366 (N_1366,In_4956,In_1197);
nand U1367 (N_1367,In_2295,In_982);
or U1368 (N_1368,In_1587,In_3508);
nor U1369 (N_1369,In_463,In_3317);
nand U1370 (N_1370,In_2905,In_1272);
and U1371 (N_1371,In_1191,In_990);
xnor U1372 (N_1372,In_999,In_349);
nand U1373 (N_1373,In_2214,In_385);
and U1374 (N_1374,In_4939,In_4436);
nor U1375 (N_1375,In_500,In_4723);
nand U1376 (N_1376,In_399,In_3381);
nand U1377 (N_1377,In_1752,In_3224);
and U1378 (N_1378,In_4429,In_2533);
xnor U1379 (N_1379,In_4080,In_2195);
or U1380 (N_1380,In_4403,In_1032);
xor U1381 (N_1381,In_556,In_1679);
and U1382 (N_1382,In_2520,In_840);
or U1383 (N_1383,In_1722,In_3277);
and U1384 (N_1384,In_3066,In_3888);
xor U1385 (N_1385,In_1494,In_250);
nor U1386 (N_1386,In_61,In_3758);
nor U1387 (N_1387,In_1638,In_4829);
and U1388 (N_1388,In_4310,In_2871);
nor U1389 (N_1389,In_2781,In_4721);
nor U1390 (N_1390,In_2169,In_4224);
nor U1391 (N_1391,In_62,In_3289);
xor U1392 (N_1392,In_842,In_168);
and U1393 (N_1393,In_913,In_2052);
or U1394 (N_1394,In_3034,In_2072);
nand U1395 (N_1395,In_4644,In_564);
xnor U1396 (N_1396,In_4329,In_3011);
nand U1397 (N_1397,In_4014,In_1422);
or U1398 (N_1398,In_148,In_66);
nor U1399 (N_1399,In_2405,In_2046);
nand U1400 (N_1400,In_4528,In_2464);
or U1401 (N_1401,In_498,In_3043);
nor U1402 (N_1402,In_2532,In_407);
xor U1403 (N_1403,In_1035,In_46);
or U1404 (N_1404,In_1187,In_3228);
and U1405 (N_1405,In_403,In_665);
and U1406 (N_1406,In_3468,In_2552);
xor U1407 (N_1407,In_256,In_4168);
and U1408 (N_1408,In_1821,In_1597);
or U1409 (N_1409,In_3798,In_3615);
nand U1410 (N_1410,In_1238,In_1072);
or U1411 (N_1411,In_1068,In_2063);
nor U1412 (N_1412,In_2732,In_4765);
or U1413 (N_1413,In_4799,In_2659);
and U1414 (N_1414,In_2886,In_4313);
and U1415 (N_1415,In_3476,In_1639);
xnor U1416 (N_1416,In_4200,In_1246);
or U1417 (N_1417,In_2728,In_4197);
and U1418 (N_1418,In_2981,In_2802);
nor U1419 (N_1419,In_993,In_4734);
or U1420 (N_1420,In_1056,In_421);
and U1421 (N_1421,In_4254,In_3754);
and U1422 (N_1422,In_4851,In_558);
nand U1423 (N_1423,In_1430,In_2472);
nor U1424 (N_1424,In_628,In_3660);
xnor U1425 (N_1425,In_853,In_4045);
or U1426 (N_1426,In_2887,In_4581);
or U1427 (N_1427,In_810,In_2594);
and U1428 (N_1428,In_1261,In_1966);
nor U1429 (N_1429,In_4492,In_10);
xor U1430 (N_1430,In_1135,In_51);
or U1431 (N_1431,In_402,In_3921);
nand U1432 (N_1432,In_2567,In_3924);
nor U1433 (N_1433,In_2138,In_1907);
or U1434 (N_1434,In_762,In_590);
nor U1435 (N_1435,In_1523,In_447);
nor U1436 (N_1436,In_2988,In_4388);
or U1437 (N_1437,In_2007,In_2324);
or U1438 (N_1438,In_2630,In_3210);
nand U1439 (N_1439,In_1902,In_2523);
and U1440 (N_1440,In_3293,In_1193);
and U1441 (N_1441,In_254,In_1989);
or U1442 (N_1442,In_4112,In_3023);
xor U1443 (N_1443,In_1549,In_3443);
nand U1444 (N_1444,In_1464,In_4318);
xnor U1445 (N_1445,In_4706,In_1099);
nor U1446 (N_1446,In_3330,In_833);
xnor U1447 (N_1447,In_341,In_3736);
xnor U1448 (N_1448,In_2661,In_3312);
nand U1449 (N_1449,In_3847,In_1992);
and U1450 (N_1450,In_4524,In_1199);
and U1451 (N_1451,In_3038,In_2954);
and U1452 (N_1452,In_673,In_1359);
and U1453 (N_1453,In_2882,In_1731);
and U1454 (N_1454,In_2801,In_4038);
or U1455 (N_1455,In_1788,In_483);
nor U1456 (N_1456,In_3585,In_1482);
nand U1457 (N_1457,In_3331,In_4998);
nor U1458 (N_1458,In_2787,In_1650);
or U1459 (N_1459,In_4544,In_2034);
or U1460 (N_1460,In_824,In_3078);
xor U1461 (N_1461,In_4984,In_1828);
or U1462 (N_1462,In_4110,In_2283);
or U1463 (N_1463,In_592,In_825);
xnor U1464 (N_1464,In_439,In_2135);
nand U1465 (N_1465,In_3744,In_3142);
or U1466 (N_1466,In_2808,In_1210);
nor U1467 (N_1467,In_4325,In_162);
and U1468 (N_1468,In_4358,In_110);
nor U1469 (N_1469,In_4821,In_2731);
or U1470 (N_1470,In_3737,In_767);
nand U1471 (N_1471,In_4772,In_560);
or U1472 (N_1472,In_4242,In_56);
nand U1473 (N_1473,In_660,In_1038);
xor U1474 (N_1474,In_3073,In_3130);
xor U1475 (N_1475,In_3695,In_1559);
xnor U1476 (N_1476,In_59,In_386);
or U1477 (N_1477,In_4027,In_2663);
xnor U1478 (N_1478,In_1316,In_4151);
nor U1479 (N_1479,In_753,In_3802);
xnor U1480 (N_1480,In_3437,In_1331);
or U1481 (N_1481,In_1031,In_4647);
and U1482 (N_1482,In_4622,In_64);
xnor U1483 (N_1483,In_2397,In_4560);
nand U1484 (N_1484,In_1702,In_2994);
nand U1485 (N_1485,In_3500,In_2701);
nand U1486 (N_1486,In_2171,In_3440);
nand U1487 (N_1487,In_87,In_3019);
nor U1488 (N_1488,In_1868,In_2908);
nor U1489 (N_1489,In_904,In_1306);
xnor U1490 (N_1490,In_2718,In_211);
xnor U1491 (N_1491,In_3631,In_2985);
xor U1492 (N_1492,In_4642,In_3489);
or U1493 (N_1493,In_4850,In_1596);
and U1494 (N_1494,In_4247,In_2968);
nor U1495 (N_1495,In_2707,In_4320);
nand U1496 (N_1496,In_1501,In_2079);
nand U1497 (N_1497,In_2304,In_4048);
nor U1498 (N_1498,In_4912,In_4165);
nor U1499 (N_1499,In_1876,In_3151);
or U1500 (N_1500,In_2280,In_4654);
or U1501 (N_1501,In_4715,In_203);
xnor U1502 (N_1502,In_3652,In_2030);
nand U1503 (N_1503,In_3964,In_4160);
and U1504 (N_1504,In_2145,In_852);
or U1505 (N_1505,In_2005,In_180);
nor U1506 (N_1506,In_639,In_915);
xor U1507 (N_1507,In_3866,In_942);
and U1508 (N_1508,In_998,In_2176);
nor U1509 (N_1509,In_33,In_4700);
xnor U1510 (N_1510,In_4185,In_2735);
xor U1511 (N_1511,In_4810,In_4531);
xnor U1512 (N_1512,In_3827,In_3985);
nor U1513 (N_1513,In_506,In_857);
xnor U1514 (N_1514,In_4147,In_4489);
and U1515 (N_1515,In_302,In_4180);
nor U1516 (N_1516,In_92,In_1488);
or U1517 (N_1517,In_4897,In_1694);
xnor U1518 (N_1518,In_2001,In_3392);
nor U1519 (N_1519,In_3272,In_2680);
xnor U1520 (N_1520,In_4161,In_275);
nand U1521 (N_1521,In_4643,In_2391);
xor U1522 (N_1522,In_4456,In_4923);
and U1523 (N_1523,In_2763,In_949);
or U1524 (N_1524,In_2437,In_3656);
nand U1525 (N_1525,In_1967,In_1729);
nor U1526 (N_1526,In_2027,In_607);
nand U1527 (N_1527,In_3222,In_3623);
nor U1528 (N_1528,In_3905,In_2530);
xnor U1529 (N_1529,In_4526,In_3494);
nor U1530 (N_1530,In_2354,In_2207);
nand U1531 (N_1531,In_476,In_1932);
or U1532 (N_1532,In_4399,In_2282);
or U1533 (N_1533,In_4847,In_2018);
and U1534 (N_1534,In_1520,In_2756);
nor U1535 (N_1535,In_1075,In_214);
or U1536 (N_1536,In_1268,In_135);
nor U1537 (N_1537,In_3276,In_3702);
or U1538 (N_1538,In_3529,In_4418);
xor U1539 (N_1539,In_220,In_2897);
and U1540 (N_1540,In_2750,In_1014);
and U1541 (N_1541,In_2358,In_1516);
nor U1542 (N_1542,In_4964,In_4880);
and U1543 (N_1543,In_2513,In_2210);
nand U1544 (N_1544,In_80,In_3230);
nand U1545 (N_1545,In_3316,In_1459);
nor U1546 (N_1546,In_4396,In_4228);
and U1547 (N_1547,In_4148,In_742);
or U1548 (N_1548,In_2104,In_4761);
nor U1549 (N_1549,In_1333,In_3952);
nand U1550 (N_1550,In_4047,In_1089);
nand U1551 (N_1551,In_4860,In_910);
nand U1552 (N_1552,In_1668,In_2686);
nor U1553 (N_1553,In_3678,In_2720);
xnor U1554 (N_1554,In_3411,In_1603);
xor U1555 (N_1555,In_2881,In_4476);
xor U1556 (N_1556,In_2691,In_4439);
nor U1557 (N_1557,In_720,In_547);
or U1558 (N_1558,In_1458,In_4422);
or U1559 (N_1559,In_2137,In_3908);
xor U1560 (N_1560,In_3096,In_322);
or U1561 (N_1561,In_4730,In_173);
nor U1562 (N_1562,In_1725,In_3150);
xor U1563 (N_1563,In_2160,In_898);
xor U1564 (N_1564,In_4295,In_187);
xor U1565 (N_1565,In_1336,In_4635);
and U1566 (N_1566,In_316,In_3093);
nor U1567 (N_1567,In_515,In_539);
xnor U1568 (N_1568,In_3648,In_3067);
xnor U1569 (N_1569,In_164,In_4118);
and U1570 (N_1570,In_4293,In_4814);
xor U1571 (N_1571,In_1521,In_4674);
nor U1572 (N_1572,In_4902,In_4856);
nand U1573 (N_1573,In_1806,In_875);
or U1574 (N_1574,In_4314,In_2937);
xor U1575 (N_1575,In_3405,In_3310);
xnor U1576 (N_1576,In_2254,In_4655);
nor U1577 (N_1577,In_4577,In_481);
xor U1578 (N_1578,In_2734,In_2286);
nand U1579 (N_1579,In_1600,In_4890);
nor U1580 (N_1580,In_3723,In_3609);
and U1581 (N_1581,In_4276,In_2961);
nand U1582 (N_1582,In_2443,In_3288);
and U1583 (N_1583,In_2215,In_2233);
nor U1584 (N_1584,In_1465,In_3070);
or U1585 (N_1585,In_2118,In_3103);
or U1586 (N_1586,In_4343,In_1517);
or U1587 (N_1587,In_1345,In_2337);
xor U1588 (N_1588,In_4620,In_2864);
xor U1589 (N_1589,In_4791,In_1943);
xnor U1590 (N_1590,In_776,In_3255);
or U1591 (N_1591,In_3795,In_620);
nand U1592 (N_1592,In_2495,In_2595);
nand U1593 (N_1593,In_4321,In_1276);
and U1594 (N_1594,In_2183,In_1727);
nand U1595 (N_1595,In_1543,In_2275);
xor U1596 (N_1596,In_2458,In_3953);
and U1597 (N_1597,In_3059,In_687);
xor U1598 (N_1598,In_3645,In_2094);
and U1599 (N_1599,In_2751,In_1946);
and U1600 (N_1600,In_1574,In_4564);
nand U1601 (N_1601,In_4819,In_2804);
nand U1602 (N_1602,In_4051,In_3771);
nand U1603 (N_1603,In_1826,In_1219);
nor U1604 (N_1604,In_308,In_4554);
or U1605 (N_1605,In_3116,In_1000);
or U1606 (N_1606,In_636,In_2201);
or U1607 (N_1607,In_3975,In_1487);
xor U1608 (N_1608,In_6,In_30);
xnor U1609 (N_1609,In_2837,In_1220);
and U1610 (N_1610,In_333,In_1867);
xor U1611 (N_1611,In_1982,In_2290);
xor U1612 (N_1612,In_1530,In_144);
and U1613 (N_1613,In_1608,In_1635);
or U1614 (N_1614,In_4117,In_2666);
and U1615 (N_1615,In_2940,In_3832);
and U1616 (N_1616,In_435,In_3545);
and U1617 (N_1617,In_75,In_1745);
xor U1618 (N_1618,In_1446,In_4614);
nor U1619 (N_1619,In_1086,In_3430);
nor U1620 (N_1620,In_4141,In_3111);
nor U1621 (N_1621,In_3356,In_3088);
or U1622 (N_1622,In_1544,In_3534);
nor U1623 (N_1623,In_2855,In_4971);
xor U1624 (N_1624,In_1759,In_2836);
xnor U1625 (N_1625,In_2246,In_4966);
and U1626 (N_1626,In_344,In_2517);
xor U1627 (N_1627,In_3155,In_748);
or U1628 (N_1628,In_2165,In_2770);
or U1629 (N_1629,In_1312,In_2561);
xor U1630 (N_1630,In_2569,In_3229);
or U1631 (N_1631,In_4302,In_3720);
and U1632 (N_1632,In_805,In_2555);
xor U1633 (N_1633,In_3527,In_2821);
and U1634 (N_1634,In_3996,In_2790);
xor U1635 (N_1635,In_2657,In_124);
nand U1636 (N_1636,In_1060,In_3054);
xnor U1637 (N_1637,In_4899,In_4872);
or U1638 (N_1638,In_4757,In_4508);
or U1639 (N_1639,In_2229,In_3600);
xor U1640 (N_1640,In_895,In_2042);
nand U1641 (N_1641,In_2345,In_3445);
nand U1642 (N_1642,In_2421,In_3442);
xor U1643 (N_1643,In_627,In_2755);
nand U1644 (N_1644,In_1153,In_4427);
xnor U1645 (N_1645,In_2450,In_140);
xor U1646 (N_1646,In_3283,In_265);
or U1647 (N_1647,In_3193,In_4075);
nor U1648 (N_1648,In_69,In_77);
or U1649 (N_1649,In_2689,In_2807);
nand U1650 (N_1650,In_3725,In_1364);
nor U1651 (N_1651,In_2459,In_1121);
and U1652 (N_1652,In_4937,In_3401);
and U1653 (N_1653,In_2117,In_501);
or U1654 (N_1654,In_3570,In_4903);
nand U1655 (N_1655,In_2854,In_4012);
xor U1656 (N_1656,In_1985,In_3382);
nand U1657 (N_1657,In_1192,In_4273);
nand U1658 (N_1658,In_1270,In_4879);
nor U1659 (N_1659,In_1904,In_4590);
nor U1660 (N_1660,In_2982,In_1136);
nand U1661 (N_1661,In_1408,In_3504);
nand U1662 (N_1662,In_2644,In_889);
nor U1663 (N_1663,In_3325,In_276);
and U1664 (N_1664,In_834,In_1143);
nor U1665 (N_1665,In_2446,In_2221);
nor U1666 (N_1666,In_3261,In_25);
and U1667 (N_1667,In_2327,In_3466);
nor U1668 (N_1668,In_2395,In_3355);
or U1669 (N_1669,In_2436,In_769);
nor U1670 (N_1670,In_2175,In_771);
and U1671 (N_1671,In_765,In_2579);
or U1672 (N_1672,In_4527,In_1818);
xnor U1673 (N_1673,In_2779,In_2116);
xor U1674 (N_1674,In_2131,In_3699);
nand U1675 (N_1675,In_671,In_2739);
and U1676 (N_1676,In_4096,In_2273);
nand U1677 (N_1677,In_4898,In_1212);
nand U1678 (N_1678,In_3796,In_1053);
and U1679 (N_1679,In_4787,In_1371);
and U1680 (N_1680,In_4363,In_3824);
xnor U1681 (N_1681,In_88,In_4298);
xor U1682 (N_1682,In_1687,In_12);
and U1683 (N_1683,In_758,In_438);
nand U1684 (N_1684,In_4265,In_4414);
nand U1685 (N_1685,In_1375,In_3934);
nor U1686 (N_1686,In_668,In_440);
nand U1687 (N_1687,In_3950,In_2602);
or U1688 (N_1688,In_2573,In_372);
and U1689 (N_1689,In_115,In_4901);
and U1690 (N_1690,In_2244,In_139);
nand U1691 (N_1691,In_836,In_524);
nand U1692 (N_1692,In_4816,In_2064);
and U1693 (N_1693,In_1865,In_2125);
xnor U1694 (N_1694,In_2627,In_2365);
and U1695 (N_1695,In_2388,In_4281);
xor U1696 (N_1696,In_2177,In_3265);
nor U1697 (N_1697,In_1262,In_2879);
xor U1698 (N_1698,In_1845,In_2862);
or U1699 (N_1699,In_4534,In_4589);
nor U1700 (N_1700,In_1915,In_2764);
and U1701 (N_1701,In_1908,In_2740);
xnor U1702 (N_1702,In_2261,In_3542);
nand U1703 (N_1703,In_436,In_3628);
or U1704 (N_1704,In_2683,In_1987);
or U1705 (N_1705,In_1999,In_4582);
and U1706 (N_1706,In_1662,In_549);
and U1707 (N_1707,In_4743,In_3713);
and U1708 (N_1708,In_2762,In_4490);
xnor U1709 (N_1709,In_1945,In_2307);
and U1710 (N_1710,In_3912,In_3243);
nor U1711 (N_1711,In_323,In_1645);
and U1712 (N_1712,In_3327,In_957);
nor U1713 (N_1713,In_4190,In_3367);
xnor U1714 (N_1714,In_2539,In_2335);
nand U1715 (N_1715,In_1116,In_2270);
and U1716 (N_1716,In_364,In_4312);
xor U1717 (N_1717,In_2328,In_2586);
or U1718 (N_1718,In_1618,In_1628);
nor U1719 (N_1719,In_686,In_1383);
xnor U1720 (N_1720,In_4832,In_2162);
and U1721 (N_1721,In_3238,In_4495);
nor U1722 (N_1722,In_2708,In_274);
or U1723 (N_1723,In_3106,In_1793);
xor U1724 (N_1724,In_4375,In_4599);
or U1725 (N_1725,In_3128,In_3719);
xnor U1726 (N_1726,In_4309,In_491);
nor U1727 (N_1727,In_527,In_3178);
and U1728 (N_1728,In_2834,In_1750);
xor U1729 (N_1729,In_3127,In_248);
nor U1730 (N_1730,In_4416,In_816);
and U1731 (N_1731,In_3206,In_4591);
xor U1732 (N_1732,In_2256,In_4754);
or U1733 (N_1733,In_2999,In_1936);
xor U1734 (N_1734,In_4861,In_676);
xor U1735 (N_1735,In_2496,In_1284);
nand U1736 (N_1736,In_4352,In_490);
nor U1737 (N_1737,In_4092,In_2037);
nand U1738 (N_1738,In_4600,In_178);
or U1739 (N_1739,In_2432,In_3520);
nor U1740 (N_1740,In_2505,In_2374);
or U1741 (N_1741,In_343,In_2753);
and U1742 (N_1742,In_4846,In_4300);
and U1743 (N_1743,In_3447,In_4332);
and U1744 (N_1744,In_4434,In_3759);
nor U1745 (N_1745,In_321,In_3823);
or U1746 (N_1746,In_684,In_3160);
or U1747 (N_1747,In_3629,In_1781);
or U1748 (N_1748,In_2190,In_2194);
or U1749 (N_1749,In_1460,In_2991);
nor U1750 (N_1750,In_819,In_917);
xor U1751 (N_1751,In_458,In_4917);
or U1752 (N_1752,In_3319,In_1678);
nand U1753 (N_1753,In_760,In_1037);
xor U1754 (N_1754,In_1236,In_3209);
nor U1755 (N_1755,In_3080,In_1814);
and U1756 (N_1756,In_454,In_5);
nand U1757 (N_1757,In_1374,In_2675);
nand U1758 (N_1758,In_4324,In_1016);
and U1759 (N_1759,In_2929,In_919);
nand U1760 (N_1760,In_4672,In_4337);
nand U1761 (N_1761,In_751,In_739);
xor U1762 (N_1762,In_4991,In_2476);
xor U1763 (N_1763,In_2912,In_1113);
nor U1764 (N_1764,In_643,In_3100);
xnor U1765 (N_1765,In_4368,In_981);
or U1766 (N_1766,In_554,In_2134);
or U1767 (N_1767,In_3640,In_552);
xor U1768 (N_1768,In_208,In_2133);
nor U1769 (N_1769,In_3287,In_1249);
or U1770 (N_1770,In_526,In_1188);
or U1771 (N_1771,In_4974,In_4580);
nand U1772 (N_1772,In_3556,In_4735);
nor U1773 (N_1773,In_2003,In_1538);
and U1774 (N_1774,In_1330,In_4636);
xor U1775 (N_1775,In_3755,In_980);
nand U1776 (N_1776,In_3674,In_4793);
or U1777 (N_1777,In_4250,In_3812);
nor U1778 (N_1778,In_2172,In_3890);
nand U1779 (N_1779,In_4612,In_4835);
xnor U1780 (N_1780,In_1726,In_1565);
nor U1781 (N_1781,In_1854,In_1378);
xnor U1782 (N_1782,In_224,In_4284);
nand U1783 (N_1783,In_2752,In_542);
nor U1784 (N_1784,In_4068,In_2723);
nand U1785 (N_1785,In_3475,In_1690);
xor U1786 (N_1786,In_3705,In_1682);
nor U1787 (N_1787,In_4289,In_1426);
nor U1788 (N_1788,In_277,In_1328);
xor U1789 (N_1789,In_1666,In_2394);
or U1790 (N_1790,In_3333,In_2979);
xnor U1791 (N_1791,In_1463,In_1036);
nor U1792 (N_1792,In_2305,In_3013);
nand U1793 (N_1793,In_743,In_1541);
nor U1794 (N_1794,In_3643,In_1952);
or U1795 (N_1795,In_4549,In_1420);
nor U1796 (N_1796,In_3837,In_757);
or U1797 (N_1797,In_766,In_232);
or U1798 (N_1798,In_4485,In_1417);
and U1799 (N_1799,In_1085,In_82);
xor U1800 (N_1800,In_4052,In_2110);
nor U1801 (N_1801,In_4007,In_2218);
and U1802 (N_1802,In_4802,In_3940);
xor U1803 (N_1803,In_1279,In_2915);
or U1804 (N_1804,In_4726,In_3854);
nor U1805 (N_1805,In_3429,In_4056);
xor U1806 (N_1806,In_947,In_1352);
or U1807 (N_1807,In_4304,In_1046);
nor U1808 (N_1808,In_3772,In_4586);
nor U1809 (N_1809,In_1020,In_772);
or U1810 (N_1810,In_2966,In_4059);
or U1811 (N_1811,In_3766,In_442);
nand U1812 (N_1812,In_1372,In_3490);
or U1813 (N_1813,In_2705,In_692);
nor U1814 (N_1814,In_2729,In_658);
xor U1815 (N_1815,In_3474,In_2029);
or U1816 (N_1816,In_1934,In_541);
nor U1817 (N_1817,In_754,In_3028);
nand U1818 (N_1818,In_4955,In_3938);
xor U1819 (N_1819,In_3014,In_4162);
nand U1820 (N_1820,In_4017,In_4470);
or U1821 (N_1821,In_2297,In_1240);
or U1822 (N_1822,In_1532,In_2357);
nand U1823 (N_1823,In_4562,In_3583);
or U1824 (N_1824,In_4060,In_397);
nor U1825 (N_1825,In_2031,In_4773);
and U1826 (N_1826,In_1150,In_4718);
and U1827 (N_1827,In_3516,In_2688);
nor U1828 (N_1828,In_3937,In_3016);
xnor U1829 (N_1829,In_4752,In_1624);
xnor U1830 (N_1830,In_336,In_2948);
xnor U1831 (N_1831,In_4906,In_3597);
xor U1832 (N_1832,In_3930,In_2112);
xor U1833 (N_1833,In_3602,In_1406);
or U1834 (N_1834,In_3118,In_3933);
and U1835 (N_1835,In_3146,In_1391);
and U1836 (N_1836,In_611,In_1033);
nor U1837 (N_1837,In_3351,In_1256);
nor U1838 (N_1838,In_3112,In_714);
nor U1839 (N_1839,In_4121,In_2186);
or U1840 (N_1840,In_3181,In_4412);
and U1841 (N_1841,In_3898,In_1795);
xor U1842 (N_1842,In_4409,In_2370);
and U1843 (N_1843,In_2209,In_801);
nor U1844 (N_1844,In_1008,In_3295);
and U1845 (N_1845,In_3865,In_2047);
xnor U1846 (N_1846,In_873,In_3416);
nor U1847 (N_1847,In_3409,In_4568);
nor U1848 (N_1848,In_2715,In_3501);
or U1849 (N_1849,In_1266,In_3722);
xor U1850 (N_1850,In_2884,In_963);
or U1851 (N_1851,In_3780,In_4753);
and U1852 (N_1852,In_2615,In_1271);
xor U1853 (N_1853,In_4392,In_535);
xnor U1854 (N_1854,In_181,In_3212);
xor U1855 (N_1855,In_567,In_1776);
nand U1856 (N_1856,In_1120,In_4900);
nor U1857 (N_1857,In_4156,In_849);
nand U1858 (N_1858,In_3560,In_2205);
or U1859 (N_1859,In_3134,In_368);
nand U1860 (N_1860,In_4775,In_406);
nor U1861 (N_1861,In_881,In_2545);
or U1862 (N_1862,In_649,In_131);
or U1863 (N_1863,In_197,In_1009);
or U1864 (N_1864,In_4929,In_443);
nand U1865 (N_1865,In_1957,In_572);
xnor U1866 (N_1866,In_332,In_2245);
nand U1867 (N_1867,In_2924,In_2010);
nor U1868 (N_1868,In_4532,In_4858);
or U1869 (N_1869,In_3380,In_4962);
and U1870 (N_1870,In_2028,In_3414);
xor U1871 (N_1871,In_1472,In_4070);
and U1872 (N_1872,In_2941,In_2084);
nor U1873 (N_1873,In_1453,In_4469);
nor U1874 (N_1874,In_1823,In_2604);
xnor U1875 (N_1875,In_4740,In_1486);
or U1876 (N_1876,In_2119,In_4557);
xor U1877 (N_1877,In_2120,In_3308);
nand U1878 (N_1878,In_1302,In_2220);
xnor U1879 (N_1879,In_3068,In_4471);
and U1880 (N_1880,In_4292,In_4424);
nand U1881 (N_1881,In_1612,In_4908);
and U1882 (N_1882,In_1927,In_505);
or U1883 (N_1883,In_3419,In_745);
nand U1884 (N_1884,In_3571,In_4128);
or U1885 (N_1885,In_71,In_2839);
nand U1886 (N_1886,In_3499,In_1923);
nor U1887 (N_1887,In_264,In_799);
xnor U1888 (N_1888,In_4256,In_1293);
nand U1889 (N_1889,In_2174,In_3469);
nand U1890 (N_1890,In_1924,In_1878);
nand U1891 (N_1891,In_1716,In_157);
nor U1892 (N_1892,In_1699,In_4400);
and U1893 (N_1893,In_2702,In_1137);
and U1894 (N_1894,In_3045,In_1858);
xor U1895 (N_1895,In_1288,In_4365);
nand U1896 (N_1896,In_4675,In_2923);
or U1897 (N_1897,In_1468,In_4946);
xnor U1898 (N_1898,In_2192,In_3989);
or U1899 (N_1899,In_2977,In_4910);
or U1900 (N_1900,In_4407,In_1161);
or U1901 (N_1901,In_2430,In_4604);
and U1902 (N_1902,In_1972,In_974);
and U1903 (N_1903,In_3675,In_3057);
nor U1904 (N_1904,In_2475,In_367);
xnor U1905 (N_1905,In_3464,In_1811);
xor U1906 (N_1906,In_2593,In_2893);
nand U1907 (N_1907,In_4990,In_1178);
nor U1908 (N_1908,In_2095,In_1226);
nand U1909 (N_1909,In_4596,In_3926);
nand U1910 (N_1910,In_1949,In_1953);
and U1911 (N_1911,In_1469,In_100);
nand U1912 (N_1912,In_4211,In_3042);
nand U1913 (N_1913,In_2129,In_1442);
or U1914 (N_1914,In_13,In_899);
and U1915 (N_1915,In_3226,In_2157);
nor U1916 (N_1916,In_412,In_1397);
and U1917 (N_1917,In_1913,In_777);
nor U1918 (N_1918,In_1159,In_4235);
nor U1919 (N_1919,In_631,In_1156);
nor U1920 (N_1920,In_366,In_4278);
xor U1921 (N_1921,In_355,In_2535);
and U1922 (N_1922,In_297,In_371);
nor U1923 (N_1923,In_235,In_3036);
or U1924 (N_1924,In_3170,In_1224);
nor U1925 (N_1925,In_3913,In_2967);
xnor U1926 (N_1926,In_4896,In_2693);
nor U1927 (N_1927,In_2616,In_4930);
nand U1928 (N_1928,In_4767,In_2936);
or U1929 (N_1929,In_2640,In_3757);
nand U1930 (N_1930,In_1623,In_3477);
or U1931 (N_1931,In_1671,In_3159);
or U1932 (N_1932,In_618,In_91);
nor U1933 (N_1933,In_2969,In_1042);
or U1934 (N_1934,In_2692,In_1259);
xnor U1935 (N_1935,In_1021,In_3279);
nand U1936 (N_1936,In_3348,In_1223);
nor U1937 (N_1937,In_724,In_4261);
or U1938 (N_1938,In_2108,In_1665);
and U1939 (N_1939,In_3983,In_496);
xor U1940 (N_1940,In_3956,In_4004);
xnor U1941 (N_1941,In_3097,In_4947);
or U1942 (N_1942,In_2853,In_1115);
xor U1943 (N_1943,In_3799,In_2149);
xnor U1944 (N_1944,In_3747,In_2399);
or U1945 (N_1945,In_2766,In_569);
or U1946 (N_1946,In_3894,In_3432);
or U1947 (N_1947,In_2566,In_3176);
nand U1948 (N_1948,In_1095,In_466);
nand U1949 (N_1949,In_1207,In_106);
or U1950 (N_1950,In_2234,In_703);
or U1951 (N_1951,In_2444,In_1701);
and U1952 (N_1952,In_2639,In_3696);
and U1953 (N_1953,In_313,In_1974);
or U1954 (N_1954,In_3523,In_876);
xnor U1955 (N_1955,In_4297,In_2455);
nand U1956 (N_1956,In_2780,In_292);
and U1957 (N_1957,In_358,In_4506);
and U1958 (N_1958,In_4732,In_3384);
or U1959 (N_1959,In_1160,In_4884);
and U1960 (N_1960,In_3461,In_1545);
nand U1961 (N_1961,In_4120,In_257);
and U1962 (N_1962,In_2187,In_307);
and U1963 (N_1963,In_1444,In_3197);
or U1964 (N_1964,In_3335,In_1387);
or U1965 (N_1965,In_2262,In_3811);
nor U1966 (N_1966,In_4646,In_1357);
xor U1967 (N_1967,In_1269,In_3730);
xor U1968 (N_1968,In_3594,In_81);
and U1969 (N_1969,In_394,In_1740);
nand U1970 (N_1970,In_2499,In_1757);
nor U1971 (N_1971,In_1572,In_4453);
nor U1972 (N_1972,In_2996,In_2127);
nor U1973 (N_1973,In_4541,In_3907);
nor U1974 (N_1974,In_782,In_301);
or U1975 (N_1975,In_3072,In_4720);
and U1976 (N_1976,In_3973,In_4214);
nor U1977 (N_1977,In_457,In_4854);
nand U1978 (N_1978,In_3554,In_3488);
nor U1979 (N_1979,In_177,In_3412);
nand U1980 (N_1980,In_1621,In_222);
nand U1981 (N_1981,In_3669,In_2382);
and U1982 (N_1982,In_4073,In_4885);
nand U1983 (N_1983,In_4094,In_3101);
xnor U1984 (N_1984,In_2554,In_3069);
nand U1985 (N_1985,In_2039,In_4762);
or U1986 (N_1986,In_3762,In_3995);
and U1987 (N_1987,In_2624,In_1124);
and U1988 (N_1988,In_2181,In_1653);
xor U1989 (N_1989,In_2865,In_2198);
or U1990 (N_1990,In_1978,In_2342);
nand U1991 (N_1991,In_3690,In_2292);
nand U1992 (N_1992,In_3083,In_3397);
or U1993 (N_1993,In_4181,In_1655);
and U1994 (N_1994,In_4377,In_4088);
nor U1995 (N_1995,In_3632,In_1354);
xnor U1996 (N_1996,In_4619,In_4770);
nor U1997 (N_1997,In_3451,In_4865);
and U1998 (N_1998,In_1741,In_4547);
xnor U1999 (N_1999,In_1576,In_3481);
or U2000 (N_2000,In_3807,In_3731);
nor U2001 (N_2001,In_1601,In_931);
and U2002 (N_2002,In_4584,In_4351);
xnor U2003 (N_2003,In_1356,In_1080);
and U2004 (N_2004,In_1948,In_4010);
and U2005 (N_2005,In_2681,In_1713);
nand U2006 (N_2006,In_4989,In_4656);
and U2007 (N_2007,In_1321,In_4245);
and U2008 (N_2008,In_2156,In_1950);
nor U2009 (N_2009,In_2665,In_1901);
and U2010 (N_2010,In_530,In_3564);
nor U2011 (N_2011,In_2147,In_4342);
nor U2012 (N_2012,In_339,In_238);
xnor U2013 (N_2013,In_3990,In_662);
nand U2014 (N_2014,In_1462,In_314);
or U2015 (N_2015,In_2408,In_409);
or U2016 (N_2016,In_2960,In_3857);
and U2017 (N_2017,In_4922,In_4206);
or U2018 (N_2018,In_3510,In_1104);
and U2019 (N_2019,In_3415,In_3861);
xnor U2020 (N_2020,In_1613,In_3603);
nor U2021 (N_2021,In_3389,In_0);
nand U2022 (N_2022,In_2758,In_2251);
and U2023 (N_2023,In_4153,In_473);
and U2024 (N_2024,In_2467,In_4146);
or U2025 (N_2025,In_243,In_270);
and U2026 (N_2026,In_3328,In_2389);
nand U2027 (N_2027,In_1303,In_3313);
nor U2028 (N_2028,In_1332,In_1599);
xor U2029 (N_2029,In_53,In_495);
and U2030 (N_2030,In_4023,In_4598);
nand U2031 (N_2031,In_384,In_2580);
xor U2032 (N_2032,In_589,In_1323);
and U2033 (N_2033,In_4667,In_2091);
xnor U2034 (N_2034,In_3169,In_3271);
and U2035 (N_2035,In_565,In_2679);
xnor U2036 (N_2036,In_3830,In_4632);
or U2037 (N_2037,In_689,In_4227);
and U2038 (N_2038,In_2492,In_4356);
nand U2039 (N_2039,In_3749,In_744);
xor U2040 (N_2040,In_3616,In_3164);
and U2041 (N_2041,In_3965,In_642);
nor U2042 (N_2042,In_79,In_4572);
nand U2043 (N_2043,In_311,In_4054);
nand U2044 (N_2044,In_932,In_2412);
nor U2045 (N_2045,In_104,In_1415);
and U2046 (N_2046,In_3465,In_1093);
or U2047 (N_2047,In_3664,In_1778);
nor U2048 (N_2048,In_3370,In_513);
or U2049 (N_2049,In_2073,In_520);
xor U2050 (N_2050,In_924,In_1329);
or U2051 (N_2051,In_2656,In_725);
nor U2052 (N_2052,In_1808,In_2906);
nor U2053 (N_2053,In_408,In_4126);
xor U2054 (N_2054,In_930,In_3378);
xor U2055 (N_2055,In_28,In_1869);
and U2056 (N_2056,In_2113,In_4493);
and U2057 (N_2057,In_874,In_2721);
nor U2058 (N_2058,In_1522,In_3048);
nor U2059 (N_2059,In_4616,In_3383);
xnor U2060 (N_2060,In_3077,In_695);
or U2061 (N_2061,In_712,In_4628);
xnor U2062 (N_2062,In_1049,In_112);
or U2063 (N_2063,In_41,In_2071);
nand U2064 (N_2064,In_2976,In_4095);
or U2065 (N_2065,In_1796,In_3280);
and U2066 (N_2066,In_3618,In_4977);
or U2067 (N_2067,In_4482,In_1112);
xor U2068 (N_2068,In_1774,In_785);
nand U2069 (N_2069,In_4249,In_1059);
xnor U2070 (N_2070,In_4941,In_3175);
or U2071 (N_2071,In_290,In_2287);
nand U2072 (N_2072,In_2451,In_2754);
or U2073 (N_2073,In_4062,In_196);
xnor U2074 (N_2074,In_4240,In_2061);
nor U2075 (N_2075,In_4594,In_3217);
xnor U2076 (N_2076,In_1751,In_431);
or U2077 (N_2077,In_3269,In_1283);
nor U2078 (N_2078,In_3189,In_586);
xor U2079 (N_2079,In_357,In_1822);
and U2080 (N_2080,In_3491,In_2041);
xor U2081 (N_2081,In_4209,In_1709);
nand U2082 (N_2082,In_2086,In_98);
nor U2083 (N_2083,In_4496,In_4798);
nor U2084 (N_2084,In_2237,In_446);
nor U2085 (N_2085,In_425,In_2588);
nor U2086 (N_2086,In_2212,In_3598);
nand U2087 (N_2087,In_1739,In_4515);
nor U2088 (N_2088,In_908,In_4020);
and U2089 (N_2089,In_3960,In_4138);
or U2090 (N_2090,In_2974,In_1083);
nand U2091 (N_2091,In_272,In_2907);
xnor U2092 (N_2092,In_2992,In_3369);
and U2093 (N_2093,In_1298,In_3270);
xnor U2094 (N_2094,In_1958,In_449);
nor U2095 (N_2095,In_1094,In_925);
or U2096 (N_2096,In_4520,In_1078);
nand U2097 (N_2097,In_897,In_1182);
nor U2098 (N_2098,In_3745,In_4692);
or U2099 (N_2099,In_3349,In_4087);
xnor U2100 (N_2100,In_4992,In_1938);
nand U2101 (N_2101,In_2783,In_4237);
or U2102 (N_2102,In_4440,In_3496);
nor U2103 (N_2103,In_2938,In_683);
nand U2104 (N_2104,In_2454,In_608);
nor U2105 (N_2105,In_4570,In_4722);
nand U2106 (N_2106,In_3133,In_1955);
nand U2107 (N_2107,In_2641,In_3340);
xor U2108 (N_2108,In_4195,In_2744);
or U2109 (N_2109,In_461,In_2745);
or U2110 (N_2110,In_4563,In_470);
xor U2111 (N_2111,In_84,In_3095);
or U2112 (N_2112,In_3741,In_1529);
nand U2113 (N_2113,In_1155,In_2903);
and U2114 (N_2114,In_3800,In_3843);
nor U2115 (N_2115,In_1447,In_2068);
and U2116 (N_2116,In_4086,In_4063);
nor U2117 (N_2117,In_2288,In_3532);
xnor U2118 (N_2118,In_4685,In_1815);
xnor U2119 (N_2119,In_163,In_2057);
and U2120 (N_2120,In_3223,In_2993);
or U2121 (N_2121,In_802,In_719);
and U2122 (N_2122,In_4859,In_2984);
or U2123 (N_2123,In_2747,In_659);
nor U2124 (N_2124,In_4825,In_3549);
or U2125 (N_2125,In_4809,In_778);
or U2126 (N_2126,In_598,In_369);
nor U2127 (N_2127,In_1214,In_2423);
and U2128 (N_2128,In_1590,In_2515);
and U2129 (N_2129,In_4768,In_959);
nand U2130 (N_2130,In_731,In_3887);
and U2131 (N_2131,In_3517,In_4166);
or U2132 (N_2132,In_822,In_1452);
nor U2133 (N_2133,In_2009,In_4191);
or U2134 (N_2134,In_1167,In_984);
and U2135 (N_2135,In_3557,In_3738);
nor U2136 (N_2136,In_246,In_1862);
and U2137 (N_2137,In_4103,In_1588);
or U2138 (N_2138,In_1860,In_3522);
nor U2139 (N_2139,In_1111,In_2343);
nor U2140 (N_2140,In_1097,In_2603);
xnor U2141 (N_2141,In_4551,In_3366);
and U2142 (N_2142,In_3423,In_892);
xnor U2143 (N_2143,In_2380,In_4874);
xor U2144 (N_2144,In_3035,In_1440);
or U2145 (N_2145,In_2858,In_4057);
nor U2146 (N_2146,In_2339,In_576);
nor U2147 (N_2147,In_4081,In_600);
and U2148 (N_2148,In_1785,In_1361);
nor U2149 (N_2149,In_677,In_4137);
nor U2150 (N_2150,In_2240,In_1029);
and U2151 (N_2151,In_652,In_194);
and U2152 (N_2152,In_2551,In_3820);
nor U2153 (N_2153,In_4085,In_969);
nor U2154 (N_2154,In_1969,In_2378);
and U2155 (N_2155,In_1409,In_718);
nand U2156 (N_2156,In_4188,In_4918);
nor U2157 (N_2157,In_3902,In_4267);
nand U2158 (N_2158,In_78,In_3353);
or U2159 (N_2159,In_3821,In_669);
xnor U2160 (N_2160,In_1198,In_4712);
or U2161 (N_2161,In_3886,In_1630);
or U2162 (N_2162,In_1229,In_2652);
xnor U2163 (N_2163,In_791,In_522);
and U2164 (N_2164,In_2200,In_3804);
and U2165 (N_2165,In_2832,In_3750);
and U2166 (N_2166,In_329,In_4812);
and U2167 (N_2167,In_4065,In_3927);
nor U2168 (N_2168,In_2997,In_3187);
or U2169 (N_2169,In_3982,In_1039);
xor U2170 (N_2170,In_4987,In_4334);
nand U2171 (N_2171,In_4624,In_4666);
or U2172 (N_2172,In_4610,In_1062);
or U2173 (N_2173,In_4959,In_331);
xor U2174 (N_2174,In_2121,In_1380);
nor U2175 (N_2175,In_2336,In_1151);
nand U2176 (N_2176,In_3945,In_884);
and U2177 (N_2177,In_381,In_2511);
and U2178 (N_2178,In_4243,In_2540);
nand U2179 (N_2179,In_1507,In_2447);
nor U2180 (N_2180,In_1841,In_2356);
nand U2181 (N_2181,In_2248,In_1177);
nand U2182 (N_2182,In_1875,In_1920);
or U2183 (N_2183,In_3925,In_3763);
xor U2184 (N_2184,In_937,In_4509);
and U2185 (N_2185,In_2309,In_405);
and U2186 (N_2186,In_961,In_2106);
nand U2187 (N_2187,In_1273,In_2460);
nand U2188 (N_2188,In_2625,In_2577);
or U2189 (N_2189,In_4797,In_3565);
or U2190 (N_2190,In_4864,In_102);
or U2191 (N_2191,In_3682,In_1762);
nor U2192 (N_2192,In_1484,In_2733);
nor U2193 (N_2193,In_1853,In_2014);
and U2194 (N_2194,In_3362,In_219);
nand U2195 (N_2195,In_2687,In_216);
or U2196 (N_2196,In_2101,In_1787);
nand U2197 (N_2197,In_4926,In_4155);
or U2198 (N_2198,In_4587,In_571);
and U2199 (N_2199,In_1040,In_94);
nand U2200 (N_2200,In_2777,In_3915);
xnor U2201 (N_2201,In_4021,In_4326);
nand U2202 (N_2202,In_266,In_3700);
nor U2203 (N_2203,In_531,In_2877);
nand U2204 (N_2204,In_2613,In_710);
nor U2205 (N_2205,In_4395,In_4731);
or U2206 (N_2206,In_3492,In_3060);
xor U2207 (N_2207,In_4372,In_2376);
xor U2208 (N_2208,In_3184,In_3903);
xnor U2209 (N_2209,In_1935,In_2153);
or U2210 (N_2210,In_3387,In_570);
and U2211 (N_2211,In_3794,In_2440);
xor U2212 (N_2212,In_1117,In_1528);
or U2213 (N_2213,In_4125,In_4182);
nor U2214 (N_2214,In_169,In_1386);
or U2215 (N_2215,In_3426,In_3482);
and U2216 (N_2216,In_4935,In_996);
or U2217 (N_2217,In_445,In_176);
or U2218 (N_2218,In_2553,In_650);
xor U2219 (N_2219,In_4957,In_1847);
xor U2220 (N_2220,In_3878,In_3676);
or U2221 (N_2221,In_4408,In_2398);
xor U2222 (N_2222,In_1542,In_1239);
nor U2223 (N_2223,In_2677,In_29);
nand U2224 (N_2224,In_4431,In_617);
xor U2225 (N_2225,In_2536,In_4404);
and U2226 (N_2226,In_4579,In_4102);
and U2227 (N_2227,In_2918,In_1147);
or U2228 (N_2228,In_1719,In_1939);
nor U2229 (N_2229,In_2601,In_1005);
xor U2230 (N_2230,In_2516,In_4238);
xor U2231 (N_2231,In_2782,In_736);
or U2232 (N_2232,In_2636,In_303);
and U2233 (N_2233,In_4189,In_861);
xnor U2234 (N_2234,In_2546,In_2473);
nor U2235 (N_2235,In_3694,In_4106);
and U2236 (N_2236,In_1563,In_4316);
xnor U2237 (N_2237,In_2626,In_4523);
or U2238 (N_2238,In_3822,In_1125);
or U2239 (N_2239,In_2373,In_143);
nor U2240 (N_2240,In_3323,In_713);
nand U2241 (N_2241,In_1977,In_1322);
or U2242 (N_2242,In_1070,In_1677);
xnor U2243 (N_2243,In_2230,In_363);
or U2244 (N_2244,In_1673,In_768);
xnor U2245 (N_2245,In_4960,In_4779);
xnor U2246 (N_2246,In_3992,In_3347);
nand U2247 (N_2247,In_2922,In_1367);
nand U2248 (N_2248,In_3785,In_4039);
xnor U2249 (N_2249,In_4140,In_1162);
nor U2250 (N_2250,In_3334,In_2066);
nand U2251 (N_2251,In_3765,In_2161);
and U2252 (N_2252,In_4704,In_4870);
and U2253 (N_2253,In_843,In_468);
nor U2254 (N_2254,In_3712,In_3438);
or U2255 (N_2255,In_4091,In_2584);
xnor U2256 (N_2256,In_747,In_2004);
xnor U2257 (N_2257,In_1874,In_1360);
and U2258 (N_2258,In_4891,In_722);
or U2259 (N_2259,In_4028,In_4697);
nand U2260 (N_2260,In_789,In_1770);
nor U2261 (N_2261,In_2301,In_4291);
and U2262 (N_2262,In_1248,In_2142);
or U2263 (N_2263,In_2193,In_2685);
nor U2264 (N_2264,In_1421,In_4979);
or U2265 (N_2265,In_504,In_2385);
or U2266 (N_2266,In_241,In_2457);
nand U2267 (N_2267,In_4025,In_1947);
or U2268 (N_2268,In_610,In_2773);
xor U2269 (N_2269,In_1341,In_4764);
and U2270 (N_2270,In_1267,In_1204);
nand U2271 (N_2271,In_3247,In_3919);
nand U2272 (N_2272,In_1166,In_3300);
nor U2273 (N_2273,In_3661,In_1777);
nor U2274 (N_2274,In_1165,In_775);
or U2275 (N_2275,In_1802,In_614);
or U2276 (N_2276,In_3567,In_255);
xnor U2277 (N_2277,In_2632,In_4919);
nor U2278 (N_2278,In_1471,In_4567);
or U2279 (N_2279,In_1894,In_4451);
nand U2280 (N_2280,In_260,In_1617);
xnor U2281 (N_2281,In_1216,In_2876);
xor U2282 (N_2282,In_1839,In_1297);
and U2283 (N_2283,In_1141,In_4980);
nor U2284 (N_2284,In_4130,In_4794);
xor U2285 (N_2285,In_3211,In_2330);
or U2286 (N_2286,In_545,In_752);
nand U2287 (N_2287,In_2132,In_3345);
and U2288 (N_2288,In_2239,In_4953);
nand U2289 (N_2289,In_204,In_4967);
xor U2290 (N_2290,In_3627,In_1055);
nand U2291 (N_2291,In_4660,In_132);
and U2292 (N_2292,In_1443,In_2428);
nor U2293 (N_2293,In_4305,In_2945);
xor U2294 (N_2294,In_1218,In_1278);
nand U2295 (N_2295,In_230,In_721);
nor U2296 (N_2296,In_3617,In_3681);
nand U2297 (N_2297,In_4671,In_960);
nor U2298 (N_2298,In_3559,In_2402);
and U2299 (N_2299,In_3900,In_4269);
nor U2300 (N_2300,In_3558,In_811);
or U2301 (N_2301,In_4338,In_1076);
nor U2302 (N_2302,In_2371,In_2128);
and U2303 (N_2303,In_2,In_641);
nor U2304 (N_2304,In_1593,In_4699);
nand U2305 (N_2305,In_1114,In_1700);
nor U2306 (N_2306,In_3040,In_859);
nor U2307 (N_2307,In_1914,In_2407);
xor U2308 (N_2308,In_2910,In_2598);
or U2309 (N_2309,In_670,In_2576);
nor U2310 (N_2310,In_2987,In_278);
nor U2311 (N_2311,In_390,In_1889);
nand U2312 (N_2312,In_2489,In_4664);
and U2313 (N_2313,In_1800,In_2439);
or U2314 (N_2314,In_2130,In_437);
nand U2315 (N_2315,In_2957,In_4629);
and U2316 (N_2316,In_362,In_4925);
nand U2317 (N_2317,In_845,In_3365);
and U2318 (N_2318,In_480,In_2950);
and U2319 (N_2319,In_448,In_1252);
and U2320 (N_2320,In_815,In_2873);
nand U2321 (N_2321,In_4367,In_521);
nor U2322 (N_2322,In_3703,In_2662);
nor U2323 (N_2323,In_2470,In_2510);
or U2324 (N_2324,In_4452,In_3997);
xnor U2325 (N_2325,In_4402,In_4255);
and U2326 (N_2326,In_2203,In_4894);
xnor U2327 (N_2327,In_4507,In_1265);
nor U2328 (N_2328,In_3966,In_1667);
or U2329 (N_2329,In_1637,In_711);
nor U2330 (N_2330,In_3810,In_538);
nor U2331 (N_2331,In_4522,In_488);
nand U2332 (N_2332,In_145,In_1684);
xnor U2333 (N_2333,In_3707,In_1001);
nor U2334 (N_2334,In_433,In_1377);
xnor U2335 (N_2335,In_1755,In_4465);
or U2336 (N_2336,In_494,In_1163);
nand U2337 (N_2337,In_2377,In_750);
xor U2338 (N_2338,In_3846,In_4975);
nor U2339 (N_2339,In_654,In_2949);
nor U2340 (N_2340,In_726,In_935);
nand U2341 (N_2341,In_1917,In_2289);
nor U2342 (N_2342,In_1994,In_3240);
nand U2343 (N_2343,In_3599,In_3998);
and U2344 (N_2344,In_970,In_4437);
or U2345 (N_2345,In_3576,In_4652);
nand U2346 (N_2346,In_1554,In_1810);
xor U2347 (N_2347,In_3521,In_1481);
xor U2348 (N_2348,In_3372,In_242);
or U2349 (N_2349,In_1195,In_890);
nand U2350 (N_2350,In_2901,In_1047);
nand U2351 (N_2351,In_2417,In_3595);
xnor U2352 (N_2352,In_3601,In_1011);
and U2353 (N_2353,In_803,In_2434);
or U2354 (N_2354,In_1736,In_1771);
and U2355 (N_2355,In_4593,In_841);
and U2356 (N_2356,In_4867,In_2557);
or U2357 (N_2357,In_3537,In_3049);
and U2358 (N_2358,In_223,In_49);
xor U2359 (N_2359,In_1024,In_3984);
nand U2360 (N_2360,In_2635,In_2479);
nand U2361 (N_2361,In_2522,In_4807);
xor U2362 (N_2362,In_419,In_3589);
or U2363 (N_2363,In_1622,In_2006);
or U2364 (N_2364,In_2857,In_1109);
nor U2365 (N_2365,In_2544,In_4542);
xor U2366 (N_2366,In_1760,In_3833);
nor U2367 (N_2367,In_365,In_3691);
nand U2368 (N_2368,In_225,In_3120);
xor U2369 (N_2369,In_1817,In_3171);
nor U2370 (N_2370,In_3850,In_3977);
xor U2371 (N_2371,In_4618,In_3196);
or U2372 (N_2372,In_3156,In_2563);
nor U2373 (N_2373,In_21,In_1830);
or U2374 (N_2374,In_1131,In_978);
xor U2375 (N_2375,In_416,In_1400);
nand U2376 (N_2376,In_108,In_4202);
nor U2377 (N_2377,In_880,In_2093);
or U2378 (N_2378,In_229,In_1434);
and U2379 (N_2379,In_4538,In_4696);
xnor U2380 (N_2380,In_2384,In_2481);
or U2381 (N_2381,In_1899,In_4477);
nand U2382 (N_2382,In_1069,In_3390);
and U2383 (N_2383,In_3044,In_146);
or U2384 (N_2384,In_1866,In_4543);
nor U2385 (N_2385,In_2166,In_3688);
xor U2386 (N_2386,In_1918,In_200);
and U2387 (N_2387,In_1310,In_1644);
and U2388 (N_2388,In_174,In_523);
and U2389 (N_2389,In_4686,In_746);
and U2390 (N_2390,In_3775,In_3923);
nor U2391 (N_2391,In_2574,In_3487);
nand U2392 (N_2392,In_1929,In_3835);
nand U2393 (N_2393,In_273,In_1756);
and U2394 (N_2394,In_878,In_3663);
and U2395 (N_2395,In_361,In_1473);
or U2396 (N_2396,In_4681,In_647);
or U2397 (N_2397,In_4778,In_1180);
or U2398 (N_2398,In_707,In_1145);
nand U2399 (N_2399,In_2202,In_3709);
xnor U2400 (N_2400,In_912,In_3396);
xor U2401 (N_2401,In_3264,In_1168);
and U2402 (N_2402,In_3976,In_1524);
xnor U2403 (N_2403,In_812,In_3959);
nor U2404 (N_2404,In_3852,In_1003);
xnor U2405 (N_2405,In_4280,In_2956);
nor U2406 (N_2406,In_1064,In_3428);
xnor U2407 (N_2407,In_2846,In_2697);
nor U2408 (N_2408,In_1546,In_487);
xor U2409 (N_2409,In_1164,In_1629);
nand U2410 (N_2410,In_4845,In_1379);
xor U2411 (N_2411,In_3050,In_2596);
xnor U2412 (N_2412,In_348,In_4344);
nor U2413 (N_2413,In_2088,In_1154);
nand U2414 (N_2414,In_279,In_813);
nor U2415 (N_2415,In_2788,In_2471);
nand U2416 (N_2416,In_2141,In_3610);
nand U2417 (N_2417,In_2847,In_1234);
nor U2418 (N_2418,In_1050,In_605);
nand U2419 (N_2419,In_244,In_732);
and U2420 (N_2420,In_1384,In_4909);
xor U2421 (N_2421,In_1674,In_4230);
xnor U2422 (N_2422,In_1625,In_1317);
nor U2423 (N_2423,In_987,In_1353);
or U2424 (N_2424,In_3590,In_694);
nor U2425 (N_2425,In_3363,In_4036);
xnor U2426 (N_2426,In_1082,In_2329);
nor U2427 (N_2427,In_1712,In_839);
nand U2428 (N_2428,In_3967,In_1743);
nor U2429 (N_2429,In_4001,In_4311);
and U2430 (N_2430,In_1681,In_4100);
and U2431 (N_2431,In_585,In_3635);
nand U2432 (N_2432,In_2528,In_3326);
or U2433 (N_2433,In_3920,In_1338);
or U2434 (N_2434,In_4183,In_663);
xnor U2435 (N_2435,In_3063,In_4244);
nand U2436 (N_2436,In_210,In_42);
or U2437 (N_2437,In_2669,In_1921);
or U2438 (N_2438,In_901,In_2299);
nor U2439 (N_2439,In_939,In_1990);
nor U2440 (N_2440,In_3436,In_4381);
or U2441 (N_2441,In_1807,In_373);
nand U2442 (N_2442,In_3258,In_2537);
nand U2443 (N_2443,In_3874,In_2682);
nor U2444 (N_2444,In_1512,In_1233);
or U2445 (N_2445,In_3805,In_4881);
or U2446 (N_2446,In_3082,In_4317);
and U2447 (N_2447,In_2845,In_4016);
xor U2448 (N_2448,In_2191,In_2507);
nand U2449 (N_2449,In_1087,In_2401);
xor U2450 (N_2450,In_1976,In_478);
nor U2451 (N_2451,In_1975,In_2986);
nand U2452 (N_2452,In_2645,In_4040);
and U2453 (N_2453,In_2247,In_1884);
and U2454 (N_2454,In_3881,In_252);
nand U2455 (N_2455,In_1250,In_4308);
nor U2456 (N_2456,In_2154,In_1693);
nor U2457 (N_2457,In_3773,In_4174);
xor U2458 (N_2458,In_4678,In_2792);
nor U2459 (N_2459,In_3005,In_2842);
nor U2460 (N_2460,In_391,In_2803);
nor U2461 (N_2461,In_3298,In_3655);
nand U2462 (N_2462,In_2518,In_3454);
and U2463 (N_2463,In_153,In_1477);
nor U2464 (N_2464,In_4711,In_3332);
or U2465 (N_2465,In_1744,In_575);
or U2466 (N_2466,In_1308,In_781);
or U2467 (N_2467,In_4658,In_2355);
nand U2468 (N_2468,In_3922,In_4253);
and U2469 (N_2469,In_2724,In_682);
nor U2470 (N_2470,In_770,In_2497);
xor U2471 (N_2471,In_4556,In_1208);
and U2472 (N_2472,In_3455,In_4782);
and U2473 (N_2473,In_2226,In_4950);
nand U2474 (N_2474,In_1560,In_534);
nor U2475 (N_2475,In_882,In_2952);
and U2476 (N_2476,In_2618,In_4464);
nor U2477 (N_2477,In_1691,In_2158);
nand U2478 (N_2478,In_1711,In_4347);
nand U2479 (N_2479,In_4179,In_4222);
xnor U2480 (N_2480,In_927,In_933);
xor U2481 (N_2481,In_1004,In_4076);
or U2482 (N_2482,In_3659,In_2252);
or U2483 (N_2483,In_1202,In_1022);
nand U2484 (N_2484,In_2294,In_63);
xnor U2485 (N_2485,In_1531,In_1394);
xnor U2486 (N_2486,In_1171,In_1200);
or U2487 (N_2487,In_3764,In_868);
and U2488 (N_2488,In_2825,In_2983);
and U2489 (N_2489,In_2589,In_599);
and U2490 (N_2490,In_2525,In_2951);
nand U2491 (N_2491,In_2633,In_1846);
and U2492 (N_2492,In_353,In_3427);
and U2493 (N_2493,In_877,In_3186);
nor U2494 (N_2494,In_2274,In_4220);
nand U2495 (N_2495,In_2805,In_2078);
nand U2496 (N_2496,In_885,In_3107);
and U2497 (N_2497,In_615,In_305);
nor U2498 (N_2498,In_2502,In_3219);
or U2499 (N_2499,In_4053,In_4024);
nor U2500 (N_2500,N_2066,N_2419);
nor U2501 (N_2501,N_2374,N_151);
nand U2502 (N_2502,N_2369,N_2156);
nand U2503 (N_2503,N_2287,N_2462);
xnor U2504 (N_2504,N_2250,N_539);
or U2505 (N_2505,N_771,N_2045);
nor U2506 (N_2506,N_140,N_2426);
or U2507 (N_2507,N_1695,N_1441);
xor U2508 (N_2508,N_2327,N_1212);
or U2509 (N_2509,N_1324,N_2433);
xor U2510 (N_2510,N_2228,N_349);
nor U2511 (N_2511,N_629,N_283);
nand U2512 (N_2512,N_847,N_264);
nand U2513 (N_2513,N_895,N_458);
and U2514 (N_2514,N_1856,N_304);
or U2515 (N_2515,N_1048,N_2447);
nand U2516 (N_2516,N_2354,N_45);
or U2517 (N_2517,N_2108,N_1613);
nor U2518 (N_2518,N_1699,N_1250);
or U2519 (N_2519,N_250,N_514);
and U2520 (N_2520,N_576,N_1591);
or U2521 (N_2521,N_1887,N_1209);
xnor U2522 (N_2522,N_125,N_647);
and U2523 (N_2523,N_1682,N_2193);
or U2524 (N_2524,N_2283,N_1336);
nand U2525 (N_2525,N_358,N_1111);
nor U2526 (N_2526,N_1127,N_2188);
xor U2527 (N_2527,N_2202,N_1744);
and U2528 (N_2528,N_957,N_1327);
nand U2529 (N_2529,N_996,N_326);
or U2530 (N_2530,N_1155,N_750);
and U2531 (N_2531,N_496,N_317);
xor U2532 (N_2532,N_880,N_2006);
nor U2533 (N_2533,N_1804,N_679);
nor U2534 (N_2534,N_1708,N_707);
nor U2535 (N_2535,N_297,N_1538);
nand U2536 (N_2536,N_1407,N_1879);
or U2537 (N_2537,N_1383,N_787);
nand U2538 (N_2538,N_2438,N_2105);
nand U2539 (N_2539,N_1476,N_2377);
xnor U2540 (N_2540,N_362,N_2449);
xor U2541 (N_2541,N_160,N_1082);
nand U2542 (N_2542,N_1663,N_1686);
nand U2543 (N_2543,N_1422,N_2382);
nor U2544 (N_2544,N_1420,N_2311);
nor U2545 (N_2545,N_25,N_294);
and U2546 (N_2546,N_240,N_1430);
and U2547 (N_2547,N_2145,N_1331);
nand U2548 (N_2548,N_1805,N_1593);
nor U2549 (N_2549,N_1845,N_1588);
or U2550 (N_2550,N_24,N_1627);
nand U2551 (N_2551,N_2097,N_2071);
xor U2552 (N_2552,N_1519,N_1330);
xor U2553 (N_2553,N_432,N_216);
nand U2554 (N_2554,N_2392,N_836);
or U2555 (N_2555,N_995,N_15);
nor U2556 (N_2556,N_614,N_1329);
and U2557 (N_2557,N_1916,N_281);
nand U2558 (N_2558,N_318,N_2139);
and U2559 (N_2559,N_1537,N_1562);
nor U2560 (N_2560,N_2185,N_422);
and U2561 (N_2561,N_584,N_99);
nand U2562 (N_2562,N_2302,N_1942);
nor U2563 (N_2563,N_2015,N_1444);
or U2564 (N_2564,N_873,N_765);
xnor U2565 (N_2565,N_1634,N_1950);
xnor U2566 (N_2566,N_319,N_2348);
nand U2567 (N_2567,N_988,N_1700);
xor U2568 (N_2568,N_1262,N_2397);
or U2569 (N_2569,N_2305,N_123);
or U2570 (N_2570,N_2220,N_2047);
and U2571 (N_2571,N_2435,N_1497);
nand U2572 (N_2572,N_1857,N_1599);
xor U2573 (N_2573,N_727,N_1689);
nand U2574 (N_2574,N_1174,N_133);
xor U2575 (N_2575,N_1450,N_1892);
and U2576 (N_2576,N_646,N_909);
or U2577 (N_2577,N_2300,N_922);
and U2578 (N_2578,N_1069,N_1360);
xor U2579 (N_2579,N_343,N_1439);
or U2580 (N_2580,N_2159,N_1506);
nand U2581 (N_2581,N_591,N_1964);
xnor U2582 (N_2582,N_2129,N_1650);
or U2583 (N_2583,N_2475,N_2352);
and U2584 (N_2584,N_2288,N_2386);
nand U2585 (N_2585,N_1211,N_2488);
xor U2586 (N_2586,N_1371,N_969);
or U2587 (N_2587,N_2445,N_2349);
or U2588 (N_2588,N_558,N_1823);
and U2589 (N_2589,N_2016,N_1995);
and U2590 (N_2590,N_144,N_1148);
nand U2591 (N_2591,N_1966,N_1931);
or U2592 (N_2592,N_1363,N_2039);
nand U2593 (N_2593,N_472,N_1306);
nand U2594 (N_2594,N_156,N_1190);
or U2595 (N_2595,N_1886,N_774);
or U2596 (N_2596,N_73,N_1577);
or U2597 (N_2597,N_1844,N_1);
nand U2598 (N_2598,N_1676,N_293);
nand U2599 (N_2599,N_876,N_1642);
or U2600 (N_2600,N_590,N_74);
nand U2601 (N_2601,N_218,N_1559);
nand U2602 (N_2602,N_1314,N_2366);
xor U2603 (N_2603,N_1935,N_2079);
and U2604 (N_2604,N_1426,N_2153);
nand U2605 (N_2605,N_824,N_286);
and U2606 (N_2606,N_639,N_2215);
or U2607 (N_2607,N_2028,N_917);
xnor U2608 (N_2608,N_1909,N_2029);
nand U2609 (N_2609,N_1630,N_738);
nand U2610 (N_2610,N_2492,N_2083);
or U2611 (N_2611,N_1761,N_26);
and U2612 (N_2612,N_812,N_903);
or U2613 (N_2613,N_1767,N_637);
nand U2614 (N_2614,N_1375,N_1685);
nor U2615 (N_2615,N_1723,N_1432);
nor U2616 (N_2616,N_2081,N_1876);
or U2617 (N_2617,N_2428,N_436);
and U2618 (N_2618,N_86,N_2424);
xnor U2619 (N_2619,N_1822,N_1645);
nand U2620 (N_2620,N_1002,N_2107);
xor U2621 (N_2621,N_385,N_1745);
or U2622 (N_2622,N_897,N_212);
nand U2623 (N_2623,N_1267,N_635);
nor U2624 (N_2624,N_2063,N_848);
xnor U2625 (N_2625,N_1080,N_656);
nand U2626 (N_2626,N_1332,N_1833);
nand U2627 (N_2627,N_1753,N_1572);
nand U2628 (N_2628,N_1527,N_731);
nor U2629 (N_2629,N_85,N_985);
nand U2630 (N_2630,N_1200,N_2058);
or U2631 (N_2631,N_1696,N_2109);
and U2632 (N_2632,N_1516,N_729);
nand U2633 (N_2633,N_2358,N_2114);
and U2634 (N_2634,N_693,N_2450);
and U2635 (N_2635,N_921,N_456);
or U2636 (N_2636,N_1567,N_2344);
and U2637 (N_2637,N_2260,N_469);
or U2638 (N_2638,N_440,N_1096);
or U2639 (N_2639,N_2399,N_538);
and U2640 (N_2640,N_1937,N_1722);
and U2641 (N_2641,N_1277,N_615);
xnor U2642 (N_2642,N_2387,N_435);
nand U2643 (N_2643,N_1166,N_583);
and U2644 (N_2644,N_136,N_1926);
nand U2645 (N_2645,N_1121,N_1883);
xor U2646 (N_2646,N_1142,N_2255);
and U2647 (N_2647,N_793,N_367);
nor U2648 (N_2648,N_1489,N_1812);
or U2649 (N_2649,N_1272,N_406);
or U2650 (N_2650,N_791,N_1756);
and U2651 (N_2651,N_509,N_288);
nor U2652 (N_2652,N_124,N_1204);
xnor U2653 (N_2653,N_2204,N_579);
or U2654 (N_2654,N_2406,N_2012);
xnor U2655 (N_2655,N_806,N_0);
nor U2656 (N_2656,N_2365,N_1421);
and U2657 (N_2657,N_1299,N_17);
xor U2658 (N_2658,N_1921,N_284);
nand U2659 (N_2659,N_1818,N_1651);
or U2660 (N_2660,N_1367,N_2163);
nand U2661 (N_2661,N_580,N_1629);
and U2662 (N_2662,N_1657,N_1618);
or U2663 (N_2663,N_723,N_2235);
nor U2664 (N_2664,N_1633,N_360);
nor U2665 (N_2665,N_519,N_1241);
nor U2666 (N_2666,N_1218,N_2431);
xor U2667 (N_2667,N_933,N_461);
and U2668 (N_2668,N_612,N_950);
xor U2669 (N_2669,N_1265,N_1092);
nor U2670 (N_2670,N_2154,N_855);
and U2671 (N_2671,N_1568,N_744);
xnor U2672 (N_2672,N_1953,N_555);
nor U2673 (N_2673,N_2142,N_947);
xor U2674 (N_2674,N_1859,N_2179);
nor U2675 (N_2675,N_1967,N_2017);
and U2676 (N_2676,N_1456,N_1674);
nand U2677 (N_2677,N_736,N_1793);
or U2678 (N_2678,N_912,N_1819);
or U2679 (N_2679,N_681,N_941);
nor U2680 (N_2680,N_2342,N_2234);
nor U2681 (N_2681,N_1714,N_1044);
xnor U2682 (N_2682,N_2379,N_1291);
and U2683 (N_2683,N_900,N_1763);
nand U2684 (N_2684,N_832,N_715);
and U2685 (N_2685,N_117,N_543);
xnor U2686 (N_2686,N_2330,N_1881);
nor U2687 (N_2687,N_2262,N_1312);
nor U2688 (N_2688,N_607,N_1298);
or U2689 (N_2689,N_1370,N_147);
xnor U2690 (N_2690,N_2242,N_2239);
nor U2691 (N_2691,N_797,N_134);
or U2692 (N_2692,N_676,N_1943);
or U2693 (N_2693,N_2138,N_1335);
xnor U2694 (N_2694,N_673,N_926);
or U2695 (N_2695,N_2044,N_976);
and U2696 (N_2696,N_2090,N_672);
nor U2697 (N_2697,N_2225,N_640);
xnor U2698 (N_2698,N_1601,N_1956);
nor U2699 (N_2699,N_739,N_9);
nand U2700 (N_2700,N_2496,N_2294);
nand U2701 (N_2701,N_2151,N_2162);
xor U2702 (N_2702,N_239,N_1374);
xor U2703 (N_2703,N_708,N_572);
or U2704 (N_2704,N_98,N_1068);
or U2705 (N_2705,N_1855,N_467);
nand U2706 (N_2706,N_405,N_1973);
xor U2707 (N_2707,N_1998,N_746);
nor U2708 (N_2708,N_2391,N_2062);
nor U2709 (N_2709,N_1194,N_2446);
nand U2710 (N_2710,N_1283,N_520);
or U2711 (N_2711,N_799,N_770);
and U2712 (N_2712,N_1436,N_2254);
nor U2713 (N_2713,N_113,N_1609);
xor U2714 (N_2714,N_153,N_998);
or U2715 (N_2715,N_1491,N_1452);
and U2716 (N_2716,N_2415,N_1032);
nor U2717 (N_2717,N_798,N_820);
and U2718 (N_2718,N_534,N_1776);
xnor U2719 (N_2719,N_1196,N_409);
xor U2720 (N_2720,N_532,N_357);
nand U2721 (N_2721,N_71,N_1488);
nand U2722 (N_2722,N_1365,N_1109);
nor U2723 (N_2723,N_227,N_1135);
nor U2724 (N_2724,N_101,N_187);
nand U2725 (N_2725,N_1631,N_1564);
nand U2726 (N_2726,N_130,N_2307);
nor U2727 (N_2727,N_1297,N_2059);
and U2728 (N_2728,N_2216,N_1052);
nor U2729 (N_2729,N_800,N_2181);
nand U2730 (N_2730,N_821,N_2346);
or U2731 (N_2731,N_1888,N_337);
nand U2732 (N_2732,N_63,N_709);
and U2733 (N_2733,N_172,N_2310);
or U2734 (N_2734,N_875,N_1992);
or U2735 (N_2735,N_1428,N_400);
or U2736 (N_2736,N_2416,N_2296);
nand U2737 (N_2737,N_1097,N_316);
nand U2738 (N_2738,N_1573,N_1120);
nor U2739 (N_2739,N_366,N_137);
or U2740 (N_2740,N_2,N_1108);
xor U2741 (N_2741,N_1731,N_403);
nand U2742 (N_2742,N_152,N_2499);
or U2743 (N_2743,N_1453,N_252);
and U2744 (N_2744,N_1758,N_546);
or U2745 (N_2745,N_974,N_1457);
and U2746 (N_2746,N_1904,N_742);
xnor U2747 (N_2747,N_1019,N_1056);
nor U2748 (N_2748,N_2130,N_650);
nand U2749 (N_2749,N_59,N_1334);
or U2750 (N_2750,N_1102,N_1947);
or U2751 (N_2751,N_1478,N_2473);
nor U2752 (N_2752,N_1028,N_831);
nand U2753 (N_2753,N_410,N_1890);
and U2754 (N_2754,N_13,N_1997);
xnor U2755 (N_2755,N_384,N_2422);
or U2756 (N_2756,N_1607,N_1153);
xor U2757 (N_2757,N_687,N_1417);
nand U2758 (N_2758,N_303,N_1081);
xor U2759 (N_2759,N_2350,N_1551);
nand U2760 (N_2760,N_1962,N_1603);
or U2761 (N_2761,N_657,N_1409);
nor U2762 (N_2762,N_291,N_75);
nor U2763 (N_2763,N_1181,N_308);
and U2764 (N_2764,N_748,N_415);
and U2765 (N_2765,N_1390,N_2295);
or U2766 (N_2766,N_1351,N_423);
and U2767 (N_2767,N_763,N_652);
nor U2768 (N_2768,N_1830,N_991);
xnor U2769 (N_2769,N_2247,N_2318);
xor U2770 (N_2770,N_953,N_2389);
nand U2771 (N_2771,N_1281,N_1934);
nand U2772 (N_2772,N_2178,N_1485);
nand U2773 (N_2773,N_1707,N_196);
and U2774 (N_2774,N_1210,N_189);
nand U2775 (N_2775,N_510,N_22);
xnor U2776 (N_2776,N_1078,N_2155);
nor U2777 (N_2777,N_2018,N_1990);
nor U2778 (N_2778,N_182,N_980);
nand U2779 (N_2779,N_1817,N_1172);
nor U2780 (N_2780,N_2413,N_478);
nor U2781 (N_2781,N_1389,N_1157);
and U2782 (N_2782,N_1798,N_192);
or U2783 (N_2783,N_524,N_2315);
or U2784 (N_2784,N_705,N_2064);
nand U2785 (N_2785,N_1680,N_1398);
xnor U2786 (N_2786,N_323,N_1625);
nand U2787 (N_2787,N_1974,N_1305);
xnor U2788 (N_2788,N_1063,N_784);
and U2789 (N_2789,N_2020,N_2308);
nor U2790 (N_2790,N_1586,N_364);
nand U2791 (N_2791,N_2189,N_1376);
nand U2792 (N_2792,N_2299,N_81);
or U2793 (N_2793,N_1893,N_331);
nor U2794 (N_2794,N_253,N_54);
nor U2795 (N_2795,N_1187,N_1946);
nor U2796 (N_2796,N_442,N_1794);
and U2797 (N_2797,N_1919,N_1341);
and U2798 (N_2798,N_649,N_1949);
and U2799 (N_2799,N_447,N_181);
nor U2800 (N_2800,N_460,N_262);
xnor U2801 (N_2801,N_307,N_2423);
or U2802 (N_2802,N_254,N_335);
or U2803 (N_2803,N_2050,N_734);
and U2804 (N_2804,N_2073,N_2152);
xor U2805 (N_2805,N_983,N_242);
nor U2806 (N_2806,N_205,N_2476);
or U2807 (N_2807,N_2201,N_1900);
and U2808 (N_2808,N_2338,N_428);
and U2809 (N_2809,N_667,N_258);
xnor U2810 (N_2810,N_982,N_1605);
xnor U2811 (N_2811,N_703,N_1350);
or U2812 (N_2812,N_222,N_50);
or U2813 (N_2813,N_2353,N_1249);
nand U2814 (N_2814,N_901,N_795);
or U2815 (N_2815,N_1199,N_1660);
or U2816 (N_2816,N_631,N_671);
xnor U2817 (N_2817,N_1023,N_87);
and U2818 (N_2818,N_854,N_527);
or U2819 (N_2819,N_320,N_2070);
nand U2820 (N_2820,N_1748,N_1922);
and U2821 (N_2821,N_1442,N_2306);
xor U2822 (N_2822,N_1510,N_867);
or U2823 (N_2823,N_1739,N_526);
nand U2824 (N_2824,N_325,N_1858);
and U2825 (N_2825,N_1550,N_565);
xor U2826 (N_2826,N_1247,N_1511);
nand U2827 (N_2827,N_382,N_1960);
or U2828 (N_2828,N_1009,N_1717);
or U2829 (N_2829,N_747,N_1936);
or U2830 (N_2830,N_1290,N_2273);
nand U2831 (N_2831,N_2171,N_2356);
or U2832 (N_2832,N_1119,N_2230);
xor U2833 (N_2833,N_488,N_2013);
nand U2834 (N_2834,N_1726,N_1523);
xor U2835 (N_2835,N_2303,N_2099);
and U2836 (N_2836,N_704,N_1141);
nor U2837 (N_2837,N_3,N_1736);
and U2838 (N_2838,N_1451,N_2370);
and U2839 (N_2839,N_159,N_1253);
xor U2840 (N_2840,N_1274,N_1612);
nand U2841 (N_2841,N_973,N_1036);
or U2842 (N_2842,N_1705,N_1825);
and U2843 (N_2843,N_497,N_2444);
or U2844 (N_2844,N_759,N_1885);
nor U2845 (N_2845,N_111,N_2376);
or U2846 (N_2846,N_167,N_1147);
xor U2847 (N_2847,N_176,N_229);
nor U2848 (N_2848,N_1649,N_1661);
nand U2849 (N_2849,N_1087,N_155);
nand U2850 (N_2850,N_1870,N_82);
or U2851 (N_2851,N_1782,N_1046);
or U2852 (N_2852,N_1178,N_619);
nor U2853 (N_2853,N_1866,N_97);
nand U2854 (N_2854,N_1801,N_962);
and U2855 (N_2855,N_2485,N_2362);
nor U2856 (N_2856,N_924,N_684);
nor U2857 (N_2857,N_1396,N_2160);
nor U2858 (N_2858,N_695,N_2463);
xnor U2859 (N_2859,N_1780,N_866);
and U2860 (N_2860,N_465,N_1160);
nand U2861 (N_2861,N_368,N_766);
and U2862 (N_2862,N_913,N_1737);
or U2863 (N_2863,N_1012,N_2493);
nand U2864 (N_2864,N_1034,N_2400);
nor U2865 (N_2865,N_668,N_1061);
nand U2866 (N_2866,N_937,N_2170);
and U2867 (N_2867,N_1923,N_945);
nor U2868 (N_2868,N_414,N_1575);
and U2869 (N_2869,N_1256,N_485);
and U2870 (N_2870,N_1810,N_1301);
nand U2871 (N_2871,N_1894,N_2326);
or U2872 (N_2872,N_2451,N_464);
or U2873 (N_2873,N_1925,N_1225);
or U2874 (N_2874,N_1668,N_892);
nor U2875 (N_2875,N_2106,N_700);
xnor U2876 (N_2876,N_480,N_1594);
xnor U2877 (N_2877,N_874,N_860);
and U2878 (N_2878,N_2208,N_1156);
xnor U2879 (N_2879,N_1742,N_990);
nor U2880 (N_2880,N_827,N_51);
nand U2881 (N_2881,N_1878,N_1706);
nand U2882 (N_2882,N_556,N_2486);
and U2883 (N_2883,N_1840,N_408);
nand U2884 (N_2884,N_446,N_2236);
nand U2885 (N_2885,N_2339,N_531);
nand U2886 (N_2886,N_691,N_2000);
nand U2887 (N_2887,N_1820,N_1161);
or U2888 (N_2888,N_2191,N_1529);
and U2889 (N_2889,N_2115,N_1560);
or U2890 (N_2890,N_2360,N_956);
or U2891 (N_2891,N_2175,N_2477);
nand U2892 (N_2892,N_1113,N_1781);
and U2893 (N_2893,N_1057,N_1610);
nand U2894 (N_2894,N_237,N_1861);
or U2895 (N_2895,N_1482,N_728);
xor U2896 (N_2896,N_999,N_632);
xnor U2897 (N_2897,N_1837,N_1502);
or U2898 (N_2898,N_2457,N_1285);
xor U2899 (N_2899,N_1924,N_849);
nor U2900 (N_2900,N_327,N_1266);
or U2901 (N_2901,N_1168,N_851);
xnor U2902 (N_2902,N_622,N_1536);
or U2903 (N_2903,N_490,N_2196);
nand U2904 (N_2904,N_533,N_1615);
and U2905 (N_2905,N_1039,N_2067);
and U2906 (N_2906,N_788,N_88);
and U2907 (N_2907,N_345,N_146);
nor U2908 (N_2908,N_2128,N_1020);
nor U2909 (N_2909,N_2317,N_2482);
and U2910 (N_2910,N_698,N_603);
nand U2911 (N_2911,N_1914,N_394);
and U2912 (N_2912,N_1743,N_1884);
xnor U2913 (N_2913,N_1110,N_570);
xnor U2914 (N_2914,N_1778,N_21);
or U2915 (N_2915,N_706,N_1655);
nand U2916 (N_2916,N_2351,N_1226);
nor U2917 (N_2917,N_322,N_2197);
nand U2918 (N_2918,N_231,N_418);
nand U2919 (N_2919,N_613,N_1850);
nand U2920 (N_2920,N_1525,N_492);
nor U2921 (N_2921,N_1616,N_722);
and U2922 (N_2922,N_1066,N_44);
nor U2923 (N_2923,N_1163,N_1540);
nor U2924 (N_2924,N_1315,N_1280);
and U2925 (N_2925,N_942,N_2388);
xor U2926 (N_2926,N_1503,N_1848);
nor U2927 (N_2927,N_1273,N_1254);
nand U2928 (N_2928,N_1385,N_642);
nand U2929 (N_2929,N_42,N_1173);
and U2930 (N_2930,N_278,N_1688);
nor U2931 (N_2931,N_689,N_2005);
nor U2932 (N_2932,N_412,N_338);
or U2933 (N_2933,N_69,N_121);
and U2934 (N_2934,N_65,N_245);
and U2935 (N_2935,N_311,N_1427);
or U2936 (N_2936,N_511,N_234);
nor U2937 (N_2937,N_525,N_2479);
nor U2938 (N_2938,N_2355,N_1115);
xnor U2939 (N_2939,N_685,N_2417);
or U2940 (N_2940,N_166,N_1985);
or U2941 (N_2941,N_1004,N_964);
xnor U2942 (N_2942,N_32,N_1321);
or U2943 (N_2943,N_845,N_2405);
nor U2944 (N_2944,N_777,N_2321);
and U2945 (N_2945,N_1725,N_1418);
or U2946 (N_2946,N_1899,N_839);
nor U2947 (N_2947,N_842,N_2432);
nor U2948 (N_2948,N_2004,N_1322);
xor U2949 (N_2949,N_2345,N_72);
or U2950 (N_2950,N_678,N_482);
xor U2951 (N_2951,N_2031,N_1309);
and U2952 (N_2952,N_1961,N_431);
nor U2953 (N_2953,N_808,N_220);
nor U2954 (N_2954,N_1667,N_2383);
and U2955 (N_2955,N_745,N_586);
xnor U2956 (N_2956,N_838,N_204);
and U2957 (N_2957,N_2157,N_1003);
nor U2958 (N_2958,N_2381,N_829);
nor U2959 (N_2959,N_499,N_761);
nand U2960 (N_2960,N_841,N_2264);
and U2961 (N_2961,N_2077,N_372);
and U2962 (N_2962,N_716,N_1463);
and U2963 (N_2963,N_1898,N_2074);
xnor U2964 (N_2964,N_1754,N_970);
nand U2965 (N_2965,N_356,N_2436);
xor U2966 (N_2966,N_2421,N_36);
and U2967 (N_2967,N_1563,N_989);
xor U2968 (N_2968,N_1815,N_1364);
xnor U2969 (N_2969,N_1552,N_207);
or U2970 (N_2970,N_434,N_1133);
nor U2971 (N_2971,N_627,N_388);
xnor U2972 (N_2972,N_1086,N_190);
and U2973 (N_2973,N_1871,N_2135);
nand U2974 (N_2974,N_180,N_1345);
xor U2975 (N_2975,N_2410,N_163);
or U2976 (N_2976,N_1996,N_127);
nor U2977 (N_2977,N_41,N_1055);
and U2978 (N_2978,N_2098,N_2023);
xnor U2979 (N_2979,N_1347,N_540);
and U2980 (N_2980,N_389,N_302);
and U2981 (N_2981,N_1864,N_946);
xor U2982 (N_2982,N_1520,N_1790);
nand U2983 (N_2983,N_1105,N_1413);
and U2984 (N_2984,N_1905,N_56);
or U2985 (N_2985,N_199,N_2136);
and U2986 (N_2986,N_486,N_1514);
xor U2987 (N_2987,N_1287,N_1522);
and U2988 (N_2988,N_1641,N_810);
and U2989 (N_2989,N_1216,N_339);
or U2990 (N_2990,N_1772,N_1681);
nor U2991 (N_2991,N_805,N_2091);
and U2992 (N_2992,N_743,N_2259);
nor U2993 (N_2993,N_1565,N_2274);
nand U2994 (N_2994,N_968,N_1860);
nor U2995 (N_2995,N_2209,N_315);
xnor U2996 (N_2996,N_992,N_2437);
xnor U2997 (N_2997,N_214,N_1531);
nor U2998 (N_2998,N_547,N_2184);
xor U2999 (N_2999,N_441,N_1944);
or U3000 (N_3000,N_1466,N_453);
xnor U3001 (N_3001,N_2104,N_1461);
nand U3002 (N_3002,N_2471,N_202);
and U3003 (N_3003,N_2341,N_1411);
nor U3004 (N_3004,N_2472,N_285);
nand U3005 (N_3005,N_1269,N_1868);
nor U3006 (N_3006,N_2285,N_236);
xnor U3007 (N_3007,N_618,N_1094);
nor U3008 (N_3008,N_2165,N_1496);
xnor U3009 (N_3009,N_1303,N_305);
or U3010 (N_3010,N_1030,N_7);
nand U3011 (N_3011,N_104,N_1675);
or U3012 (N_3012,N_1292,N_2495);
nand U3013 (N_3013,N_1795,N_1083);
and U3014 (N_3014,N_2367,N_2229);
nor U3015 (N_3015,N_2036,N_1404);
and U3016 (N_3016,N_1064,N_2340);
nor U3017 (N_3017,N_1098,N_718);
xor U3018 (N_3018,N_2222,N_280);
or U3019 (N_3019,N_1263,N_1261);
xor U3020 (N_3020,N_1175,N_1508);
and U3021 (N_3021,N_616,N_1733);
xnor U3022 (N_3022,N_1604,N_1784);
xnor U3023 (N_3023,N_758,N_981);
nand U3024 (N_3024,N_2120,N_35);
xor U3025 (N_3025,N_93,N_1487);
nand U3026 (N_3026,N_96,N_2192);
and U3027 (N_3027,N_636,N_265);
and U3028 (N_3028,N_961,N_1397);
and U3029 (N_3029,N_1991,N_741);
and U3030 (N_3030,N_512,N_1037);
and U3031 (N_3031,N_644,N_2458);
and U3032 (N_3032,N_1010,N_669);
nor U3033 (N_3033,N_730,N_2490);
nor U3034 (N_3034,N_1809,N_2252);
or U3035 (N_3035,N_1252,N_2119);
nand U3036 (N_3036,N_1001,N_314);
nand U3037 (N_3037,N_1521,N_1260);
xnor U3038 (N_3038,N_1116,N_407);
and U3039 (N_3039,N_769,N_1814);
xnor U3040 (N_3040,N_1464,N_274);
or U3041 (N_3041,N_530,N_131);
xnor U3042 (N_3042,N_1130,N_1446);
nor U3043 (N_3043,N_930,N_919);
xnor U3044 (N_3044,N_2231,N_2491);
nor U3045 (N_3045,N_2281,N_333);
or U3046 (N_3046,N_1035,N_2078);
xor U3047 (N_3047,N_633,N_886);
or U3048 (N_3048,N_1554,N_837);
nor U3049 (N_3049,N_150,N_23);
nand U3050 (N_3050,N_1355,N_168);
or U3051 (N_3051,N_177,N_452);
xor U3052 (N_3052,N_1126,N_1473);
nor U3053 (N_3053,N_471,N_246);
xnor U3054 (N_3054,N_1403,N_1392);
nor U3055 (N_3055,N_1195,N_1419);
nand U3056 (N_3056,N_2253,N_1902);
nor U3057 (N_3057,N_954,N_2335);
and U3058 (N_3058,N_889,N_395);
xnor U3059 (N_3059,N_1843,N_1728);
xor U3060 (N_3060,N_1672,N_1691);
or U3061 (N_3061,N_2088,N_2054);
or U3062 (N_3062,N_1268,N_939);
xnor U3063 (N_3063,N_1114,N_417);
nor U3064 (N_3064,N_2035,N_1244);
and U3065 (N_3065,N_2483,N_2478);
and U3066 (N_3066,N_2439,N_605);
and U3067 (N_3067,N_1539,N_1771);
xnor U3068 (N_3068,N_95,N_1959);
and U3069 (N_3069,N_2411,N_2409);
nor U3070 (N_3070,N_1755,N_623);
nor U3071 (N_3071,N_1214,N_1399);
xor U3072 (N_3072,N_1635,N_52);
xor U3073 (N_3073,N_91,N_224);
or U3074 (N_3074,N_1792,N_1765);
xor U3075 (N_3075,N_296,N_268);
nor U3076 (N_3076,N_674,N_135);
xnor U3077 (N_3077,N_1154,N_226);
or U3078 (N_3078,N_1724,N_967);
xnor U3079 (N_3079,N_299,N_2042);
nand U3080 (N_3080,N_513,N_1449);
xnor U3081 (N_3081,N_1103,N_1679);
and U3082 (N_3082,N_1400,N_811);
nor U3083 (N_3083,N_2043,N_1769);
nor U3084 (N_3084,N_1000,N_66);
xor U3085 (N_3085,N_393,N_2484);
nor U3086 (N_3086,N_1369,N_1171);
nor U3087 (N_3087,N_986,N_391);
xor U3088 (N_3088,N_49,N_2100);
xor U3089 (N_3089,N_108,N_1242);
and U3090 (N_3090,N_348,N_940);
or U3091 (N_3091,N_1874,N_1598);
or U3092 (N_3092,N_749,N_592);
and U3093 (N_3093,N_371,N_916);
nand U3094 (N_3094,N_2199,N_877);
and U3095 (N_3095,N_1143,N_321);
xor U3096 (N_3096,N_295,N_1721);
and U3097 (N_3097,N_1658,N_1186);
nand U3098 (N_3098,N_2014,N_157);
xor U3099 (N_3099,N_1546,N_2137);
nand U3100 (N_3100,N_198,N_597);
or U3101 (N_3101,N_1981,N_1104);
nand U3102 (N_3102,N_1454,N_2434);
nor U3103 (N_3103,N_132,N_2314);
nand U3104 (N_3104,N_2246,N_1971);
nand U3105 (N_3105,N_581,N_103);
xor U3106 (N_3106,N_2210,N_1913);
or U3107 (N_3107,N_1223,N_1007);
xnor U3108 (N_3108,N_235,N_1584);
xnor U3109 (N_3109,N_928,N_1697);
xnor U3110 (N_3110,N_1215,N_2249);
xor U3111 (N_3111,N_1386,N_2057);
and U3112 (N_3112,N_1951,N_260);
xor U3113 (N_3113,N_882,N_1787);
xor U3114 (N_3114,N_872,N_2218);
xnor U3115 (N_3115,N_587,N_1783);
xnor U3116 (N_3116,N_1368,N_2205);
or U3117 (N_3117,N_1678,N_1203);
nor U3118 (N_3118,N_529,N_938);
and U3119 (N_3119,N_376,N_473);
nor U3120 (N_3120,N_871,N_267);
and U3121 (N_3121,N_1185,N_772);
xnor U3122 (N_3122,N_1734,N_1646);
nor U3123 (N_3123,N_1500,N_2089);
and U3124 (N_3124,N_402,N_1807);
or U3125 (N_3125,N_495,N_2217);
nand U3126 (N_3126,N_76,N_1232);
xor U3127 (N_3127,N_624,N_2174);
nand U3128 (N_3128,N_2464,N_2122);
xnor U3129 (N_3129,N_1626,N_1167);
and U3130 (N_3130,N_1220,N_552);
nor U3131 (N_3131,N_309,N_1448);
or U3132 (N_3132,N_2390,N_944);
and U3133 (N_3133,N_1690,N_390);
xnor U3134 (N_3134,N_675,N_737);
nor U3135 (N_3135,N_2212,N_1384);
and U3136 (N_3136,N_864,N_1093);
xnor U3137 (N_3137,N_2056,N_910);
nor U3138 (N_3138,N_648,N_1005);
or U3139 (N_3139,N_1694,N_2465);
and U3140 (N_3140,N_2213,N_712);
and U3141 (N_3141,N_116,N_1278);
nand U3142 (N_3142,N_1597,N_1177);
and U3143 (N_3143,N_398,N_1683);
nor U3144 (N_3144,N_2040,N_1025);
or U3145 (N_3145,N_1372,N_1084);
xor U3146 (N_3146,N_380,N_2207);
nand U3147 (N_3147,N_651,N_817);
nor U3148 (N_3148,N_2266,N_1993);
or U3149 (N_3149,N_426,N_109);
or U3150 (N_3150,N_1797,N_149);
nor U3151 (N_3151,N_459,N_424);
nor U3152 (N_3152,N_1217,N_114);
nor U3153 (N_3153,N_1300,N_148);
and U3154 (N_3154,N_161,N_1198);
nor U3155 (N_3155,N_266,N_1665);
xor U3156 (N_3156,N_891,N_2268);
and U3157 (N_3157,N_2291,N_1053);
nand U3158 (N_3158,N_1474,N_1908);
nor U3159 (N_3159,N_1136,N_169);
nor U3160 (N_3160,N_2480,N_993);
nor U3161 (N_3161,N_1027,N_470);
nor U3162 (N_3162,N_1710,N_1880);
nor U3163 (N_3163,N_582,N_726);
xnor U3164 (N_3164,N_1467,N_861);
xnor U3165 (N_3165,N_1191,N_1712);
xnor U3166 (N_3166,N_626,N_1954);
or U3167 (N_3167,N_1041,N_2133);
and U3168 (N_3168,N_568,N_1939);
xnor U3169 (N_3169,N_2456,N_1555);
or U3170 (N_3170,N_1915,N_401);
nor U3171 (N_3171,N_1382,N_593);
xnor U3172 (N_3172,N_2025,N_425);
and U3173 (N_3173,N_379,N_814);
xor U3174 (N_3174,N_683,N_2221);
and U3175 (N_3175,N_19,N_1907);
or U3176 (N_3176,N_1124,N_574);
nand U3177 (N_3177,N_178,N_1085);
xor U3178 (N_3178,N_1854,N_2187);
xnor U3179 (N_3179,N_213,N_1077);
and U3180 (N_3180,N_102,N_1455);
xnor U3181 (N_3181,N_1090,N_1970);
and U3182 (N_3182,N_2125,N_64);
nand U3183 (N_3183,N_915,N_1556);
nor U3184 (N_3184,N_2240,N_1340);
and U3185 (N_3185,N_416,N_18);
nor U3186 (N_3186,N_2301,N_2219);
nor U3187 (N_3187,N_1632,N_1440);
and U3188 (N_3188,N_489,N_2257);
and U3189 (N_3189,N_1118,N_2244);
nand U3190 (N_3190,N_1459,N_39);
nor U3191 (N_3191,N_185,N_154);
nand U3192 (N_3192,N_1238,N_2323);
and U3193 (N_3193,N_1408,N_1768);
nand U3194 (N_3194,N_106,N_80);
nand U3195 (N_3195,N_219,N_1760);
or U3196 (N_3196,N_878,N_2272);
xor U3197 (N_3197,N_209,N_171);
or U3198 (N_3198,N_1091,N_1193);
and U3199 (N_3199,N_200,N_476);
xor U3200 (N_3200,N_536,N_1158);
nor U3201 (N_3201,N_666,N_1180);
xor U3202 (N_3202,N_535,N_1362);
nand U3203 (N_3203,N_1270,N_1518);
nand U3204 (N_3204,N_1882,N_544);
xnor U3205 (N_3205,N_563,N_1766);
and U3206 (N_3206,N_2286,N_1813);
or U3207 (N_3207,N_413,N_1654);
or U3208 (N_3208,N_2195,N_1353);
nand U3209 (N_3209,N_351,N_1841);
or U3210 (N_3210,N_1471,N_78);
and U3211 (N_3211,N_61,N_550);
and U3212 (N_3212,N_1746,N_1042);
and U3213 (N_3213,N_959,N_775);
and U3214 (N_3214,N_641,N_1138);
or U3215 (N_3215,N_1770,N_1684);
nor U3216 (N_3216,N_1891,N_1692);
xor U3217 (N_3217,N_1933,N_1507);
xor U3218 (N_3218,N_551,N_2198);
xnor U3219 (N_3219,N_1585,N_249);
and U3220 (N_3220,N_1492,N_925);
xor U3221 (N_3221,N_865,N_31);
nor U3222 (N_3222,N_191,N_1832);
xnor U3223 (N_3223,N_868,N_2233);
nand U3224 (N_3224,N_474,N_261);
nor U3225 (N_3225,N_1611,N_1773);
xnor U3226 (N_3226,N_170,N_952);
nand U3227 (N_3227,N_2332,N_569);
xnor U3228 (N_3228,N_1159,N_383);
or U3229 (N_3229,N_1821,N_1129);
nor U3230 (N_3230,N_796,N_1258);
nand U3231 (N_3231,N_363,N_1076);
or U3232 (N_3232,N_2371,N_126);
xnor U3233 (N_3233,N_670,N_100);
nand U3234 (N_3234,N_1509,N_332);
nand U3235 (N_3235,N_247,N_2194);
and U3236 (N_3236,N_887,N_1206);
and U3237 (N_3237,N_2331,N_1614);
nand U3238 (N_3238,N_1257,N_894);
and U3239 (N_3239,N_542,N_2289);
xor U3240 (N_3240,N_2248,N_585);
or U3241 (N_3241,N_870,N_201);
nand U3242 (N_3242,N_682,N_1829);
nand U3243 (N_3243,N_1965,N_328);
or U3244 (N_3244,N_1054,N_1388);
or U3245 (N_3245,N_451,N_1235);
and U3246 (N_3246,N_732,N_2459);
nor U3247 (N_3247,N_1578,N_600);
nor U3248 (N_3248,N_251,N_290);
and U3249 (N_3249,N_1800,N_2271);
and U3250 (N_3250,N_1530,N_779);
nand U3251 (N_3251,N_1255,N_677);
nor U3252 (N_3252,N_481,N_1189);
or U3253 (N_3253,N_289,N_57);
nand U3254 (N_3254,N_377,N_2095);
or U3255 (N_3255,N_1380,N_2425);
nand U3256 (N_3256,N_589,N_2442);
nand U3257 (N_3257,N_2121,N_2072);
nand U3258 (N_3258,N_857,N_16);
or U3259 (N_3259,N_753,N_856);
and U3260 (N_3260,N_813,N_1548);
nand U3261 (N_3261,N_1117,N_2022);
nand U3262 (N_3262,N_2169,N_853);
nor U3263 (N_3263,N_2033,N_659);
nand U3264 (N_3264,N_1751,N_1701);
or U3265 (N_3265,N_978,N_1276);
nand U3266 (N_3266,N_158,N_755);
nor U3267 (N_3267,N_1425,N_1192);
nor U3268 (N_3268,N_1836,N_807);
xnor U3269 (N_3269,N_336,N_105);
or U3270 (N_3270,N_1735,N_370);
nor U3271 (N_3271,N_11,N_241);
xnor U3272 (N_3272,N_740,N_2460);
or U3273 (N_3273,N_2320,N_433);
and U3274 (N_3274,N_1693,N_508);
nor U3275 (N_3275,N_1774,N_720);
xnor U3276 (N_3276,N_1975,N_927);
nor U3277 (N_3277,N_396,N_1393);
and U3278 (N_3278,N_2065,N_1636);
nor U3279 (N_3279,N_1205,N_8);
or U3280 (N_3280,N_1534,N_375);
nand U3281 (N_3281,N_439,N_1246);
or U3282 (N_3282,N_381,N_313);
nor U3283 (N_3283,N_1132,N_786);
nor U3284 (N_3284,N_2261,N_1729);
nand U3285 (N_3285,N_1307,N_573);
xnor U3286 (N_3286,N_2001,N_2116);
or U3287 (N_3287,N_1065,N_1016);
nand U3288 (N_3288,N_935,N_427);
or U3289 (N_3289,N_55,N_2373);
nor U3290 (N_3290,N_1727,N_324);
xnor U3291 (N_3291,N_518,N_862);
xor U3292 (N_3292,N_2007,N_2010);
nand U3293 (N_3293,N_1137,N_70);
and U3294 (N_3294,N_421,N_1759);
nand U3295 (N_3295,N_193,N_2440);
or U3296 (N_3296,N_2140,N_2002);
or U3297 (N_3297,N_1897,N_2061);
and U3298 (N_3298,N_768,N_1483);
or U3299 (N_3299,N_1122,N_2032);
nor U3300 (N_3300,N_2364,N_2068);
and U3301 (N_3301,N_1653,N_561);
xnor U3302 (N_3302,N_27,N_645);
and U3303 (N_3303,N_1346,N_142);
and U3304 (N_3304,N_1435,N_1320);
or U3305 (N_3305,N_1602,N_430);
xor U3306 (N_3306,N_1075,N_1581);
and U3307 (N_3307,N_184,N_1842);
nor U3308 (N_3308,N_419,N_803);
nor U3309 (N_3309,N_217,N_948);
and U3310 (N_3310,N_1145,N_754);
nand U3311 (N_3311,N_931,N_263);
or U3312 (N_3312,N_2403,N_505);
and U3313 (N_3313,N_120,N_40);
nor U3314 (N_3314,N_1088,N_575);
or U3315 (N_3315,N_654,N_1976);
or U3316 (N_3316,N_463,N_2313);
nand U3317 (N_3317,N_300,N_2393);
nand U3318 (N_3318,N_1021,N_1595);
xor U3319 (N_3319,N_221,N_553);
nand U3320 (N_3320,N_1099,N_493);
or U3321 (N_3321,N_1014,N_310);
and U3322 (N_3322,N_965,N_830);
or U3323 (N_3323,N_1481,N_1824);
or U3324 (N_3324,N_1639,N_2038);
or U3325 (N_3325,N_2238,N_2082);
nor U3326 (N_3326,N_2112,N_634);
nor U3327 (N_3327,N_1377,N_902);
and U3328 (N_3328,N_89,N_1828);
nor U3329 (N_3329,N_776,N_1058);
and U3330 (N_3330,N_818,N_1183);
and U3331 (N_3331,N_1786,N_1089);
xnor U3332 (N_3332,N_2279,N_2096);
nor U3333 (N_3333,N_479,N_699);
and U3334 (N_3334,N_359,N_1050);
nor U3335 (N_3335,N_282,N_411);
xnor U3336 (N_3336,N_1197,N_90);
or U3337 (N_3337,N_2093,N_2276);
or U3338 (N_3338,N_1207,N_1468);
and U3339 (N_3339,N_1777,N_1275);
nor U3340 (N_3340,N_1470,N_923);
or U3341 (N_3341,N_1169,N_1202);
nor U3342 (N_3342,N_1648,N_374);
nand U3343 (N_3343,N_1271,N_2177);
or U3344 (N_3344,N_143,N_2076);
nor U3345 (N_3345,N_1851,N_2146);
xnor U3346 (N_3346,N_733,N_884);
xor U3347 (N_3347,N_68,N_292);
and U3348 (N_3348,N_1526,N_1541);
xor U3349 (N_3349,N_846,N_1872);
or U3350 (N_3350,N_1557,N_2441);
nand U3351 (N_3351,N_537,N_1184);
or U3352 (N_3352,N_298,N_2452);
nor U3353 (N_3353,N_2111,N_2164);
xnor U3354 (N_3354,N_197,N_2034);
xor U3355 (N_3355,N_373,N_1912);
nand U3356 (N_3356,N_1955,N_1869);
or U3357 (N_3357,N_1149,N_1229);
xnor U3358 (N_3358,N_46,N_2086);
and U3359 (N_3359,N_1977,N_1311);
nand U3360 (N_3360,N_1969,N_1038);
xor U3361 (N_3361,N_1652,N_2041);
xnor U3362 (N_3362,N_92,N_1406);
nand U3363 (N_3363,N_175,N_598);
or U3364 (N_3364,N_1006,N_2149);
or U3365 (N_3365,N_256,N_1477);
or U3366 (N_3366,N_1553,N_1008);
nand U3367 (N_3367,N_2297,N_498);
nor U3368 (N_3368,N_2144,N_138);
and U3369 (N_3369,N_767,N_399);
nand U3370 (N_3370,N_721,N_1490);
or U3371 (N_3371,N_1239,N_1151);
or U3372 (N_3372,N_1412,N_448);
and U3373 (N_3373,N_1566,N_1901);
or U3374 (N_3374,N_760,N_2309);
nand U3375 (N_3375,N_1123,N_1401);
or U3376 (N_3376,N_2466,N_2075);
nor U3377 (N_3377,N_780,N_815);
xor U3378 (N_3378,N_271,N_2132);
nor U3379 (N_3379,N_1802,N_816);
xnor U3380 (N_3380,N_782,N_1222);
nand U3381 (N_3381,N_2429,N_994);
nand U3382 (N_3382,N_1709,N_2084);
xnor U3383 (N_3383,N_1071,N_617);
xnor U3384 (N_3384,N_1018,N_2048);
nor U3385 (N_3385,N_2182,N_2430);
and U3386 (N_3386,N_2148,N_702);
or U3387 (N_3387,N_1017,N_1352);
nor U3388 (N_3388,N_1493,N_2172);
xnor U3389 (N_3389,N_2183,N_269);
nand U3390 (N_3390,N_1415,N_2241);
nand U3391 (N_3391,N_483,N_1984);
nand U3392 (N_3392,N_255,N_1785);
xnor U3393 (N_3393,N_500,N_6);
nand U3394 (N_3394,N_58,N_2069);
nor U3395 (N_3395,N_2087,N_1227);
nor U3396 (N_3396,N_2282,N_1356);
nand U3397 (N_3397,N_48,N_966);
and U3398 (N_3398,N_643,N_714);
and U3399 (N_3399,N_883,N_2103);
and U3400 (N_3400,N_2394,N_1131);
or U3401 (N_3401,N_828,N_457);
and U3402 (N_3402,N_1698,N_1799);
or U3403 (N_3403,N_1930,N_1647);
nand U3404 (N_3404,N_1179,N_1100);
nand U3405 (N_3405,N_577,N_1106);
or U3406 (N_3406,N_653,N_2030);
nand U3407 (N_3407,N_1544,N_1150);
nand U3408 (N_3408,N_1051,N_2497);
or U3409 (N_3409,N_1979,N_717);
nor U3410 (N_3410,N_960,N_1517);
nor U3411 (N_3411,N_1987,N_1849);
nand U3412 (N_3412,N_2190,N_279);
xnor U3413 (N_3413,N_1289,N_2265);
and U3414 (N_3414,N_1357,N_1847);
nand U3415 (N_3415,N_188,N_1803);
xnor U3416 (N_3416,N_1146,N_1928);
xnor U3417 (N_3417,N_228,N_1394);
xor U3418 (N_3418,N_2474,N_2270);
xnor U3419 (N_3419,N_1125,N_437);
xor U3420 (N_3420,N_475,N_1576);
or U3421 (N_3421,N_2019,N_1932);
xor U3422 (N_3422,N_1846,N_2404);
nand U3423 (N_3423,N_203,N_277);
or U3424 (N_3424,N_2037,N_2026);
or U3425 (N_3425,N_658,N_1671);
nor U3426 (N_3426,N_1669,N_1288);
xor U3427 (N_3427,N_1713,N_833);
nand U3428 (N_3428,N_1865,N_397);
nor U3429 (N_3429,N_1504,N_5);
xnor U3430 (N_3430,N_826,N_276);
nor U3431 (N_3431,N_2380,N_2176);
nor U3432 (N_3432,N_1835,N_809);
xnor U3433 (N_3433,N_141,N_1011);
nand U3434 (N_3434,N_506,N_1128);
or U3435 (N_3435,N_1873,N_1431);
nor U3436 (N_3436,N_955,N_1015);
xnor U3437 (N_3437,N_638,N_594);
nor U3438 (N_3438,N_890,N_1664);
and U3439 (N_3439,N_1445,N_1378);
xor U3440 (N_3440,N_1533,N_1243);
xor U3441 (N_3441,N_2206,N_1582);
nand U3442 (N_3442,N_275,N_225);
nor U3443 (N_3443,N_1574,N_1259);
or U3444 (N_3444,N_2224,N_369);
or U3445 (N_3445,N_244,N_1570);
nand U3446 (N_3446,N_852,N_2498);
xnor U3447 (N_3447,N_1022,N_1596);
or U3448 (N_3448,N_2453,N_301);
nor U3449 (N_3449,N_1720,N_2008);
and U3450 (N_3450,N_819,N_1941);
nor U3451 (N_3451,N_330,N_1999);
or U3452 (N_3452,N_270,N_914);
xnor U3453 (N_3453,N_1501,N_208);
and U3454 (N_3454,N_429,N_392);
nand U3455 (N_3455,N_1738,N_2052);
and U3456 (N_3456,N_2143,N_610);
nand U3457 (N_3457,N_554,N_2384);
xor U3458 (N_3458,N_686,N_165);
nand U3459 (N_3459,N_2469,N_449);
or U3460 (N_3460,N_1512,N_77);
xnor U3461 (N_3461,N_1013,N_521);
and U3462 (N_3462,N_2333,N_1366);
or U3463 (N_3463,N_1024,N_609);
or U3464 (N_3464,N_195,N_454);
xnor U3465 (N_3465,N_1070,N_725);
nor U3466 (N_3466,N_468,N_756);
or U3467 (N_3467,N_1443,N_1201);
nor U3468 (N_3468,N_1310,N_1732);
or U3469 (N_3469,N_2414,N_934);
nor U3470 (N_3470,N_1475,N_1219);
nand U3471 (N_3471,N_2328,N_1989);
and U3472 (N_3472,N_1839,N_501);
xnor U3473 (N_3473,N_2461,N_2455);
nor U3474 (N_3474,N_129,N_2118);
or U3475 (N_3475,N_211,N_1543);
and U3476 (N_3476,N_601,N_2168);
nor U3477 (N_3477,N_1234,N_660);
or U3478 (N_3478,N_595,N_1505);
or U3479 (N_3479,N_1542,N_1337);
nand U3480 (N_3480,N_690,N_567);
nor U3481 (N_3481,N_844,N_115);
nor U3482 (N_3482,N_455,N_503);
xor U3483 (N_3483,N_2150,N_545);
xor U3484 (N_3484,N_1313,N_2147);
xnor U3485 (N_3485,N_484,N_1213);
and U3486 (N_3486,N_951,N_466);
or U3487 (N_3487,N_1750,N_2186);
xnor U3488 (N_3488,N_2359,N_2258);
nor U3489 (N_3489,N_1231,N_898);
nand U3490 (N_3490,N_112,N_1170);
or U3491 (N_3491,N_719,N_494);
nand U3492 (N_3492,N_43,N_1831);
and U3493 (N_3493,N_1983,N_1107);
and U3494 (N_3494,N_2396,N_655);
nor U3495 (N_3495,N_1494,N_1826);
and U3496 (N_3496,N_387,N_1323);
and U3497 (N_3497,N_1344,N_243);
or U3498 (N_3498,N_2009,N_1702);
xor U3499 (N_3499,N_1617,N_306);
or U3500 (N_3500,N_825,N_2134);
xnor U3501 (N_3501,N_1906,N_2060);
xor U3502 (N_3502,N_1670,N_1549);
nor U3503 (N_3503,N_1067,N_1062);
nand U3504 (N_3504,N_984,N_1662);
nor U3505 (N_3505,N_835,N_549);
and U3506 (N_3506,N_1236,N_1963);
nand U3507 (N_3507,N_1499,N_899);
and U3508 (N_3508,N_2489,N_1073);
or U3509 (N_3509,N_1354,N_1465);
nor U3510 (N_3510,N_1600,N_1952);
nor U3511 (N_3511,N_711,N_1889);
or U3512 (N_3512,N_1228,N_365);
or U3513 (N_3513,N_692,N_1424);
and U3514 (N_3514,N_2117,N_2263);
xnor U3515 (N_3515,N_1140,N_2110);
or U3516 (N_3516,N_238,N_1740);
nor U3517 (N_3517,N_2055,N_12);
nor U3518 (N_3518,N_879,N_1571);
nor U3519 (N_3519,N_896,N_1410);
nand U3520 (N_3520,N_2322,N_2454);
nand U3521 (N_3521,N_210,N_688);
and U3522 (N_3522,N_1279,N_1296);
and U3523 (N_3523,N_2053,N_1405);
and U3524 (N_3524,N_2275,N_1621);
nand U3525 (N_3525,N_2378,N_1072);
nor U3526 (N_3526,N_2003,N_1583);
nand U3527 (N_3527,N_2092,N_1379);
and U3528 (N_3528,N_2395,N_1624);
or U3529 (N_3529,N_248,N_94);
nand U3530 (N_3530,N_1423,N_1513);
and U3531 (N_3531,N_975,N_1462);
nand U3532 (N_3532,N_541,N_179);
xnor U3533 (N_3533,N_661,N_2325);
xnor U3534 (N_3534,N_905,N_1144);
xnor U3535 (N_3535,N_1535,N_843);
nand U3536 (N_3536,N_1049,N_1561);
nand U3537 (N_3537,N_1948,N_1319);
nor U3538 (N_3538,N_1447,N_2494);
nor U3539 (N_3539,N_1095,N_287);
nor U3540 (N_3540,N_885,N_1895);
nor U3541 (N_3541,N_1251,N_1164);
xnor U3542 (N_3542,N_694,N_1711);
nand U3543 (N_3543,N_2049,N_1317);
or U3544 (N_3544,N_778,N_1484);
nand U3545 (N_3545,N_1958,N_1775);
or U3546 (N_3546,N_1293,N_1677);
and U3547 (N_3547,N_206,N_361);
xor U3548 (N_3548,N_334,N_2127);
nand U3549 (N_3549,N_118,N_1808);
nor U3550 (N_3550,N_1592,N_2167);
nor U3551 (N_3551,N_1569,N_918);
and U3552 (N_3552,N_783,N_977);
or U3553 (N_3553,N_696,N_1978);
nand U3554 (N_3554,N_1730,N_2161);
or U3555 (N_3555,N_1469,N_1308);
and U3556 (N_3556,N_38,N_477);
or U3557 (N_3557,N_2101,N_502);
nor U3558 (N_3558,N_662,N_1862);
xnor U3559 (N_3559,N_1982,N_801);
or U3560 (N_3560,N_943,N_1988);
nor U3561 (N_3561,N_1715,N_1182);
or U3562 (N_3562,N_2361,N_2420);
or U3563 (N_3563,N_1134,N_881);
and U3564 (N_3564,N_223,N_2237);
and U3565 (N_3565,N_1391,N_1165);
and U3566 (N_3566,N_1074,N_566);
nand U3567 (N_3567,N_611,N_2046);
and U3568 (N_3568,N_62,N_1877);
xor U3569 (N_3569,N_2407,N_757);
or U3570 (N_3570,N_2123,N_713);
xor U3571 (N_3571,N_1587,N_2227);
or U3572 (N_3572,N_1589,N_1788);
nand U3573 (N_3573,N_273,N_599);
xor U3574 (N_3574,N_352,N_341);
nor U3575 (N_3575,N_2398,N_1579);
nor U3576 (N_3576,N_2280,N_344);
nor U3577 (N_3577,N_329,N_1079);
or U3578 (N_3578,N_1479,N_2278);
nor U3579 (N_3579,N_1920,N_588);
and U3580 (N_3580,N_1863,N_2027);
or U3581 (N_3581,N_710,N_2080);
and U3582 (N_3582,N_762,N_174);
and U3583 (N_3583,N_2024,N_1927);
nand U3584 (N_3584,N_2336,N_1619);
nand U3585 (N_3585,N_560,N_53);
and U3586 (N_3586,N_1318,N_2113);
or U3587 (N_3587,N_1929,N_350);
nor U3588 (N_3588,N_312,N_445);
or U3589 (N_3589,N_823,N_29);
nand U3590 (N_3590,N_462,N_858);
nor U3591 (N_3591,N_1325,N_1867);
nand U3592 (N_3592,N_2324,N_1047);
or U3593 (N_3593,N_1986,N_1326);
or U3594 (N_3594,N_1528,N_2021);
nor U3595 (N_3595,N_2085,N_1972);
and U3596 (N_3596,N_1957,N_971);
nor U3597 (N_3597,N_491,N_997);
or U3598 (N_3598,N_663,N_30);
nand U3599 (N_3599,N_735,N_2011);
and U3600 (N_3600,N_1348,N_516);
xor U3601 (N_3601,N_1437,N_37);
and U3602 (N_3602,N_173,N_1240);
xor U3603 (N_3603,N_664,N_1623);
and U3604 (N_3604,N_628,N_1687);
xor U3605 (N_3605,N_404,N_548);
xnor U3606 (N_3606,N_751,N_2443);
and U3607 (N_3607,N_1387,N_1188);
nand U3608 (N_3608,N_2372,N_804);
nand U3609 (N_3609,N_1373,N_562);
nor U3610 (N_3610,N_1495,N_906);
xor U3611 (N_3611,N_2292,N_2126);
nand U3612 (N_3612,N_1852,N_1659);
and U3613 (N_3613,N_1221,N_2102);
nand U3614 (N_3614,N_83,N_1994);
nor U3615 (N_3615,N_230,N_2319);
or U3616 (N_3616,N_444,N_888);
xor U3617 (N_3617,N_2166,N_1816);
nand U3618 (N_3618,N_2203,N_1968);
or U3619 (N_3619,N_2418,N_2334);
nand U3620 (N_3620,N_186,N_2312);
xnor U3621 (N_3621,N_1224,N_2180);
nor U3622 (N_3622,N_1558,N_215);
nor U3623 (N_3623,N_958,N_785);
nor U3624 (N_3624,N_354,N_2173);
and U3625 (N_3625,N_1433,N_183);
xnor U3626 (N_3626,N_1524,N_1460);
or U3627 (N_3627,N_2470,N_1580);
or U3628 (N_3628,N_84,N_128);
and U3629 (N_3629,N_904,N_1416);
or U3630 (N_3630,N_1033,N_34);
or U3631 (N_3631,N_936,N_559);
and U3632 (N_3632,N_2316,N_1045);
nor U3633 (N_3633,N_1316,N_1752);
nand U3634 (N_3634,N_2269,N_28);
nand U3635 (N_3635,N_342,N_1590);
xor U3636 (N_3636,N_2158,N_1834);
or U3637 (N_3637,N_2226,N_2214);
or U3638 (N_3638,N_1938,N_606);
xnor U3639 (N_3639,N_1622,N_139);
or U3640 (N_3640,N_625,N_2401);
and U3641 (N_3641,N_724,N_2293);
and U3642 (N_3642,N_2427,N_792);
xnor U3643 (N_3643,N_2267,N_504);
xnor U3644 (N_3644,N_1176,N_2468);
nand U3645 (N_3645,N_929,N_963);
or U3646 (N_3646,N_840,N_1666);
xor U3647 (N_3647,N_272,N_438);
nand U3648 (N_3648,N_1940,N_604);
and U3649 (N_3649,N_2481,N_2402);
nand U3650 (N_3650,N_2277,N_2223);
xor U3651 (N_3651,N_1162,N_932);
or U3652 (N_3652,N_517,N_1349);
nand U3653 (N_3653,N_972,N_1294);
and U3654 (N_3654,N_1361,N_1741);
xnor U3655 (N_3655,N_2290,N_571);
nor U3656 (N_3656,N_1747,N_1673);
or U3657 (N_3657,N_863,N_1789);
nand U3658 (N_3658,N_608,N_1295);
nand U3659 (N_3659,N_1875,N_1638);
and U3660 (N_3660,N_2211,N_701);
and U3661 (N_3661,N_1031,N_1606);
nor U3662 (N_3662,N_528,N_2408);
nand U3663 (N_3663,N_697,N_1264);
nor U3664 (N_3664,N_1338,N_907);
xnor U3665 (N_3665,N_1395,N_1230);
and U3666 (N_3666,N_145,N_386);
xnor U3667 (N_3667,N_110,N_2256);
xnor U3668 (N_3668,N_1918,N_2357);
or U3669 (N_3669,N_1911,N_1434);
nor U3670 (N_3670,N_822,N_1248);
nand U3671 (N_3671,N_355,N_869);
nand U3672 (N_3672,N_2243,N_1233);
xnor U3673 (N_3673,N_850,N_621);
nand U3674 (N_3674,N_2051,N_1532);
xnor U3675 (N_3675,N_1282,N_1043);
xor U3676 (N_3676,N_47,N_2487);
xor U3677 (N_3677,N_1339,N_20);
and U3678 (N_3678,N_1208,N_596);
nor U3679 (N_3679,N_67,N_2337);
nor U3680 (N_3680,N_1656,N_920);
or U3681 (N_3681,N_1640,N_1342);
xor U3682 (N_3682,N_522,N_1757);
xor U3683 (N_3683,N_1059,N_346);
nor U3684 (N_3684,N_2131,N_4);
or U3685 (N_3685,N_1402,N_1029);
and U3686 (N_3686,N_515,N_2368);
xnor U3687 (N_3687,N_1811,N_1498);
nand U3688 (N_3688,N_1896,N_14);
nand U3689 (N_3689,N_507,N_353);
xor U3690 (N_3690,N_1827,N_33);
xor U3691 (N_3691,N_2347,N_1703);
nand U3692 (N_3692,N_1381,N_789);
nand U3693 (N_3693,N_1486,N_2375);
and U3694 (N_3694,N_1704,N_1302);
xnor U3695 (N_3695,N_908,N_487);
or U3696 (N_3696,N_949,N_1245);
or U3697 (N_3697,N_2448,N_2363);
or U3698 (N_3698,N_2343,N_420);
or U3699 (N_3699,N_630,N_1333);
xor U3700 (N_3700,N_122,N_802);
xnor U3701 (N_3701,N_1472,N_2412);
nand U3702 (N_3702,N_119,N_1139);
nand U3703 (N_3703,N_10,N_1286);
xnor U3704 (N_3704,N_1458,N_164);
xnor U3705 (N_3705,N_1644,N_834);
nor U3706 (N_3706,N_911,N_764);
nor U3707 (N_3707,N_2124,N_1152);
nor U3708 (N_3708,N_1628,N_232);
and U3709 (N_3709,N_1620,N_2385);
nand U3710 (N_3710,N_2329,N_665);
nor U3711 (N_3711,N_1764,N_1304);
and U3712 (N_3712,N_2304,N_1547);
or U3713 (N_3713,N_1480,N_1359);
or U3714 (N_3714,N_1608,N_2467);
or U3715 (N_3715,N_2284,N_1791);
nor U3716 (N_3716,N_450,N_1545);
xor U3717 (N_3717,N_1040,N_2251);
or U3718 (N_3718,N_194,N_979);
nor U3719 (N_3719,N_107,N_2200);
and U3720 (N_3720,N_1910,N_987);
or U3721 (N_3721,N_557,N_60);
xnor U3722 (N_3722,N_162,N_340);
xor U3723 (N_3723,N_1328,N_781);
and U3724 (N_3724,N_1718,N_1945);
nand U3725 (N_3725,N_1358,N_859);
nand U3726 (N_3726,N_1838,N_602);
nand U3727 (N_3727,N_257,N_1414);
xnor U3728 (N_3728,N_79,N_1762);
nor U3729 (N_3729,N_578,N_1749);
nand U3730 (N_3730,N_1438,N_564);
and U3731 (N_3731,N_794,N_1060);
or U3732 (N_3732,N_680,N_2245);
nand U3733 (N_3733,N_347,N_752);
nor U3734 (N_3734,N_1917,N_893);
xnor U3735 (N_3735,N_523,N_1026);
nor U3736 (N_3736,N_1796,N_1515);
nand U3737 (N_3737,N_233,N_1237);
xnor U3738 (N_3738,N_1637,N_773);
or U3739 (N_3739,N_1284,N_1343);
and U3740 (N_3740,N_1806,N_378);
nand U3741 (N_3741,N_2232,N_2298);
and U3742 (N_3742,N_790,N_1853);
nor U3743 (N_3743,N_1429,N_1980);
nand U3744 (N_3744,N_2141,N_1112);
nor U3745 (N_3745,N_1716,N_2094);
nand U3746 (N_3746,N_1779,N_1719);
and U3747 (N_3747,N_1101,N_259);
nor U3748 (N_3748,N_1903,N_1643);
and U3749 (N_3749,N_620,N_443);
and U3750 (N_3750,N_132,N_1471);
xor U3751 (N_3751,N_1977,N_2364);
nand U3752 (N_3752,N_1185,N_1500);
nand U3753 (N_3753,N_1848,N_541);
xor U3754 (N_3754,N_2189,N_1051);
or U3755 (N_3755,N_2403,N_909);
and U3756 (N_3756,N_2435,N_331);
nand U3757 (N_3757,N_1213,N_385);
nor U3758 (N_3758,N_2462,N_1217);
or U3759 (N_3759,N_273,N_2025);
or U3760 (N_3760,N_211,N_136);
nor U3761 (N_3761,N_2291,N_2156);
nor U3762 (N_3762,N_1332,N_1326);
and U3763 (N_3763,N_1051,N_2013);
or U3764 (N_3764,N_1246,N_2234);
and U3765 (N_3765,N_1764,N_1426);
nor U3766 (N_3766,N_86,N_164);
and U3767 (N_3767,N_606,N_119);
and U3768 (N_3768,N_1481,N_2209);
nand U3769 (N_3769,N_2406,N_181);
nor U3770 (N_3770,N_348,N_802);
nor U3771 (N_3771,N_1266,N_50);
xnor U3772 (N_3772,N_466,N_1798);
nand U3773 (N_3773,N_1620,N_718);
xnor U3774 (N_3774,N_730,N_426);
xnor U3775 (N_3775,N_2327,N_1185);
nor U3776 (N_3776,N_622,N_1410);
xnor U3777 (N_3777,N_1554,N_427);
and U3778 (N_3778,N_490,N_447);
and U3779 (N_3779,N_381,N_2373);
nor U3780 (N_3780,N_849,N_2182);
nor U3781 (N_3781,N_1090,N_685);
nand U3782 (N_3782,N_597,N_275);
nor U3783 (N_3783,N_851,N_519);
nor U3784 (N_3784,N_315,N_196);
nand U3785 (N_3785,N_1877,N_717);
and U3786 (N_3786,N_2034,N_1219);
and U3787 (N_3787,N_2475,N_1792);
or U3788 (N_3788,N_245,N_526);
or U3789 (N_3789,N_1230,N_2389);
or U3790 (N_3790,N_2148,N_85);
nor U3791 (N_3791,N_1921,N_2238);
and U3792 (N_3792,N_562,N_966);
and U3793 (N_3793,N_2427,N_1209);
nor U3794 (N_3794,N_1211,N_716);
nor U3795 (N_3795,N_2289,N_1545);
nand U3796 (N_3796,N_163,N_1200);
or U3797 (N_3797,N_2174,N_1010);
nand U3798 (N_3798,N_1217,N_1808);
and U3799 (N_3799,N_1817,N_229);
or U3800 (N_3800,N_487,N_2300);
and U3801 (N_3801,N_1361,N_531);
nor U3802 (N_3802,N_1072,N_1379);
nand U3803 (N_3803,N_2146,N_1815);
nand U3804 (N_3804,N_1789,N_1994);
nand U3805 (N_3805,N_1281,N_1200);
nand U3806 (N_3806,N_2443,N_789);
or U3807 (N_3807,N_454,N_1429);
nor U3808 (N_3808,N_74,N_1483);
and U3809 (N_3809,N_886,N_761);
nor U3810 (N_3810,N_413,N_1826);
nand U3811 (N_3811,N_2001,N_1549);
and U3812 (N_3812,N_2007,N_494);
xnor U3813 (N_3813,N_2350,N_1859);
nor U3814 (N_3814,N_2422,N_2362);
nand U3815 (N_3815,N_2072,N_1121);
and U3816 (N_3816,N_1305,N_2132);
xor U3817 (N_3817,N_975,N_311);
and U3818 (N_3818,N_1517,N_1174);
xor U3819 (N_3819,N_705,N_640);
and U3820 (N_3820,N_1933,N_668);
or U3821 (N_3821,N_1596,N_2212);
nand U3822 (N_3822,N_1108,N_48);
nand U3823 (N_3823,N_873,N_852);
xnor U3824 (N_3824,N_2487,N_994);
or U3825 (N_3825,N_1652,N_1387);
nand U3826 (N_3826,N_902,N_1212);
and U3827 (N_3827,N_2126,N_1770);
nand U3828 (N_3828,N_1489,N_880);
or U3829 (N_3829,N_1017,N_1614);
or U3830 (N_3830,N_201,N_1936);
or U3831 (N_3831,N_2080,N_105);
xor U3832 (N_3832,N_307,N_431);
or U3833 (N_3833,N_2060,N_2214);
nor U3834 (N_3834,N_204,N_2031);
and U3835 (N_3835,N_1883,N_1044);
or U3836 (N_3836,N_791,N_2415);
and U3837 (N_3837,N_2111,N_485);
and U3838 (N_3838,N_509,N_1579);
nor U3839 (N_3839,N_1826,N_148);
nand U3840 (N_3840,N_1311,N_2435);
nand U3841 (N_3841,N_921,N_2471);
nand U3842 (N_3842,N_1362,N_1496);
or U3843 (N_3843,N_1206,N_1576);
xor U3844 (N_3844,N_1208,N_1141);
nand U3845 (N_3845,N_1431,N_637);
xnor U3846 (N_3846,N_1082,N_1081);
or U3847 (N_3847,N_2185,N_1709);
and U3848 (N_3848,N_1770,N_612);
or U3849 (N_3849,N_98,N_1145);
nor U3850 (N_3850,N_2190,N_2225);
nand U3851 (N_3851,N_1889,N_655);
xnor U3852 (N_3852,N_2077,N_1667);
nor U3853 (N_3853,N_252,N_214);
xor U3854 (N_3854,N_1300,N_2419);
nor U3855 (N_3855,N_570,N_498);
or U3856 (N_3856,N_70,N_142);
xor U3857 (N_3857,N_1490,N_933);
or U3858 (N_3858,N_1273,N_952);
or U3859 (N_3859,N_1583,N_2353);
xor U3860 (N_3860,N_1135,N_187);
xor U3861 (N_3861,N_2020,N_2352);
nand U3862 (N_3862,N_2225,N_247);
or U3863 (N_3863,N_407,N_2242);
nor U3864 (N_3864,N_1209,N_1825);
or U3865 (N_3865,N_1634,N_2038);
xnor U3866 (N_3866,N_212,N_849);
nor U3867 (N_3867,N_2359,N_1757);
nor U3868 (N_3868,N_861,N_1797);
nor U3869 (N_3869,N_355,N_841);
or U3870 (N_3870,N_634,N_361);
nand U3871 (N_3871,N_1736,N_2353);
and U3872 (N_3872,N_1845,N_713);
nand U3873 (N_3873,N_1670,N_2189);
xnor U3874 (N_3874,N_2296,N_748);
xnor U3875 (N_3875,N_2140,N_336);
nand U3876 (N_3876,N_2280,N_1478);
and U3877 (N_3877,N_1522,N_360);
nor U3878 (N_3878,N_1793,N_953);
nand U3879 (N_3879,N_539,N_2013);
nor U3880 (N_3880,N_1290,N_1566);
or U3881 (N_3881,N_937,N_1359);
nor U3882 (N_3882,N_2072,N_327);
nor U3883 (N_3883,N_373,N_150);
xnor U3884 (N_3884,N_1788,N_2131);
nor U3885 (N_3885,N_1022,N_1803);
nor U3886 (N_3886,N_1032,N_1397);
nand U3887 (N_3887,N_675,N_903);
or U3888 (N_3888,N_2357,N_2108);
xor U3889 (N_3889,N_1225,N_736);
and U3890 (N_3890,N_2427,N_2268);
and U3891 (N_3891,N_2104,N_1339);
nor U3892 (N_3892,N_1298,N_1635);
or U3893 (N_3893,N_302,N_1254);
nor U3894 (N_3894,N_2163,N_2019);
nor U3895 (N_3895,N_425,N_1260);
xnor U3896 (N_3896,N_2270,N_120);
and U3897 (N_3897,N_1560,N_778);
nand U3898 (N_3898,N_2473,N_1354);
nor U3899 (N_3899,N_2131,N_2043);
nor U3900 (N_3900,N_196,N_1436);
and U3901 (N_3901,N_2009,N_567);
or U3902 (N_3902,N_1707,N_2403);
nor U3903 (N_3903,N_1308,N_50);
xnor U3904 (N_3904,N_1152,N_1615);
nand U3905 (N_3905,N_2402,N_1160);
or U3906 (N_3906,N_79,N_591);
and U3907 (N_3907,N_46,N_1404);
and U3908 (N_3908,N_137,N_404);
and U3909 (N_3909,N_737,N_1831);
nand U3910 (N_3910,N_691,N_1711);
xnor U3911 (N_3911,N_194,N_1119);
xnor U3912 (N_3912,N_572,N_2247);
nand U3913 (N_3913,N_453,N_1674);
nand U3914 (N_3914,N_66,N_1427);
nand U3915 (N_3915,N_164,N_1596);
xor U3916 (N_3916,N_1171,N_399);
xor U3917 (N_3917,N_1628,N_2238);
or U3918 (N_3918,N_1274,N_1243);
nor U3919 (N_3919,N_138,N_736);
or U3920 (N_3920,N_281,N_2141);
nor U3921 (N_3921,N_145,N_101);
nor U3922 (N_3922,N_2212,N_1824);
and U3923 (N_3923,N_1701,N_2051);
xnor U3924 (N_3924,N_1464,N_658);
nand U3925 (N_3925,N_2147,N_550);
nor U3926 (N_3926,N_1118,N_1139);
nor U3927 (N_3927,N_1899,N_2024);
nand U3928 (N_3928,N_2055,N_1176);
nor U3929 (N_3929,N_1375,N_477);
or U3930 (N_3930,N_2380,N_1764);
nand U3931 (N_3931,N_755,N_241);
xnor U3932 (N_3932,N_1178,N_843);
nand U3933 (N_3933,N_914,N_211);
nor U3934 (N_3934,N_77,N_804);
and U3935 (N_3935,N_2336,N_2007);
xor U3936 (N_3936,N_1223,N_2017);
nand U3937 (N_3937,N_499,N_2221);
nand U3938 (N_3938,N_1295,N_30);
and U3939 (N_3939,N_2416,N_1556);
xor U3940 (N_3940,N_2245,N_2447);
nor U3941 (N_3941,N_1772,N_214);
or U3942 (N_3942,N_971,N_753);
xnor U3943 (N_3943,N_1647,N_1093);
nand U3944 (N_3944,N_1677,N_957);
and U3945 (N_3945,N_312,N_1734);
xnor U3946 (N_3946,N_923,N_1235);
and U3947 (N_3947,N_2049,N_1928);
nor U3948 (N_3948,N_558,N_331);
and U3949 (N_3949,N_637,N_1370);
nand U3950 (N_3950,N_1637,N_1715);
xor U3951 (N_3951,N_2044,N_1125);
or U3952 (N_3952,N_236,N_2062);
and U3953 (N_3953,N_1394,N_2396);
xnor U3954 (N_3954,N_2057,N_2451);
and U3955 (N_3955,N_1618,N_626);
or U3956 (N_3956,N_508,N_444);
nand U3957 (N_3957,N_1841,N_558);
nor U3958 (N_3958,N_150,N_1717);
nor U3959 (N_3959,N_386,N_745);
nand U3960 (N_3960,N_1101,N_579);
and U3961 (N_3961,N_555,N_2498);
xnor U3962 (N_3962,N_1002,N_1200);
or U3963 (N_3963,N_2289,N_1062);
or U3964 (N_3964,N_1747,N_144);
nor U3965 (N_3965,N_2237,N_801);
nand U3966 (N_3966,N_461,N_1017);
or U3967 (N_3967,N_102,N_2187);
xor U3968 (N_3968,N_616,N_2375);
and U3969 (N_3969,N_1483,N_2197);
nand U3970 (N_3970,N_1080,N_2016);
xnor U3971 (N_3971,N_1304,N_496);
nor U3972 (N_3972,N_109,N_1557);
nand U3973 (N_3973,N_2324,N_1248);
or U3974 (N_3974,N_1538,N_1161);
or U3975 (N_3975,N_1566,N_928);
or U3976 (N_3976,N_1418,N_2061);
nor U3977 (N_3977,N_1697,N_2001);
nor U3978 (N_3978,N_300,N_1477);
xnor U3979 (N_3979,N_572,N_2387);
nor U3980 (N_3980,N_1050,N_2021);
nand U3981 (N_3981,N_954,N_2130);
nor U3982 (N_3982,N_1109,N_1405);
and U3983 (N_3983,N_1937,N_347);
xor U3984 (N_3984,N_1624,N_1855);
xnor U3985 (N_3985,N_1768,N_2106);
xor U3986 (N_3986,N_1773,N_366);
nand U3987 (N_3987,N_1827,N_304);
and U3988 (N_3988,N_2170,N_2359);
xnor U3989 (N_3989,N_2281,N_982);
nand U3990 (N_3990,N_2444,N_518);
xnor U3991 (N_3991,N_490,N_897);
xnor U3992 (N_3992,N_2340,N_1450);
nand U3993 (N_3993,N_2479,N_486);
xnor U3994 (N_3994,N_1996,N_732);
or U3995 (N_3995,N_715,N_756);
and U3996 (N_3996,N_1186,N_922);
or U3997 (N_3997,N_1978,N_273);
xnor U3998 (N_3998,N_1027,N_682);
nand U3999 (N_3999,N_1797,N_1107);
and U4000 (N_4000,N_75,N_467);
nor U4001 (N_4001,N_1416,N_2095);
xnor U4002 (N_4002,N_2137,N_1105);
and U4003 (N_4003,N_731,N_1120);
nand U4004 (N_4004,N_629,N_739);
nand U4005 (N_4005,N_1602,N_640);
xor U4006 (N_4006,N_1421,N_1796);
and U4007 (N_4007,N_1599,N_1747);
nand U4008 (N_4008,N_279,N_2157);
nor U4009 (N_4009,N_1743,N_1193);
nor U4010 (N_4010,N_1770,N_716);
nor U4011 (N_4011,N_1838,N_1659);
nand U4012 (N_4012,N_186,N_2152);
xor U4013 (N_4013,N_330,N_11);
xnor U4014 (N_4014,N_1353,N_165);
xor U4015 (N_4015,N_1805,N_79);
or U4016 (N_4016,N_586,N_1456);
or U4017 (N_4017,N_1675,N_1840);
nor U4018 (N_4018,N_1164,N_457);
and U4019 (N_4019,N_927,N_1233);
xor U4020 (N_4020,N_318,N_1809);
nor U4021 (N_4021,N_1587,N_729);
or U4022 (N_4022,N_2149,N_2164);
nor U4023 (N_4023,N_610,N_302);
xnor U4024 (N_4024,N_533,N_2325);
nand U4025 (N_4025,N_922,N_1286);
or U4026 (N_4026,N_204,N_1126);
and U4027 (N_4027,N_185,N_355);
nand U4028 (N_4028,N_157,N_2333);
xnor U4029 (N_4029,N_97,N_2010);
nand U4030 (N_4030,N_402,N_156);
nor U4031 (N_4031,N_939,N_1325);
and U4032 (N_4032,N_2125,N_1790);
or U4033 (N_4033,N_2060,N_2394);
nand U4034 (N_4034,N_1896,N_2273);
xor U4035 (N_4035,N_664,N_1863);
xor U4036 (N_4036,N_513,N_304);
or U4037 (N_4037,N_1239,N_1333);
and U4038 (N_4038,N_1767,N_1077);
and U4039 (N_4039,N_1575,N_2471);
and U4040 (N_4040,N_544,N_444);
or U4041 (N_4041,N_2321,N_69);
nand U4042 (N_4042,N_2424,N_1472);
xor U4043 (N_4043,N_1013,N_868);
or U4044 (N_4044,N_1397,N_1617);
nand U4045 (N_4045,N_932,N_711);
and U4046 (N_4046,N_541,N_2040);
nand U4047 (N_4047,N_2154,N_932);
nor U4048 (N_4048,N_2397,N_1701);
xnor U4049 (N_4049,N_1520,N_650);
nand U4050 (N_4050,N_1971,N_2385);
nand U4051 (N_4051,N_892,N_20);
nor U4052 (N_4052,N_1718,N_2339);
and U4053 (N_4053,N_2446,N_28);
nand U4054 (N_4054,N_293,N_1255);
xor U4055 (N_4055,N_1899,N_1256);
nor U4056 (N_4056,N_920,N_1907);
nand U4057 (N_4057,N_1904,N_604);
or U4058 (N_4058,N_2387,N_1018);
or U4059 (N_4059,N_485,N_1439);
or U4060 (N_4060,N_378,N_933);
xnor U4061 (N_4061,N_862,N_229);
nand U4062 (N_4062,N_1320,N_492);
xnor U4063 (N_4063,N_535,N_2088);
or U4064 (N_4064,N_2371,N_2331);
xnor U4065 (N_4065,N_222,N_23);
nand U4066 (N_4066,N_515,N_2314);
nand U4067 (N_4067,N_2138,N_968);
xor U4068 (N_4068,N_9,N_2231);
and U4069 (N_4069,N_1042,N_1001);
xor U4070 (N_4070,N_314,N_246);
and U4071 (N_4071,N_299,N_1322);
or U4072 (N_4072,N_1899,N_15);
nand U4073 (N_4073,N_1639,N_2401);
and U4074 (N_4074,N_35,N_1511);
nor U4075 (N_4075,N_933,N_355);
or U4076 (N_4076,N_1915,N_1439);
or U4077 (N_4077,N_1432,N_515);
and U4078 (N_4078,N_2363,N_1013);
or U4079 (N_4079,N_1936,N_144);
xor U4080 (N_4080,N_1130,N_1841);
or U4081 (N_4081,N_665,N_92);
and U4082 (N_4082,N_1204,N_1440);
and U4083 (N_4083,N_858,N_1361);
or U4084 (N_4084,N_1745,N_770);
xor U4085 (N_4085,N_362,N_178);
and U4086 (N_4086,N_1329,N_2235);
nor U4087 (N_4087,N_2471,N_2375);
xor U4088 (N_4088,N_2112,N_1193);
or U4089 (N_4089,N_85,N_2133);
and U4090 (N_4090,N_33,N_1798);
and U4091 (N_4091,N_2161,N_1274);
xnor U4092 (N_4092,N_1020,N_128);
and U4093 (N_4093,N_2351,N_2021);
and U4094 (N_4094,N_2113,N_2098);
nor U4095 (N_4095,N_804,N_1336);
nand U4096 (N_4096,N_812,N_28);
nand U4097 (N_4097,N_1123,N_1016);
xnor U4098 (N_4098,N_749,N_1989);
nand U4099 (N_4099,N_867,N_274);
and U4100 (N_4100,N_1876,N_1901);
or U4101 (N_4101,N_26,N_1723);
or U4102 (N_4102,N_835,N_42);
nor U4103 (N_4103,N_1877,N_224);
or U4104 (N_4104,N_407,N_2063);
and U4105 (N_4105,N_329,N_1282);
and U4106 (N_4106,N_619,N_1337);
and U4107 (N_4107,N_945,N_379);
xor U4108 (N_4108,N_1343,N_1458);
nor U4109 (N_4109,N_2409,N_1516);
and U4110 (N_4110,N_1944,N_677);
xor U4111 (N_4111,N_2034,N_1184);
and U4112 (N_4112,N_1395,N_1999);
or U4113 (N_4113,N_496,N_2043);
xnor U4114 (N_4114,N_217,N_1963);
nand U4115 (N_4115,N_2024,N_1941);
nand U4116 (N_4116,N_1403,N_766);
and U4117 (N_4117,N_220,N_1622);
or U4118 (N_4118,N_1576,N_2177);
and U4119 (N_4119,N_1134,N_1392);
nand U4120 (N_4120,N_870,N_2143);
xnor U4121 (N_4121,N_1326,N_1300);
or U4122 (N_4122,N_1468,N_2030);
and U4123 (N_4123,N_2144,N_905);
nor U4124 (N_4124,N_2397,N_1589);
nand U4125 (N_4125,N_482,N_1332);
nand U4126 (N_4126,N_2018,N_2342);
nor U4127 (N_4127,N_1768,N_1435);
and U4128 (N_4128,N_2486,N_1658);
xor U4129 (N_4129,N_2214,N_580);
and U4130 (N_4130,N_593,N_957);
xor U4131 (N_4131,N_2010,N_299);
nand U4132 (N_4132,N_489,N_945);
nand U4133 (N_4133,N_1356,N_698);
nand U4134 (N_4134,N_114,N_2099);
nor U4135 (N_4135,N_1169,N_502);
nand U4136 (N_4136,N_1070,N_1293);
or U4137 (N_4137,N_2373,N_1462);
nand U4138 (N_4138,N_2105,N_975);
and U4139 (N_4139,N_922,N_1823);
nand U4140 (N_4140,N_586,N_2402);
or U4141 (N_4141,N_2010,N_1149);
and U4142 (N_4142,N_2162,N_605);
or U4143 (N_4143,N_485,N_1192);
nor U4144 (N_4144,N_1333,N_1551);
nand U4145 (N_4145,N_1261,N_1710);
and U4146 (N_4146,N_1100,N_2425);
nand U4147 (N_4147,N_51,N_560);
and U4148 (N_4148,N_1864,N_1572);
nor U4149 (N_4149,N_1647,N_1890);
and U4150 (N_4150,N_767,N_2178);
nor U4151 (N_4151,N_2175,N_1766);
and U4152 (N_4152,N_1362,N_1358);
and U4153 (N_4153,N_569,N_384);
xnor U4154 (N_4154,N_1383,N_1082);
xnor U4155 (N_4155,N_2392,N_868);
xor U4156 (N_4156,N_2242,N_1595);
xnor U4157 (N_4157,N_1250,N_2453);
and U4158 (N_4158,N_603,N_1059);
and U4159 (N_4159,N_493,N_2395);
xnor U4160 (N_4160,N_1111,N_1113);
and U4161 (N_4161,N_913,N_346);
or U4162 (N_4162,N_1366,N_1686);
nor U4163 (N_4163,N_1897,N_1935);
or U4164 (N_4164,N_241,N_2388);
and U4165 (N_4165,N_697,N_755);
or U4166 (N_4166,N_1711,N_2257);
and U4167 (N_4167,N_1468,N_236);
nor U4168 (N_4168,N_1258,N_1481);
nand U4169 (N_4169,N_2483,N_770);
nand U4170 (N_4170,N_2384,N_826);
or U4171 (N_4171,N_1163,N_791);
nand U4172 (N_4172,N_924,N_2047);
or U4173 (N_4173,N_999,N_829);
nand U4174 (N_4174,N_1765,N_1277);
nand U4175 (N_4175,N_1318,N_1274);
and U4176 (N_4176,N_635,N_103);
xnor U4177 (N_4177,N_1689,N_843);
or U4178 (N_4178,N_1182,N_1499);
or U4179 (N_4179,N_2470,N_1752);
and U4180 (N_4180,N_2433,N_1984);
or U4181 (N_4181,N_2415,N_445);
or U4182 (N_4182,N_2486,N_878);
or U4183 (N_4183,N_2433,N_1168);
or U4184 (N_4184,N_2359,N_639);
nor U4185 (N_4185,N_2098,N_1807);
xnor U4186 (N_4186,N_1142,N_158);
or U4187 (N_4187,N_1288,N_2265);
and U4188 (N_4188,N_838,N_2241);
nor U4189 (N_4189,N_1756,N_1031);
xnor U4190 (N_4190,N_309,N_947);
xor U4191 (N_4191,N_2272,N_2122);
nor U4192 (N_4192,N_1430,N_1354);
nor U4193 (N_4193,N_92,N_1481);
nor U4194 (N_4194,N_2380,N_1669);
nor U4195 (N_4195,N_2104,N_646);
nor U4196 (N_4196,N_155,N_2133);
or U4197 (N_4197,N_444,N_1897);
xnor U4198 (N_4198,N_732,N_598);
nor U4199 (N_4199,N_1630,N_1044);
nand U4200 (N_4200,N_1900,N_277);
xnor U4201 (N_4201,N_728,N_1153);
or U4202 (N_4202,N_1226,N_1052);
xor U4203 (N_4203,N_1373,N_1872);
or U4204 (N_4204,N_1737,N_2280);
nor U4205 (N_4205,N_203,N_135);
nor U4206 (N_4206,N_1927,N_2245);
nand U4207 (N_4207,N_317,N_2063);
nor U4208 (N_4208,N_204,N_1241);
nor U4209 (N_4209,N_1783,N_253);
nand U4210 (N_4210,N_1363,N_1284);
and U4211 (N_4211,N_1664,N_1310);
and U4212 (N_4212,N_558,N_906);
or U4213 (N_4213,N_1707,N_1807);
or U4214 (N_4214,N_1952,N_2252);
and U4215 (N_4215,N_452,N_1248);
nor U4216 (N_4216,N_1549,N_54);
nor U4217 (N_4217,N_612,N_1876);
xor U4218 (N_4218,N_2094,N_59);
nand U4219 (N_4219,N_700,N_1477);
nor U4220 (N_4220,N_1178,N_34);
nand U4221 (N_4221,N_1625,N_1650);
xor U4222 (N_4222,N_1394,N_746);
xnor U4223 (N_4223,N_1794,N_1194);
nand U4224 (N_4224,N_2127,N_1918);
or U4225 (N_4225,N_2047,N_387);
and U4226 (N_4226,N_958,N_727);
nor U4227 (N_4227,N_484,N_341);
or U4228 (N_4228,N_1523,N_2006);
nor U4229 (N_4229,N_495,N_30);
xnor U4230 (N_4230,N_113,N_2073);
xor U4231 (N_4231,N_2227,N_221);
nand U4232 (N_4232,N_845,N_2250);
nand U4233 (N_4233,N_1862,N_731);
nand U4234 (N_4234,N_796,N_1734);
nor U4235 (N_4235,N_1598,N_1005);
xnor U4236 (N_4236,N_2216,N_1156);
xor U4237 (N_4237,N_276,N_739);
nand U4238 (N_4238,N_1591,N_2351);
and U4239 (N_4239,N_1385,N_730);
nor U4240 (N_4240,N_2267,N_2141);
or U4241 (N_4241,N_1855,N_186);
or U4242 (N_4242,N_2066,N_2151);
nor U4243 (N_4243,N_1182,N_669);
and U4244 (N_4244,N_1579,N_927);
xnor U4245 (N_4245,N_177,N_1130);
xor U4246 (N_4246,N_307,N_543);
nand U4247 (N_4247,N_685,N_2311);
xor U4248 (N_4248,N_222,N_2069);
xor U4249 (N_4249,N_1742,N_692);
nand U4250 (N_4250,N_626,N_944);
and U4251 (N_4251,N_254,N_224);
and U4252 (N_4252,N_1174,N_1683);
and U4253 (N_4253,N_799,N_41);
xnor U4254 (N_4254,N_2,N_1084);
xnor U4255 (N_4255,N_1831,N_1949);
and U4256 (N_4256,N_1215,N_2457);
nand U4257 (N_4257,N_1599,N_1870);
or U4258 (N_4258,N_737,N_624);
nor U4259 (N_4259,N_665,N_437);
xor U4260 (N_4260,N_1287,N_951);
xnor U4261 (N_4261,N_1153,N_1363);
and U4262 (N_4262,N_2363,N_1968);
nand U4263 (N_4263,N_1148,N_106);
xor U4264 (N_4264,N_2185,N_747);
or U4265 (N_4265,N_523,N_1368);
xor U4266 (N_4266,N_1691,N_1883);
nand U4267 (N_4267,N_637,N_1968);
or U4268 (N_4268,N_1299,N_2053);
nand U4269 (N_4269,N_327,N_515);
or U4270 (N_4270,N_1493,N_1011);
nor U4271 (N_4271,N_1666,N_1683);
nand U4272 (N_4272,N_2180,N_1558);
or U4273 (N_4273,N_2221,N_1685);
xor U4274 (N_4274,N_517,N_959);
nor U4275 (N_4275,N_1664,N_1606);
or U4276 (N_4276,N_1841,N_1396);
or U4277 (N_4277,N_1651,N_1307);
or U4278 (N_4278,N_1959,N_1255);
xnor U4279 (N_4279,N_1801,N_1213);
nand U4280 (N_4280,N_1566,N_1278);
or U4281 (N_4281,N_1163,N_839);
and U4282 (N_4282,N_2479,N_110);
and U4283 (N_4283,N_899,N_2342);
xor U4284 (N_4284,N_1953,N_1379);
or U4285 (N_4285,N_794,N_313);
nand U4286 (N_4286,N_1355,N_2007);
and U4287 (N_4287,N_255,N_2139);
xor U4288 (N_4288,N_937,N_2485);
xnor U4289 (N_4289,N_2189,N_2442);
xor U4290 (N_4290,N_722,N_445);
nor U4291 (N_4291,N_247,N_1886);
nor U4292 (N_4292,N_175,N_1932);
nand U4293 (N_4293,N_1782,N_2337);
nand U4294 (N_4294,N_305,N_1545);
nand U4295 (N_4295,N_344,N_1437);
nand U4296 (N_4296,N_365,N_1958);
nand U4297 (N_4297,N_1478,N_14);
nand U4298 (N_4298,N_1744,N_2414);
nand U4299 (N_4299,N_1149,N_1923);
and U4300 (N_4300,N_2368,N_2479);
and U4301 (N_4301,N_110,N_78);
and U4302 (N_4302,N_1121,N_263);
xnor U4303 (N_4303,N_2116,N_1271);
xnor U4304 (N_4304,N_488,N_166);
nor U4305 (N_4305,N_2115,N_363);
or U4306 (N_4306,N_195,N_921);
or U4307 (N_4307,N_727,N_495);
xnor U4308 (N_4308,N_731,N_1385);
nor U4309 (N_4309,N_2290,N_1821);
and U4310 (N_4310,N_1694,N_815);
xnor U4311 (N_4311,N_2128,N_1439);
nand U4312 (N_4312,N_1519,N_851);
or U4313 (N_4313,N_2235,N_2182);
nand U4314 (N_4314,N_1459,N_2216);
xor U4315 (N_4315,N_499,N_583);
or U4316 (N_4316,N_2072,N_2001);
xnor U4317 (N_4317,N_2159,N_925);
nand U4318 (N_4318,N_1330,N_649);
nand U4319 (N_4319,N_1316,N_989);
or U4320 (N_4320,N_2107,N_2012);
nand U4321 (N_4321,N_2231,N_1297);
or U4322 (N_4322,N_1173,N_720);
nand U4323 (N_4323,N_393,N_1871);
or U4324 (N_4324,N_316,N_2396);
or U4325 (N_4325,N_941,N_437);
xnor U4326 (N_4326,N_512,N_1333);
or U4327 (N_4327,N_2086,N_87);
nor U4328 (N_4328,N_1113,N_1929);
nand U4329 (N_4329,N_388,N_468);
nand U4330 (N_4330,N_1612,N_1296);
nand U4331 (N_4331,N_2286,N_769);
xnor U4332 (N_4332,N_1156,N_2395);
nand U4333 (N_4333,N_1771,N_1293);
nor U4334 (N_4334,N_2403,N_1990);
or U4335 (N_4335,N_1921,N_2021);
xor U4336 (N_4336,N_1439,N_459);
or U4337 (N_4337,N_1334,N_1156);
nor U4338 (N_4338,N_1071,N_154);
and U4339 (N_4339,N_797,N_1298);
or U4340 (N_4340,N_494,N_85);
nor U4341 (N_4341,N_1195,N_1768);
or U4342 (N_4342,N_1010,N_1710);
and U4343 (N_4343,N_127,N_1423);
nor U4344 (N_4344,N_1867,N_931);
nand U4345 (N_4345,N_1534,N_299);
nor U4346 (N_4346,N_151,N_1517);
nand U4347 (N_4347,N_1099,N_297);
and U4348 (N_4348,N_754,N_267);
or U4349 (N_4349,N_159,N_2196);
and U4350 (N_4350,N_691,N_1963);
and U4351 (N_4351,N_68,N_1910);
and U4352 (N_4352,N_1085,N_2236);
nand U4353 (N_4353,N_1596,N_782);
nor U4354 (N_4354,N_1939,N_2477);
xor U4355 (N_4355,N_1245,N_1163);
xnor U4356 (N_4356,N_292,N_1004);
xor U4357 (N_4357,N_825,N_964);
nor U4358 (N_4358,N_596,N_1700);
or U4359 (N_4359,N_97,N_1628);
nand U4360 (N_4360,N_1578,N_562);
nand U4361 (N_4361,N_1886,N_953);
xnor U4362 (N_4362,N_1545,N_1244);
and U4363 (N_4363,N_197,N_1829);
nor U4364 (N_4364,N_1547,N_864);
xnor U4365 (N_4365,N_946,N_2434);
or U4366 (N_4366,N_1318,N_1589);
xor U4367 (N_4367,N_402,N_2012);
and U4368 (N_4368,N_1407,N_1748);
xor U4369 (N_4369,N_25,N_303);
nand U4370 (N_4370,N_614,N_1652);
and U4371 (N_4371,N_1284,N_459);
and U4372 (N_4372,N_1352,N_1427);
or U4373 (N_4373,N_1524,N_201);
xor U4374 (N_4374,N_138,N_38);
and U4375 (N_4375,N_1857,N_1509);
nor U4376 (N_4376,N_2180,N_1113);
nor U4377 (N_4377,N_2060,N_517);
or U4378 (N_4378,N_803,N_1827);
nor U4379 (N_4379,N_504,N_726);
xnor U4380 (N_4380,N_1727,N_578);
nor U4381 (N_4381,N_523,N_164);
and U4382 (N_4382,N_445,N_149);
nor U4383 (N_4383,N_927,N_2270);
nand U4384 (N_4384,N_1365,N_1966);
and U4385 (N_4385,N_1869,N_450);
and U4386 (N_4386,N_470,N_1325);
xor U4387 (N_4387,N_868,N_86);
or U4388 (N_4388,N_1382,N_2196);
xor U4389 (N_4389,N_2204,N_1914);
nand U4390 (N_4390,N_49,N_482);
xor U4391 (N_4391,N_1435,N_1702);
and U4392 (N_4392,N_683,N_270);
and U4393 (N_4393,N_2125,N_640);
or U4394 (N_4394,N_1547,N_1580);
or U4395 (N_4395,N_1467,N_937);
xnor U4396 (N_4396,N_249,N_1557);
and U4397 (N_4397,N_2408,N_727);
and U4398 (N_4398,N_737,N_301);
nand U4399 (N_4399,N_1350,N_1217);
and U4400 (N_4400,N_700,N_594);
nor U4401 (N_4401,N_76,N_2283);
nand U4402 (N_4402,N_1051,N_609);
and U4403 (N_4403,N_495,N_1847);
and U4404 (N_4404,N_2416,N_2240);
xor U4405 (N_4405,N_1791,N_1972);
and U4406 (N_4406,N_1522,N_1587);
or U4407 (N_4407,N_996,N_1682);
and U4408 (N_4408,N_1306,N_1419);
xor U4409 (N_4409,N_766,N_2129);
and U4410 (N_4410,N_2404,N_768);
xnor U4411 (N_4411,N_1015,N_2494);
nor U4412 (N_4412,N_524,N_1346);
nor U4413 (N_4413,N_526,N_2170);
or U4414 (N_4414,N_1892,N_441);
or U4415 (N_4415,N_150,N_401);
nor U4416 (N_4416,N_1438,N_2486);
nor U4417 (N_4417,N_2139,N_657);
nor U4418 (N_4418,N_503,N_110);
nor U4419 (N_4419,N_212,N_246);
or U4420 (N_4420,N_1667,N_1538);
nand U4421 (N_4421,N_1795,N_758);
or U4422 (N_4422,N_2051,N_1005);
nand U4423 (N_4423,N_474,N_2070);
xor U4424 (N_4424,N_2478,N_807);
xor U4425 (N_4425,N_2461,N_2015);
nand U4426 (N_4426,N_442,N_2081);
xor U4427 (N_4427,N_2154,N_1872);
and U4428 (N_4428,N_1856,N_1232);
xnor U4429 (N_4429,N_59,N_1576);
or U4430 (N_4430,N_1460,N_1325);
nor U4431 (N_4431,N_420,N_1420);
nor U4432 (N_4432,N_2242,N_2004);
or U4433 (N_4433,N_492,N_18);
xnor U4434 (N_4434,N_941,N_1099);
xnor U4435 (N_4435,N_980,N_1459);
and U4436 (N_4436,N_2087,N_2335);
xnor U4437 (N_4437,N_2224,N_1949);
and U4438 (N_4438,N_490,N_138);
nand U4439 (N_4439,N_1694,N_2022);
or U4440 (N_4440,N_2070,N_1490);
or U4441 (N_4441,N_2436,N_950);
and U4442 (N_4442,N_2114,N_320);
xor U4443 (N_4443,N_1783,N_45);
nand U4444 (N_4444,N_1437,N_48);
xnor U4445 (N_4445,N_1834,N_269);
and U4446 (N_4446,N_920,N_648);
xnor U4447 (N_4447,N_398,N_432);
or U4448 (N_4448,N_853,N_396);
nor U4449 (N_4449,N_1592,N_508);
nor U4450 (N_4450,N_1863,N_691);
or U4451 (N_4451,N_1886,N_678);
and U4452 (N_4452,N_2234,N_1189);
or U4453 (N_4453,N_1892,N_2079);
xor U4454 (N_4454,N_695,N_52);
xnor U4455 (N_4455,N_565,N_1157);
xnor U4456 (N_4456,N_2320,N_533);
and U4457 (N_4457,N_785,N_2205);
or U4458 (N_4458,N_726,N_2303);
nor U4459 (N_4459,N_1878,N_2333);
or U4460 (N_4460,N_2452,N_1269);
or U4461 (N_4461,N_1003,N_531);
xor U4462 (N_4462,N_2047,N_137);
xor U4463 (N_4463,N_1519,N_2177);
nand U4464 (N_4464,N_1654,N_2399);
nor U4465 (N_4465,N_200,N_1268);
and U4466 (N_4466,N_1992,N_1204);
and U4467 (N_4467,N_623,N_720);
or U4468 (N_4468,N_2458,N_2244);
nand U4469 (N_4469,N_819,N_998);
xor U4470 (N_4470,N_481,N_2328);
and U4471 (N_4471,N_2241,N_382);
nand U4472 (N_4472,N_2026,N_1145);
xnor U4473 (N_4473,N_823,N_1724);
xnor U4474 (N_4474,N_1594,N_1326);
or U4475 (N_4475,N_846,N_1317);
and U4476 (N_4476,N_194,N_1047);
and U4477 (N_4477,N_1798,N_2126);
nor U4478 (N_4478,N_475,N_2053);
or U4479 (N_4479,N_2336,N_1186);
and U4480 (N_4480,N_1818,N_855);
nand U4481 (N_4481,N_1082,N_1060);
or U4482 (N_4482,N_115,N_858);
and U4483 (N_4483,N_864,N_639);
and U4484 (N_4484,N_1146,N_490);
or U4485 (N_4485,N_626,N_1772);
nand U4486 (N_4486,N_1596,N_2053);
and U4487 (N_4487,N_618,N_321);
nor U4488 (N_4488,N_322,N_352);
and U4489 (N_4489,N_2183,N_516);
nor U4490 (N_4490,N_201,N_1614);
xnor U4491 (N_4491,N_841,N_1032);
or U4492 (N_4492,N_1449,N_868);
nand U4493 (N_4493,N_2017,N_754);
xnor U4494 (N_4494,N_827,N_140);
or U4495 (N_4495,N_418,N_330);
nor U4496 (N_4496,N_358,N_1032);
or U4497 (N_4497,N_2037,N_190);
and U4498 (N_4498,N_1577,N_886);
nor U4499 (N_4499,N_1885,N_2492);
and U4500 (N_4500,N_737,N_1667);
and U4501 (N_4501,N_35,N_1252);
and U4502 (N_4502,N_1666,N_2311);
or U4503 (N_4503,N_134,N_1285);
xnor U4504 (N_4504,N_1912,N_2002);
nand U4505 (N_4505,N_2179,N_1714);
and U4506 (N_4506,N_116,N_121);
xnor U4507 (N_4507,N_431,N_1151);
and U4508 (N_4508,N_1039,N_102);
and U4509 (N_4509,N_1780,N_457);
nand U4510 (N_4510,N_2367,N_1685);
and U4511 (N_4511,N_688,N_2458);
and U4512 (N_4512,N_499,N_194);
xor U4513 (N_4513,N_1526,N_1810);
xor U4514 (N_4514,N_212,N_2194);
nand U4515 (N_4515,N_57,N_2068);
xnor U4516 (N_4516,N_616,N_1023);
nand U4517 (N_4517,N_778,N_607);
nor U4518 (N_4518,N_367,N_1261);
nor U4519 (N_4519,N_1879,N_1083);
xor U4520 (N_4520,N_609,N_2129);
nor U4521 (N_4521,N_1634,N_2329);
or U4522 (N_4522,N_1996,N_2151);
xnor U4523 (N_4523,N_588,N_2452);
nor U4524 (N_4524,N_94,N_900);
nand U4525 (N_4525,N_822,N_2482);
nor U4526 (N_4526,N_1347,N_1642);
nand U4527 (N_4527,N_286,N_323);
or U4528 (N_4528,N_221,N_2206);
and U4529 (N_4529,N_1276,N_1908);
xnor U4530 (N_4530,N_247,N_1296);
or U4531 (N_4531,N_2412,N_845);
and U4532 (N_4532,N_2236,N_172);
or U4533 (N_4533,N_2406,N_1775);
nor U4534 (N_4534,N_89,N_405);
nand U4535 (N_4535,N_1538,N_1418);
or U4536 (N_4536,N_586,N_882);
and U4537 (N_4537,N_996,N_688);
nor U4538 (N_4538,N_741,N_1186);
nor U4539 (N_4539,N_860,N_1795);
xor U4540 (N_4540,N_2045,N_112);
nor U4541 (N_4541,N_586,N_909);
xor U4542 (N_4542,N_560,N_2214);
and U4543 (N_4543,N_674,N_869);
nor U4544 (N_4544,N_1076,N_79);
or U4545 (N_4545,N_2284,N_945);
nor U4546 (N_4546,N_1130,N_2183);
xnor U4547 (N_4547,N_641,N_2493);
nor U4548 (N_4548,N_1677,N_766);
or U4549 (N_4549,N_1354,N_2033);
and U4550 (N_4550,N_2240,N_2188);
nor U4551 (N_4551,N_750,N_66);
or U4552 (N_4552,N_296,N_1895);
xor U4553 (N_4553,N_416,N_2019);
or U4554 (N_4554,N_225,N_841);
nor U4555 (N_4555,N_1577,N_1779);
or U4556 (N_4556,N_2299,N_1598);
xnor U4557 (N_4557,N_1237,N_1178);
and U4558 (N_4558,N_1097,N_1485);
nor U4559 (N_4559,N_280,N_1813);
and U4560 (N_4560,N_1531,N_71);
or U4561 (N_4561,N_577,N_2078);
nand U4562 (N_4562,N_1179,N_487);
or U4563 (N_4563,N_241,N_459);
xor U4564 (N_4564,N_703,N_596);
and U4565 (N_4565,N_191,N_201);
xnor U4566 (N_4566,N_571,N_1895);
nand U4567 (N_4567,N_862,N_952);
and U4568 (N_4568,N_1371,N_1301);
nor U4569 (N_4569,N_545,N_1816);
nand U4570 (N_4570,N_1337,N_1516);
nor U4571 (N_4571,N_1282,N_922);
and U4572 (N_4572,N_1883,N_809);
or U4573 (N_4573,N_1859,N_916);
nand U4574 (N_4574,N_1386,N_2372);
nor U4575 (N_4575,N_190,N_2477);
or U4576 (N_4576,N_1029,N_924);
or U4577 (N_4577,N_2297,N_2344);
or U4578 (N_4578,N_2132,N_1807);
nand U4579 (N_4579,N_1690,N_2336);
nor U4580 (N_4580,N_898,N_1376);
and U4581 (N_4581,N_1796,N_1761);
or U4582 (N_4582,N_1669,N_538);
nor U4583 (N_4583,N_193,N_2237);
xnor U4584 (N_4584,N_2074,N_788);
nand U4585 (N_4585,N_1707,N_1804);
xor U4586 (N_4586,N_2130,N_481);
or U4587 (N_4587,N_1153,N_766);
nor U4588 (N_4588,N_1272,N_1888);
xor U4589 (N_4589,N_1020,N_1393);
or U4590 (N_4590,N_1994,N_1137);
and U4591 (N_4591,N_1259,N_1879);
and U4592 (N_4592,N_1858,N_45);
and U4593 (N_4593,N_1833,N_632);
and U4594 (N_4594,N_824,N_2459);
nor U4595 (N_4595,N_704,N_925);
nand U4596 (N_4596,N_1603,N_589);
or U4597 (N_4597,N_575,N_20);
and U4598 (N_4598,N_427,N_1934);
nor U4599 (N_4599,N_133,N_1563);
and U4600 (N_4600,N_829,N_1259);
nand U4601 (N_4601,N_749,N_193);
nor U4602 (N_4602,N_229,N_1192);
and U4603 (N_4603,N_840,N_1180);
nor U4604 (N_4604,N_2494,N_2189);
nor U4605 (N_4605,N_1181,N_546);
nor U4606 (N_4606,N_1945,N_1909);
nor U4607 (N_4607,N_1035,N_1157);
and U4608 (N_4608,N_172,N_1611);
nand U4609 (N_4609,N_1018,N_986);
and U4610 (N_4610,N_889,N_258);
xor U4611 (N_4611,N_1605,N_1360);
nor U4612 (N_4612,N_2032,N_1817);
or U4613 (N_4613,N_2455,N_2250);
and U4614 (N_4614,N_1292,N_632);
and U4615 (N_4615,N_1263,N_1249);
nor U4616 (N_4616,N_1249,N_218);
nand U4617 (N_4617,N_1188,N_1819);
or U4618 (N_4618,N_2174,N_1204);
nor U4619 (N_4619,N_2264,N_321);
xor U4620 (N_4620,N_245,N_1696);
nand U4621 (N_4621,N_749,N_2281);
and U4622 (N_4622,N_1114,N_1754);
or U4623 (N_4623,N_112,N_379);
nand U4624 (N_4624,N_1072,N_1491);
nor U4625 (N_4625,N_1206,N_868);
nand U4626 (N_4626,N_1872,N_1196);
nand U4627 (N_4627,N_2322,N_851);
xor U4628 (N_4628,N_1563,N_840);
nand U4629 (N_4629,N_1504,N_2155);
nand U4630 (N_4630,N_854,N_2234);
nand U4631 (N_4631,N_1165,N_494);
and U4632 (N_4632,N_2420,N_536);
nand U4633 (N_4633,N_2289,N_1147);
or U4634 (N_4634,N_1516,N_908);
xor U4635 (N_4635,N_1775,N_499);
or U4636 (N_4636,N_1912,N_504);
xnor U4637 (N_4637,N_1120,N_597);
and U4638 (N_4638,N_1821,N_331);
xor U4639 (N_4639,N_1549,N_1072);
xor U4640 (N_4640,N_823,N_1438);
or U4641 (N_4641,N_1677,N_1358);
and U4642 (N_4642,N_1361,N_569);
xnor U4643 (N_4643,N_1824,N_1253);
nor U4644 (N_4644,N_74,N_336);
xor U4645 (N_4645,N_1165,N_572);
and U4646 (N_4646,N_2389,N_684);
or U4647 (N_4647,N_909,N_1873);
and U4648 (N_4648,N_1296,N_819);
and U4649 (N_4649,N_2261,N_1430);
or U4650 (N_4650,N_2348,N_2445);
or U4651 (N_4651,N_1263,N_1477);
xor U4652 (N_4652,N_375,N_784);
and U4653 (N_4653,N_1082,N_798);
nor U4654 (N_4654,N_2407,N_353);
and U4655 (N_4655,N_927,N_2114);
nor U4656 (N_4656,N_1605,N_1051);
nor U4657 (N_4657,N_678,N_47);
or U4658 (N_4658,N_1397,N_416);
nand U4659 (N_4659,N_1370,N_1709);
or U4660 (N_4660,N_2274,N_428);
nor U4661 (N_4661,N_1624,N_1451);
and U4662 (N_4662,N_69,N_541);
xor U4663 (N_4663,N_940,N_1034);
or U4664 (N_4664,N_2165,N_1153);
or U4665 (N_4665,N_688,N_867);
nor U4666 (N_4666,N_1233,N_229);
nor U4667 (N_4667,N_1514,N_1239);
or U4668 (N_4668,N_2320,N_1703);
nor U4669 (N_4669,N_583,N_2233);
nand U4670 (N_4670,N_1064,N_426);
and U4671 (N_4671,N_204,N_679);
nand U4672 (N_4672,N_2312,N_2287);
or U4673 (N_4673,N_1091,N_1845);
nor U4674 (N_4674,N_696,N_1919);
and U4675 (N_4675,N_445,N_2033);
nor U4676 (N_4676,N_2387,N_477);
nand U4677 (N_4677,N_329,N_1833);
nand U4678 (N_4678,N_704,N_1582);
and U4679 (N_4679,N_1425,N_1723);
or U4680 (N_4680,N_658,N_1018);
or U4681 (N_4681,N_1011,N_1142);
nand U4682 (N_4682,N_764,N_2245);
nand U4683 (N_4683,N_2064,N_155);
or U4684 (N_4684,N_41,N_2317);
xor U4685 (N_4685,N_1596,N_683);
and U4686 (N_4686,N_1391,N_731);
nand U4687 (N_4687,N_2369,N_524);
and U4688 (N_4688,N_1359,N_238);
nand U4689 (N_4689,N_1695,N_633);
nor U4690 (N_4690,N_1720,N_143);
nor U4691 (N_4691,N_2403,N_2409);
nand U4692 (N_4692,N_2118,N_880);
nand U4693 (N_4693,N_1120,N_811);
and U4694 (N_4694,N_935,N_1624);
or U4695 (N_4695,N_2413,N_2254);
or U4696 (N_4696,N_1561,N_1312);
or U4697 (N_4697,N_786,N_1528);
or U4698 (N_4698,N_2085,N_649);
and U4699 (N_4699,N_2052,N_993);
or U4700 (N_4700,N_1351,N_453);
and U4701 (N_4701,N_1171,N_1031);
nor U4702 (N_4702,N_1191,N_2359);
xnor U4703 (N_4703,N_18,N_1394);
or U4704 (N_4704,N_254,N_112);
or U4705 (N_4705,N_783,N_236);
and U4706 (N_4706,N_1759,N_2314);
and U4707 (N_4707,N_1493,N_604);
nand U4708 (N_4708,N_407,N_1505);
nor U4709 (N_4709,N_286,N_2324);
and U4710 (N_4710,N_507,N_1827);
xnor U4711 (N_4711,N_2497,N_732);
and U4712 (N_4712,N_503,N_1931);
or U4713 (N_4713,N_1446,N_521);
nor U4714 (N_4714,N_96,N_2359);
or U4715 (N_4715,N_1527,N_2169);
nand U4716 (N_4716,N_1534,N_1944);
nand U4717 (N_4717,N_499,N_1110);
nor U4718 (N_4718,N_2033,N_2410);
nand U4719 (N_4719,N_731,N_734);
and U4720 (N_4720,N_1267,N_2308);
or U4721 (N_4721,N_40,N_410);
or U4722 (N_4722,N_1670,N_1310);
nand U4723 (N_4723,N_183,N_1991);
and U4724 (N_4724,N_565,N_2318);
xor U4725 (N_4725,N_2385,N_2180);
nor U4726 (N_4726,N_2430,N_2445);
nand U4727 (N_4727,N_108,N_1744);
nor U4728 (N_4728,N_628,N_73);
xor U4729 (N_4729,N_2424,N_2414);
nor U4730 (N_4730,N_1329,N_576);
and U4731 (N_4731,N_1642,N_1585);
xnor U4732 (N_4732,N_1104,N_2375);
and U4733 (N_4733,N_743,N_1706);
and U4734 (N_4734,N_2345,N_2115);
or U4735 (N_4735,N_831,N_1413);
and U4736 (N_4736,N_1601,N_368);
and U4737 (N_4737,N_1766,N_2052);
xnor U4738 (N_4738,N_389,N_1184);
xor U4739 (N_4739,N_767,N_1225);
and U4740 (N_4740,N_1674,N_833);
nor U4741 (N_4741,N_1840,N_1938);
xor U4742 (N_4742,N_1609,N_1992);
nor U4743 (N_4743,N_975,N_2473);
xnor U4744 (N_4744,N_1478,N_2130);
xnor U4745 (N_4745,N_231,N_451);
or U4746 (N_4746,N_89,N_211);
nand U4747 (N_4747,N_544,N_376);
and U4748 (N_4748,N_1413,N_2044);
nand U4749 (N_4749,N_2396,N_1193);
or U4750 (N_4750,N_70,N_1567);
nand U4751 (N_4751,N_859,N_1304);
xor U4752 (N_4752,N_1842,N_16);
nor U4753 (N_4753,N_1641,N_458);
nor U4754 (N_4754,N_16,N_2158);
or U4755 (N_4755,N_1661,N_2154);
xor U4756 (N_4756,N_933,N_0);
nor U4757 (N_4757,N_1706,N_2474);
nand U4758 (N_4758,N_711,N_2084);
xnor U4759 (N_4759,N_454,N_1848);
nand U4760 (N_4760,N_1386,N_2421);
nor U4761 (N_4761,N_2245,N_2475);
nand U4762 (N_4762,N_1651,N_37);
or U4763 (N_4763,N_208,N_1747);
xnor U4764 (N_4764,N_2477,N_2227);
xnor U4765 (N_4765,N_762,N_1365);
or U4766 (N_4766,N_1404,N_561);
and U4767 (N_4767,N_995,N_898);
xor U4768 (N_4768,N_1584,N_1324);
nand U4769 (N_4769,N_2312,N_1671);
or U4770 (N_4770,N_758,N_599);
or U4771 (N_4771,N_1765,N_2019);
nor U4772 (N_4772,N_1469,N_2161);
xor U4773 (N_4773,N_1328,N_1081);
or U4774 (N_4774,N_1129,N_1358);
or U4775 (N_4775,N_175,N_2035);
and U4776 (N_4776,N_1688,N_2337);
xnor U4777 (N_4777,N_2169,N_945);
nor U4778 (N_4778,N_188,N_1072);
xor U4779 (N_4779,N_367,N_737);
or U4780 (N_4780,N_1055,N_2345);
xor U4781 (N_4781,N_1643,N_2159);
or U4782 (N_4782,N_1504,N_1097);
or U4783 (N_4783,N_106,N_1244);
xor U4784 (N_4784,N_786,N_1580);
and U4785 (N_4785,N_505,N_2294);
nand U4786 (N_4786,N_2009,N_801);
and U4787 (N_4787,N_1731,N_662);
nand U4788 (N_4788,N_1272,N_1026);
xnor U4789 (N_4789,N_2071,N_1941);
xnor U4790 (N_4790,N_786,N_1837);
nor U4791 (N_4791,N_6,N_2231);
xnor U4792 (N_4792,N_1979,N_1535);
nand U4793 (N_4793,N_1603,N_1470);
and U4794 (N_4794,N_1465,N_1307);
nor U4795 (N_4795,N_708,N_2019);
nand U4796 (N_4796,N_737,N_1733);
nand U4797 (N_4797,N_1643,N_1454);
nor U4798 (N_4798,N_2495,N_612);
nor U4799 (N_4799,N_242,N_331);
and U4800 (N_4800,N_1621,N_1587);
nand U4801 (N_4801,N_1992,N_1056);
and U4802 (N_4802,N_1346,N_817);
xnor U4803 (N_4803,N_2428,N_2096);
or U4804 (N_4804,N_402,N_1812);
or U4805 (N_4805,N_1639,N_1867);
xnor U4806 (N_4806,N_2367,N_1857);
nand U4807 (N_4807,N_741,N_1826);
xnor U4808 (N_4808,N_1932,N_1519);
xor U4809 (N_4809,N_775,N_1475);
nor U4810 (N_4810,N_1772,N_2065);
nor U4811 (N_4811,N_561,N_2361);
or U4812 (N_4812,N_806,N_1387);
nor U4813 (N_4813,N_1818,N_111);
nor U4814 (N_4814,N_10,N_1292);
nand U4815 (N_4815,N_1087,N_403);
xnor U4816 (N_4816,N_1353,N_1582);
xnor U4817 (N_4817,N_2255,N_200);
or U4818 (N_4818,N_2133,N_1285);
nor U4819 (N_4819,N_1385,N_1233);
and U4820 (N_4820,N_1913,N_1516);
and U4821 (N_4821,N_1456,N_1117);
and U4822 (N_4822,N_2229,N_1622);
nor U4823 (N_4823,N_345,N_817);
xnor U4824 (N_4824,N_1843,N_1714);
or U4825 (N_4825,N_420,N_301);
nor U4826 (N_4826,N_508,N_107);
xor U4827 (N_4827,N_1584,N_2330);
xnor U4828 (N_4828,N_941,N_314);
or U4829 (N_4829,N_2082,N_869);
and U4830 (N_4830,N_199,N_742);
xor U4831 (N_4831,N_2091,N_829);
nor U4832 (N_4832,N_2465,N_2021);
xor U4833 (N_4833,N_1306,N_7);
or U4834 (N_4834,N_1840,N_2352);
or U4835 (N_4835,N_1174,N_430);
nor U4836 (N_4836,N_417,N_1466);
nor U4837 (N_4837,N_1540,N_2287);
nor U4838 (N_4838,N_888,N_1122);
nand U4839 (N_4839,N_1122,N_414);
nor U4840 (N_4840,N_1767,N_137);
and U4841 (N_4841,N_1439,N_1571);
or U4842 (N_4842,N_1426,N_617);
and U4843 (N_4843,N_2053,N_1645);
nand U4844 (N_4844,N_602,N_450);
or U4845 (N_4845,N_1235,N_1403);
nand U4846 (N_4846,N_2461,N_995);
nor U4847 (N_4847,N_1227,N_2223);
xnor U4848 (N_4848,N_1858,N_2167);
nand U4849 (N_4849,N_2099,N_2265);
and U4850 (N_4850,N_2167,N_547);
or U4851 (N_4851,N_257,N_459);
or U4852 (N_4852,N_1684,N_705);
nor U4853 (N_4853,N_1271,N_1186);
xnor U4854 (N_4854,N_672,N_870);
or U4855 (N_4855,N_1768,N_1037);
xnor U4856 (N_4856,N_2216,N_262);
nor U4857 (N_4857,N_656,N_1780);
xnor U4858 (N_4858,N_1088,N_2083);
and U4859 (N_4859,N_358,N_1003);
xor U4860 (N_4860,N_49,N_1989);
and U4861 (N_4861,N_853,N_2345);
and U4862 (N_4862,N_111,N_1356);
nand U4863 (N_4863,N_964,N_1573);
nor U4864 (N_4864,N_1013,N_1101);
and U4865 (N_4865,N_1841,N_1450);
nor U4866 (N_4866,N_1055,N_1599);
nor U4867 (N_4867,N_1815,N_47);
and U4868 (N_4868,N_1821,N_1680);
and U4869 (N_4869,N_458,N_18);
xnor U4870 (N_4870,N_2383,N_2136);
nand U4871 (N_4871,N_169,N_23);
and U4872 (N_4872,N_2472,N_2355);
and U4873 (N_4873,N_1135,N_1757);
and U4874 (N_4874,N_927,N_1570);
nor U4875 (N_4875,N_2122,N_1078);
and U4876 (N_4876,N_1290,N_323);
or U4877 (N_4877,N_865,N_1672);
or U4878 (N_4878,N_1289,N_2451);
nor U4879 (N_4879,N_583,N_2243);
nand U4880 (N_4880,N_7,N_2031);
or U4881 (N_4881,N_664,N_1878);
nand U4882 (N_4882,N_957,N_493);
nor U4883 (N_4883,N_637,N_18);
nand U4884 (N_4884,N_750,N_422);
and U4885 (N_4885,N_2330,N_169);
nor U4886 (N_4886,N_1853,N_1311);
xor U4887 (N_4887,N_1051,N_949);
nand U4888 (N_4888,N_1087,N_367);
or U4889 (N_4889,N_976,N_1899);
or U4890 (N_4890,N_1348,N_2069);
nand U4891 (N_4891,N_29,N_2355);
nor U4892 (N_4892,N_698,N_2033);
or U4893 (N_4893,N_734,N_1774);
xor U4894 (N_4894,N_2426,N_189);
or U4895 (N_4895,N_1062,N_179);
nand U4896 (N_4896,N_117,N_2010);
xor U4897 (N_4897,N_318,N_745);
nand U4898 (N_4898,N_904,N_2038);
or U4899 (N_4899,N_1350,N_2466);
xnor U4900 (N_4900,N_585,N_465);
nor U4901 (N_4901,N_866,N_1577);
xor U4902 (N_4902,N_708,N_121);
nor U4903 (N_4903,N_2032,N_2254);
nor U4904 (N_4904,N_271,N_1285);
or U4905 (N_4905,N_1068,N_1403);
nor U4906 (N_4906,N_1762,N_2430);
nand U4907 (N_4907,N_2333,N_1166);
nand U4908 (N_4908,N_2283,N_1951);
nor U4909 (N_4909,N_408,N_1242);
nor U4910 (N_4910,N_1033,N_554);
nor U4911 (N_4911,N_43,N_440);
or U4912 (N_4912,N_2463,N_1634);
xor U4913 (N_4913,N_998,N_986);
and U4914 (N_4914,N_2258,N_1782);
xnor U4915 (N_4915,N_740,N_1001);
and U4916 (N_4916,N_2438,N_164);
or U4917 (N_4917,N_1387,N_2115);
or U4918 (N_4918,N_587,N_449);
or U4919 (N_4919,N_1613,N_1865);
nand U4920 (N_4920,N_1114,N_693);
xor U4921 (N_4921,N_1038,N_1004);
nand U4922 (N_4922,N_1215,N_222);
nand U4923 (N_4923,N_1138,N_2273);
nor U4924 (N_4924,N_256,N_522);
nor U4925 (N_4925,N_1495,N_2472);
xnor U4926 (N_4926,N_656,N_332);
nor U4927 (N_4927,N_610,N_93);
nand U4928 (N_4928,N_925,N_1243);
and U4929 (N_4929,N_1112,N_2173);
and U4930 (N_4930,N_1219,N_1043);
nand U4931 (N_4931,N_1621,N_458);
xnor U4932 (N_4932,N_271,N_2149);
nor U4933 (N_4933,N_670,N_223);
and U4934 (N_4934,N_116,N_962);
or U4935 (N_4935,N_892,N_657);
and U4936 (N_4936,N_273,N_854);
and U4937 (N_4937,N_168,N_217);
and U4938 (N_4938,N_914,N_1811);
nand U4939 (N_4939,N_1269,N_489);
or U4940 (N_4940,N_680,N_315);
and U4941 (N_4941,N_298,N_2492);
nand U4942 (N_4942,N_237,N_1615);
nand U4943 (N_4943,N_1258,N_42);
nor U4944 (N_4944,N_1268,N_237);
or U4945 (N_4945,N_1679,N_1386);
or U4946 (N_4946,N_1129,N_2491);
nand U4947 (N_4947,N_1734,N_1675);
and U4948 (N_4948,N_1806,N_1746);
nand U4949 (N_4949,N_1306,N_481);
nand U4950 (N_4950,N_768,N_1580);
or U4951 (N_4951,N_2231,N_148);
and U4952 (N_4952,N_1418,N_1820);
or U4953 (N_4953,N_2359,N_2081);
xnor U4954 (N_4954,N_1556,N_2429);
or U4955 (N_4955,N_1740,N_432);
nand U4956 (N_4956,N_2304,N_1274);
and U4957 (N_4957,N_1858,N_1486);
nor U4958 (N_4958,N_428,N_1722);
xnor U4959 (N_4959,N_1629,N_2440);
xnor U4960 (N_4960,N_1816,N_456);
xnor U4961 (N_4961,N_1853,N_1735);
or U4962 (N_4962,N_2038,N_1356);
or U4963 (N_4963,N_2359,N_1863);
nor U4964 (N_4964,N_912,N_609);
nand U4965 (N_4965,N_1968,N_1362);
and U4966 (N_4966,N_445,N_115);
or U4967 (N_4967,N_210,N_296);
and U4968 (N_4968,N_2419,N_179);
and U4969 (N_4969,N_545,N_549);
xnor U4970 (N_4970,N_1081,N_1232);
or U4971 (N_4971,N_1246,N_1697);
nand U4972 (N_4972,N_91,N_1703);
xor U4973 (N_4973,N_980,N_484);
or U4974 (N_4974,N_157,N_1367);
or U4975 (N_4975,N_683,N_429);
nand U4976 (N_4976,N_298,N_1985);
and U4977 (N_4977,N_956,N_1279);
nor U4978 (N_4978,N_2156,N_203);
nand U4979 (N_4979,N_2343,N_1301);
and U4980 (N_4980,N_1143,N_1427);
or U4981 (N_4981,N_2270,N_1158);
nor U4982 (N_4982,N_685,N_763);
and U4983 (N_4983,N_1415,N_1698);
xnor U4984 (N_4984,N_455,N_2452);
and U4985 (N_4985,N_69,N_529);
and U4986 (N_4986,N_1553,N_1217);
nand U4987 (N_4987,N_529,N_1760);
nor U4988 (N_4988,N_1125,N_2317);
or U4989 (N_4989,N_2479,N_1463);
xnor U4990 (N_4990,N_1592,N_1582);
and U4991 (N_4991,N_2254,N_723);
and U4992 (N_4992,N_833,N_765);
and U4993 (N_4993,N_2205,N_2408);
or U4994 (N_4994,N_1530,N_2298);
nor U4995 (N_4995,N_227,N_805);
nor U4996 (N_4996,N_1365,N_1947);
and U4997 (N_4997,N_1604,N_106);
or U4998 (N_4998,N_1814,N_1861);
nand U4999 (N_4999,N_1593,N_1005);
and U5000 (N_5000,N_2734,N_3888);
nor U5001 (N_5001,N_2625,N_3455);
nor U5002 (N_5002,N_3913,N_2938);
xor U5003 (N_5003,N_4716,N_4599);
and U5004 (N_5004,N_3757,N_3309);
nor U5005 (N_5005,N_4153,N_4732);
or U5006 (N_5006,N_4268,N_3687);
and U5007 (N_5007,N_3993,N_4965);
and U5008 (N_5008,N_3895,N_2699);
and U5009 (N_5009,N_3586,N_3353);
nand U5010 (N_5010,N_3062,N_3192);
xor U5011 (N_5011,N_4162,N_3034);
xnor U5012 (N_5012,N_3686,N_4607);
or U5013 (N_5013,N_3810,N_3580);
or U5014 (N_5014,N_3963,N_4029);
nor U5015 (N_5015,N_3197,N_4438);
xnor U5016 (N_5016,N_4368,N_4609);
and U5017 (N_5017,N_4027,N_3612);
or U5018 (N_5018,N_2793,N_4072);
and U5019 (N_5019,N_2941,N_2729);
xor U5020 (N_5020,N_3097,N_4325);
nor U5021 (N_5021,N_3003,N_4650);
xor U5022 (N_5022,N_4316,N_3106);
xor U5023 (N_5023,N_4206,N_2668);
xnor U5024 (N_5024,N_3819,N_4718);
nor U5025 (N_5025,N_4581,N_4661);
xnor U5026 (N_5026,N_2897,N_4390);
or U5027 (N_5027,N_3500,N_4935);
xor U5028 (N_5028,N_4568,N_2577);
nand U5029 (N_5029,N_3211,N_2836);
and U5030 (N_5030,N_3666,N_3536);
and U5031 (N_5031,N_3294,N_3893);
nor U5032 (N_5032,N_3037,N_4047);
or U5033 (N_5033,N_4647,N_3743);
nor U5034 (N_5034,N_4913,N_3007);
nand U5035 (N_5035,N_3951,N_3774);
xor U5036 (N_5036,N_2531,N_4817);
nand U5037 (N_5037,N_2979,N_4656);
xor U5038 (N_5038,N_4906,N_2722);
xor U5039 (N_5039,N_3877,N_2865);
nand U5040 (N_5040,N_4509,N_3730);
or U5041 (N_5041,N_3792,N_2900);
nor U5042 (N_5042,N_4749,N_3480);
or U5043 (N_5043,N_4256,N_3864);
and U5044 (N_5044,N_3136,N_4665);
nand U5045 (N_5045,N_4202,N_3179);
nor U5046 (N_5046,N_2679,N_3983);
and U5047 (N_5047,N_3701,N_3558);
xnor U5048 (N_5048,N_2864,N_4981);
nand U5049 (N_5049,N_4366,N_4057);
nand U5050 (N_5050,N_4613,N_3869);
or U5051 (N_5051,N_3145,N_4333);
and U5052 (N_5052,N_3191,N_3549);
and U5053 (N_5053,N_4804,N_4184);
or U5054 (N_5054,N_3640,N_3632);
nand U5055 (N_5055,N_4401,N_2942);
nor U5056 (N_5056,N_4707,N_4694);
nand U5057 (N_5057,N_3978,N_4840);
or U5058 (N_5058,N_4264,N_2918);
nor U5059 (N_5059,N_2984,N_3052);
and U5060 (N_5060,N_3302,N_4944);
nor U5061 (N_5061,N_3525,N_4045);
nand U5062 (N_5062,N_4999,N_2891);
and U5063 (N_5063,N_4920,N_4631);
nor U5064 (N_5064,N_3321,N_3867);
xor U5065 (N_5065,N_2527,N_3912);
xnor U5066 (N_5066,N_4957,N_3273);
nand U5067 (N_5067,N_3655,N_3183);
or U5068 (N_5068,N_2766,N_3493);
xor U5069 (N_5069,N_3671,N_3881);
nand U5070 (N_5070,N_3844,N_3826);
and U5071 (N_5071,N_3048,N_4200);
or U5072 (N_5072,N_4159,N_3679);
nand U5073 (N_5073,N_2676,N_3892);
nand U5074 (N_5074,N_4077,N_4942);
nand U5075 (N_5075,N_3718,N_2610);
or U5076 (N_5076,N_3617,N_3470);
nand U5077 (N_5077,N_3138,N_3680);
or U5078 (N_5078,N_2686,N_3648);
or U5079 (N_5079,N_4593,N_2930);
nor U5080 (N_5080,N_3456,N_4535);
nand U5081 (N_5081,N_3256,N_4224);
nor U5082 (N_5082,N_3749,N_4422);
xnor U5083 (N_5083,N_3661,N_4423);
nor U5084 (N_5084,N_3340,N_4721);
nand U5085 (N_5085,N_2619,N_4808);
or U5086 (N_5086,N_3180,N_4834);
and U5087 (N_5087,N_3738,N_3409);
or U5088 (N_5088,N_3146,N_3673);
nand U5089 (N_5089,N_2852,N_2923);
and U5090 (N_5090,N_3334,N_4432);
and U5091 (N_5091,N_3002,N_4505);
nand U5092 (N_5092,N_4270,N_2694);
nand U5093 (N_5093,N_4652,N_4524);
or U5094 (N_5094,N_3204,N_3440);
xor U5095 (N_5095,N_2517,N_4044);
nor U5096 (N_5096,N_3025,N_3071);
xnor U5097 (N_5097,N_2949,N_3290);
and U5098 (N_5098,N_2583,N_4802);
nand U5099 (N_5099,N_4191,N_4570);
nor U5100 (N_5100,N_4812,N_4140);
nand U5101 (N_5101,N_4000,N_2704);
nand U5102 (N_5102,N_4078,N_3605);
and U5103 (N_5103,N_4888,N_4063);
nand U5104 (N_5104,N_4755,N_3221);
nand U5105 (N_5105,N_3501,N_3144);
nand U5106 (N_5106,N_4218,N_2901);
xnor U5107 (N_5107,N_3719,N_2662);
and U5108 (N_5108,N_4810,N_3324);
xnor U5109 (N_5109,N_3459,N_3117);
nor U5110 (N_5110,N_4692,N_4389);
nand U5111 (N_5111,N_2961,N_4091);
and U5112 (N_5112,N_4878,N_4742);
nand U5113 (N_5113,N_4427,N_4708);
xor U5114 (N_5114,N_3156,N_3759);
nand U5115 (N_5115,N_4939,N_3150);
nor U5116 (N_5116,N_4596,N_3153);
or U5117 (N_5117,N_3652,N_2929);
xor U5118 (N_5118,N_2603,N_4618);
xor U5119 (N_5119,N_4553,N_4457);
and U5120 (N_5120,N_3862,N_3254);
or U5121 (N_5121,N_3889,N_2565);
xnor U5122 (N_5122,N_2654,N_4883);
and U5123 (N_5123,N_3027,N_2940);
and U5124 (N_5124,N_3061,N_3429);
xor U5125 (N_5125,N_3331,N_3781);
and U5126 (N_5126,N_2586,N_4624);
and U5127 (N_5127,N_4569,N_4238);
and U5128 (N_5128,N_2711,N_3842);
and U5129 (N_5129,N_3159,N_3975);
nor U5130 (N_5130,N_3289,N_4858);
or U5131 (N_5131,N_3430,N_4658);
and U5132 (N_5132,N_3597,N_3843);
nand U5133 (N_5133,N_2811,N_3506);
nand U5134 (N_5134,N_2713,N_2671);
nor U5135 (N_5135,N_4709,N_3234);
nor U5136 (N_5136,N_3777,N_4467);
nor U5137 (N_5137,N_3583,N_4125);
or U5138 (N_5138,N_4600,N_4902);
or U5139 (N_5139,N_4411,N_4862);
or U5140 (N_5140,N_3207,N_4937);
nor U5141 (N_5141,N_3499,N_4085);
and U5142 (N_5142,N_3075,N_4821);
nand U5143 (N_5143,N_2697,N_4466);
nor U5144 (N_5144,N_4365,N_3858);
and U5145 (N_5145,N_2876,N_2685);
and U5146 (N_5146,N_2636,N_4550);
and U5147 (N_5147,N_2844,N_4105);
xor U5148 (N_5148,N_3389,N_2580);
nor U5149 (N_5149,N_4557,N_3532);
nand U5150 (N_5150,N_2601,N_3291);
or U5151 (N_5151,N_2665,N_3885);
nor U5152 (N_5152,N_3190,N_4727);
and U5153 (N_5153,N_4781,N_4969);
nor U5154 (N_5154,N_4725,N_3335);
nor U5155 (N_5155,N_3036,N_3059);
and U5156 (N_5156,N_4379,N_4783);
nand U5157 (N_5157,N_4204,N_3964);
xor U5158 (N_5158,N_2510,N_2791);
xnor U5159 (N_5159,N_3988,N_3974);
nor U5160 (N_5160,N_4818,N_3836);
or U5161 (N_5161,N_2796,N_4038);
nand U5162 (N_5162,N_4831,N_4070);
or U5163 (N_5163,N_3521,N_3057);
and U5164 (N_5164,N_3930,N_4479);
and U5165 (N_5165,N_4852,N_4470);
and U5166 (N_5166,N_4940,N_4385);
or U5167 (N_5167,N_4829,N_4927);
and U5168 (N_5168,N_4860,N_4436);
nor U5169 (N_5169,N_2725,N_3039);
and U5170 (N_5170,N_4100,N_3219);
nor U5171 (N_5171,N_4219,N_3265);
nand U5172 (N_5172,N_3123,N_4369);
xnor U5173 (N_5173,N_2672,N_2630);
xor U5174 (N_5174,N_3228,N_3905);
nand U5175 (N_5175,N_3396,N_2994);
nor U5176 (N_5176,N_2954,N_3803);
nor U5177 (N_5177,N_4426,N_2647);
or U5178 (N_5178,N_4075,N_3884);
nor U5179 (N_5179,N_3364,N_2969);
or U5180 (N_5180,N_2605,N_4552);
nor U5181 (N_5181,N_4211,N_3972);
or U5182 (N_5182,N_4779,N_2670);
nor U5183 (N_5183,N_3181,N_3275);
and U5184 (N_5184,N_4726,N_4059);
nor U5185 (N_5185,N_3543,N_2526);
xor U5186 (N_5186,N_2569,N_4740);
xor U5187 (N_5187,N_3947,N_3984);
xnor U5188 (N_5188,N_4869,N_2810);
nor U5189 (N_5189,N_4118,N_3997);
or U5190 (N_5190,N_4155,N_2664);
nand U5191 (N_5191,N_3615,N_2945);
nor U5192 (N_5192,N_4166,N_3727);
and U5193 (N_5193,N_4336,N_4290);
nand U5194 (N_5194,N_4022,N_3473);
xnor U5195 (N_5195,N_3613,N_4214);
nand U5196 (N_5196,N_3088,N_2588);
nor U5197 (N_5197,N_4982,N_2785);
nand U5198 (N_5198,N_3220,N_2736);
and U5199 (N_5199,N_4034,N_3789);
nand U5200 (N_5200,N_4803,N_3314);
or U5201 (N_5201,N_3943,N_3526);
nand U5202 (N_5202,N_4510,N_4226);
nand U5203 (N_5203,N_4321,N_3641);
xnor U5204 (N_5204,N_3629,N_4949);
or U5205 (N_5205,N_3255,N_4754);
or U5206 (N_5206,N_3780,N_4319);
nand U5207 (N_5207,N_2747,N_3371);
nor U5208 (N_5208,N_4433,N_4547);
and U5209 (N_5209,N_2626,N_3203);
and U5210 (N_5210,N_4501,N_3315);
nand U5211 (N_5211,N_4586,N_3405);
nand U5212 (N_5212,N_3556,N_3927);
xor U5213 (N_5213,N_2617,N_3401);
nand U5214 (N_5214,N_3354,N_4441);
xor U5215 (N_5215,N_2576,N_3591);
xnor U5216 (N_5216,N_4496,N_3910);
nor U5217 (N_5217,N_2997,N_4203);
and U5218 (N_5218,N_3808,N_4189);
nor U5219 (N_5219,N_3977,N_3938);
nor U5220 (N_5220,N_2982,N_3298);
and U5221 (N_5221,N_4683,N_3735);
or U5222 (N_5222,N_4777,N_4201);
nand U5223 (N_5223,N_4341,N_4799);
or U5224 (N_5224,N_3028,N_2587);
nor U5225 (N_5225,N_4623,N_3702);
or U5226 (N_5226,N_4946,N_2532);
nand U5227 (N_5227,N_3518,N_3288);
or U5228 (N_5228,N_4216,N_3546);
and U5229 (N_5229,N_3009,N_3299);
and U5230 (N_5230,N_4789,N_4048);
nor U5231 (N_5231,N_3259,N_2656);
nor U5232 (N_5232,N_4752,N_4239);
nor U5233 (N_5233,N_4388,N_3274);
or U5234 (N_5234,N_3896,N_3987);
and U5235 (N_5235,N_3797,N_3073);
nand U5236 (N_5236,N_4938,N_3320);
nand U5237 (N_5237,N_3451,N_4901);
or U5238 (N_5238,N_3596,N_3045);
xor U5239 (N_5239,N_3876,N_3338);
nand U5240 (N_5240,N_4086,N_3644);
xnor U5241 (N_5241,N_4187,N_2981);
and U5242 (N_5242,N_2883,N_3721);
and U5243 (N_5243,N_2519,N_2553);
xor U5244 (N_5244,N_2880,N_4970);
or U5245 (N_5245,N_4157,N_4882);
nor U5246 (N_5246,N_4364,N_2540);
or U5247 (N_5247,N_2618,N_4655);
or U5248 (N_5248,N_3021,N_3973);
and U5249 (N_5249,N_3787,N_4830);
or U5250 (N_5250,N_4353,N_3194);
and U5251 (N_5251,N_3066,N_3301);
and U5252 (N_5252,N_3871,N_3713);
nand U5253 (N_5253,N_3817,N_3609);
nor U5254 (N_5254,N_4639,N_2936);
or U5255 (N_5255,N_4629,N_4909);
and U5256 (N_5256,N_4691,N_4450);
xnor U5257 (N_5257,N_3300,N_2655);
and U5258 (N_5258,N_3418,N_4720);
nand U5259 (N_5259,N_3832,N_3756);
nand U5260 (N_5260,N_4061,N_4916);
nand U5261 (N_5261,N_2559,N_4538);
nor U5262 (N_5262,N_3232,N_3860);
nor U5263 (N_5263,N_4855,N_3731);
nand U5264 (N_5264,N_4773,N_2955);
nor U5265 (N_5265,N_2541,N_4357);
and U5266 (N_5266,N_3247,N_4293);
nand U5267 (N_5267,N_4877,N_3950);
nand U5268 (N_5268,N_4486,N_3511);
nand U5269 (N_5269,N_4334,N_4659);
nor U5270 (N_5270,N_4367,N_3688);
or U5271 (N_5271,N_3070,N_4625);
xor U5272 (N_5272,N_4128,N_4642);
and U5273 (N_5273,N_4371,N_3033);
xor U5274 (N_5274,N_2989,N_3257);
xor U5275 (N_5275,N_2505,N_4948);
nand U5276 (N_5276,N_2888,N_3707);
and U5277 (N_5277,N_4136,N_3698);
nor U5278 (N_5278,N_3261,N_2873);
nor U5279 (N_5279,N_2925,N_4657);
xor U5280 (N_5280,N_4512,N_2896);
nand U5281 (N_5281,N_2751,N_3816);
or U5282 (N_5282,N_4199,N_4572);
and U5283 (N_5283,N_3189,N_4278);
and U5284 (N_5284,N_3084,N_3995);
xnor U5285 (N_5285,N_4442,N_3579);
xor U5286 (N_5286,N_3530,N_3098);
nand U5287 (N_5287,N_3236,N_4523);
nand U5288 (N_5288,N_4491,N_3026);
xnor U5289 (N_5289,N_4339,N_3811);
or U5290 (N_5290,N_3260,N_4513);
or U5291 (N_5291,N_3434,N_4879);
or U5292 (N_5292,N_4469,N_4687);
nor U5293 (N_5293,N_2786,N_2534);
and U5294 (N_5294,N_2872,N_2764);
nor U5295 (N_5295,N_2874,N_3216);
nand U5296 (N_5296,N_3775,N_3667);
xnor U5297 (N_5297,N_4014,N_2608);
xor U5298 (N_5298,N_4266,N_4456);
xor U5299 (N_5299,N_4996,N_3435);
or U5300 (N_5300,N_4355,N_2803);
nor U5301 (N_5301,N_3773,N_3820);
and U5302 (N_5302,N_3252,N_2965);
nand U5303 (N_5303,N_2783,N_4787);
or U5304 (N_5304,N_4306,N_4471);
or U5305 (N_5305,N_4864,N_2644);
or U5306 (N_5306,N_3672,N_4734);
xor U5307 (N_5307,N_3861,N_3740);
nor U5308 (N_5308,N_2996,N_3961);
nor U5309 (N_5309,N_3105,N_3802);
and U5310 (N_5310,N_2757,N_4228);
or U5311 (N_5311,N_4932,N_3414);
and U5312 (N_5312,N_2732,N_3751);
nand U5313 (N_5313,N_3072,N_4528);
or U5314 (N_5314,N_3834,N_3092);
nand U5315 (N_5315,N_4300,N_3282);
and U5316 (N_5316,N_2986,N_3598);
nor U5317 (N_5317,N_3494,N_3996);
nor U5318 (N_5318,N_3737,N_4033);
or U5319 (N_5319,N_3668,N_4251);
xor U5320 (N_5320,N_3639,N_3618);
or U5321 (N_5321,N_3250,N_4076);
xor U5322 (N_5322,N_2794,N_4575);
and U5323 (N_5323,N_2728,N_3465);
xnor U5324 (N_5324,N_3573,N_4229);
xor U5325 (N_5325,N_4792,N_4952);
or U5326 (N_5326,N_3280,N_3894);
xor U5327 (N_5327,N_3942,N_4784);
xor U5328 (N_5328,N_4042,N_4519);
nand U5329 (N_5329,N_3363,N_3642);
nor U5330 (N_5330,N_4884,N_2775);
nor U5331 (N_5331,N_4271,N_4870);
or U5332 (N_5332,N_4260,N_4252);
and U5333 (N_5333,N_3746,N_4881);
nand U5334 (N_5334,N_4542,N_3931);
or U5335 (N_5335,N_2584,N_3436);
nor U5336 (N_5336,N_3528,N_4430);
or U5337 (N_5337,N_4717,N_4102);
and U5338 (N_5338,N_3263,N_4120);
and U5339 (N_5339,N_2910,N_2703);
and U5340 (N_5340,N_3878,N_3638);
nand U5341 (N_5341,N_3424,N_3030);
and U5342 (N_5342,N_2518,N_4876);
nand U5343 (N_5343,N_3732,N_4092);
xnor U5344 (N_5344,N_3229,N_3023);
xor U5345 (N_5345,N_3083,N_4416);
or U5346 (N_5346,N_3237,N_3578);
nand U5347 (N_5347,N_3574,N_3091);
nor U5348 (N_5348,N_4998,N_3800);
nand U5349 (N_5349,N_3133,N_2542);
xor U5350 (N_5350,N_3555,N_3182);
and U5351 (N_5351,N_4654,N_3481);
and U5352 (N_5352,N_4517,N_3361);
nand U5353 (N_5353,N_4898,N_2769);
or U5354 (N_5354,N_3010,N_4477);
nand U5355 (N_5355,N_3919,N_3019);
nor U5356 (N_5356,N_3659,N_3572);
nand U5357 (N_5357,N_2770,N_4158);
nand U5358 (N_5358,N_2629,N_3121);
nor U5359 (N_5359,N_3457,N_3319);
nand U5360 (N_5360,N_3104,N_3352);
or U5361 (N_5361,N_4208,N_2507);
nor U5362 (N_5362,N_3427,N_4871);
xor U5363 (N_5363,N_2849,N_3770);
nand U5364 (N_5364,N_4580,N_3475);
xnor U5365 (N_5365,N_3148,N_2538);
nor U5366 (N_5366,N_4507,N_2934);
and U5367 (N_5367,N_4774,N_3482);
and U5368 (N_5368,N_4284,N_4504);
nand U5369 (N_5369,N_4354,N_4019);
nand U5370 (N_5370,N_2815,N_4445);
and U5371 (N_5371,N_4213,N_2855);
or U5372 (N_5372,N_4112,N_3576);
nand U5373 (N_5373,N_2513,N_4680);
and U5374 (N_5374,N_3411,N_3697);
and U5375 (N_5375,N_2529,N_4588);
and U5376 (N_5376,N_3538,N_4488);
or U5377 (N_5377,N_3080,N_3769);
nand U5378 (N_5378,N_2882,N_2566);
and U5379 (N_5379,N_4084,N_4713);
nor U5380 (N_5380,N_3087,N_3503);
nand U5381 (N_5381,N_3491,N_4782);
xnor U5382 (N_5382,N_4358,N_4793);
and U5383 (N_5383,N_3096,N_4980);
and U5384 (N_5384,N_3859,N_3227);
nor U5385 (N_5385,N_4452,N_4037);
and U5386 (N_5386,N_4663,N_2980);
and U5387 (N_5387,N_3267,N_4904);
or U5388 (N_5388,N_4443,N_4925);
nand U5389 (N_5389,N_3330,N_2556);
nor U5390 (N_5390,N_3917,N_3502);
and U5391 (N_5391,N_4729,N_3733);
nand U5392 (N_5392,N_3239,N_2787);
nand U5393 (N_5393,N_2778,N_2909);
nand U5394 (N_5394,N_4558,N_3225);
xnor U5395 (N_5395,N_4074,N_3637);
and U5396 (N_5396,N_2845,N_4997);
or U5397 (N_5397,N_4108,N_4298);
nand U5398 (N_5398,N_3492,N_3868);
nor U5399 (N_5399,N_3649,N_2834);
nand U5400 (N_5400,N_3040,N_4719);
and U5401 (N_5401,N_3449,N_3420);
xnor U5402 (N_5402,N_4280,N_4258);
nor U5403 (N_5403,N_4622,N_4724);
nor U5404 (N_5404,N_4093,N_3195);
and U5405 (N_5405,N_4710,N_4344);
nand U5406 (N_5406,N_4978,N_4832);
nor U5407 (N_5407,N_3113,N_2717);
or U5408 (N_5408,N_2806,N_3162);
nor U5409 (N_5409,N_3514,N_2831);
nand U5410 (N_5410,N_3377,N_2726);
nand U5411 (N_5411,N_3017,N_4246);
nor U5412 (N_5412,N_2710,N_3253);
nand U5413 (N_5413,N_3067,N_3628);
xor U5414 (N_5414,N_2939,N_3214);
or U5415 (N_5415,N_4801,N_4276);
xor U5416 (N_5416,N_4966,N_4705);
nand U5417 (N_5417,N_4960,N_3468);
xnor U5418 (N_5418,N_3281,N_3336);
xor U5419 (N_5419,N_4738,N_4972);
nor U5420 (N_5420,N_2842,N_3368);
nor U5421 (N_5421,N_2857,N_4404);
nand U5422 (N_5422,N_3662,N_3969);
nand U5423 (N_5423,N_2678,N_4257);
or U5424 (N_5424,N_3399,N_3085);
nor U5425 (N_5425,N_4378,N_3378);
or U5426 (N_5426,N_3674,N_3012);
nor U5427 (N_5427,N_2760,N_4492);
or U5428 (N_5428,N_2755,N_3241);
and U5429 (N_5429,N_2899,N_3825);
or U5430 (N_5430,N_4689,N_3297);
or U5431 (N_5431,N_4731,N_4921);
and U5432 (N_5432,N_2666,N_3185);
nand U5433 (N_5433,N_4988,N_3870);
xor U5434 (N_5434,N_3140,N_2879);
xor U5435 (N_5435,N_4577,N_4824);
nand U5436 (N_5436,N_2761,N_2707);
nand U5437 (N_5437,N_2690,N_4820);
and U5438 (N_5438,N_4924,N_3723);
nand U5439 (N_5439,N_3665,N_3313);
and U5440 (N_5440,N_4139,N_3130);
and U5441 (N_5441,N_3188,N_4950);
nor U5442 (N_5442,N_3522,N_4233);
xor U5443 (N_5443,N_4923,N_4069);
nand U5444 (N_5444,N_3355,N_4302);
nor U5445 (N_5445,N_4060,N_2887);
nand U5446 (N_5446,N_4054,N_2968);
or U5447 (N_5447,N_4016,N_3956);
xnor U5448 (N_5448,N_4886,N_2854);
xor U5449 (N_5449,N_4733,N_4123);
and U5450 (N_5450,N_4791,N_4017);
or U5451 (N_5451,N_2801,N_3829);
or U5452 (N_5452,N_4317,N_2863);
xnor U5453 (N_5453,N_3477,N_2781);
nand U5454 (N_5454,N_2607,N_4833);
or U5455 (N_5455,N_2784,N_4420);
nor U5456 (N_5456,N_2841,N_3897);
nand U5457 (N_5457,N_2738,N_2592);
xor U5458 (N_5458,N_4845,N_3714);
and U5459 (N_5459,N_3478,N_4160);
xnor U5460 (N_5460,N_3218,N_3542);
and U5461 (N_5461,N_3032,N_2602);
and U5462 (N_5462,N_3170,N_3126);
xor U5463 (N_5463,N_4197,N_4406);
and U5464 (N_5464,N_4514,N_2881);
nand U5465 (N_5465,N_4458,N_2702);
nand U5466 (N_5466,N_3342,N_4299);
nor U5467 (N_5467,N_2611,N_4180);
or U5468 (N_5468,N_3554,N_4351);
nor U5469 (N_5469,N_3137,N_3244);
nand U5470 (N_5470,N_3582,N_2953);
or U5471 (N_5471,N_2823,N_2992);
and U5472 (N_5472,N_3607,N_3163);
nor U5473 (N_5473,N_3142,N_4583);
nand U5474 (N_5474,N_3544,N_3959);
and U5475 (N_5475,N_4638,N_3461);
xnor U5476 (N_5476,N_4343,N_3110);
or U5477 (N_5477,N_3082,N_2999);
and U5478 (N_5478,N_2916,N_4097);
xnor U5479 (N_5479,N_4002,N_4453);
or U5480 (N_5480,N_3184,N_2683);
nand U5481 (N_5481,N_4277,N_4332);
xor U5482 (N_5482,N_3922,N_2645);
or U5483 (N_5483,N_2906,N_3957);
nand U5484 (N_5484,N_2904,N_3968);
or U5485 (N_5485,N_3328,N_4460);
xor U5486 (N_5486,N_4764,N_4392);
xor U5487 (N_5487,N_4854,N_3437);
or U5488 (N_5488,N_4677,N_3074);
nand U5489 (N_5489,N_3439,N_4541);
xor U5490 (N_5490,N_2829,N_4152);
or U5491 (N_5491,N_4326,N_2744);
nand U5492 (N_5492,N_3595,N_4030);
xnor U5493 (N_5493,N_4963,N_4800);
xnor U5494 (N_5494,N_2533,N_4674);
nand U5495 (N_5495,N_3994,N_3285);
or U5496 (N_5496,N_4329,N_4892);
nor U5497 (N_5497,N_4324,N_3308);
or U5498 (N_5498,N_2709,N_4759);
nand U5499 (N_5499,N_3102,N_3734);
nand U5500 (N_5500,N_3660,N_4011);
and U5501 (N_5501,N_3100,N_4262);
nor U5502 (N_5502,N_4941,N_2635);
and U5503 (N_5503,N_2727,N_4672);
and U5504 (N_5504,N_4737,N_4912);
nand U5505 (N_5505,N_2895,N_3520);
and U5506 (N_5506,N_3531,N_4221);
nand U5507 (N_5507,N_3201,N_3068);
nand U5508 (N_5508,N_4169,N_4761);
nand U5509 (N_5509,N_3276,N_3423);
nand U5510 (N_5510,N_4018,N_3046);
or U5511 (N_5511,N_2753,N_2643);
nor U5512 (N_5512,N_4846,N_3381);
nand U5513 (N_5513,N_2959,N_4062);
nor U5514 (N_5514,N_2501,N_2640);
and U5515 (N_5515,N_2698,N_4653);
nand U5516 (N_5516,N_3408,N_4150);
nor U5517 (N_5517,N_4554,N_3443);
or U5518 (N_5518,N_2637,N_2554);
nor U5519 (N_5519,N_3898,N_3001);
nand U5520 (N_5520,N_4396,N_3305);
or U5521 (N_5521,N_4254,N_3421);
nor U5522 (N_5522,N_3921,N_4359);
nand U5523 (N_5523,N_4915,N_3814);
nand U5524 (N_5524,N_4220,N_3772);
nor U5525 (N_5525,N_3278,N_3173);
nand U5526 (N_5526,N_3426,N_3675);
nand U5527 (N_5527,N_3099,N_3134);
nor U5528 (N_5528,N_2884,N_2835);
nand U5529 (N_5529,N_3193,N_4853);
or U5530 (N_5530,N_3647,N_2822);
xnor U5531 (N_5531,N_2522,N_2756);
or U5532 (N_5532,N_3882,N_4373);
xor U5533 (N_5533,N_3955,N_4098);
xnor U5534 (N_5534,N_3387,N_3784);
xnor U5535 (N_5535,N_3630,N_2562);
nor U5536 (N_5536,N_4106,N_3374);
xor U5537 (N_5537,N_4498,N_3177);
and U5538 (N_5538,N_4318,N_3622);
nor U5539 (N_5539,N_2998,N_2682);
nand U5540 (N_5540,N_3619,N_3985);
nor U5541 (N_5541,N_4099,N_4807);
or U5542 (N_5542,N_2837,N_2604);
nand U5543 (N_5543,N_3485,N_4698);
or U5544 (N_5544,N_4043,N_3928);
or U5545 (N_5545,N_4255,N_4990);
nand U5546 (N_5546,N_4750,N_3958);
nand U5547 (N_5547,N_3801,N_4237);
xor U5548 (N_5548,N_3212,N_4567);
nor U5549 (N_5549,N_4168,N_3873);
and U5550 (N_5550,N_4338,N_3681);
xor U5551 (N_5551,N_3833,N_3690);
nor U5552 (N_5552,N_2609,N_3060);
or U5553 (N_5553,N_4346,N_3534);
or U5554 (N_5554,N_3999,N_3366);
and U5555 (N_5555,N_4796,N_4314);
nand U5556 (N_5556,N_3535,N_3608);
nand U5557 (N_5557,N_4408,N_3742);
or U5558 (N_5558,N_4728,N_2701);
nand U5559 (N_5559,N_3112,N_3016);
nand U5560 (N_5560,N_4770,N_3744);
xnor U5561 (N_5561,N_2827,N_2589);
and U5562 (N_5562,N_4143,N_2771);
nand U5563 (N_5563,N_4826,N_3900);
nor U5564 (N_5564,N_4788,N_3386);
and U5565 (N_5565,N_3223,N_4849);
nor U5566 (N_5566,N_3516,N_3262);
nor U5567 (N_5567,N_4985,N_3965);
and U5568 (N_5568,N_4578,N_2870);
xor U5569 (N_5569,N_3933,N_3786);
xor U5570 (N_5570,N_3487,N_3264);
xor U5571 (N_5571,N_4363,N_3390);
and U5572 (N_5572,N_4887,N_2731);
nand U5573 (N_5573,N_2733,N_4762);
nand U5574 (N_5574,N_4001,N_4413);
xnor U5575 (N_5575,N_4847,N_4560);
nor U5576 (N_5576,N_3095,N_3627);
and U5577 (N_5577,N_4195,N_4207);
or U5578 (N_5578,N_3726,N_3277);
xor U5579 (N_5579,N_2578,N_3293);
nand U5580 (N_5580,N_2748,N_2649);
and U5581 (N_5581,N_4115,N_2991);
nor U5582 (N_5582,N_3107,N_4865);
xnor U5583 (N_5583,N_4171,N_3272);
nor U5584 (N_5584,N_2721,N_4806);
xor U5585 (N_5585,N_3614,N_4756);
and U5586 (N_5586,N_4073,N_4447);
or U5587 (N_5587,N_3739,N_2521);
nor U5588 (N_5588,N_3908,N_3828);
or U5589 (N_5589,N_4595,N_2850);
nor U5590 (N_5590,N_3446,N_4117);
nand U5591 (N_5591,N_4417,N_3857);
and U5592 (N_5592,N_2878,N_3200);
and U5593 (N_5593,N_4867,N_4911);
nand U5594 (N_5594,N_4621,N_3512);
or U5595 (N_5595,N_4684,N_4602);
nor U5596 (N_5596,N_4089,N_3118);
and U5597 (N_5597,N_3550,N_3720);
and U5598 (N_5598,N_2724,N_3348);
or U5599 (N_5599,N_4984,N_4297);
xnor U5600 (N_5600,N_4863,N_2563);
and U5601 (N_5601,N_4751,N_2869);
nand U5602 (N_5602,N_4476,N_3926);
and U5603 (N_5603,N_2759,N_3120);
or U5604 (N_5604,N_3709,N_2877);
nand U5605 (N_5605,N_3699,N_2838);
and U5606 (N_5606,N_3899,N_4272);
nand U5607 (N_5607,N_4485,N_3903);
nand U5608 (N_5608,N_2798,N_3767);
and U5609 (N_5609,N_4064,N_4785);
nor U5610 (N_5610,N_4039,N_3565);
xor U5611 (N_5611,N_2741,N_3589);
xnor U5612 (N_5612,N_4975,N_4475);
and U5613 (N_5613,N_3271,N_4451);
and U5614 (N_5614,N_4473,N_3693);
xor U5615 (N_5615,N_2921,N_3924);
or U5616 (N_5616,N_2919,N_4530);
nand U5617 (N_5617,N_4244,N_4522);
nand U5618 (N_5618,N_3620,N_4340);
xnor U5619 (N_5619,N_4574,N_3116);
or U5620 (N_5620,N_4636,N_2614);
nand U5621 (N_5621,N_2848,N_3490);
or U5622 (N_5622,N_4415,N_4702);
nor U5623 (N_5623,N_4555,N_3419);
and U5624 (N_5624,N_4926,N_3966);
and U5625 (N_5625,N_4612,N_4670);
and U5626 (N_5626,N_4914,N_3631);
nand U5627 (N_5627,N_3486,N_4489);
xor U5628 (N_5628,N_4540,N_4585);
or U5629 (N_5629,N_4741,N_3076);
nor U5630 (N_5630,N_4403,N_4440);
or U5631 (N_5631,N_4381,N_4107);
nand U5632 (N_5632,N_2606,N_2596);
nand U5633 (N_5633,N_4243,N_2572);
nor U5634 (N_5634,N_4281,N_3109);
xnor U5635 (N_5635,N_2612,N_4402);
and U5636 (N_5636,N_3450,N_4163);
nor U5637 (N_5637,N_4532,N_4533);
nor U5638 (N_5638,N_4814,N_3577);
or U5639 (N_5639,N_3054,N_3284);
xnor U5640 (N_5640,N_3846,N_2898);
xor U5641 (N_5641,N_4976,N_3013);
and U5642 (N_5642,N_3643,N_3907);
and U5643 (N_5643,N_2673,N_3507);
nand U5644 (N_5644,N_3139,N_4225);
and U5645 (N_5645,N_4444,N_3600);
or U5646 (N_5646,N_4497,N_3914);
nor U5647 (N_5647,N_3838,N_3174);
xnor U5648 (N_5648,N_4186,N_2508);
and U5649 (N_5649,N_2890,N_2546);
and U5650 (N_5650,N_4431,N_3329);
nand U5651 (N_5651,N_3323,N_3206);
nand U5652 (N_5652,N_2659,N_4837);
nor U5653 (N_5653,N_3934,N_3616);
nor U5654 (N_5654,N_3989,N_4055);
and U5655 (N_5655,N_2502,N_4352);
nand U5656 (N_5656,N_4405,N_4885);
or U5657 (N_5657,N_3763,N_3160);
xnor U5658 (N_5658,N_3849,N_2820);
nand U5659 (N_5659,N_3822,N_4977);
and U5660 (N_5660,N_3654,N_3360);
or U5661 (N_5661,N_4215,N_4161);
xnor U5662 (N_5662,N_4979,N_2623);
nand U5663 (N_5663,N_2653,N_2817);
nand U5664 (N_5664,N_4303,N_4760);
or U5665 (N_5665,N_3458,N_4662);
nand U5666 (N_5666,N_3215,N_4715);
nand U5667 (N_5667,N_4579,N_2967);
nor U5668 (N_5668,N_3393,N_2544);
and U5669 (N_5669,N_3762,N_4131);
or U5670 (N_5670,N_4137,N_3000);
or U5671 (N_5671,N_4521,N_3441);
nand U5672 (N_5672,N_2651,N_3691);
nor U5673 (N_5673,N_4418,N_4046);
nand U5674 (N_5674,N_4337,N_4474);
nor U5675 (N_5675,N_3304,N_4087);
xor U5676 (N_5676,N_3132,N_3587);
or U5677 (N_5677,N_3243,N_3658);
nor U5678 (N_5678,N_3915,N_4549);
and U5679 (N_5679,N_2695,N_3447);
nor U5680 (N_5680,N_4908,N_3135);
nand U5681 (N_5681,N_2780,N_3761);
or U5682 (N_5682,N_3416,N_3428);
or U5683 (N_5683,N_2933,N_3410);
nor U5684 (N_5684,N_3312,N_4502);
nor U5685 (N_5685,N_4958,N_2931);
or U5686 (N_5686,N_2975,N_3504);
or U5687 (N_5687,N_2735,N_3911);
nor U5688 (N_5688,N_4435,N_2641);
nand U5689 (N_5689,N_4259,N_4464);
xor U5690 (N_5690,N_4190,N_4209);
or U5691 (N_5691,N_4114,N_2579);
and U5692 (N_5692,N_4576,N_2693);
and U5693 (N_5693,N_2983,N_4628);
and U5694 (N_5694,N_4472,N_4518);
nand U5695 (N_5695,N_4088,N_4548);
nor U5696 (N_5696,N_4856,N_2892);
or U5697 (N_5697,N_3935,N_4748);
nor U5698 (N_5698,N_4561,N_4394);
nand U5699 (N_5699,N_2912,N_3069);
nand U5700 (N_5700,N_2689,N_3115);
xor U5701 (N_5701,N_2730,N_4372);
or U5702 (N_5702,N_2993,N_3413);
xor U5703 (N_5703,N_4240,N_2763);
nor U5704 (N_5704,N_4040,N_3677);
nor U5705 (N_5705,N_3796,N_3729);
nand U5706 (N_5706,N_4265,N_4015);
xnor U5707 (N_5707,N_3855,N_3382);
or U5708 (N_5708,N_3990,N_4875);
xor U5709 (N_5709,N_4632,N_4964);
and U5710 (N_5710,N_3890,N_4232);
nand U5711 (N_5711,N_3398,N_4330);
nand U5712 (N_5712,N_4428,N_4003);
xnor U5713 (N_5713,N_3954,N_3610);
nor U5714 (N_5714,N_3240,N_4174);
and U5715 (N_5715,N_4130,N_2908);
nand U5716 (N_5716,N_4210,N_2809);
nor U5717 (N_5717,N_4962,N_4110);
and U5718 (N_5718,N_4414,N_3929);
and U5719 (N_5719,N_3711,N_4028);
xnor U5720 (N_5720,N_4973,N_3551);
nor U5721 (N_5721,N_3079,N_4129);
nand U5722 (N_5722,N_3422,N_2765);
and U5723 (N_5723,N_2742,N_2774);
nor U5724 (N_5724,N_3559,N_4605);
or U5725 (N_5725,N_3728,N_2813);
and U5726 (N_5726,N_3676,N_3840);
xnor U5727 (N_5727,N_4866,N_4696);
and U5728 (N_5728,N_3187,N_2927);
nor U5729 (N_5729,N_4176,N_2598);
nor U5730 (N_5730,N_3863,N_3799);
and U5731 (N_5731,N_4899,N_3008);
or U5732 (N_5732,N_3540,N_2705);
and U5733 (N_5733,N_4714,N_4900);
xor U5734 (N_5734,N_3581,N_3402);
or U5735 (N_5735,N_3790,N_3479);
xnor U5736 (N_5736,N_3710,N_3851);
and U5737 (N_5737,N_2960,N_3056);
nor U5738 (N_5738,N_4678,N_4983);
or U5739 (N_5739,N_4619,N_4395);
nor U5740 (N_5740,N_3523,N_4603);
nand U5741 (N_5741,N_3590,N_4119);
nand U5742 (N_5742,N_3347,N_3233);
nand U5743 (N_5743,N_3031,N_2548);
nor U5744 (N_5744,N_4328,N_4676);
nand U5745 (N_5745,N_3725,N_2560);
and U5746 (N_5746,N_4267,N_4604);
and U5747 (N_5747,N_2528,N_4036);
or U5748 (N_5748,N_3835,N_4669);
xnor U5749 (N_5749,N_3650,N_3708);
or U5750 (N_5750,N_3208,N_4695);
nor U5751 (N_5751,N_3552,N_3444);
nor U5752 (N_5752,N_4376,N_4026);
nor U5753 (N_5753,N_4090,N_4173);
or U5754 (N_5754,N_3108,N_4104);
and U5755 (N_5755,N_4004,N_3902);
or U5756 (N_5756,N_2804,N_3783);
nor U5757 (N_5757,N_3656,N_2825);
nand U5758 (N_5758,N_4134,N_3041);
nand U5759 (N_5759,N_4024,N_4310);
or U5760 (N_5760,N_2558,N_2962);
nand U5761 (N_5761,N_4590,N_4361);
or U5762 (N_5762,N_4223,N_2570);
xor U5763 (N_5763,N_2946,N_2520);
and U5764 (N_5764,N_3852,N_4516);
and U5765 (N_5765,N_2639,N_4391);
nor U5766 (N_5766,N_4247,N_4701);
nand U5767 (N_5767,N_3891,N_3238);
or U5768 (N_5768,N_2687,N_3412);
nor U5769 (N_5769,N_3375,N_4455);
nand U5770 (N_5770,N_4167,N_3178);
nor U5771 (N_5771,N_4842,N_4484);
nor U5772 (N_5772,N_2847,N_4231);
or U5773 (N_5773,N_4079,N_3695);
nand U5774 (N_5774,N_3509,N_3625);
and U5775 (N_5775,N_2638,N_3670);
or U5776 (N_5776,N_3663,N_3745);
or U5777 (N_5777,N_3251,N_3495);
and U5778 (N_5778,N_4461,N_4601);
or U5779 (N_5779,N_4013,N_3505);
xor U5780 (N_5780,N_3078,N_3515);
nor U5781 (N_5781,N_2723,N_4971);
nand U5782 (N_5782,N_2715,N_3634);
or U5783 (N_5783,N_4943,N_3562);
and U5784 (N_5784,N_3460,N_2720);
nand U5785 (N_5785,N_4327,N_3593);
nand U5786 (N_5786,N_2902,N_4311);
or U5787 (N_5787,N_3768,N_2990);
or U5788 (N_5788,N_4508,N_4068);
xnor U5789 (N_5789,N_3821,N_3292);
xor U5790 (N_5790,N_4529,N_3196);
nand U5791 (N_5791,N_4758,N_3175);
nor U5792 (N_5792,N_3024,N_2537);
nand U5793 (N_5793,N_4172,N_3127);
and U5794 (N_5794,N_2585,N_4931);
or U5795 (N_5795,N_4308,N_3379);
nand U5796 (N_5796,N_4175,N_3570);
or U5797 (N_5797,N_3442,N_2633);
xor U5798 (N_5798,N_4614,N_3705);
and U5799 (N_5799,N_3776,N_4360);
xor U5800 (N_5800,N_3372,N_2843);
or U5801 (N_5801,N_4424,N_3350);
nand U5802 (N_5802,N_2832,N_3417);
and U5803 (N_5803,N_4571,N_4049);
nor U5804 (N_5804,N_2777,N_3785);
or U5805 (N_5805,N_4766,N_3886);
or U5806 (N_5806,N_4007,N_4640);
or U5807 (N_5807,N_3553,N_3937);
or U5808 (N_5808,N_4666,N_3269);
nand U5809 (N_5809,N_3129,N_4775);
or U5810 (N_5810,N_3433,N_4797);
nor U5811 (N_5811,N_3406,N_2582);
nand U5812 (N_5812,N_3141,N_4757);
or U5813 (N_5813,N_4673,N_2597);
and U5814 (N_5814,N_2800,N_3053);
nand U5815 (N_5815,N_2500,N_3058);
xor U5816 (N_5816,N_2846,N_4798);
or U5817 (N_5817,N_4992,N_2964);
xor U5818 (N_5818,N_3778,N_4598);
and U5819 (N_5819,N_4145,N_4515);
nand U5820 (N_5820,N_3741,N_3463);
or U5821 (N_5821,N_4083,N_4309);
nor U5822 (N_5822,N_4819,N_4697);
and U5823 (N_5823,N_2802,N_2646);
nor U5824 (N_5824,N_4188,N_3469);
or U5825 (N_5825,N_3621,N_4465);
or U5826 (N_5826,N_3754,N_4811);
nand U5827 (N_5827,N_2808,N_2963);
or U5828 (N_5828,N_4335,N_4565);
nand U5829 (N_5829,N_2995,N_4816);
nor U5830 (N_5830,N_2970,N_4989);
nor U5831 (N_5831,N_4109,N_3210);
and U5832 (N_5832,N_4133,N_4425);
nor U5833 (N_5833,N_2875,N_4616);
nand U5834 (N_5834,N_4142,N_4006);
nand U5835 (N_5835,N_2739,N_4951);
and U5836 (N_5836,N_4611,N_4345);
nor U5837 (N_5837,N_3226,N_3636);
nor U5838 (N_5838,N_4227,N_3022);
nand U5839 (N_5839,N_2658,N_3563);
nor U5840 (N_5840,N_4805,N_3357);
or U5841 (N_5841,N_4880,N_2889);
nand U5842 (N_5842,N_3601,N_3548);
nor U5843 (N_5843,N_4947,N_3004);
and U5844 (N_5844,N_3202,N_3474);
nor U5845 (N_5845,N_2669,N_4776);
nor U5846 (N_5846,N_2971,N_2661);
nor U5847 (N_5847,N_2826,N_4597);
nor U5848 (N_5848,N_3747,N_3462);
nor U5849 (N_5849,N_2905,N_4954);
xnor U5850 (N_5850,N_3736,N_3883);
and U5851 (N_5851,N_3327,N_2767);
and U5852 (N_5852,N_4956,N_2754);
xor U5853 (N_5853,N_2779,N_4537);
nor U5854 (N_5854,N_3568,N_3818);
or U5855 (N_5855,N_2591,N_3920);
xnor U5856 (N_5856,N_4929,N_3089);
xor U5857 (N_5857,N_4056,N_4671);
or U5858 (N_5858,N_4894,N_4872);
nand U5859 (N_5859,N_4768,N_4543);
and U5860 (N_5860,N_3047,N_4682);
nor U5861 (N_5861,N_4675,N_2657);
nor U5862 (N_5862,N_3205,N_4645);
nand U5863 (N_5863,N_2950,N_4905);
or U5864 (N_5864,N_4285,N_3199);
nor U5865 (N_5865,N_2947,N_4483);
xnor U5866 (N_5866,N_4294,N_3635);
nand U5867 (N_5867,N_4331,N_3764);
or U5868 (N_5868,N_3604,N_3962);
nand U5869 (N_5869,N_4370,N_4790);
xnor U5870 (N_5870,N_4375,N_3149);
and U5871 (N_5871,N_2749,N_4304);
or U5872 (N_5872,N_2922,N_4934);
or U5873 (N_5873,N_3722,N_4051);
nand U5874 (N_5874,N_3782,N_2914);
xor U5875 (N_5875,N_4082,N_4559);
and U5876 (N_5876,N_4463,N_4292);
nand U5877 (N_5877,N_3944,N_4919);
or U5878 (N_5878,N_4744,N_3683);
nor U5879 (N_5879,N_2600,N_3044);
nand U5880 (N_5880,N_4591,N_2768);
nand U5881 (N_5881,N_3750,N_3584);
and U5882 (N_5882,N_3266,N_2812);
and U5883 (N_5883,N_4005,N_4374);
and U5884 (N_5884,N_2509,N_3606);
nand U5885 (N_5885,N_3564,N_4825);
xor U5886 (N_5886,N_3077,N_2737);
nor U5887 (N_5887,N_3866,N_2706);
nand U5888 (N_5888,N_4961,N_4116);
and U5889 (N_5889,N_3760,N_4245);
nor U5890 (N_5890,N_4686,N_3152);
and U5891 (N_5891,N_3249,N_4103);
xnor U5892 (N_5892,N_4429,N_2714);
nor U5893 (N_5893,N_2506,N_4889);
nor U5894 (N_5894,N_3940,N_4050);
nor U5895 (N_5895,N_3114,N_3326);
xnor U5896 (N_5896,N_2663,N_3065);
nor U5897 (N_5897,N_3837,N_2833);
and U5898 (N_5898,N_4995,N_4287);
or U5899 (N_5899,N_4058,N_3176);
and U5900 (N_5900,N_2867,N_4147);
nor U5901 (N_5901,N_4126,N_4348);
xor U5902 (N_5902,N_3795,N_2818);
and U5903 (N_5903,N_4706,N_3038);
and U5904 (N_5904,N_3766,N_4301);
or U5905 (N_5905,N_2976,N_4384);
or U5906 (N_5906,N_3939,N_3051);
xnor U5907 (N_5907,N_3848,N_3524);
or U5908 (N_5908,N_3824,N_2564);
nand U5909 (N_5909,N_2911,N_3310);
and U5910 (N_5910,N_3971,N_2913);
xnor U5911 (N_5911,N_4703,N_3367);
nor U5912 (N_5912,N_4286,N_3345);
nor U5913 (N_5913,N_3560,N_2858);
nor U5914 (N_5914,N_3164,N_3498);
or U5915 (N_5915,N_3483,N_3043);
and U5916 (N_5916,N_4735,N_3689);
nor U5917 (N_5917,N_3879,N_3369);
xor U5918 (N_5918,N_3998,N_4347);
nand U5919 (N_5919,N_2859,N_4587);
nand U5920 (N_5920,N_3383,N_3124);
and U5921 (N_5921,N_4462,N_4009);
and U5922 (N_5922,N_3125,N_4634);
nand U5923 (N_5923,N_4021,N_4610);
or U5924 (N_5924,N_3603,N_2634);
nor U5925 (N_5925,N_2788,N_4815);
and U5926 (N_5926,N_3384,N_3050);
and U5927 (N_5927,N_3700,N_3151);
and U5928 (N_5928,N_2856,N_4080);
or U5929 (N_5929,N_2593,N_4419);
nand U5930 (N_5930,N_4562,N_4291);
nand U5931 (N_5931,N_4198,N_4564);
nor U5932 (N_5932,N_4500,N_4809);
nand U5933 (N_5933,N_3575,N_3946);
and U5934 (N_5934,N_2642,N_4688);
nand U5935 (N_5935,N_3397,N_4181);
nor U5936 (N_5936,N_4936,N_2985);
or U5937 (N_5937,N_3351,N_4273);
nand U5938 (N_5938,N_2543,N_3519);
or U5939 (N_5939,N_4289,N_4421);
or U5940 (N_5940,N_3980,N_2853);
nand U5941 (N_5941,N_4794,N_3812);
or U5942 (N_5942,N_3932,N_3830);
or U5943 (N_5943,N_3484,N_3623);
and U5944 (N_5944,N_2525,N_3343);
nor U5945 (N_5945,N_4182,N_3154);
or U5946 (N_5946,N_3166,N_4235);
or U5947 (N_5947,N_4312,N_4968);
nand U5948 (N_5948,N_2691,N_3346);
nor U5949 (N_5949,N_2551,N_2557);
and U5950 (N_5950,N_2894,N_4868);
and U5951 (N_5951,N_3143,N_2652);
xnor U5952 (N_5952,N_4897,N_3682);
xor U5953 (N_5953,N_3268,N_3472);
nor U5954 (N_5954,N_3906,N_4448);
nor U5955 (N_5955,N_3602,N_3703);
and U5956 (N_5956,N_3448,N_2944);
or U5957 (N_5957,N_4032,N_4930);
and U5958 (N_5958,N_4643,N_3901);
xor U5959 (N_5959,N_4953,N_2547);
xor U5960 (N_5960,N_4895,N_4994);
or U5961 (N_5961,N_4813,N_2511);
xor U5962 (N_5962,N_4315,N_2974);
or U5963 (N_5963,N_3476,N_2648);
xor U5964 (N_5964,N_4362,N_3806);
or U5965 (N_5965,N_2515,N_4493);
and U5966 (N_5966,N_3537,N_4307);
nand U5967 (N_5967,N_3005,N_4349);
nand U5968 (N_5968,N_4165,N_3165);
nand U5969 (N_5969,N_4248,N_3209);
nand U5970 (N_5970,N_3952,N_4627);
nand U5971 (N_5971,N_3035,N_3791);
nor U5972 (N_5972,N_4679,N_3286);
nor U5973 (N_5973,N_4179,N_4454);
or U5974 (N_5974,N_3167,N_2595);
xnor U5975 (N_5975,N_4573,N_4608);
xnor U5976 (N_5976,N_4836,N_2790);
and U5977 (N_5977,N_3432,N_4178);
nor U5978 (N_5978,N_4212,N_2504);
and U5979 (N_5979,N_2977,N_3545);
or U5980 (N_5980,N_2674,N_4437);
or U5981 (N_5981,N_4279,N_4217);
xor U5982 (N_5982,N_2792,N_3344);
nor U5983 (N_5983,N_3633,N_4387);
and U5984 (N_5984,N_3986,N_4539);
xor U5985 (N_5985,N_3015,N_3388);
and U5986 (N_5986,N_3669,N_2632);
nor U5987 (N_5987,N_4778,N_4236);
nor U5988 (N_5988,N_2719,N_2821);
or U5989 (N_5989,N_4873,N_3712);
or U5990 (N_5990,N_3991,N_2932);
nand U5991 (N_5991,N_4124,N_3157);
xor U5992 (N_5992,N_3283,N_3875);
nor U5993 (N_5993,N_2851,N_3318);
and U5994 (N_5994,N_3403,N_3793);
or U5995 (N_5995,N_3147,N_4711);
or U5996 (N_5996,N_3029,N_4196);
and U5997 (N_5997,N_4263,N_4874);
nor U5998 (N_5998,N_3794,N_4035);
and U5999 (N_5999,N_2745,N_2807);
and U6000 (N_6000,N_3296,N_3011);
nand U6001 (N_6001,N_3186,N_3404);
and U6002 (N_6002,N_4848,N_3557);
xnor U6003 (N_6003,N_4843,N_3466);
nand U6004 (N_6004,N_3385,N_4907);
nand U6005 (N_6005,N_3813,N_4780);
or U6006 (N_6006,N_3171,N_4933);
nand U6007 (N_6007,N_4487,N_4546);
and U6008 (N_6008,N_3322,N_4660);
nor U6009 (N_6009,N_3452,N_3231);
xor U6010 (N_6010,N_4633,N_3303);
xor U6011 (N_6011,N_2920,N_2924);
and U6012 (N_6012,N_3081,N_4827);
and U6013 (N_6013,N_3704,N_3356);
or U6014 (N_6014,N_2512,N_2696);
nand U6015 (N_6015,N_3370,N_4275);
or U6016 (N_6016,N_4582,N_3539);
and U6017 (N_6017,N_3230,N_4020);
or U6018 (N_6018,N_4839,N_4651);
or U6019 (N_6019,N_3599,N_2773);
nor U6020 (N_6020,N_3945,N_4393);
nand U6021 (N_6021,N_4138,N_4747);
xnor U6022 (N_6022,N_3592,N_3431);
and U6023 (N_6023,N_4841,N_4503);
nand U6024 (N_6024,N_3706,N_4646);
or U6025 (N_6025,N_3279,N_3805);
nor U6026 (N_6026,N_4478,N_3779);
xor U6027 (N_6027,N_2684,N_3941);
and U6028 (N_6028,N_4615,N_4991);
and U6029 (N_6029,N_4261,N_3979);
and U6030 (N_6030,N_4891,N_4641);
xor U6031 (N_6031,N_4242,N_2622);
and U6032 (N_6032,N_2746,N_3753);
nor U6033 (N_6033,N_3809,N_4681);
or U6034 (N_6034,N_4397,N_4398);
and U6035 (N_6035,N_2624,N_4156);
xnor U6036 (N_6036,N_4928,N_3316);
and U6037 (N_6037,N_3752,N_3119);
nor U6038 (N_6038,N_2987,N_2758);
nand U6039 (N_6039,N_4594,N_2523);
and U6040 (N_6040,N_3872,N_4468);
xor U6041 (N_6041,N_2797,N_2805);
and U6042 (N_6042,N_4342,N_4193);
and U6043 (N_6043,N_3306,N_3245);
or U6044 (N_6044,N_3445,N_3567);
or U6045 (N_6045,N_4850,N_3645);
nand U6046 (N_6046,N_4113,N_2743);
nand U6047 (N_6047,N_3158,N_3341);
or U6048 (N_6048,N_4739,N_3845);
nand U6049 (N_6049,N_3585,N_3807);
xnor U6050 (N_6050,N_4012,N_3850);
and U6051 (N_6051,N_2552,N_4617);
nand U6052 (N_6052,N_4704,N_4606);
nor U6053 (N_6053,N_2628,N_4861);
xnor U6054 (N_6054,N_3664,N_2692);
nand U6055 (N_6055,N_3561,N_3128);
xor U6056 (N_6056,N_3287,N_4743);
nor U6057 (N_6057,N_3981,N_4644);
xor U6058 (N_6058,N_4122,N_3438);
nor U6059 (N_6059,N_4736,N_3533);
and U6060 (N_6060,N_2866,N_3765);
xnor U6061 (N_6061,N_2567,N_2943);
xor U6062 (N_6062,N_2937,N_3376);
xor U6063 (N_6063,N_4205,N_4127);
or U6064 (N_6064,N_4531,N_3856);
and U6065 (N_6065,N_3976,N_3464);
nor U6066 (N_6066,N_2871,N_3489);
or U6067 (N_6067,N_3982,N_3425);
nor U6068 (N_6068,N_4955,N_4065);
nand U6069 (N_6069,N_2772,N_4534);
or U6070 (N_6070,N_4322,N_3224);
and U6071 (N_6071,N_2712,N_3594);
or U6072 (N_6072,N_3529,N_4544);
nand U6073 (N_6073,N_3925,N_3936);
xnor U6074 (N_6074,N_2885,N_2700);
and U6075 (N_6075,N_4031,N_3571);
nor U6076 (N_6076,N_4828,N_4177);
and U6077 (N_6077,N_3358,N_4434);
xnor U6078 (N_6078,N_4323,N_3365);
xnor U6079 (N_6079,N_4786,N_4234);
nor U6080 (N_6080,N_4723,N_2718);
and U6081 (N_6081,N_4230,N_2555);
or U6082 (N_6082,N_2886,N_3337);
nand U6083 (N_6083,N_4584,N_3359);
or U6084 (N_6084,N_2550,N_2972);
xnor U6085 (N_6085,N_3527,N_3827);
nor U6086 (N_6086,N_4010,N_3333);
nand U6087 (N_6087,N_2681,N_4712);
or U6088 (N_6088,N_3624,N_4896);
xnor U6089 (N_6089,N_3949,N_4269);
or U6090 (N_6090,N_4480,N_3865);
or U6091 (N_6091,N_3566,N_3394);
or U6092 (N_6092,N_3006,N_3887);
and U6093 (N_6093,N_3467,N_4893);
or U6094 (N_6094,N_4506,N_4890);
nor U6095 (N_6095,N_4446,N_4295);
xnor U6096 (N_6096,N_3960,N_3918);
and U6097 (N_6097,N_2828,N_3063);
nand U6098 (N_6098,N_3380,N_2539);
xnor U6099 (N_6099,N_4566,N_2574);
xor U6100 (N_6100,N_2716,N_2903);
nor U6101 (N_6101,N_2627,N_4987);
nand U6102 (N_6102,N_4637,N_4052);
and U6103 (N_6103,N_2928,N_4386);
and U6104 (N_6104,N_4096,N_4356);
and U6105 (N_6105,N_2915,N_4399);
and U6106 (N_6106,N_4693,N_3295);
nand U6107 (N_6107,N_3541,N_4041);
or U6108 (N_6108,N_3198,N_4763);
or U6109 (N_6109,N_4380,N_4668);
nand U6110 (N_6110,N_3122,N_2514);
and U6111 (N_6111,N_3014,N_2907);
nor U6112 (N_6112,N_2840,N_3270);
xnor U6113 (N_6113,N_2957,N_2816);
nor U6114 (N_6114,N_3090,N_4746);
nor U6115 (N_6115,N_4769,N_4410);
nand U6116 (N_6116,N_4407,N_2688);
or U6117 (N_6117,N_2616,N_3248);
or U6118 (N_6118,N_4851,N_3513);
nand U6119 (N_6119,N_4767,N_3692);
and U6120 (N_6120,N_3948,N_3653);
nor U6121 (N_6121,N_4095,N_4635);
and U6122 (N_6122,N_3724,N_4649);
xnor U6123 (N_6123,N_3349,N_4132);
and U6124 (N_6124,N_4690,N_3172);
xnor U6125 (N_6125,N_4412,N_2935);
xnor U6126 (N_6126,N_4545,N_4400);
or U6127 (N_6127,N_2650,N_4648);
nor U6128 (N_6128,N_4917,N_4149);
xor U6129 (N_6129,N_4745,N_3967);
or U6130 (N_6130,N_4313,N_3392);
xnor U6131 (N_6131,N_4449,N_3311);
or U6132 (N_6132,N_4563,N_4495);
and U6133 (N_6133,N_4859,N_2978);
xor U6134 (N_6134,N_4823,N_3839);
xor U6135 (N_6135,N_4241,N_3103);
nand U6136 (N_6136,N_4274,N_2549);
or U6137 (N_6137,N_4377,N_2958);
or U6138 (N_6138,N_2952,N_4986);
xnor U6139 (N_6139,N_2575,N_3798);
nor U6140 (N_6140,N_4305,N_3042);
xnor U6141 (N_6141,N_3049,N_3454);
xnor U6142 (N_6142,N_3804,N_3909);
nor U6143 (N_6143,N_3222,N_2545);
xnor U6144 (N_6144,N_3471,N_4382);
and U6145 (N_6145,N_3788,N_3916);
and U6146 (N_6146,N_4023,N_2599);
xor U6147 (N_6147,N_3657,N_4838);
xor U6148 (N_6148,N_2503,N_3696);
xor U6149 (N_6149,N_3953,N_3094);
nor U6150 (N_6150,N_3258,N_2795);
nand U6151 (N_6151,N_4148,N_2762);
and U6152 (N_6152,N_4918,N_4288);
or U6153 (N_6153,N_4067,N_2893);
nor U6154 (N_6154,N_2631,N_4730);
xnor U6155 (N_6155,N_3853,N_4700);
or U6156 (N_6156,N_3823,N_4722);
nor U6157 (N_6157,N_4630,N_2620);
and U6158 (N_6158,N_4589,N_4439);
nand U6159 (N_6159,N_3717,N_2861);
and U6160 (N_6160,N_3626,N_4183);
nand U6161 (N_6161,N_2524,N_4772);
nor U6162 (N_6162,N_2675,N_4526);
nand U6163 (N_6163,N_3332,N_4154);
xor U6164 (N_6164,N_2799,N_4685);
xnor U6165 (N_6165,N_3854,N_2613);
or U6166 (N_6166,N_3325,N_3904);
and U6167 (N_6167,N_4667,N_3020);
nand U6168 (N_6168,N_4081,N_3131);
or U6169 (N_6169,N_2814,N_2862);
xnor U6170 (N_6170,N_2973,N_3400);
nand U6171 (N_6171,N_4482,N_3992);
nor U6172 (N_6172,N_2830,N_3064);
nand U6173 (N_6173,N_4499,N_2581);
nor U6174 (N_6174,N_3970,N_2568);
xnor U6175 (N_6175,N_2860,N_4664);
nand U6176 (N_6176,N_2750,N_4844);
nor U6177 (N_6177,N_4144,N_4170);
and U6178 (N_6178,N_3488,N_2926);
and U6179 (N_6179,N_4296,N_2615);
and U6180 (N_6180,N_2988,N_4481);
nor U6181 (N_6181,N_3510,N_3569);
nand U6182 (N_6182,N_3831,N_4974);
xor U6183 (N_6183,N_4556,N_3874);
or U6184 (N_6184,N_4620,N_2868);
nor U6185 (N_6185,N_3086,N_3611);
or U6186 (N_6186,N_3168,N_3923);
nor U6187 (N_6187,N_3880,N_3841);
and U6188 (N_6188,N_4066,N_3111);
or U6189 (N_6189,N_4282,N_4795);
xnor U6190 (N_6190,N_4008,N_2740);
and U6191 (N_6191,N_3758,N_3588);
xor U6192 (N_6192,N_3161,N_2680);
nand U6193 (N_6193,N_4141,N_2530);
nor U6194 (N_6194,N_3685,N_4525);
or U6195 (N_6195,N_3684,N_3407);
or U6196 (N_6196,N_2776,N_4945);
or U6197 (N_6197,N_2956,N_3391);
xnor U6198 (N_6198,N_4350,N_2677);
nor U6199 (N_6199,N_4383,N_3771);
nor U6200 (N_6200,N_4490,N_4249);
nor U6201 (N_6201,N_4536,N_4494);
nor U6202 (N_6202,N_4520,N_4967);
nand U6203 (N_6203,N_4857,N_2594);
nor U6204 (N_6204,N_2708,N_4071);
nand U6205 (N_6205,N_4094,N_3055);
nand U6206 (N_6206,N_4922,N_3093);
and U6207 (N_6207,N_3646,N_4835);
and U6208 (N_6208,N_3317,N_4903);
nand U6209 (N_6209,N_2948,N_4822);
or U6210 (N_6210,N_3815,N_3242);
or U6211 (N_6211,N_4527,N_2561);
xnor U6212 (N_6212,N_2782,N_2752);
and U6213 (N_6213,N_3307,N_4253);
xnor U6214 (N_6214,N_2789,N_4101);
nor U6215 (N_6215,N_3217,N_3246);
and U6216 (N_6216,N_2819,N_2660);
nand U6217 (N_6217,N_4151,N_4121);
or U6218 (N_6218,N_2621,N_4250);
nor U6219 (N_6219,N_3716,N_2824);
xor U6220 (N_6220,N_4459,N_3155);
or U6221 (N_6221,N_3213,N_4283);
xnor U6222 (N_6222,N_4111,N_2536);
nor U6223 (N_6223,N_3496,N_4699);
and U6224 (N_6224,N_4771,N_4320);
or U6225 (N_6225,N_4164,N_3508);
xnor U6226 (N_6226,N_3018,N_4626);
xor U6227 (N_6227,N_4551,N_4194);
nor U6228 (N_6228,N_3517,N_3101);
xnor U6229 (N_6229,N_4053,N_4592);
and U6230 (N_6230,N_3694,N_3395);
and U6231 (N_6231,N_2839,N_4765);
nand U6232 (N_6232,N_4185,N_2535);
nand U6233 (N_6233,N_3235,N_3715);
or U6234 (N_6234,N_4753,N_3362);
xnor U6235 (N_6235,N_3547,N_3651);
and U6236 (N_6236,N_2516,N_3415);
nor U6237 (N_6237,N_2917,N_4146);
nand U6238 (N_6238,N_4993,N_2573);
nor U6239 (N_6239,N_2590,N_4192);
xnor U6240 (N_6240,N_4409,N_3169);
nor U6241 (N_6241,N_3755,N_4959);
xnor U6242 (N_6242,N_2951,N_4135);
and U6243 (N_6243,N_4222,N_4511);
or U6244 (N_6244,N_2966,N_3339);
nor U6245 (N_6245,N_3748,N_4025);
and U6246 (N_6246,N_2571,N_3678);
nand U6247 (N_6247,N_2667,N_3373);
xnor U6248 (N_6248,N_3847,N_3497);
nand U6249 (N_6249,N_4910,N_3453);
xnor U6250 (N_6250,N_3974,N_3305);
and U6251 (N_6251,N_4637,N_4174);
nor U6252 (N_6252,N_2595,N_2827);
nand U6253 (N_6253,N_3035,N_4985);
and U6254 (N_6254,N_4133,N_4043);
nand U6255 (N_6255,N_3391,N_3922);
nor U6256 (N_6256,N_2506,N_4662);
nor U6257 (N_6257,N_4718,N_2840);
and U6258 (N_6258,N_4606,N_3847);
or U6259 (N_6259,N_4291,N_3067);
xor U6260 (N_6260,N_3285,N_3784);
nand U6261 (N_6261,N_4537,N_4669);
nor U6262 (N_6262,N_3880,N_3176);
or U6263 (N_6263,N_3953,N_3806);
xnor U6264 (N_6264,N_4998,N_3110);
xnor U6265 (N_6265,N_3662,N_3880);
or U6266 (N_6266,N_2829,N_4792);
xor U6267 (N_6267,N_2915,N_3804);
xnor U6268 (N_6268,N_3095,N_2805);
or U6269 (N_6269,N_3114,N_4365);
nor U6270 (N_6270,N_3635,N_3329);
nor U6271 (N_6271,N_3412,N_3773);
nor U6272 (N_6272,N_4767,N_3496);
or U6273 (N_6273,N_3790,N_3472);
and U6274 (N_6274,N_3752,N_3596);
and U6275 (N_6275,N_3785,N_4488);
and U6276 (N_6276,N_2831,N_4080);
and U6277 (N_6277,N_2705,N_3265);
nand U6278 (N_6278,N_3041,N_4767);
or U6279 (N_6279,N_3269,N_4264);
nor U6280 (N_6280,N_4039,N_4956);
nor U6281 (N_6281,N_4632,N_3711);
and U6282 (N_6282,N_4723,N_3443);
xor U6283 (N_6283,N_2696,N_3928);
nand U6284 (N_6284,N_3583,N_3184);
nor U6285 (N_6285,N_4648,N_3828);
nand U6286 (N_6286,N_4588,N_3000);
xor U6287 (N_6287,N_3804,N_3817);
nor U6288 (N_6288,N_4211,N_2970);
and U6289 (N_6289,N_3388,N_4455);
nand U6290 (N_6290,N_3779,N_4113);
xnor U6291 (N_6291,N_2580,N_2673);
nand U6292 (N_6292,N_3060,N_3217);
xnor U6293 (N_6293,N_2613,N_2848);
nand U6294 (N_6294,N_4716,N_3092);
xor U6295 (N_6295,N_3411,N_3260);
xor U6296 (N_6296,N_4947,N_4130);
or U6297 (N_6297,N_4092,N_4752);
nor U6298 (N_6298,N_4408,N_4469);
nand U6299 (N_6299,N_4373,N_4977);
xnor U6300 (N_6300,N_2895,N_4040);
or U6301 (N_6301,N_2531,N_2658);
nand U6302 (N_6302,N_3847,N_3265);
xor U6303 (N_6303,N_3097,N_3013);
nand U6304 (N_6304,N_3933,N_4669);
nand U6305 (N_6305,N_3524,N_3827);
and U6306 (N_6306,N_4308,N_4762);
xor U6307 (N_6307,N_4601,N_4627);
xor U6308 (N_6308,N_2968,N_3310);
xor U6309 (N_6309,N_4541,N_2730);
and U6310 (N_6310,N_4844,N_4753);
nor U6311 (N_6311,N_3182,N_3824);
nor U6312 (N_6312,N_3354,N_3248);
and U6313 (N_6313,N_2695,N_2879);
nand U6314 (N_6314,N_4583,N_4717);
and U6315 (N_6315,N_2523,N_3313);
or U6316 (N_6316,N_2671,N_4008);
nand U6317 (N_6317,N_2797,N_4303);
or U6318 (N_6318,N_4784,N_2849);
and U6319 (N_6319,N_3251,N_4215);
xnor U6320 (N_6320,N_4479,N_4802);
nor U6321 (N_6321,N_3853,N_3191);
nor U6322 (N_6322,N_3010,N_3585);
and U6323 (N_6323,N_4617,N_2822);
nor U6324 (N_6324,N_4426,N_3243);
or U6325 (N_6325,N_2955,N_3001);
xor U6326 (N_6326,N_4678,N_4137);
and U6327 (N_6327,N_3199,N_4113);
nand U6328 (N_6328,N_4502,N_3001);
and U6329 (N_6329,N_2699,N_3887);
and U6330 (N_6330,N_4482,N_3047);
nand U6331 (N_6331,N_3768,N_4291);
and U6332 (N_6332,N_2927,N_3671);
or U6333 (N_6333,N_3710,N_3927);
nor U6334 (N_6334,N_4384,N_3431);
nor U6335 (N_6335,N_4033,N_2927);
nor U6336 (N_6336,N_2587,N_3920);
or U6337 (N_6337,N_3765,N_2634);
and U6338 (N_6338,N_2662,N_2670);
nor U6339 (N_6339,N_2527,N_3186);
nor U6340 (N_6340,N_3845,N_4066);
and U6341 (N_6341,N_3308,N_4759);
xnor U6342 (N_6342,N_3913,N_3387);
or U6343 (N_6343,N_2718,N_4939);
nor U6344 (N_6344,N_4788,N_2865);
and U6345 (N_6345,N_2847,N_2854);
nand U6346 (N_6346,N_2762,N_2945);
and U6347 (N_6347,N_4752,N_2696);
xor U6348 (N_6348,N_4472,N_3997);
and U6349 (N_6349,N_2871,N_4428);
nor U6350 (N_6350,N_3531,N_4839);
and U6351 (N_6351,N_3282,N_4280);
and U6352 (N_6352,N_4207,N_4806);
or U6353 (N_6353,N_3983,N_4299);
nor U6354 (N_6354,N_3039,N_2924);
or U6355 (N_6355,N_3359,N_4085);
xnor U6356 (N_6356,N_2688,N_3649);
and U6357 (N_6357,N_4407,N_4877);
nor U6358 (N_6358,N_4428,N_2802);
nor U6359 (N_6359,N_4105,N_2832);
nand U6360 (N_6360,N_3629,N_3310);
or U6361 (N_6361,N_3182,N_3761);
and U6362 (N_6362,N_2752,N_2715);
xor U6363 (N_6363,N_4170,N_4326);
and U6364 (N_6364,N_4141,N_3879);
xnor U6365 (N_6365,N_4893,N_4998);
xnor U6366 (N_6366,N_3855,N_4647);
xor U6367 (N_6367,N_3662,N_4592);
or U6368 (N_6368,N_2707,N_2977);
xor U6369 (N_6369,N_2729,N_2720);
and U6370 (N_6370,N_2546,N_4209);
or U6371 (N_6371,N_3409,N_3673);
or U6372 (N_6372,N_4383,N_3692);
nor U6373 (N_6373,N_3233,N_3494);
nor U6374 (N_6374,N_3424,N_4337);
and U6375 (N_6375,N_2997,N_4283);
nor U6376 (N_6376,N_3534,N_4383);
or U6377 (N_6377,N_4051,N_3365);
or U6378 (N_6378,N_3956,N_3105);
nor U6379 (N_6379,N_3314,N_3067);
xor U6380 (N_6380,N_3630,N_3591);
or U6381 (N_6381,N_4879,N_3256);
nor U6382 (N_6382,N_3511,N_3984);
or U6383 (N_6383,N_4021,N_3537);
or U6384 (N_6384,N_4987,N_2740);
or U6385 (N_6385,N_4751,N_2639);
nand U6386 (N_6386,N_4567,N_4549);
and U6387 (N_6387,N_3502,N_4200);
nand U6388 (N_6388,N_3667,N_4193);
nor U6389 (N_6389,N_4604,N_3754);
nand U6390 (N_6390,N_2919,N_3110);
or U6391 (N_6391,N_2705,N_4188);
nand U6392 (N_6392,N_4079,N_3021);
xnor U6393 (N_6393,N_2577,N_4695);
nor U6394 (N_6394,N_4765,N_3360);
and U6395 (N_6395,N_3179,N_3257);
nand U6396 (N_6396,N_4733,N_3822);
xor U6397 (N_6397,N_3922,N_4088);
and U6398 (N_6398,N_4552,N_4613);
or U6399 (N_6399,N_4443,N_2657);
xnor U6400 (N_6400,N_3802,N_3963);
xnor U6401 (N_6401,N_3364,N_3173);
or U6402 (N_6402,N_4008,N_3271);
and U6403 (N_6403,N_2532,N_3000);
nor U6404 (N_6404,N_4097,N_4879);
nand U6405 (N_6405,N_4569,N_2925);
or U6406 (N_6406,N_3794,N_2985);
or U6407 (N_6407,N_4732,N_2546);
or U6408 (N_6408,N_4649,N_3288);
and U6409 (N_6409,N_4873,N_3403);
xnor U6410 (N_6410,N_2773,N_2702);
and U6411 (N_6411,N_4072,N_4572);
nand U6412 (N_6412,N_2518,N_4955);
xnor U6413 (N_6413,N_4860,N_2631);
nand U6414 (N_6414,N_4137,N_3856);
xor U6415 (N_6415,N_4354,N_3668);
xor U6416 (N_6416,N_2987,N_3534);
or U6417 (N_6417,N_4988,N_3217);
or U6418 (N_6418,N_4282,N_2564);
nand U6419 (N_6419,N_4805,N_3133);
and U6420 (N_6420,N_4976,N_3081);
nor U6421 (N_6421,N_4321,N_3370);
nand U6422 (N_6422,N_3523,N_4877);
or U6423 (N_6423,N_4288,N_3621);
nor U6424 (N_6424,N_4737,N_3375);
nor U6425 (N_6425,N_3334,N_3280);
nand U6426 (N_6426,N_4136,N_3891);
nand U6427 (N_6427,N_3127,N_4330);
nand U6428 (N_6428,N_4824,N_3785);
xor U6429 (N_6429,N_3759,N_3592);
nor U6430 (N_6430,N_4644,N_3877);
nor U6431 (N_6431,N_3373,N_4386);
nand U6432 (N_6432,N_3308,N_4078);
nor U6433 (N_6433,N_4697,N_4946);
nor U6434 (N_6434,N_2949,N_4537);
xor U6435 (N_6435,N_3062,N_4464);
nor U6436 (N_6436,N_4303,N_2934);
xor U6437 (N_6437,N_4579,N_3173);
and U6438 (N_6438,N_4514,N_3797);
nor U6439 (N_6439,N_4288,N_3195);
and U6440 (N_6440,N_3619,N_3522);
xnor U6441 (N_6441,N_2814,N_4275);
and U6442 (N_6442,N_2853,N_3222);
xor U6443 (N_6443,N_3998,N_2637);
and U6444 (N_6444,N_2950,N_4526);
nand U6445 (N_6445,N_4133,N_4890);
and U6446 (N_6446,N_2760,N_4238);
nand U6447 (N_6447,N_3915,N_2604);
xnor U6448 (N_6448,N_4924,N_2974);
nand U6449 (N_6449,N_2638,N_4380);
nand U6450 (N_6450,N_3402,N_4495);
xor U6451 (N_6451,N_3291,N_3528);
nand U6452 (N_6452,N_2964,N_4877);
and U6453 (N_6453,N_2883,N_3152);
xor U6454 (N_6454,N_3826,N_4153);
nor U6455 (N_6455,N_4027,N_3549);
or U6456 (N_6456,N_2720,N_4343);
or U6457 (N_6457,N_3430,N_4307);
nand U6458 (N_6458,N_2942,N_4387);
and U6459 (N_6459,N_3824,N_3960);
or U6460 (N_6460,N_2518,N_3933);
nor U6461 (N_6461,N_4764,N_4475);
nand U6462 (N_6462,N_2673,N_4972);
and U6463 (N_6463,N_2867,N_4615);
nor U6464 (N_6464,N_4601,N_4175);
xor U6465 (N_6465,N_2800,N_3975);
or U6466 (N_6466,N_3763,N_3950);
nor U6467 (N_6467,N_3227,N_3188);
nand U6468 (N_6468,N_3189,N_4020);
nor U6469 (N_6469,N_2641,N_3437);
xnor U6470 (N_6470,N_3731,N_3656);
nand U6471 (N_6471,N_4864,N_4148);
nand U6472 (N_6472,N_4657,N_2663);
nor U6473 (N_6473,N_4632,N_4922);
and U6474 (N_6474,N_2823,N_3740);
xor U6475 (N_6475,N_3994,N_2835);
nand U6476 (N_6476,N_4195,N_3390);
nor U6477 (N_6477,N_4629,N_4260);
nor U6478 (N_6478,N_3768,N_2624);
xor U6479 (N_6479,N_2894,N_4054);
nor U6480 (N_6480,N_4424,N_4195);
or U6481 (N_6481,N_3457,N_3810);
xor U6482 (N_6482,N_2983,N_3556);
and U6483 (N_6483,N_2805,N_4942);
and U6484 (N_6484,N_2866,N_3111);
or U6485 (N_6485,N_4212,N_3080);
and U6486 (N_6486,N_4732,N_3718);
and U6487 (N_6487,N_3513,N_3336);
and U6488 (N_6488,N_3778,N_4725);
and U6489 (N_6489,N_4971,N_3637);
and U6490 (N_6490,N_4117,N_4913);
and U6491 (N_6491,N_2809,N_3512);
and U6492 (N_6492,N_3823,N_4254);
and U6493 (N_6493,N_4554,N_4942);
nor U6494 (N_6494,N_3941,N_2769);
and U6495 (N_6495,N_2839,N_4218);
xor U6496 (N_6496,N_2812,N_4916);
and U6497 (N_6497,N_3313,N_4327);
nand U6498 (N_6498,N_3661,N_3617);
nand U6499 (N_6499,N_3579,N_3501);
xor U6500 (N_6500,N_3072,N_4497);
or U6501 (N_6501,N_4584,N_3600);
or U6502 (N_6502,N_3510,N_2689);
or U6503 (N_6503,N_2691,N_3720);
or U6504 (N_6504,N_3932,N_4945);
nand U6505 (N_6505,N_3219,N_4726);
or U6506 (N_6506,N_3354,N_3921);
nor U6507 (N_6507,N_4503,N_4354);
and U6508 (N_6508,N_2805,N_3467);
xnor U6509 (N_6509,N_4379,N_2658);
xnor U6510 (N_6510,N_4614,N_4817);
nand U6511 (N_6511,N_2684,N_4704);
and U6512 (N_6512,N_3828,N_3206);
or U6513 (N_6513,N_4066,N_4134);
nand U6514 (N_6514,N_3743,N_2983);
or U6515 (N_6515,N_3906,N_4411);
xnor U6516 (N_6516,N_3135,N_2819);
nor U6517 (N_6517,N_4176,N_4891);
or U6518 (N_6518,N_2972,N_3483);
xor U6519 (N_6519,N_4854,N_4918);
and U6520 (N_6520,N_4313,N_4903);
xor U6521 (N_6521,N_2806,N_3856);
and U6522 (N_6522,N_3743,N_3671);
and U6523 (N_6523,N_4171,N_2687);
nor U6524 (N_6524,N_2512,N_4505);
xnor U6525 (N_6525,N_4637,N_4240);
nand U6526 (N_6526,N_2684,N_4933);
or U6527 (N_6527,N_4653,N_4144);
and U6528 (N_6528,N_4891,N_3307);
and U6529 (N_6529,N_3957,N_2969);
xnor U6530 (N_6530,N_2513,N_4231);
xnor U6531 (N_6531,N_3145,N_4036);
nor U6532 (N_6532,N_4408,N_2796);
or U6533 (N_6533,N_2709,N_4113);
nor U6534 (N_6534,N_4011,N_4354);
and U6535 (N_6535,N_4200,N_4497);
xnor U6536 (N_6536,N_4141,N_2612);
or U6537 (N_6537,N_3227,N_4950);
xnor U6538 (N_6538,N_3377,N_2733);
nand U6539 (N_6539,N_4257,N_3798);
or U6540 (N_6540,N_3471,N_3952);
nand U6541 (N_6541,N_3985,N_3787);
nand U6542 (N_6542,N_3544,N_3276);
and U6543 (N_6543,N_4729,N_2681);
and U6544 (N_6544,N_4405,N_3502);
and U6545 (N_6545,N_4273,N_4284);
xor U6546 (N_6546,N_4592,N_3009);
or U6547 (N_6547,N_3101,N_2614);
or U6548 (N_6548,N_2680,N_2596);
or U6549 (N_6549,N_4745,N_3821);
xor U6550 (N_6550,N_3550,N_3191);
or U6551 (N_6551,N_4561,N_4810);
or U6552 (N_6552,N_3160,N_3081);
nor U6553 (N_6553,N_3572,N_3145);
or U6554 (N_6554,N_4987,N_3728);
or U6555 (N_6555,N_3765,N_4465);
nor U6556 (N_6556,N_2798,N_4224);
xor U6557 (N_6557,N_3844,N_4475);
nand U6558 (N_6558,N_3703,N_3559);
xnor U6559 (N_6559,N_3353,N_2601);
or U6560 (N_6560,N_4528,N_4886);
or U6561 (N_6561,N_3110,N_3835);
nor U6562 (N_6562,N_4206,N_4847);
xor U6563 (N_6563,N_4933,N_4268);
and U6564 (N_6564,N_4231,N_3528);
nor U6565 (N_6565,N_2836,N_4359);
xor U6566 (N_6566,N_4389,N_4787);
and U6567 (N_6567,N_3790,N_4001);
xnor U6568 (N_6568,N_2746,N_4678);
nor U6569 (N_6569,N_2583,N_3533);
nand U6570 (N_6570,N_3535,N_3432);
nor U6571 (N_6571,N_2841,N_4962);
or U6572 (N_6572,N_4043,N_3486);
or U6573 (N_6573,N_3220,N_2863);
and U6574 (N_6574,N_4171,N_3808);
nor U6575 (N_6575,N_2970,N_3323);
xnor U6576 (N_6576,N_4702,N_4796);
or U6577 (N_6577,N_4443,N_3386);
nor U6578 (N_6578,N_2809,N_3285);
or U6579 (N_6579,N_4362,N_3601);
or U6580 (N_6580,N_4605,N_3486);
and U6581 (N_6581,N_3829,N_3995);
xor U6582 (N_6582,N_4874,N_2774);
or U6583 (N_6583,N_4600,N_3479);
nor U6584 (N_6584,N_4753,N_4097);
or U6585 (N_6585,N_3775,N_2559);
or U6586 (N_6586,N_3100,N_2924);
xnor U6587 (N_6587,N_4574,N_4200);
and U6588 (N_6588,N_2906,N_2528);
and U6589 (N_6589,N_2521,N_3867);
nor U6590 (N_6590,N_3403,N_3184);
xor U6591 (N_6591,N_4886,N_3138);
or U6592 (N_6592,N_2869,N_2839);
or U6593 (N_6593,N_3662,N_2722);
and U6594 (N_6594,N_4523,N_4958);
xnor U6595 (N_6595,N_2800,N_3349);
or U6596 (N_6596,N_4695,N_2809);
or U6597 (N_6597,N_2673,N_3701);
nor U6598 (N_6598,N_2733,N_3614);
and U6599 (N_6599,N_4017,N_4867);
or U6600 (N_6600,N_3957,N_4764);
nor U6601 (N_6601,N_4651,N_4732);
nand U6602 (N_6602,N_4315,N_2810);
nand U6603 (N_6603,N_4281,N_4904);
and U6604 (N_6604,N_3611,N_2589);
nand U6605 (N_6605,N_3268,N_3586);
nor U6606 (N_6606,N_4086,N_2568);
or U6607 (N_6607,N_3632,N_2924);
xnor U6608 (N_6608,N_3910,N_4845);
or U6609 (N_6609,N_3894,N_3608);
xnor U6610 (N_6610,N_4740,N_3869);
xnor U6611 (N_6611,N_4611,N_4630);
or U6612 (N_6612,N_4740,N_4604);
nand U6613 (N_6613,N_3029,N_2537);
or U6614 (N_6614,N_4221,N_3343);
nor U6615 (N_6615,N_3046,N_2530);
xnor U6616 (N_6616,N_3577,N_4415);
nor U6617 (N_6617,N_2618,N_4027);
or U6618 (N_6618,N_3018,N_4436);
nor U6619 (N_6619,N_3637,N_4622);
and U6620 (N_6620,N_2821,N_3685);
or U6621 (N_6621,N_2680,N_3231);
or U6622 (N_6622,N_4077,N_4631);
nor U6623 (N_6623,N_3805,N_3748);
nor U6624 (N_6624,N_4420,N_2768);
or U6625 (N_6625,N_3181,N_4263);
xnor U6626 (N_6626,N_3546,N_3820);
and U6627 (N_6627,N_4864,N_3250);
nand U6628 (N_6628,N_4996,N_3895);
nand U6629 (N_6629,N_4494,N_4169);
nor U6630 (N_6630,N_3347,N_2718);
nand U6631 (N_6631,N_3090,N_2950);
or U6632 (N_6632,N_2706,N_2667);
xor U6633 (N_6633,N_4852,N_4491);
nor U6634 (N_6634,N_4710,N_4329);
xnor U6635 (N_6635,N_4134,N_3721);
or U6636 (N_6636,N_4203,N_2938);
and U6637 (N_6637,N_4533,N_3643);
and U6638 (N_6638,N_4853,N_4659);
and U6639 (N_6639,N_2893,N_2686);
nand U6640 (N_6640,N_4277,N_4816);
or U6641 (N_6641,N_4086,N_3117);
or U6642 (N_6642,N_4636,N_3692);
nand U6643 (N_6643,N_3101,N_3364);
nand U6644 (N_6644,N_4457,N_2684);
and U6645 (N_6645,N_3747,N_4847);
and U6646 (N_6646,N_3400,N_3989);
or U6647 (N_6647,N_4718,N_3670);
nor U6648 (N_6648,N_4387,N_4576);
xor U6649 (N_6649,N_3249,N_3178);
nor U6650 (N_6650,N_2605,N_3629);
and U6651 (N_6651,N_3775,N_4581);
and U6652 (N_6652,N_4613,N_3290);
and U6653 (N_6653,N_3345,N_3927);
or U6654 (N_6654,N_3749,N_3091);
nor U6655 (N_6655,N_2513,N_3119);
nor U6656 (N_6656,N_4468,N_4639);
or U6657 (N_6657,N_3232,N_3520);
xor U6658 (N_6658,N_4148,N_2937);
nand U6659 (N_6659,N_3818,N_3885);
or U6660 (N_6660,N_2701,N_3396);
nand U6661 (N_6661,N_4973,N_3396);
xnor U6662 (N_6662,N_4931,N_3796);
and U6663 (N_6663,N_3372,N_3300);
xnor U6664 (N_6664,N_4081,N_2726);
nor U6665 (N_6665,N_3695,N_3872);
or U6666 (N_6666,N_2744,N_4462);
xnor U6667 (N_6667,N_3820,N_4468);
or U6668 (N_6668,N_3784,N_3696);
nor U6669 (N_6669,N_3975,N_4820);
and U6670 (N_6670,N_2568,N_4818);
nand U6671 (N_6671,N_4420,N_4217);
nor U6672 (N_6672,N_4326,N_4258);
nand U6673 (N_6673,N_4974,N_4628);
and U6674 (N_6674,N_4657,N_3319);
nor U6675 (N_6675,N_3899,N_3526);
nor U6676 (N_6676,N_3773,N_4450);
and U6677 (N_6677,N_4408,N_2848);
nand U6678 (N_6678,N_3666,N_4660);
and U6679 (N_6679,N_4898,N_2867);
nor U6680 (N_6680,N_4425,N_4673);
and U6681 (N_6681,N_2801,N_4437);
or U6682 (N_6682,N_4503,N_4461);
nor U6683 (N_6683,N_4920,N_3400);
nor U6684 (N_6684,N_4414,N_3065);
nand U6685 (N_6685,N_4309,N_4256);
nor U6686 (N_6686,N_2507,N_3456);
or U6687 (N_6687,N_2801,N_4075);
and U6688 (N_6688,N_2923,N_4202);
nand U6689 (N_6689,N_3138,N_2791);
xnor U6690 (N_6690,N_4617,N_2835);
or U6691 (N_6691,N_4405,N_3027);
or U6692 (N_6692,N_4335,N_3153);
or U6693 (N_6693,N_3139,N_3707);
xnor U6694 (N_6694,N_4474,N_4039);
and U6695 (N_6695,N_4111,N_2686);
nor U6696 (N_6696,N_2831,N_3458);
nor U6697 (N_6697,N_4758,N_4445);
nand U6698 (N_6698,N_2999,N_2871);
xor U6699 (N_6699,N_2612,N_2931);
or U6700 (N_6700,N_4203,N_2921);
and U6701 (N_6701,N_3993,N_3737);
or U6702 (N_6702,N_2658,N_4292);
xnor U6703 (N_6703,N_3757,N_4600);
and U6704 (N_6704,N_3099,N_4375);
xor U6705 (N_6705,N_3992,N_4049);
nand U6706 (N_6706,N_2643,N_3293);
and U6707 (N_6707,N_3217,N_4707);
nand U6708 (N_6708,N_3399,N_4205);
xnor U6709 (N_6709,N_3479,N_4258);
or U6710 (N_6710,N_3792,N_4278);
or U6711 (N_6711,N_3409,N_3244);
nand U6712 (N_6712,N_2722,N_4336);
and U6713 (N_6713,N_4350,N_4020);
and U6714 (N_6714,N_4634,N_3610);
or U6715 (N_6715,N_3170,N_2729);
xor U6716 (N_6716,N_3824,N_4043);
nor U6717 (N_6717,N_3083,N_3161);
xnor U6718 (N_6718,N_3503,N_3833);
xor U6719 (N_6719,N_3599,N_4909);
or U6720 (N_6720,N_3496,N_2602);
and U6721 (N_6721,N_4770,N_2923);
nand U6722 (N_6722,N_2954,N_3452);
and U6723 (N_6723,N_2849,N_3768);
nor U6724 (N_6724,N_2872,N_4688);
and U6725 (N_6725,N_3911,N_3278);
nor U6726 (N_6726,N_3839,N_4308);
or U6727 (N_6727,N_3592,N_4572);
or U6728 (N_6728,N_3366,N_2986);
xnor U6729 (N_6729,N_4295,N_3586);
nand U6730 (N_6730,N_2639,N_4792);
nand U6731 (N_6731,N_2788,N_4768);
nand U6732 (N_6732,N_3717,N_3418);
nand U6733 (N_6733,N_3662,N_3678);
and U6734 (N_6734,N_4426,N_4901);
xor U6735 (N_6735,N_4955,N_4362);
and U6736 (N_6736,N_3597,N_4310);
nand U6737 (N_6737,N_3422,N_4899);
nor U6738 (N_6738,N_3446,N_4755);
or U6739 (N_6739,N_3721,N_4587);
nor U6740 (N_6740,N_2670,N_3101);
nand U6741 (N_6741,N_4206,N_3224);
xor U6742 (N_6742,N_3997,N_3567);
nor U6743 (N_6743,N_4309,N_2538);
xor U6744 (N_6744,N_3050,N_3472);
or U6745 (N_6745,N_2773,N_4699);
or U6746 (N_6746,N_4116,N_4864);
xnor U6747 (N_6747,N_2614,N_4719);
nand U6748 (N_6748,N_2932,N_3925);
xnor U6749 (N_6749,N_2947,N_4915);
nor U6750 (N_6750,N_4251,N_4039);
or U6751 (N_6751,N_3419,N_2783);
nor U6752 (N_6752,N_3141,N_4368);
nor U6753 (N_6753,N_2973,N_3515);
nor U6754 (N_6754,N_3942,N_3769);
and U6755 (N_6755,N_2932,N_4761);
or U6756 (N_6756,N_3502,N_2769);
xnor U6757 (N_6757,N_4754,N_3511);
nand U6758 (N_6758,N_3609,N_4060);
nor U6759 (N_6759,N_3126,N_3461);
and U6760 (N_6760,N_4947,N_4725);
and U6761 (N_6761,N_3756,N_4564);
or U6762 (N_6762,N_4543,N_3457);
xnor U6763 (N_6763,N_4656,N_4688);
nor U6764 (N_6764,N_3623,N_4961);
xor U6765 (N_6765,N_4944,N_2872);
or U6766 (N_6766,N_2607,N_4309);
and U6767 (N_6767,N_3103,N_2552);
nand U6768 (N_6768,N_4997,N_4124);
or U6769 (N_6769,N_4224,N_3681);
nand U6770 (N_6770,N_3126,N_3540);
and U6771 (N_6771,N_4861,N_4102);
xor U6772 (N_6772,N_3898,N_3762);
xnor U6773 (N_6773,N_3023,N_3188);
nand U6774 (N_6774,N_4831,N_4927);
and U6775 (N_6775,N_3271,N_3822);
nor U6776 (N_6776,N_4535,N_4845);
xnor U6777 (N_6777,N_4562,N_2513);
or U6778 (N_6778,N_3436,N_2602);
nand U6779 (N_6779,N_3355,N_4882);
nand U6780 (N_6780,N_3490,N_3068);
nand U6781 (N_6781,N_3829,N_2666);
and U6782 (N_6782,N_4025,N_4891);
and U6783 (N_6783,N_3155,N_4222);
xor U6784 (N_6784,N_3435,N_2538);
nand U6785 (N_6785,N_4113,N_3635);
xor U6786 (N_6786,N_3032,N_2883);
or U6787 (N_6787,N_4580,N_3892);
nor U6788 (N_6788,N_2953,N_3073);
nand U6789 (N_6789,N_4700,N_4496);
or U6790 (N_6790,N_3336,N_3616);
xnor U6791 (N_6791,N_3753,N_3391);
and U6792 (N_6792,N_2634,N_2719);
and U6793 (N_6793,N_2905,N_4607);
and U6794 (N_6794,N_4520,N_4323);
xnor U6795 (N_6795,N_4069,N_4981);
nand U6796 (N_6796,N_2949,N_4111);
nand U6797 (N_6797,N_4036,N_3616);
nor U6798 (N_6798,N_3858,N_3603);
or U6799 (N_6799,N_2874,N_3359);
nand U6800 (N_6800,N_4191,N_2542);
nor U6801 (N_6801,N_3356,N_3872);
or U6802 (N_6802,N_2969,N_4358);
or U6803 (N_6803,N_4769,N_2822);
nand U6804 (N_6804,N_4228,N_4196);
or U6805 (N_6805,N_4203,N_2596);
or U6806 (N_6806,N_3506,N_4071);
and U6807 (N_6807,N_3619,N_4921);
nand U6808 (N_6808,N_4794,N_3533);
or U6809 (N_6809,N_4161,N_4314);
and U6810 (N_6810,N_2819,N_3874);
nand U6811 (N_6811,N_4587,N_3273);
nand U6812 (N_6812,N_4587,N_4874);
or U6813 (N_6813,N_4395,N_4731);
and U6814 (N_6814,N_3844,N_3129);
nand U6815 (N_6815,N_4857,N_4994);
and U6816 (N_6816,N_3955,N_3566);
nand U6817 (N_6817,N_2714,N_4842);
nor U6818 (N_6818,N_3973,N_3481);
or U6819 (N_6819,N_2684,N_3328);
xnor U6820 (N_6820,N_3754,N_3272);
xnor U6821 (N_6821,N_2700,N_3383);
xor U6822 (N_6822,N_4762,N_3898);
nor U6823 (N_6823,N_4589,N_3965);
xor U6824 (N_6824,N_4644,N_2770);
and U6825 (N_6825,N_3435,N_4342);
xor U6826 (N_6826,N_4407,N_4220);
xor U6827 (N_6827,N_3482,N_4275);
xor U6828 (N_6828,N_4072,N_4399);
nor U6829 (N_6829,N_2762,N_4426);
or U6830 (N_6830,N_3815,N_3023);
and U6831 (N_6831,N_3320,N_3422);
nand U6832 (N_6832,N_3528,N_4243);
xor U6833 (N_6833,N_3859,N_4904);
nand U6834 (N_6834,N_3778,N_3457);
or U6835 (N_6835,N_3004,N_4441);
xnor U6836 (N_6836,N_3550,N_4466);
or U6837 (N_6837,N_3633,N_2745);
nor U6838 (N_6838,N_4838,N_4110);
nor U6839 (N_6839,N_3269,N_3619);
and U6840 (N_6840,N_3970,N_3187);
nand U6841 (N_6841,N_4409,N_3868);
nor U6842 (N_6842,N_3433,N_4739);
nor U6843 (N_6843,N_2846,N_4102);
or U6844 (N_6844,N_2569,N_2513);
and U6845 (N_6845,N_2575,N_4872);
xnor U6846 (N_6846,N_4970,N_3745);
nand U6847 (N_6847,N_2766,N_3112);
nand U6848 (N_6848,N_3536,N_3973);
xnor U6849 (N_6849,N_2572,N_4498);
nand U6850 (N_6850,N_3558,N_3566);
nor U6851 (N_6851,N_3095,N_3215);
or U6852 (N_6852,N_4063,N_4951);
xor U6853 (N_6853,N_2579,N_4438);
nand U6854 (N_6854,N_4701,N_4748);
nand U6855 (N_6855,N_4144,N_3151);
and U6856 (N_6856,N_3282,N_2682);
xnor U6857 (N_6857,N_3084,N_4189);
or U6858 (N_6858,N_3914,N_4776);
or U6859 (N_6859,N_4951,N_4862);
xnor U6860 (N_6860,N_3908,N_3659);
xor U6861 (N_6861,N_4677,N_3429);
and U6862 (N_6862,N_4357,N_3952);
or U6863 (N_6863,N_3691,N_3710);
nor U6864 (N_6864,N_2504,N_2803);
xnor U6865 (N_6865,N_3451,N_3629);
or U6866 (N_6866,N_2711,N_4041);
or U6867 (N_6867,N_3983,N_3646);
xor U6868 (N_6868,N_4066,N_4760);
nor U6869 (N_6869,N_2618,N_4038);
xnor U6870 (N_6870,N_4258,N_3446);
xor U6871 (N_6871,N_4049,N_2649);
or U6872 (N_6872,N_4575,N_3062);
and U6873 (N_6873,N_3586,N_4872);
and U6874 (N_6874,N_2686,N_3279);
or U6875 (N_6875,N_3217,N_4360);
nor U6876 (N_6876,N_3509,N_4144);
or U6877 (N_6877,N_2880,N_2741);
nand U6878 (N_6878,N_4988,N_3907);
and U6879 (N_6879,N_3731,N_3800);
nor U6880 (N_6880,N_3139,N_3204);
or U6881 (N_6881,N_4537,N_4563);
or U6882 (N_6882,N_4300,N_2663);
nand U6883 (N_6883,N_4457,N_4577);
xor U6884 (N_6884,N_4260,N_2620);
xnor U6885 (N_6885,N_4675,N_3013);
nand U6886 (N_6886,N_3137,N_4974);
xor U6887 (N_6887,N_3139,N_4525);
nand U6888 (N_6888,N_3212,N_4209);
nor U6889 (N_6889,N_2876,N_4677);
nand U6890 (N_6890,N_3800,N_4755);
or U6891 (N_6891,N_3938,N_3872);
nor U6892 (N_6892,N_4013,N_4110);
and U6893 (N_6893,N_4052,N_4671);
xor U6894 (N_6894,N_3648,N_3204);
nor U6895 (N_6895,N_3482,N_4857);
xor U6896 (N_6896,N_4952,N_4055);
or U6897 (N_6897,N_3182,N_4586);
nand U6898 (N_6898,N_4366,N_3029);
xor U6899 (N_6899,N_3935,N_4386);
and U6900 (N_6900,N_3893,N_3227);
nor U6901 (N_6901,N_4000,N_4399);
or U6902 (N_6902,N_2923,N_4233);
or U6903 (N_6903,N_3461,N_3683);
nor U6904 (N_6904,N_2722,N_2976);
xnor U6905 (N_6905,N_3664,N_4890);
nor U6906 (N_6906,N_3750,N_2873);
nand U6907 (N_6907,N_3850,N_2784);
or U6908 (N_6908,N_3365,N_4473);
nand U6909 (N_6909,N_3274,N_2693);
xor U6910 (N_6910,N_2697,N_2501);
xnor U6911 (N_6911,N_2708,N_4577);
or U6912 (N_6912,N_3719,N_3607);
xnor U6913 (N_6913,N_4575,N_3421);
or U6914 (N_6914,N_2661,N_4619);
and U6915 (N_6915,N_3926,N_4616);
and U6916 (N_6916,N_3813,N_3997);
or U6917 (N_6917,N_4720,N_3186);
xor U6918 (N_6918,N_3338,N_4392);
or U6919 (N_6919,N_3028,N_4588);
xnor U6920 (N_6920,N_3332,N_4500);
or U6921 (N_6921,N_2935,N_4657);
xor U6922 (N_6922,N_3412,N_3165);
and U6923 (N_6923,N_3912,N_2810);
nand U6924 (N_6924,N_4045,N_4811);
xor U6925 (N_6925,N_3693,N_4298);
nor U6926 (N_6926,N_2737,N_2687);
nor U6927 (N_6927,N_2507,N_3651);
nand U6928 (N_6928,N_4179,N_2936);
xnor U6929 (N_6929,N_2998,N_3281);
or U6930 (N_6930,N_2599,N_3989);
nand U6931 (N_6931,N_4899,N_4176);
nand U6932 (N_6932,N_3436,N_4312);
and U6933 (N_6933,N_2859,N_3147);
nand U6934 (N_6934,N_3092,N_3418);
and U6935 (N_6935,N_3860,N_4367);
nor U6936 (N_6936,N_3963,N_4652);
xnor U6937 (N_6937,N_4350,N_3084);
and U6938 (N_6938,N_2506,N_4050);
nor U6939 (N_6939,N_3094,N_3148);
nor U6940 (N_6940,N_4775,N_4912);
and U6941 (N_6941,N_4136,N_2607);
and U6942 (N_6942,N_2720,N_2651);
nor U6943 (N_6943,N_4191,N_4604);
nand U6944 (N_6944,N_3670,N_3068);
nand U6945 (N_6945,N_4326,N_4793);
and U6946 (N_6946,N_3327,N_2769);
and U6947 (N_6947,N_3813,N_3856);
and U6948 (N_6948,N_4227,N_2793);
and U6949 (N_6949,N_3134,N_2908);
nand U6950 (N_6950,N_4319,N_2624);
xnor U6951 (N_6951,N_2985,N_4391);
nand U6952 (N_6952,N_3810,N_2656);
and U6953 (N_6953,N_2885,N_4299);
xor U6954 (N_6954,N_3352,N_4883);
xnor U6955 (N_6955,N_4210,N_4691);
nand U6956 (N_6956,N_3141,N_3081);
and U6957 (N_6957,N_3307,N_4568);
or U6958 (N_6958,N_2972,N_4257);
nor U6959 (N_6959,N_3489,N_4332);
xor U6960 (N_6960,N_4962,N_4907);
nor U6961 (N_6961,N_2907,N_4975);
xor U6962 (N_6962,N_4535,N_4039);
nand U6963 (N_6963,N_3872,N_4055);
or U6964 (N_6964,N_3343,N_3483);
nor U6965 (N_6965,N_3742,N_3728);
nor U6966 (N_6966,N_2834,N_3606);
or U6967 (N_6967,N_3302,N_3419);
nand U6968 (N_6968,N_3878,N_4503);
nand U6969 (N_6969,N_4079,N_3156);
and U6970 (N_6970,N_2634,N_4778);
nand U6971 (N_6971,N_4546,N_4324);
or U6972 (N_6972,N_3585,N_2898);
or U6973 (N_6973,N_2670,N_3710);
xnor U6974 (N_6974,N_2991,N_2544);
and U6975 (N_6975,N_4928,N_3733);
or U6976 (N_6976,N_4431,N_2916);
nor U6977 (N_6977,N_3822,N_4187);
or U6978 (N_6978,N_4951,N_4999);
or U6979 (N_6979,N_3415,N_4886);
nor U6980 (N_6980,N_3510,N_3477);
xnor U6981 (N_6981,N_2926,N_3813);
and U6982 (N_6982,N_4624,N_4411);
nand U6983 (N_6983,N_2885,N_3741);
or U6984 (N_6984,N_3058,N_4037);
xor U6985 (N_6985,N_3829,N_2655);
xor U6986 (N_6986,N_4705,N_3976);
nor U6987 (N_6987,N_2647,N_3916);
xnor U6988 (N_6988,N_4850,N_3563);
xnor U6989 (N_6989,N_2527,N_4597);
and U6990 (N_6990,N_3869,N_3612);
and U6991 (N_6991,N_4815,N_3787);
or U6992 (N_6992,N_2868,N_2623);
nand U6993 (N_6993,N_3572,N_4739);
nor U6994 (N_6994,N_2829,N_3389);
xnor U6995 (N_6995,N_2821,N_3938);
or U6996 (N_6996,N_3800,N_3758);
nor U6997 (N_6997,N_4536,N_3010);
xor U6998 (N_6998,N_4326,N_3996);
nor U6999 (N_6999,N_4711,N_3323);
nand U7000 (N_7000,N_3927,N_3637);
nand U7001 (N_7001,N_3621,N_3279);
and U7002 (N_7002,N_3083,N_3541);
xor U7003 (N_7003,N_3174,N_3496);
and U7004 (N_7004,N_2763,N_3666);
and U7005 (N_7005,N_2657,N_3004);
and U7006 (N_7006,N_4190,N_3075);
xnor U7007 (N_7007,N_3167,N_3011);
xor U7008 (N_7008,N_4403,N_2835);
nor U7009 (N_7009,N_4000,N_4897);
or U7010 (N_7010,N_3259,N_3195);
nor U7011 (N_7011,N_4918,N_4732);
nor U7012 (N_7012,N_2603,N_2800);
and U7013 (N_7013,N_3219,N_3600);
and U7014 (N_7014,N_2579,N_4244);
or U7015 (N_7015,N_2822,N_3667);
nand U7016 (N_7016,N_3756,N_4775);
nand U7017 (N_7017,N_3888,N_3565);
nor U7018 (N_7018,N_3466,N_4797);
nor U7019 (N_7019,N_3487,N_4539);
nand U7020 (N_7020,N_3837,N_3609);
or U7021 (N_7021,N_2501,N_2649);
nor U7022 (N_7022,N_3503,N_4275);
and U7023 (N_7023,N_3928,N_4911);
or U7024 (N_7024,N_3777,N_3026);
and U7025 (N_7025,N_3887,N_3397);
and U7026 (N_7026,N_2634,N_2982);
nand U7027 (N_7027,N_4872,N_4285);
nor U7028 (N_7028,N_4136,N_3576);
nand U7029 (N_7029,N_3136,N_4781);
nand U7030 (N_7030,N_3243,N_3462);
or U7031 (N_7031,N_3802,N_4723);
xnor U7032 (N_7032,N_4503,N_3638);
nand U7033 (N_7033,N_3511,N_3319);
xnor U7034 (N_7034,N_3457,N_2775);
xnor U7035 (N_7035,N_4781,N_4986);
nand U7036 (N_7036,N_3628,N_4158);
nor U7037 (N_7037,N_2613,N_2836);
nor U7038 (N_7038,N_2806,N_4799);
nor U7039 (N_7039,N_3352,N_2688);
nand U7040 (N_7040,N_3562,N_2590);
xnor U7041 (N_7041,N_3775,N_4730);
nor U7042 (N_7042,N_4653,N_3064);
xnor U7043 (N_7043,N_4394,N_3076);
and U7044 (N_7044,N_3723,N_2659);
nand U7045 (N_7045,N_4848,N_3516);
nand U7046 (N_7046,N_2976,N_3360);
or U7047 (N_7047,N_3268,N_3476);
or U7048 (N_7048,N_3885,N_2689);
nand U7049 (N_7049,N_3247,N_4808);
and U7050 (N_7050,N_4808,N_3025);
nand U7051 (N_7051,N_3653,N_2533);
nor U7052 (N_7052,N_4309,N_2545);
xnor U7053 (N_7053,N_2696,N_4396);
xor U7054 (N_7054,N_4155,N_4507);
nor U7055 (N_7055,N_4655,N_4048);
xnor U7056 (N_7056,N_4766,N_2625);
or U7057 (N_7057,N_3574,N_4828);
nor U7058 (N_7058,N_3875,N_3768);
or U7059 (N_7059,N_3564,N_4576);
and U7060 (N_7060,N_3500,N_4973);
or U7061 (N_7061,N_3295,N_3424);
or U7062 (N_7062,N_3896,N_4823);
xor U7063 (N_7063,N_2845,N_3621);
nand U7064 (N_7064,N_3372,N_2978);
nor U7065 (N_7065,N_2797,N_3440);
or U7066 (N_7066,N_2748,N_4230);
nor U7067 (N_7067,N_4944,N_2770);
xor U7068 (N_7068,N_4567,N_4600);
or U7069 (N_7069,N_4023,N_4944);
and U7070 (N_7070,N_3259,N_3724);
and U7071 (N_7071,N_4048,N_4016);
nand U7072 (N_7072,N_4318,N_3072);
nand U7073 (N_7073,N_4301,N_3445);
xnor U7074 (N_7074,N_4903,N_3195);
xnor U7075 (N_7075,N_4403,N_3174);
nor U7076 (N_7076,N_4311,N_3336);
nor U7077 (N_7077,N_3328,N_2735);
xor U7078 (N_7078,N_4480,N_4111);
and U7079 (N_7079,N_4090,N_2615);
and U7080 (N_7080,N_4973,N_3688);
and U7081 (N_7081,N_3163,N_2604);
nor U7082 (N_7082,N_4874,N_4325);
nand U7083 (N_7083,N_3592,N_3681);
nor U7084 (N_7084,N_4818,N_3175);
nand U7085 (N_7085,N_4710,N_4114);
nand U7086 (N_7086,N_2577,N_2986);
nor U7087 (N_7087,N_4719,N_3440);
nor U7088 (N_7088,N_4027,N_4913);
xnor U7089 (N_7089,N_4590,N_2538);
or U7090 (N_7090,N_4480,N_2739);
nor U7091 (N_7091,N_4671,N_3868);
and U7092 (N_7092,N_4990,N_4775);
xnor U7093 (N_7093,N_2698,N_2708);
nor U7094 (N_7094,N_3133,N_3777);
nand U7095 (N_7095,N_2931,N_4724);
nor U7096 (N_7096,N_4120,N_3988);
and U7097 (N_7097,N_3589,N_4655);
or U7098 (N_7098,N_2630,N_2899);
xnor U7099 (N_7099,N_4008,N_2670);
xnor U7100 (N_7100,N_2652,N_4763);
xor U7101 (N_7101,N_2678,N_2590);
nand U7102 (N_7102,N_3566,N_3894);
nand U7103 (N_7103,N_4791,N_2937);
nor U7104 (N_7104,N_4817,N_3703);
and U7105 (N_7105,N_4909,N_4154);
xor U7106 (N_7106,N_2706,N_4664);
and U7107 (N_7107,N_3622,N_4839);
nor U7108 (N_7108,N_4344,N_2635);
nor U7109 (N_7109,N_3746,N_2696);
xnor U7110 (N_7110,N_4324,N_4164);
nor U7111 (N_7111,N_2859,N_4879);
and U7112 (N_7112,N_2747,N_4843);
nor U7113 (N_7113,N_4748,N_2692);
nand U7114 (N_7114,N_4275,N_2878);
or U7115 (N_7115,N_3855,N_4874);
and U7116 (N_7116,N_4573,N_2838);
xnor U7117 (N_7117,N_4735,N_4412);
xor U7118 (N_7118,N_3252,N_4050);
xnor U7119 (N_7119,N_4710,N_4918);
nand U7120 (N_7120,N_4792,N_4012);
and U7121 (N_7121,N_3652,N_3095);
xnor U7122 (N_7122,N_2881,N_4971);
and U7123 (N_7123,N_3829,N_4903);
or U7124 (N_7124,N_3116,N_3014);
and U7125 (N_7125,N_4921,N_4179);
or U7126 (N_7126,N_3651,N_3599);
nand U7127 (N_7127,N_4916,N_4361);
nand U7128 (N_7128,N_3947,N_3811);
xnor U7129 (N_7129,N_4421,N_3888);
or U7130 (N_7130,N_3107,N_2642);
nand U7131 (N_7131,N_4511,N_3281);
nand U7132 (N_7132,N_3786,N_3220);
or U7133 (N_7133,N_3836,N_2750);
nor U7134 (N_7134,N_4962,N_3110);
and U7135 (N_7135,N_4822,N_2655);
nand U7136 (N_7136,N_3219,N_3997);
nand U7137 (N_7137,N_2609,N_4246);
nor U7138 (N_7138,N_3228,N_2818);
nand U7139 (N_7139,N_3192,N_4596);
xnor U7140 (N_7140,N_3671,N_4724);
nand U7141 (N_7141,N_4040,N_2847);
or U7142 (N_7142,N_4966,N_2926);
and U7143 (N_7143,N_2639,N_3640);
nand U7144 (N_7144,N_3243,N_3094);
and U7145 (N_7145,N_3436,N_4138);
xor U7146 (N_7146,N_3187,N_3384);
nor U7147 (N_7147,N_3570,N_3320);
nor U7148 (N_7148,N_4609,N_4156);
nand U7149 (N_7149,N_4700,N_2627);
nand U7150 (N_7150,N_2942,N_4939);
xnor U7151 (N_7151,N_3122,N_3959);
nor U7152 (N_7152,N_4749,N_4482);
or U7153 (N_7153,N_3983,N_4999);
xnor U7154 (N_7154,N_3789,N_4895);
nor U7155 (N_7155,N_3730,N_2842);
nand U7156 (N_7156,N_3879,N_3049);
nand U7157 (N_7157,N_2544,N_3519);
nor U7158 (N_7158,N_3998,N_3798);
nand U7159 (N_7159,N_4889,N_3482);
xnor U7160 (N_7160,N_4726,N_3304);
and U7161 (N_7161,N_3419,N_3400);
xnor U7162 (N_7162,N_2956,N_4346);
nor U7163 (N_7163,N_2899,N_4612);
nor U7164 (N_7164,N_4447,N_4871);
xor U7165 (N_7165,N_2843,N_3582);
nor U7166 (N_7166,N_3397,N_4120);
and U7167 (N_7167,N_3742,N_4591);
nor U7168 (N_7168,N_2682,N_3901);
nor U7169 (N_7169,N_3807,N_3490);
xnor U7170 (N_7170,N_3283,N_2833);
xor U7171 (N_7171,N_4941,N_3707);
nand U7172 (N_7172,N_3656,N_2598);
xnor U7173 (N_7173,N_3194,N_4041);
nor U7174 (N_7174,N_2542,N_4722);
nor U7175 (N_7175,N_3648,N_4924);
and U7176 (N_7176,N_3274,N_2679);
or U7177 (N_7177,N_3883,N_3529);
and U7178 (N_7178,N_3934,N_3009);
xnor U7179 (N_7179,N_3408,N_3274);
or U7180 (N_7180,N_3287,N_4418);
xnor U7181 (N_7181,N_3160,N_3604);
xnor U7182 (N_7182,N_2971,N_2694);
and U7183 (N_7183,N_4197,N_4749);
xnor U7184 (N_7184,N_3648,N_3718);
xor U7185 (N_7185,N_4677,N_4861);
nand U7186 (N_7186,N_3757,N_4113);
and U7187 (N_7187,N_2553,N_4081);
nor U7188 (N_7188,N_3521,N_4355);
or U7189 (N_7189,N_3583,N_4536);
xnor U7190 (N_7190,N_3806,N_3159);
nor U7191 (N_7191,N_2822,N_4624);
or U7192 (N_7192,N_2895,N_3962);
nor U7193 (N_7193,N_3231,N_4434);
xnor U7194 (N_7194,N_3643,N_4677);
nor U7195 (N_7195,N_4785,N_3695);
and U7196 (N_7196,N_3323,N_2901);
xor U7197 (N_7197,N_4872,N_4679);
nand U7198 (N_7198,N_2579,N_3424);
nor U7199 (N_7199,N_3719,N_4954);
and U7200 (N_7200,N_4952,N_2643);
and U7201 (N_7201,N_3030,N_4228);
and U7202 (N_7202,N_4656,N_4337);
and U7203 (N_7203,N_4196,N_3031);
and U7204 (N_7204,N_2799,N_2809);
xor U7205 (N_7205,N_3115,N_4822);
and U7206 (N_7206,N_4846,N_3091);
xnor U7207 (N_7207,N_2654,N_4707);
xnor U7208 (N_7208,N_3236,N_3074);
or U7209 (N_7209,N_4868,N_4527);
nand U7210 (N_7210,N_3835,N_4252);
nor U7211 (N_7211,N_3867,N_2769);
nor U7212 (N_7212,N_3251,N_4090);
and U7213 (N_7213,N_3618,N_4408);
or U7214 (N_7214,N_4791,N_2905);
and U7215 (N_7215,N_3930,N_3387);
or U7216 (N_7216,N_3564,N_4201);
nand U7217 (N_7217,N_4492,N_3766);
xor U7218 (N_7218,N_3362,N_2941);
nor U7219 (N_7219,N_3185,N_4887);
or U7220 (N_7220,N_3081,N_4216);
nor U7221 (N_7221,N_4100,N_2860);
and U7222 (N_7222,N_4970,N_4436);
or U7223 (N_7223,N_3263,N_4292);
or U7224 (N_7224,N_4074,N_4806);
or U7225 (N_7225,N_4602,N_4124);
or U7226 (N_7226,N_2982,N_3051);
nor U7227 (N_7227,N_2755,N_4420);
nand U7228 (N_7228,N_4697,N_4072);
xor U7229 (N_7229,N_2510,N_4564);
and U7230 (N_7230,N_3916,N_3963);
nand U7231 (N_7231,N_4476,N_3324);
or U7232 (N_7232,N_3249,N_3537);
xor U7233 (N_7233,N_3923,N_4339);
and U7234 (N_7234,N_3100,N_3324);
and U7235 (N_7235,N_3176,N_4241);
or U7236 (N_7236,N_2629,N_4750);
nor U7237 (N_7237,N_4310,N_4876);
nand U7238 (N_7238,N_3921,N_2860);
xor U7239 (N_7239,N_3419,N_3681);
xnor U7240 (N_7240,N_3292,N_2821);
and U7241 (N_7241,N_4988,N_2623);
nand U7242 (N_7242,N_2516,N_3938);
or U7243 (N_7243,N_4308,N_4627);
xor U7244 (N_7244,N_3066,N_3832);
xor U7245 (N_7245,N_3589,N_4922);
nor U7246 (N_7246,N_4398,N_4632);
nor U7247 (N_7247,N_4669,N_4138);
nand U7248 (N_7248,N_3680,N_4299);
nor U7249 (N_7249,N_3048,N_2691);
and U7250 (N_7250,N_3216,N_2680);
nor U7251 (N_7251,N_4224,N_2721);
nor U7252 (N_7252,N_4457,N_3697);
nor U7253 (N_7253,N_4388,N_3223);
and U7254 (N_7254,N_4954,N_2508);
xnor U7255 (N_7255,N_2715,N_3361);
nor U7256 (N_7256,N_3907,N_2609);
nor U7257 (N_7257,N_3097,N_3739);
nor U7258 (N_7258,N_3043,N_2870);
and U7259 (N_7259,N_4237,N_4655);
and U7260 (N_7260,N_2605,N_4975);
and U7261 (N_7261,N_3525,N_3399);
xnor U7262 (N_7262,N_4813,N_4147);
and U7263 (N_7263,N_4219,N_2654);
or U7264 (N_7264,N_4025,N_4183);
nand U7265 (N_7265,N_4820,N_3532);
and U7266 (N_7266,N_3347,N_4694);
or U7267 (N_7267,N_2920,N_3425);
nand U7268 (N_7268,N_4987,N_4608);
nor U7269 (N_7269,N_4566,N_3267);
nor U7270 (N_7270,N_4269,N_4332);
nand U7271 (N_7271,N_4185,N_4099);
and U7272 (N_7272,N_4414,N_4277);
nor U7273 (N_7273,N_2687,N_2823);
nor U7274 (N_7274,N_4100,N_2594);
and U7275 (N_7275,N_4143,N_2639);
nor U7276 (N_7276,N_4363,N_3131);
nor U7277 (N_7277,N_2811,N_3413);
or U7278 (N_7278,N_3926,N_3372);
or U7279 (N_7279,N_3455,N_4712);
nand U7280 (N_7280,N_3120,N_2647);
nor U7281 (N_7281,N_2558,N_4260);
xnor U7282 (N_7282,N_3605,N_3795);
and U7283 (N_7283,N_3842,N_4714);
nand U7284 (N_7284,N_4113,N_3242);
nand U7285 (N_7285,N_3469,N_4470);
nor U7286 (N_7286,N_3398,N_4244);
or U7287 (N_7287,N_3412,N_4064);
nand U7288 (N_7288,N_3569,N_3551);
and U7289 (N_7289,N_2936,N_4557);
and U7290 (N_7290,N_2719,N_3055);
nor U7291 (N_7291,N_3457,N_3775);
or U7292 (N_7292,N_3296,N_2992);
xnor U7293 (N_7293,N_4577,N_2693);
nand U7294 (N_7294,N_3799,N_4585);
xor U7295 (N_7295,N_4413,N_3909);
nand U7296 (N_7296,N_2558,N_3513);
xnor U7297 (N_7297,N_4537,N_3221);
or U7298 (N_7298,N_2967,N_4467);
nor U7299 (N_7299,N_3987,N_4648);
or U7300 (N_7300,N_4231,N_4486);
and U7301 (N_7301,N_3839,N_4001);
nor U7302 (N_7302,N_3718,N_4224);
nand U7303 (N_7303,N_2602,N_3529);
xor U7304 (N_7304,N_3053,N_3455);
and U7305 (N_7305,N_2726,N_3748);
or U7306 (N_7306,N_3801,N_4264);
or U7307 (N_7307,N_4332,N_4873);
and U7308 (N_7308,N_4923,N_3459);
or U7309 (N_7309,N_3352,N_3103);
and U7310 (N_7310,N_4437,N_2715);
or U7311 (N_7311,N_3700,N_2728);
or U7312 (N_7312,N_3403,N_4499);
xor U7313 (N_7313,N_4678,N_4336);
xor U7314 (N_7314,N_2590,N_4885);
nor U7315 (N_7315,N_4732,N_2735);
or U7316 (N_7316,N_3955,N_3469);
and U7317 (N_7317,N_3708,N_3559);
nand U7318 (N_7318,N_4720,N_3515);
nand U7319 (N_7319,N_3174,N_4243);
or U7320 (N_7320,N_4520,N_2738);
and U7321 (N_7321,N_4803,N_4984);
xor U7322 (N_7322,N_4857,N_3483);
nor U7323 (N_7323,N_3338,N_2701);
nor U7324 (N_7324,N_3032,N_3407);
nand U7325 (N_7325,N_2580,N_3391);
nand U7326 (N_7326,N_4259,N_4290);
xnor U7327 (N_7327,N_3935,N_3222);
and U7328 (N_7328,N_2629,N_3898);
xor U7329 (N_7329,N_4367,N_2588);
nor U7330 (N_7330,N_4934,N_3883);
xnor U7331 (N_7331,N_3472,N_3942);
nand U7332 (N_7332,N_4842,N_4977);
or U7333 (N_7333,N_4976,N_3825);
nor U7334 (N_7334,N_3273,N_3837);
nand U7335 (N_7335,N_4772,N_2820);
nor U7336 (N_7336,N_4160,N_2956);
nand U7337 (N_7337,N_4222,N_4245);
or U7338 (N_7338,N_3070,N_3659);
and U7339 (N_7339,N_4346,N_3106);
nand U7340 (N_7340,N_4704,N_4041);
nand U7341 (N_7341,N_2554,N_4240);
and U7342 (N_7342,N_4031,N_4177);
xor U7343 (N_7343,N_4565,N_4635);
or U7344 (N_7344,N_3974,N_3391);
nand U7345 (N_7345,N_3014,N_4184);
or U7346 (N_7346,N_3554,N_3586);
nor U7347 (N_7347,N_4855,N_3242);
nand U7348 (N_7348,N_2547,N_2611);
nand U7349 (N_7349,N_4929,N_4902);
nor U7350 (N_7350,N_2858,N_2869);
xor U7351 (N_7351,N_4013,N_3273);
nand U7352 (N_7352,N_2802,N_3982);
and U7353 (N_7353,N_4893,N_3191);
and U7354 (N_7354,N_3904,N_2617);
nand U7355 (N_7355,N_4872,N_3767);
or U7356 (N_7356,N_3995,N_3288);
and U7357 (N_7357,N_3720,N_4177);
xor U7358 (N_7358,N_3392,N_4929);
or U7359 (N_7359,N_4014,N_4077);
nand U7360 (N_7360,N_3627,N_4104);
xor U7361 (N_7361,N_4110,N_3540);
and U7362 (N_7362,N_3350,N_3478);
xor U7363 (N_7363,N_3707,N_2882);
nor U7364 (N_7364,N_4482,N_4602);
and U7365 (N_7365,N_3783,N_3827);
xnor U7366 (N_7366,N_4143,N_3740);
and U7367 (N_7367,N_2607,N_3794);
nand U7368 (N_7368,N_3213,N_4396);
and U7369 (N_7369,N_3710,N_2908);
xor U7370 (N_7370,N_3031,N_3310);
xnor U7371 (N_7371,N_3659,N_3956);
and U7372 (N_7372,N_4198,N_4340);
nor U7373 (N_7373,N_4099,N_2654);
nand U7374 (N_7374,N_2966,N_3526);
or U7375 (N_7375,N_3826,N_4826);
nor U7376 (N_7376,N_4796,N_4695);
xnor U7377 (N_7377,N_4003,N_3750);
nor U7378 (N_7378,N_3723,N_3389);
or U7379 (N_7379,N_4191,N_4896);
nor U7380 (N_7380,N_3241,N_3026);
xnor U7381 (N_7381,N_2592,N_4929);
nand U7382 (N_7382,N_4850,N_2915);
nand U7383 (N_7383,N_4332,N_2899);
or U7384 (N_7384,N_2645,N_2582);
nand U7385 (N_7385,N_4174,N_3512);
nor U7386 (N_7386,N_4673,N_3294);
or U7387 (N_7387,N_3248,N_2695);
and U7388 (N_7388,N_3114,N_2919);
xor U7389 (N_7389,N_3405,N_2714);
and U7390 (N_7390,N_3723,N_4834);
and U7391 (N_7391,N_4383,N_4872);
xnor U7392 (N_7392,N_3606,N_3370);
xor U7393 (N_7393,N_3556,N_3332);
or U7394 (N_7394,N_4364,N_4975);
or U7395 (N_7395,N_3733,N_2678);
nor U7396 (N_7396,N_2810,N_4211);
nand U7397 (N_7397,N_3878,N_3796);
and U7398 (N_7398,N_4673,N_4075);
xor U7399 (N_7399,N_3033,N_2985);
nor U7400 (N_7400,N_4960,N_3292);
nand U7401 (N_7401,N_3432,N_3944);
xnor U7402 (N_7402,N_4001,N_3474);
xor U7403 (N_7403,N_3602,N_2733);
nor U7404 (N_7404,N_2969,N_4577);
xor U7405 (N_7405,N_4062,N_4165);
xor U7406 (N_7406,N_4815,N_3286);
and U7407 (N_7407,N_2730,N_3383);
or U7408 (N_7408,N_4193,N_4993);
nand U7409 (N_7409,N_3343,N_4264);
nand U7410 (N_7410,N_4420,N_2766);
and U7411 (N_7411,N_4242,N_2999);
and U7412 (N_7412,N_3881,N_4643);
nand U7413 (N_7413,N_4169,N_3439);
xnor U7414 (N_7414,N_2974,N_4019);
nand U7415 (N_7415,N_4200,N_3050);
and U7416 (N_7416,N_3843,N_3101);
xor U7417 (N_7417,N_4969,N_4510);
and U7418 (N_7418,N_2574,N_3612);
and U7419 (N_7419,N_3269,N_3200);
or U7420 (N_7420,N_2606,N_4356);
and U7421 (N_7421,N_4789,N_4939);
or U7422 (N_7422,N_4132,N_3912);
nand U7423 (N_7423,N_4289,N_2979);
or U7424 (N_7424,N_2610,N_3817);
or U7425 (N_7425,N_4920,N_2741);
nor U7426 (N_7426,N_4765,N_2825);
xnor U7427 (N_7427,N_2845,N_4639);
or U7428 (N_7428,N_3677,N_2689);
and U7429 (N_7429,N_3205,N_3758);
or U7430 (N_7430,N_3905,N_4691);
nand U7431 (N_7431,N_4901,N_3554);
and U7432 (N_7432,N_4906,N_2520);
and U7433 (N_7433,N_2799,N_4895);
or U7434 (N_7434,N_3938,N_4531);
or U7435 (N_7435,N_2953,N_4551);
or U7436 (N_7436,N_4741,N_4804);
nor U7437 (N_7437,N_3482,N_4564);
or U7438 (N_7438,N_3624,N_4211);
and U7439 (N_7439,N_3680,N_3817);
and U7440 (N_7440,N_4418,N_2747);
xor U7441 (N_7441,N_3401,N_3128);
nor U7442 (N_7442,N_3203,N_4233);
nand U7443 (N_7443,N_2552,N_4591);
xor U7444 (N_7444,N_3604,N_4293);
and U7445 (N_7445,N_2807,N_4926);
or U7446 (N_7446,N_4459,N_2566);
and U7447 (N_7447,N_3356,N_3110);
or U7448 (N_7448,N_3044,N_3131);
nand U7449 (N_7449,N_3019,N_3824);
nor U7450 (N_7450,N_4255,N_4262);
xnor U7451 (N_7451,N_2786,N_3424);
and U7452 (N_7452,N_4462,N_3892);
nor U7453 (N_7453,N_4606,N_4717);
and U7454 (N_7454,N_4394,N_4333);
and U7455 (N_7455,N_4168,N_3561);
nor U7456 (N_7456,N_2864,N_3577);
or U7457 (N_7457,N_3745,N_4066);
nand U7458 (N_7458,N_4357,N_3178);
or U7459 (N_7459,N_4493,N_4628);
or U7460 (N_7460,N_2806,N_2914);
or U7461 (N_7461,N_3155,N_3499);
xnor U7462 (N_7462,N_3933,N_2671);
nand U7463 (N_7463,N_4339,N_3272);
xnor U7464 (N_7464,N_3534,N_3178);
and U7465 (N_7465,N_3680,N_3900);
or U7466 (N_7466,N_4896,N_3136);
nand U7467 (N_7467,N_2517,N_4791);
and U7468 (N_7468,N_4606,N_2889);
xnor U7469 (N_7469,N_3449,N_2967);
or U7470 (N_7470,N_3619,N_4663);
and U7471 (N_7471,N_2930,N_3310);
nor U7472 (N_7472,N_3756,N_4923);
xnor U7473 (N_7473,N_4139,N_3332);
or U7474 (N_7474,N_3338,N_3816);
and U7475 (N_7475,N_2851,N_4064);
nand U7476 (N_7476,N_2974,N_3245);
nor U7477 (N_7477,N_3387,N_3028);
or U7478 (N_7478,N_4772,N_2917);
xnor U7479 (N_7479,N_2682,N_3534);
nor U7480 (N_7480,N_4174,N_2768);
nor U7481 (N_7481,N_3093,N_4572);
nor U7482 (N_7482,N_3557,N_3988);
nand U7483 (N_7483,N_3605,N_4788);
xor U7484 (N_7484,N_3633,N_3458);
nand U7485 (N_7485,N_2812,N_3226);
nor U7486 (N_7486,N_3693,N_2676);
and U7487 (N_7487,N_3563,N_2857);
nor U7488 (N_7488,N_3856,N_2724);
xor U7489 (N_7489,N_3706,N_4856);
or U7490 (N_7490,N_3925,N_3912);
and U7491 (N_7491,N_4835,N_3299);
nor U7492 (N_7492,N_3522,N_3569);
nand U7493 (N_7493,N_3664,N_3940);
nor U7494 (N_7494,N_4123,N_2969);
nand U7495 (N_7495,N_3551,N_4890);
xor U7496 (N_7496,N_4007,N_3480);
nor U7497 (N_7497,N_3822,N_3684);
nor U7498 (N_7498,N_4323,N_4456);
nor U7499 (N_7499,N_4228,N_4725);
or U7500 (N_7500,N_5714,N_7300);
nor U7501 (N_7501,N_6039,N_6111);
nand U7502 (N_7502,N_6407,N_5899);
nand U7503 (N_7503,N_7354,N_5344);
nand U7504 (N_7504,N_6623,N_5825);
nor U7505 (N_7505,N_6310,N_5522);
nor U7506 (N_7506,N_6506,N_6068);
and U7507 (N_7507,N_5517,N_5771);
nand U7508 (N_7508,N_6665,N_6867);
xnor U7509 (N_7509,N_5859,N_5911);
nor U7510 (N_7510,N_6852,N_6544);
nor U7511 (N_7511,N_6466,N_5726);
and U7512 (N_7512,N_6619,N_5834);
nor U7513 (N_7513,N_5286,N_7419);
and U7514 (N_7514,N_5419,N_7049);
nand U7515 (N_7515,N_7236,N_6204);
or U7516 (N_7516,N_7175,N_7367);
and U7517 (N_7517,N_5040,N_6315);
xor U7518 (N_7518,N_5501,N_7349);
nor U7519 (N_7519,N_6216,N_5083);
nand U7520 (N_7520,N_6255,N_5128);
and U7521 (N_7521,N_7075,N_5959);
nand U7522 (N_7522,N_6313,N_6300);
or U7523 (N_7523,N_5023,N_6803);
or U7524 (N_7524,N_6819,N_6613);
and U7525 (N_7525,N_7216,N_5743);
nor U7526 (N_7526,N_6228,N_5674);
xnor U7527 (N_7527,N_6994,N_6515);
and U7528 (N_7528,N_7228,N_7151);
xnor U7529 (N_7529,N_7482,N_6692);
nor U7530 (N_7530,N_5394,N_7293);
nand U7531 (N_7531,N_6268,N_5373);
nand U7532 (N_7532,N_7222,N_5681);
or U7533 (N_7533,N_6545,N_6184);
xnor U7534 (N_7534,N_6316,N_6185);
xor U7535 (N_7535,N_5875,N_5695);
nand U7536 (N_7536,N_6174,N_5592);
xnor U7537 (N_7537,N_7043,N_5229);
nand U7538 (N_7538,N_6909,N_5043);
xor U7539 (N_7539,N_6723,N_5256);
or U7540 (N_7540,N_6259,N_7009);
and U7541 (N_7541,N_7291,N_5576);
xnor U7542 (N_7542,N_7240,N_5379);
and U7543 (N_7543,N_5730,N_5417);
xnor U7544 (N_7544,N_5577,N_6203);
and U7545 (N_7545,N_5526,N_5039);
nor U7546 (N_7546,N_7350,N_7424);
nand U7547 (N_7547,N_5182,N_7427);
nand U7548 (N_7548,N_7429,N_5346);
and U7549 (N_7549,N_6575,N_5782);
and U7550 (N_7550,N_5766,N_5369);
nor U7551 (N_7551,N_6114,N_7130);
xnor U7552 (N_7552,N_5007,N_6304);
nand U7553 (N_7553,N_6060,N_6085);
or U7554 (N_7554,N_7341,N_7188);
and U7555 (N_7555,N_6705,N_7003);
and U7556 (N_7556,N_5560,N_6420);
or U7557 (N_7557,N_5388,N_5786);
nor U7558 (N_7558,N_6715,N_6726);
nand U7559 (N_7559,N_6707,N_7452);
xnor U7560 (N_7560,N_6886,N_6498);
xnor U7561 (N_7561,N_6598,N_6195);
xor U7562 (N_7562,N_6198,N_6235);
xor U7563 (N_7563,N_7475,N_5655);
nand U7564 (N_7564,N_6532,N_6236);
and U7565 (N_7565,N_6211,N_5846);
or U7566 (N_7566,N_6059,N_6131);
xor U7567 (N_7567,N_6787,N_5968);
nor U7568 (N_7568,N_5324,N_5853);
or U7569 (N_7569,N_5937,N_7356);
xor U7570 (N_7570,N_6221,N_6344);
nor U7571 (N_7571,N_6824,N_6234);
nor U7572 (N_7572,N_5964,N_6584);
xor U7573 (N_7573,N_7466,N_6943);
xor U7574 (N_7574,N_5066,N_5919);
or U7575 (N_7575,N_5126,N_7468);
and U7576 (N_7576,N_6642,N_6999);
or U7577 (N_7577,N_6468,N_5842);
nand U7578 (N_7578,N_5248,N_7083);
nand U7579 (N_7579,N_5198,N_5262);
or U7580 (N_7580,N_7239,N_5214);
or U7581 (N_7581,N_5979,N_6434);
nor U7582 (N_7582,N_6731,N_7262);
or U7583 (N_7583,N_7290,N_5824);
nand U7584 (N_7584,N_7160,N_6855);
nand U7585 (N_7585,N_5057,N_6166);
and U7586 (N_7586,N_6423,N_5226);
and U7587 (N_7587,N_5191,N_5787);
and U7588 (N_7588,N_7401,N_5727);
nor U7589 (N_7589,N_5200,N_5861);
xor U7590 (N_7590,N_7076,N_7062);
and U7591 (N_7591,N_5199,N_7000);
xnor U7592 (N_7592,N_5579,N_6997);
and U7593 (N_7593,N_6249,N_5272);
nand U7594 (N_7594,N_5116,N_5996);
or U7595 (N_7595,N_7238,N_5733);
and U7596 (N_7596,N_5235,N_6818);
or U7597 (N_7597,N_5542,N_5048);
or U7598 (N_7598,N_5932,N_5147);
nor U7599 (N_7599,N_5012,N_5016);
nor U7600 (N_7600,N_6158,N_7321);
xor U7601 (N_7601,N_7057,N_7232);
nor U7602 (N_7602,N_7071,N_6928);
and U7603 (N_7603,N_5575,N_5459);
nand U7604 (N_7604,N_5564,N_6321);
nor U7605 (N_7605,N_5600,N_6154);
and U7606 (N_7606,N_7423,N_6858);
and U7607 (N_7607,N_7324,N_5947);
xor U7608 (N_7608,N_5990,N_5018);
nor U7609 (N_7609,N_6581,N_5682);
or U7610 (N_7610,N_6242,N_5967);
or U7611 (N_7611,N_6412,N_6795);
nor U7612 (N_7612,N_5294,N_6295);
and U7613 (N_7613,N_7444,N_5120);
and U7614 (N_7614,N_6853,N_5903);
xnor U7615 (N_7615,N_6654,N_6659);
nor U7616 (N_7616,N_7348,N_5829);
nand U7617 (N_7617,N_6934,N_6605);
or U7618 (N_7618,N_6695,N_7085);
and U7619 (N_7619,N_5372,N_5547);
or U7620 (N_7620,N_5339,N_6370);
or U7621 (N_7621,N_5512,N_5795);
xnor U7622 (N_7622,N_5744,N_7335);
xor U7623 (N_7623,N_6611,N_7019);
nor U7624 (N_7624,N_6820,N_5506);
nand U7625 (N_7625,N_6979,N_6981);
xnor U7626 (N_7626,N_6583,N_5046);
nand U7627 (N_7627,N_6212,N_7089);
nand U7628 (N_7628,N_7208,N_6920);
nor U7629 (N_7629,N_6708,N_5411);
nand U7630 (N_7630,N_6067,N_6922);
xor U7631 (N_7631,N_7060,N_7244);
and U7632 (N_7632,N_7394,N_5127);
or U7633 (N_7633,N_6863,N_5953);
or U7634 (N_7634,N_5789,N_6021);
and U7635 (N_7635,N_5431,N_6157);
nor U7636 (N_7636,N_6938,N_7195);
and U7637 (N_7637,N_6500,N_5240);
nand U7638 (N_7638,N_5595,N_6163);
nand U7639 (N_7639,N_6082,N_6034);
and U7640 (N_7640,N_7385,N_6550);
or U7641 (N_7641,N_5383,N_6908);
nor U7642 (N_7642,N_5278,N_5654);
and U7643 (N_7643,N_5275,N_6594);
and U7644 (N_7644,N_7231,N_5849);
xor U7645 (N_7645,N_5347,N_6509);
nor U7646 (N_7646,N_6200,N_5180);
nor U7647 (N_7647,N_5923,N_5397);
and U7648 (N_7648,N_6856,N_7126);
and U7649 (N_7649,N_6124,N_6366);
or U7650 (N_7650,N_5669,N_5203);
or U7651 (N_7651,N_5683,N_6520);
nand U7652 (N_7652,N_5457,N_5939);
or U7653 (N_7653,N_5644,N_7458);
xnor U7654 (N_7654,N_5178,N_5585);
xor U7655 (N_7655,N_5319,N_5905);
and U7656 (N_7656,N_5772,N_7398);
nand U7657 (N_7657,N_5101,N_5831);
and U7658 (N_7658,N_5232,N_7146);
and U7659 (N_7659,N_5086,N_7357);
or U7660 (N_7660,N_5550,N_5282);
nand U7661 (N_7661,N_5307,N_5629);
or U7662 (N_7662,N_6456,N_6968);
and U7663 (N_7663,N_6209,N_6368);
and U7664 (N_7664,N_6190,N_6260);
and U7665 (N_7665,N_6971,N_6005);
or U7666 (N_7666,N_5426,N_5395);
nor U7667 (N_7667,N_7337,N_6254);
or U7668 (N_7668,N_7194,N_7097);
nand U7669 (N_7669,N_6749,N_6038);
and U7670 (N_7670,N_6877,N_5804);
nor U7671 (N_7671,N_7391,N_7001);
xor U7672 (N_7672,N_6391,N_6066);
and U7673 (N_7673,N_6014,N_6961);
and U7674 (N_7674,N_5944,N_7039);
nand U7675 (N_7675,N_5409,N_6698);
nor U7676 (N_7676,N_5485,N_6006);
xor U7677 (N_7677,N_6686,N_6789);
or U7678 (N_7678,N_5455,N_6057);
xnor U7679 (N_7679,N_5099,N_5796);
xnor U7680 (N_7680,N_7338,N_5156);
nand U7681 (N_7681,N_6670,N_5357);
xnor U7682 (N_7682,N_6663,N_5895);
or U7683 (N_7683,N_5341,N_6574);
or U7684 (N_7684,N_6828,N_7305);
nor U7685 (N_7685,N_6278,N_6056);
nand U7686 (N_7686,N_6411,N_7055);
nand U7687 (N_7687,N_6972,N_5640);
xnor U7688 (N_7688,N_5537,N_6293);
xor U7689 (N_7689,N_5152,N_6556);
nand U7690 (N_7690,N_5111,N_5699);
nor U7691 (N_7691,N_6524,N_7371);
or U7692 (N_7692,N_5225,N_7311);
or U7693 (N_7693,N_6587,N_7431);
and U7694 (N_7694,N_5260,N_5231);
and U7695 (N_7695,N_5352,N_6284);
and U7696 (N_7696,N_5348,N_6491);
and U7697 (N_7697,N_5428,N_6948);
xor U7698 (N_7698,N_6340,N_6449);
xor U7699 (N_7699,N_6873,N_5025);
and U7700 (N_7700,N_5195,N_6135);
nor U7701 (N_7701,N_5488,N_5193);
or U7702 (N_7702,N_5252,N_6764);
xnor U7703 (N_7703,N_5927,N_6075);
xor U7704 (N_7704,N_5472,N_7428);
or U7705 (N_7705,N_7246,N_6120);
nor U7706 (N_7706,N_5407,N_5499);
or U7707 (N_7707,N_5885,N_6936);
xor U7708 (N_7708,N_6826,N_5423);
and U7709 (N_7709,N_6843,N_5335);
nand U7710 (N_7710,N_5219,N_5138);
nor U7711 (N_7711,N_5597,N_5429);
nor U7712 (N_7712,N_7045,N_7140);
and U7713 (N_7713,N_6088,N_7110);
or U7714 (N_7714,N_6722,N_5011);
nand U7715 (N_7715,N_7365,N_5561);
and U7716 (N_7716,N_5239,N_5777);
xor U7717 (N_7717,N_5509,N_6232);
nand U7718 (N_7718,N_6586,N_7027);
or U7719 (N_7719,N_5162,N_7221);
or U7720 (N_7720,N_5545,N_6918);
nand U7721 (N_7721,N_5773,N_5345);
nand U7722 (N_7722,N_6339,N_6808);
nand U7723 (N_7723,N_5943,N_5500);
and U7724 (N_7724,N_6213,N_5211);
nand U7725 (N_7725,N_5879,N_5053);
xnor U7726 (N_7726,N_6274,N_7199);
and U7727 (N_7727,N_5461,N_7494);
nor U7728 (N_7728,N_5438,N_6827);
nor U7729 (N_7729,N_6342,N_6256);
nor U7730 (N_7730,N_5364,N_7281);
xnor U7731 (N_7731,N_5360,N_6530);
nand U7732 (N_7732,N_7314,N_5150);
nor U7733 (N_7733,N_7414,N_6777);
or U7734 (N_7734,N_5481,N_7181);
nor U7735 (N_7735,N_6429,N_7326);
or U7736 (N_7736,N_5737,N_5188);
and U7737 (N_7737,N_6016,N_5452);
nand U7738 (N_7738,N_6071,N_6878);
and U7739 (N_7739,N_5008,N_5054);
xnor U7740 (N_7740,N_7416,N_5848);
nor U7741 (N_7741,N_6964,N_5015);
nand U7742 (N_7742,N_7355,N_6298);
xnor U7743 (N_7743,N_6164,N_5062);
or U7744 (N_7744,N_6589,N_6288);
nor U7745 (N_7745,N_7380,N_7041);
nor U7746 (N_7746,N_6849,N_5762);
nor U7747 (N_7747,N_5873,N_5986);
xor U7748 (N_7748,N_6165,N_6664);
or U7749 (N_7749,N_6469,N_5857);
and U7750 (N_7750,N_6739,N_6330);
xor U7751 (N_7751,N_7488,N_6261);
nand U7752 (N_7752,N_5724,N_6635);
and U7753 (N_7753,N_7363,N_7167);
xnor U7754 (N_7754,N_7172,N_6489);
nor U7755 (N_7755,N_6568,N_7226);
nor U7756 (N_7756,N_7455,N_6769);
xor U7757 (N_7757,N_5165,N_5814);
and U7758 (N_7758,N_7020,N_5504);
and U7759 (N_7759,N_6326,N_6167);
xnor U7760 (N_7760,N_5149,N_6650);
xor U7761 (N_7761,N_6810,N_5807);
nand U7762 (N_7762,N_6329,N_7498);
xor U7763 (N_7763,N_6813,N_6176);
and U7764 (N_7764,N_7058,N_6269);
or U7765 (N_7765,N_7042,N_5440);
or U7766 (N_7766,N_6450,N_7315);
or U7767 (N_7767,N_6227,N_6406);
xnor U7768 (N_7768,N_5616,N_6360);
nand U7769 (N_7769,N_7472,N_5261);
or U7770 (N_7770,N_5569,N_5869);
nand U7771 (N_7771,N_6998,N_7190);
nand U7772 (N_7772,N_7292,N_5477);
nor U7773 (N_7773,N_5708,N_5233);
or U7774 (N_7774,N_5338,N_5966);
or U7775 (N_7775,N_6473,N_6779);
nor U7776 (N_7776,N_7400,N_5247);
nor U7777 (N_7777,N_6788,N_5478);
nor U7778 (N_7778,N_7440,N_6404);
nand U7779 (N_7779,N_5572,N_7191);
nand U7780 (N_7780,N_6400,N_5552);
xnor U7781 (N_7781,N_5755,N_7285);
xor U7782 (N_7782,N_6662,N_6570);
and U7783 (N_7783,N_7344,N_5029);
and U7784 (N_7784,N_5113,N_6751);
or U7785 (N_7785,N_6446,N_5776);
and U7786 (N_7786,N_6554,N_7170);
nand U7787 (N_7787,N_6015,N_6512);
and U7788 (N_7788,N_7013,N_7277);
or U7789 (N_7789,N_6730,N_6929);
nand U7790 (N_7790,N_6323,N_5001);
nor U7791 (N_7791,N_5168,N_5610);
and U7792 (N_7792,N_6561,N_6864);
xor U7793 (N_7793,N_5562,N_6035);
nor U7794 (N_7794,N_6175,N_5328);
xor U7795 (N_7795,N_5502,N_5874);
nor U7796 (N_7796,N_5798,N_6053);
or U7797 (N_7797,N_6794,N_5377);
or U7798 (N_7798,N_5183,N_7180);
xor U7799 (N_7799,N_7374,N_5672);
or U7800 (N_7800,N_6384,N_5822);
and U7801 (N_7801,N_5535,N_7064);
or U7802 (N_7802,N_5624,N_5693);
or U7803 (N_7803,N_6651,N_7050);
or U7804 (N_7804,N_5622,N_6762);
nor U7805 (N_7805,N_5516,N_7405);
or U7806 (N_7806,N_7382,N_6048);
nor U7807 (N_7807,N_6714,N_6237);
xor U7808 (N_7808,N_7259,N_6866);
xor U7809 (N_7809,N_5055,N_5720);
nor U7810 (N_7810,N_5482,N_6387);
xor U7811 (N_7811,N_6292,N_5618);
and U7812 (N_7812,N_6092,N_5106);
nor U7813 (N_7813,N_5729,N_6697);
and U7814 (N_7814,N_5034,N_6311);
nand U7815 (N_7815,N_6258,N_5003);
nand U7816 (N_7816,N_5525,N_5531);
nand U7817 (N_7817,N_5074,N_7462);
and U7818 (N_7818,N_5258,N_6403);
xor U7819 (N_7819,N_6266,N_6986);
xnor U7820 (N_7820,N_7063,N_5659);
nor U7821 (N_7821,N_7031,N_7411);
and U7822 (N_7822,N_5541,N_6952);
nor U7823 (N_7823,N_6746,N_6193);
and U7824 (N_7824,N_5738,N_6752);
and U7825 (N_7825,N_7250,N_7484);
nor U7826 (N_7826,N_5573,N_7052);
nand U7827 (N_7827,N_7212,N_6540);
xor U7828 (N_7828,N_6401,N_5170);
xor U7829 (N_7829,N_6253,N_6481);
nand U7830 (N_7830,N_6433,N_6263);
and U7831 (N_7831,N_6634,N_5378);
nor U7832 (N_7832,N_5255,N_6478);
nor U7833 (N_7833,N_6600,N_5942);
nor U7834 (N_7834,N_5089,N_5356);
nor U7835 (N_7835,N_7093,N_5920);
or U7836 (N_7836,N_5746,N_5975);
and U7837 (N_7837,N_5420,N_5507);
and U7838 (N_7838,N_7164,N_6501);
nor U7839 (N_7839,N_6197,N_6012);
and U7840 (N_7840,N_6771,N_7119);
and U7841 (N_7841,N_6703,N_6086);
or U7842 (N_7842,N_5632,N_6628);
xor U7843 (N_7843,N_6632,N_6917);
xnor U7844 (N_7844,N_7149,N_6748);
nor U7845 (N_7845,N_6815,N_5320);
and U7846 (N_7846,N_5004,N_6439);
xnor U7847 (N_7847,N_6912,N_6743);
or U7848 (N_7848,N_5835,N_5530);
nor U7849 (N_7849,N_6924,N_5483);
and U7850 (N_7850,N_5940,N_5072);
nand U7851 (N_7851,N_6693,N_7456);
nand U7852 (N_7852,N_5279,N_5867);
nand U7853 (N_7853,N_7322,N_7378);
xnor U7854 (N_7854,N_6658,N_6606);
or U7855 (N_7855,N_6050,N_7198);
and U7856 (N_7856,N_7123,N_5930);
nor U7857 (N_7857,N_5056,N_5151);
or U7858 (N_7858,N_7430,N_5936);
nor U7859 (N_7859,N_7490,N_5910);
xnor U7860 (N_7860,N_7203,N_5578);
and U7861 (N_7861,N_6095,N_6438);
xor U7862 (N_7862,N_5172,N_6685);
nor U7863 (N_7863,N_7446,N_6537);
or U7864 (N_7864,N_7032,N_7028);
xnor U7865 (N_7865,N_5756,N_5900);
and U7866 (N_7866,N_6508,N_5163);
nor U7867 (N_7867,N_5337,N_6440);
and U7868 (N_7868,N_5297,N_6499);
nor U7869 (N_7869,N_5623,N_5761);
and U7870 (N_7870,N_5995,N_6962);
and U7871 (N_7871,N_7183,N_7156);
nor U7872 (N_7872,N_5238,N_6025);
nand U7873 (N_7873,N_5989,N_6416);
or U7874 (N_7874,N_6895,N_6425);
xor U7875 (N_7875,N_5021,N_7451);
and U7876 (N_7876,N_5480,N_7131);
xor U7877 (N_7877,N_7016,N_6062);
and U7878 (N_7878,N_5157,N_5104);
nor U7879 (N_7879,N_7068,N_6987);
or U7880 (N_7880,N_6797,N_7496);
and U7881 (N_7881,N_7359,N_5915);
nor U7882 (N_7882,N_6270,N_6458);
xor U7883 (N_7883,N_5177,N_5608);
or U7884 (N_7884,N_6527,N_6984);
or U7885 (N_7885,N_7454,N_5148);
or U7886 (N_7886,N_5076,N_6139);
and U7887 (N_7887,N_5811,N_6955);
xor U7888 (N_7888,N_5747,N_7173);
xnor U7889 (N_7889,N_6474,N_5665);
nor U7890 (N_7890,N_6620,N_6141);
nor U7891 (N_7891,N_5223,N_6428);
and U7892 (N_7892,N_5768,N_7258);
xnor U7893 (N_7893,N_5167,N_6100);
nand U7894 (N_7894,N_5902,N_7495);
xnor U7895 (N_7895,N_6890,N_6960);
xnor U7896 (N_7896,N_7092,N_7395);
nor U7897 (N_7897,N_7298,N_7105);
xor U7898 (N_7898,N_5553,N_6279);
nand U7899 (N_7899,N_6381,N_6098);
and U7900 (N_7900,N_7121,N_5767);
and U7901 (N_7901,N_7426,N_6893);
nand U7902 (N_7902,N_6152,N_7267);
xor U7903 (N_7903,N_5636,N_6225);
or U7904 (N_7904,N_6365,N_7485);
nand U7905 (N_7905,N_6240,N_5268);
or U7906 (N_7906,N_5494,N_7421);
xor U7907 (N_7907,N_6622,N_6982);
nor U7908 (N_7908,N_6364,N_5589);
or U7909 (N_7909,N_6954,N_5391);
xor U7910 (N_7910,N_6402,N_7487);
or U7911 (N_7911,N_7215,N_6717);
xor U7912 (N_7912,N_5121,N_5605);
and U7913 (N_7913,N_7408,N_6709);
nand U7914 (N_7914,N_6023,N_5131);
xor U7915 (N_7915,N_5792,N_6729);
nand U7916 (N_7916,N_7409,N_6058);
and U7917 (N_7917,N_6689,N_7320);
nand U7918 (N_7918,N_5412,N_5715);
nor U7919 (N_7919,N_5628,N_6410);
or U7920 (N_7920,N_5489,N_7393);
and U7921 (N_7921,N_6345,N_6539);
nor U7922 (N_7922,N_5006,N_5449);
nand U7923 (N_7923,N_5565,N_5122);
xor U7924 (N_7924,N_6522,N_6367);
nand U7925 (N_7925,N_6244,N_5549);
nand U7926 (N_7926,N_7273,N_6140);
xor U7927 (N_7927,N_5241,N_5141);
nand U7928 (N_7928,N_5495,N_5819);
nor U7929 (N_7929,N_5087,N_6105);
xor U7930 (N_7930,N_7390,N_7008);
nand U7931 (N_7931,N_6842,N_7345);
nand U7932 (N_7932,N_6335,N_5706);
nor U7933 (N_7933,N_5118,N_5047);
or U7934 (N_7934,N_5556,N_5581);
and U7935 (N_7935,N_5991,N_6201);
nand U7936 (N_7936,N_5090,N_6396);
nor U7937 (N_7937,N_6923,N_5791);
nand U7938 (N_7938,N_7274,N_5441);
or U7939 (N_7939,N_6621,N_5709);
and U7940 (N_7940,N_5263,N_6042);
xnor U7941 (N_7941,N_6661,N_5559);
and U7942 (N_7942,N_5361,N_5974);
nand U7943 (N_7943,N_6459,N_7422);
nor U7944 (N_7944,N_5336,N_5664);
nor U7945 (N_7945,N_5958,N_5688);
nor U7946 (N_7946,N_6040,N_6302);
or U7947 (N_7947,N_5886,N_6845);
or U7948 (N_7948,N_6182,N_6250);
or U7949 (N_7949,N_6393,N_7383);
and U7950 (N_7950,N_6355,N_6590);
nor U7951 (N_7951,N_5742,N_6711);
nand U7952 (N_7952,N_5826,N_5137);
or U7953 (N_7953,N_7251,N_5458);
nand U7954 (N_7954,N_7152,N_6445);
and U7955 (N_7955,N_7272,N_5926);
or U7956 (N_7956,N_7330,N_5197);
nor U7957 (N_7957,N_7325,N_7117);
xor U7958 (N_7958,N_5933,N_5566);
or U7959 (N_7959,N_6737,N_5080);
and U7960 (N_7960,N_6388,N_6690);
and U7961 (N_7961,N_7286,N_5368);
xnor U7962 (N_7962,N_6937,N_6102);
nor U7963 (N_7963,N_6875,N_5856);
nand U7964 (N_7964,N_5702,N_6353);
nor U7965 (N_7965,N_6980,N_5471);
and U7966 (N_7966,N_5365,N_6636);
and U7967 (N_7967,N_7005,N_7189);
and U7968 (N_7968,N_6989,N_5060);
or U7969 (N_7969,N_7201,N_6538);
nor U7970 (N_7970,N_5901,N_5928);
and U7971 (N_7971,N_7474,N_5684);
and U7972 (N_7972,N_5273,N_5434);
or U7973 (N_7973,N_6966,N_5703);
nand U7974 (N_7974,N_5298,N_7407);
nor U7975 (N_7975,N_5783,N_7479);
nor U7976 (N_7976,N_5960,N_5073);
and U7977 (N_7977,N_7271,N_6517);
or U7978 (N_7978,N_6065,N_5265);
or U7979 (N_7979,N_5408,N_6780);
or U7980 (N_7980,N_7051,N_6026);
nor U7981 (N_7981,N_6683,N_7403);
xor U7982 (N_7982,N_5031,N_5518);
or U7983 (N_7983,N_5643,N_6694);
or U7984 (N_7984,N_6983,N_6900);
or U7985 (N_7985,N_6944,N_5027);
nor U7986 (N_7986,N_6325,N_6493);
nand U7987 (N_7987,N_6847,N_6626);
nand U7988 (N_7988,N_6533,N_5567);
or U7989 (N_7989,N_5888,N_5650);
nand U7990 (N_7990,N_7415,N_6884);
and U7991 (N_7991,N_6881,N_6108);
xnor U7992 (N_7992,N_5267,N_6734);
or U7993 (N_7993,N_7059,N_5405);
and U7994 (N_7994,N_6080,N_7388);
xnor U7995 (N_7995,N_5951,N_5770);
and U7996 (N_7996,N_5571,N_5082);
nor U7997 (N_7997,N_5588,N_5295);
and U7998 (N_7998,N_5350,N_7284);
nor U7999 (N_7999,N_5467,N_6186);
or U8000 (N_8000,N_6147,N_5310);
or U8001 (N_8001,N_5583,N_7230);
nand U8002 (N_8002,N_5963,N_5515);
nor U8003 (N_8003,N_7288,N_6482);
xor U8004 (N_8004,N_6348,N_5555);
nor U8005 (N_8005,N_7214,N_5897);
xor U8006 (N_8006,N_7030,N_6338);
nor U8007 (N_8007,N_5815,N_5002);
and U8008 (N_8008,N_6888,N_7247);
nor U8009 (N_8009,N_6671,N_6931);
xnor U8010 (N_8010,N_6432,N_5331);
or U8011 (N_8011,N_6170,N_7346);
and U8012 (N_8012,N_7477,N_6541);
nand U8013 (N_8013,N_6032,N_6076);
nor U8014 (N_8014,N_5889,N_6871);
and U8015 (N_8015,N_6118,N_6578);
nor U8016 (N_8016,N_6046,N_6872);
nor U8017 (N_8017,N_5833,N_5318);
or U8018 (N_8018,N_5642,N_6914);
nand U8019 (N_8019,N_6514,N_7373);
or U8020 (N_8020,N_5717,N_7497);
and U8021 (N_8021,N_7480,N_5539);
nor U8022 (N_8022,N_6666,N_6816);
and U8023 (N_8023,N_6985,N_6935);
or U8024 (N_8024,N_6319,N_6463);
or U8025 (N_8025,N_6418,N_7006);
nand U8026 (N_8026,N_6303,N_5802);
nand U8027 (N_8027,N_6835,N_6899);
xnor U8028 (N_8028,N_7361,N_7033);
nor U8029 (N_8029,N_6798,N_5329);
nand U8030 (N_8030,N_5700,N_6639);
xnor U8031 (N_8031,N_7307,N_6146);
xor U8032 (N_8032,N_7243,N_5266);
xor U8033 (N_8033,N_6030,N_5317);
nor U8034 (N_8034,N_6320,N_6129);
xor U8035 (N_8035,N_7370,N_6691);
nor U8036 (N_8036,N_6510,N_7264);
or U8037 (N_8037,N_7137,N_5723);
or U8038 (N_8038,N_5332,N_5460);
or U8039 (N_8039,N_7220,N_7372);
nor U8040 (N_8040,N_6281,N_5257);
and U8041 (N_8041,N_6959,N_5051);
nor U8042 (N_8042,N_5067,N_6045);
nor U8043 (N_8043,N_5330,N_7148);
xnor U8044 (N_8044,N_7491,N_7025);
nor U8045 (N_8045,N_5443,N_7011);
or U8046 (N_8046,N_5399,N_7319);
or U8047 (N_8047,N_5841,N_6887);
nor U8048 (N_8048,N_6471,N_6003);
nand U8049 (N_8049,N_5732,N_5558);
nor U8050 (N_8050,N_5028,N_5865);
xor U8051 (N_8051,N_5037,N_5221);
nor U8052 (N_8052,N_5403,N_5679);
xor U8053 (N_8053,N_5353,N_7317);
xor U8054 (N_8054,N_6248,N_5992);
and U8055 (N_8055,N_5251,N_5680);
nor U8056 (N_8056,N_6728,N_7309);
xnor U8057 (N_8057,N_5097,N_7099);
nand U8058 (N_8058,N_6783,N_5444);
nand U8059 (N_8059,N_5845,N_5314);
nor U8060 (N_8060,N_7369,N_6906);
nor U8061 (N_8061,N_6812,N_5620);
nor U8062 (N_8062,N_5342,N_6460);
nand U8063 (N_8063,N_7169,N_6868);
nor U8064 (N_8064,N_6051,N_7332);
nand U8065 (N_8065,N_6307,N_6667);
xor U8066 (N_8066,N_5827,N_5625);
and U8067 (N_8067,N_6609,N_7275);
nor U8068 (N_8068,N_6566,N_6825);
xor U8069 (N_8069,N_6317,N_5019);
nand U8070 (N_8070,N_5918,N_5862);
or U8071 (N_8071,N_5748,N_5883);
xnor U8072 (N_8072,N_5741,N_5249);
xnor U8073 (N_8073,N_5977,N_6882);
or U8074 (N_8074,N_5400,N_6245);
and U8075 (N_8075,N_5705,N_7268);
xor U8076 (N_8076,N_6097,N_5830);
nor U8077 (N_8077,N_5590,N_6072);
xor U8078 (N_8078,N_6821,N_5631);
or U8079 (N_8079,N_6916,N_5102);
nand U8080 (N_8080,N_5646,N_6738);
xor U8081 (N_8081,N_7360,N_5645);
xor U8082 (N_8082,N_5095,N_5637);
nor U8083 (N_8083,N_7182,N_5769);
or U8084 (N_8084,N_5010,N_5925);
or U8085 (N_8085,N_6552,N_5586);
nor U8086 (N_8086,N_5366,N_7023);
nor U8087 (N_8087,N_6484,N_6949);
and U8088 (N_8088,N_6133,N_5921);
or U8089 (N_8089,N_7340,N_6945);
and U8090 (N_8090,N_6442,N_5981);
nand U8091 (N_8091,N_6331,N_6010);
and U8092 (N_8092,N_6419,N_6024);
xnor U8093 (N_8093,N_5511,N_5326);
and U8094 (N_8094,N_6103,N_6940);
and U8095 (N_8095,N_5492,N_5949);
nand U8096 (N_8096,N_7095,N_5957);
xnor U8097 (N_8097,N_6155,N_6398);
nand U8098 (N_8098,N_6956,N_6207);
nor U8099 (N_8099,N_7193,N_6421);
and U8100 (N_8100,N_7046,N_6294);
and U8101 (N_8101,N_6297,N_5956);
xor U8102 (N_8102,N_5532,N_6905);
nand U8103 (N_8103,N_6678,N_5433);
nand U8104 (N_8104,N_5253,N_6385);
and U8105 (N_8105,N_5988,N_5496);
or U8106 (N_8106,N_5917,N_5064);
nand U8107 (N_8107,N_5976,N_5662);
or U8108 (N_8108,N_5005,N_7015);
nor U8109 (N_8109,N_5134,N_5685);
or U8110 (N_8110,N_6631,N_7242);
nor U8111 (N_8111,N_6549,N_7417);
and U8112 (N_8112,N_5626,N_5315);
nor U8113 (N_8113,N_6246,N_7145);
and U8114 (N_8114,N_6377,N_5098);
nor U8115 (N_8115,N_6782,N_5017);
xor U8116 (N_8116,N_6090,N_7397);
nor U8117 (N_8117,N_5882,N_6375);
or U8118 (N_8118,N_6461,N_6031);
nor U8119 (N_8119,N_6553,N_6272);
nor U8120 (N_8120,N_5538,N_5159);
nor U8121 (N_8121,N_7205,N_6957);
or U8122 (N_8122,N_7459,N_6518);
xor U8123 (N_8123,N_5657,N_5978);
nand U8124 (N_8124,N_5712,N_7227);
and U8125 (N_8125,N_6121,N_6503);
xor U8126 (N_8126,N_5757,N_6926);
or U8127 (N_8127,N_6681,N_6573);
or U8128 (N_8128,N_5316,N_6755);
or U8129 (N_8129,N_5065,N_5190);
nand U8130 (N_8130,N_5362,N_5922);
nor U8131 (N_8131,N_6529,N_7186);
and U8132 (N_8132,N_7328,N_7461);
and U8133 (N_8133,N_7252,N_6837);
xor U8134 (N_8134,N_5969,N_6488);
nor U8135 (N_8135,N_7406,N_5453);
nand U8136 (N_8136,N_6977,N_6444);
and U8137 (N_8137,N_5469,N_6464);
and U8138 (N_8138,N_7287,N_5084);
nand U8139 (N_8139,N_6110,N_6083);
or U8140 (N_8140,N_7029,N_7445);
nor U8141 (N_8141,N_5851,N_5731);
xnor U8142 (N_8142,N_7122,N_6180);
xor U8143 (N_8143,N_7302,N_6976);
nand U8144 (N_8144,N_6205,N_5667);
nor U8145 (N_8145,N_5914,N_5764);
or U8146 (N_8146,N_7473,N_5540);
or U8147 (N_8147,N_5658,N_7263);
nand U8148 (N_8148,N_6130,N_6903);
nor U8149 (N_8149,N_6801,N_5740);
or U8150 (N_8150,N_5752,N_6911);
xnor U8151 (N_8151,N_5302,N_7418);
nand U8152 (N_8152,N_7073,N_6397);
and U8153 (N_8153,N_7161,N_6970);
nand U8154 (N_8154,N_6308,N_6369);
xnor U8155 (N_8155,N_5524,N_6625);
nand U8156 (N_8156,N_6682,N_6470);
and U8157 (N_8157,N_6357,N_7048);
or U8158 (N_8158,N_5718,N_6383);
and U8159 (N_8159,N_5997,N_7040);
nand U8160 (N_8160,N_7065,N_6283);
nand U8161 (N_8161,N_7399,N_7077);
nand U8162 (N_8162,N_7103,N_6150);
and U8163 (N_8163,N_5075,N_5801);
and U8164 (N_8164,N_5184,N_7237);
xor U8165 (N_8165,N_6993,N_7112);
xor U8166 (N_8166,N_5146,N_5668);
xnor U8167 (N_8167,N_5523,N_6910);
nor U8168 (N_8168,N_7336,N_6061);
xnor U8169 (N_8169,N_7218,N_7124);
nand U8170 (N_8170,N_6804,N_5735);
and U8171 (N_8171,N_5243,N_5140);
nand U8172 (N_8172,N_7014,N_5638);
nand U8173 (N_8173,N_6504,N_6765);
nand U8174 (N_8174,N_7438,N_6602);
xor U8175 (N_8175,N_5704,N_7269);
and U8176 (N_8176,N_5442,N_5941);
xnor U8177 (N_8177,N_7425,N_5529);
nor U8178 (N_8178,N_6523,N_5779);
nor U8179 (N_8179,N_6995,N_6564);
and U8180 (N_8180,N_6580,N_5711);
or U8181 (N_8181,N_7132,N_7125);
nand U8182 (N_8182,N_6567,N_7379);
nand U8183 (N_8183,N_5793,N_6679);
nand U8184 (N_8184,N_7082,N_6089);
nor U8185 (N_8185,N_6351,N_5139);
and U8186 (N_8186,N_6716,N_5745);
and U8187 (N_8187,N_6595,N_6572);
nor U8188 (N_8188,N_5676,N_6571);
nor U8189 (N_8189,N_7443,N_5935);
and U8190 (N_8190,N_6649,N_5863);
nor U8191 (N_8191,N_6836,N_6822);
and U8192 (N_8192,N_5671,N_5207);
nand U8193 (N_8193,N_5785,N_5784);
nor U8194 (N_8194,N_6560,N_5220);
xnor U8195 (N_8195,N_7436,N_6767);
xor U8196 (N_8196,N_5652,N_7206);
or U8197 (N_8197,N_5858,N_5061);
nand U8198 (N_8198,N_5389,N_6563);
nand U8199 (N_8199,N_5114,N_6229);
or U8200 (N_8200,N_6454,N_6451);
and U8201 (N_8201,N_5276,N_5661);
nor U8202 (N_8202,N_6712,N_7449);
xnor U8203 (N_8203,N_6336,N_6638);
and U8204 (N_8204,N_6044,N_7081);
and U8205 (N_8205,N_6112,N_6719);
nor U8206 (N_8206,N_5871,N_6991);
nor U8207 (N_8207,N_6208,N_6479);
and U8208 (N_8208,N_5059,N_7229);
and U8209 (N_8209,N_5870,N_6378);
nand U8210 (N_8210,N_7413,N_5602);
xnor U8211 (N_8211,N_5024,N_6220);
or U8212 (N_8212,N_7396,N_6676);
or U8213 (N_8213,N_5970,N_7476);
or U8214 (N_8214,N_7113,N_5009);
or U8215 (N_8215,N_5304,N_5078);
nor U8216 (N_8216,N_7481,N_5813);
nand U8217 (N_8217,N_5349,N_7303);
nor U8218 (N_8218,N_6790,N_6390);
nor U8219 (N_8219,N_5955,N_5049);
xnor U8220 (N_8220,N_6939,N_6226);
or U8221 (N_8221,N_5828,N_6122);
nor U8222 (N_8222,N_5818,N_7210);
and U8223 (N_8223,N_7260,N_5202);
nor U8224 (N_8224,N_6772,N_5884);
xnor U8225 (N_8225,N_5430,N_6020);
nand U8226 (N_8226,N_5891,N_5574);
nand U8227 (N_8227,N_7107,N_5519);
or U8228 (N_8228,N_6363,N_5691);
or U8229 (N_8229,N_5633,N_6091);
or U8230 (N_8230,N_5404,N_7248);
and U8231 (N_8231,N_6543,N_6879);
or U8232 (N_8232,N_5410,N_5660);
and U8233 (N_8233,N_5604,N_5596);
xor U8234 (N_8234,N_6817,N_6104);
and U8235 (N_8235,N_7007,N_5621);
xnor U8236 (N_8236,N_5912,N_5809);
or U8237 (N_8237,N_5728,N_6477);
nor U8238 (N_8238,N_6222,N_5041);
or U8239 (N_8239,N_6191,N_7158);
nand U8240 (N_8240,N_5647,N_7434);
or U8241 (N_8241,N_5543,N_7492);
or U8242 (N_8242,N_5775,N_5751);
nand U8243 (N_8243,N_6669,N_7088);
xnor U8244 (N_8244,N_7283,N_6333);
or U8245 (N_8245,N_6930,N_5103);
nand U8246 (N_8246,N_5110,N_5599);
nor U8247 (N_8247,N_6655,N_7070);
and U8248 (N_8248,N_6291,N_5503);
nor U8249 (N_8249,N_7127,N_7171);
and U8250 (N_8250,N_5312,N_7053);
nand U8251 (N_8251,N_6883,N_6160);
nand U8252 (N_8252,N_6832,N_6521);
xor U8253 (N_8253,N_6049,N_6531);
xnor U8254 (N_8254,N_6492,N_5363);
nor U8255 (N_8255,N_6047,N_6027);
xnor U8256 (N_8256,N_5036,N_6603);
nand U8257 (N_8257,N_6004,N_5962);
or U8258 (N_8258,N_5528,N_6992);
or U8259 (N_8259,N_7155,N_5422);
and U8260 (N_8260,N_6389,N_7256);
nor U8261 (N_8261,N_6776,N_6786);
or U8262 (N_8262,N_5079,N_5293);
nand U8263 (N_8263,N_6684,N_5439);
and U8264 (N_8264,N_5993,N_7366);
and U8265 (N_8265,N_5694,N_5864);
nor U8266 (N_8266,N_5305,N_5913);
or U8267 (N_8267,N_6177,N_5381);
xor U8268 (N_8268,N_6084,N_5948);
and U8269 (N_8269,N_6171,N_7211);
nor U8270 (N_8270,N_6668,N_6448);
xor U8271 (N_8271,N_5468,N_6125);
nand U8272 (N_8272,N_7368,N_7376);
xnor U8273 (N_8273,N_7402,N_5952);
nor U8274 (N_8274,N_6380,N_5812);
nor U8275 (N_8275,N_5321,N_5701);
nor U8276 (N_8276,N_5563,N_5938);
and U8277 (N_8277,N_6644,N_7162);
nand U8278 (N_8278,N_7266,N_7120);
nor U8279 (N_8279,N_6231,N_6178);
and U8280 (N_8280,N_5663,N_6760);
xnor U8281 (N_8281,N_6660,N_6546);
or U8282 (N_8282,N_6000,N_6646);
xor U8283 (N_8283,N_5205,N_6919);
nand U8284 (N_8284,N_5215,N_6974);
nand U8285 (N_8285,N_5115,N_5582);
xor U8286 (N_8286,N_5570,N_6373);
and U8287 (N_8287,N_6009,N_5508);
nor U8288 (N_8288,N_7257,N_6640);
xor U8289 (N_8289,N_6753,N_6946);
nor U8290 (N_8290,N_6526,N_7072);
and U8291 (N_8291,N_5402,N_5192);
xnor U8292 (N_8292,N_5736,N_5414);
or U8293 (N_8293,N_6073,N_5185);
or U8294 (N_8294,N_5803,N_5355);
xnor U8295 (N_8295,N_5274,N_7114);
nor U8296 (N_8296,N_5656,N_5832);
and U8297 (N_8297,N_7280,N_6202);
xor U8298 (N_8298,N_6958,N_7432);
and U8299 (N_8299,N_6846,N_6975);
xor U8300 (N_8300,N_5270,N_6829);
nor U8301 (N_8301,N_6932,N_5999);
and U8302 (N_8302,N_7202,N_6688);
or U8303 (N_8303,N_6142,N_5085);
xor U8304 (N_8304,N_7090,N_5797);
nor U8305 (N_8305,N_5301,N_5872);
nand U8306 (N_8306,N_6610,N_6674);
xor U8307 (N_8307,N_6747,N_6823);
or U8308 (N_8308,N_6744,N_7347);
nand U8309 (N_8309,N_5451,N_6558);
and U8310 (N_8310,N_6437,N_6896);
nor U8311 (N_8311,N_7312,N_5208);
and U8312 (N_8312,N_6870,N_5107);
nor U8313 (N_8313,N_5587,N_6455);
or U8314 (N_8314,N_5171,N_6588);
xnor U8315 (N_8315,N_7086,N_7079);
nor U8316 (N_8316,N_7200,N_5890);
nor U8317 (N_8317,N_5194,N_5759);
and U8318 (N_8318,N_6358,N_5269);
nor U8319 (N_8319,N_5081,N_6770);
nand U8320 (N_8320,N_6399,N_5734);
nor U8321 (N_8321,N_5760,N_5908);
and U8322 (N_8322,N_6314,N_5415);
xnor U8323 (N_8323,N_5686,N_6740);
nand U8324 (N_8324,N_6885,N_6973);
and U8325 (N_8325,N_5781,N_7448);
nand U8326 (N_8326,N_6275,N_6392);
nor U8327 (N_8327,N_6309,N_6301);
and U8328 (N_8328,N_6128,N_5311);
nor U8329 (N_8329,N_7386,N_7318);
nor U8330 (N_8330,N_6630,N_5924);
or U8331 (N_8331,N_6774,N_6548);
and U8332 (N_8332,N_7035,N_7299);
nor U8333 (N_8333,N_5794,N_5259);
nor U8334 (N_8334,N_5145,N_6505);
xnor U8335 (N_8335,N_6029,N_6341);
and U8336 (N_8336,N_6577,N_6844);
nor U8337 (N_8337,N_5892,N_5614);
or U8338 (N_8338,N_6217,N_5179);
and U8339 (N_8339,N_5068,N_5898);
nand U8340 (N_8340,N_5973,N_5670);
nand U8341 (N_8341,N_6285,N_6257);
nor U8342 (N_8342,N_7174,N_5598);
nand U8343 (N_8343,N_5799,N_6187);
nand U8344 (N_8344,N_7467,N_5447);
nand U8345 (N_8345,N_7197,N_5187);
and U8346 (N_8346,N_7153,N_5164);
xnor U8347 (N_8347,N_5844,N_6892);
xor U8348 (N_8348,N_5020,N_6079);
and U8349 (N_8349,N_6070,N_7087);
and U8350 (N_8350,N_7381,N_6238);
nand U8351 (N_8351,N_7109,N_7159);
and U8352 (N_8352,N_5498,N_6941);
nor U8353 (N_8353,N_5806,N_5514);
or U8354 (N_8354,N_5463,N_5069);
or U8355 (N_8355,N_5606,N_5385);
or U8356 (N_8356,N_6386,N_7331);
xor U8357 (N_8357,N_6811,N_5130);
or U8358 (N_8358,N_5493,N_7101);
nand U8359 (N_8359,N_5931,N_6008);
nand U8360 (N_8360,N_7078,N_6415);
xor U8361 (N_8361,N_5639,N_6206);
and U8362 (N_8362,N_5425,N_6831);
xnor U8363 (N_8363,N_7056,N_6830);
nand U8364 (N_8364,N_7437,N_6840);
nand U8365 (N_8365,N_6615,N_7364);
nor U8366 (N_8366,N_7447,N_5907);
xor U8367 (N_8367,N_5109,N_6417);
xnor U8368 (N_8368,N_5212,N_5371);
and U8369 (N_8369,N_5765,N_6612);
and U8370 (N_8370,N_5965,N_6276);
nand U8371 (N_8371,N_6462,N_6267);
xor U8372 (N_8372,N_5521,N_5413);
xor U8373 (N_8373,N_6324,N_6214);
and U8374 (N_8374,N_5788,N_6247);
and U8375 (N_8375,N_5725,N_7096);
nand U8376 (N_8376,N_7118,N_7460);
or U8377 (N_8377,N_7389,N_5186);
nor U8378 (N_8378,N_5868,N_5370);
xnor U8379 (N_8379,N_5906,N_5359);
nand U8380 (N_8380,N_5224,N_6149);
and U8381 (N_8381,N_6582,N_5982);
xor U8382 (N_8382,N_7334,N_6921);
nand U8383 (N_8383,N_5236,N_6475);
nor U8384 (N_8384,N_5124,N_6699);
and U8385 (N_8385,N_5013,N_5491);
and U8386 (N_8386,N_7106,N_5454);
or U8387 (N_8387,N_6273,N_6834);
and U8388 (N_8388,N_6144,N_5677);
and U8389 (N_8389,N_6223,N_6136);
or U8390 (N_8390,N_5050,N_5852);
xor U8391 (N_8391,N_5893,N_7224);
nor U8392 (N_8392,N_6435,N_7241);
or U8393 (N_8393,N_6687,N_6727);
xor U8394 (N_8394,N_6347,N_6116);
nor U8395 (N_8395,N_6758,N_6756);
and U8396 (N_8396,N_6718,N_5244);
xor U8397 (N_8397,N_6704,N_5306);
nor U8398 (N_8398,N_7306,N_5354);
nand U8399 (N_8399,N_6796,N_7135);
nand U8400 (N_8400,N_6037,N_5351);
nor U8401 (N_8401,N_6148,N_6528);
or U8402 (N_8402,N_5479,N_6013);
nand U8403 (N_8403,N_7358,N_6597);
xor U8404 (N_8404,N_6183,N_6179);
xnor U8405 (N_8405,N_5557,N_5396);
or U8406 (N_8406,N_6346,N_7333);
nand U8407 (N_8407,N_5603,N_6750);
or U8408 (N_8408,N_6535,N_6645);
or U8409 (N_8409,N_5816,N_7219);
nand U8410 (N_8410,N_6452,N_6282);
or U8411 (N_8411,N_6096,N_6637);
or U8412 (N_8412,N_6001,N_5204);
nor U8413 (N_8413,N_6028,N_5367);
and U8414 (N_8414,N_6902,N_7223);
and U8415 (N_8415,N_6519,N_5166);
or U8416 (N_8416,N_5296,N_5580);
xor U8417 (N_8417,N_5476,N_7270);
or U8418 (N_8418,N_7387,N_7037);
and U8419 (N_8419,N_5125,N_6443);
nand U8420 (N_8420,N_5972,N_6511);
xor U8421 (N_8421,N_7410,N_5790);
nand U8422 (N_8422,N_5456,N_5510);
nor U8423 (N_8423,N_7327,N_5774);
nand U8424 (N_8424,N_5998,N_5201);
nor U8425 (N_8425,N_7245,N_5242);
or U8426 (N_8426,N_6860,N_5465);
nand U8427 (N_8427,N_6596,N_5778);
nor U8428 (N_8428,N_6601,N_6143);
xor U8429 (N_8429,N_7069,N_6607);
xor U8430 (N_8430,N_6617,N_5611);
or U8431 (N_8431,N_6172,N_5292);
nor U8432 (N_8432,N_5380,N_6710);
xor U8433 (N_8433,N_5601,N_5527);
nor U8434 (N_8434,N_5591,N_7018);
or U8435 (N_8435,N_6262,N_7010);
nor U8436 (N_8436,N_6099,N_6978);
nor U8437 (N_8437,N_7128,N_5406);
xnor U8438 (N_8438,N_6372,N_6210);
or U8439 (N_8439,N_6362,N_5520);
xnor U8440 (N_8440,N_5474,N_5289);
nand U8441 (N_8441,N_5129,N_6161);
nor U8442 (N_8442,N_6159,N_5810);
nor U8443 (N_8443,N_7276,N_6395);
and U8444 (N_8444,N_5376,N_6117);
xnor U8445 (N_8445,N_5303,N_7133);
nand U8446 (N_8446,N_6305,N_6465);
nand U8447 (N_8447,N_7352,N_5254);
xor U8448 (N_8448,N_5435,N_6988);
or U8449 (N_8449,N_6942,N_7295);
nor U8450 (N_8450,N_5698,N_7144);
or U8451 (N_8451,N_7351,N_5854);
xnor U8452 (N_8452,N_5641,N_6618);
nand U8453 (N_8453,N_5071,N_6913);
or U8454 (N_8454,N_5143,N_6593);
nand U8455 (N_8455,N_7047,N_7094);
xnor U8456 (N_8456,N_6534,N_6405);
nor U8457 (N_8457,N_5994,N_7184);
and U8458 (N_8458,N_5384,N_5401);
xnor U8459 (N_8459,N_6427,N_6579);
or U8460 (N_8460,N_6898,N_6483);
or U8461 (N_8461,N_7192,N_6990);
or U8462 (N_8462,N_5739,N_6542);
nor U8463 (N_8463,N_5754,N_6706);
xnor U8464 (N_8464,N_5689,N_6799);
and U8465 (N_8465,N_6354,N_6677);
xnor U8466 (N_8466,N_7235,N_7067);
and U8467 (N_8467,N_6585,N_5108);
xnor U8468 (N_8468,N_6915,N_6525);
or U8469 (N_8469,N_7091,N_5196);
or U8470 (N_8470,N_5374,N_6656);
nor U8471 (N_8471,N_5285,N_6951);
or U8472 (N_8472,N_6745,N_5153);
nor U8473 (N_8473,N_5505,N_6241);
and U8474 (N_8474,N_6424,N_7157);
nand U8475 (N_8475,N_6127,N_6778);
or U8476 (N_8476,N_5821,N_7254);
and U8477 (N_8477,N_6243,N_5327);
or U8478 (N_8478,N_6054,N_7404);
or U8479 (N_8479,N_5390,N_6022);
or U8480 (N_8480,N_6647,N_5896);
or U8481 (N_8481,N_5954,N_6265);
or U8482 (N_8482,N_6862,N_6430);
nor U8483 (N_8483,N_5176,N_6408);
or U8484 (N_8484,N_6880,N_6773);
xnor U8485 (N_8485,N_6289,N_5880);
nor U8486 (N_8486,N_6675,N_7282);
or U8487 (N_8487,N_6696,N_5228);
xnor U8488 (N_8488,N_6290,N_5246);
nand U8489 (N_8489,N_5092,N_6841);
or U8490 (N_8490,N_7080,N_5615);
nand U8491 (N_8491,N_6833,N_7499);
or U8492 (N_8492,N_6562,N_5971);
nor U8493 (N_8493,N_7034,N_7142);
and U8494 (N_8494,N_5690,N_7465);
and U8495 (N_8495,N_7478,N_5210);
xnor U8496 (N_8496,N_6516,N_5464);
and U8497 (N_8497,N_7297,N_6732);
and U8498 (N_8498,N_5308,N_6350);
nor U8499 (N_8499,N_6436,N_5264);
or U8500 (N_8500,N_7054,N_6793);
nand U8501 (N_8501,N_7392,N_5206);
nor U8502 (N_8502,N_5593,N_7486);
nand U8503 (N_8503,N_5387,N_7022);
nand U8504 (N_8504,N_6230,N_6807);
nand U8505 (N_8505,N_5466,N_6007);
and U8506 (N_8506,N_7163,N_6865);
and U8507 (N_8507,N_6713,N_5112);
nand U8508 (N_8508,N_7463,N_5209);
nor U8509 (N_8509,N_6113,N_5398);
nand U8510 (N_8510,N_7279,N_7134);
nand U8511 (N_8511,N_5544,N_5393);
and U8512 (N_8512,N_6328,N_5839);
nor U8513 (N_8513,N_6551,N_6052);
or U8514 (N_8514,N_5820,N_6145);
nor U8515 (N_8515,N_5840,N_7384);
nor U8516 (N_8516,N_5070,N_5250);
or U8517 (N_8517,N_5551,N_5300);
nand U8518 (N_8518,N_5627,N_6162);
and U8519 (N_8519,N_7294,N_6359);
and U8520 (N_8520,N_7021,N_7233);
nand U8521 (N_8521,N_6555,N_6608);
or U8522 (N_8522,N_6287,N_6318);
xor U8523 (N_8523,N_6653,N_6781);
and U8524 (N_8524,N_5119,N_6033);
nor U8525 (N_8525,N_5707,N_7234);
nand U8526 (N_8526,N_5281,N_5823);
xnor U8527 (N_8527,N_6002,N_5763);
nor U8528 (N_8528,N_7177,N_5484);
and U8529 (N_8529,N_6925,N_7308);
or U8530 (N_8530,N_5142,N_6851);
nand U8531 (N_8531,N_6106,N_6371);
xnor U8532 (N_8532,N_7002,N_5866);
or U8533 (N_8533,N_7296,N_6507);
nor U8534 (N_8534,N_7412,N_5284);
or U8535 (N_8535,N_6356,N_5035);
nand U8536 (N_8536,N_6721,N_6967);
and U8537 (N_8537,N_5838,N_6306);
or U8538 (N_8538,N_7450,N_6576);
nor U8539 (N_8539,N_6559,N_6702);
or U8540 (N_8540,N_5980,N_6219);
or U8541 (N_8541,N_6806,N_7115);
and U8542 (N_8542,N_6775,N_5094);
and U8543 (N_8543,N_6547,N_6701);
nor U8544 (N_8544,N_6280,N_5696);
or U8545 (N_8545,N_6724,N_5934);
and U8546 (N_8546,N_7012,N_6996);
and U8547 (N_8547,N_6673,N_7165);
xor U8548 (N_8548,N_6334,N_7196);
or U8549 (N_8549,N_7471,N_6889);
xor U8550 (N_8550,N_6413,N_6907);
or U8551 (N_8551,N_6019,N_6441);
nor U8552 (N_8552,N_5135,N_5271);
nand U8553 (N_8553,N_6768,N_6109);
nor U8554 (N_8554,N_5534,N_5245);
xnor U8555 (N_8555,N_5847,N_6741);
nand U8556 (N_8556,N_5322,N_7217);
and U8557 (N_8557,N_6838,N_5230);
xnor U8558 (N_8558,N_6277,N_6239);
xnor U8559 (N_8559,N_5000,N_5155);
and U8560 (N_8560,N_5946,N_5470);
or U8561 (N_8561,N_6322,N_6218);
xnor U8562 (N_8562,N_6742,N_7329);
nand U8563 (N_8563,N_6876,N_5648);
and U8564 (N_8564,N_5710,N_6134);
or U8565 (N_8565,N_6337,N_6616);
and U8566 (N_8566,N_7141,N_6409);
or U8567 (N_8567,N_7470,N_6641);
xor U8568 (N_8568,N_6614,N_5750);
xor U8569 (N_8569,N_5678,N_5030);
nand U8570 (N_8570,N_6081,N_5594);
and U8571 (N_8571,N_6453,N_6485);
nor U8572 (N_8572,N_6869,N_6126);
and U8573 (N_8573,N_6299,N_5032);
nand U8574 (N_8574,N_7453,N_6809);
nor U8575 (N_8575,N_6332,N_6192);
or U8576 (N_8576,N_5697,N_6017);
and U8577 (N_8577,N_7044,N_7017);
nand U8578 (N_8578,N_5630,N_6850);
xor U8579 (N_8579,N_6414,N_5473);
nand U8580 (N_8580,N_5634,N_5358);
nand U8581 (N_8581,N_5687,N_7150);
nand U8582 (N_8582,N_5436,N_5416);
nand U8583 (N_8583,N_5160,N_6680);
or U8584 (N_8584,N_7483,N_6074);
or U8585 (N_8585,N_6947,N_6480);
or U8586 (N_8586,N_5045,N_6115);
or U8587 (N_8587,N_7116,N_5375);
nor U8588 (N_8588,N_7310,N_6857);
nor U8589 (N_8589,N_5136,N_7100);
or U8590 (N_8590,N_6735,N_7179);
or U8591 (N_8591,N_5929,N_6861);
nand U8592 (N_8592,N_6169,N_7420);
nor U8593 (N_8593,N_7493,N_5216);
nor U8594 (N_8594,N_6188,N_5093);
xor U8595 (N_8595,N_5719,N_6754);
or U8596 (N_8596,N_5692,N_6327);
and U8597 (N_8597,N_5753,N_6848);
xor U8598 (N_8598,N_5876,N_7435);
or U8599 (N_8599,N_7061,N_7129);
nor U8600 (N_8600,N_7464,N_7313);
and U8601 (N_8601,N_6763,N_6194);
nand U8602 (N_8602,N_6153,N_6629);
nor U8603 (N_8603,N_6457,N_6382);
or U8604 (N_8604,N_5800,N_5175);
nand U8605 (N_8605,N_5058,N_6805);
and U8606 (N_8606,N_6173,N_5077);
xor U8607 (N_8607,N_5617,N_7209);
nor U8608 (N_8608,N_6969,N_5780);
nor U8609 (N_8609,N_5334,N_5287);
or U8610 (N_8610,N_5805,N_5945);
nor U8611 (N_8611,N_5063,N_6854);
and U8612 (N_8612,N_5237,N_5837);
nor U8613 (N_8613,N_5022,N_5462);
or U8614 (N_8614,N_7289,N_6497);
xor U8615 (N_8615,N_5432,N_5983);
nand U8616 (N_8616,N_6536,N_6502);
nor U8617 (N_8617,N_6093,N_5343);
nor U8618 (N_8618,N_6591,N_5612);
nand U8619 (N_8619,N_7176,N_7265);
xor U8620 (N_8620,N_5283,N_7362);
nor U8621 (N_8621,N_5386,N_6138);
xnor U8622 (N_8622,N_6565,N_5568);
or U8623 (N_8623,N_6286,N_5291);
or U8624 (N_8624,N_5290,N_5123);
xnor U8625 (N_8625,N_7111,N_6119);
xor U8626 (N_8626,N_6374,N_6592);
or U8627 (N_8627,N_6271,N_6761);
nand U8628 (N_8628,N_5546,N_6604);
nand U8629 (N_8629,N_6181,N_5042);
or U8630 (N_8630,N_6839,N_6055);
xor U8631 (N_8631,N_6036,N_6251);
nand U8632 (N_8632,N_6215,N_7204);
nor U8633 (N_8633,N_6094,N_5280);
or U8634 (N_8634,N_5424,N_5105);
nand U8635 (N_8635,N_6672,N_7316);
xor U8636 (N_8636,N_5234,N_5169);
or U8637 (N_8637,N_6490,N_6725);
nand U8638 (N_8638,N_6394,N_5749);
or U8639 (N_8639,N_5189,N_7339);
or U8640 (N_8640,N_7225,N_6624);
and U8641 (N_8641,N_7154,N_5635);
nand U8642 (N_8642,N_5288,N_6189);
and U8643 (N_8643,N_5533,N_6224);
or U8644 (N_8644,N_7489,N_5340);
xnor U8645 (N_8645,N_5985,N_5144);
and U8646 (N_8646,N_6041,N_7249);
and U8647 (N_8647,N_5323,N_6137);
or U8648 (N_8648,N_6652,N_5421);
and U8649 (N_8649,N_5916,N_6648);
nor U8650 (N_8650,N_6426,N_7255);
and U8651 (N_8651,N_5894,N_6132);
nand U8652 (N_8652,N_7084,N_5382);
nor U8653 (N_8653,N_5758,N_6859);
and U8654 (N_8654,N_6011,N_5950);
nand U8655 (N_8655,N_5309,N_5088);
and U8656 (N_8656,N_5987,N_7323);
nand U8657 (N_8657,N_5446,N_5651);
or U8658 (N_8658,N_6063,N_7004);
nor U8659 (N_8659,N_5808,N_7353);
nor U8660 (N_8660,N_7138,N_5333);
nand U8661 (N_8661,N_6376,N_6950);
xor U8662 (N_8662,N_5497,N_7301);
and U8663 (N_8663,N_6233,N_6472);
nor U8664 (N_8664,N_7147,N_6123);
or U8665 (N_8665,N_6904,N_5675);
xnor U8666 (N_8666,N_5607,N_7026);
nor U8667 (N_8667,N_6168,N_6087);
and U8668 (N_8668,N_5213,N_6196);
and U8669 (N_8669,N_7375,N_5033);
nor U8670 (N_8670,N_7036,N_7213);
xnor U8671 (N_8671,N_5613,N_5038);
nor U8672 (N_8672,N_6486,N_6107);
nor U8673 (N_8673,N_6784,N_6078);
nor U8674 (N_8674,N_6422,N_5877);
nor U8675 (N_8675,N_6933,N_5909);
xor U8676 (N_8676,N_7136,N_6800);
xor U8677 (N_8677,N_5554,N_5313);
nand U8678 (N_8678,N_5860,N_6963);
nand U8679 (N_8679,N_5722,N_6476);
xnor U8680 (N_8680,N_7108,N_5513);
nand U8681 (N_8681,N_7377,N_5418);
and U8682 (N_8682,N_5486,N_5154);
and U8683 (N_8683,N_5227,N_7187);
nand U8684 (N_8684,N_6792,N_6264);
and U8685 (N_8685,N_5014,N_6627);
nand U8686 (N_8686,N_7442,N_6759);
or U8687 (N_8687,N_7278,N_5445);
nor U8688 (N_8688,N_6312,N_7104);
and U8689 (N_8689,N_5984,N_5850);
or U8690 (N_8690,N_5299,N_6814);
xnor U8691 (N_8691,N_6296,N_5392);
and U8692 (N_8692,N_5117,N_5653);
nand U8693 (N_8693,N_6151,N_7469);
nand U8694 (N_8694,N_7038,N_6494);
or U8695 (N_8695,N_6557,N_5044);
and U8696 (N_8696,N_5437,N_7439);
and U8697 (N_8697,N_5713,N_6379);
nand U8698 (N_8698,N_6757,N_5649);
and U8699 (N_8699,N_7098,N_7207);
or U8700 (N_8700,N_7074,N_5158);
and U8701 (N_8701,N_7102,N_6791);
nor U8702 (N_8702,N_5222,N_7253);
xor U8703 (N_8703,N_6927,N_5904);
or U8704 (N_8704,N_5721,N_6513);
xnor U8705 (N_8705,N_7342,N_5218);
nand U8706 (N_8706,N_7024,N_6766);
xnor U8707 (N_8707,N_5487,N_6467);
or U8708 (N_8708,N_6495,N_5817);
nor U8709 (N_8709,N_5536,N_7185);
nand U8710 (N_8710,N_6352,N_5666);
nand U8711 (N_8711,N_6901,N_6897);
xnor U8712 (N_8712,N_6894,N_7261);
xnor U8713 (N_8713,N_5843,N_6101);
xnor U8714 (N_8714,N_6700,N_6953);
nor U8715 (N_8715,N_6733,N_5673);
nor U8716 (N_8716,N_6736,N_6657);
nand U8717 (N_8717,N_5716,N_5132);
xnor U8718 (N_8718,N_7178,N_7304);
or U8719 (N_8719,N_5052,N_5609);
or U8720 (N_8720,N_6891,N_7066);
and U8721 (N_8721,N_5548,N_5181);
xnor U8722 (N_8722,N_5133,N_6156);
xor U8723 (N_8723,N_5475,N_6077);
xor U8724 (N_8724,N_5619,N_7139);
nand U8725 (N_8725,N_6569,N_6064);
xnor U8726 (N_8726,N_5100,N_6643);
or U8727 (N_8727,N_5584,N_6361);
or U8728 (N_8728,N_6447,N_5448);
and U8729 (N_8729,N_7441,N_6496);
nor U8730 (N_8730,N_6720,N_6785);
nand U8731 (N_8731,N_6874,N_5091);
or U8732 (N_8732,N_5096,N_7168);
or U8733 (N_8733,N_6018,N_5217);
nor U8734 (N_8734,N_5961,N_6965);
and U8735 (N_8735,N_5490,N_5878);
or U8736 (N_8736,N_7143,N_5427);
xor U8737 (N_8737,N_6599,N_5887);
xor U8738 (N_8738,N_6199,N_6343);
and U8739 (N_8739,N_5173,N_7166);
nor U8740 (N_8740,N_5174,N_5325);
xnor U8741 (N_8741,N_6043,N_6487);
nand U8742 (N_8742,N_7433,N_5855);
nand U8743 (N_8743,N_5161,N_6349);
nand U8744 (N_8744,N_5026,N_6802);
nor U8745 (N_8745,N_5881,N_6069);
nand U8746 (N_8746,N_7457,N_6252);
xor U8747 (N_8747,N_5450,N_6431);
nor U8748 (N_8748,N_5277,N_7343);
and U8749 (N_8749,N_6633,N_5836);
and U8750 (N_8750,N_6882,N_6590);
or U8751 (N_8751,N_5240,N_5023);
or U8752 (N_8752,N_7082,N_7166);
nor U8753 (N_8753,N_6383,N_6999);
or U8754 (N_8754,N_7382,N_5412);
nand U8755 (N_8755,N_6896,N_5029);
and U8756 (N_8756,N_6131,N_5405);
nor U8757 (N_8757,N_7429,N_6811);
or U8758 (N_8758,N_6642,N_6568);
or U8759 (N_8759,N_5068,N_6144);
xor U8760 (N_8760,N_5858,N_5479);
nor U8761 (N_8761,N_6897,N_7210);
nor U8762 (N_8762,N_6008,N_5118);
nand U8763 (N_8763,N_6631,N_6651);
and U8764 (N_8764,N_6416,N_5015);
nor U8765 (N_8765,N_5099,N_6280);
xor U8766 (N_8766,N_6980,N_5915);
or U8767 (N_8767,N_7314,N_7404);
or U8768 (N_8768,N_6264,N_6355);
and U8769 (N_8769,N_6755,N_7214);
nand U8770 (N_8770,N_7102,N_5492);
nand U8771 (N_8771,N_7450,N_6319);
and U8772 (N_8772,N_6132,N_6803);
nor U8773 (N_8773,N_6932,N_5243);
xor U8774 (N_8774,N_6596,N_6910);
nand U8775 (N_8775,N_5513,N_5452);
or U8776 (N_8776,N_5652,N_5552);
xnor U8777 (N_8777,N_6555,N_7332);
or U8778 (N_8778,N_7140,N_6161);
nand U8779 (N_8779,N_6292,N_5873);
and U8780 (N_8780,N_7100,N_5206);
xnor U8781 (N_8781,N_6433,N_5899);
xnor U8782 (N_8782,N_5454,N_5484);
nand U8783 (N_8783,N_6826,N_7284);
and U8784 (N_8784,N_7414,N_5601);
nor U8785 (N_8785,N_6980,N_5051);
xnor U8786 (N_8786,N_6501,N_7122);
xnor U8787 (N_8787,N_6001,N_7258);
xnor U8788 (N_8788,N_5866,N_7286);
and U8789 (N_8789,N_7456,N_6332);
or U8790 (N_8790,N_6061,N_5889);
or U8791 (N_8791,N_5734,N_7192);
nand U8792 (N_8792,N_5836,N_7319);
nand U8793 (N_8793,N_6373,N_5869);
and U8794 (N_8794,N_6397,N_6033);
xnor U8795 (N_8795,N_7125,N_6700);
or U8796 (N_8796,N_6384,N_5958);
xnor U8797 (N_8797,N_6939,N_5345);
xnor U8798 (N_8798,N_5987,N_5051);
xor U8799 (N_8799,N_6651,N_5016);
xor U8800 (N_8800,N_6887,N_6311);
xnor U8801 (N_8801,N_6248,N_5969);
nor U8802 (N_8802,N_5511,N_5166);
nand U8803 (N_8803,N_7120,N_5840);
and U8804 (N_8804,N_5258,N_6710);
and U8805 (N_8805,N_6775,N_6062);
or U8806 (N_8806,N_7315,N_5638);
or U8807 (N_8807,N_6612,N_5712);
nor U8808 (N_8808,N_5014,N_6569);
nor U8809 (N_8809,N_6533,N_6352);
and U8810 (N_8810,N_5599,N_6447);
or U8811 (N_8811,N_5017,N_7447);
nand U8812 (N_8812,N_6427,N_6465);
xor U8813 (N_8813,N_5628,N_5925);
or U8814 (N_8814,N_6711,N_6341);
xor U8815 (N_8815,N_7404,N_6972);
nand U8816 (N_8816,N_6567,N_5524);
nand U8817 (N_8817,N_5231,N_5240);
and U8818 (N_8818,N_5686,N_5424);
nand U8819 (N_8819,N_6713,N_5886);
nand U8820 (N_8820,N_7011,N_5904);
xnor U8821 (N_8821,N_5623,N_5055);
nand U8822 (N_8822,N_6752,N_5351);
nand U8823 (N_8823,N_5965,N_6115);
xnor U8824 (N_8824,N_6799,N_5112);
or U8825 (N_8825,N_7314,N_5918);
nand U8826 (N_8826,N_6014,N_5759);
and U8827 (N_8827,N_7317,N_6991);
or U8828 (N_8828,N_5469,N_6888);
nand U8829 (N_8829,N_5777,N_5411);
xor U8830 (N_8830,N_6509,N_6163);
nor U8831 (N_8831,N_5024,N_6956);
nor U8832 (N_8832,N_5849,N_6732);
xnor U8833 (N_8833,N_6448,N_5028);
xor U8834 (N_8834,N_5013,N_5521);
xor U8835 (N_8835,N_6429,N_6028);
xnor U8836 (N_8836,N_7190,N_5416);
xor U8837 (N_8837,N_6964,N_5751);
xor U8838 (N_8838,N_5486,N_5254);
and U8839 (N_8839,N_6168,N_5701);
xnor U8840 (N_8840,N_7464,N_6702);
xnor U8841 (N_8841,N_7063,N_7129);
xor U8842 (N_8842,N_6173,N_5889);
and U8843 (N_8843,N_5987,N_5342);
nor U8844 (N_8844,N_6176,N_7209);
or U8845 (N_8845,N_7165,N_6345);
xor U8846 (N_8846,N_5519,N_6495);
and U8847 (N_8847,N_6101,N_5122);
nor U8848 (N_8848,N_7412,N_5227);
or U8849 (N_8849,N_5316,N_6663);
nor U8850 (N_8850,N_6148,N_5942);
xor U8851 (N_8851,N_5161,N_5031);
xor U8852 (N_8852,N_7076,N_6583);
or U8853 (N_8853,N_6671,N_6289);
or U8854 (N_8854,N_6814,N_5508);
nand U8855 (N_8855,N_7414,N_6649);
nand U8856 (N_8856,N_5238,N_5440);
nand U8857 (N_8857,N_5409,N_5160);
or U8858 (N_8858,N_6298,N_6067);
and U8859 (N_8859,N_5469,N_6611);
nor U8860 (N_8860,N_7033,N_7248);
nand U8861 (N_8861,N_6306,N_7071);
or U8862 (N_8862,N_7074,N_6637);
nand U8863 (N_8863,N_6380,N_7208);
nor U8864 (N_8864,N_6109,N_7413);
or U8865 (N_8865,N_5630,N_7433);
nand U8866 (N_8866,N_6001,N_7129);
nor U8867 (N_8867,N_5358,N_5659);
xnor U8868 (N_8868,N_5683,N_5156);
nor U8869 (N_8869,N_6608,N_5265);
nor U8870 (N_8870,N_6636,N_5653);
nor U8871 (N_8871,N_6226,N_6153);
xnor U8872 (N_8872,N_7343,N_6885);
nor U8873 (N_8873,N_6565,N_6166);
nor U8874 (N_8874,N_7464,N_6042);
xnor U8875 (N_8875,N_5310,N_6914);
or U8876 (N_8876,N_5901,N_5318);
xor U8877 (N_8877,N_6853,N_6375);
xnor U8878 (N_8878,N_7167,N_5221);
and U8879 (N_8879,N_5236,N_6519);
nand U8880 (N_8880,N_5525,N_5033);
nand U8881 (N_8881,N_6511,N_5515);
xor U8882 (N_8882,N_5998,N_5855);
and U8883 (N_8883,N_5467,N_5052);
nand U8884 (N_8884,N_6411,N_6884);
nor U8885 (N_8885,N_6429,N_7370);
nor U8886 (N_8886,N_5866,N_5446);
and U8887 (N_8887,N_5701,N_7160);
nand U8888 (N_8888,N_5237,N_5592);
or U8889 (N_8889,N_7231,N_6115);
or U8890 (N_8890,N_5419,N_6831);
and U8891 (N_8891,N_6819,N_6933);
nand U8892 (N_8892,N_5675,N_6286);
nand U8893 (N_8893,N_5668,N_6638);
xor U8894 (N_8894,N_7369,N_6903);
nor U8895 (N_8895,N_7068,N_6413);
nor U8896 (N_8896,N_6962,N_6139);
or U8897 (N_8897,N_5625,N_6503);
nand U8898 (N_8898,N_6489,N_7112);
and U8899 (N_8899,N_6046,N_6468);
xnor U8900 (N_8900,N_5704,N_6509);
xor U8901 (N_8901,N_6418,N_5483);
xor U8902 (N_8902,N_5254,N_7215);
xnor U8903 (N_8903,N_5063,N_6496);
xor U8904 (N_8904,N_7374,N_7186);
nor U8905 (N_8905,N_7218,N_7152);
xnor U8906 (N_8906,N_5213,N_7481);
and U8907 (N_8907,N_7480,N_6715);
xnor U8908 (N_8908,N_5360,N_5073);
or U8909 (N_8909,N_6590,N_6074);
nor U8910 (N_8910,N_7244,N_5470);
nand U8911 (N_8911,N_5388,N_5615);
xor U8912 (N_8912,N_7171,N_5621);
or U8913 (N_8913,N_5303,N_5070);
nor U8914 (N_8914,N_5167,N_5165);
or U8915 (N_8915,N_7183,N_6811);
or U8916 (N_8916,N_7425,N_7257);
nor U8917 (N_8917,N_5451,N_7303);
nand U8918 (N_8918,N_7485,N_6424);
nor U8919 (N_8919,N_6159,N_6381);
and U8920 (N_8920,N_5303,N_6836);
xnor U8921 (N_8921,N_5405,N_5799);
nor U8922 (N_8922,N_6415,N_5313);
or U8923 (N_8923,N_5370,N_6826);
or U8924 (N_8924,N_6134,N_5140);
nor U8925 (N_8925,N_6898,N_5672);
xor U8926 (N_8926,N_5950,N_7406);
nand U8927 (N_8927,N_5460,N_5388);
or U8928 (N_8928,N_6321,N_5463);
xnor U8929 (N_8929,N_6470,N_5093);
nand U8930 (N_8930,N_6969,N_6464);
or U8931 (N_8931,N_7163,N_5483);
and U8932 (N_8932,N_6901,N_6367);
nor U8933 (N_8933,N_6692,N_6177);
xnor U8934 (N_8934,N_7482,N_6969);
xnor U8935 (N_8935,N_5361,N_6351);
nand U8936 (N_8936,N_6364,N_7227);
nor U8937 (N_8937,N_6548,N_7274);
nand U8938 (N_8938,N_5155,N_6206);
or U8939 (N_8939,N_6553,N_6890);
nand U8940 (N_8940,N_6356,N_5172);
or U8941 (N_8941,N_6803,N_7288);
and U8942 (N_8942,N_7247,N_7224);
or U8943 (N_8943,N_5508,N_6089);
and U8944 (N_8944,N_7038,N_5154);
xor U8945 (N_8945,N_5633,N_5569);
and U8946 (N_8946,N_6169,N_6608);
and U8947 (N_8947,N_5803,N_7276);
and U8948 (N_8948,N_6029,N_6891);
or U8949 (N_8949,N_7211,N_6982);
or U8950 (N_8950,N_7031,N_6322);
nand U8951 (N_8951,N_6671,N_6307);
and U8952 (N_8952,N_5355,N_6418);
xnor U8953 (N_8953,N_7406,N_6185);
nor U8954 (N_8954,N_5741,N_5591);
or U8955 (N_8955,N_6239,N_5016);
nor U8956 (N_8956,N_7387,N_7163);
and U8957 (N_8957,N_6378,N_6123);
and U8958 (N_8958,N_5866,N_5123);
nor U8959 (N_8959,N_6982,N_6923);
nand U8960 (N_8960,N_7348,N_6426);
nand U8961 (N_8961,N_7246,N_5320);
nor U8962 (N_8962,N_7445,N_6586);
nand U8963 (N_8963,N_6974,N_5734);
nand U8964 (N_8964,N_5071,N_7319);
and U8965 (N_8965,N_6751,N_6142);
and U8966 (N_8966,N_5341,N_6444);
nor U8967 (N_8967,N_5093,N_5845);
nor U8968 (N_8968,N_6836,N_5348);
or U8969 (N_8969,N_6978,N_6399);
and U8970 (N_8970,N_5623,N_5180);
or U8971 (N_8971,N_7147,N_6080);
nand U8972 (N_8972,N_5799,N_6483);
xnor U8973 (N_8973,N_5707,N_6922);
and U8974 (N_8974,N_6554,N_6096);
xor U8975 (N_8975,N_7499,N_6769);
or U8976 (N_8976,N_5089,N_6810);
xor U8977 (N_8977,N_6813,N_5386);
nor U8978 (N_8978,N_5113,N_6721);
or U8979 (N_8979,N_6717,N_6245);
nor U8980 (N_8980,N_7304,N_7383);
nand U8981 (N_8981,N_6815,N_5752);
xnor U8982 (N_8982,N_5781,N_5408);
xnor U8983 (N_8983,N_6300,N_5259);
and U8984 (N_8984,N_6010,N_6838);
nor U8985 (N_8985,N_6774,N_7279);
and U8986 (N_8986,N_6182,N_5523);
nand U8987 (N_8987,N_5190,N_6973);
nand U8988 (N_8988,N_6426,N_5037);
xnor U8989 (N_8989,N_5988,N_7041);
xor U8990 (N_8990,N_6612,N_5371);
and U8991 (N_8991,N_6487,N_6911);
and U8992 (N_8992,N_7466,N_5904);
and U8993 (N_8993,N_6178,N_6194);
nand U8994 (N_8994,N_6760,N_6028);
and U8995 (N_8995,N_7294,N_6084);
nand U8996 (N_8996,N_5110,N_7149);
and U8997 (N_8997,N_6521,N_7135);
xnor U8998 (N_8998,N_5310,N_5812);
and U8999 (N_8999,N_6304,N_5069);
or U9000 (N_9000,N_6788,N_6901);
nand U9001 (N_9001,N_6949,N_5924);
nand U9002 (N_9002,N_5944,N_6247);
nor U9003 (N_9003,N_5418,N_5266);
or U9004 (N_9004,N_6042,N_7318);
xnor U9005 (N_9005,N_5221,N_5011);
and U9006 (N_9006,N_6952,N_5681);
or U9007 (N_9007,N_5864,N_7327);
or U9008 (N_9008,N_7177,N_6352);
or U9009 (N_9009,N_7480,N_7050);
or U9010 (N_9010,N_6135,N_6710);
nand U9011 (N_9011,N_6536,N_7097);
xor U9012 (N_9012,N_6642,N_7453);
nor U9013 (N_9013,N_6754,N_6814);
nor U9014 (N_9014,N_5599,N_6561);
nand U9015 (N_9015,N_5552,N_5678);
or U9016 (N_9016,N_6178,N_5302);
nand U9017 (N_9017,N_5333,N_7152);
or U9018 (N_9018,N_7450,N_5281);
nor U9019 (N_9019,N_7346,N_7233);
and U9020 (N_9020,N_5789,N_5804);
nand U9021 (N_9021,N_7463,N_5678);
and U9022 (N_9022,N_5189,N_7492);
nand U9023 (N_9023,N_6531,N_5670);
nand U9024 (N_9024,N_6948,N_6413);
or U9025 (N_9025,N_6788,N_6332);
or U9026 (N_9026,N_5447,N_7269);
nand U9027 (N_9027,N_5117,N_5719);
nand U9028 (N_9028,N_5838,N_5536);
xor U9029 (N_9029,N_6132,N_6724);
and U9030 (N_9030,N_5645,N_5696);
xnor U9031 (N_9031,N_7368,N_7070);
or U9032 (N_9032,N_6993,N_6937);
or U9033 (N_9033,N_6199,N_6463);
xnor U9034 (N_9034,N_5493,N_5772);
nand U9035 (N_9035,N_5986,N_5428);
xor U9036 (N_9036,N_6898,N_6444);
and U9037 (N_9037,N_6872,N_5554);
xnor U9038 (N_9038,N_5256,N_5840);
or U9039 (N_9039,N_5972,N_7035);
nor U9040 (N_9040,N_5067,N_7488);
or U9041 (N_9041,N_5396,N_6763);
nor U9042 (N_9042,N_5286,N_6081);
nand U9043 (N_9043,N_6973,N_6475);
nor U9044 (N_9044,N_6366,N_5202);
nand U9045 (N_9045,N_6152,N_7084);
and U9046 (N_9046,N_6385,N_5512);
and U9047 (N_9047,N_7084,N_5465);
or U9048 (N_9048,N_7403,N_6576);
nand U9049 (N_9049,N_6069,N_5828);
nand U9050 (N_9050,N_6289,N_6269);
nor U9051 (N_9051,N_5965,N_7379);
xor U9052 (N_9052,N_6219,N_6768);
nand U9053 (N_9053,N_5253,N_6941);
and U9054 (N_9054,N_5170,N_6467);
xor U9055 (N_9055,N_6308,N_6537);
and U9056 (N_9056,N_5908,N_5987);
xnor U9057 (N_9057,N_6459,N_5707);
xor U9058 (N_9058,N_6067,N_6665);
nor U9059 (N_9059,N_7048,N_6780);
nor U9060 (N_9060,N_5681,N_6125);
nand U9061 (N_9061,N_5629,N_6877);
xnor U9062 (N_9062,N_5613,N_6565);
or U9063 (N_9063,N_5451,N_7493);
nor U9064 (N_9064,N_5089,N_7326);
nor U9065 (N_9065,N_7426,N_6593);
and U9066 (N_9066,N_6058,N_6168);
nor U9067 (N_9067,N_5115,N_6093);
xor U9068 (N_9068,N_6510,N_7424);
and U9069 (N_9069,N_5756,N_6697);
and U9070 (N_9070,N_6511,N_5332);
and U9071 (N_9071,N_7125,N_6010);
nand U9072 (N_9072,N_6826,N_6885);
nand U9073 (N_9073,N_5820,N_5596);
and U9074 (N_9074,N_7358,N_6196);
nand U9075 (N_9075,N_5663,N_5368);
and U9076 (N_9076,N_6949,N_5072);
and U9077 (N_9077,N_7078,N_6430);
and U9078 (N_9078,N_5225,N_7291);
nor U9079 (N_9079,N_5105,N_5220);
nand U9080 (N_9080,N_6047,N_6346);
or U9081 (N_9081,N_5246,N_5434);
nand U9082 (N_9082,N_5104,N_6809);
nand U9083 (N_9083,N_6509,N_7481);
or U9084 (N_9084,N_6831,N_6324);
xnor U9085 (N_9085,N_5163,N_5952);
nand U9086 (N_9086,N_6291,N_7069);
nand U9087 (N_9087,N_5319,N_6780);
or U9088 (N_9088,N_5469,N_6274);
nor U9089 (N_9089,N_7219,N_7239);
xnor U9090 (N_9090,N_7302,N_7310);
nand U9091 (N_9091,N_5488,N_6985);
or U9092 (N_9092,N_5041,N_5209);
and U9093 (N_9093,N_7016,N_6121);
xnor U9094 (N_9094,N_5504,N_5596);
nand U9095 (N_9095,N_7366,N_5095);
nor U9096 (N_9096,N_5368,N_5997);
nor U9097 (N_9097,N_5386,N_5879);
xor U9098 (N_9098,N_5573,N_6621);
nand U9099 (N_9099,N_7084,N_7335);
and U9100 (N_9100,N_6828,N_7124);
nand U9101 (N_9101,N_5268,N_6825);
nor U9102 (N_9102,N_5627,N_7127);
nand U9103 (N_9103,N_6843,N_6800);
nand U9104 (N_9104,N_5349,N_5840);
xor U9105 (N_9105,N_7312,N_5714);
nor U9106 (N_9106,N_5368,N_6613);
and U9107 (N_9107,N_5790,N_6125);
nand U9108 (N_9108,N_7271,N_5387);
or U9109 (N_9109,N_6617,N_5375);
nand U9110 (N_9110,N_6469,N_6242);
xnor U9111 (N_9111,N_6765,N_5177);
nor U9112 (N_9112,N_5201,N_6011);
nor U9113 (N_9113,N_5373,N_5872);
and U9114 (N_9114,N_5329,N_5272);
or U9115 (N_9115,N_5984,N_6961);
and U9116 (N_9116,N_6889,N_6566);
nand U9117 (N_9117,N_5983,N_7033);
nor U9118 (N_9118,N_6197,N_7200);
nand U9119 (N_9119,N_6430,N_5599);
and U9120 (N_9120,N_6418,N_7218);
nand U9121 (N_9121,N_5891,N_5855);
nor U9122 (N_9122,N_5760,N_5470);
or U9123 (N_9123,N_5567,N_6513);
or U9124 (N_9124,N_7121,N_7434);
xnor U9125 (N_9125,N_7037,N_6633);
xor U9126 (N_9126,N_6301,N_7012);
nand U9127 (N_9127,N_6762,N_5067);
xor U9128 (N_9128,N_5062,N_6930);
xor U9129 (N_9129,N_7151,N_6615);
or U9130 (N_9130,N_6677,N_6148);
xnor U9131 (N_9131,N_7196,N_5876);
and U9132 (N_9132,N_5223,N_5573);
nor U9133 (N_9133,N_6520,N_7197);
nand U9134 (N_9134,N_5741,N_7345);
and U9135 (N_9135,N_6557,N_5206);
and U9136 (N_9136,N_6340,N_6528);
nand U9137 (N_9137,N_7269,N_5092);
and U9138 (N_9138,N_5307,N_5067);
and U9139 (N_9139,N_6245,N_6269);
xor U9140 (N_9140,N_6049,N_5250);
and U9141 (N_9141,N_5218,N_5766);
and U9142 (N_9142,N_5579,N_6266);
nor U9143 (N_9143,N_7240,N_5407);
and U9144 (N_9144,N_5536,N_7340);
xnor U9145 (N_9145,N_6592,N_7323);
nand U9146 (N_9146,N_5055,N_6957);
xnor U9147 (N_9147,N_6361,N_6217);
and U9148 (N_9148,N_6413,N_5650);
nor U9149 (N_9149,N_5103,N_5280);
nor U9150 (N_9150,N_6137,N_6079);
nand U9151 (N_9151,N_6107,N_7093);
nand U9152 (N_9152,N_5767,N_5512);
and U9153 (N_9153,N_5798,N_7058);
nand U9154 (N_9154,N_5108,N_7256);
xor U9155 (N_9155,N_5810,N_5117);
nand U9156 (N_9156,N_5988,N_6530);
or U9157 (N_9157,N_6117,N_6512);
nor U9158 (N_9158,N_5674,N_7445);
or U9159 (N_9159,N_7313,N_7026);
nand U9160 (N_9160,N_5882,N_5206);
xnor U9161 (N_9161,N_7122,N_5324);
nor U9162 (N_9162,N_5314,N_6000);
xnor U9163 (N_9163,N_6470,N_5276);
or U9164 (N_9164,N_7326,N_7444);
and U9165 (N_9165,N_6869,N_6726);
xnor U9166 (N_9166,N_6715,N_6561);
and U9167 (N_9167,N_5564,N_5576);
or U9168 (N_9168,N_5186,N_5033);
nand U9169 (N_9169,N_5753,N_6203);
nand U9170 (N_9170,N_5992,N_5936);
xor U9171 (N_9171,N_6512,N_6324);
or U9172 (N_9172,N_5511,N_6290);
or U9173 (N_9173,N_6621,N_5712);
nand U9174 (N_9174,N_6831,N_6868);
xor U9175 (N_9175,N_6868,N_6699);
or U9176 (N_9176,N_5882,N_7225);
xnor U9177 (N_9177,N_5628,N_7453);
or U9178 (N_9178,N_5011,N_7068);
nor U9179 (N_9179,N_5747,N_5309);
nand U9180 (N_9180,N_6482,N_5803);
or U9181 (N_9181,N_6368,N_6831);
nor U9182 (N_9182,N_5650,N_6005);
nand U9183 (N_9183,N_7236,N_5909);
and U9184 (N_9184,N_5730,N_6492);
nor U9185 (N_9185,N_5584,N_7201);
nor U9186 (N_9186,N_5048,N_5267);
nor U9187 (N_9187,N_7031,N_6889);
nand U9188 (N_9188,N_6063,N_6573);
nand U9189 (N_9189,N_6221,N_5212);
nor U9190 (N_9190,N_5813,N_6650);
nand U9191 (N_9191,N_5611,N_6370);
xnor U9192 (N_9192,N_5727,N_6366);
nor U9193 (N_9193,N_5787,N_6870);
nand U9194 (N_9194,N_6103,N_5722);
xor U9195 (N_9195,N_5856,N_7310);
or U9196 (N_9196,N_5509,N_5188);
nor U9197 (N_9197,N_6600,N_5320);
nor U9198 (N_9198,N_7291,N_5231);
nand U9199 (N_9199,N_5306,N_6183);
or U9200 (N_9200,N_6396,N_6355);
or U9201 (N_9201,N_5961,N_6717);
or U9202 (N_9202,N_5595,N_6521);
nor U9203 (N_9203,N_7196,N_6186);
nor U9204 (N_9204,N_5298,N_6101);
and U9205 (N_9205,N_6307,N_5396);
nand U9206 (N_9206,N_6323,N_6753);
xnor U9207 (N_9207,N_6144,N_6450);
or U9208 (N_9208,N_7295,N_6282);
nand U9209 (N_9209,N_7254,N_5106);
nand U9210 (N_9210,N_5102,N_7207);
and U9211 (N_9211,N_7395,N_5697);
nand U9212 (N_9212,N_5627,N_7488);
or U9213 (N_9213,N_6157,N_5112);
xor U9214 (N_9214,N_6467,N_7325);
nor U9215 (N_9215,N_5228,N_6537);
nor U9216 (N_9216,N_6336,N_5021);
and U9217 (N_9217,N_7378,N_5422);
or U9218 (N_9218,N_5847,N_6815);
nand U9219 (N_9219,N_6843,N_6679);
or U9220 (N_9220,N_6640,N_5432);
and U9221 (N_9221,N_6767,N_5612);
and U9222 (N_9222,N_7080,N_6640);
and U9223 (N_9223,N_6192,N_6919);
nor U9224 (N_9224,N_5644,N_5960);
nor U9225 (N_9225,N_5538,N_5114);
xor U9226 (N_9226,N_6157,N_5119);
nor U9227 (N_9227,N_5727,N_5199);
nand U9228 (N_9228,N_7211,N_6519);
xnor U9229 (N_9229,N_6216,N_5879);
nand U9230 (N_9230,N_5642,N_6254);
and U9231 (N_9231,N_6748,N_6185);
nand U9232 (N_9232,N_6347,N_6270);
or U9233 (N_9233,N_5292,N_5237);
xor U9234 (N_9234,N_6122,N_6548);
and U9235 (N_9235,N_6782,N_7352);
nor U9236 (N_9236,N_5879,N_5236);
and U9237 (N_9237,N_6282,N_6188);
xnor U9238 (N_9238,N_6252,N_5352);
nor U9239 (N_9239,N_5736,N_7375);
nor U9240 (N_9240,N_6973,N_5795);
and U9241 (N_9241,N_6062,N_6046);
or U9242 (N_9242,N_5451,N_7336);
xor U9243 (N_9243,N_5245,N_7409);
or U9244 (N_9244,N_7396,N_6017);
nor U9245 (N_9245,N_5466,N_5564);
xnor U9246 (N_9246,N_5038,N_5582);
nand U9247 (N_9247,N_7367,N_5595);
and U9248 (N_9248,N_6023,N_7060);
or U9249 (N_9249,N_6431,N_7003);
or U9250 (N_9250,N_5091,N_6765);
nor U9251 (N_9251,N_6972,N_6111);
xnor U9252 (N_9252,N_5943,N_6034);
xnor U9253 (N_9253,N_5773,N_5998);
and U9254 (N_9254,N_5518,N_5280);
xor U9255 (N_9255,N_5754,N_7435);
xor U9256 (N_9256,N_5227,N_5330);
and U9257 (N_9257,N_7377,N_7422);
or U9258 (N_9258,N_6430,N_6659);
nor U9259 (N_9259,N_7239,N_6841);
xor U9260 (N_9260,N_6768,N_6560);
and U9261 (N_9261,N_5521,N_5020);
nand U9262 (N_9262,N_6089,N_5256);
and U9263 (N_9263,N_6273,N_6288);
nor U9264 (N_9264,N_5865,N_6695);
and U9265 (N_9265,N_5704,N_6698);
and U9266 (N_9266,N_7389,N_6697);
xnor U9267 (N_9267,N_6656,N_6911);
nand U9268 (N_9268,N_5092,N_7158);
nor U9269 (N_9269,N_6751,N_7019);
nor U9270 (N_9270,N_5873,N_6303);
nor U9271 (N_9271,N_7147,N_7002);
xor U9272 (N_9272,N_5345,N_7259);
or U9273 (N_9273,N_5915,N_6669);
xnor U9274 (N_9274,N_7343,N_5415);
or U9275 (N_9275,N_5510,N_7354);
nor U9276 (N_9276,N_5257,N_7054);
and U9277 (N_9277,N_6959,N_5669);
nand U9278 (N_9278,N_6227,N_7161);
nand U9279 (N_9279,N_6256,N_6273);
nand U9280 (N_9280,N_6508,N_6418);
nand U9281 (N_9281,N_6739,N_6097);
nand U9282 (N_9282,N_5170,N_6714);
or U9283 (N_9283,N_5610,N_5666);
xnor U9284 (N_9284,N_6783,N_6906);
or U9285 (N_9285,N_7474,N_6343);
xor U9286 (N_9286,N_6139,N_7181);
or U9287 (N_9287,N_6989,N_6064);
or U9288 (N_9288,N_5190,N_6479);
and U9289 (N_9289,N_6877,N_7223);
xor U9290 (N_9290,N_6600,N_5871);
nor U9291 (N_9291,N_6677,N_5685);
and U9292 (N_9292,N_5508,N_5920);
xor U9293 (N_9293,N_5599,N_6220);
nand U9294 (N_9294,N_6072,N_5907);
nor U9295 (N_9295,N_6132,N_5956);
nand U9296 (N_9296,N_5730,N_7318);
and U9297 (N_9297,N_5918,N_6382);
or U9298 (N_9298,N_5407,N_5424);
and U9299 (N_9299,N_7397,N_6017);
or U9300 (N_9300,N_5174,N_7469);
or U9301 (N_9301,N_6575,N_5555);
nand U9302 (N_9302,N_6094,N_6496);
nor U9303 (N_9303,N_6274,N_5232);
and U9304 (N_9304,N_7081,N_5608);
nand U9305 (N_9305,N_6031,N_6464);
xor U9306 (N_9306,N_5433,N_7130);
xnor U9307 (N_9307,N_6473,N_5136);
or U9308 (N_9308,N_5532,N_6779);
nand U9309 (N_9309,N_7186,N_7103);
or U9310 (N_9310,N_7497,N_7104);
nor U9311 (N_9311,N_5717,N_5871);
nand U9312 (N_9312,N_6725,N_5595);
and U9313 (N_9313,N_5989,N_5244);
xor U9314 (N_9314,N_5416,N_5257);
and U9315 (N_9315,N_7437,N_6555);
nor U9316 (N_9316,N_6828,N_6726);
and U9317 (N_9317,N_7216,N_5462);
xnor U9318 (N_9318,N_6427,N_5806);
and U9319 (N_9319,N_7130,N_6431);
or U9320 (N_9320,N_5263,N_5248);
or U9321 (N_9321,N_5912,N_6440);
nor U9322 (N_9322,N_7014,N_7301);
xnor U9323 (N_9323,N_5678,N_5128);
nand U9324 (N_9324,N_5329,N_7372);
nand U9325 (N_9325,N_5007,N_5765);
nand U9326 (N_9326,N_5905,N_7441);
or U9327 (N_9327,N_6405,N_6768);
nand U9328 (N_9328,N_6549,N_6762);
xnor U9329 (N_9329,N_5281,N_7050);
or U9330 (N_9330,N_6271,N_7429);
xor U9331 (N_9331,N_6947,N_5980);
or U9332 (N_9332,N_5770,N_7133);
and U9333 (N_9333,N_5997,N_6752);
or U9334 (N_9334,N_6151,N_5687);
nor U9335 (N_9335,N_5413,N_5595);
nor U9336 (N_9336,N_6409,N_7272);
xor U9337 (N_9337,N_7196,N_5475);
and U9338 (N_9338,N_6835,N_6249);
or U9339 (N_9339,N_5689,N_6481);
nand U9340 (N_9340,N_5948,N_5503);
nor U9341 (N_9341,N_6969,N_6933);
and U9342 (N_9342,N_6624,N_7376);
xor U9343 (N_9343,N_6942,N_5217);
nor U9344 (N_9344,N_6527,N_6386);
nor U9345 (N_9345,N_5073,N_5056);
nand U9346 (N_9346,N_5160,N_7319);
and U9347 (N_9347,N_5379,N_6933);
and U9348 (N_9348,N_6222,N_5768);
and U9349 (N_9349,N_5395,N_5081);
nor U9350 (N_9350,N_5255,N_5659);
and U9351 (N_9351,N_7259,N_7305);
nand U9352 (N_9352,N_7276,N_5232);
nand U9353 (N_9353,N_6658,N_5229);
nand U9354 (N_9354,N_7293,N_7276);
nand U9355 (N_9355,N_6137,N_6128);
nor U9356 (N_9356,N_6823,N_5397);
or U9357 (N_9357,N_7190,N_5637);
xnor U9358 (N_9358,N_6268,N_6549);
xnor U9359 (N_9359,N_5319,N_7139);
and U9360 (N_9360,N_6101,N_5752);
nand U9361 (N_9361,N_5060,N_6455);
xor U9362 (N_9362,N_5879,N_6407);
or U9363 (N_9363,N_7024,N_5233);
or U9364 (N_9364,N_5581,N_5635);
nor U9365 (N_9365,N_5320,N_5949);
xor U9366 (N_9366,N_6412,N_7136);
xnor U9367 (N_9367,N_6428,N_7317);
nand U9368 (N_9368,N_5055,N_6518);
xnor U9369 (N_9369,N_7225,N_6272);
nand U9370 (N_9370,N_5948,N_7001);
nand U9371 (N_9371,N_7000,N_7404);
xor U9372 (N_9372,N_7052,N_7438);
and U9373 (N_9373,N_6463,N_5394);
and U9374 (N_9374,N_5811,N_6072);
or U9375 (N_9375,N_5915,N_7212);
and U9376 (N_9376,N_5357,N_5503);
or U9377 (N_9377,N_6499,N_5645);
nor U9378 (N_9378,N_5327,N_6046);
nor U9379 (N_9379,N_5796,N_7182);
nand U9380 (N_9380,N_5602,N_5423);
or U9381 (N_9381,N_7232,N_5032);
or U9382 (N_9382,N_6004,N_7078);
and U9383 (N_9383,N_6697,N_5874);
and U9384 (N_9384,N_5736,N_6341);
xnor U9385 (N_9385,N_6219,N_5530);
or U9386 (N_9386,N_6846,N_5634);
xor U9387 (N_9387,N_6704,N_6088);
nor U9388 (N_9388,N_7228,N_5558);
nor U9389 (N_9389,N_6751,N_6356);
nand U9390 (N_9390,N_5818,N_6532);
or U9391 (N_9391,N_7158,N_7328);
or U9392 (N_9392,N_5512,N_7314);
xnor U9393 (N_9393,N_6648,N_5045);
and U9394 (N_9394,N_5714,N_5147);
xnor U9395 (N_9395,N_5203,N_5138);
xnor U9396 (N_9396,N_6210,N_6883);
or U9397 (N_9397,N_6555,N_5550);
and U9398 (N_9398,N_5960,N_6024);
xor U9399 (N_9399,N_5422,N_5893);
nand U9400 (N_9400,N_5738,N_6677);
and U9401 (N_9401,N_5512,N_5373);
and U9402 (N_9402,N_7038,N_7309);
nand U9403 (N_9403,N_5293,N_5060);
nor U9404 (N_9404,N_5019,N_6445);
and U9405 (N_9405,N_7336,N_5912);
and U9406 (N_9406,N_5744,N_5751);
nand U9407 (N_9407,N_5144,N_6132);
and U9408 (N_9408,N_5863,N_5292);
and U9409 (N_9409,N_7130,N_5001);
or U9410 (N_9410,N_5035,N_6924);
and U9411 (N_9411,N_6956,N_6154);
nor U9412 (N_9412,N_6739,N_6243);
nand U9413 (N_9413,N_7342,N_5238);
or U9414 (N_9414,N_6416,N_6934);
xor U9415 (N_9415,N_7439,N_5654);
xnor U9416 (N_9416,N_6396,N_5836);
nor U9417 (N_9417,N_6118,N_6866);
or U9418 (N_9418,N_7449,N_6928);
nor U9419 (N_9419,N_7035,N_5874);
and U9420 (N_9420,N_6954,N_6564);
xor U9421 (N_9421,N_5252,N_6971);
or U9422 (N_9422,N_6842,N_6095);
nand U9423 (N_9423,N_5932,N_7241);
xor U9424 (N_9424,N_6451,N_5744);
xnor U9425 (N_9425,N_6543,N_7116);
xnor U9426 (N_9426,N_5762,N_6204);
xnor U9427 (N_9427,N_6265,N_5424);
and U9428 (N_9428,N_7354,N_6320);
or U9429 (N_9429,N_6381,N_7363);
nand U9430 (N_9430,N_5858,N_5661);
or U9431 (N_9431,N_6894,N_7363);
nor U9432 (N_9432,N_5290,N_7249);
and U9433 (N_9433,N_6164,N_7454);
and U9434 (N_9434,N_7088,N_7092);
xor U9435 (N_9435,N_7152,N_5646);
nor U9436 (N_9436,N_5093,N_7029);
xnor U9437 (N_9437,N_5829,N_5402);
xor U9438 (N_9438,N_6253,N_7310);
xnor U9439 (N_9439,N_6630,N_6463);
or U9440 (N_9440,N_6589,N_5996);
or U9441 (N_9441,N_7201,N_7089);
and U9442 (N_9442,N_7306,N_5902);
nand U9443 (N_9443,N_6745,N_6969);
or U9444 (N_9444,N_5173,N_7459);
nand U9445 (N_9445,N_7002,N_6181);
nand U9446 (N_9446,N_5395,N_5228);
xor U9447 (N_9447,N_6396,N_6077);
nand U9448 (N_9448,N_5489,N_6304);
xnor U9449 (N_9449,N_7395,N_7488);
nand U9450 (N_9450,N_6663,N_7173);
and U9451 (N_9451,N_5662,N_5159);
xor U9452 (N_9452,N_7248,N_6556);
nor U9453 (N_9453,N_7175,N_5976);
and U9454 (N_9454,N_6361,N_6435);
or U9455 (N_9455,N_6156,N_6306);
nor U9456 (N_9456,N_5042,N_6706);
nor U9457 (N_9457,N_6358,N_6634);
xnor U9458 (N_9458,N_7487,N_7161);
or U9459 (N_9459,N_5990,N_5041);
nor U9460 (N_9460,N_7323,N_7026);
xnor U9461 (N_9461,N_6111,N_6010);
xnor U9462 (N_9462,N_7003,N_5701);
nor U9463 (N_9463,N_6248,N_6029);
or U9464 (N_9464,N_5261,N_6345);
nand U9465 (N_9465,N_5468,N_6473);
nand U9466 (N_9466,N_6775,N_6888);
nand U9467 (N_9467,N_5886,N_6312);
nor U9468 (N_9468,N_6109,N_6932);
and U9469 (N_9469,N_7410,N_7132);
xnor U9470 (N_9470,N_7346,N_5774);
or U9471 (N_9471,N_5752,N_6212);
nor U9472 (N_9472,N_6749,N_6657);
and U9473 (N_9473,N_6792,N_5403);
nand U9474 (N_9474,N_6591,N_7034);
xor U9475 (N_9475,N_6739,N_5416);
nand U9476 (N_9476,N_5686,N_5382);
nand U9477 (N_9477,N_6594,N_6702);
and U9478 (N_9478,N_6118,N_5824);
and U9479 (N_9479,N_6198,N_5176);
nand U9480 (N_9480,N_7137,N_5280);
nand U9481 (N_9481,N_7374,N_7323);
nand U9482 (N_9482,N_5460,N_6222);
xnor U9483 (N_9483,N_5785,N_6330);
and U9484 (N_9484,N_6562,N_7407);
xor U9485 (N_9485,N_6355,N_5039);
and U9486 (N_9486,N_6825,N_6272);
or U9487 (N_9487,N_5123,N_6283);
nand U9488 (N_9488,N_5413,N_5669);
nor U9489 (N_9489,N_5175,N_6521);
nand U9490 (N_9490,N_7438,N_5588);
nor U9491 (N_9491,N_5286,N_6453);
and U9492 (N_9492,N_5532,N_6541);
nand U9493 (N_9493,N_6995,N_6758);
xor U9494 (N_9494,N_6953,N_5154);
and U9495 (N_9495,N_7105,N_5427);
nand U9496 (N_9496,N_7028,N_6053);
or U9497 (N_9497,N_5280,N_5154);
or U9498 (N_9498,N_6527,N_6773);
nand U9499 (N_9499,N_6111,N_5036);
and U9500 (N_9500,N_6171,N_6377);
and U9501 (N_9501,N_7084,N_6803);
or U9502 (N_9502,N_5049,N_6901);
nand U9503 (N_9503,N_6594,N_6801);
nor U9504 (N_9504,N_5890,N_5330);
and U9505 (N_9505,N_7351,N_5497);
xnor U9506 (N_9506,N_5620,N_6824);
xnor U9507 (N_9507,N_5046,N_6423);
or U9508 (N_9508,N_5639,N_5242);
or U9509 (N_9509,N_5561,N_5246);
nor U9510 (N_9510,N_6892,N_6062);
nand U9511 (N_9511,N_5166,N_7200);
xor U9512 (N_9512,N_6405,N_6913);
or U9513 (N_9513,N_6218,N_6372);
or U9514 (N_9514,N_5749,N_5361);
nand U9515 (N_9515,N_5010,N_7030);
nand U9516 (N_9516,N_6099,N_6488);
and U9517 (N_9517,N_5470,N_6916);
nor U9518 (N_9518,N_7162,N_6983);
xnor U9519 (N_9519,N_6032,N_6907);
or U9520 (N_9520,N_5749,N_6311);
or U9521 (N_9521,N_5191,N_5085);
or U9522 (N_9522,N_7367,N_7364);
nor U9523 (N_9523,N_6096,N_5901);
xnor U9524 (N_9524,N_7303,N_6618);
nand U9525 (N_9525,N_5829,N_6662);
and U9526 (N_9526,N_6387,N_6507);
xnor U9527 (N_9527,N_6358,N_6915);
nand U9528 (N_9528,N_5795,N_5140);
xnor U9529 (N_9529,N_6507,N_5798);
nand U9530 (N_9530,N_6267,N_6544);
and U9531 (N_9531,N_5378,N_7065);
xor U9532 (N_9532,N_6327,N_6981);
xor U9533 (N_9533,N_7120,N_5946);
nand U9534 (N_9534,N_5360,N_5557);
nor U9535 (N_9535,N_5903,N_5062);
and U9536 (N_9536,N_7356,N_6734);
and U9537 (N_9537,N_5692,N_6250);
nor U9538 (N_9538,N_5053,N_5871);
nand U9539 (N_9539,N_6201,N_7076);
or U9540 (N_9540,N_6749,N_6525);
or U9541 (N_9541,N_6604,N_6972);
or U9542 (N_9542,N_5551,N_6364);
or U9543 (N_9543,N_7131,N_5066);
and U9544 (N_9544,N_6394,N_6352);
nand U9545 (N_9545,N_6824,N_6063);
or U9546 (N_9546,N_6783,N_7222);
nand U9547 (N_9547,N_7441,N_6652);
or U9548 (N_9548,N_6032,N_5579);
nand U9549 (N_9549,N_6584,N_7160);
nor U9550 (N_9550,N_5084,N_5265);
xor U9551 (N_9551,N_7317,N_5939);
xnor U9552 (N_9552,N_6206,N_5471);
nand U9553 (N_9553,N_5994,N_6192);
nor U9554 (N_9554,N_6394,N_5940);
or U9555 (N_9555,N_6848,N_6703);
nand U9556 (N_9556,N_5605,N_5595);
nor U9557 (N_9557,N_6849,N_5536);
or U9558 (N_9558,N_7056,N_6253);
xor U9559 (N_9559,N_5829,N_5273);
and U9560 (N_9560,N_6130,N_7386);
nand U9561 (N_9561,N_5355,N_6584);
nand U9562 (N_9562,N_5472,N_5771);
nor U9563 (N_9563,N_6714,N_6157);
xnor U9564 (N_9564,N_5725,N_7365);
or U9565 (N_9565,N_7346,N_7403);
or U9566 (N_9566,N_5401,N_7276);
and U9567 (N_9567,N_7404,N_5393);
or U9568 (N_9568,N_6958,N_6631);
nor U9569 (N_9569,N_6445,N_7162);
nor U9570 (N_9570,N_7135,N_6217);
nor U9571 (N_9571,N_5295,N_6386);
xnor U9572 (N_9572,N_6688,N_7067);
nor U9573 (N_9573,N_5766,N_5908);
nor U9574 (N_9574,N_7028,N_7084);
nand U9575 (N_9575,N_6781,N_5992);
nor U9576 (N_9576,N_7092,N_6483);
and U9577 (N_9577,N_6874,N_6226);
nand U9578 (N_9578,N_6335,N_5519);
nor U9579 (N_9579,N_6615,N_6737);
or U9580 (N_9580,N_5876,N_6183);
nand U9581 (N_9581,N_5946,N_7132);
nor U9582 (N_9582,N_6275,N_5304);
or U9583 (N_9583,N_5255,N_6538);
nand U9584 (N_9584,N_5564,N_6668);
and U9585 (N_9585,N_6096,N_7194);
nor U9586 (N_9586,N_6128,N_6678);
nor U9587 (N_9587,N_6060,N_5458);
xnor U9588 (N_9588,N_7404,N_5277);
nand U9589 (N_9589,N_6233,N_7004);
or U9590 (N_9590,N_7087,N_6493);
nor U9591 (N_9591,N_5553,N_7214);
xnor U9592 (N_9592,N_6263,N_6877);
nor U9593 (N_9593,N_7286,N_6413);
nand U9594 (N_9594,N_5437,N_5469);
or U9595 (N_9595,N_6360,N_7308);
xor U9596 (N_9596,N_6093,N_6445);
nand U9597 (N_9597,N_5395,N_7441);
nand U9598 (N_9598,N_6396,N_5715);
xor U9599 (N_9599,N_5748,N_7382);
nor U9600 (N_9600,N_6382,N_6277);
nand U9601 (N_9601,N_5314,N_6531);
nand U9602 (N_9602,N_6400,N_6826);
and U9603 (N_9603,N_5460,N_5691);
nor U9604 (N_9604,N_5817,N_5306);
or U9605 (N_9605,N_6012,N_7138);
and U9606 (N_9606,N_5601,N_5631);
xor U9607 (N_9607,N_5702,N_5102);
and U9608 (N_9608,N_5740,N_7053);
nand U9609 (N_9609,N_5225,N_5866);
nand U9610 (N_9610,N_6223,N_5856);
and U9611 (N_9611,N_5780,N_5794);
or U9612 (N_9612,N_6455,N_5641);
nor U9613 (N_9613,N_6738,N_5359);
or U9614 (N_9614,N_7438,N_5619);
or U9615 (N_9615,N_5161,N_5814);
and U9616 (N_9616,N_5364,N_5490);
or U9617 (N_9617,N_6110,N_7220);
nand U9618 (N_9618,N_6630,N_5053);
and U9619 (N_9619,N_6265,N_7488);
or U9620 (N_9620,N_5085,N_6613);
or U9621 (N_9621,N_7223,N_7122);
or U9622 (N_9622,N_5666,N_5819);
nand U9623 (N_9623,N_5924,N_6279);
nor U9624 (N_9624,N_7199,N_6063);
and U9625 (N_9625,N_5038,N_6691);
or U9626 (N_9626,N_6112,N_6466);
nor U9627 (N_9627,N_5608,N_6570);
and U9628 (N_9628,N_7106,N_5745);
nor U9629 (N_9629,N_5229,N_5374);
and U9630 (N_9630,N_5696,N_6006);
and U9631 (N_9631,N_6194,N_6307);
nor U9632 (N_9632,N_6491,N_5342);
or U9633 (N_9633,N_7047,N_5121);
xnor U9634 (N_9634,N_5759,N_6934);
nand U9635 (N_9635,N_5947,N_5993);
nand U9636 (N_9636,N_6923,N_5989);
or U9637 (N_9637,N_6442,N_6766);
nor U9638 (N_9638,N_5288,N_7254);
nand U9639 (N_9639,N_6623,N_7238);
and U9640 (N_9640,N_7481,N_6989);
xnor U9641 (N_9641,N_7220,N_5640);
nand U9642 (N_9642,N_5374,N_5050);
or U9643 (N_9643,N_6169,N_6995);
or U9644 (N_9644,N_6927,N_7381);
or U9645 (N_9645,N_6592,N_7083);
nand U9646 (N_9646,N_6661,N_5279);
nor U9647 (N_9647,N_6960,N_5306);
nand U9648 (N_9648,N_7209,N_7107);
nand U9649 (N_9649,N_5592,N_5446);
and U9650 (N_9650,N_5313,N_7072);
xnor U9651 (N_9651,N_6602,N_7248);
nand U9652 (N_9652,N_6790,N_6063);
or U9653 (N_9653,N_7072,N_6485);
nand U9654 (N_9654,N_5566,N_7447);
or U9655 (N_9655,N_5713,N_6568);
xnor U9656 (N_9656,N_5263,N_6420);
and U9657 (N_9657,N_5604,N_6860);
nand U9658 (N_9658,N_5482,N_5144);
and U9659 (N_9659,N_7140,N_6099);
nand U9660 (N_9660,N_6326,N_5852);
nand U9661 (N_9661,N_5857,N_7370);
xnor U9662 (N_9662,N_5324,N_7071);
nor U9663 (N_9663,N_6260,N_7242);
and U9664 (N_9664,N_5237,N_5497);
nand U9665 (N_9665,N_7061,N_7191);
nand U9666 (N_9666,N_6371,N_5567);
and U9667 (N_9667,N_5695,N_7217);
or U9668 (N_9668,N_5455,N_6511);
or U9669 (N_9669,N_6124,N_7343);
and U9670 (N_9670,N_6396,N_6851);
nand U9671 (N_9671,N_5339,N_6261);
xor U9672 (N_9672,N_7088,N_5271);
or U9673 (N_9673,N_6775,N_6378);
and U9674 (N_9674,N_5533,N_5161);
xnor U9675 (N_9675,N_6041,N_5870);
nor U9676 (N_9676,N_6096,N_5472);
or U9677 (N_9677,N_7410,N_5666);
nor U9678 (N_9678,N_6658,N_5656);
xor U9679 (N_9679,N_7210,N_5134);
xor U9680 (N_9680,N_6604,N_6264);
and U9681 (N_9681,N_6079,N_6894);
nand U9682 (N_9682,N_5209,N_7093);
or U9683 (N_9683,N_5045,N_7373);
nor U9684 (N_9684,N_5035,N_6650);
nor U9685 (N_9685,N_6904,N_5479);
nor U9686 (N_9686,N_6403,N_6918);
or U9687 (N_9687,N_6956,N_7378);
nand U9688 (N_9688,N_5293,N_7202);
xnor U9689 (N_9689,N_7326,N_7475);
and U9690 (N_9690,N_5347,N_6781);
nand U9691 (N_9691,N_5565,N_6006);
or U9692 (N_9692,N_6027,N_5851);
or U9693 (N_9693,N_5087,N_5247);
or U9694 (N_9694,N_6448,N_5567);
or U9695 (N_9695,N_6438,N_6739);
or U9696 (N_9696,N_5260,N_6862);
and U9697 (N_9697,N_5245,N_7149);
nand U9698 (N_9698,N_7340,N_5801);
xnor U9699 (N_9699,N_7276,N_6407);
or U9700 (N_9700,N_6046,N_6352);
nand U9701 (N_9701,N_6311,N_5586);
or U9702 (N_9702,N_5296,N_7366);
xnor U9703 (N_9703,N_5017,N_5500);
xnor U9704 (N_9704,N_6617,N_6845);
xor U9705 (N_9705,N_6917,N_6826);
and U9706 (N_9706,N_7116,N_7469);
xor U9707 (N_9707,N_6212,N_5329);
nor U9708 (N_9708,N_6342,N_7104);
and U9709 (N_9709,N_5199,N_6776);
nand U9710 (N_9710,N_6988,N_5679);
or U9711 (N_9711,N_5023,N_6863);
xnor U9712 (N_9712,N_5577,N_6656);
xor U9713 (N_9713,N_6765,N_7205);
or U9714 (N_9714,N_5237,N_6667);
and U9715 (N_9715,N_6062,N_6163);
nand U9716 (N_9716,N_6448,N_6121);
or U9717 (N_9717,N_6401,N_5382);
xor U9718 (N_9718,N_7074,N_5869);
or U9719 (N_9719,N_7429,N_5040);
xnor U9720 (N_9720,N_6684,N_5263);
nand U9721 (N_9721,N_5333,N_6834);
and U9722 (N_9722,N_5317,N_7179);
xor U9723 (N_9723,N_6930,N_5569);
or U9724 (N_9724,N_5787,N_6221);
nand U9725 (N_9725,N_5667,N_7482);
nand U9726 (N_9726,N_6408,N_5002);
or U9727 (N_9727,N_6583,N_7129);
or U9728 (N_9728,N_6979,N_7441);
nor U9729 (N_9729,N_5444,N_6697);
or U9730 (N_9730,N_7003,N_6938);
and U9731 (N_9731,N_5971,N_5078);
and U9732 (N_9732,N_6232,N_6661);
nand U9733 (N_9733,N_6179,N_5687);
xnor U9734 (N_9734,N_6590,N_6297);
or U9735 (N_9735,N_5869,N_7425);
and U9736 (N_9736,N_6890,N_6209);
or U9737 (N_9737,N_5504,N_6134);
or U9738 (N_9738,N_5430,N_6227);
nor U9739 (N_9739,N_5571,N_6560);
and U9740 (N_9740,N_5568,N_6292);
nor U9741 (N_9741,N_5813,N_7400);
or U9742 (N_9742,N_5681,N_6527);
or U9743 (N_9743,N_7390,N_6543);
nor U9744 (N_9744,N_6673,N_6400);
nor U9745 (N_9745,N_5749,N_6765);
xnor U9746 (N_9746,N_7355,N_7044);
xor U9747 (N_9747,N_6359,N_5486);
nand U9748 (N_9748,N_5408,N_6712);
nor U9749 (N_9749,N_6952,N_5080);
or U9750 (N_9750,N_7446,N_5467);
or U9751 (N_9751,N_6628,N_6492);
and U9752 (N_9752,N_5560,N_5452);
nor U9753 (N_9753,N_7013,N_5687);
or U9754 (N_9754,N_6574,N_5765);
nor U9755 (N_9755,N_5662,N_5869);
or U9756 (N_9756,N_6106,N_6532);
nor U9757 (N_9757,N_7400,N_5413);
and U9758 (N_9758,N_7406,N_6797);
xnor U9759 (N_9759,N_6137,N_5111);
and U9760 (N_9760,N_5666,N_7062);
xor U9761 (N_9761,N_6911,N_5328);
xnor U9762 (N_9762,N_5362,N_5447);
nor U9763 (N_9763,N_5225,N_5691);
and U9764 (N_9764,N_5494,N_6530);
nor U9765 (N_9765,N_6204,N_5994);
or U9766 (N_9766,N_5898,N_5021);
and U9767 (N_9767,N_6560,N_5010);
or U9768 (N_9768,N_5421,N_5976);
nand U9769 (N_9769,N_7239,N_6986);
nor U9770 (N_9770,N_5096,N_5661);
nor U9771 (N_9771,N_5933,N_7069);
or U9772 (N_9772,N_6149,N_6246);
nor U9773 (N_9773,N_6961,N_5696);
or U9774 (N_9774,N_5213,N_5953);
or U9775 (N_9775,N_6904,N_7083);
or U9776 (N_9776,N_6993,N_7223);
nand U9777 (N_9777,N_5506,N_6951);
nor U9778 (N_9778,N_7400,N_6746);
and U9779 (N_9779,N_5181,N_6403);
and U9780 (N_9780,N_7069,N_6532);
nand U9781 (N_9781,N_5576,N_6417);
or U9782 (N_9782,N_7486,N_7228);
xnor U9783 (N_9783,N_5849,N_6882);
nand U9784 (N_9784,N_7442,N_6979);
and U9785 (N_9785,N_5668,N_5640);
xor U9786 (N_9786,N_6170,N_6712);
and U9787 (N_9787,N_5130,N_6821);
nand U9788 (N_9788,N_6179,N_6332);
and U9789 (N_9789,N_5014,N_6819);
and U9790 (N_9790,N_5711,N_7099);
and U9791 (N_9791,N_5192,N_6581);
nand U9792 (N_9792,N_5304,N_6606);
nor U9793 (N_9793,N_7462,N_5899);
and U9794 (N_9794,N_6884,N_7363);
or U9795 (N_9795,N_7314,N_6173);
or U9796 (N_9796,N_7195,N_6123);
and U9797 (N_9797,N_7072,N_5072);
xnor U9798 (N_9798,N_6873,N_7064);
nand U9799 (N_9799,N_5782,N_6348);
nand U9800 (N_9800,N_5443,N_7276);
nor U9801 (N_9801,N_6585,N_6171);
nand U9802 (N_9802,N_5043,N_5349);
nor U9803 (N_9803,N_6752,N_5875);
and U9804 (N_9804,N_6787,N_7333);
or U9805 (N_9805,N_7201,N_7146);
or U9806 (N_9806,N_5008,N_6675);
or U9807 (N_9807,N_6742,N_6131);
xor U9808 (N_9808,N_5317,N_6619);
xnor U9809 (N_9809,N_5523,N_5980);
nand U9810 (N_9810,N_5708,N_6768);
and U9811 (N_9811,N_6919,N_5098);
and U9812 (N_9812,N_5149,N_5264);
xnor U9813 (N_9813,N_5180,N_6494);
and U9814 (N_9814,N_7062,N_5498);
or U9815 (N_9815,N_5814,N_6881);
xnor U9816 (N_9816,N_5045,N_7377);
and U9817 (N_9817,N_6250,N_5501);
or U9818 (N_9818,N_7186,N_6435);
or U9819 (N_9819,N_5560,N_5279);
or U9820 (N_9820,N_6728,N_6462);
nand U9821 (N_9821,N_5452,N_5096);
or U9822 (N_9822,N_6254,N_7039);
nand U9823 (N_9823,N_5808,N_6043);
or U9824 (N_9824,N_5495,N_5255);
xnor U9825 (N_9825,N_6592,N_7426);
nor U9826 (N_9826,N_6655,N_7167);
and U9827 (N_9827,N_6018,N_7002);
nor U9828 (N_9828,N_6286,N_6150);
and U9829 (N_9829,N_5355,N_6508);
or U9830 (N_9830,N_7111,N_5874);
nor U9831 (N_9831,N_5371,N_7023);
nor U9832 (N_9832,N_6119,N_6120);
xnor U9833 (N_9833,N_5815,N_5483);
xor U9834 (N_9834,N_6260,N_6358);
xor U9835 (N_9835,N_7442,N_6285);
or U9836 (N_9836,N_6590,N_6691);
and U9837 (N_9837,N_7064,N_5527);
nand U9838 (N_9838,N_5064,N_6735);
nor U9839 (N_9839,N_7311,N_6617);
nor U9840 (N_9840,N_6227,N_7075);
and U9841 (N_9841,N_5449,N_6469);
and U9842 (N_9842,N_5823,N_5388);
xnor U9843 (N_9843,N_6432,N_6523);
nand U9844 (N_9844,N_5547,N_6785);
nand U9845 (N_9845,N_7332,N_7281);
nand U9846 (N_9846,N_5418,N_7311);
nor U9847 (N_9847,N_6944,N_5588);
or U9848 (N_9848,N_6945,N_7239);
nor U9849 (N_9849,N_7116,N_7388);
and U9850 (N_9850,N_6807,N_5665);
nor U9851 (N_9851,N_6541,N_6787);
nor U9852 (N_9852,N_5069,N_6975);
nor U9853 (N_9853,N_6554,N_6008);
or U9854 (N_9854,N_5455,N_6063);
xnor U9855 (N_9855,N_5969,N_5634);
or U9856 (N_9856,N_5467,N_7321);
xnor U9857 (N_9857,N_5638,N_6392);
or U9858 (N_9858,N_7401,N_6250);
and U9859 (N_9859,N_5931,N_7260);
and U9860 (N_9860,N_7291,N_7421);
and U9861 (N_9861,N_5087,N_7041);
or U9862 (N_9862,N_6710,N_6187);
nand U9863 (N_9863,N_6363,N_5863);
nor U9864 (N_9864,N_5793,N_6882);
or U9865 (N_9865,N_6131,N_5575);
and U9866 (N_9866,N_7130,N_5228);
or U9867 (N_9867,N_6313,N_6598);
nor U9868 (N_9868,N_6433,N_5725);
nor U9869 (N_9869,N_6795,N_6834);
or U9870 (N_9870,N_5640,N_5545);
or U9871 (N_9871,N_7059,N_5237);
or U9872 (N_9872,N_7215,N_6660);
or U9873 (N_9873,N_6447,N_5055);
or U9874 (N_9874,N_7481,N_5067);
or U9875 (N_9875,N_7400,N_6488);
nand U9876 (N_9876,N_5842,N_5903);
and U9877 (N_9877,N_5450,N_7368);
or U9878 (N_9878,N_5163,N_6241);
and U9879 (N_9879,N_6936,N_6413);
xnor U9880 (N_9880,N_6295,N_6569);
nand U9881 (N_9881,N_6837,N_5709);
xor U9882 (N_9882,N_5373,N_5590);
xnor U9883 (N_9883,N_5987,N_6619);
or U9884 (N_9884,N_5138,N_5576);
nand U9885 (N_9885,N_5789,N_6309);
and U9886 (N_9886,N_5652,N_5689);
or U9887 (N_9887,N_7235,N_7239);
or U9888 (N_9888,N_7204,N_7143);
xnor U9889 (N_9889,N_6762,N_6974);
or U9890 (N_9890,N_6527,N_7321);
and U9891 (N_9891,N_6277,N_6908);
xnor U9892 (N_9892,N_6034,N_5391);
nand U9893 (N_9893,N_7488,N_6644);
nor U9894 (N_9894,N_6297,N_6332);
xor U9895 (N_9895,N_5618,N_6835);
nand U9896 (N_9896,N_5702,N_5571);
nand U9897 (N_9897,N_7028,N_6775);
nand U9898 (N_9898,N_5906,N_5746);
nor U9899 (N_9899,N_5743,N_5137);
nand U9900 (N_9900,N_5287,N_5928);
or U9901 (N_9901,N_5692,N_6448);
nand U9902 (N_9902,N_6306,N_6713);
nor U9903 (N_9903,N_5758,N_5807);
nor U9904 (N_9904,N_7435,N_5778);
and U9905 (N_9905,N_6073,N_6275);
nor U9906 (N_9906,N_5266,N_5470);
or U9907 (N_9907,N_5151,N_5357);
xor U9908 (N_9908,N_5472,N_6867);
nand U9909 (N_9909,N_5369,N_7316);
and U9910 (N_9910,N_5423,N_6939);
nand U9911 (N_9911,N_6763,N_6661);
or U9912 (N_9912,N_6567,N_6185);
nor U9913 (N_9913,N_5384,N_7283);
or U9914 (N_9914,N_5769,N_6970);
xnor U9915 (N_9915,N_5826,N_5671);
nand U9916 (N_9916,N_5023,N_5848);
or U9917 (N_9917,N_6124,N_6581);
and U9918 (N_9918,N_6120,N_6053);
nand U9919 (N_9919,N_6675,N_6324);
nand U9920 (N_9920,N_5562,N_7417);
xor U9921 (N_9921,N_6878,N_5403);
nand U9922 (N_9922,N_5599,N_5580);
nor U9923 (N_9923,N_7256,N_5544);
nand U9924 (N_9924,N_7287,N_6294);
nand U9925 (N_9925,N_6727,N_7126);
xnor U9926 (N_9926,N_5601,N_5146);
or U9927 (N_9927,N_5111,N_5458);
xnor U9928 (N_9928,N_5137,N_7382);
nor U9929 (N_9929,N_6565,N_6950);
nor U9930 (N_9930,N_7201,N_5545);
and U9931 (N_9931,N_6530,N_6747);
or U9932 (N_9932,N_6376,N_7458);
nand U9933 (N_9933,N_5776,N_5390);
xor U9934 (N_9934,N_5510,N_6661);
nand U9935 (N_9935,N_5157,N_6682);
nor U9936 (N_9936,N_7345,N_6175);
xor U9937 (N_9937,N_6458,N_7106);
xor U9938 (N_9938,N_7323,N_6966);
nand U9939 (N_9939,N_5352,N_6612);
or U9940 (N_9940,N_5716,N_6345);
nor U9941 (N_9941,N_6965,N_6566);
and U9942 (N_9942,N_6974,N_5317);
nand U9943 (N_9943,N_5710,N_6458);
or U9944 (N_9944,N_5031,N_5968);
or U9945 (N_9945,N_7463,N_6630);
nor U9946 (N_9946,N_7148,N_7499);
nand U9947 (N_9947,N_5224,N_6283);
nand U9948 (N_9948,N_7355,N_7225);
nand U9949 (N_9949,N_5054,N_6535);
nor U9950 (N_9950,N_7050,N_5838);
and U9951 (N_9951,N_6299,N_7222);
nor U9952 (N_9952,N_6974,N_5009);
and U9953 (N_9953,N_6469,N_7098);
and U9954 (N_9954,N_5647,N_7349);
nor U9955 (N_9955,N_5965,N_6450);
and U9956 (N_9956,N_7102,N_5190);
or U9957 (N_9957,N_5266,N_6426);
nand U9958 (N_9958,N_6909,N_5312);
xor U9959 (N_9959,N_6559,N_6851);
or U9960 (N_9960,N_5349,N_7371);
xor U9961 (N_9961,N_5787,N_5489);
or U9962 (N_9962,N_7197,N_5545);
or U9963 (N_9963,N_6107,N_6019);
or U9964 (N_9964,N_5458,N_6231);
nand U9965 (N_9965,N_6445,N_7339);
nor U9966 (N_9966,N_5937,N_5113);
nand U9967 (N_9967,N_5172,N_5168);
or U9968 (N_9968,N_7286,N_6323);
xnor U9969 (N_9969,N_6328,N_6993);
nor U9970 (N_9970,N_7449,N_6528);
nor U9971 (N_9971,N_6461,N_6117);
xnor U9972 (N_9972,N_7447,N_6118);
nand U9973 (N_9973,N_6268,N_5578);
and U9974 (N_9974,N_6764,N_6009);
xor U9975 (N_9975,N_7444,N_6408);
xor U9976 (N_9976,N_5341,N_5440);
xor U9977 (N_9977,N_6224,N_7112);
nor U9978 (N_9978,N_5000,N_6700);
or U9979 (N_9979,N_5955,N_6245);
xor U9980 (N_9980,N_7086,N_6383);
and U9981 (N_9981,N_7341,N_7103);
and U9982 (N_9982,N_5649,N_5606);
nand U9983 (N_9983,N_7495,N_6088);
or U9984 (N_9984,N_7365,N_5671);
or U9985 (N_9985,N_6445,N_6051);
nor U9986 (N_9986,N_5288,N_7164);
nand U9987 (N_9987,N_6936,N_5608);
nor U9988 (N_9988,N_6149,N_5147);
nor U9989 (N_9989,N_6778,N_7415);
and U9990 (N_9990,N_6324,N_6309);
xnor U9991 (N_9991,N_6708,N_6473);
nor U9992 (N_9992,N_6856,N_7265);
or U9993 (N_9993,N_5297,N_6552);
or U9994 (N_9994,N_5706,N_6187);
or U9995 (N_9995,N_6377,N_6023);
nand U9996 (N_9996,N_6112,N_7141);
nand U9997 (N_9997,N_5617,N_5210);
xor U9998 (N_9998,N_5760,N_5799);
and U9999 (N_9999,N_7192,N_6682);
nand U10000 (N_10000,N_8068,N_8853);
xor U10001 (N_10001,N_8022,N_9280);
nand U10002 (N_10002,N_8042,N_8516);
or U10003 (N_10003,N_7995,N_9239);
xnor U10004 (N_10004,N_7606,N_7773);
nor U10005 (N_10005,N_9989,N_8844);
nand U10006 (N_10006,N_7749,N_9268);
nor U10007 (N_10007,N_9799,N_8429);
nor U10008 (N_10008,N_9534,N_7878);
nand U10009 (N_10009,N_8017,N_8778);
xnor U10010 (N_10010,N_8032,N_8897);
and U10011 (N_10011,N_8054,N_9889);
xor U10012 (N_10012,N_9862,N_9964);
nor U10013 (N_10013,N_8795,N_8999);
or U10014 (N_10014,N_8988,N_9297);
and U10015 (N_10015,N_8189,N_7691);
nand U10016 (N_10016,N_8887,N_7640);
nor U10017 (N_10017,N_9871,N_7513);
xor U10018 (N_10018,N_7521,N_7659);
and U10019 (N_10019,N_9109,N_8784);
or U10020 (N_10020,N_7619,N_9609);
nand U10021 (N_10021,N_9475,N_8125);
and U10022 (N_10022,N_7949,N_7567);
or U10023 (N_10023,N_9911,N_9221);
or U10024 (N_10024,N_7656,N_8761);
nand U10025 (N_10025,N_8615,N_9669);
and U10026 (N_10026,N_8435,N_9749);
nand U10027 (N_10027,N_7776,N_9736);
and U10028 (N_10028,N_8446,N_8820);
and U10029 (N_10029,N_8319,N_9107);
nor U10030 (N_10030,N_8771,N_9070);
and U10031 (N_10031,N_9357,N_7875);
and U10032 (N_10032,N_8779,N_9287);
xor U10033 (N_10033,N_9563,N_8324);
xor U10034 (N_10034,N_8184,N_8078);
xnor U10035 (N_10035,N_9513,N_9652);
nand U10036 (N_10036,N_7715,N_9433);
nor U10037 (N_10037,N_9486,N_7789);
xor U10038 (N_10038,N_9796,N_8722);
nand U10039 (N_10039,N_7660,N_9810);
or U10040 (N_10040,N_8901,N_7708);
nand U10041 (N_10041,N_8418,N_8013);
and U10042 (N_10042,N_9467,N_8342);
nor U10043 (N_10043,N_9815,N_8097);
xnor U10044 (N_10044,N_9996,N_8862);
nand U10045 (N_10045,N_7533,N_9015);
nor U10046 (N_10046,N_8952,N_7870);
and U10047 (N_10047,N_8646,N_8548);
and U10048 (N_10048,N_7566,N_9708);
or U10049 (N_10049,N_8698,N_9668);
or U10050 (N_10050,N_9979,N_9778);
xor U10051 (N_10051,N_9640,N_8824);
xor U10052 (N_10052,N_8743,N_9775);
nor U10053 (N_10053,N_9530,N_7586);
nand U10054 (N_10054,N_8444,N_9085);
nor U10055 (N_10055,N_7718,N_8663);
nor U10056 (N_10056,N_9406,N_9637);
xor U10057 (N_10057,N_8832,N_8536);
nor U10058 (N_10058,N_9629,N_8105);
and U10059 (N_10059,N_8938,N_8221);
nor U10060 (N_10060,N_8488,N_8461);
or U10061 (N_10061,N_8482,N_8742);
or U10062 (N_10062,N_7679,N_7832);
or U10063 (N_10063,N_8472,N_8349);
nor U10064 (N_10064,N_9502,N_9762);
or U10065 (N_10065,N_9728,N_9900);
or U10066 (N_10066,N_8785,N_8400);
and U10067 (N_10067,N_9589,N_7827);
or U10068 (N_10068,N_9188,N_8168);
or U10069 (N_10069,N_8193,N_9392);
xnor U10070 (N_10070,N_9352,N_8948);
and U10071 (N_10071,N_9332,N_9365);
and U10072 (N_10072,N_8334,N_9388);
nand U10073 (N_10073,N_7503,N_8129);
xor U10074 (N_10074,N_7535,N_8109);
or U10075 (N_10075,N_8328,N_7743);
xnor U10076 (N_10076,N_8509,N_8960);
nor U10077 (N_10077,N_9586,N_7671);
or U10078 (N_10078,N_7585,N_9145);
nand U10079 (N_10079,N_9108,N_9564);
nor U10080 (N_10080,N_9315,N_8464);
or U10081 (N_10081,N_9879,N_7784);
nand U10082 (N_10082,N_9910,N_9643);
or U10083 (N_10083,N_9569,N_9274);
nand U10084 (N_10084,N_8558,N_7849);
or U10085 (N_10085,N_9638,N_9197);
and U10086 (N_10086,N_9349,N_7696);
or U10087 (N_10087,N_8187,N_9581);
nand U10088 (N_10088,N_8493,N_8805);
nand U10089 (N_10089,N_8374,N_8411);
nor U10090 (N_10090,N_8563,N_9020);
and U10091 (N_10091,N_8906,N_7959);
xor U10092 (N_10092,N_9237,N_7903);
or U10093 (N_10093,N_9304,N_8043);
xor U10094 (N_10094,N_8589,N_7665);
nand U10095 (N_10095,N_8401,N_9848);
nor U10096 (N_10096,N_9580,N_8882);
nor U10097 (N_10097,N_9617,N_7511);
nand U10098 (N_10098,N_9273,N_9149);
nand U10099 (N_10099,N_8837,N_8269);
and U10100 (N_10100,N_9945,N_9947);
and U10101 (N_10101,N_9831,N_7859);
xnor U10102 (N_10102,N_8749,N_8059);
and U10103 (N_10103,N_9263,N_9307);
xnor U10104 (N_10104,N_8503,N_7865);
xor U10105 (N_10105,N_9094,N_7582);
xnor U10106 (N_10106,N_7605,N_7962);
xor U10107 (N_10107,N_8531,N_9380);
nand U10108 (N_10108,N_9679,N_8593);
nand U10109 (N_10109,N_9173,N_9376);
xor U10110 (N_10110,N_7615,N_8552);
and U10111 (N_10111,N_7620,N_8875);
or U10112 (N_10112,N_9892,N_7922);
xnor U10113 (N_10113,N_7633,N_9299);
or U10114 (N_10114,N_7873,N_9251);
nor U10115 (N_10115,N_9322,N_9393);
nand U10116 (N_10116,N_7617,N_9037);
xnor U10117 (N_10117,N_8085,N_8997);
xor U10118 (N_10118,N_8029,N_9847);
or U10119 (N_10119,N_9485,N_7795);
or U10120 (N_10120,N_8460,N_9191);
or U10121 (N_10121,N_8855,N_8904);
nor U10122 (N_10122,N_9285,N_8336);
or U10123 (N_10123,N_9827,N_8953);
and U10124 (N_10124,N_8793,N_8712);
or U10125 (N_10125,N_9805,N_9861);
nand U10126 (N_10126,N_9435,N_8188);
nor U10127 (N_10127,N_9972,N_9545);
or U10128 (N_10128,N_9182,N_9938);
xor U10129 (N_10129,N_8362,N_9175);
nand U10130 (N_10130,N_8836,N_9860);
nand U10131 (N_10131,N_8266,N_8280);
xor U10132 (N_10132,N_8725,N_8512);
nand U10133 (N_10133,N_8919,N_9087);
or U10134 (N_10134,N_8327,N_9849);
xnor U10135 (N_10135,N_8494,N_9992);
nand U10136 (N_10136,N_8641,N_9676);
or U10137 (N_10137,N_8684,N_9325);
and U10138 (N_10138,N_7687,N_8827);
nand U10139 (N_10139,N_9309,N_8404);
nor U10140 (N_10140,N_7993,N_9624);
nor U10141 (N_10141,N_9417,N_9187);
xor U10142 (N_10142,N_9231,N_9014);
or U10143 (N_10143,N_8647,N_7532);
xor U10144 (N_10144,N_8412,N_8858);
nand U10145 (N_10145,N_7531,N_9368);
nor U10146 (N_10146,N_9326,N_8640);
or U10147 (N_10147,N_8380,N_8087);
nand U10148 (N_10148,N_8961,N_9528);
and U10149 (N_10149,N_7830,N_9543);
nand U10150 (N_10150,N_8240,N_9704);
nor U10151 (N_10151,N_7926,N_9659);
or U10152 (N_10152,N_7732,N_9712);
nand U10153 (N_10153,N_9006,N_9803);
nand U10154 (N_10154,N_8958,N_9294);
and U10155 (N_10155,N_7952,N_8477);
or U10156 (N_10156,N_9601,N_8654);
xnor U10157 (N_10157,N_7597,N_7602);
or U10158 (N_10158,N_8309,N_9412);
xor U10159 (N_10159,N_9963,N_8406);
nand U10160 (N_10160,N_8682,N_7756);
xnor U10161 (N_10161,N_8851,N_9786);
and U10162 (N_10162,N_8185,N_8293);
nand U10163 (N_10163,N_7909,N_8247);
and U10164 (N_10164,N_9698,N_7982);
and U10165 (N_10165,N_8983,N_9126);
xnor U10166 (N_10166,N_8826,N_8979);
and U10167 (N_10167,N_7751,N_8448);
and U10168 (N_10168,N_8976,N_8772);
nand U10169 (N_10169,N_8471,N_7860);
nor U10170 (N_10170,N_8726,N_8700);
and U10171 (N_10171,N_9573,N_7885);
xnor U10172 (N_10172,N_9469,N_9714);
xor U10173 (N_10173,N_9374,N_8172);
nand U10174 (N_10174,N_8922,N_8326);
or U10175 (N_10175,N_9940,N_8614);
nor U10176 (N_10176,N_7757,N_9804);
or U10177 (N_10177,N_8816,N_8994);
and U10178 (N_10178,N_8756,N_9907);
or U10179 (N_10179,N_9010,N_7824);
and U10180 (N_10180,N_8203,N_8223);
or U10181 (N_10181,N_9092,N_8182);
nor U10182 (N_10182,N_8996,N_9766);
nor U10183 (N_10183,N_8718,N_7558);
or U10184 (N_10184,N_7645,N_8288);
or U10185 (N_10185,N_7825,N_9451);
xor U10186 (N_10186,N_8658,N_9250);
and U10187 (N_10187,N_8524,N_9228);
nand U10188 (N_10188,N_8605,N_7848);
and U10189 (N_10189,N_7628,N_9410);
nor U10190 (N_10190,N_8877,N_8932);
xor U10191 (N_10191,N_9257,N_8272);
or U10192 (N_10192,N_7923,N_8450);
or U10193 (N_10193,N_9444,N_8764);
and U10194 (N_10194,N_9635,N_9032);
nand U10195 (N_10195,N_8693,N_7596);
nand U10196 (N_10196,N_9781,N_8110);
nand U10197 (N_10197,N_8335,N_9355);
nor U10198 (N_10198,N_8166,N_9503);
or U10199 (N_10199,N_9636,N_8703);
and U10200 (N_10200,N_7507,N_8368);
nand U10201 (N_10201,N_8316,N_8856);
and U10202 (N_10202,N_8917,N_8214);
nand U10203 (N_10203,N_9887,N_7933);
nor U10204 (N_10204,N_8408,N_8470);
or U10205 (N_10205,N_9955,N_9578);
xor U10206 (N_10206,N_9324,N_7540);
nand U10207 (N_10207,N_7599,N_8145);
xor U10208 (N_10208,N_9480,N_7955);
xor U10209 (N_10209,N_8005,N_8798);
nor U10210 (N_10210,N_9153,N_8220);
xor U10211 (N_10211,N_8091,N_9612);
xnor U10212 (N_10212,N_7935,N_9007);
or U10213 (N_10213,N_8817,N_9870);
and U10214 (N_10214,N_8530,N_8128);
xor U10215 (N_10215,N_9536,N_9905);
xnor U10216 (N_10216,N_7838,N_8332);
xnor U10217 (N_10217,N_8676,N_9050);
or U10218 (N_10218,N_9138,N_9873);
nand U10219 (N_10219,N_9575,N_8545);
nand U10220 (N_10220,N_7747,N_8179);
nor U10221 (N_10221,N_9592,N_8839);
nand U10222 (N_10222,N_9248,N_9419);
nor U10223 (N_10223,N_8681,N_7774);
and U10224 (N_10224,N_9524,N_8748);
xnor U10225 (N_10225,N_8982,N_8517);
xor U10226 (N_10226,N_9764,N_8161);
and U10227 (N_10227,N_8197,N_9943);
nor U10228 (N_10228,N_9398,N_9067);
nand U10229 (N_10229,N_7501,N_8273);
and U10230 (N_10230,N_8510,N_9912);
nand U10231 (N_10231,N_8040,N_7562);
nor U10232 (N_10232,N_7733,N_9991);
or U10233 (N_10233,N_8403,N_9544);
nor U10234 (N_10234,N_9837,N_8802);
or U10235 (N_10235,N_9041,N_7777);
and U10236 (N_10236,N_9794,N_8148);
xnor U10237 (N_10237,N_8532,N_9090);
nor U10238 (N_10238,N_8644,N_7871);
nand U10239 (N_10239,N_9328,N_8351);
and U10240 (N_10240,N_9724,N_8719);
nand U10241 (N_10241,N_7919,N_8064);
or U10242 (N_10242,N_9771,N_9481);
nand U10243 (N_10243,N_9995,N_8439);
or U10244 (N_10244,N_9272,N_8965);
nor U10245 (N_10245,N_7664,N_8370);
nand U10246 (N_10246,N_7702,N_8434);
xnor U10247 (N_10247,N_7810,N_8706);
nand U10248 (N_10248,N_9993,N_9261);
nor U10249 (N_10249,N_8883,N_8320);
and U10250 (N_10250,N_9715,N_7775);
nor U10251 (N_10251,N_9292,N_9628);
or U10252 (N_10252,N_9282,N_9474);
nor U10253 (N_10253,N_8705,N_9243);
nor U10254 (N_10254,N_9401,N_9987);
nor U10255 (N_10255,N_9854,N_9664);
xnor U10256 (N_10256,N_7934,N_8709);
nor U10257 (N_10257,N_7731,N_7816);
nor U10258 (N_10258,N_8050,N_7555);
xnor U10259 (N_10259,N_8767,N_9049);
and U10260 (N_10260,N_9484,N_9779);
and U10261 (N_10261,N_8198,N_8590);
nor U10262 (N_10262,N_8300,N_9852);
nand U10263 (N_10263,N_7793,N_8632);
nand U10264 (N_10264,N_9427,N_8118);
xnor U10265 (N_10265,N_8101,N_8970);
xnor U10266 (N_10266,N_7630,N_9678);
nor U10267 (N_10267,N_8468,N_8800);
xor U10268 (N_10268,N_8123,N_8549);
nand U10269 (N_10269,N_8356,N_9023);
nor U10270 (N_10270,N_8484,N_8670);
and U10271 (N_10271,N_8021,N_9168);
xnor U10272 (N_10272,N_7549,N_7670);
xor U10273 (N_10273,N_7697,N_9776);
nand U10274 (N_10274,N_9622,N_8609);
and U10275 (N_10275,N_9447,N_8860);
xor U10276 (N_10276,N_8313,N_7791);
xor U10277 (N_10277,N_7735,N_7945);
or U10278 (N_10278,N_9224,N_8803);
nand U10279 (N_10279,N_7704,N_7768);
nand U10280 (N_10280,N_8207,N_9855);
nor U10281 (N_10281,N_7509,N_9232);
or U10282 (N_10282,N_8151,N_8141);
and U10283 (N_10283,N_7724,N_8556);
xor U10284 (N_10284,N_8942,N_9496);
xnor U10285 (N_10285,N_9179,N_7802);
and U10286 (N_10286,N_9650,N_8416);
nand U10287 (N_10287,N_9933,N_8135);
nor U10288 (N_10288,N_9161,N_8292);
nor U10289 (N_10289,N_9117,N_7676);
nand U10290 (N_10290,N_9789,N_9075);
nor U10291 (N_10291,N_8539,N_8498);
xor U10292 (N_10292,N_8916,N_8736);
nand U10293 (N_10293,N_7713,N_7598);
and U10294 (N_10294,N_9978,N_8271);
xor U10295 (N_10295,N_7764,N_8980);
nand U10296 (N_10296,N_8016,N_9761);
nor U10297 (N_10297,N_9162,N_8047);
nor U10298 (N_10298,N_9048,N_8191);
nor U10299 (N_10299,N_8012,N_8208);
nand U10300 (N_10300,N_9780,N_7884);
nand U10301 (N_10301,N_8741,N_9695);
or U10302 (N_10302,N_9974,N_9465);
or U10303 (N_10303,N_9362,N_8576);
and U10304 (N_10304,N_8603,N_9823);
and U10305 (N_10305,N_8098,N_8004);
and U10306 (N_10306,N_8250,N_9448);
nand U10307 (N_10307,N_8463,N_9747);
or U10308 (N_10308,N_9529,N_8788);
nand U10309 (N_10309,N_8631,N_9363);
xnor U10310 (N_10310,N_8410,N_9036);
and U10311 (N_10311,N_9450,N_9449);
xnor U10312 (N_10312,N_8571,N_9763);
xor U10313 (N_10313,N_8371,N_8655);
xnor U10314 (N_10314,N_7877,N_8111);
and U10315 (N_10315,N_9455,N_8325);
xor U10316 (N_10316,N_9167,N_7556);
xor U10317 (N_10317,N_9491,N_8194);
or U10318 (N_10318,N_7646,N_8030);
and U10319 (N_10319,N_9262,N_9562);
nand U10320 (N_10320,N_9206,N_9183);
xnor U10321 (N_10321,N_7753,N_7961);
and U10322 (N_10322,N_9785,N_7744);
or U10323 (N_10323,N_7680,N_7709);
nand U10324 (N_10324,N_9812,N_8879);
and U10325 (N_10325,N_8481,N_7843);
nor U10326 (N_10326,N_9512,N_7991);
nand U10327 (N_10327,N_9745,N_8398);
nand U10328 (N_10328,N_7560,N_8528);
xor U10329 (N_10329,N_7576,N_8001);
xor U10330 (N_10330,N_7856,N_8205);
and U10331 (N_10331,N_9792,N_9115);
nor U10332 (N_10332,N_8390,N_9002);
nand U10333 (N_10333,N_9160,N_9341);
nand U10334 (N_10334,N_8964,N_8913);
nor U10335 (N_10335,N_9645,N_8865);
nand U10336 (N_10336,N_8947,N_9639);
or U10337 (N_10337,N_8559,N_9354);
nand U10338 (N_10338,N_8483,N_8925);
nor U10339 (N_10339,N_7739,N_7797);
nor U10340 (N_10340,N_7817,N_9915);
or U10341 (N_10341,N_7506,N_9884);
and U10342 (N_10342,N_8515,N_9705);
nand U10343 (N_10343,N_8588,N_7631);
and U10344 (N_10344,N_9220,N_9195);
nand U10345 (N_10345,N_9056,N_8765);
nand U10346 (N_10346,N_9260,N_9641);
nand U10347 (N_10347,N_8264,N_8635);
xor U10348 (N_10348,N_7545,N_9603);
or U10349 (N_10349,N_8209,N_8583);
or U10350 (N_10350,N_9219,N_9557);
nand U10351 (N_10351,N_9648,N_9256);
nand U10352 (N_10352,N_8734,N_8167);
or U10353 (N_10353,N_8661,N_7639);
xnor U10354 (N_10354,N_8625,N_9735);
nand U10355 (N_10355,N_7692,N_8155);
xor U10356 (N_10356,N_7570,N_8677);
and U10357 (N_10357,N_9136,N_7745);
or U10358 (N_10358,N_9523,N_7834);
and U10359 (N_10359,N_8228,N_7572);
or U10360 (N_10360,N_8139,N_9507);
and U10361 (N_10361,N_8830,N_9553);
xnor U10362 (N_10362,N_7904,N_7520);
nand U10363 (N_10363,N_8808,N_7828);
nor U10364 (N_10364,N_7728,N_9180);
xnor U10365 (N_10365,N_9356,N_8720);
or U10366 (N_10366,N_7901,N_9956);
nand U10367 (N_10367,N_9495,N_8089);
nor U10368 (N_10368,N_8317,N_8233);
nand U10369 (N_10369,N_9426,N_8386);
or U10370 (N_10370,N_9443,N_9962);
nor U10371 (N_10371,N_9247,N_9430);
nor U10372 (N_10372,N_9017,N_8842);
or U10373 (N_10373,N_9806,N_9906);
and U10374 (N_10374,N_8971,N_8954);
nor U10375 (N_10375,N_7693,N_9760);
xnor U10376 (N_10376,N_8537,N_8610);
or U10377 (N_10377,N_7968,N_7893);
nor U10378 (N_10378,N_8683,N_8415);
nor U10379 (N_10379,N_8792,N_8164);
and U10380 (N_10380,N_9208,N_8294);
xor U10381 (N_10381,N_8224,N_9446);
xor U10382 (N_10382,N_9868,N_8660);
or U10383 (N_10383,N_7761,N_7730);
and U10384 (N_10384,N_9865,N_9080);
xnor U10385 (N_10385,N_9240,N_9694);
or U10386 (N_10386,N_7988,N_9620);
xor U10387 (N_10387,N_7841,N_7557);
or U10388 (N_10388,N_8737,N_9391);
nand U10389 (N_10389,N_9672,N_8083);
and U10390 (N_10390,N_9044,N_8870);
nor U10391 (N_10391,N_9801,N_9721);
nand U10392 (N_10392,N_9984,N_9074);
and U10393 (N_10393,N_9881,N_9336);
or U10394 (N_10394,N_8146,N_8192);
xor U10395 (N_10395,N_9515,N_7519);
nor U10396 (N_10396,N_9774,N_8518);
nand U10397 (N_10397,N_8505,N_8405);
nand U10398 (N_10398,N_9600,N_7609);
and U10399 (N_10399,N_9464,N_9318);
nor U10400 (N_10400,N_9245,N_9730);
nand U10401 (N_10401,N_9314,N_8715);
and U10402 (N_10402,N_8926,N_9917);
and U10403 (N_10403,N_9101,N_8159);
or U10404 (N_10404,N_9560,N_8375);
and U10405 (N_10405,N_7648,N_8200);
or U10406 (N_10406,N_9880,N_7771);
and U10407 (N_10407,N_8673,N_7786);
or U10408 (N_10408,N_9510,N_9019);
or U10409 (N_10409,N_8449,N_7547);
xor U10410 (N_10410,N_8669,N_7880);
nand U10411 (N_10411,N_8747,N_9066);
nor U10412 (N_10412,N_9893,N_9867);
and U10413 (N_10413,N_9539,N_9896);
nand U10414 (N_10414,N_9949,N_8373);
or U10415 (N_10415,N_8818,N_9919);
and U10416 (N_10416,N_8854,N_9308);
nand U10417 (N_10417,N_9086,N_8383);
or U10418 (N_10418,N_9331,N_7887);
nand U10419 (N_10419,N_9113,N_8131);
nor U10420 (N_10420,N_9063,N_7882);
xor U10421 (N_10421,N_9859,N_9651);
xor U10422 (N_10422,N_9259,N_8529);
or U10423 (N_10423,N_8107,N_9018);
nand U10424 (N_10424,N_8773,N_9671);
and U10425 (N_10425,N_8033,N_9429);
nand U10426 (N_10426,N_8442,N_9817);
or U10427 (N_10427,N_9720,N_8768);
nor U10428 (N_10428,N_9016,N_9627);
nand U10429 (N_10429,N_7649,N_7623);
and U10430 (N_10430,N_9830,N_9744);
or U10431 (N_10431,N_9926,N_7833);
and U10432 (N_10432,N_7826,N_9967);
nor U10433 (N_10433,N_8621,N_8597);
nor U10434 (N_10434,N_8358,N_8829);
nor U10435 (N_10435,N_7726,N_7979);
xnor U10436 (N_10436,N_9696,N_8685);
nand U10437 (N_10437,N_8093,N_9784);
and U10438 (N_10438,N_8133,N_7782);
nor U10439 (N_10439,N_9439,N_9874);
nand U10440 (N_10440,N_8438,N_8710);
nor U10441 (N_10441,N_7932,N_9039);
xnor U10442 (N_10442,N_7818,N_7569);
or U10443 (N_10443,N_9768,N_8094);
nand U10444 (N_10444,N_8459,N_7790);
and U10445 (N_10445,N_7965,N_9959);
nand U10446 (N_10446,N_9303,N_9546);
nor U10447 (N_10447,N_9091,N_8868);
xor U10448 (N_10448,N_8846,N_8986);
and U10449 (N_10449,N_9819,N_7766);
and U10450 (N_10450,N_9667,N_8170);
nor U10451 (N_10451,N_9857,N_7722);
nand U10452 (N_10452,N_8453,N_9691);
xnor U10453 (N_10453,N_8216,N_7647);
nand U10454 (N_10454,N_7502,N_8389);
nor U10455 (N_10455,N_8859,N_9205);
xnor U10456 (N_10456,N_8372,N_9997);
nand U10457 (N_10457,N_8023,N_9004);
and U10458 (N_10458,N_8217,N_9833);
xnor U10459 (N_10459,N_8786,N_9828);
xor U10460 (N_10460,N_8507,N_8874);
and U10461 (N_10461,N_7537,N_9681);
xor U10462 (N_10462,N_9405,N_9283);
xor U10463 (N_10463,N_8648,N_9150);
and U10464 (N_10464,N_7546,N_7568);
nand U10465 (N_10465,N_7673,N_8259);
nor U10466 (N_10466,N_7593,N_9550);
xnor U10467 (N_10467,N_9965,N_8045);
nor U10468 (N_10468,N_7505,N_8254);
or U10469 (N_10469,N_9269,N_9618);
xnor U10470 (N_10470,N_8345,N_9661);
xnor U10471 (N_10471,N_8944,N_7845);
nor U10472 (N_10472,N_8144,N_9824);
or U10473 (N_10473,N_9061,N_8027);
and U10474 (N_10474,N_9098,N_8431);
or U10475 (N_10475,N_8253,N_8809);
and U10476 (N_10476,N_7658,N_9716);
and U10477 (N_10477,N_7588,N_8981);
nand U10478 (N_10478,N_9932,N_9252);
and U10479 (N_10479,N_7940,N_8935);
or U10480 (N_10480,N_9311,N_9754);
and U10481 (N_10481,N_8766,N_9428);
or U10482 (N_10482,N_7796,N_9505);
and U10483 (N_10483,N_8797,N_8567);
and U10484 (N_10484,N_9533,N_9255);
nor U10485 (N_10485,N_7986,N_8791);
nor U10486 (N_10486,N_9982,N_9000);
or U10487 (N_10487,N_8227,N_9918);
xnor U10488 (N_10488,N_9317,N_7953);
or U10489 (N_10489,N_8657,N_9741);
nor U10490 (N_10490,N_9408,N_8031);
and U10491 (N_10491,N_8279,N_7840);
xnor U10492 (N_10492,N_9369,N_8491);
and U10493 (N_10493,N_9165,N_7883);
or U10494 (N_10494,N_9946,N_7711);
or U10495 (N_10495,N_9367,N_9171);
xor U10496 (N_10496,N_9937,N_9390);
nor U10497 (N_10497,N_8361,N_8562);
and U10498 (N_10498,N_8478,N_8365);
nor U10499 (N_10499,N_9807,N_9029);
nor U10500 (N_10500,N_8616,N_7976);
xor U10501 (N_10501,N_9777,N_8092);
nor U10502 (N_10502,N_9024,N_9399);
and U10503 (N_10503,N_8572,N_8758);
nor U10504 (N_10504,N_9218,N_8624);
nor U10505 (N_10505,N_7815,N_9330);
xnor U10506 (N_10506,N_7652,N_8946);
nor U10507 (N_10507,N_8759,N_9683);
or U10508 (N_10508,N_7651,N_8987);
or U10509 (N_10509,N_9504,N_8469);
nand U10510 (N_10510,N_8880,N_8540);
nor U10511 (N_10511,N_8473,N_9460);
and U10512 (N_10512,N_9499,N_9462);
nor U10513 (N_10513,N_8399,N_9366);
nand U10514 (N_10514,N_9611,N_7574);
or U10515 (N_10515,N_8154,N_8462);
xnor U10516 (N_10516,N_9675,N_8520);
nor U10517 (N_10517,N_8521,N_8283);
and U10518 (N_10518,N_8267,N_9276);
and U10519 (N_10519,N_7754,N_8619);
or U10520 (N_10520,N_9229,N_7927);
or U10521 (N_10521,N_9470,N_8969);
nand U10522 (N_10522,N_9003,N_8312);
nor U10523 (N_10523,N_9800,N_8513);
xor U10524 (N_10524,N_9477,N_9878);
xor U10525 (N_10525,N_9835,N_8395);
nand U10526 (N_10526,N_9073,N_8420);
xor U10527 (N_10527,N_7994,N_9687);
and U10528 (N_10528,N_9904,N_9348);
and U10529 (N_10529,N_8433,N_9630);
nor U10530 (N_10530,N_9966,N_7734);
or U10531 (N_10531,N_9387,N_8781);
nand U10532 (N_10532,N_9337,N_8343);
nor U10533 (N_10533,N_9452,N_9270);
and U10534 (N_10534,N_8291,N_9414);
or U10535 (N_10535,N_8062,N_8081);
nor U10536 (N_10536,N_9522,N_8303);
nor U10537 (N_10537,N_8841,N_9194);
and U10538 (N_10538,N_9596,N_8263);
or U10539 (N_10539,N_9432,N_7769);
xnor U10540 (N_10540,N_8740,N_9454);
nor U10541 (N_10541,N_8789,N_7948);
or U10542 (N_10542,N_9323,N_9456);
and U10543 (N_10543,N_8183,N_9159);
nor U10544 (N_10544,N_9594,N_8028);
nand U10545 (N_10545,N_9541,N_9970);
or U10546 (N_10546,N_9302,N_8555);
xor U10547 (N_10547,N_8397,N_9345);
xnor U10548 (N_10548,N_9404,N_8894);
and U10549 (N_10549,N_7667,N_8950);
and U10550 (N_10550,N_9459,N_7767);
nor U10551 (N_10551,N_8311,N_8330);
nor U10552 (N_10552,N_8840,N_7536);
and U10553 (N_10553,N_8249,N_7974);
or U10554 (N_10554,N_8451,N_7780);
nor U10555 (N_10555,N_8923,N_9588);
xnor U10556 (N_10556,N_7892,N_7954);
xor U10557 (N_10557,N_9631,N_7799);
xor U10558 (N_10558,N_7595,N_7740);
xnor U10559 (N_10559,N_8366,N_8285);
or U10560 (N_10560,N_8231,N_8968);
nor U10561 (N_10561,N_9656,N_8955);
nand U10562 (N_10562,N_9953,N_9339);
nor U10563 (N_10563,N_9210,N_8308);
nor U10564 (N_10564,N_8519,N_8959);
xnor U10565 (N_10565,N_9494,N_9146);
nor U10566 (N_10566,N_9277,N_8881);
nor U10567 (N_10567,N_8871,N_9384);
xnor U10568 (N_10568,N_7842,N_9185);
nand U10569 (N_10569,N_8298,N_8173);
or U10570 (N_10570,N_8591,N_8122);
xor U10571 (N_10571,N_9954,N_7785);
or U10572 (N_10572,N_7902,N_8833);
or U10573 (N_10573,N_8222,N_7748);
or U10574 (N_10574,N_9511,N_9990);
xor U10575 (N_10575,N_9346,N_9060);
and U10576 (N_10576,N_8242,N_8359);
and U10577 (N_10577,N_8260,N_9296);
nor U10578 (N_10578,N_8268,N_7746);
nor U10579 (N_10579,N_7858,N_9425);
xor U10580 (N_10580,N_8000,N_8845);
or U10581 (N_10581,N_9209,N_8704);
nor U10582 (N_10582,N_9119,N_7717);
nor U10583 (N_10583,N_9765,N_8810);
nor U10584 (N_10584,N_8323,N_7690);
nor U10585 (N_10585,N_8977,N_8566);
nor U10586 (N_10586,N_8126,N_9709);
and U10587 (N_10587,N_8666,N_7973);
or U10588 (N_10588,N_9808,N_9466);
or U10589 (N_10589,N_8665,N_9062);
or U10590 (N_10590,N_7943,N_8367);
nand U10591 (N_10591,N_9012,N_8723);
nand U10592 (N_10592,N_8495,N_8834);
and U10593 (N_10593,N_7925,N_9525);
and U10594 (N_10594,N_8504,N_9021);
and U10595 (N_10595,N_8595,N_9623);
or U10596 (N_10596,N_9851,N_8413);
and U10597 (N_10597,N_7636,N_7552);
nor U10598 (N_10598,N_8314,N_7992);
nor U10599 (N_10599,N_8344,N_9551);
or U10600 (N_10600,N_9028,N_7705);
nand U10601 (N_10601,N_8746,N_9516);
nor U10602 (N_10602,N_9244,N_7930);
or U10603 (N_10603,N_9071,N_8007);
and U10604 (N_10604,N_7750,N_7759);
xor U10605 (N_10605,N_8113,N_8627);
or U10606 (N_10606,N_8825,N_8812);
xnor U10607 (N_10607,N_8057,N_9184);
and U10608 (N_10608,N_9373,N_8653);
or U10609 (N_10609,N_9207,N_8811);
nand U10610 (N_10610,N_7737,N_8891);
xor U10611 (N_10611,N_7663,N_7872);
nor U10612 (N_10612,N_8423,N_9396);
and U10613 (N_10613,N_9999,N_9597);
nor U10614 (N_10614,N_9157,N_7527);
xor U10615 (N_10615,N_8578,N_9181);
and U10616 (N_10616,N_8219,N_8455);
or U10617 (N_10617,N_9532,N_9359);
or U10618 (N_10618,N_8754,N_8490);
or U10619 (N_10619,N_8750,N_8662);
or U10620 (N_10620,N_8634,N_7894);
nand U10621 (N_10621,N_9193,N_8522);
and U10622 (N_10622,N_8777,N_7950);
or U10623 (N_10623,N_9124,N_7541);
and U10624 (N_10624,N_9027,N_8931);
xnor U10625 (N_10625,N_7508,N_8496);
xor U10626 (N_10626,N_7762,N_7822);
or U10627 (N_10627,N_8190,N_8905);
or U10628 (N_10628,N_7851,N_8287);
nor U10629 (N_10629,N_8069,N_8246);
and U10630 (N_10630,N_9079,N_7675);
xnor U10631 (N_10631,N_7804,N_9114);
nor U10632 (N_10632,N_7621,N_9400);
and U10633 (N_10633,N_9732,N_9135);
nor U10634 (N_10634,N_8127,N_7891);
nor U10635 (N_10635,N_9832,N_9929);
nand U10636 (N_10636,N_7551,N_7758);
and U10637 (N_10637,N_9201,N_9291);
and U10638 (N_10638,N_7707,N_9344);
or U10639 (N_10639,N_8206,N_9409);
or U10640 (N_10640,N_9750,N_9674);
or U10641 (N_10641,N_9570,N_8058);
nand U10642 (N_10642,N_8229,N_9547);
xnor U10643 (N_10643,N_8714,N_8036);
or U10644 (N_10644,N_7811,N_9253);
or U10645 (N_10645,N_9100,N_8675);
and U10646 (N_10646,N_9985,N_7504);
xor U10647 (N_10647,N_9839,N_8599);
and U10648 (N_10648,N_7912,N_7669);
or U10649 (N_10649,N_8432,N_8077);
nand U10650 (N_10650,N_8533,N_9418);
and U10651 (N_10651,N_9519,N_7914);
and U10652 (N_10652,N_8204,N_9139);
xnor U10653 (N_10653,N_9438,N_9131);
nor U10654 (N_10654,N_8236,N_9152);
xor U10655 (N_10655,N_8581,N_9176);
or U10656 (N_10656,N_8301,N_9733);
or U10657 (N_10657,N_9351,N_8119);
or U10658 (N_10658,N_9305,N_7755);
nand U10659 (N_10659,N_8071,N_9127);
and U10660 (N_10660,N_7798,N_8770);
nand U10661 (N_10661,N_9531,N_9293);
or U10662 (N_10662,N_7829,N_9973);
nor U10663 (N_10663,N_9431,N_9163);
and U10664 (N_10664,N_9614,N_9773);
nor U10665 (N_10665,N_8526,N_8352);
or U10666 (N_10666,N_9442,N_8850);
nand U10667 (N_10667,N_7938,N_8422);
or U10668 (N_10668,N_9706,N_8447);
or U10669 (N_10669,N_8617,N_8903);
nor U10670 (N_10670,N_9701,N_8339);
nand U10671 (N_10671,N_8396,N_8985);
xor U10672 (N_10672,N_9920,N_9089);
and U10673 (N_10673,N_9670,N_9540);
or U10674 (N_10674,N_8620,N_8304);
and U10675 (N_10675,N_9548,N_7844);
or U10676 (N_10676,N_9613,N_7688);
and U10677 (N_10677,N_8121,N_8643);
xor U10678 (N_10678,N_8893,N_9876);
nand U10679 (N_10679,N_8108,N_8180);
and U10680 (N_10680,N_8394,N_8427);
and U10681 (N_10681,N_7969,N_9555);
or U10682 (N_10682,N_8783,N_8456);
nor U10683 (N_10683,N_8594,N_9011);
and U10684 (N_10684,N_9838,N_8899);
nor U10685 (N_10685,N_9122,N_8708);
nand U10686 (N_10686,N_8943,N_9105);
nor U10687 (N_10687,N_7853,N_8014);
xnor U10688 (N_10688,N_8888,N_8322);
xnor U10689 (N_10689,N_9068,N_8244);
nor U10690 (N_10690,N_8711,N_9818);
and U10691 (N_10691,N_7998,N_9064);
and U10692 (N_10692,N_8608,N_7852);
or U10693 (N_10693,N_9213,N_8186);
xor U10694 (N_10694,N_9654,N_8385);
nor U10695 (N_10695,N_7522,N_9321);
nand U10696 (N_10696,N_8611,N_9961);
xnor U10697 (N_10697,N_9595,N_8633);
xnor U10698 (N_10698,N_9520,N_8918);
and U10699 (N_10699,N_9151,N_9440);
nor U10700 (N_10700,N_7876,N_9289);
or U10701 (N_10701,N_7581,N_8909);
nor U10702 (N_10702,N_7895,N_9802);
nand U10703 (N_10703,N_8176,N_7685);
nor U10704 (N_10704,N_9342,N_8066);
xor U10705 (N_10705,N_7863,N_8636);
nand U10706 (N_10706,N_8598,N_8290);
nor U10707 (N_10707,N_8914,N_9758);
and U10708 (N_10708,N_9238,N_8602);
nor U10709 (N_10709,N_9649,N_7888);
xor U10710 (N_10710,N_8348,N_8835);
and U10711 (N_10711,N_8941,N_8790);
or U10712 (N_10712,N_9606,N_8707);
xor U10713 (N_10713,N_8100,N_8138);
and U10714 (N_10714,N_8051,N_9501);
nor U10715 (N_10715,N_8664,N_9891);
xnor U10716 (N_10716,N_7770,N_9096);
nor U10717 (N_10717,N_9692,N_9316);
xor U10718 (N_10718,N_7975,N_9983);
and U10719 (N_10719,N_9572,N_9902);
nor U10720 (N_10720,N_8134,N_9254);
or U10721 (N_10721,N_8652,N_8849);
xnor U10722 (N_10722,N_8152,N_7600);
xnor U10723 (N_10723,N_7626,N_9923);
xnor U10724 (N_10724,N_8044,N_8695);
nand U10725 (N_10725,N_8574,N_9725);
or U10726 (N_10726,N_8090,N_9759);
or U10727 (N_10727,N_7951,N_9358);
and U10728 (N_10728,N_9610,N_9890);
xor U10729 (N_10729,N_9482,N_7999);
nand U10730 (N_10730,N_7963,N_8592);
nor U10731 (N_10731,N_9952,N_8838);
nor U10732 (N_10732,N_8174,N_8995);
nor U10733 (N_10733,N_9106,N_8295);
nand U10734 (N_10734,N_7957,N_8920);
or U10735 (N_10735,N_9249,N_9748);
nand U10736 (N_10736,N_9155,N_8639);
nand U10737 (N_10737,N_9719,N_8506);
nor U10738 (N_10738,N_8940,N_7529);
or U10739 (N_10739,N_8466,N_8315);
and U10740 (N_10740,N_9756,N_7783);
nor U10741 (N_10741,N_8177,N_9436);
nor U10742 (N_10742,N_8690,N_7812);
xnor U10743 (N_10743,N_9040,N_9568);
nand U10744 (N_10744,N_8116,N_7559);
xnor U10745 (N_10745,N_8347,N_9927);
xor U10746 (N_10746,N_8511,N_8171);
or U10747 (N_10747,N_8237,N_8689);
nor U10748 (N_10748,N_8041,N_9140);
xor U10749 (N_10749,N_8243,N_9403);
nand U10750 (N_10750,N_9058,N_9312);
nand U10751 (N_10751,N_9770,N_7879);
or U10752 (N_10752,N_9083,N_9055);
or U10753 (N_10753,N_7654,N_8329);
or U10754 (N_10754,N_8132,N_9492);
and U10755 (N_10755,N_8252,N_7897);
or U10756 (N_10756,N_8003,N_9264);
nand U10757 (N_10757,N_9141,N_9825);
nand U10758 (N_10758,N_8212,N_7805);
xnor U10759 (N_10759,N_8613,N_9582);
nand U10760 (N_10760,N_8020,N_7996);
and U10761 (N_10761,N_8821,N_7823);
nand U10762 (N_10762,N_8245,N_8934);
nand U10763 (N_10763,N_9211,N_9869);
nand U10764 (N_10764,N_8426,N_9821);
xor U10765 (N_10765,N_7725,N_9976);
nand U10766 (N_10766,N_8388,N_9204);
nor U10767 (N_10767,N_9782,N_7956);
nor U10768 (N_10768,N_7918,N_9909);
xnor U10769 (N_10769,N_8232,N_9300);
or U10770 (N_10770,N_9216,N_7635);
nand U10771 (N_10771,N_8140,N_7530);
xnor U10772 (N_10772,N_8476,N_7668);
and U10773 (N_10773,N_8357,N_8769);
and U10774 (N_10774,N_9942,N_8436);
nor U10775 (N_10775,N_9621,N_8391);
and U10776 (N_10776,N_8445,N_8753);
xnor U10777 (N_10777,N_9413,N_9517);
xnor U10778 (N_10778,N_7990,N_9673);
or U10779 (N_10779,N_8992,N_8937);
nand U10780 (N_10780,N_8892,N_8103);
nand U10781 (N_10781,N_9743,N_8006);
xor U10782 (N_10782,N_8195,N_9633);
nand U10783 (N_10783,N_9082,N_7868);
nand U10784 (N_10784,N_7960,N_9133);
nand U10785 (N_10785,N_9948,N_8697);
and U10786 (N_10786,N_7862,N_8497);
or U10787 (N_10787,N_8201,N_8847);
nor U10788 (N_10788,N_9001,N_7716);
nand U10789 (N_10789,N_7899,N_8360);
and U10790 (N_10790,N_9863,N_8501);
nand U10791 (N_10791,N_7661,N_9116);
nor U10792 (N_10792,N_7763,N_7604);
or U10793 (N_10793,N_8070,N_9046);
nor U10794 (N_10794,N_9301,N_8306);
xnor U10795 (N_10795,N_8895,N_7915);
and U10796 (N_10796,N_8573,N_9816);
and U10797 (N_10797,N_8305,N_8699);
nand U10798 (N_10798,N_7765,N_8049);
and U10799 (N_10799,N_7634,N_8008);
nor U10800 (N_10800,N_8230,N_9914);
or U10801 (N_10801,N_9402,N_7543);
and U10802 (N_10802,N_8378,N_7727);
nand U10803 (N_10803,N_8686,N_9497);
nor U10804 (N_10804,N_9158,N_9894);
xor U10805 (N_10805,N_9866,N_8048);
or U10806 (N_10806,N_9458,N_8284);
xor U10807 (N_10807,N_8508,N_8073);
or U10808 (N_10808,N_8623,N_9657);
or U10809 (N_10809,N_9958,N_8618);
or U10810 (N_10810,N_9717,N_7980);
or U10811 (N_10811,N_9042,N_7989);
xor U10812 (N_10812,N_8861,N_7855);
nand U10813 (N_10813,N_7689,N_8543);
nand U10814 (N_10814,N_8485,N_7864);
nor U10815 (N_10815,N_7937,N_9123);
nor U10816 (N_10816,N_9177,N_9102);
xor U10817 (N_10817,N_7683,N_7510);
and U10818 (N_10818,N_9156,N_9663);
nor U10819 (N_10819,N_7987,N_7889);
or U10820 (N_10820,N_8630,N_8165);
xor U10821 (N_10821,N_9713,N_9076);
and U10822 (N_10822,N_8554,N_8600);
nor U10823 (N_10823,N_7686,N_8831);
nor U10824 (N_10824,N_9587,N_9059);
nand U10825 (N_10825,N_9662,N_8579);
xnor U10826 (N_10826,N_9898,N_9875);
nand U10827 (N_10827,N_8265,N_9591);
or U10828 (N_10828,N_8124,N_8546);
nand U10829 (N_10829,N_8651,N_9526);
nor U10830 (N_10830,N_9130,N_7594);
or U10831 (N_10831,N_8696,N_9577);
and U10832 (N_10832,N_8972,N_8514);
or U10833 (N_10833,N_9099,N_9500);
nand U10834 (N_10834,N_8088,N_9602);
nand U10835 (N_10835,N_9288,N_9542);
and U10836 (N_10836,N_8046,N_8024);
nand U10837 (N_10837,N_8104,N_7936);
nor U10838 (N_10838,N_7997,N_8392);
nand U10839 (N_10839,N_9521,N_9950);
and U10840 (N_10840,N_9112,N_9916);
nor U10841 (N_10841,N_9072,N_8762);
nand U10842 (N_10842,N_9619,N_9598);
xor U10843 (N_10843,N_9203,N_8310);
nor U10844 (N_10844,N_7613,N_8534);
xor U10845 (N_10845,N_9371,N_9549);
nand U10846 (N_10846,N_9729,N_9353);
or U10847 (N_10847,N_7526,N_8568);
or U10848 (N_10848,N_8458,N_9265);
nand U10849 (N_10849,N_9381,N_9129);
and U10850 (N_10850,N_8270,N_9407);
and U10851 (N_10851,N_9795,N_7821);
and U10852 (N_10852,N_9561,N_8915);
and U10853 (N_10853,N_9478,N_8499);
and U10854 (N_10854,N_7861,N_8055);
and U10855 (N_10855,N_9599,N_8732);
nor U10856 (N_10856,N_8900,N_9751);
nor U10857 (N_10857,N_8553,N_8106);
nand U10858 (N_10858,N_9077,N_7625);
nor U10859 (N_10859,N_8065,N_7584);
or U10860 (N_10860,N_9490,N_8601);
nand U10861 (N_10861,N_9726,N_8076);
nand U10862 (N_10862,N_8467,N_9275);
or U10863 (N_10863,N_8550,N_8814);
and U10864 (N_10864,N_9653,N_9535);
xor U10865 (N_10865,N_9968,N_8929);
nand U10866 (N_10866,N_7813,N_7583);
or U10867 (N_10867,N_9222,N_8728);
nor U10868 (N_10868,N_9791,N_7524);
or U10869 (N_10869,N_8873,N_9279);
nand U10870 (N_10870,N_7787,N_7779);
or U10871 (N_10871,N_9723,N_8162);
and U10872 (N_10872,N_8884,N_9319);
nand U10873 (N_10873,N_9172,N_9647);
xor U10874 (N_10874,N_9934,N_9845);
nor U10875 (N_10875,N_7929,N_9986);
xnor U10876 (N_10876,N_9217,N_8523);
xor U10877 (N_10877,N_7701,N_9395);
and U10878 (N_10878,N_9343,N_7908);
or U10879 (N_10879,N_7629,N_9225);
nor U10880 (N_10880,N_8160,N_9718);
and U10881 (N_10881,N_7972,N_8331);
or U10882 (N_10882,N_9148,N_9688);
and U10883 (N_10883,N_7857,N_7516);
and U10884 (N_10884,N_8815,N_7752);
or U10885 (N_10885,N_9045,N_9559);
xor U10886 (N_10886,N_9364,N_7622);
nand U10887 (N_10887,N_8796,N_8585);
nor U10888 (N_10888,N_7618,N_8776);
nor U10889 (N_10889,N_9811,N_9975);
and U10890 (N_10890,N_9820,N_9120);
nor U10891 (N_10891,N_9605,N_8402);
or U10892 (N_10892,N_7565,N_8307);
or U10893 (N_10893,N_9737,N_9615);
nand U10894 (N_10894,N_8967,N_8755);
and U10895 (N_10895,N_9334,N_8890);
nor U10896 (N_10896,N_9397,N_9767);
or U10897 (N_10897,N_9788,N_9095);
and U10898 (N_10898,N_7947,N_8169);
or U10899 (N_10899,N_8072,N_7637);
and U10900 (N_10900,N_7590,N_9538);
and U10901 (N_10901,N_9215,N_9137);
and U10902 (N_10902,N_9234,N_9054);
or U10903 (N_10903,N_7983,N_8500);
xor U10904 (N_10904,N_9574,N_9711);
or U10905 (N_10905,N_9843,N_9684);
nand U10906 (N_10906,N_9361,N_8966);
nor U10907 (N_10907,N_9936,N_8680);
xnor U10908 (N_10908,N_8607,N_9814);
and U10909 (N_10909,N_9329,N_9576);
nand U10910 (N_10910,N_7515,N_7571);
nor U10911 (N_10911,N_7638,N_8628);
and U10912 (N_10912,N_7573,N_8885);
nand U10913 (N_10913,N_7580,N_7607);
and U10914 (N_10914,N_7579,N_7577);
nand U10915 (N_10915,N_8060,N_8163);
and U10916 (N_10916,N_9033,N_7611);
nor U10917 (N_10917,N_8037,N_8278);
nand U10918 (N_10918,N_9038,N_8525);
nor U10919 (N_10919,N_8015,N_9772);
nand U10920 (N_10920,N_8889,N_9487);
nand U10921 (N_10921,N_7528,N_9338);
nor U10922 (N_10922,N_7869,N_8276);
nand U10923 (N_10923,N_9340,N_9226);
nor U10924 (N_10924,N_8479,N_8612);
and U10925 (N_10925,N_9434,N_7523);
or U10926 (N_10926,N_7881,N_8998);
and U10927 (N_10927,N_9877,N_9941);
or U10928 (N_10928,N_8274,N_8975);
or U10929 (N_10929,N_9313,N_7839);
and U10930 (N_10930,N_8650,N_9509);
nand U10931 (N_10931,N_9051,N_9769);
xor U10932 (N_10932,N_8852,N_8137);
nor U10933 (N_10933,N_8261,N_8691);
nand U10934 (N_10934,N_7575,N_8480);
and U10935 (N_10935,N_8213,N_8927);
nor U10936 (N_10936,N_8866,N_9722);
nor U10937 (N_10937,N_7921,N_9842);
nor U10938 (N_10938,N_9025,N_7587);
nor U10939 (N_10939,N_7703,N_9142);
xor U10940 (N_10940,N_9383,N_8018);
nor U10941 (N_10941,N_8486,N_8430);
nand U10942 (N_10942,N_8716,N_8727);
and U10943 (N_10943,N_9078,N_8738);
or U10944 (N_10944,N_9424,N_7847);
or U10945 (N_10945,N_8056,N_9925);
and U10946 (N_10946,N_9632,N_7589);
and U10947 (N_10947,N_9518,N_7641);
nor U10948 (N_10948,N_9214,N_8580);
xor U10949 (N_10949,N_7837,N_8009);
and U10950 (N_10950,N_9147,N_9170);
nor U10951 (N_10951,N_9200,N_8694);
or U10952 (N_10952,N_7700,N_8801);
and U10953 (N_10953,N_8080,N_9378);
or U10954 (N_10954,N_8951,N_8262);
or U10955 (N_10955,N_9230,N_9286);
and U10956 (N_10956,N_9335,N_9472);
xor U10957 (N_10957,N_7653,N_8551);
xnor U10958 (N_10958,N_8735,N_9537);
or U10959 (N_10959,N_7710,N_8724);
nand U10960 (N_10960,N_8302,N_8541);
nor U10961 (N_10961,N_8752,N_7928);
nor U10962 (N_10962,N_7550,N_8626);
nand U10963 (N_10963,N_8130,N_7677);
xnor U10964 (N_10964,N_7721,N_9488);
xnor U10965 (N_10965,N_8381,N_9957);
nand U10966 (N_10966,N_9885,N_9258);
or U10967 (N_10967,N_9710,N_9241);
or U10968 (N_10968,N_8407,N_7674);
xor U10969 (N_10969,N_8760,N_9739);
nand U10970 (N_10970,N_8721,N_8443);
xnor U10971 (N_10971,N_9554,N_8886);
or U10972 (N_10972,N_9882,N_7800);
xnor U10973 (N_10973,N_7803,N_9423);
or U10974 (N_10974,N_8713,N_8318);
xor U10975 (N_10975,N_9379,N_9506);
nand U10976 (N_10976,N_8872,N_8649);
nor U10977 (N_10977,N_7814,N_8659);
or U10978 (N_10978,N_9693,N_9453);
and U10979 (N_10979,N_9888,N_7518);
nor U10980 (N_10980,N_8289,N_8281);
nand U10981 (N_10981,N_7632,N_9310);
xor U10982 (N_10982,N_8156,N_8475);
nand U10983 (N_10983,N_7525,N_8823);
xor U10984 (N_10984,N_9235,N_8112);
xor U10985 (N_10985,N_8340,N_8993);
nor U10986 (N_10986,N_9853,N_9856);
nand U10987 (N_10987,N_7924,N_7984);
nand U10988 (N_10988,N_9284,N_9154);
nor U10989 (N_10989,N_9689,N_9281);
or U10990 (N_10990,N_9267,N_7539);
and U10991 (N_10991,N_9677,N_8067);
and U10992 (N_10992,N_8428,N_8569);
nand U10993 (N_10993,N_7627,N_8384);
xor U10994 (N_10994,N_9858,N_8120);
and U10995 (N_10995,N_7642,N_7517);
nor U10996 (N_10996,N_8061,N_7917);
and U10997 (N_10997,N_9132,N_8035);
nor U10998 (N_10998,N_9386,N_9081);
and U10999 (N_10999,N_8596,N_8086);
or U11000 (N_11000,N_8688,N_9584);
or U11001 (N_11001,N_9266,N_9088);
and U11002 (N_11002,N_8804,N_9295);
nand U11003 (N_11003,N_8454,N_7672);
and U11004 (N_11004,N_9468,N_7723);
or U11005 (N_11005,N_9921,N_7854);
nand U11006 (N_11006,N_9583,N_9841);
and U11007 (N_11007,N_9608,N_9798);
nor U11008 (N_11008,N_7538,N_8828);
xnor U11009 (N_11009,N_9616,N_7714);
xnor U11010 (N_11010,N_8587,N_8282);
xnor U11011 (N_11011,N_8255,N_8052);
or U11012 (N_11012,N_7808,N_9864);
nor U11013 (N_11013,N_8642,N_9125);
or U11014 (N_11014,N_8744,N_9969);
nor U11015 (N_11015,N_7603,N_9922);
xnor U11016 (N_11016,N_9236,N_8745);
xnor U11017 (N_11017,N_7500,N_7678);
and U11018 (N_11018,N_8063,N_8547);
nor U11019 (N_11019,N_8258,N_8667);
nor U11020 (N_11020,N_8489,N_9604);
nor U11021 (N_11021,N_7699,N_8002);
nor U11022 (N_11022,N_8096,N_9793);
xor U11023 (N_11023,N_9734,N_9473);
nand U11024 (N_11024,N_9886,N_9394);
nor U11025 (N_11025,N_9646,N_9971);
nor U11026 (N_11026,N_8876,N_7931);
and U11027 (N_11027,N_8679,N_8843);
and U11028 (N_11028,N_9186,N_9757);
or U11029 (N_11029,N_8933,N_9644);
nand U11030 (N_11030,N_8794,N_8136);
xor U11031 (N_11031,N_7729,N_8175);
and U11032 (N_11032,N_7781,N_8928);
or U11033 (N_11033,N_8377,N_8010);
and U11034 (N_11034,N_9022,N_8153);
xnor U11035 (N_11035,N_9212,N_8296);
and U11036 (N_11036,N_7807,N_9585);
and U11037 (N_11037,N_8991,N_8674);
and U11038 (N_11038,N_8656,N_9552);
nor U11039 (N_11039,N_8421,N_8898);
nor U11040 (N_11040,N_9626,N_9166);
and U11041 (N_11041,N_9742,N_8084);
or U11042 (N_11042,N_8147,N_7820);
or U11043 (N_11043,N_9415,N_8819);
xor U11044 (N_11044,N_9939,N_7772);
xor U11045 (N_11045,N_9836,N_9829);
nor U11046 (N_11046,N_9883,N_7514);
or U11047 (N_11047,N_8582,N_8025);
xor U11048 (N_11048,N_8672,N_8215);
xnor U11049 (N_11049,N_8257,N_8896);
or U11050 (N_11050,N_9928,N_9913);
nor U11051 (N_11051,N_9590,N_8930);
nor U11052 (N_11052,N_8369,N_8074);
nand U11053 (N_11053,N_8424,N_8238);
or U11054 (N_11054,N_7806,N_8973);
nor U11055 (N_11055,N_7616,N_9897);
and U11056 (N_11056,N_9233,N_8150);
and U11057 (N_11057,N_8730,N_8717);
and U11058 (N_11058,N_7544,N_9278);
xnor U11059 (N_11059,N_8414,N_7760);
and U11060 (N_11060,N_8277,N_8974);
xnor U11061 (N_11061,N_9746,N_7898);
nor U11062 (N_11062,N_8564,N_8869);
xor U11063 (N_11063,N_8234,N_8502);
nor U11064 (N_11064,N_9483,N_8637);
or U11065 (N_11065,N_8908,N_9988);
xnor U11066 (N_11066,N_9463,N_7601);
xnor U11067 (N_11067,N_8202,N_8775);
and U11068 (N_11068,N_9457,N_8011);
nand U11069 (N_11069,N_7719,N_9846);
nor U11070 (N_11070,N_9347,N_9660);
nor U11071 (N_11071,N_8782,N_8911);
nand U11072 (N_11072,N_7819,N_7554);
xor U11073 (N_11073,N_8157,N_7911);
and U11074 (N_11074,N_9797,N_8668);
nor U11075 (N_11075,N_9899,N_9111);
and U11076 (N_11076,N_9385,N_8346);
nand U11077 (N_11077,N_8196,N_9508);
nand U11078 (N_11078,N_8606,N_7967);
and U11079 (N_11079,N_9441,N_7591);
or U11080 (N_11080,N_7835,N_9826);
xnor U11081 (N_11081,N_9202,N_8962);
nand U11082 (N_11082,N_9935,N_8350);
nor U11083 (N_11083,N_8990,N_8465);
and U11084 (N_11084,N_8731,N_9306);
and U11085 (N_11085,N_7794,N_9567);
nor U11086 (N_11086,N_7809,N_8102);
nor U11087 (N_11087,N_7916,N_7944);
nor U11088 (N_11088,N_8286,N_7738);
and U11089 (N_11089,N_9658,N_9731);
nand U11090 (N_11090,N_8867,N_8604);
nor U11091 (N_11091,N_8535,N_8241);
xor U11092 (N_11092,N_7977,N_8275);
or U11093 (N_11093,N_9065,N_8363);
xnor U11094 (N_11094,N_7906,N_9740);
xor U11095 (N_11095,N_9290,N_8586);
nor U11096 (N_11096,N_7698,N_8210);
and U11097 (N_11097,N_9901,N_9634);
or U11098 (N_11098,N_9370,N_8577);
xnor U11099 (N_11099,N_9752,N_9057);
or U11100 (N_11100,N_9333,N_8321);
nand U11101 (N_11101,N_8787,N_9121);
nand U11102 (N_11102,N_7695,N_9034);
and U11103 (N_11103,N_7706,N_7662);
or U11104 (N_11104,N_9476,N_9223);
nor U11105 (N_11105,N_8978,N_7970);
xor U11106 (N_11106,N_8863,N_8417);
xor U11107 (N_11107,N_7666,N_7966);
nand U11108 (N_11108,N_8957,N_8936);
or U11109 (N_11109,N_8142,N_7614);
xnor U11110 (N_11110,N_7650,N_7578);
and U11111 (N_11111,N_9903,N_9872);
nand U11112 (N_11112,N_9445,N_9103);
or U11113 (N_11113,N_7985,N_7561);
nor U11114 (N_11114,N_7512,N_9579);
xor U11115 (N_11115,N_8218,N_8956);
or U11116 (N_11116,N_8751,N_9844);
nor U11117 (N_11117,N_9005,N_9607);
and U11118 (N_11118,N_8487,N_7682);
xor U11119 (N_11119,N_7612,N_8095);
or U11120 (N_11120,N_9169,N_7890);
xnor U11121 (N_11121,N_8984,N_9924);
or U11122 (N_11122,N_9738,N_8542);
and U11123 (N_11123,N_8143,N_8692);
xor U11124 (N_11124,N_9790,N_8457);
and U11125 (N_11125,N_7742,N_7684);
xor U11126 (N_11126,N_9043,N_9327);
xnor U11127 (N_11127,N_9422,N_9164);
nand U11128 (N_11128,N_9178,N_7971);
xnor U11129 (N_11129,N_9069,N_8575);
xnor U11130 (N_11130,N_9144,N_9666);
or U11131 (N_11131,N_9377,N_8178);
nor U11132 (N_11132,N_9727,N_7741);
nand U11133 (N_11133,N_8739,N_8671);
xnor U11134 (N_11134,N_8251,N_9461);
nand U11135 (N_11135,N_9128,N_9686);
nand U11136 (N_11136,N_7981,N_7643);
nand U11137 (N_11137,N_7896,N_8440);
and U11138 (N_11138,N_9951,N_9787);
and U11139 (N_11139,N_9566,N_9700);
or U11140 (N_11140,N_8687,N_9655);
xor U11141 (N_11141,N_7958,N_7831);
and U11142 (N_11142,N_7910,N_9809);
and U11143 (N_11143,N_7624,N_8921);
and U11144 (N_11144,N_8379,N_8763);
nand U11145 (N_11145,N_8565,N_8924);
nand U11146 (N_11146,N_9697,N_9479);
xnor U11147 (N_11147,N_8544,N_9571);
and U11148 (N_11148,N_8075,N_8848);
or U11149 (N_11149,N_8149,N_9840);
and U11150 (N_11150,N_9498,N_8117);
nand U11151 (N_11151,N_9030,N_9035);
xnor U11152 (N_11152,N_8034,N_8053);
nand U11153 (N_11153,N_8338,N_9372);
nand U11154 (N_11154,N_7553,N_8425);
nand U11155 (N_11155,N_9242,N_7610);
or U11156 (N_11156,N_9084,N_8409);
nand U11157 (N_11157,N_8645,N_9097);
or U11158 (N_11158,N_8364,N_9755);
or U11159 (N_11159,N_9707,N_9702);
or U11160 (N_11160,N_9416,N_7850);
nor U11161 (N_11161,N_8354,N_9196);
and U11162 (N_11162,N_7548,N_9703);
xor U11163 (N_11163,N_9246,N_8557);
or U11164 (N_11164,N_8799,N_8353);
and U11165 (N_11165,N_8701,N_9944);
xnor U11166 (N_11166,N_9375,N_7712);
xnor U11167 (N_11167,N_9134,N_8702);
nand U11168 (N_11168,N_9931,N_8297);
nor U11169 (N_11169,N_7920,N_7846);
xnor U11170 (N_11170,N_8114,N_8419);
nand U11171 (N_11171,N_7563,N_9665);
xnor U11172 (N_11172,N_7720,N_8235);
nor U11173 (N_11173,N_8026,N_9822);
and U11174 (N_11174,N_9753,N_9625);
nand U11175 (N_11175,N_7866,N_8857);
nor U11176 (N_11176,N_8226,N_9981);
nor U11177 (N_11177,N_9690,N_8902);
xnor U11178 (N_11178,N_8822,N_8878);
xor U11179 (N_11179,N_9118,N_9271);
or U11180 (N_11180,N_9960,N_8813);
and U11181 (N_11181,N_8538,N_9680);
nand U11182 (N_11182,N_9421,N_8256);
nor U11183 (N_11183,N_9189,N_9699);
xnor U11184 (N_11184,N_7736,N_7946);
and U11185 (N_11185,N_8181,N_8225);
nor U11186 (N_11186,N_9998,N_8622);
and U11187 (N_11187,N_8299,N_8355);
nand U11188 (N_11188,N_8949,N_8115);
xnor U11189 (N_11189,N_8199,N_8910);
and U11190 (N_11190,N_8019,N_9199);
nand U11191 (N_11191,N_7939,N_7657);
nand U11192 (N_11192,N_8560,N_7694);
or U11193 (N_11193,N_8437,N_9382);
nor U11194 (N_11194,N_9685,N_9143);
or U11195 (N_11195,N_7978,N_8570);
xor U11196 (N_11196,N_7867,N_7644);
nor U11197 (N_11197,N_9514,N_9565);
xnor U11198 (N_11198,N_8239,N_9190);
xor U11199 (N_11199,N_9047,N_9198);
xnor U11200 (N_11200,N_9980,N_8963);
or U11201 (N_11201,N_9977,N_7788);
and U11202 (N_11202,N_9895,N_9834);
or U11203 (N_11203,N_9994,N_8341);
or U11204 (N_11204,N_9053,N_8082);
or U11205 (N_11205,N_9593,N_7907);
or U11206 (N_11206,N_9420,N_7913);
nor U11207 (N_11207,N_7836,N_7874);
xor U11208 (N_11208,N_8729,N_8561);
nor U11209 (N_11209,N_8382,N_8211);
nand U11210 (N_11210,N_7534,N_9008);
and U11211 (N_11211,N_8474,N_8387);
nand U11212 (N_11212,N_8248,N_8945);
xor U11213 (N_11213,N_9031,N_7900);
nor U11214 (N_11214,N_8864,N_7941);
nor U11215 (N_11215,N_9813,N_8629);
and U11216 (N_11216,N_8527,N_9389);
or U11217 (N_11217,N_8939,N_8989);
or U11218 (N_11218,N_8733,N_9930);
nand U11219 (N_11219,N_8038,N_9320);
and U11220 (N_11220,N_8158,N_9556);
nor U11221 (N_11221,N_8678,N_9110);
nand U11222 (N_11222,N_7542,N_8333);
or U11223 (N_11223,N_8807,N_8638);
or U11224 (N_11224,N_8376,N_9437);
xor U11225 (N_11225,N_7778,N_8907);
nor U11226 (N_11226,N_8774,N_7792);
xnor U11227 (N_11227,N_7942,N_9093);
nor U11228 (N_11228,N_9489,N_9850);
or U11229 (N_11229,N_9227,N_9642);
and U11230 (N_11230,N_7564,N_8780);
xor U11231 (N_11231,N_9009,N_9104);
nand U11232 (N_11232,N_9558,N_8099);
and U11233 (N_11233,N_9411,N_9298);
xor U11234 (N_11234,N_8337,N_7592);
xor U11235 (N_11235,N_9682,N_7801);
nor U11236 (N_11236,N_9360,N_7681);
xor U11237 (N_11237,N_9013,N_9527);
nor U11238 (N_11238,N_7964,N_9174);
and U11239 (N_11239,N_8452,N_7655);
nand U11240 (N_11240,N_7886,N_9350);
and U11241 (N_11241,N_8806,N_9783);
or U11242 (N_11242,N_9052,N_8393);
or U11243 (N_11243,N_7905,N_8039);
or U11244 (N_11244,N_8757,N_8079);
nor U11245 (N_11245,N_7608,N_9026);
nand U11246 (N_11246,N_8492,N_9908);
nor U11247 (N_11247,N_9192,N_8441);
or U11248 (N_11248,N_9471,N_9493);
nand U11249 (N_11249,N_8584,N_8912);
nand U11250 (N_11250,N_8367,N_9676);
and U11251 (N_11251,N_7508,N_8970);
and U11252 (N_11252,N_9176,N_8832);
and U11253 (N_11253,N_9428,N_8435);
nand U11254 (N_11254,N_7633,N_7612);
nor U11255 (N_11255,N_9253,N_8500);
nand U11256 (N_11256,N_8668,N_8883);
or U11257 (N_11257,N_8859,N_8421);
nand U11258 (N_11258,N_8465,N_7989);
nand U11259 (N_11259,N_8967,N_9796);
nand U11260 (N_11260,N_9479,N_8576);
nor U11261 (N_11261,N_7685,N_8134);
and U11262 (N_11262,N_8708,N_9382);
and U11263 (N_11263,N_8736,N_8160);
xnor U11264 (N_11264,N_8235,N_7742);
and U11265 (N_11265,N_9641,N_9543);
xnor U11266 (N_11266,N_9084,N_8761);
xor U11267 (N_11267,N_9714,N_8433);
and U11268 (N_11268,N_7634,N_9367);
nor U11269 (N_11269,N_8590,N_8557);
xnor U11270 (N_11270,N_8627,N_9881);
or U11271 (N_11271,N_7869,N_8933);
and U11272 (N_11272,N_8041,N_9587);
or U11273 (N_11273,N_8509,N_8717);
or U11274 (N_11274,N_9256,N_7512);
or U11275 (N_11275,N_7811,N_7805);
nor U11276 (N_11276,N_8774,N_8616);
xnor U11277 (N_11277,N_9052,N_9901);
xor U11278 (N_11278,N_8506,N_7521);
nor U11279 (N_11279,N_8941,N_9900);
nor U11280 (N_11280,N_9966,N_9722);
and U11281 (N_11281,N_9001,N_7638);
and U11282 (N_11282,N_7546,N_8256);
and U11283 (N_11283,N_9991,N_9158);
nand U11284 (N_11284,N_8008,N_8289);
xor U11285 (N_11285,N_8542,N_9465);
and U11286 (N_11286,N_7778,N_8407);
or U11287 (N_11287,N_9035,N_8923);
nor U11288 (N_11288,N_9350,N_7881);
or U11289 (N_11289,N_8918,N_8053);
and U11290 (N_11290,N_8483,N_8929);
xnor U11291 (N_11291,N_9329,N_8340);
nor U11292 (N_11292,N_9211,N_8661);
xnor U11293 (N_11293,N_9858,N_8169);
nor U11294 (N_11294,N_8065,N_8222);
or U11295 (N_11295,N_9708,N_7884);
and U11296 (N_11296,N_7952,N_7702);
xnor U11297 (N_11297,N_8279,N_7862);
nor U11298 (N_11298,N_8828,N_9688);
nor U11299 (N_11299,N_8255,N_8049);
and U11300 (N_11300,N_7598,N_8427);
and U11301 (N_11301,N_8037,N_8375);
nand U11302 (N_11302,N_8974,N_8467);
and U11303 (N_11303,N_8940,N_8350);
nand U11304 (N_11304,N_9911,N_8951);
nor U11305 (N_11305,N_7971,N_9857);
nand U11306 (N_11306,N_7872,N_7803);
and U11307 (N_11307,N_9389,N_9184);
xor U11308 (N_11308,N_8006,N_9105);
nor U11309 (N_11309,N_9607,N_9644);
and U11310 (N_11310,N_8952,N_8048);
or U11311 (N_11311,N_7903,N_8080);
nor U11312 (N_11312,N_9261,N_9943);
or U11313 (N_11313,N_9417,N_9432);
nand U11314 (N_11314,N_9698,N_9077);
and U11315 (N_11315,N_8412,N_9649);
and U11316 (N_11316,N_9921,N_9635);
and U11317 (N_11317,N_8604,N_8035);
or U11318 (N_11318,N_9908,N_8843);
nand U11319 (N_11319,N_8190,N_8051);
or U11320 (N_11320,N_8570,N_9118);
nand U11321 (N_11321,N_8630,N_9201);
nand U11322 (N_11322,N_8828,N_8593);
nor U11323 (N_11323,N_7950,N_8047);
or U11324 (N_11324,N_7848,N_9046);
or U11325 (N_11325,N_8479,N_9500);
xor U11326 (N_11326,N_7561,N_8341);
xor U11327 (N_11327,N_9198,N_7681);
or U11328 (N_11328,N_9180,N_8381);
nand U11329 (N_11329,N_9664,N_8229);
nand U11330 (N_11330,N_8427,N_9972);
xnor U11331 (N_11331,N_9210,N_9063);
or U11332 (N_11332,N_9262,N_9810);
xnor U11333 (N_11333,N_8780,N_8682);
nand U11334 (N_11334,N_9836,N_8402);
xor U11335 (N_11335,N_9592,N_9808);
or U11336 (N_11336,N_9665,N_9344);
or U11337 (N_11337,N_8735,N_9125);
or U11338 (N_11338,N_7718,N_8365);
nor U11339 (N_11339,N_8598,N_9820);
and U11340 (N_11340,N_9514,N_9712);
and U11341 (N_11341,N_9354,N_8439);
nand U11342 (N_11342,N_7517,N_9336);
and U11343 (N_11343,N_9683,N_8473);
nor U11344 (N_11344,N_8101,N_7700);
or U11345 (N_11345,N_7585,N_9178);
nand U11346 (N_11346,N_9837,N_9800);
xnor U11347 (N_11347,N_7580,N_8872);
or U11348 (N_11348,N_9126,N_9437);
or U11349 (N_11349,N_8298,N_7614);
and U11350 (N_11350,N_7991,N_8055);
xnor U11351 (N_11351,N_9100,N_8452);
and U11352 (N_11352,N_9754,N_7934);
nor U11353 (N_11353,N_8510,N_8068);
nand U11354 (N_11354,N_8963,N_9483);
xor U11355 (N_11355,N_8670,N_9604);
nand U11356 (N_11356,N_8673,N_7531);
or U11357 (N_11357,N_8501,N_8119);
or U11358 (N_11358,N_8998,N_8959);
nor U11359 (N_11359,N_7820,N_8195);
xor U11360 (N_11360,N_8906,N_8061);
and U11361 (N_11361,N_7721,N_7994);
xor U11362 (N_11362,N_9527,N_9786);
nand U11363 (N_11363,N_8115,N_9181);
or U11364 (N_11364,N_8716,N_9512);
nand U11365 (N_11365,N_9661,N_8111);
and U11366 (N_11366,N_7729,N_7724);
nor U11367 (N_11367,N_8685,N_9505);
nand U11368 (N_11368,N_8296,N_8553);
and U11369 (N_11369,N_7987,N_8441);
xor U11370 (N_11370,N_8401,N_7943);
nand U11371 (N_11371,N_8835,N_9818);
or U11372 (N_11372,N_7954,N_8183);
xnor U11373 (N_11373,N_8400,N_7736);
and U11374 (N_11374,N_8648,N_8668);
or U11375 (N_11375,N_9234,N_8575);
nand U11376 (N_11376,N_7777,N_9942);
or U11377 (N_11377,N_9373,N_8842);
or U11378 (N_11378,N_8981,N_9777);
and U11379 (N_11379,N_7890,N_7974);
and U11380 (N_11380,N_7548,N_8325);
nor U11381 (N_11381,N_8699,N_9167);
and U11382 (N_11382,N_9878,N_8503);
nor U11383 (N_11383,N_8928,N_8242);
xnor U11384 (N_11384,N_8498,N_9546);
and U11385 (N_11385,N_8619,N_8671);
and U11386 (N_11386,N_9287,N_8516);
nor U11387 (N_11387,N_8715,N_8245);
nor U11388 (N_11388,N_9977,N_9359);
nor U11389 (N_11389,N_8173,N_7913);
nand U11390 (N_11390,N_8643,N_8682);
or U11391 (N_11391,N_8246,N_8366);
xnor U11392 (N_11392,N_9492,N_8608);
and U11393 (N_11393,N_8512,N_9211);
or U11394 (N_11394,N_8266,N_8780);
nand U11395 (N_11395,N_8009,N_8826);
nand U11396 (N_11396,N_8979,N_9857);
and U11397 (N_11397,N_9161,N_9854);
or U11398 (N_11398,N_8832,N_9611);
nand U11399 (N_11399,N_7919,N_8410);
or U11400 (N_11400,N_8160,N_8840);
or U11401 (N_11401,N_7518,N_9861);
nand U11402 (N_11402,N_7966,N_7977);
and U11403 (N_11403,N_8549,N_7651);
and U11404 (N_11404,N_7770,N_9683);
and U11405 (N_11405,N_8095,N_9425);
or U11406 (N_11406,N_8039,N_8788);
xor U11407 (N_11407,N_9673,N_8492);
nand U11408 (N_11408,N_9328,N_9166);
xor U11409 (N_11409,N_7622,N_9575);
and U11410 (N_11410,N_8499,N_9207);
or U11411 (N_11411,N_7546,N_9655);
nor U11412 (N_11412,N_9286,N_8213);
or U11413 (N_11413,N_7604,N_9910);
nor U11414 (N_11414,N_7543,N_7684);
nor U11415 (N_11415,N_9134,N_7520);
nand U11416 (N_11416,N_9385,N_7704);
nand U11417 (N_11417,N_8882,N_9216);
or U11418 (N_11418,N_9876,N_8358);
and U11419 (N_11419,N_8393,N_8960);
and U11420 (N_11420,N_9571,N_8094);
and U11421 (N_11421,N_8957,N_8640);
or U11422 (N_11422,N_7679,N_7945);
nor U11423 (N_11423,N_7645,N_8149);
and U11424 (N_11424,N_7886,N_7651);
and U11425 (N_11425,N_9115,N_8569);
xnor U11426 (N_11426,N_7964,N_8267);
nand U11427 (N_11427,N_9360,N_8823);
nand U11428 (N_11428,N_9528,N_8556);
nand U11429 (N_11429,N_9973,N_9167);
nand U11430 (N_11430,N_8599,N_9940);
xnor U11431 (N_11431,N_9833,N_7526);
xnor U11432 (N_11432,N_8504,N_8552);
and U11433 (N_11433,N_8019,N_9504);
nand U11434 (N_11434,N_9121,N_9181);
or U11435 (N_11435,N_7823,N_8527);
and U11436 (N_11436,N_8372,N_9025);
and U11437 (N_11437,N_8879,N_8194);
nand U11438 (N_11438,N_8214,N_8629);
nor U11439 (N_11439,N_7503,N_8055);
nand U11440 (N_11440,N_8164,N_9446);
xnor U11441 (N_11441,N_9878,N_9721);
and U11442 (N_11442,N_7591,N_9114);
nand U11443 (N_11443,N_8788,N_9555);
or U11444 (N_11444,N_9234,N_8979);
nor U11445 (N_11445,N_9627,N_8819);
nor U11446 (N_11446,N_7642,N_9812);
nand U11447 (N_11447,N_9064,N_7703);
xnor U11448 (N_11448,N_8187,N_9335);
or U11449 (N_11449,N_9577,N_9071);
xnor U11450 (N_11450,N_8172,N_9786);
and U11451 (N_11451,N_7951,N_9141);
xnor U11452 (N_11452,N_9094,N_8415);
nand U11453 (N_11453,N_8682,N_7704);
or U11454 (N_11454,N_7780,N_7906);
and U11455 (N_11455,N_9539,N_8772);
and U11456 (N_11456,N_9382,N_7659);
and U11457 (N_11457,N_7625,N_9659);
nand U11458 (N_11458,N_7845,N_9131);
nand U11459 (N_11459,N_7657,N_9657);
or U11460 (N_11460,N_8974,N_9806);
and U11461 (N_11461,N_9168,N_9374);
or U11462 (N_11462,N_7904,N_7531);
nor U11463 (N_11463,N_9657,N_8619);
nand U11464 (N_11464,N_7971,N_8978);
or U11465 (N_11465,N_7721,N_9927);
xnor U11466 (N_11466,N_8344,N_8844);
nand U11467 (N_11467,N_8516,N_9878);
or U11468 (N_11468,N_9916,N_8300);
and U11469 (N_11469,N_9335,N_8717);
and U11470 (N_11470,N_9451,N_9559);
xor U11471 (N_11471,N_8733,N_7927);
nand U11472 (N_11472,N_8754,N_8250);
nor U11473 (N_11473,N_9505,N_9139);
nor U11474 (N_11474,N_9418,N_9487);
xor U11475 (N_11475,N_8763,N_7610);
nor U11476 (N_11476,N_7997,N_9514);
and U11477 (N_11477,N_9848,N_7693);
and U11478 (N_11478,N_8083,N_7584);
nand U11479 (N_11479,N_8495,N_8645);
xor U11480 (N_11480,N_9979,N_8000);
nand U11481 (N_11481,N_9817,N_7556);
nor U11482 (N_11482,N_8993,N_7802);
nor U11483 (N_11483,N_7888,N_9174);
nor U11484 (N_11484,N_8289,N_9899);
nand U11485 (N_11485,N_8777,N_7961);
xor U11486 (N_11486,N_8945,N_8371);
and U11487 (N_11487,N_8210,N_8955);
xnor U11488 (N_11488,N_7706,N_8345);
xnor U11489 (N_11489,N_7640,N_8363);
or U11490 (N_11490,N_9023,N_8896);
and U11491 (N_11491,N_7772,N_7867);
xor U11492 (N_11492,N_9140,N_8773);
or U11493 (N_11493,N_8115,N_9681);
or U11494 (N_11494,N_7994,N_9764);
nor U11495 (N_11495,N_7988,N_7691);
or U11496 (N_11496,N_7865,N_8861);
xnor U11497 (N_11497,N_7886,N_9617);
and U11498 (N_11498,N_9791,N_8831);
xnor U11499 (N_11499,N_9802,N_8422);
xor U11500 (N_11500,N_9381,N_8571);
or U11501 (N_11501,N_9953,N_8656);
xnor U11502 (N_11502,N_8373,N_8097);
nand U11503 (N_11503,N_8266,N_9863);
nor U11504 (N_11504,N_9834,N_7717);
nand U11505 (N_11505,N_8094,N_7808);
nor U11506 (N_11506,N_9976,N_7556);
and U11507 (N_11507,N_8454,N_8991);
nand U11508 (N_11508,N_8234,N_9685);
or U11509 (N_11509,N_7698,N_9071);
nand U11510 (N_11510,N_9553,N_8386);
xor U11511 (N_11511,N_8594,N_8878);
nor U11512 (N_11512,N_9652,N_7670);
or U11513 (N_11513,N_9796,N_8374);
and U11514 (N_11514,N_7964,N_8834);
or U11515 (N_11515,N_8143,N_7681);
and U11516 (N_11516,N_8200,N_8327);
or U11517 (N_11517,N_9152,N_8956);
and U11518 (N_11518,N_7887,N_9110);
nand U11519 (N_11519,N_8381,N_8631);
xor U11520 (N_11520,N_7569,N_9392);
nand U11521 (N_11521,N_9215,N_8060);
xnor U11522 (N_11522,N_8271,N_8921);
nand U11523 (N_11523,N_8843,N_7525);
nor U11524 (N_11524,N_9173,N_9427);
and U11525 (N_11525,N_8609,N_9504);
or U11526 (N_11526,N_9643,N_7908);
nor U11527 (N_11527,N_8941,N_9403);
or U11528 (N_11528,N_8339,N_9120);
nand U11529 (N_11529,N_8447,N_9879);
nor U11530 (N_11530,N_7549,N_7889);
or U11531 (N_11531,N_8707,N_8882);
and U11532 (N_11532,N_9942,N_9129);
and U11533 (N_11533,N_8251,N_9083);
nand U11534 (N_11534,N_8815,N_8028);
nor U11535 (N_11535,N_8363,N_8187);
and U11536 (N_11536,N_7901,N_8961);
nor U11537 (N_11537,N_7500,N_9665);
nor U11538 (N_11538,N_7798,N_8226);
and U11539 (N_11539,N_7578,N_9415);
xnor U11540 (N_11540,N_7805,N_9393);
xor U11541 (N_11541,N_9429,N_9497);
xnor U11542 (N_11542,N_9832,N_8086);
xnor U11543 (N_11543,N_8305,N_8904);
and U11544 (N_11544,N_9716,N_7882);
xor U11545 (N_11545,N_9284,N_7586);
nand U11546 (N_11546,N_9722,N_9134);
nor U11547 (N_11547,N_9809,N_9582);
and U11548 (N_11548,N_9343,N_9573);
nand U11549 (N_11549,N_9547,N_7523);
and U11550 (N_11550,N_8694,N_8019);
nor U11551 (N_11551,N_8252,N_9892);
nand U11552 (N_11552,N_8068,N_8310);
nor U11553 (N_11553,N_7899,N_8773);
or U11554 (N_11554,N_9900,N_9195);
or U11555 (N_11555,N_8986,N_9564);
xnor U11556 (N_11556,N_7950,N_9023);
nor U11557 (N_11557,N_8662,N_9202);
xor U11558 (N_11558,N_9150,N_9360);
nor U11559 (N_11559,N_7633,N_9362);
xor U11560 (N_11560,N_8604,N_9311);
or U11561 (N_11561,N_8124,N_9228);
and U11562 (N_11562,N_9887,N_8872);
xor U11563 (N_11563,N_9783,N_8489);
nand U11564 (N_11564,N_8104,N_8669);
or U11565 (N_11565,N_9721,N_9169);
nand U11566 (N_11566,N_8311,N_9673);
xnor U11567 (N_11567,N_7946,N_9262);
nand U11568 (N_11568,N_9649,N_7535);
and U11569 (N_11569,N_8848,N_7548);
nand U11570 (N_11570,N_8011,N_9661);
nand U11571 (N_11571,N_8967,N_7673);
nand U11572 (N_11572,N_8624,N_8141);
nor U11573 (N_11573,N_9721,N_7741);
xnor U11574 (N_11574,N_7711,N_7954);
nand U11575 (N_11575,N_8276,N_8074);
nor U11576 (N_11576,N_8359,N_8068);
nand U11577 (N_11577,N_9002,N_8858);
nand U11578 (N_11578,N_8601,N_8021);
xor U11579 (N_11579,N_9461,N_7504);
xor U11580 (N_11580,N_8168,N_8910);
or U11581 (N_11581,N_9072,N_7673);
and U11582 (N_11582,N_7634,N_7582);
and U11583 (N_11583,N_9196,N_8897);
nand U11584 (N_11584,N_8773,N_9664);
nand U11585 (N_11585,N_9353,N_8889);
xnor U11586 (N_11586,N_9832,N_8398);
and U11587 (N_11587,N_7737,N_7587);
xor U11588 (N_11588,N_7600,N_7783);
xnor U11589 (N_11589,N_8010,N_8026);
nand U11590 (N_11590,N_8061,N_7587);
nand U11591 (N_11591,N_8585,N_7939);
nand U11592 (N_11592,N_9933,N_7739);
nand U11593 (N_11593,N_7732,N_9860);
nand U11594 (N_11594,N_9323,N_8899);
nor U11595 (N_11595,N_7907,N_8633);
xnor U11596 (N_11596,N_7547,N_8737);
and U11597 (N_11597,N_7790,N_9188);
or U11598 (N_11598,N_8469,N_9337);
or U11599 (N_11599,N_7503,N_9993);
xnor U11600 (N_11600,N_8742,N_8475);
or U11601 (N_11601,N_7698,N_7563);
and U11602 (N_11602,N_7501,N_9226);
nand U11603 (N_11603,N_7962,N_8178);
or U11604 (N_11604,N_8097,N_8627);
nand U11605 (N_11605,N_7844,N_7700);
nor U11606 (N_11606,N_8319,N_8816);
nand U11607 (N_11607,N_8387,N_8799);
nand U11608 (N_11608,N_7765,N_8956);
xnor U11609 (N_11609,N_8155,N_9806);
nor U11610 (N_11610,N_8567,N_8965);
or U11611 (N_11611,N_9913,N_9284);
or U11612 (N_11612,N_9704,N_8934);
xor U11613 (N_11613,N_8904,N_9062);
or U11614 (N_11614,N_9646,N_8704);
xor U11615 (N_11615,N_9479,N_9066);
nor U11616 (N_11616,N_9934,N_8168);
and U11617 (N_11617,N_8796,N_9837);
nand U11618 (N_11618,N_9646,N_9392);
nor U11619 (N_11619,N_8192,N_8108);
nand U11620 (N_11620,N_8075,N_9940);
and U11621 (N_11621,N_7704,N_8670);
or U11622 (N_11622,N_9260,N_9143);
nand U11623 (N_11623,N_9703,N_7749);
or U11624 (N_11624,N_7912,N_8758);
xor U11625 (N_11625,N_7749,N_9877);
or U11626 (N_11626,N_9951,N_9508);
nor U11627 (N_11627,N_9093,N_8296);
or U11628 (N_11628,N_9954,N_9731);
or U11629 (N_11629,N_7854,N_8913);
or U11630 (N_11630,N_7824,N_8207);
nor U11631 (N_11631,N_9155,N_9610);
nor U11632 (N_11632,N_9690,N_8720);
and U11633 (N_11633,N_8542,N_7801);
xor U11634 (N_11634,N_7540,N_8181);
nand U11635 (N_11635,N_7998,N_8752);
xnor U11636 (N_11636,N_9067,N_8085);
xnor U11637 (N_11637,N_7841,N_8469);
nor U11638 (N_11638,N_7936,N_7776);
nor U11639 (N_11639,N_7531,N_8668);
xor U11640 (N_11640,N_7895,N_8260);
xor U11641 (N_11641,N_9724,N_8362);
xnor U11642 (N_11642,N_8479,N_9253);
xnor U11643 (N_11643,N_9087,N_8187);
nor U11644 (N_11644,N_7896,N_9205);
or U11645 (N_11645,N_8217,N_7886);
nand U11646 (N_11646,N_9165,N_8168);
nand U11647 (N_11647,N_8958,N_8496);
nor U11648 (N_11648,N_7769,N_8233);
nand U11649 (N_11649,N_9687,N_7925);
nor U11650 (N_11650,N_9661,N_8519);
nor U11651 (N_11651,N_9905,N_7678);
xor U11652 (N_11652,N_9494,N_7645);
and U11653 (N_11653,N_8250,N_8242);
nor U11654 (N_11654,N_8759,N_8795);
xnor U11655 (N_11655,N_7764,N_8141);
nor U11656 (N_11656,N_8982,N_8624);
or U11657 (N_11657,N_8084,N_9719);
nand U11658 (N_11658,N_8192,N_8640);
nand U11659 (N_11659,N_9533,N_7848);
nor U11660 (N_11660,N_7775,N_9530);
or U11661 (N_11661,N_8547,N_9191);
or U11662 (N_11662,N_8210,N_8260);
nand U11663 (N_11663,N_9216,N_9561);
nand U11664 (N_11664,N_8081,N_9383);
xor U11665 (N_11665,N_9830,N_7574);
nor U11666 (N_11666,N_7889,N_8153);
nand U11667 (N_11667,N_8330,N_7949);
nor U11668 (N_11668,N_9076,N_8766);
and U11669 (N_11669,N_9103,N_9504);
nand U11670 (N_11670,N_8588,N_9526);
nand U11671 (N_11671,N_8840,N_7844);
or U11672 (N_11672,N_7556,N_9177);
and U11673 (N_11673,N_9576,N_9624);
and U11674 (N_11674,N_8492,N_8340);
xnor U11675 (N_11675,N_8743,N_7893);
nor U11676 (N_11676,N_8072,N_8911);
or U11677 (N_11677,N_8456,N_8545);
or U11678 (N_11678,N_8507,N_9291);
nor U11679 (N_11679,N_8739,N_8255);
or U11680 (N_11680,N_7871,N_9030);
nor U11681 (N_11681,N_9167,N_8725);
xor U11682 (N_11682,N_8632,N_9252);
xor U11683 (N_11683,N_8948,N_7803);
nor U11684 (N_11684,N_8102,N_7768);
and U11685 (N_11685,N_8746,N_7841);
or U11686 (N_11686,N_8618,N_8908);
or U11687 (N_11687,N_8074,N_8646);
or U11688 (N_11688,N_9736,N_8199);
nand U11689 (N_11689,N_8235,N_9417);
or U11690 (N_11690,N_8748,N_8234);
and U11691 (N_11691,N_9408,N_9948);
xnor U11692 (N_11692,N_9024,N_7880);
xnor U11693 (N_11693,N_8612,N_8865);
nand U11694 (N_11694,N_7724,N_7849);
nand U11695 (N_11695,N_9167,N_7862);
xnor U11696 (N_11696,N_8137,N_9907);
xnor U11697 (N_11697,N_8091,N_8504);
nand U11698 (N_11698,N_9667,N_8309);
nand U11699 (N_11699,N_8818,N_8842);
xor U11700 (N_11700,N_9460,N_9949);
nand U11701 (N_11701,N_9200,N_8553);
or U11702 (N_11702,N_9750,N_8185);
or U11703 (N_11703,N_9892,N_7629);
nor U11704 (N_11704,N_9646,N_8428);
nor U11705 (N_11705,N_9608,N_9612);
and U11706 (N_11706,N_8855,N_8487);
nand U11707 (N_11707,N_9535,N_9441);
nand U11708 (N_11708,N_9499,N_9560);
or U11709 (N_11709,N_9862,N_7723);
xor U11710 (N_11710,N_9111,N_8914);
nand U11711 (N_11711,N_8204,N_8643);
and U11712 (N_11712,N_7620,N_8828);
xor U11713 (N_11713,N_9495,N_7877);
nand U11714 (N_11714,N_8867,N_7789);
nand U11715 (N_11715,N_9878,N_8011);
nand U11716 (N_11716,N_9967,N_8169);
and U11717 (N_11717,N_8330,N_8576);
or U11718 (N_11718,N_9098,N_7555);
or U11719 (N_11719,N_8370,N_9910);
or U11720 (N_11720,N_7777,N_8050);
nor U11721 (N_11721,N_8846,N_9161);
and U11722 (N_11722,N_8941,N_7993);
nor U11723 (N_11723,N_8197,N_8263);
nor U11724 (N_11724,N_9707,N_9204);
nor U11725 (N_11725,N_9760,N_8629);
xor U11726 (N_11726,N_9799,N_9963);
xor U11727 (N_11727,N_9087,N_8266);
and U11728 (N_11728,N_9343,N_8558);
nand U11729 (N_11729,N_8704,N_8389);
or U11730 (N_11730,N_7903,N_9658);
nor U11731 (N_11731,N_7841,N_8666);
nor U11732 (N_11732,N_8179,N_9894);
and U11733 (N_11733,N_8370,N_7699);
and U11734 (N_11734,N_8622,N_8288);
nand U11735 (N_11735,N_9630,N_8865);
xnor U11736 (N_11736,N_9174,N_8452);
or U11737 (N_11737,N_8047,N_9622);
nor U11738 (N_11738,N_9041,N_7872);
or U11739 (N_11739,N_7833,N_8188);
nand U11740 (N_11740,N_7597,N_9464);
or U11741 (N_11741,N_9616,N_8644);
or U11742 (N_11742,N_9102,N_8209);
nand U11743 (N_11743,N_8721,N_9220);
and U11744 (N_11744,N_9830,N_7632);
and U11745 (N_11745,N_7716,N_9384);
nor U11746 (N_11746,N_9023,N_8877);
and U11747 (N_11747,N_9212,N_8179);
or U11748 (N_11748,N_8309,N_9327);
xnor U11749 (N_11749,N_8816,N_8400);
nor U11750 (N_11750,N_9197,N_8527);
or U11751 (N_11751,N_7634,N_9829);
nand U11752 (N_11752,N_8217,N_9797);
or U11753 (N_11753,N_8678,N_8170);
nor U11754 (N_11754,N_8112,N_7609);
xnor U11755 (N_11755,N_9218,N_7601);
and U11756 (N_11756,N_9754,N_8289);
or U11757 (N_11757,N_9706,N_7795);
xnor U11758 (N_11758,N_8608,N_7863);
nand U11759 (N_11759,N_9670,N_9591);
nor U11760 (N_11760,N_8768,N_9554);
nor U11761 (N_11761,N_7793,N_8424);
nand U11762 (N_11762,N_7622,N_8902);
xnor U11763 (N_11763,N_7604,N_9880);
nor U11764 (N_11764,N_7975,N_9016);
nor U11765 (N_11765,N_9880,N_8348);
or U11766 (N_11766,N_8211,N_8237);
nor U11767 (N_11767,N_8145,N_9572);
or U11768 (N_11768,N_8577,N_8221);
and U11769 (N_11769,N_8748,N_8977);
nor U11770 (N_11770,N_9980,N_8075);
nand U11771 (N_11771,N_9044,N_9318);
nor U11772 (N_11772,N_8133,N_9057);
or U11773 (N_11773,N_9749,N_7830);
and U11774 (N_11774,N_9285,N_9857);
nor U11775 (N_11775,N_9666,N_9891);
nor U11776 (N_11776,N_9488,N_9868);
xnor U11777 (N_11777,N_8071,N_8445);
nand U11778 (N_11778,N_7541,N_8732);
nand U11779 (N_11779,N_9315,N_9475);
or U11780 (N_11780,N_7890,N_8446);
nand U11781 (N_11781,N_8226,N_8872);
or U11782 (N_11782,N_8287,N_9029);
nor U11783 (N_11783,N_8789,N_8486);
nand U11784 (N_11784,N_9974,N_9504);
xor U11785 (N_11785,N_9816,N_9804);
and U11786 (N_11786,N_9399,N_9978);
nand U11787 (N_11787,N_8642,N_9482);
nor U11788 (N_11788,N_8068,N_8396);
and U11789 (N_11789,N_8431,N_9734);
and U11790 (N_11790,N_9076,N_8407);
nor U11791 (N_11791,N_9450,N_8338);
xor U11792 (N_11792,N_8705,N_8996);
xor U11793 (N_11793,N_7722,N_7801);
nand U11794 (N_11794,N_9060,N_8414);
and U11795 (N_11795,N_7969,N_7917);
xor U11796 (N_11796,N_9160,N_9878);
and U11797 (N_11797,N_9436,N_8301);
and U11798 (N_11798,N_9745,N_9371);
xnor U11799 (N_11799,N_9005,N_7795);
xor U11800 (N_11800,N_9063,N_8906);
or U11801 (N_11801,N_7856,N_9626);
nor U11802 (N_11802,N_7819,N_8914);
xnor U11803 (N_11803,N_7732,N_9702);
nand U11804 (N_11804,N_8477,N_9350);
and U11805 (N_11805,N_9776,N_9268);
nor U11806 (N_11806,N_7776,N_9471);
and U11807 (N_11807,N_8029,N_8501);
nand U11808 (N_11808,N_8718,N_9126);
xnor U11809 (N_11809,N_8093,N_8354);
or U11810 (N_11810,N_8435,N_8528);
xor U11811 (N_11811,N_9338,N_9168);
nor U11812 (N_11812,N_9204,N_7566);
or U11813 (N_11813,N_8213,N_8359);
and U11814 (N_11814,N_7674,N_9688);
nand U11815 (N_11815,N_7598,N_9849);
or U11816 (N_11816,N_9457,N_7574);
and U11817 (N_11817,N_9242,N_9626);
or U11818 (N_11818,N_8152,N_9422);
xor U11819 (N_11819,N_8244,N_9312);
nand U11820 (N_11820,N_7706,N_9870);
nand U11821 (N_11821,N_8328,N_8548);
or U11822 (N_11822,N_7920,N_8599);
and U11823 (N_11823,N_8968,N_8094);
or U11824 (N_11824,N_8880,N_7608);
and U11825 (N_11825,N_8047,N_9828);
and U11826 (N_11826,N_9608,N_9745);
xnor U11827 (N_11827,N_8729,N_8644);
nand U11828 (N_11828,N_9777,N_9854);
nor U11829 (N_11829,N_8222,N_9934);
nor U11830 (N_11830,N_8282,N_9840);
nor U11831 (N_11831,N_9693,N_7629);
xnor U11832 (N_11832,N_9797,N_9842);
nand U11833 (N_11833,N_7742,N_8516);
or U11834 (N_11834,N_7624,N_7560);
nor U11835 (N_11835,N_8398,N_8995);
nand U11836 (N_11836,N_7717,N_9438);
xnor U11837 (N_11837,N_8828,N_9173);
xor U11838 (N_11838,N_7724,N_9380);
nand U11839 (N_11839,N_7506,N_9804);
nor U11840 (N_11840,N_9613,N_9985);
nand U11841 (N_11841,N_9552,N_9361);
nand U11842 (N_11842,N_9825,N_7507);
or U11843 (N_11843,N_8619,N_9467);
nand U11844 (N_11844,N_9347,N_9928);
and U11845 (N_11845,N_8469,N_7911);
nor U11846 (N_11846,N_8166,N_8522);
or U11847 (N_11847,N_8133,N_8380);
nor U11848 (N_11848,N_7579,N_8941);
or U11849 (N_11849,N_9272,N_9710);
xnor U11850 (N_11850,N_7840,N_9406);
or U11851 (N_11851,N_9323,N_8579);
nor U11852 (N_11852,N_9374,N_9304);
and U11853 (N_11853,N_8482,N_8887);
nand U11854 (N_11854,N_8697,N_8112);
xor U11855 (N_11855,N_9066,N_7969);
and U11856 (N_11856,N_9472,N_8978);
or U11857 (N_11857,N_7782,N_7810);
and U11858 (N_11858,N_8720,N_7862);
nor U11859 (N_11859,N_9823,N_9936);
nand U11860 (N_11860,N_8808,N_9613);
or U11861 (N_11861,N_9475,N_8452);
and U11862 (N_11862,N_7641,N_9533);
xor U11863 (N_11863,N_9475,N_9017);
or U11864 (N_11864,N_7959,N_9965);
nor U11865 (N_11865,N_8919,N_9611);
nor U11866 (N_11866,N_9266,N_9461);
nor U11867 (N_11867,N_7975,N_9766);
nor U11868 (N_11868,N_8101,N_9713);
or U11869 (N_11869,N_9645,N_9420);
or U11870 (N_11870,N_9573,N_8866);
nor U11871 (N_11871,N_9682,N_8871);
nor U11872 (N_11872,N_9005,N_9271);
or U11873 (N_11873,N_8412,N_9879);
and U11874 (N_11874,N_8561,N_7679);
or U11875 (N_11875,N_9698,N_9927);
nor U11876 (N_11876,N_8702,N_9090);
or U11877 (N_11877,N_9395,N_8405);
nor U11878 (N_11878,N_9525,N_8650);
nand U11879 (N_11879,N_7806,N_7644);
or U11880 (N_11880,N_8497,N_8383);
nor U11881 (N_11881,N_9804,N_9641);
and U11882 (N_11882,N_8673,N_7950);
or U11883 (N_11883,N_8973,N_8446);
nor U11884 (N_11884,N_8516,N_9754);
or U11885 (N_11885,N_8843,N_7627);
and U11886 (N_11886,N_8793,N_9373);
xor U11887 (N_11887,N_7870,N_9944);
xnor U11888 (N_11888,N_9524,N_8943);
nand U11889 (N_11889,N_9422,N_9666);
nand U11890 (N_11890,N_8689,N_8500);
nand U11891 (N_11891,N_9907,N_8901);
and U11892 (N_11892,N_8014,N_7500);
or U11893 (N_11893,N_7891,N_9544);
nand U11894 (N_11894,N_8752,N_8279);
xor U11895 (N_11895,N_7834,N_9091);
nand U11896 (N_11896,N_8601,N_8827);
or U11897 (N_11897,N_8518,N_8663);
nand U11898 (N_11898,N_8329,N_8953);
or U11899 (N_11899,N_7868,N_8063);
nand U11900 (N_11900,N_7781,N_8815);
xnor U11901 (N_11901,N_8031,N_7916);
or U11902 (N_11902,N_9091,N_7826);
and U11903 (N_11903,N_9895,N_9765);
nand U11904 (N_11904,N_9419,N_9166);
nand U11905 (N_11905,N_9982,N_9395);
and U11906 (N_11906,N_9251,N_7501);
xnor U11907 (N_11907,N_8396,N_9030);
xor U11908 (N_11908,N_9366,N_7503);
xor U11909 (N_11909,N_7569,N_9561);
nor U11910 (N_11910,N_9892,N_8573);
xnor U11911 (N_11911,N_9330,N_7845);
or U11912 (N_11912,N_8019,N_9561);
xnor U11913 (N_11913,N_9966,N_8314);
nor U11914 (N_11914,N_9149,N_8729);
and U11915 (N_11915,N_8652,N_8577);
and U11916 (N_11916,N_8659,N_9699);
nor U11917 (N_11917,N_8716,N_7558);
nand U11918 (N_11918,N_7764,N_7808);
nor U11919 (N_11919,N_9085,N_8425);
or U11920 (N_11920,N_8711,N_9215);
xor U11921 (N_11921,N_8074,N_9809);
xnor U11922 (N_11922,N_7621,N_8862);
nand U11923 (N_11923,N_7715,N_9641);
or U11924 (N_11924,N_7835,N_7594);
nor U11925 (N_11925,N_9651,N_9706);
or U11926 (N_11926,N_9961,N_8636);
nand U11927 (N_11927,N_9910,N_7521);
xor U11928 (N_11928,N_7872,N_8448);
nor U11929 (N_11929,N_9490,N_9714);
and U11930 (N_11930,N_8257,N_9619);
nor U11931 (N_11931,N_9776,N_9203);
nor U11932 (N_11932,N_8548,N_7536);
nand U11933 (N_11933,N_8754,N_9492);
or U11934 (N_11934,N_7834,N_7813);
or U11935 (N_11935,N_8606,N_8130);
nor U11936 (N_11936,N_9643,N_9500);
and U11937 (N_11937,N_9659,N_9846);
xnor U11938 (N_11938,N_7892,N_7741);
or U11939 (N_11939,N_7860,N_8396);
or U11940 (N_11940,N_9933,N_9507);
and U11941 (N_11941,N_9223,N_8845);
xnor U11942 (N_11942,N_7561,N_8227);
or U11943 (N_11943,N_8308,N_9041);
and U11944 (N_11944,N_7580,N_9486);
nand U11945 (N_11945,N_8229,N_9971);
or U11946 (N_11946,N_8211,N_8581);
nor U11947 (N_11947,N_8975,N_9989);
nand U11948 (N_11948,N_8078,N_9070);
nand U11949 (N_11949,N_8583,N_9808);
nand U11950 (N_11950,N_8490,N_7768);
xor U11951 (N_11951,N_8832,N_9334);
xnor U11952 (N_11952,N_8008,N_8049);
nand U11953 (N_11953,N_8563,N_9514);
or U11954 (N_11954,N_8930,N_9244);
nand U11955 (N_11955,N_9622,N_9296);
and U11956 (N_11956,N_7919,N_7753);
or U11957 (N_11957,N_8742,N_9135);
nor U11958 (N_11958,N_7778,N_7561);
nand U11959 (N_11959,N_8865,N_9928);
nand U11960 (N_11960,N_9153,N_8391);
and U11961 (N_11961,N_8479,N_8346);
nor U11962 (N_11962,N_8086,N_9001);
nand U11963 (N_11963,N_9498,N_8024);
nor U11964 (N_11964,N_9086,N_8269);
and U11965 (N_11965,N_9732,N_9177);
xnor U11966 (N_11966,N_9755,N_9556);
and U11967 (N_11967,N_8134,N_8815);
nor U11968 (N_11968,N_9587,N_9331);
nor U11969 (N_11969,N_7501,N_8832);
or U11970 (N_11970,N_8149,N_8377);
and U11971 (N_11971,N_9615,N_7539);
nand U11972 (N_11972,N_8774,N_8170);
xor U11973 (N_11973,N_8698,N_9732);
and U11974 (N_11974,N_9305,N_9987);
or U11975 (N_11975,N_9099,N_9903);
or U11976 (N_11976,N_8912,N_8948);
xnor U11977 (N_11977,N_9140,N_8775);
or U11978 (N_11978,N_9990,N_9642);
nor U11979 (N_11979,N_9681,N_9137);
xnor U11980 (N_11980,N_9815,N_8574);
nor U11981 (N_11981,N_7615,N_9641);
nand U11982 (N_11982,N_9219,N_9724);
nor U11983 (N_11983,N_7918,N_9529);
and U11984 (N_11984,N_9816,N_9165);
nand U11985 (N_11985,N_9138,N_9158);
nor U11986 (N_11986,N_9609,N_7586);
and U11987 (N_11987,N_9141,N_9336);
nor U11988 (N_11988,N_8956,N_9728);
xnor U11989 (N_11989,N_9697,N_9889);
nor U11990 (N_11990,N_7758,N_8464);
or U11991 (N_11991,N_8510,N_8146);
xor U11992 (N_11992,N_9216,N_8569);
nor U11993 (N_11993,N_8170,N_9342);
nand U11994 (N_11994,N_7999,N_8211);
nor U11995 (N_11995,N_8292,N_8110);
xnor U11996 (N_11996,N_7921,N_9580);
and U11997 (N_11997,N_8983,N_8458);
xnor U11998 (N_11998,N_9014,N_7612);
and U11999 (N_11999,N_9170,N_9727);
nor U12000 (N_12000,N_7660,N_7701);
xnor U12001 (N_12001,N_8885,N_9420);
or U12002 (N_12002,N_8876,N_8562);
or U12003 (N_12003,N_9407,N_7833);
xnor U12004 (N_12004,N_8192,N_8772);
nand U12005 (N_12005,N_8536,N_9621);
and U12006 (N_12006,N_9911,N_9331);
nand U12007 (N_12007,N_8013,N_8344);
or U12008 (N_12008,N_9192,N_7672);
xor U12009 (N_12009,N_9790,N_8603);
nand U12010 (N_12010,N_9530,N_9745);
nand U12011 (N_12011,N_9117,N_9407);
and U12012 (N_12012,N_7811,N_8764);
or U12013 (N_12013,N_8047,N_8275);
or U12014 (N_12014,N_8888,N_7991);
or U12015 (N_12015,N_8419,N_8382);
nor U12016 (N_12016,N_8049,N_9248);
or U12017 (N_12017,N_9100,N_9315);
nand U12018 (N_12018,N_9123,N_9542);
or U12019 (N_12019,N_8979,N_9572);
or U12020 (N_12020,N_8980,N_7927);
and U12021 (N_12021,N_9231,N_9282);
or U12022 (N_12022,N_7673,N_8319);
and U12023 (N_12023,N_8114,N_7972);
nand U12024 (N_12024,N_8458,N_9139);
or U12025 (N_12025,N_9788,N_8360);
nand U12026 (N_12026,N_9551,N_9263);
or U12027 (N_12027,N_9530,N_7705);
nand U12028 (N_12028,N_8571,N_8646);
or U12029 (N_12029,N_9782,N_8050);
or U12030 (N_12030,N_7520,N_7793);
xor U12031 (N_12031,N_8857,N_8489);
nor U12032 (N_12032,N_9417,N_7720);
nand U12033 (N_12033,N_8883,N_7575);
nand U12034 (N_12034,N_8577,N_9530);
xor U12035 (N_12035,N_9558,N_8403);
xor U12036 (N_12036,N_8176,N_7776);
xor U12037 (N_12037,N_7838,N_9535);
or U12038 (N_12038,N_9324,N_7668);
and U12039 (N_12039,N_9311,N_9038);
and U12040 (N_12040,N_9490,N_7917);
xor U12041 (N_12041,N_9064,N_9798);
and U12042 (N_12042,N_9787,N_9721);
or U12043 (N_12043,N_8616,N_9194);
nand U12044 (N_12044,N_7858,N_7672);
or U12045 (N_12045,N_7921,N_8323);
and U12046 (N_12046,N_8668,N_8590);
nor U12047 (N_12047,N_8629,N_8827);
nor U12048 (N_12048,N_8474,N_7783);
nand U12049 (N_12049,N_8937,N_9396);
and U12050 (N_12050,N_9289,N_8743);
and U12051 (N_12051,N_9649,N_9924);
or U12052 (N_12052,N_9758,N_9148);
xor U12053 (N_12053,N_9278,N_8801);
nand U12054 (N_12054,N_8285,N_7960);
and U12055 (N_12055,N_7617,N_8165);
and U12056 (N_12056,N_8044,N_8042);
nor U12057 (N_12057,N_9221,N_9596);
xnor U12058 (N_12058,N_8073,N_7501);
nor U12059 (N_12059,N_8597,N_9615);
xnor U12060 (N_12060,N_9732,N_9230);
nand U12061 (N_12061,N_9148,N_9753);
nor U12062 (N_12062,N_9476,N_7659);
nor U12063 (N_12063,N_8919,N_7554);
nor U12064 (N_12064,N_9543,N_8451);
and U12065 (N_12065,N_9626,N_9655);
nor U12066 (N_12066,N_8310,N_9967);
nor U12067 (N_12067,N_9304,N_8063);
and U12068 (N_12068,N_8804,N_9793);
nor U12069 (N_12069,N_8957,N_9162);
and U12070 (N_12070,N_9030,N_9841);
nand U12071 (N_12071,N_8174,N_8421);
nand U12072 (N_12072,N_9328,N_8948);
nand U12073 (N_12073,N_8379,N_8327);
nand U12074 (N_12074,N_8901,N_7684);
xnor U12075 (N_12075,N_9389,N_7589);
and U12076 (N_12076,N_8812,N_8424);
nor U12077 (N_12077,N_9963,N_8980);
and U12078 (N_12078,N_9457,N_9533);
nand U12079 (N_12079,N_9526,N_8415);
xor U12080 (N_12080,N_8025,N_9706);
nand U12081 (N_12081,N_9706,N_8630);
nand U12082 (N_12082,N_8896,N_7804);
nor U12083 (N_12083,N_8719,N_8281);
nand U12084 (N_12084,N_8051,N_9655);
xor U12085 (N_12085,N_9614,N_8343);
xor U12086 (N_12086,N_7665,N_9262);
xnor U12087 (N_12087,N_8942,N_9581);
nand U12088 (N_12088,N_8833,N_8542);
or U12089 (N_12089,N_8831,N_8358);
xor U12090 (N_12090,N_8501,N_7707);
nand U12091 (N_12091,N_9240,N_7687);
and U12092 (N_12092,N_9609,N_7646);
nor U12093 (N_12093,N_9923,N_9196);
and U12094 (N_12094,N_9951,N_8390);
and U12095 (N_12095,N_8663,N_7764);
or U12096 (N_12096,N_8449,N_9304);
xor U12097 (N_12097,N_8109,N_9927);
xnor U12098 (N_12098,N_8081,N_9585);
and U12099 (N_12099,N_9617,N_9358);
nor U12100 (N_12100,N_9237,N_9998);
nor U12101 (N_12101,N_9061,N_9620);
nand U12102 (N_12102,N_8587,N_7928);
or U12103 (N_12103,N_9449,N_7526);
nand U12104 (N_12104,N_9403,N_9109);
nand U12105 (N_12105,N_7620,N_8062);
or U12106 (N_12106,N_8609,N_9870);
or U12107 (N_12107,N_8305,N_7975);
or U12108 (N_12108,N_9031,N_7694);
nor U12109 (N_12109,N_8630,N_8958);
nand U12110 (N_12110,N_8392,N_9512);
and U12111 (N_12111,N_7595,N_8514);
xor U12112 (N_12112,N_8004,N_9401);
nor U12113 (N_12113,N_7763,N_8739);
nor U12114 (N_12114,N_7531,N_7596);
or U12115 (N_12115,N_7697,N_8118);
nand U12116 (N_12116,N_7834,N_7810);
and U12117 (N_12117,N_8910,N_9846);
nor U12118 (N_12118,N_8814,N_9288);
and U12119 (N_12119,N_8497,N_8458);
nor U12120 (N_12120,N_9484,N_8030);
nand U12121 (N_12121,N_8662,N_9595);
and U12122 (N_12122,N_8758,N_8534);
nor U12123 (N_12123,N_8645,N_8718);
xor U12124 (N_12124,N_8344,N_8758);
nand U12125 (N_12125,N_9809,N_9855);
or U12126 (N_12126,N_8203,N_9089);
xnor U12127 (N_12127,N_8081,N_9832);
and U12128 (N_12128,N_7881,N_7948);
xnor U12129 (N_12129,N_8605,N_8795);
nand U12130 (N_12130,N_8782,N_9704);
or U12131 (N_12131,N_9761,N_7894);
or U12132 (N_12132,N_9723,N_8408);
nor U12133 (N_12133,N_8459,N_9201);
and U12134 (N_12134,N_8910,N_9254);
xor U12135 (N_12135,N_7759,N_8101);
or U12136 (N_12136,N_9461,N_8085);
xor U12137 (N_12137,N_8626,N_8559);
nor U12138 (N_12138,N_8075,N_8084);
and U12139 (N_12139,N_8547,N_9272);
and U12140 (N_12140,N_9719,N_9463);
xnor U12141 (N_12141,N_9577,N_9509);
and U12142 (N_12142,N_9805,N_8057);
or U12143 (N_12143,N_9943,N_7869);
nand U12144 (N_12144,N_8790,N_8340);
and U12145 (N_12145,N_7666,N_9334);
and U12146 (N_12146,N_9966,N_7908);
xnor U12147 (N_12147,N_8796,N_8611);
or U12148 (N_12148,N_8262,N_8881);
nand U12149 (N_12149,N_8418,N_8099);
xor U12150 (N_12150,N_8340,N_8263);
nand U12151 (N_12151,N_9759,N_9150);
xnor U12152 (N_12152,N_7836,N_9266);
and U12153 (N_12153,N_8632,N_7687);
and U12154 (N_12154,N_9167,N_9279);
nor U12155 (N_12155,N_7856,N_7586);
nor U12156 (N_12156,N_9559,N_9720);
nor U12157 (N_12157,N_8762,N_9805);
and U12158 (N_12158,N_8418,N_7752);
and U12159 (N_12159,N_7693,N_9330);
nor U12160 (N_12160,N_8471,N_9011);
or U12161 (N_12161,N_8565,N_9248);
xor U12162 (N_12162,N_9590,N_7907);
xnor U12163 (N_12163,N_9950,N_8817);
and U12164 (N_12164,N_9043,N_9941);
and U12165 (N_12165,N_9742,N_9610);
and U12166 (N_12166,N_7600,N_8295);
xnor U12167 (N_12167,N_9554,N_8323);
xor U12168 (N_12168,N_7521,N_9368);
nand U12169 (N_12169,N_8930,N_8387);
nand U12170 (N_12170,N_8356,N_7738);
nand U12171 (N_12171,N_9444,N_9901);
nor U12172 (N_12172,N_9433,N_8417);
nor U12173 (N_12173,N_9545,N_7691);
xor U12174 (N_12174,N_8047,N_7596);
nand U12175 (N_12175,N_7975,N_9419);
nor U12176 (N_12176,N_8277,N_7878);
and U12177 (N_12177,N_7543,N_9240);
or U12178 (N_12178,N_9070,N_7733);
or U12179 (N_12179,N_8681,N_8711);
nor U12180 (N_12180,N_9064,N_9917);
xnor U12181 (N_12181,N_9341,N_8310);
or U12182 (N_12182,N_8264,N_8572);
nor U12183 (N_12183,N_9192,N_9519);
or U12184 (N_12184,N_8125,N_8257);
nand U12185 (N_12185,N_9902,N_9878);
nor U12186 (N_12186,N_8864,N_9857);
or U12187 (N_12187,N_9777,N_7891);
or U12188 (N_12188,N_7604,N_7583);
xor U12189 (N_12189,N_7732,N_9463);
nand U12190 (N_12190,N_9928,N_8191);
nor U12191 (N_12191,N_9552,N_8847);
xnor U12192 (N_12192,N_9020,N_8840);
nand U12193 (N_12193,N_8642,N_8265);
or U12194 (N_12194,N_9160,N_8876);
or U12195 (N_12195,N_9796,N_8391);
nor U12196 (N_12196,N_9217,N_8147);
xnor U12197 (N_12197,N_8115,N_7955);
nor U12198 (N_12198,N_9671,N_8037);
xnor U12199 (N_12199,N_8724,N_9547);
nor U12200 (N_12200,N_8879,N_9089);
nand U12201 (N_12201,N_9314,N_7930);
nand U12202 (N_12202,N_8406,N_7937);
and U12203 (N_12203,N_8719,N_8092);
or U12204 (N_12204,N_8995,N_8361);
and U12205 (N_12205,N_9764,N_8379);
and U12206 (N_12206,N_9320,N_7672);
xnor U12207 (N_12207,N_7741,N_8009);
and U12208 (N_12208,N_8556,N_9855);
nor U12209 (N_12209,N_9913,N_7993);
nand U12210 (N_12210,N_7964,N_8487);
and U12211 (N_12211,N_7770,N_7806);
nor U12212 (N_12212,N_8619,N_9505);
nor U12213 (N_12213,N_7708,N_7654);
xor U12214 (N_12214,N_8719,N_8924);
xnor U12215 (N_12215,N_9876,N_9492);
and U12216 (N_12216,N_8409,N_9826);
nor U12217 (N_12217,N_9819,N_8725);
xor U12218 (N_12218,N_7839,N_8858);
or U12219 (N_12219,N_9294,N_7884);
nor U12220 (N_12220,N_9034,N_8193);
and U12221 (N_12221,N_7829,N_9251);
xnor U12222 (N_12222,N_9218,N_8497);
and U12223 (N_12223,N_8818,N_9803);
or U12224 (N_12224,N_9893,N_7526);
xnor U12225 (N_12225,N_9850,N_9593);
nand U12226 (N_12226,N_9911,N_9508);
and U12227 (N_12227,N_9714,N_8799);
nand U12228 (N_12228,N_7723,N_9342);
nand U12229 (N_12229,N_7733,N_7998);
nor U12230 (N_12230,N_9653,N_9219);
nand U12231 (N_12231,N_8592,N_8266);
xnor U12232 (N_12232,N_8879,N_7916);
nand U12233 (N_12233,N_7702,N_9647);
xor U12234 (N_12234,N_8787,N_8909);
nor U12235 (N_12235,N_9378,N_7539);
xor U12236 (N_12236,N_7805,N_9450);
and U12237 (N_12237,N_7541,N_8366);
nor U12238 (N_12238,N_9835,N_7856);
and U12239 (N_12239,N_9764,N_8031);
or U12240 (N_12240,N_8842,N_8797);
nor U12241 (N_12241,N_8179,N_9872);
or U12242 (N_12242,N_7920,N_8213);
nand U12243 (N_12243,N_9363,N_9579);
nand U12244 (N_12244,N_9123,N_9267);
or U12245 (N_12245,N_8547,N_9725);
and U12246 (N_12246,N_7767,N_9561);
or U12247 (N_12247,N_9583,N_9535);
and U12248 (N_12248,N_8703,N_9609);
nor U12249 (N_12249,N_7540,N_8847);
nor U12250 (N_12250,N_8227,N_8928);
xor U12251 (N_12251,N_8464,N_8100);
nor U12252 (N_12252,N_8989,N_9169);
and U12253 (N_12253,N_7768,N_8248);
nor U12254 (N_12254,N_8430,N_9859);
and U12255 (N_12255,N_8697,N_8469);
or U12256 (N_12256,N_9601,N_8402);
xor U12257 (N_12257,N_8445,N_8693);
and U12258 (N_12258,N_7811,N_9382);
and U12259 (N_12259,N_9203,N_9155);
and U12260 (N_12260,N_9366,N_7802);
xor U12261 (N_12261,N_7939,N_9318);
or U12262 (N_12262,N_8986,N_8091);
or U12263 (N_12263,N_8693,N_9321);
xor U12264 (N_12264,N_8869,N_9432);
nor U12265 (N_12265,N_8595,N_9893);
xor U12266 (N_12266,N_8108,N_7604);
and U12267 (N_12267,N_8792,N_9953);
nor U12268 (N_12268,N_9911,N_7588);
and U12269 (N_12269,N_7572,N_9691);
xnor U12270 (N_12270,N_7962,N_9981);
xor U12271 (N_12271,N_8962,N_9319);
and U12272 (N_12272,N_9384,N_8487);
or U12273 (N_12273,N_7633,N_8694);
xnor U12274 (N_12274,N_9864,N_9186);
and U12275 (N_12275,N_9157,N_9890);
nor U12276 (N_12276,N_8612,N_9228);
xnor U12277 (N_12277,N_8610,N_8156);
and U12278 (N_12278,N_7813,N_8242);
nand U12279 (N_12279,N_9133,N_8779);
nor U12280 (N_12280,N_8223,N_9213);
nand U12281 (N_12281,N_9113,N_8351);
nand U12282 (N_12282,N_8058,N_8054);
and U12283 (N_12283,N_7669,N_9858);
nand U12284 (N_12284,N_9506,N_8939);
and U12285 (N_12285,N_9121,N_8690);
xor U12286 (N_12286,N_8424,N_9698);
or U12287 (N_12287,N_9542,N_8003);
or U12288 (N_12288,N_8141,N_8805);
xnor U12289 (N_12289,N_8118,N_9764);
or U12290 (N_12290,N_9108,N_9314);
nand U12291 (N_12291,N_9168,N_8007);
nor U12292 (N_12292,N_9128,N_7784);
xnor U12293 (N_12293,N_8983,N_8272);
nand U12294 (N_12294,N_7947,N_7735);
and U12295 (N_12295,N_9457,N_8575);
nand U12296 (N_12296,N_8820,N_8432);
and U12297 (N_12297,N_8684,N_9356);
nor U12298 (N_12298,N_8033,N_8285);
and U12299 (N_12299,N_9704,N_9124);
and U12300 (N_12300,N_8300,N_9635);
nor U12301 (N_12301,N_7601,N_7646);
xor U12302 (N_12302,N_8222,N_8072);
or U12303 (N_12303,N_9598,N_8751);
and U12304 (N_12304,N_8671,N_7799);
and U12305 (N_12305,N_7697,N_9275);
xor U12306 (N_12306,N_7886,N_8535);
nand U12307 (N_12307,N_9066,N_8970);
and U12308 (N_12308,N_7988,N_9447);
nor U12309 (N_12309,N_8795,N_9393);
or U12310 (N_12310,N_9513,N_9597);
or U12311 (N_12311,N_8550,N_7836);
nand U12312 (N_12312,N_8608,N_8933);
nand U12313 (N_12313,N_8460,N_9346);
nand U12314 (N_12314,N_8952,N_9845);
nand U12315 (N_12315,N_9049,N_7767);
or U12316 (N_12316,N_7552,N_8907);
nor U12317 (N_12317,N_8926,N_8798);
and U12318 (N_12318,N_8145,N_8193);
and U12319 (N_12319,N_8063,N_9105);
or U12320 (N_12320,N_8462,N_8871);
nand U12321 (N_12321,N_9871,N_8113);
or U12322 (N_12322,N_8777,N_9952);
xor U12323 (N_12323,N_9305,N_8874);
or U12324 (N_12324,N_7600,N_8335);
nand U12325 (N_12325,N_8791,N_8034);
nor U12326 (N_12326,N_9396,N_8013);
or U12327 (N_12327,N_7775,N_9831);
xor U12328 (N_12328,N_8103,N_8794);
nand U12329 (N_12329,N_8685,N_9673);
and U12330 (N_12330,N_8008,N_9078);
or U12331 (N_12331,N_8995,N_9873);
nor U12332 (N_12332,N_9560,N_9625);
xor U12333 (N_12333,N_9595,N_8265);
nor U12334 (N_12334,N_9440,N_9969);
or U12335 (N_12335,N_9698,N_9075);
or U12336 (N_12336,N_8614,N_9737);
xnor U12337 (N_12337,N_8353,N_8372);
nor U12338 (N_12338,N_8698,N_9120);
nand U12339 (N_12339,N_9932,N_7506);
xor U12340 (N_12340,N_9042,N_7636);
nor U12341 (N_12341,N_8643,N_8358);
xnor U12342 (N_12342,N_8121,N_8529);
nand U12343 (N_12343,N_9811,N_9397);
and U12344 (N_12344,N_8428,N_8487);
or U12345 (N_12345,N_8381,N_8082);
or U12346 (N_12346,N_9627,N_7959);
xnor U12347 (N_12347,N_8865,N_9863);
xnor U12348 (N_12348,N_9955,N_7816);
nand U12349 (N_12349,N_8919,N_8593);
nor U12350 (N_12350,N_9440,N_8705);
or U12351 (N_12351,N_8963,N_9369);
xnor U12352 (N_12352,N_7617,N_8736);
and U12353 (N_12353,N_8935,N_8766);
nand U12354 (N_12354,N_7855,N_9126);
nand U12355 (N_12355,N_8527,N_9878);
and U12356 (N_12356,N_9665,N_9817);
and U12357 (N_12357,N_9606,N_8050);
nand U12358 (N_12358,N_9330,N_9925);
nand U12359 (N_12359,N_8982,N_8773);
nor U12360 (N_12360,N_7964,N_9168);
nand U12361 (N_12361,N_8743,N_9394);
nand U12362 (N_12362,N_9763,N_7522);
nand U12363 (N_12363,N_7887,N_8931);
or U12364 (N_12364,N_8064,N_8039);
or U12365 (N_12365,N_9557,N_9993);
nand U12366 (N_12366,N_8389,N_8402);
nor U12367 (N_12367,N_8019,N_9912);
nand U12368 (N_12368,N_7887,N_8686);
and U12369 (N_12369,N_9058,N_7967);
or U12370 (N_12370,N_8658,N_9505);
and U12371 (N_12371,N_8479,N_8543);
nor U12372 (N_12372,N_9332,N_8239);
xnor U12373 (N_12373,N_8274,N_9664);
and U12374 (N_12374,N_9799,N_9627);
or U12375 (N_12375,N_7543,N_8371);
xnor U12376 (N_12376,N_8051,N_7925);
nor U12377 (N_12377,N_9914,N_9654);
nor U12378 (N_12378,N_9167,N_9992);
nand U12379 (N_12379,N_7955,N_9825);
and U12380 (N_12380,N_7870,N_8065);
xnor U12381 (N_12381,N_8275,N_9328);
nor U12382 (N_12382,N_9844,N_8354);
and U12383 (N_12383,N_9890,N_7559);
nand U12384 (N_12384,N_8028,N_8947);
nor U12385 (N_12385,N_9499,N_8222);
nor U12386 (N_12386,N_9617,N_7608);
and U12387 (N_12387,N_8018,N_8696);
and U12388 (N_12388,N_8132,N_8557);
or U12389 (N_12389,N_9607,N_7676);
xor U12390 (N_12390,N_9811,N_8397);
and U12391 (N_12391,N_9380,N_8554);
nor U12392 (N_12392,N_8746,N_9101);
or U12393 (N_12393,N_7506,N_8588);
nand U12394 (N_12394,N_9388,N_9392);
nand U12395 (N_12395,N_9755,N_8403);
or U12396 (N_12396,N_7626,N_7961);
and U12397 (N_12397,N_8986,N_9065);
nor U12398 (N_12398,N_7955,N_7795);
and U12399 (N_12399,N_9292,N_8092);
xor U12400 (N_12400,N_7809,N_9262);
or U12401 (N_12401,N_8568,N_7869);
xor U12402 (N_12402,N_8113,N_9330);
xor U12403 (N_12403,N_9256,N_8083);
nand U12404 (N_12404,N_9463,N_9052);
nor U12405 (N_12405,N_8160,N_8909);
xnor U12406 (N_12406,N_8295,N_8374);
nor U12407 (N_12407,N_9612,N_8138);
and U12408 (N_12408,N_9291,N_8168);
nor U12409 (N_12409,N_8701,N_9043);
nand U12410 (N_12410,N_9868,N_7749);
and U12411 (N_12411,N_8012,N_9498);
xor U12412 (N_12412,N_7676,N_8967);
and U12413 (N_12413,N_9531,N_8748);
nand U12414 (N_12414,N_8937,N_8459);
or U12415 (N_12415,N_7506,N_7728);
nand U12416 (N_12416,N_8254,N_7745);
and U12417 (N_12417,N_7712,N_8517);
xor U12418 (N_12418,N_8158,N_8357);
nor U12419 (N_12419,N_9940,N_9354);
and U12420 (N_12420,N_7782,N_9982);
xor U12421 (N_12421,N_8080,N_8178);
or U12422 (N_12422,N_9691,N_9167);
xnor U12423 (N_12423,N_7930,N_8558);
and U12424 (N_12424,N_8308,N_9879);
nand U12425 (N_12425,N_8237,N_8554);
or U12426 (N_12426,N_8260,N_8952);
nor U12427 (N_12427,N_9452,N_9388);
nand U12428 (N_12428,N_7773,N_9542);
and U12429 (N_12429,N_7920,N_8676);
and U12430 (N_12430,N_9557,N_8812);
nor U12431 (N_12431,N_9699,N_7855);
nor U12432 (N_12432,N_9257,N_8011);
xor U12433 (N_12433,N_9238,N_7554);
or U12434 (N_12434,N_8430,N_8104);
or U12435 (N_12435,N_9773,N_8006);
nor U12436 (N_12436,N_9433,N_7650);
and U12437 (N_12437,N_8269,N_7899);
nor U12438 (N_12438,N_9815,N_8683);
nor U12439 (N_12439,N_8707,N_9865);
or U12440 (N_12440,N_8337,N_8093);
nand U12441 (N_12441,N_9291,N_8423);
nand U12442 (N_12442,N_7797,N_9377);
nor U12443 (N_12443,N_9284,N_9505);
xor U12444 (N_12444,N_9560,N_9223);
or U12445 (N_12445,N_7769,N_8670);
nor U12446 (N_12446,N_7567,N_7695);
or U12447 (N_12447,N_9151,N_8443);
or U12448 (N_12448,N_8288,N_8289);
xor U12449 (N_12449,N_8021,N_9187);
nand U12450 (N_12450,N_9983,N_8368);
xnor U12451 (N_12451,N_7629,N_9274);
xnor U12452 (N_12452,N_8789,N_7629);
nor U12453 (N_12453,N_8187,N_8332);
nor U12454 (N_12454,N_8492,N_7665);
nor U12455 (N_12455,N_9203,N_8277);
nand U12456 (N_12456,N_8458,N_8669);
nand U12457 (N_12457,N_8347,N_7647);
xnor U12458 (N_12458,N_8886,N_9991);
nand U12459 (N_12459,N_8322,N_8764);
or U12460 (N_12460,N_8677,N_7914);
and U12461 (N_12461,N_8214,N_7715);
nor U12462 (N_12462,N_7712,N_8093);
and U12463 (N_12463,N_9463,N_9451);
nor U12464 (N_12464,N_7945,N_9995);
and U12465 (N_12465,N_8758,N_9746);
nor U12466 (N_12466,N_9820,N_8343);
nor U12467 (N_12467,N_8561,N_8031);
and U12468 (N_12468,N_8433,N_7637);
nand U12469 (N_12469,N_9333,N_7961);
or U12470 (N_12470,N_7586,N_8604);
xor U12471 (N_12471,N_8350,N_8871);
or U12472 (N_12472,N_8416,N_8878);
nor U12473 (N_12473,N_7973,N_8925);
nand U12474 (N_12474,N_8620,N_8572);
xnor U12475 (N_12475,N_9587,N_8193);
and U12476 (N_12476,N_9219,N_8242);
nor U12477 (N_12477,N_9860,N_8075);
xnor U12478 (N_12478,N_9957,N_9569);
nand U12479 (N_12479,N_9875,N_9595);
nor U12480 (N_12480,N_9535,N_7888);
and U12481 (N_12481,N_9727,N_8894);
xnor U12482 (N_12482,N_8918,N_8080);
and U12483 (N_12483,N_8903,N_7876);
or U12484 (N_12484,N_9933,N_7725);
nor U12485 (N_12485,N_9844,N_8371);
xor U12486 (N_12486,N_8561,N_9711);
and U12487 (N_12487,N_9368,N_8409);
or U12488 (N_12488,N_9434,N_8679);
and U12489 (N_12489,N_9415,N_9082);
or U12490 (N_12490,N_9046,N_9335);
xnor U12491 (N_12491,N_9702,N_8455);
or U12492 (N_12492,N_9953,N_9881);
or U12493 (N_12493,N_8037,N_9285);
or U12494 (N_12494,N_7936,N_8179);
or U12495 (N_12495,N_9413,N_9597);
and U12496 (N_12496,N_7909,N_7785);
and U12497 (N_12497,N_9564,N_7740);
xor U12498 (N_12498,N_8755,N_7991);
nand U12499 (N_12499,N_7642,N_8810);
or U12500 (N_12500,N_10126,N_12231);
and U12501 (N_12501,N_11627,N_11989);
or U12502 (N_12502,N_12402,N_11946);
nor U12503 (N_12503,N_12264,N_10605);
or U12504 (N_12504,N_11022,N_10957);
and U12505 (N_12505,N_11529,N_10028);
or U12506 (N_12506,N_11703,N_11241);
nor U12507 (N_12507,N_11737,N_12092);
or U12508 (N_12508,N_12493,N_10435);
nand U12509 (N_12509,N_11897,N_11564);
nand U12510 (N_12510,N_11363,N_11834);
or U12511 (N_12511,N_11601,N_11464);
or U12512 (N_12512,N_12437,N_12066);
xor U12513 (N_12513,N_12495,N_10763);
or U12514 (N_12514,N_11644,N_10679);
nand U12515 (N_12515,N_12232,N_11863);
xnor U12516 (N_12516,N_12431,N_11711);
or U12517 (N_12517,N_11284,N_11632);
nor U12518 (N_12518,N_12332,N_11626);
nand U12519 (N_12519,N_12413,N_10498);
and U12520 (N_12520,N_10318,N_10439);
xor U12521 (N_12521,N_10352,N_10405);
xnor U12522 (N_12522,N_11650,N_11871);
nand U12523 (N_12523,N_12456,N_10750);
xnor U12524 (N_12524,N_12147,N_11069);
nor U12525 (N_12525,N_11215,N_10102);
or U12526 (N_12526,N_11572,N_12399);
nor U12527 (N_12527,N_11079,N_10298);
xor U12528 (N_12528,N_11164,N_11036);
and U12529 (N_12529,N_11090,N_10644);
nand U12530 (N_12530,N_11893,N_10741);
nor U12531 (N_12531,N_10351,N_10768);
nor U12532 (N_12532,N_10683,N_10146);
nand U12533 (N_12533,N_11672,N_12283);
xor U12534 (N_12534,N_11991,N_10471);
nand U12535 (N_12535,N_12131,N_12139);
and U12536 (N_12536,N_10185,N_12115);
nand U12537 (N_12537,N_12320,N_12268);
xor U12538 (N_12538,N_11294,N_11110);
xor U12539 (N_12539,N_10365,N_10936);
or U12540 (N_12540,N_11092,N_10717);
xnor U12541 (N_12541,N_10534,N_11046);
xnor U12542 (N_12542,N_10560,N_12289);
nor U12543 (N_12543,N_11362,N_10444);
and U12544 (N_12544,N_12427,N_12164);
nand U12545 (N_12545,N_11148,N_10490);
xor U12546 (N_12546,N_11059,N_10867);
nor U12547 (N_12547,N_11903,N_11189);
and U12548 (N_12548,N_11651,N_11274);
nor U12549 (N_12549,N_10825,N_11055);
nand U12550 (N_12550,N_11376,N_10826);
nand U12551 (N_12551,N_12329,N_11123);
xor U12552 (N_12552,N_11722,N_12248);
nor U12553 (N_12553,N_11965,N_10850);
or U12554 (N_12554,N_10890,N_11887);
xnor U12555 (N_12555,N_11083,N_10985);
and U12556 (N_12556,N_10424,N_11899);
nand U12557 (N_12557,N_10576,N_11548);
nor U12558 (N_12558,N_10015,N_12208);
xor U12559 (N_12559,N_10227,N_11454);
nor U12560 (N_12560,N_11996,N_11925);
xnor U12561 (N_12561,N_12022,N_11697);
nand U12562 (N_12562,N_12260,N_12040);
xor U12563 (N_12563,N_11789,N_10607);
nand U12564 (N_12564,N_11875,N_10504);
nand U12565 (N_12565,N_11931,N_11203);
or U12566 (N_12566,N_11417,N_10017);
or U12567 (N_12567,N_12154,N_10061);
or U12568 (N_12568,N_10319,N_11020);
xor U12569 (N_12569,N_12256,N_10288);
or U12570 (N_12570,N_12193,N_11790);
nand U12571 (N_12571,N_10037,N_10198);
nand U12572 (N_12572,N_12309,N_10955);
xor U12573 (N_12573,N_10987,N_12235);
and U12574 (N_12574,N_11128,N_10445);
xnor U12575 (N_12575,N_10843,N_11616);
nand U12576 (N_12576,N_10321,N_12265);
and U12577 (N_12577,N_10054,N_12042);
nor U12578 (N_12578,N_10267,N_10802);
or U12579 (N_12579,N_11485,N_10143);
nor U12580 (N_12580,N_10509,N_10497);
or U12581 (N_12581,N_11589,N_11543);
xor U12582 (N_12582,N_12168,N_11013);
xor U12583 (N_12583,N_11579,N_11990);
xor U12584 (N_12584,N_10645,N_11967);
xnor U12585 (N_12585,N_10005,N_10511);
and U12586 (N_12586,N_12420,N_10093);
and U12587 (N_12587,N_11701,N_12481);
xor U12588 (N_12588,N_10858,N_10252);
nand U12589 (N_12589,N_10922,N_11161);
nor U12590 (N_12590,N_10572,N_10415);
nor U12591 (N_12591,N_12450,N_11436);
nand U12592 (N_12592,N_12475,N_11157);
xnor U12593 (N_12593,N_10519,N_12060);
xor U12594 (N_12594,N_11388,N_11620);
xor U12595 (N_12595,N_11745,N_12061);
or U12596 (N_12596,N_12227,N_12156);
or U12597 (N_12597,N_10262,N_12225);
nand U12598 (N_12598,N_10673,N_10244);
or U12599 (N_12599,N_11209,N_10730);
xnor U12600 (N_12600,N_12093,N_10530);
xor U12601 (N_12601,N_11999,N_10708);
xnor U12602 (N_12602,N_10959,N_12343);
nor U12603 (N_12603,N_10510,N_12284);
or U12604 (N_12604,N_11142,N_12369);
and U12605 (N_12605,N_11320,N_10080);
nand U12606 (N_12606,N_10368,N_10207);
xnor U12607 (N_12607,N_10499,N_12118);
or U12608 (N_12608,N_12301,N_11188);
and U12609 (N_12609,N_11918,N_11257);
or U12610 (N_12610,N_10148,N_11151);
and U12611 (N_12611,N_12001,N_11732);
and U12612 (N_12612,N_10931,N_10817);
xnor U12613 (N_12613,N_11242,N_11207);
xnor U12614 (N_12614,N_10894,N_11104);
or U12615 (N_12615,N_12078,N_10513);
or U12616 (N_12616,N_10529,N_10698);
xnor U12617 (N_12617,N_11520,N_12465);
nand U12618 (N_12618,N_11815,N_10761);
nand U12619 (N_12619,N_10729,N_10749);
xnor U12620 (N_12620,N_11686,N_11920);
or U12621 (N_12621,N_10003,N_12352);
or U12622 (N_12622,N_12355,N_11125);
and U12623 (N_12623,N_10229,N_10819);
and U12624 (N_12624,N_11445,N_11682);
and U12625 (N_12625,N_10789,N_11523);
nand U12626 (N_12626,N_10793,N_10664);
nand U12627 (N_12627,N_10544,N_10440);
or U12628 (N_12628,N_11374,N_11258);
nor U12629 (N_12629,N_11237,N_10870);
nor U12630 (N_12630,N_10614,N_11714);
nor U12631 (N_12631,N_11959,N_11660);
nand U12632 (N_12632,N_10928,N_11533);
xnor U12633 (N_12633,N_11972,N_12238);
and U12634 (N_12634,N_12491,N_11421);
or U12635 (N_12635,N_11927,N_11071);
nand U12636 (N_12636,N_11534,N_11057);
xor U12637 (N_12637,N_10871,N_11021);
nand U12638 (N_12638,N_11120,N_10141);
nand U12639 (N_12639,N_10191,N_12432);
or U12640 (N_12640,N_10091,N_12057);
and U12641 (N_12641,N_12149,N_12104);
or U12642 (N_12642,N_11721,N_11962);
nand U12643 (N_12643,N_10205,N_11657);
nand U12644 (N_12644,N_12342,N_10376);
and U12645 (N_12645,N_10626,N_12009);
xor U12646 (N_12646,N_10864,N_10578);
and U12647 (N_12647,N_10349,N_10924);
nand U12648 (N_12648,N_11921,N_10417);
nand U12649 (N_12649,N_10014,N_11429);
or U12650 (N_12650,N_10981,N_12348);
nand U12651 (N_12651,N_10488,N_10755);
xnor U12652 (N_12652,N_10790,N_11352);
xnor U12653 (N_12653,N_11668,N_10570);
xor U12654 (N_12654,N_11587,N_11233);
and U12655 (N_12655,N_11825,N_10627);
nand U12656 (N_12656,N_12218,N_11604);
and U12657 (N_12657,N_12414,N_11526);
and U12658 (N_12658,N_11438,N_11032);
or U12659 (N_12659,N_11116,N_10006);
or U12660 (N_12660,N_12426,N_11185);
nand U12661 (N_12661,N_10587,N_11357);
or U12662 (N_12662,N_11412,N_11295);
nand U12663 (N_12663,N_10394,N_10428);
xor U12664 (N_12664,N_12429,N_12424);
and U12665 (N_12665,N_12261,N_12055);
or U12666 (N_12666,N_10580,N_10839);
xor U12667 (N_12667,N_10581,N_11709);
xor U12668 (N_12668,N_12359,N_12379);
nor U12669 (N_12669,N_11939,N_12137);
nor U12670 (N_12670,N_10187,N_10167);
nor U12671 (N_12671,N_11111,N_10737);
and U12672 (N_12672,N_10044,N_11095);
xor U12673 (N_12673,N_11905,N_12254);
nand U12674 (N_12674,N_11957,N_11670);
or U12675 (N_12675,N_11439,N_10340);
and U12676 (N_12676,N_10619,N_10838);
nand U12677 (N_12677,N_11419,N_10886);
nor U12678 (N_12678,N_10674,N_10844);
nand U12679 (N_12679,N_11030,N_11776);
nor U12680 (N_12680,N_11818,N_10121);
nand U12681 (N_12681,N_10726,N_10050);
nand U12682 (N_12682,N_10114,N_11353);
or U12683 (N_12683,N_12085,N_10625);
or U12684 (N_12684,N_12070,N_10773);
or U12685 (N_12685,N_10590,N_11528);
nor U12686 (N_12686,N_10742,N_10450);
xor U12687 (N_12687,N_11612,N_10129);
and U12688 (N_12688,N_12230,N_10618);
xor U12689 (N_12689,N_12006,N_10232);
xnor U12690 (N_12690,N_11309,N_12313);
xor U12691 (N_12691,N_11935,N_10408);
nor U12692 (N_12692,N_12051,N_11930);
xor U12693 (N_12693,N_11836,N_12498);
or U12694 (N_12694,N_10180,N_11853);
nand U12695 (N_12695,N_10778,N_10263);
nor U12696 (N_12696,N_11740,N_11679);
and U12697 (N_12697,N_10221,N_10961);
nor U12698 (N_12698,N_11248,N_10923);
nand U12699 (N_12699,N_10182,N_11968);
and U12700 (N_12700,N_12434,N_12269);
nand U12701 (N_12701,N_12328,N_11008);
or U12702 (N_12702,N_11727,N_10881);
or U12703 (N_12703,N_12296,N_11724);
nor U12704 (N_12704,N_11786,N_11846);
and U12705 (N_12705,N_11743,N_10254);
or U12706 (N_12706,N_10370,N_10958);
nor U12707 (N_12707,N_10941,N_12141);
xnor U12708 (N_12708,N_10233,N_12444);
and U12709 (N_12709,N_11498,N_10700);
and U12710 (N_12710,N_12191,N_10592);
and U12711 (N_12711,N_11435,N_11719);
and U12712 (N_12712,N_10413,N_10975);
xor U12713 (N_12713,N_12086,N_12270);
and U12714 (N_12714,N_10548,N_10366);
or U12715 (N_12715,N_11854,N_11546);
nand U12716 (N_12716,N_12170,N_11243);
and U12717 (N_12717,N_10788,N_12396);
and U12718 (N_12718,N_10395,N_12084);
or U12719 (N_12719,N_10677,N_10361);
nor U12720 (N_12720,N_11377,N_10381);
and U12721 (N_12721,N_10703,N_10585);
xor U12722 (N_12722,N_10947,N_11103);
or U12723 (N_12723,N_11923,N_12076);
nor U12724 (N_12724,N_10308,N_11788);
nor U12725 (N_12725,N_11787,N_11593);
xor U12726 (N_12726,N_12169,N_10725);
or U12727 (N_12727,N_12449,N_12463);
xor U12728 (N_12728,N_11986,N_12178);
nor U12729 (N_12729,N_12455,N_11170);
xor U12730 (N_12730,N_10709,N_11254);
or U12731 (N_12731,N_10983,N_10995);
xnor U12732 (N_12732,N_11677,N_10083);
nand U12733 (N_12733,N_10637,N_12157);
xor U12734 (N_12734,N_11524,N_11859);
nand U12735 (N_12735,N_12204,N_12024);
and U12736 (N_12736,N_12435,N_11251);
nand U12737 (N_12737,N_12462,N_10678);
or U12738 (N_12738,N_12198,N_11810);
or U12739 (N_12739,N_11441,N_11468);
nor U12740 (N_12740,N_10926,N_12173);
and U12741 (N_12741,N_11898,N_11463);
and U12742 (N_12742,N_10069,N_10807);
nand U12743 (N_12743,N_10702,N_10097);
nor U12744 (N_12744,N_10942,N_11094);
and U12745 (N_12745,N_11652,N_10549);
xnor U12746 (N_12746,N_10294,N_10816);
or U12747 (N_12747,N_10203,N_11282);
and U12748 (N_12748,N_11025,N_12063);
nand U12749 (N_12749,N_12326,N_10606);
and U12750 (N_12750,N_11039,N_12389);
nor U12751 (N_12751,N_10039,N_11004);
nand U12752 (N_12752,N_12111,N_10347);
nand U12753 (N_12753,N_10032,N_11914);
and U12754 (N_12754,N_10136,N_10713);
and U12755 (N_12755,N_11843,N_11566);
and U12756 (N_12756,N_10887,N_11019);
nand U12757 (N_12757,N_10669,N_10655);
or U12758 (N_12758,N_10400,N_12219);
nor U12759 (N_12759,N_12171,N_10139);
and U12760 (N_12760,N_10165,N_10064);
and U12761 (N_12761,N_10665,N_11746);
xor U12762 (N_12762,N_10599,N_11916);
xnor U12763 (N_12763,N_12215,N_12217);
nor U12764 (N_12764,N_11635,N_10118);
xor U12765 (N_12765,N_12182,N_12321);
or U12766 (N_12766,N_12210,N_12019);
nor U12767 (N_12767,N_10506,N_11394);
nand U12768 (N_12768,N_11423,N_10927);
or U12769 (N_12769,N_10989,N_11430);
nand U12770 (N_12770,N_11347,N_10010);
or U12771 (N_12771,N_10646,N_12257);
nor U12772 (N_12772,N_11645,N_11304);
or U12773 (N_12773,N_12467,N_11698);
or U12774 (N_12774,N_12083,N_11637);
and U12775 (N_12775,N_12387,N_12186);
nand U12776 (N_12776,N_11121,N_10345);
xnor U12777 (N_12777,N_12452,N_10896);
nor U12778 (N_12778,N_11545,N_11639);
nand U12779 (N_12779,N_10225,N_10324);
nand U12780 (N_12780,N_10798,N_12487);
nand U12781 (N_12781,N_11560,N_11872);
xnor U12782 (N_12782,N_11945,N_11176);
nand U12783 (N_12783,N_10668,N_11433);
and U12784 (N_12784,N_11915,N_10623);
xor U12785 (N_12785,N_10567,N_10951);
nand U12786 (N_12786,N_11360,N_10293);
or U12787 (N_12787,N_12106,N_11559);
and U12788 (N_12788,N_10489,N_11663);
nand U12789 (N_12789,N_10505,N_11487);
xor U12790 (N_12790,N_12479,N_11206);
and U12791 (N_12791,N_11135,N_12029);
and U12792 (N_12792,N_10418,N_10214);
or U12793 (N_12793,N_12206,N_11625);
nand U12794 (N_12794,N_10174,N_11200);
xnor U12795 (N_12795,N_10374,N_11144);
nor U12796 (N_12796,N_11778,N_11301);
or U12797 (N_12797,N_11707,N_10043);
and U12798 (N_12798,N_11693,N_11926);
or U12799 (N_12799,N_10339,N_11061);
xnor U12800 (N_12800,N_11948,N_11310);
or U12801 (N_12801,N_10586,N_12004);
or U12802 (N_12802,N_11177,N_12130);
and U12803 (N_12803,N_10212,N_12382);
or U12804 (N_12804,N_11045,N_11594);
nand U12805 (N_12805,N_11232,N_11043);
nand U12806 (N_12806,N_11149,N_10150);
and U12807 (N_12807,N_11864,N_10155);
nand U12808 (N_12808,N_11443,N_11488);
nor U12809 (N_12809,N_11501,N_11107);
or U12810 (N_12810,N_11784,N_11580);
xnor U12811 (N_12811,N_11782,N_10264);
and U12812 (N_12812,N_10797,N_10888);
xor U12813 (N_12813,N_10904,N_11199);
and U12814 (N_12814,N_10893,N_10234);
and U12815 (N_12815,N_11797,N_11422);
and U12816 (N_12816,N_11431,N_10055);
nand U12817 (N_12817,N_10704,N_12159);
nor U12818 (N_12818,N_10494,N_11671);
and U12819 (N_12819,N_11253,N_10722);
nand U12820 (N_12820,N_10023,N_10138);
nor U12821 (N_12821,N_10119,N_10107);
and U12822 (N_12822,N_12319,N_12152);
or U12823 (N_12823,N_10243,N_11610);
nand U12824 (N_12824,N_10905,N_12233);
nand U12825 (N_12825,N_12318,N_10159);
and U12826 (N_12826,N_12197,N_10170);
nand U12827 (N_12827,N_11221,N_11770);
and U12828 (N_12828,N_11553,N_11075);
nand U12829 (N_12829,N_11122,N_10663);
xnor U12830 (N_12830,N_11150,N_11570);
or U12831 (N_12831,N_10579,N_12499);
nor U12832 (N_12832,N_11499,N_10152);
xor U12833 (N_12833,N_10818,N_10215);
nor U12834 (N_12834,N_10082,N_10157);
and U12835 (N_12835,N_12041,N_12489);
nand U12836 (N_12836,N_11131,N_10634);
nor U12837 (N_12837,N_11456,N_10186);
or U12838 (N_12838,N_11117,N_11665);
xnor U12839 (N_12839,N_11583,N_11870);
nand U12840 (N_12840,N_11829,N_12300);
nand U12841 (N_12841,N_10769,N_10456);
or U12842 (N_12842,N_12110,N_10588);
xor U12843 (N_12843,N_10382,N_10036);
nand U12844 (N_12844,N_10348,N_10598);
nor U12845 (N_12845,N_12145,N_10701);
and U12846 (N_12846,N_12108,N_10681);
or U12847 (N_12847,N_12393,N_10086);
or U12848 (N_12848,N_10156,N_11855);
xnor U12849 (N_12849,N_11392,N_11434);
nand U12850 (N_12850,N_11980,N_12294);
nor U12851 (N_12851,N_10379,N_11344);
nand U12852 (N_12852,N_10528,N_10323);
nand U12853 (N_12853,N_10142,N_10392);
nor U12854 (N_12854,N_10181,N_10582);
or U12855 (N_12855,N_12453,N_10992);
nand U12856 (N_12856,N_12026,N_11406);
xnor U12857 (N_12857,N_10209,N_12401);
nor U12858 (N_12858,N_10390,N_10829);
nor U12859 (N_12859,N_12419,N_11078);
nor U12860 (N_12860,N_12439,N_11837);
nand U12861 (N_12861,N_11571,N_12114);
nor U12862 (N_12862,N_11619,N_10442);
xnor U12863 (N_12863,N_10782,N_10486);
nor U12864 (N_12864,N_12079,N_10973);
nor U12865 (N_12865,N_10502,N_12161);
nand U12866 (N_12866,N_10422,N_11832);
nor U12867 (N_12867,N_11190,N_10688);
nand U12868 (N_12868,N_10879,N_10780);
nor U12869 (N_12869,N_12365,N_10539);
xor U12870 (N_12870,N_10643,N_10980);
or U12871 (N_12871,N_10612,N_11729);
and U12872 (N_12872,N_11067,N_11889);
or U12873 (N_12873,N_10049,N_10103);
xnor U12874 (N_12874,N_11226,N_11324);
nor U12875 (N_12875,N_10747,N_12408);
xnor U12876 (N_12876,N_11692,N_12285);
and U12877 (N_12877,N_10020,N_12043);
nand U12878 (N_12878,N_10393,N_12459);
nor U12879 (N_12879,N_10033,N_12388);
xnor U12880 (N_12880,N_11471,N_11910);
or U12881 (N_12881,N_10076,N_10998);
nand U12882 (N_12882,N_12391,N_10785);
nor U12883 (N_12883,N_11066,N_10237);
nor U12884 (N_12884,N_11082,N_10787);
or U12885 (N_12885,N_12018,N_10806);
or U12886 (N_12886,N_12017,N_12211);
and U12887 (N_12887,N_10994,N_11093);
or U12888 (N_12888,N_10657,N_10196);
nand U12889 (N_12889,N_12371,N_12027);
and U12890 (N_12890,N_11895,N_11849);
and U12891 (N_12891,N_11005,N_12199);
and U12892 (N_12892,N_11947,N_10759);
nor U12893 (N_12893,N_12179,N_11425);
nor U12894 (N_12894,N_11115,N_10963);
xor U12895 (N_12895,N_10265,N_10060);
nor U12896 (N_12896,N_11288,N_12375);
nand U12897 (N_12897,N_12331,N_11827);
xor U12898 (N_12898,N_10120,N_12174);
nor U12899 (N_12899,N_11051,N_12036);
or U12900 (N_12900,N_10822,N_12202);
xor U12901 (N_12901,N_11291,N_10177);
or U12902 (N_12902,N_12222,N_11048);
nor U12903 (N_12903,N_11276,N_11563);
nand U12904 (N_12904,N_11646,N_10429);
xnor U12905 (N_12905,N_11678,N_11494);
nor U12906 (N_12906,N_12010,N_12400);
xor U12907 (N_12907,N_12150,N_12088);
and U12908 (N_12908,N_10711,N_10401);
and U12909 (N_12909,N_11821,N_11766);
xor U12910 (N_12910,N_11602,N_11882);
nand U12911 (N_12911,N_10112,N_11712);
nor U12912 (N_12912,N_12436,N_11249);
nand U12913 (N_12913,N_10594,N_10559);
or U12914 (N_12914,N_11358,N_11942);
nand U12915 (N_12915,N_10949,N_11953);
nor U12916 (N_12916,N_11230,N_12203);
nand U12917 (N_12917,N_12207,N_11245);
and U12918 (N_12918,N_10641,N_10460);
or U12919 (N_12919,N_11934,N_11259);
nor U12920 (N_12920,N_12160,N_10168);
or U12921 (N_12921,N_12370,N_10783);
nor U12922 (N_12922,N_12445,N_10411);
and U12923 (N_12923,N_10868,N_11919);
or U12924 (N_12924,N_10132,N_12236);
or U12925 (N_12925,N_10096,N_11012);
xnor U12926 (N_12926,N_12165,N_11018);
nor U12927 (N_12927,N_11750,N_10013);
or U12928 (N_12928,N_12028,N_11857);
nor U12929 (N_12929,N_10380,N_11510);
and U12930 (N_12930,N_11816,N_10228);
or U12931 (N_12931,N_11197,N_12000);
xor U12932 (N_12932,N_10451,N_11072);
xnor U12933 (N_12933,N_10770,N_11447);
xnor U12934 (N_12934,N_12395,N_12302);
nand U12935 (N_12935,N_10877,N_11405);
xor U12936 (N_12936,N_12056,N_11186);
or U12937 (N_12937,N_12047,N_11466);
or U12938 (N_12938,N_10518,N_11541);
nand U12939 (N_12939,N_10303,N_11015);
or U12940 (N_12940,N_11623,N_12188);
xor U12941 (N_12941,N_11641,N_10289);
or U12942 (N_12942,N_12275,N_11314);
xor U12943 (N_12943,N_10301,N_10903);
xnor U12944 (N_12944,N_11806,N_10145);
xor U12945 (N_12945,N_11256,N_10122);
nand U12946 (N_12946,N_12443,N_11756);
xor U12947 (N_12947,N_11076,N_12460);
and U12948 (N_12948,N_10151,N_10048);
and U12949 (N_12949,N_11845,N_11955);
or U12950 (N_12950,N_12122,N_10406);
and U12951 (N_12951,N_11640,N_12129);
nor U12952 (N_12952,N_11329,N_12101);
nand U12953 (N_12953,N_10041,N_10734);
xnor U12954 (N_12954,N_11717,N_12213);
or U12955 (N_12955,N_11280,N_12229);
or U12956 (N_12956,N_11054,N_11588);
nor U12957 (N_12957,N_11193,N_10706);
xor U12958 (N_12958,N_10088,N_10464);
nor U12959 (N_12959,N_10837,N_11210);
nor U12960 (N_12960,N_11852,N_10326);
and U12961 (N_12961,N_10477,N_10661);
or U12962 (N_12962,N_10946,N_11042);
and U12963 (N_12963,N_12461,N_12472);
and U12964 (N_12964,N_11263,N_11516);
or U12965 (N_12965,N_10953,N_11356);
xnor U12966 (N_12966,N_11633,N_11191);
nand U12967 (N_12967,N_11047,N_11317);
or U12968 (N_12968,N_12335,N_12094);
xnor U12969 (N_12969,N_10094,N_10840);
nand U12970 (N_12970,N_12337,N_10169);
xor U12971 (N_12971,N_12125,N_11970);
nand U12972 (N_12972,N_10042,N_12358);
and U12973 (N_12973,N_11536,N_12340);
or U12974 (N_12974,N_10633,N_11537);
and U12975 (N_12975,N_11772,N_11550);
nand U12976 (N_12976,N_12220,N_10322);
and U12977 (N_12977,N_11653,N_10194);
and U12978 (N_12978,N_12067,N_10784);
xor U12979 (N_12979,N_11708,N_12205);
nor U12980 (N_12980,N_10235,N_12409);
nand U12981 (N_12981,N_10848,N_12080);
nand U12982 (N_12982,N_10311,N_11542);
nor U12983 (N_12983,N_10106,N_12003);
or U12984 (N_12984,N_10948,N_11993);
xnor U12985 (N_12985,N_12410,N_12038);
nand U12986 (N_12986,N_12336,N_10371);
xor U12987 (N_12987,N_10735,N_12077);
nand U12988 (N_12988,N_11346,N_10555);
nor U12989 (N_12989,N_11631,N_12128);
nor U12990 (N_12990,N_12405,N_11390);
or U12991 (N_12991,N_10873,N_11361);
xnor U12992 (N_12992,N_10176,N_12404);
nand U12993 (N_12993,N_10079,N_10596);
and U12994 (N_12994,N_10462,N_11759);
xnor U12995 (N_12995,N_10457,N_11555);
xnor U12996 (N_12996,N_10478,N_11687);
and U12997 (N_12997,N_11613,N_10786);
nand U12998 (N_12998,N_11733,N_10740);
and U12999 (N_12999,N_11608,N_12185);
nand U13000 (N_13000,N_11507,N_10409);
nand U13001 (N_13001,N_11337,N_11844);
or U13002 (N_13002,N_11465,N_11383);
xnor U13003 (N_13003,N_12316,N_11913);
and U13004 (N_13004,N_12458,N_11217);
or U13005 (N_13005,N_11586,N_10332);
xnor U13006 (N_13006,N_10387,N_10680);
xor U13007 (N_13007,N_10158,N_10184);
and U13008 (N_13008,N_10416,N_12135);
nor U13009 (N_13009,N_11380,N_12425);
xor U13010 (N_13010,N_11449,N_12143);
xnor U13011 (N_13011,N_12314,N_11674);
nand U13012 (N_13012,N_11366,N_10052);
or U13013 (N_13013,N_11567,N_10835);
and U13014 (N_13014,N_10694,N_10117);
nor U13015 (N_13015,N_10527,N_11909);
and U13016 (N_13016,N_10346,N_11050);
xnor U13017 (N_13017,N_12357,N_10153);
nand U13018 (N_13018,N_11688,N_11742);
or U13019 (N_13019,N_11381,N_11486);
or U13020 (N_13020,N_11154,N_12305);
xnor U13021 (N_13021,N_10068,N_10656);
and U13022 (N_13022,N_12184,N_11162);
nand U13023 (N_13023,N_11860,N_10448);
nor U13024 (N_13024,N_10402,N_10917);
xnor U13025 (N_13025,N_10330,N_10705);
nand U13026 (N_13026,N_11908,N_10760);
nand U13027 (N_13027,N_10752,N_11219);
xnor U13028 (N_13028,N_11382,N_10131);
xnor U13029 (N_13029,N_11658,N_10046);
xnor U13030 (N_13030,N_12276,N_11178);
nor U13031 (N_13031,N_11917,N_11293);
or U13032 (N_13032,N_10075,N_10913);
or U13033 (N_13033,N_10271,N_10831);
or U13034 (N_13034,N_11180,N_11007);
nand U13035 (N_13035,N_10996,N_10373);
xor U13036 (N_13036,N_10410,N_11216);
or U13037 (N_13037,N_10240,N_11876);
xor U13038 (N_13038,N_11963,N_10419);
and U13039 (N_13039,N_10135,N_10222);
and U13040 (N_13040,N_10874,N_11595);
and U13041 (N_13041,N_11166,N_12064);
xor U13042 (N_13042,N_11063,N_12306);
and U13043 (N_13043,N_10960,N_10100);
and U13044 (N_13044,N_11342,N_12494);
nand U13045 (N_13045,N_10256,N_11861);
xor U13046 (N_13046,N_11139,N_11736);
nand U13047 (N_13047,N_12212,N_11685);
xor U13048 (N_13048,N_11683,N_11028);
xnor U13049 (N_13049,N_11747,N_10270);
xnor U13050 (N_13050,N_11643,N_11089);
and U13051 (N_13051,N_11814,N_11371);
and U13052 (N_13052,N_11630,N_11977);
xor U13053 (N_13053,N_10566,N_10557);
and U13054 (N_13054,N_12119,N_11393);
nand U13055 (N_13055,N_12423,N_10845);
or U13056 (N_13056,N_12034,N_12255);
nor U13057 (N_13057,N_12380,N_10716);
or U13058 (N_13058,N_11398,N_11819);
and U13059 (N_13059,N_10437,N_10248);
or U13060 (N_13060,N_10281,N_10147);
xor U13061 (N_13061,N_12065,N_11281);
and U13062 (N_13062,N_12251,N_10902);
nor U13063 (N_13063,N_12397,N_11462);
xor U13064 (N_13064,N_11086,N_10183);
xor U13065 (N_13065,N_11868,N_10423);
or U13066 (N_13066,N_10508,N_10891);
xor U13067 (N_13067,N_10745,N_12278);
and U13068 (N_13068,N_12155,N_10446);
or U13069 (N_13069,N_11803,N_11275);
xor U13070 (N_13070,N_10801,N_10172);
and U13071 (N_13071,N_10781,N_12324);
nand U13072 (N_13072,N_11053,N_11525);
nand U13073 (N_13073,N_11774,N_11350);
nor U13074 (N_13074,N_12023,N_11041);
nand U13075 (N_13075,N_12117,N_11765);
nor U13076 (N_13076,N_12267,N_11303);
or U13077 (N_13077,N_11482,N_10962);
or U13078 (N_13078,N_12105,N_12492);
and U13079 (N_13079,N_10642,N_11192);
nand U13080 (N_13080,N_11751,N_11557);
or U13081 (N_13081,N_11300,N_10404);
and U13082 (N_13082,N_10651,N_11762);
and U13083 (N_13083,N_10213,N_12090);
and U13084 (N_13084,N_12490,N_10935);
xor U13085 (N_13085,N_11710,N_11334);
and U13086 (N_13086,N_11937,N_12062);
nor U13087 (N_13087,N_11754,N_11598);
or U13088 (N_13088,N_11410,N_12442);
and U13089 (N_13089,N_10883,N_10342);
or U13090 (N_13090,N_10911,N_11027);
xnor U13091 (N_13091,N_10282,N_11472);
nor U13092 (N_13092,N_11305,N_12372);
xor U13093 (N_13093,N_10525,N_11723);
xor U13094 (N_13094,N_10639,N_11944);
nor U13095 (N_13095,N_10483,N_10589);
or U13096 (N_13096,N_10175,N_10660);
nand U13097 (N_13097,N_10693,N_10774);
nor U13098 (N_13098,N_12291,N_12454);
and U13099 (N_13099,N_10466,N_10480);
nor U13100 (N_13100,N_12447,N_10261);
xor U13101 (N_13101,N_10622,N_11605);
nor U13102 (N_13102,N_11218,N_10290);
nand U13103 (N_13103,N_10128,N_10743);
and U13104 (N_13104,N_11133,N_12097);
nor U13105 (N_13105,N_10236,N_11364);
and U13106 (N_13106,N_10856,N_11460);
or U13107 (N_13107,N_11212,N_12364);
xor U13108 (N_13108,N_11659,N_11058);
xor U13109 (N_13109,N_10384,N_11584);
and U13110 (N_13110,N_12354,N_10388);
xnor U13111 (N_13111,N_10855,N_10872);
and U13112 (N_13112,N_10540,N_10299);
nor U13113 (N_13113,N_11119,N_10550);
or U13114 (N_13114,N_12044,N_10921);
xnor U13115 (N_13115,N_10775,N_11530);
or U13116 (N_13116,N_12304,N_10601);
and U13117 (N_13117,N_11590,N_10426);
xor U13118 (N_13118,N_10939,N_11318);
or U13119 (N_13119,N_10149,N_12166);
and U13120 (N_13120,N_12073,N_10662);
nor U13121 (N_13121,N_10815,N_10964);
nand U13122 (N_13122,N_12249,N_11877);
nor U13123 (N_13123,N_11098,N_11974);
or U13124 (N_13124,N_11205,N_10111);
nand U13125 (N_13125,N_10524,N_12045);
nand U13126 (N_13126,N_11960,N_12383);
nor U13127 (N_13127,N_11675,N_11888);
nand U13128 (N_13128,N_11785,N_12158);
xor U13129 (N_13129,N_12020,N_11805);
nand U13130 (N_13130,N_10986,N_11938);
and U13131 (N_13131,N_10000,N_10173);
or U13132 (N_13132,N_12196,N_10966);
and U13133 (N_13133,N_11949,N_11173);
and U13134 (N_13134,N_11720,N_10613);
or U13135 (N_13135,N_10564,N_12098);
nor U13136 (N_13136,N_10968,N_10335);
and U13137 (N_13137,N_11368,N_10011);
xor U13138 (N_13138,N_11540,N_12406);
xnor U13139 (N_13139,N_12322,N_10284);
or U13140 (N_13140,N_12226,N_11480);
nor U13141 (N_13141,N_11582,N_11780);
xor U13142 (N_13142,N_10876,N_11880);
nand U13143 (N_13143,N_11547,N_11416);
and U13144 (N_13144,N_12466,N_11969);
nor U13145 (N_13145,N_11556,N_11009);
nor U13146 (N_13146,N_11229,N_12351);
and U13147 (N_13147,N_12407,N_11088);
nor U13148 (N_13148,N_10495,N_10313);
nor U13149 (N_13149,N_10830,N_12244);
or U13150 (N_13150,N_11681,N_11255);
nand U13151 (N_13151,N_10930,N_11184);
and U13152 (N_13152,N_11299,N_11552);
xnor U13153 (N_13153,N_10820,N_11512);
or U13154 (N_13154,N_10860,N_10472);
xor U13155 (N_13155,N_11629,N_10714);
xor U13156 (N_13156,N_10407,N_11049);
nand U13157 (N_13157,N_11673,N_11705);
xor U13158 (N_13158,N_12016,N_12245);
or U13159 (N_13159,N_10231,N_11316);
xor U13160 (N_13160,N_10556,N_11549);
nor U13161 (N_13161,N_10648,N_12310);
xor U13162 (N_13162,N_11348,N_11455);
or U13163 (N_13163,N_12428,N_10073);
xor U13164 (N_13164,N_10239,N_11984);
and U13165 (N_13165,N_12192,N_11822);
nand U13166 (N_13166,N_10353,N_10226);
and U13167 (N_13167,N_10638,N_10260);
xnor U13168 (N_13168,N_11322,N_10253);
xnor U13169 (N_13169,N_11521,N_10597);
nor U13170 (N_13170,N_10123,N_11424);
xnor U13171 (N_13171,N_11246,N_10800);
nand U13172 (N_13172,N_10616,N_11461);
nor U13173 (N_13173,N_12430,N_10171);
and U13174 (N_13174,N_10443,N_11375);
nor U13175 (N_13175,N_12496,N_10219);
nor U13176 (N_13176,N_12250,N_10794);
xnor U13177 (N_13177,N_10554,N_10360);
nand U13178 (N_13178,N_10059,N_11509);
nor U13179 (N_13179,N_11691,N_12398);
xnor U13180 (N_13180,N_10575,N_12201);
nand U13181 (N_13181,N_10766,N_12100);
xnor U13182 (N_13182,N_12247,N_10018);
nor U13183 (N_13183,N_11900,N_11147);
xnor U13184 (N_13184,N_11793,N_10919);
and U13185 (N_13185,N_11985,N_12486);
nand U13186 (N_13186,N_10389,N_11867);
and U13187 (N_13187,N_12344,N_11181);
xnor U13188 (N_13188,N_10115,N_10045);
nor U13189 (N_13189,N_11378,N_11730);
nand U13190 (N_13190,N_10433,N_11420);
or U13191 (N_13191,N_10696,N_12099);
xor U13192 (N_13192,N_10685,N_11208);
nand U13193 (N_13193,N_11715,N_10636);
nand U13194 (N_13194,N_10841,N_12438);
nor U13195 (N_13195,N_10016,N_12471);
or U13196 (N_13196,N_11427,N_12163);
nor U13197 (N_13197,N_10449,N_10732);
and U13198 (N_13198,N_12120,N_11551);
nor U13199 (N_13199,N_11138,N_11885);
nand U13200 (N_13200,N_10189,N_11731);
and U13201 (N_13201,N_10629,N_10160);
nor U13202 (N_13202,N_10255,N_11077);
and U13203 (N_13203,N_10081,N_11734);
nand U13204 (N_13204,N_10878,N_11313);
or U13205 (N_13205,N_10982,N_11656);
nand U13206 (N_13206,N_10934,N_12035);
nor U13207 (N_13207,N_11978,N_11016);
nor U13208 (N_13208,N_12172,N_12058);
nor U13209 (N_13209,N_11479,N_12107);
and U13210 (N_13210,N_11958,N_11896);
or U13211 (N_13211,N_12448,N_11143);
or U13212 (N_13212,N_10916,N_11437);
nor U13213 (N_13213,N_12298,N_11323);
xor U13214 (N_13214,N_11865,N_10659);
nand U13215 (N_13215,N_11911,N_10095);
nand U13216 (N_13216,N_10166,N_10811);
nor U13217 (N_13217,N_10190,N_11272);
or U13218 (N_13218,N_10337,N_10628);
nand U13219 (N_13219,N_10521,N_11798);
or U13220 (N_13220,N_10071,N_11114);
xnor U13221 (N_13221,N_11395,N_10940);
nand U13222 (N_13222,N_12470,N_10687);
xnor U13223 (N_13223,N_10216,N_10715);
nor U13224 (N_13224,N_10805,N_12368);
or U13225 (N_13225,N_12422,N_10431);
nor U13226 (N_13226,N_10350,N_12127);
xnor U13227 (N_13227,N_10162,N_11666);
nor U13228 (N_13228,N_11262,N_11811);
or U13229 (N_13229,N_11807,N_10316);
nor U13230 (N_13230,N_11389,N_11385);
xnor U13231 (N_13231,N_10072,N_11952);
or U13232 (N_13232,N_10029,N_12069);
or U13233 (N_13233,N_11321,N_10414);
and U13234 (N_13234,N_12292,N_10412);
nand U13235 (N_13235,N_10479,N_11179);
nand U13236 (N_13236,N_11183,N_12446);
nand U13237 (N_13237,N_10130,N_11753);
nand U13238 (N_13238,N_12007,N_11874);
xor U13239 (N_13239,N_11642,N_10537);
nand U13240 (N_13240,N_10277,N_11172);
nor U13241 (N_13241,N_11129,N_11738);
or U13242 (N_13242,N_11614,N_10900);
and U13243 (N_13243,N_11446,N_12350);
nor U13244 (N_13244,N_11981,N_10803);
xnor U13245 (N_13245,N_12046,N_11890);
nor U13246 (N_13246,N_12273,N_11023);
or U13247 (N_13247,N_10372,N_10810);
nand U13248 (N_13248,N_10438,N_12412);
or U13249 (N_13249,N_12183,N_11628);
and U13250 (N_13250,N_11725,N_12288);
or U13251 (N_13251,N_10019,N_12325);
nor U13252 (N_13252,N_10470,N_12282);
nor U13253 (N_13253,N_11330,N_10468);
nor U13254 (N_13254,N_10328,N_11539);
or U13255 (N_13255,N_10427,N_11922);
nor U13256 (N_13256,N_11779,N_10611);
or U13257 (N_13257,N_10558,N_11634);
or U13258 (N_13258,N_11307,N_12272);
xor U13259 (N_13259,N_10492,N_11809);
xor U13260 (N_13260,N_12146,N_10503);
nand U13261 (N_13261,N_11174,N_11791);
nor U13262 (N_13262,N_11268,N_12071);
nor U13263 (N_13263,N_11669,N_10978);
xor U13264 (N_13264,N_11354,N_10875);
and U13265 (N_13265,N_12346,N_12059);
xnor U13266 (N_13266,N_10791,N_12239);
xor U13267 (N_13267,N_10776,N_11992);
or U13268 (N_13268,N_10546,N_10571);
and U13269 (N_13269,N_11768,N_11029);
nor U13270 (N_13270,N_12136,N_10568);
or U13271 (N_13271,N_11167,N_11343);
xnor U13272 (N_13272,N_10474,N_10652);
nand U13273 (N_13273,N_10880,N_10430);
xor U13274 (N_13274,N_10320,N_10202);
or U13275 (N_13275,N_10024,N_10718);
nand U13276 (N_13276,N_12033,N_10224);
nor U13277 (N_13277,N_12246,N_12195);
nand U13278 (N_13278,N_10292,N_10475);
and U13279 (N_13279,N_11484,N_10918);
nor U13280 (N_13280,N_11792,N_10569);
nand U13281 (N_13281,N_10733,N_10063);
nor U13282 (N_13282,N_12482,N_11824);
nor U13283 (N_13283,N_10283,N_11573);
and U13284 (N_13284,N_12240,N_11987);
xor U13285 (N_13285,N_11554,N_10109);
and U13286 (N_13286,N_10812,N_10833);
and U13287 (N_13287,N_10908,N_10542);
and U13288 (N_13288,N_10327,N_11728);
xnor U13289 (N_13289,N_10543,N_10454);
or U13290 (N_13290,N_10920,N_12366);
xor U13291 (N_13291,N_11664,N_11187);
xnor U13292 (N_13292,N_10329,N_11535);
xor U13293 (N_13293,N_11879,N_10420);
nor U13294 (N_13294,N_10004,N_10898);
nor U13295 (N_13295,N_11982,N_11618);
and U13296 (N_13296,N_11286,N_11839);
nor U13297 (N_13297,N_10280,N_12334);
and U13298 (N_13298,N_11038,N_10676);
or U13299 (N_13299,N_12014,N_11695);
and U13300 (N_13300,N_10259,N_10901);
and U13301 (N_13301,N_11769,N_10970);
and U13302 (N_13302,N_10533,N_12216);
xnor U13303 (N_13303,N_12048,N_12457);
nor U13304 (N_13304,N_12234,N_11396);
xnor U13305 (N_13305,N_10515,N_10312);
or U13306 (N_13306,N_10796,N_10485);
nand U13307 (N_13307,N_12451,N_11024);
xnor U13308 (N_13308,N_12039,N_11428);
nor U13309 (N_13309,N_11426,N_10507);
and U13310 (N_13310,N_11081,N_12095);
nand U13311 (N_13311,N_11214,N_11369);
nand U13312 (N_13312,N_10777,N_11153);
nand U13313 (N_13313,N_11817,N_11296);
nor U13314 (N_13314,N_12209,N_11513);
nand U13315 (N_13315,N_11840,N_10631);
nand U13316 (N_13316,N_10754,N_12441);
or U13317 (N_13317,N_11267,N_11037);
xor U13318 (N_13318,N_10836,N_11833);
nor U13319 (N_13319,N_11831,N_10574);
and U13320 (N_13320,N_10101,N_10545);
and U13321 (N_13321,N_12297,N_11448);
and U13322 (N_13322,N_10383,N_10099);
and U13323 (N_13323,N_10038,N_11489);
xor U13324 (N_13324,N_10436,N_11247);
or U13325 (N_13325,N_11370,N_10125);
or U13326 (N_13326,N_10724,N_10223);
or U13327 (N_13327,N_10553,N_10653);
nand U13328 (N_13328,N_11596,N_12138);
xnor U13329 (N_13329,N_11518,N_11469);
xor U13330 (N_13330,N_12473,N_10021);
or U13331 (N_13331,N_11126,N_11068);
nand U13332 (N_13332,N_11475,N_10744);
and U13333 (N_13333,N_12012,N_12237);
nor U13334 (N_13334,N_11983,N_11607);
nor U13335 (N_13335,N_10317,N_11236);
nor U13336 (N_13336,N_10707,N_11224);
or U13337 (N_13337,N_11070,N_10988);
xnor U13338 (N_13338,N_11132,N_11764);
nand U13339 (N_13339,N_10847,N_11033);
xor U13340 (N_13340,N_12376,N_10296);
nand U13341 (N_13341,N_11040,N_11718);
nand U13342 (N_13342,N_10285,N_11340);
xor U13343 (N_13343,N_10465,N_11662);
nand U13344 (N_13344,N_10832,N_10859);
nor U13345 (N_13345,N_10600,N_11886);
nand U13346 (N_13346,N_10309,N_10241);
nor U13347 (N_13347,N_11932,N_12286);
and U13348 (N_13348,N_11379,N_11222);
and U13349 (N_13349,N_12180,N_10910);
or U13350 (N_13350,N_11384,N_11097);
and U13351 (N_13351,N_10952,N_10813);
and U13352 (N_13352,N_11976,N_12081);
xor U13353 (N_13353,N_11238,N_12403);
and U13354 (N_13354,N_10690,N_10272);
nand U13355 (N_13355,N_12005,N_10461);
nor U13356 (N_13356,N_11600,N_12312);
nand U13357 (N_13357,N_11505,N_11741);
nor U13358 (N_13358,N_11936,N_10757);
and U13359 (N_13359,N_11477,N_12243);
or U13360 (N_13360,N_10359,N_11994);
xor U13361 (N_13361,N_11113,N_10291);
nor U13362 (N_13362,N_11349,N_10670);
nor U13363 (N_13363,N_12262,N_11964);
nand U13364 (N_13364,N_11289,N_12089);
nand U13365 (N_13365,N_10257,N_10608);
nor U13366 (N_13366,N_11585,N_11458);
nor U13367 (N_13367,N_12287,N_11101);
and U13368 (N_13368,N_10814,N_10362);
or U13369 (N_13369,N_12082,N_11108);
xnor U13370 (N_13370,N_10739,N_12113);
xnor U13371 (N_13371,N_10035,N_10375);
nand U13372 (N_13372,N_10487,N_12476);
and U13373 (N_13373,N_10697,N_11823);
nor U13374 (N_13374,N_11562,N_11568);
nor U13375 (N_13375,N_11940,N_11997);
and U13376 (N_13376,N_10008,N_10098);
or U13377 (N_13377,N_11760,N_10595);
and U13378 (N_13378,N_11175,N_11271);
nor U13379 (N_13379,N_11878,N_11838);
nor U13380 (N_13380,N_10302,N_11667);
xnor U13381 (N_13381,N_11862,N_10609);
xnor U13382 (N_13382,N_10541,N_11869);
or U13383 (N_13383,N_11726,N_10217);
xor U13384 (N_13384,N_12074,N_10025);
and U13385 (N_13385,N_10134,N_11328);
nand U13386 (N_13386,N_11907,N_11336);
and U13387 (N_13387,N_11802,N_11655);
or U13388 (N_13388,N_10493,N_10315);
nor U13389 (N_13389,N_10331,N_11158);
or U13390 (N_13390,N_12176,N_10565);
or U13391 (N_13391,N_12032,N_10602);
and U13392 (N_13392,N_12190,N_11749);
nor U13393 (N_13393,N_10710,N_10925);
and U13394 (N_13394,N_11661,N_11609);
or U13395 (N_13395,N_12187,N_10649);
nor U13396 (N_13396,N_11490,N_10343);
or U13397 (N_13397,N_11136,N_11773);
xnor U13398 (N_13398,N_11194,N_11901);
xor U13399 (N_13399,N_12259,N_11775);
nor U13400 (N_13400,N_11235,N_12485);
xor U13401 (N_13401,N_11404,N_10246);
nor U13402 (N_13402,N_10022,N_12252);
and U13403 (N_13403,N_11495,N_11403);
nor U13404 (N_13404,N_10675,N_10199);
and U13405 (N_13405,N_10247,N_11234);
nand U13406 (N_13406,N_10666,N_10085);
or U13407 (N_13407,N_10040,N_11085);
nor U13408 (N_13408,N_10325,N_11891);
and U13409 (N_13409,N_12068,N_10767);
nand U13410 (N_13410,N_10459,N_10809);
or U13411 (N_13411,N_11099,N_11283);
nor U13412 (N_13412,N_11597,N_12194);
nor U13413 (N_13413,N_12279,N_10937);
nor U13414 (N_13414,N_10615,N_10496);
or U13415 (N_13415,N_10993,N_10610);
or U13416 (N_13416,N_10884,N_11702);
xor U13417 (N_13417,N_11574,N_12308);
xnor U13418 (N_13418,N_11156,N_11694);
xnor U13419 (N_13419,N_10206,N_10824);
and U13420 (N_13420,N_10929,N_12338);
xnor U13421 (N_13421,N_10808,N_10058);
xor U13422 (N_13422,N_11165,N_11014);
xor U13423 (N_13423,N_10369,N_10862);
or U13424 (N_13424,N_11706,N_12315);
or U13425 (N_13425,N_11452,N_11603);
nand U13426 (N_13426,N_11060,N_11956);
and U13427 (N_13427,N_10396,N_10274);
xor U13428 (N_13428,N_10484,N_12483);
xnor U13429 (N_13429,N_12103,N_10719);
and U13430 (N_13430,N_11003,N_10047);
and U13431 (N_13431,N_11820,N_12167);
or U13432 (N_13432,N_10852,N_12341);
xor U13433 (N_13433,N_10861,N_10795);
nand U13434 (N_13434,N_10821,N_11306);
nand U13435 (N_13435,N_12274,N_10276);
or U13436 (N_13436,N_11951,N_11577);
and U13437 (N_13437,N_11763,N_10210);
or U13438 (N_13438,N_12121,N_11444);
nor U13439 (N_13439,N_12417,N_11312);
nor U13440 (N_13440,N_11141,N_11591);
nor U13441 (N_13441,N_10238,N_11450);
nand U13442 (N_13442,N_10799,N_12421);
xor U13443 (N_13443,N_12497,N_11481);
nor U13444 (N_13444,N_11519,N_11064);
nand U13445 (N_13445,N_10363,N_10278);
and U13446 (N_13446,N_10144,N_11010);
xor U13447 (N_13447,N_11168,N_10482);
nor U13448 (N_13448,N_10307,N_10621);
and U13449 (N_13449,N_10991,N_12242);
or U13450 (N_13450,N_10007,N_12381);
nor U13451 (N_13451,N_10204,N_10971);
or U13452 (N_13452,N_10230,N_12349);
nor U13453 (N_13453,N_10846,N_10727);
nand U13454 (N_13454,N_11716,N_10909);
nand U13455 (N_13455,N_10603,N_10604);
nand U13456 (N_13456,N_11483,N_11569);
xnor U13457 (N_13457,N_10728,N_10056);
xnor U13458 (N_13458,N_11290,N_10731);
xnor U13459 (N_13459,N_10933,N_11250);
xor U13460 (N_13460,N_10895,N_10976);
nor U13461 (N_13461,N_10990,N_11575);
xor U13462 (N_13462,N_11228,N_12290);
nor U13463 (N_13463,N_10584,N_11690);
xnor U13464 (N_13464,N_10956,N_11493);
nor U13465 (N_13465,N_10354,N_12140);
nor U13466 (N_13466,N_12362,N_10712);
nand U13467 (N_13467,N_10577,N_11924);
or U13468 (N_13468,N_10758,N_12109);
nor U13469 (N_13469,N_11418,N_11470);
nand U13470 (N_13470,N_11752,N_11453);
or U13471 (N_13471,N_11884,N_11140);
nand U13472 (N_13472,N_10378,N_11961);
and U13473 (N_13473,N_10074,N_10640);
nand U13474 (N_13474,N_10065,N_10164);
xor U13475 (N_13475,N_10067,N_11704);
or U13476 (N_13476,N_10273,N_10869);
xnor U13477 (N_13477,N_10385,N_11904);
and U13478 (N_13478,N_12374,N_10721);
nand U13479 (N_13479,N_12151,N_10218);
nor U13480 (N_13480,N_11906,N_11223);
or U13481 (N_13481,N_10364,N_10538);
xor U13482 (N_13482,N_12263,N_10885);
xnor U13483 (N_13483,N_11971,N_10338);
nor U13484 (N_13484,N_12223,N_10447);
xnor U13485 (N_13485,N_11408,N_11367);
or U13486 (N_13486,N_10654,N_10333);
and U13487 (N_13487,N_12415,N_10090);
and U13488 (N_13488,N_11372,N_10027);
nand U13489 (N_13489,N_10092,N_10425);
and U13490 (N_13490,N_12021,N_11735);
xnor U13491 (N_13491,N_11826,N_10686);
nand U13492 (N_13492,N_10915,N_10834);
nor U13493 (N_13493,N_10251,N_11298);
xor U13494 (N_13494,N_11073,N_12464);
nor U13495 (N_13495,N_11277,N_10526);
nor U13496 (N_13496,N_10467,N_11373);
nor U13497 (N_13497,N_12087,N_12333);
nor U13498 (N_13498,N_10455,N_10517);
nor U13499 (N_13499,N_11001,N_10854);
xor U13500 (N_13500,N_11160,N_10682);
nor U13501 (N_13501,N_11409,N_11325);
nand U13502 (N_13502,N_10476,N_12323);
nand U13503 (N_13503,N_11576,N_10154);
nand U13504 (N_13504,N_11391,N_10906);
nor U13505 (N_13505,N_10699,N_10738);
or U13506 (N_13506,N_11100,N_11858);
xnor U13507 (N_13507,N_10857,N_11699);
and U13508 (N_13508,N_12049,N_10954);
xnor U13509 (N_13509,N_12480,N_10635);
nor U13510 (N_13510,N_10536,N_11202);
xnor U13511 (N_13511,N_10720,N_12241);
xnor U13512 (N_13512,N_12124,N_11266);
nor U13513 (N_13513,N_11700,N_11397);
or U13514 (N_13514,N_10031,N_12144);
nand U13515 (N_13515,N_10516,N_11941);
nor U13516 (N_13516,N_11988,N_10469);
or U13517 (N_13517,N_11252,N_12390);
or U13518 (N_13518,N_12416,N_11812);
or U13519 (N_13519,N_11467,N_12367);
nand U13520 (N_13520,N_11813,N_11544);
and U13521 (N_13521,N_11883,N_10208);
nor U13522 (N_13522,N_10828,N_10889);
or U13523 (N_13523,N_10501,N_11261);
xor U13524 (N_13524,N_11451,N_10999);
nand U13525 (N_13525,N_11581,N_11387);
and U13526 (N_13526,N_10772,N_12050);
or U13527 (N_13527,N_12385,N_12363);
and U13528 (N_13528,N_12116,N_11841);
nor U13529 (N_13529,N_10053,N_10689);
xnor U13530 (N_13530,N_10441,N_11017);
and U13531 (N_13531,N_12013,N_12277);
or U13532 (N_13532,N_10358,N_12330);
or U13533 (N_13533,N_10552,N_10104);
and U13534 (N_13534,N_11163,N_11995);
nor U13535 (N_13535,N_12295,N_12311);
or U13536 (N_13536,N_12011,N_11954);
nor U13537 (N_13537,N_11091,N_12281);
nor U13538 (N_13538,N_11124,N_11459);
nand U13539 (N_13539,N_10334,N_11062);
or U13540 (N_13540,N_11302,N_12378);
and U13541 (N_13541,N_10520,N_10398);
xnor U13542 (N_13542,N_11338,N_10684);
and U13543 (N_13543,N_11473,N_12175);
nor U13544 (N_13544,N_10736,N_11504);
and U13545 (N_13545,N_10907,N_10779);
xor U13546 (N_13546,N_11808,N_10950);
nand U13547 (N_13547,N_12153,N_10078);
nand U13548 (N_13548,N_11415,N_10765);
and U13549 (N_13549,N_11866,N_12339);
and U13550 (N_13550,N_10193,N_11638);
xnor U13551 (N_13551,N_10110,N_11648);
or U13552 (N_13552,N_10723,N_11848);
xor U13553 (N_13553,N_11102,N_12054);
or U13554 (N_13554,N_11341,N_10624);
or U13555 (N_13555,N_10523,N_11929);
nor U13556 (N_13556,N_11801,N_11308);
xor U13557 (N_13557,N_11227,N_11531);
and U13558 (N_13558,N_11713,N_10899);
nand U13559 (N_13559,N_12214,N_12132);
or U13560 (N_13560,N_10762,N_11011);
nand U13561 (N_13561,N_11402,N_12384);
or U13562 (N_13562,N_10967,N_12392);
xnor U13563 (N_13563,N_10804,N_12360);
and U13564 (N_13564,N_11796,N_10583);
or U13565 (N_13565,N_12356,N_12488);
or U13566 (N_13566,N_10421,N_12258);
nor U13567 (N_13567,N_11558,N_11106);
xnor U13568 (N_13568,N_10304,N_10617);
or U13569 (N_13569,N_11514,N_11680);
xnor U13570 (N_13570,N_11928,N_11359);
nor U13571 (N_13571,N_10211,N_12134);
nor U13572 (N_13572,N_11026,N_11311);
and U13573 (N_13573,N_10658,N_11169);
nand U13574 (N_13574,N_10897,N_11118);
and U13575 (N_13575,N_11478,N_10620);
xnor U13576 (N_13576,N_11881,N_10827);
nor U13577 (N_13577,N_10026,N_10748);
and U13578 (N_13578,N_12177,N_10692);
or U13579 (N_13579,N_10453,N_10314);
nor U13580 (N_13580,N_10532,N_11758);
xnor U13581 (N_13581,N_10452,N_10853);
or U13582 (N_13582,N_11696,N_10977);
nand U13583 (N_13583,N_11975,N_11351);
or U13584 (N_13584,N_11457,N_10367);
nor U13585 (N_13585,N_11000,N_11979);
or U13586 (N_13586,N_11414,N_10671);
or U13587 (N_13587,N_11035,N_10077);
nor U13588 (N_13588,N_11260,N_10399);
and U13589 (N_13589,N_11748,N_11440);
xnor U13590 (N_13590,N_10997,N_11847);
xnor U13591 (N_13591,N_10341,N_10051);
xnor U13592 (N_13592,N_11335,N_10984);
nor U13593 (N_13593,N_12386,N_12053);
and U13594 (N_13594,N_11326,N_11624);
nand U13595 (N_13595,N_10245,N_10179);
nand U13596 (N_13596,N_12411,N_11084);
nand U13597 (N_13597,N_11532,N_10842);
and U13598 (N_13598,N_12112,N_12148);
and U13599 (N_13599,N_11647,N_11400);
nand U13600 (N_13600,N_11503,N_10944);
xor U13601 (N_13601,N_10849,N_10691);
xnor U13602 (N_13602,N_11112,N_10851);
xnor U13603 (N_13603,N_10305,N_10965);
or U13604 (N_13604,N_10057,N_11152);
nand U13605 (N_13605,N_10938,N_10667);
or U13606 (N_13606,N_12123,N_11339);
and U13607 (N_13607,N_11065,N_11496);
and U13608 (N_13608,N_10220,N_11676);
xnor U13609 (N_13609,N_12307,N_10377);
xnor U13610 (N_13610,N_11134,N_11578);
or U13611 (N_13611,N_10269,N_10356);
xnor U13612 (N_13612,N_12037,N_11204);
nand U13613 (N_13613,N_10250,N_10001);
or U13614 (N_13614,N_11835,N_11225);
xor U13615 (N_13615,N_11842,N_11933);
or U13616 (N_13616,N_11331,N_11851);
nand U13617 (N_13617,N_10945,N_10551);
nor U13618 (N_13618,N_11155,N_10573);
or U13619 (N_13619,N_11830,N_10087);
or U13620 (N_13620,N_12052,N_10969);
or U13621 (N_13621,N_11273,N_11087);
nor U13622 (N_13622,N_11617,N_11892);
and U13623 (N_13623,N_11781,N_11739);
nor U13624 (N_13624,N_11515,N_11771);
nor U13625 (N_13625,N_10562,N_10458);
or U13626 (N_13626,N_10163,N_12478);
or U13627 (N_13627,N_11355,N_10535);
xor U13628 (N_13628,N_10792,N_10892);
nand U13629 (N_13629,N_10192,N_11109);
xor U13630 (N_13630,N_11327,N_10632);
xnor U13631 (N_13631,N_11270,N_11800);
xor U13632 (N_13632,N_10066,N_12015);
xor U13633 (N_13633,N_12440,N_11239);
and U13634 (N_13634,N_12072,N_10650);
or U13635 (N_13635,N_10344,N_10463);
nand U13636 (N_13636,N_11492,N_12327);
or U13637 (N_13637,N_11850,N_11527);
and U13638 (N_13638,N_11130,N_12303);
xnor U13639 (N_13639,N_10197,N_10522);
xnor U13640 (N_13640,N_11240,N_10062);
xor U13641 (N_13641,N_11442,N_11074);
and U13642 (N_13642,N_10201,N_10200);
or U13643 (N_13643,N_12377,N_11943);
and U13644 (N_13644,N_10070,N_10297);
xor U13645 (N_13645,N_11783,N_11319);
xnor U13646 (N_13646,N_10397,N_11006);
nand U13647 (N_13647,N_12091,N_12361);
xor U13648 (N_13648,N_12126,N_10295);
and U13649 (N_13649,N_11973,N_11511);
or U13650 (N_13650,N_12142,N_11411);
xor U13651 (N_13651,N_11127,N_11767);
nor U13652 (N_13652,N_10124,N_10753);
nor U13653 (N_13653,N_12266,N_10514);
nand U13654 (N_13654,N_11538,N_10751);
or U13655 (N_13655,N_10914,N_12221);
xnor U13656 (N_13656,N_10306,N_10108);
xnor U13657 (N_13657,N_10764,N_11998);
nor U13658 (N_13658,N_12224,N_11636);
nor U13659 (N_13659,N_11873,N_11894);
nand U13660 (N_13660,N_12484,N_11474);
nand U13661 (N_13661,N_11795,N_12133);
nand U13662 (N_13662,N_10823,N_11213);
xor U13663 (N_13663,N_10310,N_11761);
xor U13664 (N_13664,N_11522,N_10882);
xor U13665 (N_13665,N_10593,N_11105);
or U13666 (N_13666,N_10133,N_10034);
nor U13667 (N_13667,N_10105,N_11146);
or U13668 (N_13668,N_12469,N_11137);
nor U13669 (N_13669,N_12096,N_10336);
and U13670 (N_13670,N_11279,N_10672);
xor U13671 (N_13671,N_11345,N_12468);
or U13672 (N_13672,N_11828,N_10188);
nand U13673 (N_13673,N_10979,N_11856);
and U13674 (N_13674,N_11592,N_11052);
nor U13675 (N_13675,N_11508,N_10286);
nor U13676 (N_13676,N_10089,N_11599);
nand U13677 (N_13677,N_12317,N_11002);
nand U13678 (N_13678,N_10195,N_10258);
xnor U13679 (N_13679,N_11401,N_11365);
nand U13680 (N_13680,N_10012,N_10932);
xnor U13681 (N_13681,N_10178,N_11287);
nand U13682 (N_13682,N_10287,N_10161);
or U13683 (N_13683,N_10863,N_11606);
nor U13684 (N_13684,N_12181,N_11432);
nand U13685 (N_13685,N_11804,N_11757);
nor U13686 (N_13686,N_11622,N_12433);
or U13687 (N_13687,N_11145,N_10591);
nand U13688 (N_13688,N_11755,N_12353);
or U13689 (N_13689,N_10030,N_12373);
or U13690 (N_13690,N_10943,N_10512);
nand U13691 (N_13691,N_11333,N_11615);
nand U13692 (N_13692,N_12031,N_10561);
xnor U13693 (N_13693,N_11517,N_11292);
nand U13694 (N_13694,N_10630,N_10391);
nor U13695 (N_13695,N_11198,N_12189);
xnor U13696 (N_13696,N_10127,N_10300);
xnor U13697 (N_13697,N_10432,N_10695);
nor U13698 (N_13698,N_11689,N_12299);
nand U13699 (N_13699,N_11500,N_11502);
xnor U13700 (N_13700,N_11044,N_11654);
and U13701 (N_13701,N_11611,N_12280);
nand U13702 (N_13702,N_12162,N_11231);
and U13703 (N_13703,N_11244,N_12008);
nand U13704 (N_13704,N_10242,N_10113);
or U13705 (N_13705,N_12271,N_10972);
or U13706 (N_13706,N_11332,N_11171);
or U13707 (N_13707,N_10974,N_11195);
nand U13708 (N_13708,N_11285,N_11966);
and U13709 (N_13709,N_10547,N_11912);
xnor U13710 (N_13710,N_11096,N_11265);
xor U13711 (N_13711,N_10434,N_10275);
and U13712 (N_13712,N_12293,N_12418);
or U13713 (N_13713,N_11476,N_11264);
nand U13714 (N_13714,N_12253,N_12394);
or U13715 (N_13715,N_11777,N_11794);
nor U13716 (N_13716,N_10137,N_12030);
nor U13717 (N_13717,N_12474,N_10386);
nor U13718 (N_13718,N_11386,N_11278);
xor U13719 (N_13719,N_11056,N_11413);
nand U13720 (N_13720,N_10249,N_10355);
xnor U13721 (N_13721,N_11201,N_10357);
nor U13722 (N_13722,N_10756,N_11297);
or U13723 (N_13723,N_12477,N_11744);
or U13724 (N_13724,N_11497,N_12345);
and U13725 (N_13725,N_10771,N_11159);
xnor U13726 (N_13726,N_10531,N_10266);
xnor U13727 (N_13727,N_12102,N_11799);
nand U13728 (N_13728,N_12228,N_10002);
nor U13729 (N_13729,N_10279,N_11080);
and U13730 (N_13730,N_12200,N_11565);
nand U13731 (N_13731,N_11491,N_11269);
nand U13732 (N_13732,N_11031,N_10912);
or U13733 (N_13733,N_12075,N_10500);
nor U13734 (N_13734,N_11684,N_11902);
nand U13735 (N_13735,N_11506,N_11407);
or U13736 (N_13736,N_10084,N_11561);
and U13737 (N_13737,N_10268,N_12025);
nand U13738 (N_13738,N_10009,N_10866);
xnor U13739 (N_13739,N_11950,N_10473);
nor U13740 (N_13740,N_10865,N_10647);
or U13741 (N_13741,N_10116,N_11182);
nor U13742 (N_13742,N_11034,N_11211);
xor U13743 (N_13743,N_10403,N_11399);
xor U13744 (N_13744,N_12347,N_10481);
and U13745 (N_13745,N_10563,N_12002);
nor U13746 (N_13746,N_11220,N_11196);
and U13747 (N_13747,N_10491,N_11621);
nor U13748 (N_13748,N_11649,N_10140);
nor U13749 (N_13749,N_10746,N_11315);
xnor U13750 (N_13750,N_11044,N_11319);
and U13751 (N_13751,N_12140,N_11230);
or U13752 (N_13752,N_11739,N_12174);
nand U13753 (N_13753,N_11962,N_10562);
nand U13754 (N_13754,N_11822,N_12073);
nor U13755 (N_13755,N_10295,N_10415);
and U13756 (N_13756,N_11744,N_11492);
or U13757 (N_13757,N_11845,N_11855);
nand U13758 (N_13758,N_12161,N_11800);
nor U13759 (N_13759,N_10494,N_11822);
nand U13760 (N_13760,N_11346,N_11182);
nand U13761 (N_13761,N_11220,N_11708);
and U13762 (N_13762,N_10427,N_10914);
nor U13763 (N_13763,N_11977,N_11474);
or U13764 (N_13764,N_10400,N_12269);
nor U13765 (N_13765,N_10892,N_11586);
and U13766 (N_13766,N_11217,N_11797);
nand U13767 (N_13767,N_12167,N_12401);
or U13768 (N_13768,N_11329,N_12092);
xor U13769 (N_13769,N_11875,N_12019);
xor U13770 (N_13770,N_12358,N_11561);
nor U13771 (N_13771,N_10180,N_10573);
xor U13772 (N_13772,N_10450,N_10363);
xor U13773 (N_13773,N_10459,N_12260);
or U13774 (N_13774,N_12143,N_11107);
and U13775 (N_13775,N_10545,N_11231);
nand U13776 (N_13776,N_12273,N_10799);
nor U13777 (N_13777,N_12417,N_12486);
xor U13778 (N_13778,N_11277,N_10596);
or U13779 (N_13779,N_11457,N_11315);
and U13780 (N_13780,N_11345,N_10080);
xnor U13781 (N_13781,N_10298,N_11352);
nand U13782 (N_13782,N_12124,N_11392);
nand U13783 (N_13783,N_11331,N_12095);
nand U13784 (N_13784,N_12232,N_10732);
and U13785 (N_13785,N_11735,N_12205);
nand U13786 (N_13786,N_10410,N_10391);
nand U13787 (N_13787,N_11357,N_10560);
xor U13788 (N_13788,N_11857,N_12107);
nand U13789 (N_13789,N_12346,N_10013);
nor U13790 (N_13790,N_12182,N_11009);
nor U13791 (N_13791,N_10078,N_12124);
or U13792 (N_13792,N_11362,N_12050);
and U13793 (N_13793,N_12396,N_12482);
and U13794 (N_13794,N_11488,N_11626);
or U13795 (N_13795,N_11351,N_10237);
nor U13796 (N_13796,N_10648,N_10969);
nand U13797 (N_13797,N_11842,N_11398);
and U13798 (N_13798,N_11260,N_10428);
nor U13799 (N_13799,N_10483,N_11244);
and U13800 (N_13800,N_11902,N_11341);
and U13801 (N_13801,N_10613,N_12469);
xnor U13802 (N_13802,N_12330,N_11693);
xnor U13803 (N_13803,N_11952,N_11402);
nand U13804 (N_13804,N_10932,N_10602);
or U13805 (N_13805,N_11555,N_10539);
nand U13806 (N_13806,N_11456,N_10117);
or U13807 (N_13807,N_10077,N_11934);
and U13808 (N_13808,N_11782,N_11036);
nor U13809 (N_13809,N_11075,N_11458);
or U13810 (N_13810,N_11819,N_10992);
nor U13811 (N_13811,N_11943,N_12309);
or U13812 (N_13812,N_12267,N_11713);
and U13813 (N_13813,N_11843,N_10422);
and U13814 (N_13814,N_11805,N_10855);
and U13815 (N_13815,N_11954,N_11874);
nand U13816 (N_13816,N_10675,N_11725);
or U13817 (N_13817,N_12158,N_11564);
and U13818 (N_13818,N_11842,N_11244);
nor U13819 (N_13819,N_11766,N_10298);
nor U13820 (N_13820,N_12111,N_10066);
and U13821 (N_13821,N_10051,N_11813);
or U13822 (N_13822,N_10170,N_11515);
or U13823 (N_13823,N_12141,N_10319);
and U13824 (N_13824,N_11369,N_12044);
xor U13825 (N_13825,N_11524,N_10952);
xnor U13826 (N_13826,N_12333,N_10901);
nand U13827 (N_13827,N_12460,N_11255);
nor U13828 (N_13828,N_11521,N_11105);
nand U13829 (N_13829,N_12400,N_12174);
nand U13830 (N_13830,N_11859,N_10368);
nand U13831 (N_13831,N_10146,N_12491);
xor U13832 (N_13832,N_10952,N_11433);
or U13833 (N_13833,N_12264,N_10373);
nor U13834 (N_13834,N_10960,N_11051);
xor U13835 (N_13835,N_11430,N_10149);
or U13836 (N_13836,N_11995,N_11336);
and U13837 (N_13837,N_12012,N_11294);
and U13838 (N_13838,N_10759,N_11848);
xor U13839 (N_13839,N_11048,N_12331);
or U13840 (N_13840,N_10681,N_10302);
and U13841 (N_13841,N_11050,N_10434);
and U13842 (N_13842,N_10316,N_11638);
or U13843 (N_13843,N_12378,N_10059);
or U13844 (N_13844,N_11893,N_10819);
nor U13845 (N_13845,N_10666,N_10151);
xnor U13846 (N_13846,N_12195,N_11607);
or U13847 (N_13847,N_10602,N_10887);
xnor U13848 (N_13848,N_11310,N_12221);
or U13849 (N_13849,N_11740,N_12438);
nor U13850 (N_13850,N_12377,N_11982);
and U13851 (N_13851,N_12060,N_10370);
nor U13852 (N_13852,N_10206,N_10616);
nand U13853 (N_13853,N_11754,N_11735);
or U13854 (N_13854,N_11618,N_11734);
nand U13855 (N_13855,N_11471,N_12118);
and U13856 (N_13856,N_12398,N_11847);
nand U13857 (N_13857,N_10651,N_11544);
or U13858 (N_13858,N_11713,N_10424);
xor U13859 (N_13859,N_11346,N_10435);
xnor U13860 (N_13860,N_12343,N_11780);
nand U13861 (N_13861,N_10079,N_12272);
and U13862 (N_13862,N_10239,N_10953);
xor U13863 (N_13863,N_11706,N_11536);
xor U13864 (N_13864,N_12016,N_11061);
and U13865 (N_13865,N_10232,N_11296);
nor U13866 (N_13866,N_10179,N_10454);
xor U13867 (N_13867,N_10924,N_10643);
or U13868 (N_13868,N_10733,N_11743);
nor U13869 (N_13869,N_10384,N_10853);
xor U13870 (N_13870,N_10765,N_10947);
nor U13871 (N_13871,N_10615,N_11338);
and U13872 (N_13872,N_10214,N_11523);
or U13873 (N_13873,N_10526,N_10633);
nand U13874 (N_13874,N_10904,N_11832);
xor U13875 (N_13875,N_10743,N_11033);
or U13876 (N_13876,N_10770,N_11431);
or U13877 (N_13877,N_10714,N_10335);
or U13878 (N_13878,N_12052,N_10080);
nor U13879 (N_13879,N_12262,N_10270);
xnor U13880 (N_13880,N_10149,N_12432);
or U13881 (N_13881,N_11468,N_12365);
and U13882 (N_13882,N_11620,N_10268);
nand U13883 (N_13883,N_12404,N_12486);
or U13884 (N_13884,N_11089,N_12133);
and U13885 (N_13885,N_10542,N_11142);
xnor U13886 (N_13886,N_11346,N_11834);
nand U13887 (N_13887,N_11988,N_12420);
or U13888 (N_13888,N_10972,N_11187);
or U13889 (N_13889,N_11159,N_10934);
xor U13890 (N_13890,N_10215,N_10084);
xnor U13891 (N_13891,N_10206,N_10502);
and U13892 (N_13892,N_10637,N_11830);
nor U13893 (N_13893,N_10875,N_12021);
nor U13894 (N_13894,N_11295,N_12072);
nor U13895 (N_13895,N_11812,N_10577);
nand U13896 (N_13896,N_12059,N_10784);
xor U13897 (N_13897,N_11471,N_11678);
nand U13898 (N_13898,N_12432,N_10172);
nor U13899 (N_13899,N_10443,N_10718);
and U13900 (N_13900,N_12041,N_10374);
xor U13901 (N_13901,N_10768,N_10217);
or U13902 (N_13902,N_10152,N_11232);
xnor U13903 (N_13903,N_10242,N_10108);
or U13904 (N_13904,N_11936,N_10390);
xnor U13905 (N_13905,N_10867,N_11637);
and U13906 (N_13906,N_10704,N_11620);
xnor U13907 (N_13907,N_11512,N_11886);
xnor U13908 (N_13908,N_10798,N_12031);
nand U13909 (N_13909,N_12152,N_10198);
nor U13910 (N_13910,N_10508,N_12282);
xnor U13911 (N_13911,N_11965,N_10986);
and U13912 (N_13912,N_12316,N_12238);
nand U13913 (N_13913,N_12073,N_11806);
xor U13914 (N_13914,N_10080,N_11132);
and U13915 (N_13915,N_11591,N_11943);
nor U13916 (N_13916,N_10536,N_11708);
xnor U13917 (N_13917,N_10523,N_11551);
and U13918 (N_13918,N_10177,N_11239);
nor U13919 (N_13919,N_10304,N_10114);
nand U13920 (N_13920,N_11515,N_12268);
nor U13921 (N_13921,N_11625,N_11475);
or U13922 (N_13922,N_12432,N_12060);
nand U13923 (N_13923,N_12050,N_10859);
and U13924 (N_13924,N_11146,N_11902);
and U13925 (N_13925,N_10293,N_12173);
and U13926 (N_13926,N_10240,N_10472);
xor U13927 (N_13927,N_11726,N_11679);
or U13928 (N_13928,N_10141,N_11756);
xor U13929 (N_13929,N_12282,N_10040);
or U13930 (N_13930,N_10152,N_11670);
and U13931 (N_13931,N_12211,N_12193);
xnor U13932 (N_13932,N_11277,N_11906);
nor U13933 (N_13933,N_11451,N_11020);
and U13934 (N_13934,N_11669,N_10212);
nand U13935 (N_13935,N_12254,N_10126);
and U13936 (N_13936,N_11832,N_11654);
or U13937 (N_13937,N_11985,N_10342);
or U13938 (N_13938,N_12052,N_10403);
or U13939 (N_13939,N_10914,N_10907);
or U13940 (N_13940,N_12261,N_12018);
nand U13941 (N_13941,N_11245,N_11867);
xnor U13942 (N_13942,N_10582,N_10172);
xor U13943 (N_13943,N_10826,N_11815);
nor U13944 (N_13944,N_10473,N_11482);
xor U13945 (N_13945,N_11206,N_12093);
xnor U13946 (N_13946,N_11259,N_10107);
xnor U13947 (N_13947,N_12295,N_10285);
xor U13948 (N_13948,N_11984,N_10705);
xnor U13949 (N_13949,N_10072,N_10731);
nand U13950 (N_13950,N_10721,N_10020);
or U13951 (N_13951,N_10103,N_12049);
nor U13952 (N_13952,N_10564,N_11512);
and U13953 (N_13953,N_10027,N_10103);
and U13954 (N_13954,N_12137,N_11843);
or U13955 (N_13955,N_10874,N_10151);
nand U13956 (N_13956,N_10757,N_11043);
nor U13957 (N_13957,N_10358,N_10286);
nor U13958 (N_13958,N_11718,N_12365);
xnor U13959 (N_13959,N_10085,N_11030);
and U13960 (N_13960,N_10533,N_10134);
or U13961 (N_13961,N_10198,N_12487);
and U13962 (N_13962,N_10761,N_10050);
nor U13963 (N_13963,N_12294,N_10880);
xor U13964 (N_13964,N_10104,N_12345);
nand U13965 (N_13965,N_10520,N_12270);
and U13966 (N_13966,N_10189,N_12312);
or U13967 (N_13967,N_11937,N_12172);
nor U13968 (N_13968,N_11139,N_10727);
nor U13969 (N_13969,N_12440,N_11647);
nor U13970 (N_13970,N_10493,N_11722);
and U13971 (N_13971,N_11693,N_10477);
nor U13972 (N_13972,N_10143,N_11913);
or U13973 (N_13973,N_10710,N_11952);
and U13974 (N_13974,N_11694,N_11454);
or U13975 (N_13975,N_12023,N_11610);
or U13976 (N_13976,N_11266,N_10470);
xor U13977 (N_13977,N_11600,N_11228);
and U13978 (N_13978,N_11114,N_10552);
or U13979 (N_13979,N_10041,N_11912);
or U13980 (N_13980,N_11842,N_10042);
or U13981 (N_13981,N_10380,N_11317);
nand U13982 (N_13982,N_12490,N_10395);
nand U13983 (N_13983,N_11268,N_11004);
nand U13984 (N_13984,N_11800,N_11793);
nand U13985 (N_13985,N_10674,N_11486);
nand U13986 (N_13986,N_12466,N_10481);
or U13987 (N_13987,N_10601,N_10645);
nor U13988 (N_13988,N_10263,N_11694);
and U13989 (N_13989,N_10582,N_10094);
nand U13990 (N_13990,N_11977,N_11743);
or U13991 (N_13991,N_11800,N_11446);
nand U13992 (N_13992,N_11487,N_11305);
and U13993 (N_13993,N_10630,N_11792);
or U13994 (N_13994,N_11938,N_11001);
nand U13995 (N_13995,N_11892,N_10266);
nand U13996 (N_13996,N_12057,N_10622);
and U13997 (N_13997,N_11098,N_12107);
or U13998 (N_13998,N_10028,N_12396);
nand U13999 (N_13999,N_11073,N_11013);
and U14000 (N_14000,N_10289,N_11360);
xor U14001 (N_14001,N_12289,N_12288);
and U14002 (N_14002,N_12253,N_10419);
nor U14003 (N_14003,N_12385,N_10467);
nand U14004 (N_14004,N_10195,N_10644);
and U14005 (N_14005,N_11939,N_11033);
xor U14006 (N_14006,N_11653,N_12256);
nand U14007 (N_14007,N_11826,N_11508);
nand U14008 (N_14008,N_11204,N_11280);
xor U14009 (N_14009,N_10483,N_11271);
nand U14010 (N_14010,N_10506,N_10923);
nand U14011 (N_14011,N_10488,N_11446);
and U14012 (N_14012,N_10238,N_12309);
nor U14013 (N_14013,N_10420,N_10077);
nor U14014 (N_14014,N_10263,N_10196);
nand U14015 (N_14015,N_10427,N_12230);
or U14016 (N_14016,N_11575,N_12322);
nor U14017 (N_14017,N_12226,N_10588);
or U14018 (N_14018,N_11278,N_11907);
and U14019 (N_14019,N_10082,N_11956);
or U14020 (N_14020,N_12308,N_10085);
and U14021 (N_14021,N_11829,N_12394);
nor U14022 (N_14022,N_10509,N_11469);
and U14023 (N_14023,N_11520,N_10068);
xor U14024 (N_14024,N_10617,N_10118);
or U14025 (N_14025,N_10018,N_11062);
and U14026 (N_14026,N_12162,N_12468);
and U14027 (N_14027,N_11913,N_11169);
nand U14028 (N_14028,N_11323,N_10561);
and U14029 (N_14029,N_10544,N_11183);
nor U14030 (N_14030,N_11549,N_10997);
or U14031 (N_14031,N_12135,N_11549);
nand U14032 (N_14032,N_10923,N_10742);
and U14033 (N_14033,N_10045,N_10913);
xnor U14034 (N_14034,N_10887,N_10169);
and U14035 (N_14035,N_10321,N_10292);
nor U14036 (N_14036,N_11562,N_11427);
or U14037 (N_14037,N_10232,N_11685);
xnor U14038 (N_14038,N_10528,N_10408);
nand U14039 (N_14039,N_10508,N_10405);
xnor U14040 (N_14040,N_10885,N_10664);
nand U14041 (N_14041,N_11836,N_10322);
nand U14042 (N_14042,N_12112,N_11589);
xor U14043 (N_14043,N_10318,N_11668);
and U14044 (N_14044,N_10979,N_11518);
xor U14045 (N_14045,N_11796,N_11149);
xor U14046 (N_14046,N_11429,N_11443);
xnor U14047 (N_14047,N_12214,N_12179);
or U14048 (N_14048,N_11298,N_11884);
and U14049 (N_14049,N_12075,N_12371);
and U14050 (N_14050,N_11409,N_11508);
and U14051 (N_14051,N_10804,N_10870);
nor U14052 (N_14052,N_12071,N_12077);
nand U14053 (N_14053,N_11688,N_12388);
or U14054 (N_14054,N_11067,N_11795);
and U14055 (N_14055,N_11859,N_11201);
xnor U14056 (N_14056,N_10365,N_11967);
and U14057 (N_14057,N_11844,N_11269);
or U14058 (N_14058,N_10877,N_10596);
nor U14059 (N_14059,N_10537,N_12406);
or U14060 (N_14060,N_11213,N_10529);
or U14061 (N_14061,N_11453,N_11297);
xor U14062 (N_14062,N_11953,N_12403);
or U14063 (N_14063,N_10110,N_12321);
nor U14064 (N_14064,N_10753,N_10206);
xnor U14065 (N_14065,N_11679,N_11721);
and U14066 (N_14066,N_12283,N_10606);
xor U14067 (N_14067,N_10958,N_10262);
nor U14068 (N_14068,N_11745,N_11761);
xor U14069 (N_14069,N_10895,N_10691);
nor U14070 (N_14070,N_12436,N_10599);
xnor U14071 (N_14071,N_11865,N_10992);
and U14072 (N_14072,N_10575,N_11911);
nand U14073 (N_14073,N_11443,N_10475);
nand U14074 (N_14074,N_10233,N_12244);
and U14075 (N_14075,N_10949,N_11194);
nor U14076 (N_14076,N_12150,N_12296);
xor U14077 (N_14077,N_11030,N_10734);
nor U14078 (N_14078,N_11561,N_11554);
nand U14079 (N_14079,N_10876,N_10277);
and U14080 (N_14080,N_11110,N_11663);
nand U14081 (N_14081,N_10328,N_12460);
xor U14082 (N_14082,N_10510,N_10802);
and U14083 (N_14083,N_10566,N_11558);
nand U14084 (N_14084,N_12026,N_11039);
and U14085 (N_14085,N_11652,N_12475);
or U14086 (N_14086,N_11326,N_11568);
nand U14087 (N_14087,N_11848,N_11854);
or U14088 (N_14088,N_11028,N_11909);
xor U14089 (N_14089,N_10418,N_11862);
xor U14090 (N_14090,N_12114,N_10280);
nand U14091 (N_14091,N_11606,N_11882);
nand U14092 (N_14092,N_10138,N_11119);
nor U14093 (N_14093,N_10175,N_10140);
or U14094 (N_14094,N_11882,N_10428);
nor U14095 (N_14095,N_10494,N_11160);
nor U14096 (N_14096,N_10641,N_10235);
xnor U14097 (N_14097,N_11639,N_10235);
nand U14098 (N_14098,N_10883,N_11607);
nand U14099 (N_14099,N_12008,N_11777);
and U14100 (N_14100,N_11609,N_11053);
or U14101 (N_14101,N_12000,N_11892);
and U14102 (N_14102,N_10480,N_12221);
nand U14103 (N_14103,N_11290,N_12466);
nand U14104 (N_14104,N_12381,N_11962);
xor U14105 (N_14105,N_10848,N_10499);
xor U14106 (N_14106,N_11425,N_12176);
xnor U14107 (N_14107,N_10770,N_11403);
xor U14108 (N_14108,N_10112,N_12398);
xnor U14109 (N_14109,N_10555,N_10942);
or U14110 (N_14110,N_10291,N_12058);
or U14111 (N_14111,N_10366,N_11186);
xnor U14112 (N_14112,N_10487,N_11827);
xnor U14113 (N_14113,N_11495,N_11938);
or U14114 (N_14114,N_12249,N_10381);
or U14115 (N_14115,N_10486,N_10160);
nand U14116 (N_14116,N_10817,N_10506);
nand U14117 (N_14117,N_10828,N_12043);
or U14118 (N_14118,N_10936,N_11191);
and U14119 (N_14119,N_10760,N_11068);
nand U14120 (N_14120,N_11252,N_10683);
nor U14121 (N_14121,N_12363,N_10724);
xor U14122 (N_14122,N_11266,N_11668);
nor U14123 (N_14123,N_11984,N_10459);
xnor U14124 (N_14124,N_11621,N_10591);
nor U14125 (N_14125,N_10888,N_12162);
nor U14126 (N_14126,N_12287,N_12318);
nor U14127 (N_14127,N_11580,N_12355);
nand U14128 (N_14128,N_10405,N_11094);
xor U14129 (N_14129,N_12208,N_10739);
or U14130 (N_14130,N_11266,N_11763);
xor U14131 (N_14131,N_11614,N_10549);
and U14132 (N_14132,N_10369,N_10234);
nand U14133 (N_14133,N_10507,N_10968);
nand U14134 (N_14134,N_11743,N_11621);
and U14135 (N_14135,N_10546,N_10427);
nor U14136 (N_14136,N_11778,N_11113);
or U14137 (N_14137,N_11719,N_10336);
or U14138 (N_14138,N_10394,N_10437);
nor U14139 (N_14139,N_12163,N_10039);
and U14140 (N_14140,N_10105,N_10325);
or U14141 (N_14141,N_11908,N_12359);
nand U14142 (N_14142,N_11159,N_11559);
or U14143 (N_14143,N_12046,N_11027);
or U14144 (N_14144,N_11559,N_12408);
nor U14145 (N_14145,N_11929,N_11742);
or U14146 (N_14146,N_11053,N_11063);
nand U14147 (N_14147,N_10665,N_11554);
xor U14148 (N_14148,N_11026,N_10448);
xor U14149 (N_14149,N_12414,N_11719);
or U14150 (N_14150,N_11026,N_11222);
or U14151 (N_14151,N_10965,N_10062);
or U14152 (N_14152,N_12258,N_11862);
or U14153 (N_14153,N_10269,N_10887);
xnor U14154 (N_14154,N_12290,N_10280);
or U14155 (N_14155,N_11365,N_10954);
or U14156 (N_14156,N_10097,N_11903);
or U14157 (N_14157,N_12126,N_12217);
nor U14158 (N_14158,N_11319,N_10217);
nor U14159 (N_14159,N_11012,N_11419);
and U14160 (N_14160,N_11659,N_11252);
xnor U14161 (N_14161,N_11952,N_11922);
or U14162 (N_14162,N_11663,N_10895);
and U14163 (N_14163,N_10520,N_11073);
nor U14164 (N_14164,N_11376,N_11420);
xnor U14165 (N_14165,N_11418,N_11650);
nor U14166 (N_14166,N_11338,N_10105);
and U14167 (N_14167,N_11275,N_10843);
xor U14168 (N_14168,N_11712,N_11135);
and U14169 (N_14169,N_12071,N_11948);
and U14170 (N_14170,N_10051,N_12454);
and U14171 (N_14171,N_12000,N_10318);
and U14172 (N_14172,N_12011,N_11914);
nand U14173 (N_14173,N_10303,N_11565);
and U14174 (N_14174,N_12335,N_10110);
or U14175 (N_14175,N_11005,N_10297);
xor U14176 (N_14176,N_10076,N_10255);
or U14177 (N_14177,N_10041,N_12359);
xor U14178 (N_14178,N_10817,N_11198);
nand U14179 (N_14179,N_11799,N_11981);
nor U14180 (N_14180,N_10163,N_11247);
nand U14181 (N_14181,N_10429,N_10896);
and U14182 (N_14182,N_10330,N_10135);
xnor U14183 (N_14183,N_12273,N_11511);
xor U14184 (N_14184,N_10716,N_10937);
or U14185 (N_14185,N_10468,N_12490);
xor U14186 (N_14186,N_11842,N_11572);
or U14187 (N_14187,N_12116,N_10645);
nand U14188 (N_14188,N_10467,N_10446);
or U14189 (N_14189,N_10269,N_12494);
and U14190 (N_14190,N_10548,N_11831);
nand U14191 (N_14191,N_12347,N_11196);
nor U14192 (N_14192,N_10298,N_10677);
or U14193 (N_14193,N_12301,N_12033);
or U14194 (N_14194,N_10745,N_10733);
xnor U14195 (N_14195,N_10197,N_10490);
and U14196 (N_14196,N_11240,N_11781);
or U14197 (N_14197,N_11917,N_11166);
nand U14198 (N_14198,N_11799,N_10345);
nand U14199 (N_14199,N_10407,N_12408);
nor U14200 (N_14200,N_11388,N_11023);
nor U14201 (N_14201,N_10843,N_10103);
and U14202 (N_14202,N_12154,N_12221);
or U14203 (N_14203,N_10090,N_11484);
nor U14204 (N_14204,N_11965,N_11745);
and U14205 (N_14205,N_11753,N_11022);
nand U14206 (N_14206,N_11769,N_12484);
xnor U14207 (N_14207,N_12114,N_12275);
and U14208 (N_14208,N_11936,N_10273);
nand U14209 (N_14209,N_11240,N_10772);
nor U14210 (N_14210,N_10424,N_12221);
or U14211 (N_14211,N_10699,N_10926);
xor U14212 (N_14212,N_10873,N_11554);
or U14213 (N_14213,N_12240,N_11102);
xnor U14214 (N_14214,N_12128,N_11930);
nor U14215 (N_14215,N_10428,N_11540);
xnor U14216 (N_14216,N_10159,N_10288);
nand U14217 (N_14217,N_11299,N_12091);
xnor U14218 (N_14218,N_11954,N_11794);
and U14219 (N_14219,N_10548,N_12049);
nor U14220 (N_14220,N_11479,N_11141);
or U14221 (N_14221,N_11302,N_10016);
and U14222 (N_14222,N_10732,N_11970);
nor U14223 (N_14223,N_11660,N_12040);
or U14224 (N_14224,N_11833,N_11857);
and U14225 (N_14225,N_10329,N_11724);
nor U14226 (N_14226,N_12060,N_11438);
and U14227 (N_14227,N_12424,N_11575);
nor U14228 (N_14228,N_11241,N_10908);
nand U14229 (N_14229,N_12493,N_11746);
nor U14230 (N_14230,N_10813,N_10817);
xor U14231 (N_14231,N_11301,N_10161);
nand U14232 (N_14232,N_12379,N_11438);
nand U14233 (N_14233,N_12315,N_11746);
nor U14234 (N_14234,N_11826,N_10299);
or U14235 (N_14235,N_11177,N_12357);
nand U14236 (N_14236,N_12243,N_10936);
nand U14237 (N_14237,N_10819,N_10323);
nand U14238 (N_14238,N_12388,N_10617);
nor U14239 (N_14239,N_11250,N_11222);
or U14240 (N_14240,N_12333,N_12097);
nor U14241 (N_14241,N_12168,N_11974);
nand U14242 (N_14242,N_11798,N_12183);
nand U14243 (N_14243,N_10023,N_12158);
xor U14244 (N_14244,N_11495,N_10298);
and U14245 (N_14245,N_11197,N_10319);
and U14246 (N_14246,N_11004,N_10225);
or U14247 (N_14247,N_11498,N_11035);
nor U14248 (N_14248,N_12138,N_12063);
or U14249 (N_14249,N_12008,N_10180);
xor U14250 (N_14250,N_10357,N_12359);
or U14251 (N_14251,N_10448,N_11987);
and U14252 (N_14252,N_10769,N_11298);
and U14253 (N_14253,N_11108,N_11995);
and U14254 (N_14254,N_11283,N_10542);
xnor U14255 (N_14255,N_10479,N_10959);
or U14256 (N_14256,N_10291,N_10321);
nand U14257 (N_14257,N_11773,N_10000);
xor U14258 (N_14258,N_11700,N_10597);
nor U14259 (N_14259,N_11974,N_11679);
nand U14260 (N_14260,N_10630,N_10552);
xnor U14261 (N_14261,N_11212,N_10121);
or U14262 (N_14262,N_11559,N_12142);
and U14263 (N_14263,N_11285,N_10840);
or U14264 (N_14264,N_12137,N_12209);
nor U14265 (N_14265,N_12001,N_11680);
nor U14266 (N_14266,N_12029,N_12217);
nand U14267 (N_14267,N_10806,N_11339);
nand U14268 (N_14268,N_10382,N_10967);
nand U14269 (N_14269,N_10610,N_11171);
and U14270 (N_14270,N_11707,N_10058);
nor U14271 (N_14271,N_10455,N_10482);
or U14272 (N_14272,N_11385,N_10074);
and U14273 (N_14273,N_11831,N_12203);
and U14274 (N_14274,N_12474,N_11329);
xnor U14275 (N_14275,N_10414,N_11712);
nand U14276 (N_14276,N_10861,N_11139);
nand U14277 (N_14277,N_12458,N_12369);
and U14278 (N_14278,N_11856,N_10712);
and U14279 (N_14279,N_10587,N_11858);
nor U14280 (N_14280,N_12348,N_10929);
and U14281 (N_14281,N_10000,N_10050);
or U14282 (N_14282,N_11631,N_12138);
nand U14283 (N_14283,N_11303,N_11173);
and U14284 (N_14284,N_10402,N_10109);
or U14285 (N_14285,N_10333,N_11900);
xor U14286 (N_14286,N_11525,N_11295);
xor U14287 (N_14287,N_10178,N_10578);
or U14288 (N_14288,N_12211,N_12050);
nand U14289 (N_14289,N_11948,N_11611);
or U14290 (N_14290,N_10560,N_11260);
and U14291 (N_14291,N_10985,N_12269);
nand U14292 (N_14292,N_10030,N_10958);
or U14293 (N_14293,N_11419,N_11945);
nand U14294 (N_14294,N_11130,N_11609);
xnor U14295 (N_14295,N_12404,N_10445);
xnor U14296 (N_14296,N_11818,N_11895);
and U14297 (N_14297,N_11019,N_11692);
nor U14298 (N_14298,N_11213,N_12414);
xnor U14299 (N_14299,N_11327,N_10428);
or U14300 (N_14300,N_10002,N_11277);
or U14301 (N_14301,N_10565,N_12073);
or U14302 (N_14302,N_11105,N_10032);
xnor U14303 (N_14303,N_12402,N_12241);
or U14304 (N_14304,N_11970,N_12490);
xnor U14305 (N_14305,N_10955,N_12023);
nand U14306 (N_14306,N_11767,N_11215);
nand U14307 (N_14307,N_10478,N_12146);
xnor U14308 (N_14308,N_10386,N_10219);
or U14309 (N_14309,N_10615,N_11950);
nor U14310 (N_14310,N_11780,N_11863);
or U14311 (N_14311,N_12073,N_11051);
nor U14312 (N_14312,N_10784,N_11358);
and U14313 (N_14313,N_11709,N_10641);
or U14314 (N_14314,N_11478,N_11796);
or U14315 (N_14315,N_11054,N_11019);
xor U14316 (N_14316,N_12267,N_11557);
and U14317 (N_14317,N_11443,N_10785);
nor U14318 (N_14318,N_11754,N_10949);
nor U14319 (N_14319,N_10635,N_12112);
nor U14320 (N_14320,N_12111,N_11914);
xnor U14321 (N_14321,N_12388,N_11006);
xor U14322 (N_14322,N_11160,N_10478);
or U14323 (N_14323,N_10108,N_10223);
or U14324 (N_14324,N_11400,N_11803);
or U14325 (N_14325,N_12206,N_11357);
and U14326 (N_14326,N_11779,N_10359);
or U14327 (N_14327,N_11211,N_10981);
nor U14328 (N_14328,N_10282,N_11664);
nor U14329 (N_14329,N_11348,N_10849);
or U14330 (N_14330,N_11182,N_10019);
nor U14331 (N_14331,N_11292,N_10133);
xor U14332 (N_14332,N_11176,N_10521);
xnor U14333 (N_14333,N_11663,N_12314);
or U14334 (N_14334,N_10754,N_11433);
and U14335 (N_14335,N_10917,N_10315);
or U14336 (N_14336,N_12416,N_11264);
nor U14337 (N_14337,N_11395,N_10317);
xor U14338 (N_14338,N_11801,N_11679);
nor U14339 (N_14339,N_10016,N_10420);
nand U14340 (N_14340,N_10607,N_11957);
nor U14341 (N_14341,N_10002,N_10745);
and U14342 (N_14342,N_10444,N_11530);
or U14343 (N_14343,N_11697,N_11271);
nand U14344 (N_14344,N_11643,N_11825);
nand U14345 (N_14345,N_11596,N_10122);
and U14346 (N_14346,N_11848,N_12352);
and U14347 (N_14347,N_10541,N_10604);
and U14348 (N_14348,N_10844,N_10429);
and U14349 (N_14349,N_10748,N_10088);
xnor U14350 (N_14350,N_10694,N_11927);
or U14351 (N_14351,N_12386,N_11580);
nand U14352 (N_14352,N_11006,N_10874);
xnor U14353 (N_14353,N_12457,N_11732);
and U14354 (N_14354,N_12004,N_11081);
or U14355 (N_14355,N_12148,N_11550);
xor U14356 (N_14356,N_10191,N_12306);
nand U14357 (N_14357,N_10107,N_10905);
xnor U14358 (N_14358,N_11719,N_10203);
nand U14359 (N_14359,N_10087,N_10753);
xnor U14360 (N_14360,N_10884,N_10805);
xor U14361 (N_14361,N_12427,N_10720);
nor U14362 (N_14362,N_10011,N_11726);
and U14363 (N_14363,N_12038,N_10668);
or U14364 (N_14364,N_10901,N_12196);
and U14365 (N_14365,N_10739,N_12001);
nor U14366 (N_14366,N_10810,N_10214);
xor U14367 (N_14367,N_10443,N_10485);
nand U14368 (N_14368,N_10008,N_11117);
nand U14369 (N_14369,N_10229,N_11093);
or U14370 (N_14370,N_10768,N_11800);
or U14371 (N_14371,N_10429,N_10423);
xor U14372 (N_14372,N_11907,N_11571);
nand U14373 (N_14373,N_12062,N_10519);
nor U14374 (N_14374,N_10650,N_10716);
and U14375 (N_14375,N_11207,N_11539);
nand U14376 (N_14376,N_11253,N_12282);
and U14377 (N_14377,N_11778,N_10219);
nand U14378 (N_14378,N_10745,N_12125);
or U14379 (N_14379,N_12142,N_12300);
or U14380 (N_14380,N_12107,N_12344);
or U14381 (N_14381,N_10081,N_11735);
xor U14382 (N_14382,N_10011,N_10986);
and U14383 (N_14383,N_12081,N_12239);
nand U14384 (N_14384,N_12340,N_11699);
nor U14385 (N_14385,N_12493,N_11470);
and U14386 (N_14386,N_11646,N_10147);
and U14387 (N_14387,N_11755,N_10014);
xor U14388 (N_14388,N_12092,N_12390);
nand U14389 (N_14389,N_10612,N_10507);
or U14390 (N_14390,N_10854,N_12455);
xnor U14391 (N_14391,N_11891,N_11953);
and U14392 (N_14392,N_10687,N_10825);
or U14393 (N_14393,N_11660,N_10997);
or U14394 (N_14394,N_11383,N_10355);
or U14395 (N_14395,N_12061,N_12294);
nor U14396 (N_14396,N_10264,N_10213);
or U14397 (N_14397,N_11904,N_11886);
nand U14398 (N_14398,N_12266,N_11101);
or U14399 (N_14399,N_11320,N_11957);
and U14400 (N_14400,N_10485,N_11374);
and U14401 (N_14401,N_10549,N_10935);
nand U14402 (N_14402,N_12356,N_11308);
xor U14403 (N_14403,N_10853,N_12425);
nand U14404 (N_14404,N_10991,N_10052);
and U14405 (N_14405,N_11766,N_11149);
xor U14406 (N_14406,N_12000,N_10599);
and U14407 (N_14407,N_10988,N_10552);
and U14408 (N_14408,N_10384,N_12430);
or U14409 (N_14409,N_12205,N_12375);
xor U14410 (N_14410,N_11741,N_12491);
nand U14411 (N_14411,N_10161,N_12075);
nand U14412 (N_14412,N_11646,N_12398);
nor U14413 (N_14413,N_11739,N_11907);
nand U14414 (N_14414,N_10440,N_10528);
or U14415 (N_14415,N_10588,N_11993);
xnor U14416 (N_14416,N_11332,N_10621);
nand U14417 (N_14417,N_11284,N_11447);
nand U14418 (N_14418,N_11578,N_11461);
nand U14419 (N_14419,N_10861,N_12193);
xnor U14420 (N_14420,N_12429,N_11690);
and U14421 (N_14421,N_10415,N_12471);
xnor U14422 (N_14422,N_12243,N_12097);
xnor U14423 (N_14423,N_10768,N_10181);
nor U14424 (N_14424,N_11169,N_11376);
nor U14425 (N_14425,N_10984,N_12351);
nor U14426 (N_14426,N_11719,N_12477);
nor U14427 (N_14427,N_11507,N_11258);
nand U14428 (N_14428,N_11525,N_10660);
or U14429 (N_14429,N_11515,N_10450);
nor U14430 (N_14430,N_10923,N_11548);
xor U14431 (N_14431,N_12181,N_12314);
nor U14432 (N_14432,N_10513,N_11756);
xnor U14433 (N_14433,N_10097,N_12423);
or U14434 (N_14434,N_11934,N_10685);
or U14435 (N_14435,N_12002,N_10374);
nor U14436 (N_14436,N_12059,N_10728);
or U14437 (N_14437,N_10553,N_10868);
or U14438 (N_14438,N_11341,N_11805);
xor U14439 (N_14439,N_10217,N_11324);
xor U14440 (N_14440,N_11104,N_11005);
xor U14441 (N_14441,N_10185,N_12461);
nor U14442 (N_14442,N_10306,N_11569);
and U14443 (N_14443,N_12167,N_11271);
or U14444 (N_14444,N_10675,N_12093);
nor U14445 (N_14445,N_10806,N_11631);
nor U14446 (N_14446,N_10964,N_10697);
and U14447 (N_14447,N_12438,N_11746);
and U14448 (N_14448,N_10490,N_11780);
and U14449 (N_14449,N_11411,N_11345);
xor U14450 (N_14450,N_11700,N_10508);
or U14451 (N_14451,N_12275,N_10238);
nor U14452 (N_14452,N_10825,N_12224);
or U14453 (N_14453,N_12367,N_10928);
nand U14454 (N_14454,N_11355,N_10092);
and U14455 (N_14455,N_11867,N_11015);
and U14456 (N_14456,N_10238,N_10786);
nand U14457 (N_14457,N_10576,N_11642);
nor U14458 (N_14458,N_10854,N_11467);
xor U14459 (N_14459,N_10015,N_11032);
and U14460 (N_14460,N_10996,N_10934);
xnor U14461 (N_14461,N_10929,N_12241);
or U14462 (N_14462,N_11120,N_11610);
or U14463 (N_14463,N_11058,N_11100);
and U14464 (N_14464,N_10473,N_10893);
and U14465 (N_14465,N_10272,N_10247);
or U14466 (N_14466,N_10139,N_11897);
xor U14467 (N_14467,N_11991,N_11046);
nand U14468 (N_14468,N_12268,N_10150);
xor U14469 (N_14469,N_10967,N_10903);
and U14470 (N_14470,N_10876,N_12155);
xnor U14471 (N_14471,N_11775,N_10632);
nand U14472 (N_14472,N_10413,N_10020);
nand U14473 (N_14473,N_10120,N_10721);
or U14474 (N_14474,N_11328,N_12040);
xnor U14475 (N_14475,N_10347,N_10757);
or U14476 (N_14476,N_12294,N_10300);
and U14477 (N_14477,N_11029,N_12003);
xor U14478 (N_14478,N_10179,N_11380);
and U14479 (N_14479,N_10297,N_11878);
or U14480 (N_14480,N_10537,N_11224);
nor U14481 (N_14481,N_10297,N_12463);
or U14482 (N_14482,N_11346,N_11923);
nor U14483 (N_14483,N_11165,N_10656);
and U14484 (N_14484,N_11083,N_10443);
nand U14485 (N_14485,N_10305,N_10847);
xnor U14486 (N_14486,N_12286,N_11482);
or U14487 (N_14487,N_11268,N_10454);
and U14488 (N_14488,N_10031,N_11118);
and U14489 (N_14489,N_11232,N_10897);
or U14490 (N_14490,N_11632,N_11668);
and U14491 (N_14491,N_11986,N_11091);
nor U14492 (N_14492,N_11384,N_10377);
xor U14493 (N_14493,N_12065,N_11055);
nand U14494 (N_14494,N_11972,N_11482);
nand U14495 (N_14495,N_12021,N_11744);
nor U14496 (N_14496,N_11403,N_11846);
xor U14497 (N_14497,N_11619,N_10358);
xnor U14498 (N_14498,N_11788,N_10800);
nor U14499 (N_14499,N_11311,N_12383);
xor U14500 (N_14500,N_10541,N_10603);
or U14501 (N_14501,N_10678,N_11015);
xnor U14502 (N_14502,N_10446,N_11705);
nand U14503 (N_14503,N_11421,N_10558);
nand U14504 (N_14504,N_11879,N_10653);
and U14505 (N_14505,N_11461,N_12392);
or U14506 (N_14506,N_11222,N_10276);
or U14507 (N_14507,N_11070,N_10130);
xnor U14508 (N_14508,N_10482,N_10550);
or U14509 (N_14509,N_10904,N_12132);
nand U14510 (N_14510,N_10664,N_11447);
xor U14511 (N_14511,N_11644,N_10882);
nand U14512 (N_14512,N_11335,N_10034);
nor U14513 (N_14513,N_10991,N_10585);
nor U14514 (N_14514,N_10425,N_11660);
xor U14515 (N_14515,N_11834,N_11948);
or U14516 (N_14516,N_11725,N_11792);
nand U14517 (N_14517,N_10622,N_11913);
nor U14518 (N_14518,N_10386,N_12253);
nor U14519 (N_14519,N_11198,N_11306);
and U14520 (N_14520,N_10807,N_11075);
nand U14521 (N_14521,N_12498,N_10417);
xor U14522 (N_14522,N_10259,N_11887);
and U14523 (N_14523,N_11720,N_10799);
nor U14524 (N_14524,N_12338,N_11820);
and U14525 (N_14525,N_11915,N_10779);
nand U14526 (N_14526,N_11417,N_10207);
nand U14527 (N_14527,N_11347,N_10131);
xnor U14528 (N_14528,N_10955,N_11815);
xnor U14529 (N_14529,N_10050,N_11117);
and U14530 (N_14530,N_11748,N_10647);
xor U14531 (N_14531,N_11449,N_10527);
or U14532 (N_14532,N_10443,N_12051);
nand U14533 (N_14533,N_11081,N_10350);
nand U14534 (N_14534,N_11266,N_11801);
or U14535 (N_14535,N_10542,N_11720);
or U14536 (N_14536,N_11456,N_12287);
nor U14537 (N_14537,N_11660,N_11841);
xnor U14538 (N_14538,N_10535,N_10840);
and U14539 (N_14539,N_10219,N_11818);
or U14540 (N_14540,N_11972,N_11802);
xor U14541 (N_14541,N_12043,N_10055);
or U14542 (N_14542,N_12335,N_12147);
and U14543 (N_14543,N_10805,N_12158);
nand U14544 (N_14544,N_11810,N_10511);
nor U14545 (N_14545,N_10800,N_12482);
nand U14546 (N_14546,N_10245,N_12206);
xor U14547 (N_14547,N_12079,N_10315);
and U14548 (N_14548,N_10501,N_11534);
xnor U14549 (N_14549,N_11056,N_11548);
and U14550 (N_14550,N_11153,N_12195);
nand U14551 (N_14551,N_10757,N_10750);
xnor U14552 (N_14552,N_11021,N_11270);
and U14553 (N_14553,N_10330,N_10508);
and U14554 (N_14554,N_10484,N_11509);
and U14555 (N_14555,N_11822,N_11012);
xnor U14556 (N_14556,N_10585,N_10780);
or U14557 (N_14557,N_11887,N_12476);
and U14558 (N_14558,N_10492,N_10580);
or U14559 (N_14559,N_10901,N_11713);
nand U14560 (N_14560,N_11081,N_10539);
and U14561 (N_14561,N_12473,N_10229);
nor U14562 (N_14562,N_11466,N_10056);
xor U14563 (N_14563,N_10298,N_11696);
nor U14564 (N_14564,N_10727,N_12298);
xnor U14565 (N_14565,N_11486,N_12293);
nor U14566 (N_14566,N_10765,N_11667);
nor U14567 (N_14567,N_11826,N_11619);
nor U14568 (N_14568,N_10831,N_12036);
nor U14569 (N_14569,N_11391,N_11606);
or U14570 (N_14570,N_11199,N_10810);
nand U14571 (N_14571,N_11648,N_10385);
xnor U14572 (N_14572,N_10229,N_10835);
or U14573 (N_14573,N_11640,N_10260);
xor U14574 (N_14574,N_11216,N_10137);
xnor U14575 (N_14575,N_10225,N_11229);
nand U14576 (N_14576,N_10886,N_10226);
xor U14577 (N_14577,N_11133,N_12435);
and U14578 (N_14578,N_11246,N_11647);
nor U14579 (N_14579,N_10889,N_11165);
nand U14580 (N_14580,N_11659,N_10960);
xor U14581 (N_14581,N_10988,N_10951);
and U14582 (N_14582,N_10508,N_12257);
nor U14583 (N_14583,N_11883,N_10191);
or U14584 (N_14584,N_11424,N_10965);
or U14585 (N_14585,N_12028,N_10202);
or U14586 (N_14586,N_11618,N_10315);
xor U14587 (N_14587,N_10168,N_11701);
xnor U14588 (N_14588,N_11512,N_11980);
nor U14589 (N_14589,N_11505,N_10790);
nor U14590 (N_14590,N_12380,N_11830);
nand U14591 (N_14591,N_12311,N_10402);
nor U14592 (N_14592,N_10965,N_11947);
or U14593 (N_14593,N_12134,N_10852);
nand U14594 (N_14594,N_11679,N_10531);
nor U14595 (N_14595,N_11083,N_10368);
xnor U14596 (N_14596,N_12127,N_10104);
nand U14597 (N_14597,N_10737,N_11755);
nand U14598 (N_14598,N_11191,N_12480);
or U14599 (N_14599,N_10454,N_11523);
or U14600 (N_14600,N_10371,N_11726);
or U14601 (N_14601,N_11105,N_11370);
xnor U14602 (N_14602,N_12077,N_10961);
and U14603 (N_14603,N_12258,N_11604);
nor U14604 (N_14604,N_11764,N_10888);
or U14605 (N_14605,N_11520,N_12262);
nor U14606 (N_14606,N_11811,N_10726);
nand U14607 (N_14607,N_10735,N_11481);
or U14608 (N_14608,N_10080,N_10239);
nor U14609 (N_14609,N_11835,N_11124);
nor U14610 (N_14610,N_11979,N_11895);
nor U14611 (N_14611,N_10127,N_12121);
nand U14612 (N_14612,N_12446,N_12357);
xnor U14613 (N_14613,N_10401,N_10613);
nand U14614 (N_14614,N_11553,N_11158);
or U14615 (N_14615,N_11343,N_11241);
xnor U14616 (N_14616,N_11490,N_10012);
or U14617 (N_14617,N_11209,N_10569);
xor U14618 (N_14618,N_11280,N_12269);
nand U14619 (N_14619,N_11495,N_10138);
or U14620 (N_14620,N_10558,N_11535);
nand U14621 (N_14621,N_10840,N_11327);
nand U14622 (N_14622,N_10915,N_11060);
nor U14623 (N_14623,N_12403,N_12491);
nand U14624 (N_14624,N_10747,N_10925);
or U14625 (N_14625,N_11926,N_12156);
nand U14626 (N_14626,N_12293,N_10902);
nor U14627 (N_14627,N_10525,N_10834);
and U14628 (N_14628,N_11082,N_10196);
or U14629 (N_14629,N_11578,N_10277);
nand U14630 (N_14630,N_10031,N_11382);
nor U14631 (N_14631,N_11170,N_11469);
xor U14632 (N_14632,N_11534,N_12301);
nor U14633 (N_14633,N_10902,N_10883);
nor U14634 (N_14634,N_11544,N_11386);
nand U14635 (N_14635,N_10575,N_10604);
xnor U14636 (N_14636,N_12434,N_11265);
or U14637 (N_14637,N_11027,N_11946);
or U14638 (N_14638,N_10221,N_11219);
nor U14639 (N_14639,N_11570,N_12475);
nor U14640 (N_14640,N_11470,N_12461);
nand U14641 (N_14641,N_11882,N_11016);
and U14642 (N_14642,N_10338,N_12487);
and U14643 (N_14643,N_11225,N_12417);
nor U14644 (N_14644,N_11426,N_11717);
nor U14645 (N_14645,N_12081,N_10089);
xnor U14646 (N_14646,N_10269,N_12165);
xnor U14647 (N_14647,N_12466,N_11968);
nor U14648 (N_14648,N_11462,N_11053);
xnor U14649 (N_14649,N_10624,N_12363);
or U14650 (N_14650,N_12093,N_11767);
or U14651 (N_14651,N_10514,N_10251);
nand U14652 (N_14652,N_11147,N_11382);
xor U14653 (N_14653,N_10156,N_10040);
and U14654 (N_14654,N_10785,N_10114);
nand U14655 (N_14655,N_11393,N_10691);
or U14656 (N_14656,N_10701,N_11691);
nand U14657 (N_14657,N_12028,N_10554);
and U14658 (N_14658,N_10272,N_11720);
and U14659 (N_14659,N_12158,N_10417);
or U14660 (N_14660,N_12029,N_10552);
xnor U14661 (N_14661,N_11772,N_11312);
nand U14662 (N_14662,N_11727,N_10871);
or U14663 (N_14663,N_10111,N_11189);
nor U14664 (N_14664,N_11175,N_11732);
or U14665 (N_14665,N_11620,N_10782);
and U14666 (N_14666,N_11077,N_10251);
nor U14667 (N_14667,N_10378,N_10616);
nand U14668 (N_14668,N_11784,N_12234);
and U14669 (N_14669,N_11622,N_12374);
or U14670 (N_14670,N_10048,N_10043);
nand U14671 (N_14671,N_11963,N_12418);
nand U14672 (N_14672,N_10370,N_10907);
nor U14673 (N_14673,N_10441,N_12084);
or U14674 (N_14674,N_12330,N_12192);
nor U14675 (N_14675,N_10371,N_11851);
and U14676 (N_14676,N_10808,N_10729);
and U14677 (N_14677,N_10081,N_10543);
nand U14678 (N_14678,N_10554,N_10250);
and U14679 (N_14679,N_11850,N_11434);
xnor U14680 (N_14680,N_10227,N_11715);
xnor U14681 (N_14681,N_11206,N_10752);
and U14682 (N_14682,N_11657,N_11232);
or U14683 (N_14683,N_10571,N_10082);
and U14684 (N_14684,N_10918,N_11655);
nor U14685 (N_14685,N_12057,N_10443);
and U14686 (N_14686,N_10413,N_11851);
xnor U14687 (N_14687,N_12476,N_11704);
xor U14688 (N_14688,N_11643,N_12276);
nand U14689 (N_14689,N_12483,N_10903);
xor U14690 (N_14690,N_10226,N_10647);
nand U14691 (N_14691,N_11205,N_12068);
or U14692 (N_14692,N_10367,N_10116);
xor U14693 (N_14693,N_11619,N_10999);
nand U14694 (N_14694,N_10986,N_10348);
xor U14695 (N_14695,N_11833,N_12016);
xor U14696 (N_14696,N_10979,N_12167);
xnor U14697 (N_14697,N_10065,N_11294);
xnor U14698 (N_14698,N_12234,N_10789);
nor U14699 (N_14699,N_10771,N_12102);
and U14700 (N_14700,N_11510,N_12480);
or U14701 (N_14701,N_10835,N_11761);
nor U14702 (N_14702,N_10992,N_11357);
nor U14703 (N_14703,N_10823,N_10099);
nor U14704 (N_14704,N_12090,N_10517);
and U14705 (N_14705,N_10922,N_10190);
nand U14706 (N_14706,N_10753,N_11138);
and U14707 (N_14707,N_10510,N_11134);
nand U14708 (N_14708,N_11302,N_11247);
and U14709 (N_14709,N_11883,N_10834);
xor U14710 (N_14710,N_10857,N_10476);
or U14711 (N_14711,N_11166,N_10438);
or U14712 (N_14712,N_11079,N_11717);
nand U14713 (N_14713,N_12479,N_11501);
and U14714 (N_14714,N_10134,N_11597);
xor U14715 (N_14715,N_11666,N_10187);
nor U14716 (N_14716,N_12462,N_10300);
nor U14717 (N_14717,N_10466,N_11290);
nand U14718 (N_14718,N_10415,N_11036);
nand U14719 (N_14719,N_11992,N_11690);
and U14720 (N_14720,N_11679,N_10034);
nand U14721 (N_14721,N_11785,N_11434);
xnor U14722 (N_14722,N_12154,N_11777);
nand U14723 (N_14723,N_10829,N_10495);
and U14724 (N_14724,N_12490,N_11053);
nand U14725 (N_14725,N_11366,N_10878);
nand U14726 (N_14726,N_11681,N_10183);
xor U14727 (N_14727,N_12401,N_11875);
nor U14728 (N_14728,N_11863,N_11356);
nor U14729 (N_14729,N_11370,N_10231);
xnor U14730 (N_14730,N_12380,N_10112);
or U14731 (N_14731,N_12197,N_10569);
xor U14732 (N_14732,N_10670,N_10765);
nand U14733 (N_14733,N_12496,N_10113);
nand U14734 (N_14734,N_11547,N_11535);
or U14735 (N_14735,N_11913,N_10060);
nor U14736 (N_14736,N_12126,N_11466);
nand U14737 (N_14737,N_10396,N_11367);
nor U14738 (N_14738,N_11781,N_12439);
xor U14739 (N_14739,N_11545,N_12078);
and U14740 (N_14740,N_10026,N_12269);
xor U14741 (N_14741,N_10805,N_10914);
xnor U14742 (N_14742,N_10568,N_11267);
or U14743 (N_14743,N_11125,N_11393);
or U14744 (N_14744,N_11972,N_10912);
xnor U14745 (N_14745,N_11087,N_11315);
or U14746 (N_14746,N_10104,N_11918);
or U14747 (N_14747,N_10288,N_12361);
or U14748 (N_14748,N_11863,N_11878);
xnor U14749 (N_14749,N_10512,N_12279);
or U14750 (N_14750,N_10147,N_10014);
nor U14751 (N_14751,N_11835,N_12414);
xnor U14752 (N_14752,N_11095,N_11854);
xor U14753 (N_14753,N_12228,N_11976);
nand U14754 (N_14754,N_12274,N_10075);
or U14755 (N_14755,N_11885,N_11911);
and U14756 (N_14756,N_11789,N_12248);
or U14757 (N_14757,N_12204,N_10437);
and U14758 (N_14758,N_11487,N_11397);
nor U14759 (N_14759,N_10598,N_11854);
or U14760 (N_14760,N_11112,N_11279);
nand U14761 (N_14761,N_10459,N_10364);
and U14762 (N_14762,N_11358,N_12283);
or U14763 (N_14763,N_10853,N_10192);
and U14764 (N_14764,N_11706,N_10991);
or U14765 (N_14765,N_11663,N_12417);
nor U14766 (N_14766,N_10806,N_11350);
xnor U14767 (N_14767,N_11736,N_10916);
nand U14768 (N_14768,N_11418,N_11682);
or U14769 (N_14769,N_12467,N_10851);
and U14770 (N_14770,N_12258,N_11977);
nand U14771 (N_14771,N_11136,N_10227);
nor U14772 (N_14772,N_10463,N_12227);
xor U14773 (N_14773,N_10379,N_10630);
xnor U14774 (N_14774,N_12392,N_12375);
and U14775 (N_14775,N_10500,N_11374);
or U14776 (N_14776,N_11885,N_10722);
nand U14777 (N_14777,N_11840,N_10172);
and U14778 (N_14778,N_12364,N_11812);
nor U14779 (N_14779,N_11721,N_11638);
nor U14780 (N_14780,N_12450,N_12105);
and U14781 (N_14781,N_11759,N_11559);
xnor U14782 (N_14782,N_10243,N_10273);
nand U14783 (N_14783,N_12313,N_11879);
and U14784 (N_14784,N_10802,N_10895);
nor U14785 (N_14785,N_10956,N_10006);
xor U14786 (N_14786,N_11674,N_12064);
nand U14787 (N_14787,N_11068,N_10398);
xnor U14788 (N_14788,N_10867,N_11651);
or U14789 (N_14789,N_11767,N_11219);
or U14790 (N_14790,N_11579,N_12144);
and U14791 (N_14791,N_11196,N_11150);
xor U14792 (N_14792,N_12194,N_12064);
nand U14793 (N_14793,N_11524,N_12069);
nor U14794 (N_14794,N_10335,N_12404);
or U14795 (N_14795,N_12250,N_10310);
nand U14796 (N_14796,N_11380,N_12439);
xnor U14797 (N_14797,N_10726,N_11368);
xnor U14798 (N_14798,N_10592,N_11174);
or U14799 (N_14799,N_11741,N_10459);
and U14800 (N_14800,N_10473,N_10389);
and U14801 (N_14801,N_10177,N_10904);
nor U14802 (N_14802,N_11651,N_11481);
nand U14803 (N_14803,N_12436,N_10362);
or U14804 (N_14804,N_10366,N_10268);
nor U14805 (N_14805,N_10343,N_10959);
nand U14806 (N_14806,N_10276,N_11592);
and U14807 (N_14807,N_12005,N_11094);
nand U14808 (N_14808,N_11792,N_10908);
nor U14809 (N_14809,N_11418,N_11869);
nand U14810 (N_14810,N_11086,N_10478);
and U14811 (N_14811,N_12165,N_10592);
nand U14812 (N_14812,N_10328,N_11510);
nand U14813 (N_14813,N_11905,N_12387);
nor U14814 (N_14814,N_10101,N_10894);
nor U14815 (N_14815,N_10713,N_11050);
or U14816 (N_14816,N_10038,N_10125);
and U14817 (N_14817,N_11587,N_11274);
nor U14818 (N_14818,N_11441,N_12349);
nor U14819 (N_14819,N_11878,N_12330);
nand U14820 (N_14820,N_11279,N_12328);
and U14821 (N_14821,N_11728,N_12077);
xnor U14822 (N_14822,N_11717,N_10635);
or U14823 (N_14823,N_10818,N_10075);
xnor U14824 (N_14824,N_11033,N_10496);
xnor U14825 (N_14825,N_10404,N_11570);
and U14826 (N_14826,N_10430,N_11785);
or U14827 (N_14827,N_11886,N_10774);
or U14828 (N_14828,N_11577,N_11770);
and U14829 (N_14829,N_10889,N_10446);
or U14830 (N_14830,N_11221,N_11632);
xnor U14831 (N_14831,N_12021,N_11399);
or U14832 (N_14832,N_11946,N_10040);
xnor U14833 (N_14833,N_11114,N_10481);
xor U14834 (N_14834,N_11482,N_10065);
or U14835 (N_14835,N_10317,N_11976);
and U14836 (N_14836,N_10886,N_10843);
or U14837 (N_14837,N_11719,N_12306);
nand U14838 (N_14838,N_11792,N_12123);
xnor U14839 (N_14839,N_10397,N_11775);
and U14840 (N_14840,N_12436,N_10354);
nand U14841 (N_14841,N_11978,N_10399);
or U14842 (N_14842,N_11198,N_11897);
xnor U14843 (N_14843,N_10754,N_11653);
or U14844 (N_14844,N_10279,N_10753);
xor U14845 (N_14845,N_11316,N_10966);
and U14846 (N_14846,N_12099,N_11357);
xor U14847 (N_14847,N_11631,N_10862);
or U14848 (N_14848,N_11651,N_11498);
nor U14849 (N_14849,N_11080,N_12077);
or U14850 (N_14850,N_10838,N_11606);
nor U14851 (N_14851,N_10385,N_10979);
and U14852 (N_14852,N_11683,N_10391);
nand U14853 (N_14853,N_11575,N_12494);
nor U14854 (N_14854,N_11311,N_10538);
and U14855 (N_14855,N_11733,N_10465);
nand U14856 (N_14856,N_11364,N_12138);
nor U14857 (N_14857,N_10544,N_12326);
nor U14858 (N_14858,N_11744,N_12383);
or U14859 (N_14859,N_11719,N_11299);
nor U14860 (N_14860,N_11973,N_10680);
nand U14861 (N_14861,N_10144,N_10058);
or U14862 (N_14862,N_10893,N_12219);
or U14863 (N_14863,N_10848,N_10552);
or U14864 (N_14864,N_11444,N_10941);
xnor U14865 (N_14865,N_10509,N_11647);
xnor U14866 (N_14866,N_11392,N_10171);
nand U14867 (N_14867,N_11427,N_11515);
nand U14868 (N_14868,N_10376,N_11977);
nand U14869 (N_14869,N_11203,N_11467);
and U14870 (N_14870,N_11691,N_11393);
xor U14871 (N_14871,N_10411,N_12308);
xnor U14872 (N_14872,N_10366,N_11859);
nand U14873 (N_14873,N_11388,N_12139);
and U14874 (N_14874,N_11194,N_11170);
or U14875 (N_14875,N_12492,N_12468);
or U14876 (N_14876,N_11703,N_10467);
nor U14877 (N_14877,N_10275,N_12484);
nor U14878 (N_14878,N_10651,N_10731);
nand U14879 (N_14879,N_12369,N_11894);
or U14880 (N_14880,N_12046,N_11702);
or U14881 (N_14881,N_12390,N_11986);
nor U14882 (N_14882,N_10199,N_12017);
nand U14883 (N_14883,N_11759,N_11722);
nand U14884 (N_14884,N_10351,N_10213);
and U14885 (N_14885,N_12063,N_10921);
nand U14886 (N_14886,N_11353,N_11772);
nor U14887 (N_14887,N_12197,N_11429);
or U14888 (N_14888,N_10977,N_11300);
xor U14889 (N_14889,N_10453,N_11491);
or U14890 (N_14890,N_10936,N_10201);
or U14891 (N_14891,N_10493,N_12452);
nor U14892 (N_14892,N_11368,N_12194);
xor U14893 (N_14893,N_11113,N_12099);
and U14894 (N_14894,N_10732,N_10479);
or U14895 (N_14895,N_11615,N_12274);
and U14896 (N_14896,N_10520,N_10183);
nor U14897 (N_14897,N_12223,N_10160);
or U14898 (N_14898,N_11288,N_10655);
or U14899 (N_14899,N_11129,N_11043);
xnor U14900 (N_14900,N_11040,N_12488);
xor U14901 (N_14901,N_10941,N_10270);
xnor U14902 (N_14902,N_10012,N_10007);
or U14903 (N_14903,N_10987,N_10816);
nand U14904 (N_14904,N_12398,N_10074);
or U14905 (N_14905,N_12035,N_11459);
and U14906 (N_14906,N_11655,N_12375);
or U14907 (N_14907,N_11833,N_12419);
xor U14908 (N_14908,N_10555,N_12223);
nand U14909 (N_14909,N_12394,N_11210);
and U14910 (N_14910,N_10992,N_12486);
xor U14911 (N_14911,N_11654,N_12346);
nor U14912 (N_14912,N_10488,N_11963);
nor U14913 (N_14913,N_10958,N_10741);
or U14914 (N_14914,N_10656,N_12080);
xnor U14915 (N_14915,N_12216,N_10401);
nand U14916 (N_14916,N_11469,N_11846);
or U14917 (N_14917,N_10247,N_12112);
xor U14918 (N_14918,N_10957,N_11890);
xnor U14919 (N_14919,N_10556,N_11209);
and U14920 (N_14920,N_10384,N_11042);
or U14921 (N_14921,N_10085,N_11124);
nand U14922 (N_14922,N_10387,N_11054);
xnor U14923 (N_14923,N_10465,N_10446);
nor U14924 (N_14924,N_11311,N_11541);
and U14925 (N_14925,N_10203,N_11201);
or U14926 (N_14926,N_11481,N_10708);
nand U14927 (N_14927,N_11017,N_10473);
and U14928 (N_14928,N_12325,N_10578);
nor U14929 (N_14929,N_11139,N_11217);
and U14930 (N_14930,N_10320,N_10887);
nor U14931 (N_14931,N_11483,N_10796);
xnor U14932 (N_14932,N_10386,N_12201);
nand U14933 (N_14933,N_12172,N_12039);
xnor U14934 (N_14934,N_10107,N_11691);
or U14935 (N_14935,N_11330,N_10816);
nor U14936 (N_14936,N_10022,N_11444);
nand U14937 (N_14937,N_11774,N_10571);
or U14938 (N_14938,N_12410,N_10096);
xnor U14939 (N_14939,N_10769,N_11966);
xor U14940 (N_14940,N_10288,N_11442);
xnor U14941 (N_14941,N_11495,N_11675);
nand U14942 (N_14942,N_12413,N_11414);
and U14943 (N_14943,N_10811,N_10362);
and U14944 (N_14944,N_12400,N_10788);
xor U14945 (N_14945,N_12431,N_11686);
nand U14946 (N_14946,N_10292,N_11885);
nand U14947 (N_14947,N_11696,N_11021);
xor U14948 (N_14948,N_11762,N_10728);
nor U14949 (N_14949,N_11816,N_10362);
nor U14950 (N_14950,N_11708,N_12094);
and U14951 (N_14951,N_12175,N_10593);
xor U14952 (N_14952,N_10214,N_11249);
nor U14953 (N_14953,N_12496,N_11443);
nor U14954 (N_14954,N_12189,N_10383);
nand U14955 (N_14955,N_10680,N_11591);
nand U14956 (N_14956,N_12307,N_11930);
nor U14957 (N_14957,N_11181,N_11013);
or U14958 (N_14958,N_11884,N_12387);
nor U14959 (N_14959,N_11151,N_10274);
and U14960 (N_14960,N_10821,N_11757);
or U14961 (N_14961,N_11507,N_10252);
or U14962 (N_14962,N_12434,N_10617);
or U14963 (N_14963,N_10754,N_10933);
and U14964 (N_14964,N_10802,N_10463);
nor U14965 (N_14965,N_10150,N_10674);
xnor U14966 (N_14966,N_11464,N_12217);
xor U14967 (N_14967,N_11137,N_10178);
nor U14968 (N_14968,N_10265,N_11554);
nand U14969 (N_14969,N_11553,N_10016);
nand U14970 (N_14970,N_11322,N_10239);
nor U14971 (N_14971,N_12330,N_12023);
and U14972 (N_14972,N_11462,N_11018);
nand U14973 (N_14973,N_10958,N_11150);
or U14974 (N_14974,N_10233,N_10672);
nor U14975 (N_14975,N_10433,N_12292);
xor U14976 (N_14976,N_11892,N_10652);
and U14977 (N_14977,N_10291,N_11837);
or U14978 (N_14978,N_10948,N_11115);
nand U14979 (N_14979,N_12048,N_12332);
xor U14980 (N_14980,N_10444,N_11059);
nor U14981 (N_14981,N_11403,N_10983);
xnor U14982 (N_14982,N_11246,N_10311);
nand U14983 (N_14983,N_11190,N_12115);
nor U14984 (N_14984,N_12096,N_10926);
and U14985 (N_14985,N_11294,N_11213);
nor U14986 (N_14986,N_12420,N_11147);
or U14987 (N_14987,N_10596,N_11699);
or U14988 (N_14988,N_12021,N_12453);
nor U14989 (N_14989,N_11849,N_12468);
and U14990 (N_14990,N_12322,N_11796);
nor U14991 (N_14991,N_11616,N_12095);
and U14992 (N_14992,N_11595,N_10362);
nand U14993 (N_14993,N_12095,N_10399);
or U14994 (N_14994,N_10782,N_10767);
and U14995 (N_14995,N_12340,N_11401);
xnor U14996 (N_14996,N_11051,N_11588);
or U14997 (N_14997,N_10038,N_11609);
and U14998 (N_14998,N_10499,N_12139);
and U14999 (N_14999,N_10898,N_11351);
xor U15000 (N_15000,N_14997,N_13875);
nor U15001 (N_15001,N_13786,N_14735);
xnor U15002 (N_15002,N_13282,N_14726);
or U15003 (N_15003,N_13395,N_14132);
nor U15004 (N_15004,N_14544,N_14933);
nand U15005 (N_15005,N_14700,N_14439);
xnor U15006 (N_15006,N_13207,N_14667);
nand U15007 (N_15007,N_12911,N_12530);
nor U15008 (N_15008,N_13757,N_14660);
or U15009 (N_15009,N_14902,N_13359);
and U15010 (N_15010,N_13179,N_14119);
and U15011 (N_15011,N_12847,N_13271);
xnor U15012 (N_15012,N_13176,N_14067);
or U15013 (N_15013,N_14755,N_14225);
nor U15014 (N_15014,N_14800,N_14303);
nor U15015 (N_15015,N_13639,N_12739);
xor U15016 (N_15016,N_13522,N_13364);
nand U15017 (N_15017,N_13361,N_13495);
and U15018 (N_15018,N_14390,N_14602);
or U15019 (N_15019,N_13314,N_13248);
or U15020 (N_15020,N_12827,N_14992);
xnor U15021 (N_15021,N_14190,N_12955);
or U15022 (N_15022,N_14071,N_14236);
and U15023 (N_15023,N_12543,N_13962);
and U15024 (N_15024,N_12695,N_12604);
xor U15025 (N_15025,N_14978,N_14287);
xnor U15026 (N_15026,N_14682,N_13329);
or U15027 (N_15027,N_13113,N_13706);
nor U15028 (N_15028,N_13840,N_12879);
or U15029 (N_15029,N_13820,N_14603);
or U15030 (N_15030,N_13990,N_14825);
and U15031 (N_15031,N_14569,N_14763);
or U15032 (N_15032,N_12786,N_14799);
nor U15033 (N_15033,N_13237,N_13803);
or U15034 (N_15034,N_13251,N_14771);
nand U15035 (N_15035,N_13685,N_13942);
nand U15036 (N_15036,N_13457,N_12779);
and U15037 (N_15037,N_13755,N_14724);
or U15038 (N_15038,N_14080,N_14969);
or U15039 (N_15039,N_13273,N_13376);
and U15040 (N_15040,N_14211,N_12658);
nand U15041 (N_15041,N_14989,N_14470);
nor U15042 (N_15042,N_14112,N_12965);
nand U15043 (N_15043,N_13426,N_14055);
nor U15044 (N_15044,N_12523,N_14916);
nor U15045 (N_15045,N_13069,N_13167);
xnor U15046 (N_15046,N_13869,N_14806);
nor U15047 (N_15047,N_14084,N_14379);
or U15048 (N_15048,N_14123,N_13164);
nand U15049 (N_15049,N_12634,N_13897);
nand U15050 (N_15050,N_14391,N_13455);
xor U15051 (N_15051,N_12657,N_12930);
or U15052 (N_15052,N_13267,N_14954);
nor U15053 (N_15053,N_14296,N_14894);
xnor U15054 (N_15054,N_13527,N_14418);
xnor U15055 (N_15055,N_13230,N_12961);
and U15056 (N_15056,N_14448,N_14374);
xnor U15057 (N_15057,N_14893,N_14666);
and U15058 (N_15058,N_13648,N_14903);
or U15059 (N_15059,N_12748,N_12871);
and U15060 (N_15060,N_13078,N_13265);
nor U15061 (N_15061,N_13913,N_13168);
nor U15062 (N_15062,N_13301,N_13507);
nand U15063 (N_15063,N_14113,N_13851);
nor U15064 (N_15064,N_14051,N_14594);
and U15065 (N_15065,N_13630,N_14298);
nor U15066 (N_15066,N_14986,N_12937);
or U15067 (N_15067,N_13319,N_14573);
and U15068 (N_15068,N_12607,N_13310);
and U15069 (N_15069,N_13831,N_13041);
or U15070 (N_15070,N_13701,N_13155);
and U15071 (N_15071,N_14713,N_12639);
nand U15072 (N_15072,N_13605,N_14496);
and U15073 (N_15073,N_13946,N_13590);
nand U15074 (N_15074,N_13599,N_13083);
nand U15075 (N_15075,N_14446,N_14212);
and U15076 (N_15076,N_14467,N_14261);
nor U15077 (N_15077,N_12694,N_13817);
nor U15078 (N_15078,N_13969,N_12712);
xnor U15079 (N_15079,N_13974,N_12551);
and U15080 (N_15080,N_12941,N_14353);
or U15081 (N_15081,N_13064,N_12790);
xor U15082 (N_15082,N_14527,N_13186);
and U15083 (N_15083,N_12898,N_13438);
nand U15084 (N_15084,N_14128,N_13569);
or U15085 (N_15085,N_14759,N_13858);
nand U15086 (N_15086,N_14737,N_13657);
or U15087 (N_15087,N_13613,N_13995);
and U15088 (N_15088,N_12969,N_14455);
nor U15089 (N_15089,N_14622,N_14795);
nand U15090 (N_15090,N_12725,N_14090);
nand U15091 (N_15091,N_13369,N_13478);
xnor U15092 (N_15092,N_13012,N_13610);
nand U15093 (N_15093,N_13857,N_14677);
or U15094 (N_15094,N_13254,N_12570);
and U15095 (N_15095,N_14299,N_13790);
and U15096 (N_15096,N_12959,N_14230);
xnor U15097 (N_15097,N_13245,N_13025);
or U15098 (N_15098,N_13299,N_12726);
nor U15099 (N_15099,N_12841,N_14535);
nand U15100 (N_15100,N_12706,N_13703);
xor U15101 (N_15101,N_13306,N_12684);
or U15102 (N_15102,N_13655,N_13277);
nor U15103 (N_15103,N_13019,N_14440);
and U15104 (N_15104,N_13042,N_13980);
and U15105 (N_15105,N_14073,N_12799);
xnor U15106 (N_15106,N_14166,N_14510);
nor U15107 (N_15107,N_12599,N_13414);
nand U15108 (N_15108,N_13286,N_13988);
or U15109 (N_15109,N_12980,N_13429);
and U15110 (N_15110,N_14665,N_13567);
or U15111 (N_15111,N_12615,N_12766);
nand U15112 (N_15112,N_14635,N_12801);
and U15113 (N_15113,N_13046,N_14729);
or U15114 (N_15114,N_12782,N_14886);
or U15115 (N_15115,N_12508,N_13094);
or U15116 (N_15116,N_14864,N_13449);
and U15117 (N_15117,N_14576,N_13353);
or U15118 (N_15118,N_14250,N_13462);
nor U15119 (N_15119,N_13589,N_12992);
xor U15120 (N_15120,N_13724,N_14953);
and U15121 (N_15121,N_13062,N_13795);
and U15122 (N_15122,N_13998,N_12518);
nand U15123 (N_15123,N_13366,N_13354);
and U15124 (N_15124,N_13746,N_14523);
or U15125 (N_15125,N_14692,N_13415);
nor U15126 (N_15126,N_13228,N_13517);
and U15127 (N_15127,N_14497,N_13138);
and U15128 (N_15128,N_14215,N_14408);
xor U15129 (N_15129,N_14689,N_12683);
nor U15130 (N_15130,N_12531,N_14063);
and U15131 (N_15131,N_13134,N_14895);
nand U15132 (N_15132,N_13075,N_14740);
xor U15133 (N_15133,N_14445,N_12920);
nor U15134 (N_15134,N_14449,N_13890);
and U15135 (N_15135,N_13016,N_12892);
nor U15136 (N_15136,N_14384,N_13100);
and U15137 (N_15137,N_12951,N_14377);
nor U15138 (N_15138,N_14637,N_14872);
xnor U15139 (N_15139,N_13206,N_14174);
nor U15140 (N_15140,N_14792,N_14963);
xor U15141 (N_15141,N_13994,N_13793);
or U15142 (N_15142,N_13939,N_12534);
or U15143 (N_15143,N_13997,N_13351);
or U15144 (N_15144,N_14307,N_13597);
nor U15145 (N_15145,N_13761,N_14078);
nor U15146 (N_15146,N_14186,N_12734);
or U15147 (N_15147,N_14828,N_14490);
and U15148 (N_15148,N_14779,N_14278);
or U15149 (N_15149,N_14885,N_14350);
nand U15150 (N_15150,N_12882,N_14820);
xor U15151 (N_15151,N_13203,N_12652);
or U15152 (N_15152,N_14362,N_14965);
or U15153 (N_15153,N_13692,N_13472);
xor U15154 (N_15154,N_13022,N_14253);
nor U15155 (N_15155,N_13652,N_13384);
and U15156 (N_15156,N_14505,N_13882);
and U15157 (N_15157,N_12504,N_14781);
and U15158 (N_15158,N_13895,N_14009);
nand U15159 (N_15159,N_14109,N_13911);
xnor U15160 (N_15160,N_14699,N_12632);
or U15161 (N_15161,N_14185,N_13975);
and U15162 (N_15162,N_13082,N_13323);
nand U15163 (N_15163,N_12737,N_14932);
nor U15164 (N_15164,N_14949,N_13493);
nand U15165 (N_15165,N_13289,N_12563);
nor U15166 (N_15166,N_14896,N_13564);
or U15167 (N_15167,N_12957,N_13051);
nand U15168 (N_15168,N_14231,N_14574);
nand U15169 (N_15169,N_12869,N_13506);
nor U15170 (N_15170,N_13201,N_14214);
nor U15171 (N_15171,N_13432,N_13367);
nand U15172 (N_15172,N_12738,N_13782);
nor U15173 (N_15173,N_13643,N_13850);
nand U15174 (N_15174,N_14366,N_14457);
xnor U15175 (N_15175,N_13777,N_13127);
nor U15176 (N_15176,N_13914,N_13656);
nand U15177 (N_15177,N_12721,N_13872);
or U15178 (N_15178,N_13806,N_14783);
nor U15179 (N_15179,N_13119,N_14014);
nand U15180 (N_15180,N_13611,N_13433);
and U15181 (N_15181,N_14942,N_14855);
nor U15182 (N_15182,N_14675,N_14077);
nand U15183 (N_15183,N_13192,N_13787);
and U15184 (N_15184,N_14036,N_13157);
or U15185 (N_15185,N_12881,N_13389);
or U15186 (N_15186,N_13215,N_12773);
xnor U15187 (N_15187,N_14169,N_12752);
nand U15188 (N_15188,N_14027,N_12716);
or U15189 (N_15189,N_13208,N_14846);
and U15190 (N_15190,N_13607,N_12928);
xnor U15191 (N_15191,N_13001,N_14308);
and U15192 (N_15192,N_14427,N_13244);
xor U15193 (N_15193,N_12500,N_14579);
nand U15194 (N_15194,N_13198,N_13349);
nand U15195 (N_15195,N_13832,N_14615);
nor U15196 (N_15196,N_13204,N_13154);
xor U15197 (N_15197,N_13796,N_14605);
and U15198 (N_15198,N_14034,N_13676);
and U15199 (N_15199,N_14008,N_14106);
and U15200 (N_15200,N_13629,N_12846);
nand U15201 (N_15201,N_14450,N_13765);
or U15202 (N_15202,N_13241,N_14901);
nand U15203 (N_15203,N_13823,N_14757);
and U15204 (N_15204,N_14183,N_13712);
nor U15205 (N_15205,N_12741,N_14939);
or U15206 (N_15206,N_13090,N_12884);
nand U15207 (N_15207,N_13234,N_13532);
nor U15208 (N_15208,N_12587,N_14748);
xnor U15209 (N_15209,N_12850,N_14094);
and U15210 (N_15210,N_13054,N_12768);
xnor U15211 (N_15211,N_12876,N_13169);
xor U15212 (N_15212,N_14007,N_14608);
nand U15213 (N_15213,N_14581,N_14679);
nand U15214 (N_15214,N_13702,N_14500);
or U15215 (N_15215,N_13915,N_12536);
nor U15216 (N_15216,N_14884,N_12763);
nor U15217 (N_15217,N_14356,N_13683);
nor U15218 (N_15218,N_14281,N_14426);
or U15219 (N_15219,N_13693,N_13573);
and U15220 (N_15220,N_13191,N_14575);
or U15221 (N_15221,N_12594,N_13818);
or U15222 (N_15222,N_13774,N_13592);
and U15223 (N_15223,N_12525,N_13726);
and U15224 (N_15224,N_13344,N_14772);
nor U15225 (N_15225,N_12544,N_13152);
or U15226 (N_15226,N_13189,N_12901);
xor U15227 (N_15227,N_13822,N_13688);
nand U15228 (N_15228,N_12624,N_14956);
xor U15229 (N_15229,N_14599,N_12538);
and U15230 (N_15230,N_14260,N_14591);
xnor U15231 (N_15231,N_13993,N_12978);
and U15232 (N_15232,N_14566,N_12910);
nor U15233 (N_15233,N_13212,N_14354);
and U15234 (N_15234,N_14201,N_13742);
and U15235 (N_15235,N_14518,N_14826);
or U15236 (N_15236,N_14597,N_14263);
nor U15237 (N_15237,N_12714,N_13149);
nor U15238 (N_15238,N_13531,N_14054);
and U15239 (N_15239,N_13931,N_14829);
and U15240 (N_15240,N_12550,N_13516);
or U15241 (N_15241,N_14035,N_14313);
nand U15242 (N_15242,N_12601,N_13085);
or U15243 (N_15243,N_13442,N_13868);
nand U15244 (N_15244,N_13756,N_14327);
nand U15245 (N_15245,N_14385,N_14802);
or U15246 (N_15246,N_13560,N_12924);
nor U15247 (N_15247,N_14640,N_14911);
nand U15248 (N_15248,N_14013,N_13340);
or U15249 (N_15249,N_13562,N_13233);
and U15250 (N_15250,N_14310,N_14405);
and U15251 (N_15251,N_12511,N_13338);
and U15252 (N_15252,N_12717,N_13794);
and U15253 (N_15253,N_14482,N_14220);
nand U15254 (N_15254,N_14661,N_12557);
nor U15255 (N_15255,N_13576,N_12885);
xor U15256 (N_15256,N_14403,N_14559);
or U15257 (N_15257,N_14223,N_14728);
nor U15258 (N_15258,N_12713,N_12635);
or U15259 (N_15259,N_13469,N_12516);
nor U15260 (N_15260,N_13582,N_14474);
or U15261 (N_15261,N_13031,N_13920);
nor U15262 (N_15262,N_14709,N_13381);
nor U15263 (N_15263,N_14655,N_13659);
nor U15264 (N_15264,N_14380,N_13258);
nor U15265 (N_15265,N_13036,N_14477);
xnor U15266 (N_15266,N_12619,N_13139);
xnor U15267 (N_15267,N_14419,N_14152);
nor U15268 (N_15268,N_12583,N_14842);
nand U15269 (N_15269,N_12993,N_14424);
or U15270 (N_15270,N_13718,N_12997);
and U15271 (N_15271,N_13320,N_13973);
and U15272 (N_15272,N_13866,N_14471);
nand U15273 (N_15273,N_14971,N_13220);
nor U15274 (N_15274,N_14337,N_12715);
or U15275 (N_15275,N_14164,N_14684);
xor U15276 (N_15276,N_12533,N_14756);
xor U15277 (N_15277,N_13135,N_14256);
and U15278 (N_15278,N_14139,N_12872);
nand U15279 (N_15279,N_13346,N_13651);
nor U15280 (N_15280,N_12705,N_14540);
xor U15281 (N_15281,N_13679,N_13935);
xnor U15282 (N_15282,N_13422,N_13977);
or U15283 (N_15283,N_14836,N_13476);
nand U15284 (N_15284,N_12912,N_13654);
nor U15285 (N_15285,N_12784,N_14442);
xnor U15286 (N_15286,N_13072,N_13067);
xnor U15287 (N_15287,N_13484,N_13898);
xor U15288 (N_15288,N_12507,N_14780);
nor U15289 (N_15289,N_12862,N_14782);
nand U15290 (N_15290,N_13081,N_14632);
and U15291 (N_15291,N_13543,N_13918);
or U15292 (N_15292,N_13393,N_13750);
nor U15293 (N_15293,N_14498,N_14791);
nand U15294 (N_15294,N_13190,N_14875);
nor U15295 (N_15295,N_13080,N_12861);
and U15296 (N_15296,N_13884,N_12864);
nand U15297 (N_15297,N_14147,N_13728);
xnor U15298 (N_15298,N_13399,N_14839);
and U15299 (N_15299,N_13956,N_13185);
nor U15300 (N_15300,N_14121,N_13537);
and U15301 (N_15301,N_12711,N_14503);
xnor U15302 (N_15302,N_14217,N_12838);
and U15303 (N_15303,N_13363,N_12877);
nand U15304 (N_15304,N_13644,N_13565);
or U15305 (N_15305,N_14480,N_13128);
or U15306 (N_15306,N_12857,N_12932);
and U15307 (N_15307,N_12939,N_13714);
xor U15308 (N_15308,N_12995,N_14808);
xnor U15309 (N_15309,N_13725,N_14068);
xor U15310 (N_15310,N_12628,N_14393);
nand U15311 (N_15311,N_14987,N_13281);
nand U15312 (N_15312,N_12787,N_14582);
nand U15313 (N_15313,N_13837,N_14821);
nand U15314 (N_15314,N_14289,N_14716);
or U15315 (N_15315,N_13071,N_13934);
nor U15316 (N_15316,N_14598,N_13847);
nor U15317 (N_15317,N_12842,N_12791);
and U15318 (N_15318,N_12769,N_13122);
nand U15319 (N_15319,N_13930,N_13653);
nor U15320 (N_15320,N_14506,N_12584);
or U15321 (N_15321,N_12613,N_13183);
nor U15322 (N_15322,N_14741,N_12775);
xnor U15323 (N_15323,N_12848,N_12627);
nor U15324 (N_15324,N_13156,N_13325);
or U15325 (N_15325,N_14926,N_14601);
and U15326 (N_15326,N_13663,N_14447);
nand U15327 (N_15327,N_13841,N_14562);
xnor U15328 (N_15328,N_13076,N_13261);
nand U15329 (N_15329,N_12761,N_12603);
nand U15330 (N_15330,N_13779,N_13842);
nand U15331 (N_15331,N_14466,N_14056);
nand U15332 (N_15332,N_12960,N_14823);
xnor U15333 (N_15333,N_13058,N_14227);
nor U15334 (N_15334,N_13752,N_13616);
xnor U15335 (N_15335,N_12641,N_14423);
nand U15336 (N_15336,N_13177,N_12863);
xnor U15337 (N_15337,N_13330,N_13408);
or U15338 (N_15338,N_14273,N_14088);
nand U15339 (N_15339,N_14395,N_14941);
xor U15340 (N_15340,N_13465,N_13836);
nand U15341 (N_15341,N_12727,N_14673);
or U15342 (N_15342,N_13955,N_13545);
and U15343 (N_15343,N_13510,N_13419);
xnor U15344 (N_15344,N_14085,N_14845);
or U15345 (N_15345,N_14493,N_14589);
nor U15346 (N_15346,N_13209,N_13691);
nor U15347 (N_15347,N_13747,N_14041);
and U15348 (N_15348,N_12891,N_13754);
nor U15349 (N_15349,N_13073,N_13948);
nand U15350 (N_15350,N_12945,N_12800);
and U15351 (N_15351,N_13514,N_13050);
or U15352 (N_15352,N_14722,N_13958);
nand U15353 (N_15353,N_14696,N_13403);
and U15354 (N_15354,N_14134,N_14137);
xnor U15355 (N_15355,N_13461,N_13608);
xor U15356 (N_15356,N_13987,N_12854);
or U15357 (N_15357,N_13909,N_13061);
nor U15358 (N_15358,N_13385,N_13638);
nand U15359 (N_15359,N_13161,N_14628);
and U15360 (N_15360,N_14315,N_13326);
nor U15361 (N_15361,N_13846,N_12510);
nand U15362 (N_15362,N_14398,N_14465);
nor U15363 (N_15363,N_14421,N_12540);
or U15364 (N_15364,N_14338,N_13680);
nand U15365 (N_15365,N_12580,N_13769);
nand U15366 (N_15366,N_14483,N_13238);
xor U15367 (N_15367,N_13632,N_13398);
and U15368 (N_15368,N_12571,N_12558);
nor U15369 (N_15369,N_14560,N_14999);
and U15370 (N_15370,N_12917,N_13242);
and U15371 (N_15371,N_13813,N_13048);
or U15372 (N_15372,N_14148,N_13658);
nand U15373 (N_15373,N_14010,N_12889);
and U15374 (N_15374,N_13059,N_12923);
and U15375 (N_15375,N_13929,N_14943);
nor U15376 (N_15376,N_14948,N_13887);
xor U15377 (N_15377,N_13079,N_13144);
xor U15378 (N_15378,N_14409,N_12807);
and U15379 (N_15379,N_14822,N_14991);
or U15380 (N_15380,N_14951,N_14351);
xor U15381 (N_15381,N_14837,N_12825);
and U15382 (N_15382,N_14768,N_12865);
or U15383 (N_15383,N_13312,N_14072);
xor U15384 (N_15384,N_12815,N_12699);
nand U15385 (N_15385,N_12593,N_14270);
and U15386 (N_15386,N_14114,N_13454);
nand U15387 (N_15387,N_13473,N_14863);
xnor U15388 (N_15388,N_14208,N_13900);
and U15389 (N_15389,N_14304,N_12781);
nand U15390 (N_15390,N_12692,N_13917);
xor U15391 (N_15391,N_13172,N_14357);
or U15392 (N_15392,N_13810,N_14004);
nand U15393 (N_15393,N_14024,N_14793);
nand U15394 (N_15394,N_14401,N_13165);
and U15395 (N_15395,N_13088,N_14154);
nor U15396 (N_15396,N_14509,N_13766);
and U15397 (N_15397,N_14021,N_13290);
nor U15398 (N_15398,N_13174,N_14751);
or U15399 (N_15399,N_13184,N_12818);
and U15400 (N_15400,N_14146,N_13322);
nor U15401 (N_15401,N_14202,N_14508);
or U15402 (N_15402,N_13269,N_14815);
nor U15403 (N_15403,N_13225,N_12757);
nor U15404 (N_15404,N_14698,N_14070);
nand U15405 (N_15405,N_14542,N_14868);
or U15406 (N_15406,N_14302,N_14025);
xnor U15407 (N_15407,N_14382,N_14974);
nor U15408 (N_15408,N_13358,N_14738);
xnor U15409 (N_15409,N_14539,N_13957);
xnor U15410 (N_15410,N_14428,N_13425);
or U15411 (N_15411,N_12954,N_12823);
and U15412 (N_15412,N_13483,N_12927);
xor U15413 (N_15413,N_12561,N_14180);
nand U15414 (N_15414,N_12883,N_14631);
and U15415 (N_15415,N_14001,N_13740);
xor U15416 (N_15416,N_13421,N_13068);
or U15417 (N_15417,N_14979,N_14288);
xnor U15418 (N_15418,N_14019,N_13137);
xnor U15419 (N_15419,N_14835,N_13451);
or U15420 (N_15420,N_14141,N_13182);
or U15421 (N_15421,N_14099,N_13731);
and U15422 (N_15422,N_13908,N_13949);
nor U15423 (N_15423,N_13318,N_14750);
and U15424 (N_15424,N_14329,N_14163);
or U15425 (N_15425,N_13551,N_14871);
nand U15426 (N_15426,N_14909,N_12909);
and U15427 (N_15427,N_14588,N_13466);
xor U15428 (N_15428,N_12897,N_14411);
nand U15429 (N_15429,N_14649,N_13456);
nor U15430 (N_15430,N_14300,N_13409);
and U15431 (N_15431,N_12868,N_13332);
xor U15432 (N_15432,N_13047,N_14925);
and U15433 (N_15433,N_13760,N_13280);
and U15434 (N_15434,N_13328,N_13240);
and U15435 (N_15435,N_13533,N_12732);
nor U15436 (N_15436,N_13111,N_13053);
and U15437 (N_15437,N_14293,N_14623);
or U15438 (N_15438,N_13523,N_13854);
or U15439 (N_15439,N_12858,N_12546);
and U15440 (N_15440,N_14514,N_13867);
nand U15441 (N_15441,N_12708,N_13453);
nor U15442 (N_15442,N_14468,N_13798);
nor U15443 (N_15443,N_13448,N_12855);
or U15444 (N_15444,N_12703,N_13379);
xor U15445 (N_15445,N_13252,N_13697);
and U15446 (N_15446,N_14914,N_13158);
and U15447 (N_15447,N_12964,N_14235);
xor U15448 (N_15448,N_13427,N_13606);
or U15449 (N_15449,N_14558,N_14504);
nand U15450 (N_15450,N_13859,N_14697);
xor U15451 (N_15451,N_13776,N_14057);
nand U15452 (N_15452,N_14921,N_14340);
and U15453 (N_15453,N_13166,N_12780);
and U15454 (N_15454,N_13479,N_14282);
nor U15455 (N_15455,N_13350,N_14720);
nor U15456 (N_15456,N_13396,N_13243);
and U15457 (N_15457,N_12985,N_13305);
nand U15458 (N_15458,N_14066,N_13650);
or U15459 (N_15459,N_13501,N_12811);
or U15460 (N_15460,N_12777,N_12890);
xnor U15461 (N_15461,N_14228,N_12894);
xnor U15462 (N_15462,N_13197,N_13378);
xor U15463 (N_15463,N_14274,N_12709);
xor U15464 (N_15464,N_14785,N_13260);
nand U15465 (N_15465,N_13450,N_12524);
and U15466 (N_15466,N_14259,N_14478);
and U15467 (N_15467,N_12794,N_14593);
nand U15468 (N_15468,N_12931,N_13646);
xnor U15469 (N_15469,N_14316,N_13043);
or U15470 (N_15470,N_13696,N_12903);
nand U15471 (N_15471,N_13907,N_12754);
and U15472 (N_15472,N_13675,N_13151);
nand U15473 (N_15473,N_14096,N_12968);
nor U15474 (N_15474,N_13812,N_13216);
nor U15475 (N_15475,N_14538,N_14548);
nand U15476 (N_15476,N_14272,N_14120);
and U15477 (N_15477,N_14485,N_14564);
nand U15478 (N_15478,N_13819,N_13721);
xnor U15479 (N_15479,N_13767,N_14511);
and U15480 (N_15480,N_12532,N_13744);
nor U15481 (N_15481,N_12663,N_14714);
and U15482 (N_15482,N_13045,N_12940);
nand U15483 (N_15483,N_13631,N_13097);
nor U15484 (N_15484,N_13581,N_14378);
xor U15485 (N_15485,N_13287,N_12574);
or U15486 (N_15486,N_12866,N_14743);
or U15487 (N_15487,N_12926,N_13263);
or U15488 (N_15488,N_12919,N_14827);
and U15489 (N_15489,N_13536,N_12637);
xor U15490 (N_15490,N_12680,N_12682);
xnor U15491 (N_15491,N_13196,N_14326);
nand U15492 (N_15492,N_12849,N_14335);
nor U15493 (N_15493,N_13377,N_12810);
nor U15494 (N_15494,N_14853,N_14861);
or U15495 (N_15495,N_12674,N_12595);
nand U15496 (N_15496,N_14767,N_14461);
nor U15497 (N_15497,N_14171,N_14079);
nor U15498 (N_15498,N_13849,N_13594);
or U15499 (N_15499,N_14258,N_14422);
nor U15500 (N_15500,N_12772,N_14196);
xnor U15501 (N_15501,N_13499,N_12902);
or U15502 (N_15502,N_12806,N_14881);
nand U15503 (N_15503,N_14050,N_13785);
nand U15504 (N_15504,N_13333,N_14194);
nand U15505 (N_15505,N_12758,N_13110);
or U15506 (N_15506,N_14671,N_14363);
nand U15507 (N_15507,N_13026,N_12696);
or U15508 (N_15508,N_12873,N_14552);
nor U15509 (N_15509,N_14150,N_13732);
xor U15510 (N_15510,N_14416,N_13392);
or U15511 (N_15511,N_12502,N_12614);
nand U15512 (N_15512,N_14923,N_13441);
xor U15513 (N_15513,N_13485,N_13905);
nor U15514 (N_15514,N_12759,N_13259);
xnor U15515 (N_15515,N_14890,N_14040);
xor U15516 (N_15516,N_13649,N_13894);
nand U15517 (N_15517,N_14499,N_13627);
xor U15518 (N_15518,N_13405,N_13246);
xnor U15519 (N_15519,N_14459,N_12552);
and U15520 (N_15520,N_13029,N_14852);
xnor U15521 (N_15521,N_13512,N_12728);
or U15522 (N_15522,N_14131,N_14229);
and U15523 (N_15523,N_14028,N_14117);
xnor U15524 (N_15524,N_13807,N_14805);
or U15525 (N_15525,N_13034,N_14908);
or U15526 (N_15526,N_12554,N_14657);
or U15527 (N_15527,N_14922,N_14676);
xor U15528 (N_15528,N_14929,N_14711);
nor U15529 (N_15529,N_13959,N_12906);
nor U15530 (N_15530,N_14794,N_13788);
nor U15531 (N_15531,N_14678,N_14502);
nor U15532 (N_15532,N_14016,N_13491);
and U15533 (N_15533,N_13255,N_14484);
nand U15534 (N_15534,N_12701,N_14819);
nor U15535 (N_15535,N_14453,N_12675);
nor U15536 (N_15536,N_13596,N_12631);
and U15537 (N_15537,N_13521,N_13130);
nor U15538 (N_15538,N_12812,N_13748);
or U15539 (N_15539,N_14520,N_14436);
and U15540 (N_15540,N_14988,N_13687);
xnor U15541 (N_15541,N_14370,N_12522);
and U15542 (N_15542,N_12859,N_13768);
and U15543 (N_15543,N_14892,N_12589);
xor U15544 (N_15544,N_14317,N_12633);
and U15545 (N_15545,N_12556,N_12623);
nor U15546 (N_15546,N_12527,N_13435);
and U15547 (N_15547,N_13538,N_12987);
and U15548 (N_15548,N_13925,N_14766);
and U15549 (N_15549,N_14680,N_13181);
and U15550 (N_15550,N_13609,N_14381);
nor U15551 (N_15551,N_13095,N_13224);
nand U15552 (N_15552,N_12569,N_14249);
or U15553 (N_15553,N_13826,N_12653);
xor U15554 (N_15554,N_13556,N_14849);
xor U15555 (N_15555,N_14107,N_13437);
xor U15556 (N_15556,N_14874,N_14530);
and U15557 (N_15557,N_13542,N_13984);
or U15558 (N_15558,N_13316,N_14417);
or U15559 (N_15559,N_12860,N_13227);
xnor U15560 (N_15560,N_12778,N_14998);
or U15561 (N_15561,N_13960,N_13295);
or U15562 (N_15562,N_13274,N_13716);
xnor U15563 (N_15563,N_14905,N_13365);
and U15564 (N_15564,N_13808,N_13729);
nand U15565 (N_15565,N_13579,N_14161);
and U15566 (N_15566,N_14824,N_13300);
nor U15567 (N_15567,N_13881,N_14642);
xor U15568 (N_15568,N_14207,N_12689);
and U15569 (N_15569,N_13871,N_14891);
or U15570 (N_15570,N_14648,N_14332);
xnor U15571 (N_15571,N_13136,N_14143);
or U15572 (N_15572,N_14990,N_13296);
nand U15573 (N_15573,N_14060,N_13084);
and U15574 (N_15574,N_14246,N_13040);
and U15575 (N_15575,N_12649,N_14882);
and U15576 (N_15576,N_14869,N_12592);
and U15577 (N_15577,N_13580,N_13694);
and U15578 (N_15578,N_13736,N_13383);
and U15579 (N_15579,N_13440,N_14817);
nand U15580 (N_15580,N_14159,N_14026);
xnor U15581 (N_15581,N_12817,N_14850);
and U15582 (N_15582,N_13520,N_12608);
nor U15583 (N_15583,N_14269,N_13671);
nor U15584 (N_15584,N_14683,N_12662);
nor U15585 (N_15585,N_14749,N_12655);
nand U15586 (N_15586,N_13839,N_12991);
and U15587 (N_15587,N_13480,N_12996);
and U15588 (N_15588,N_13781,N_14184);
nor U15589 (N_15589,N_14633,N_14092);
xor U15590 (N_15590,N_14476,N_13066);
and U15591 (N_15591,N_13153,N_13210);
and U15592 (N_15592,N_13011,N_13335);
nor U15593 (N_15593,N_13715,N_14873);
and U15594 (N_15594,N_13751,N_13528);
or U15595 (N_15595,N_14481,N_14451);
and U15596 (N_15596,N_14646,N_13912);
xnor U15597 (N_15597,N_14162,N_14854);
nor U15598 (N_15598,N_13339,N_13063);
or U15599 (N_15599,N_14807,N_13213);
nor U15600 (N_15600,N_12743,N_13519);
nor U15601 (N_15601,N_14616,N_14023);
nand U15602 (N_15602,N_13730,N_14571);
and U15603 (N_15603,N_12989,N_12821);
nor U15604 (N_15604,N_14938,N_14584);
nand U15605 (N_15605,N_14945,N_12938);
nand U15606 (N_15606,N_14140,N_13007);
or U15607 (N_15607,N_13352,N_14167);
nand U15608 (N_15608,N_14277,N_13922);
nor U15609 (N_15609,N_13999,N_14460);
xnor U15610 (N_15610,N_12609,N_12774);
and U15611 (N_15611,N_14456,N_14005);
and U15612 (N_15612,N_14101,N_13666);
nor U15613 (N_15613,N_14127,N_13809);
nand U15614 (N_15614,N_13226,N_14022);
or U15615 (N_15615,N_13825,N_12667);
or U15616 (N_15616,N_14816,N_12990);
xor U15617 (N_15617,N_14803,N_14076);
or U15618 (N_15618,N_14145,N_12568);
nand U15619 (N_15619,N_14318,N_14730);
or U15620 (N_15620,N_14639,N_14432);
nand U15621 (N_15621,N_14406,N_14856);
nor U15622 (N_15622,N_14279,N_12612);
xnor U15623 (N_15623,N_12742,N_12814);
and U15624 (N_15624,N_14108,N_14376);
nand U15625 (N_15625,N_12756,N_14924);
nor U15626 (N_15626,N_12822,N_14347);
xnor U15627 (N_15627,N_14797,N_14454);
or U15628 (N_15628,N_13636,N_14039);
or U15629 (N_15629,N_12856,N_14664);
xor U15630 (N_15630,N_14151,N_14629);
xnor U15631 (N_15631,N_13417,N_14912);
and U15632 (N_15632,N_13923,N_13669);
xnor U15633 (N_15633,N_12971,N_12509);
nand U15634 (N_15634,N_14065,N_13991);
or U15635 (N_15635,N_13291,N_14388);
nand U15636 (N_15636,N_14074,N_14030);
xnor U15637 (N_15637,N_14551,N_13575);
xor U15638 (N_15638,N_13024,N_12914);
nor U15639 (N_15639,N_14486,N_12598);
nand U15640 (N_15640,N_12529,N_14801);
or U15641 (N_15641,N_14179,N_12542);
and U15642 (N_15642,N_12943,N_14103);
xor U15643 (N_15643,N_14862,N_13901);
or U15644 (N_15644,N_14973,N_13424);
nand U15645 (N_15645,N_12832,N_14786);
or U15646 (N_15646,N_14276,N_14472);
and U15647 (N_15647,N_12630,N_13665);
nor U15648 (N_15648,N_14919,N_12578);
xor U15649 (N_15649,N_13943,N_14812);
xnor U15650 (N_15650,N_13170,N_13223);
nand U15651 (N_15651,N_13317,N_13647);
and U15652 (N_15652,N_14777,N_13103);
nand U15653 (N_15653,N_14790,N_14906);
nand U15654 (N_15654,N_12702,N_12918);
nor U15655 (N_15655,N_13140,N_13574);
nor U15656 (N_15656,N_14547,N_14283);
nand U15657 (N_15657,N_13634,N_14061);
and U15658 (N_15658,N_13540,N_13002);
xor U15659 (N_15659,N_13315,N_12982);
xnor U15660 (N_15660,N_13711,N_13200);
or U15661 (N_15661,N_12676,N_14967);
nand U15662 (N_15662,N_14210,N_14098);
nand U15663 (N_15663,N_14592,N_14138);
nand U15664 (N_15664,N_14075,N_13039);
xnor U15665 (N_15665,N_14764,N_12562);
nand U15666 (N_15666,N_12539,N_14244);
or U15667 (N_15667,N_14972,N_12640);
and U15668 (N_15668,N_12528,N_14323);
xnor U15669 (N_15669,N_14443,N_14434);
nand U15670 (N_15670,N_13633,N_12893);
and U15671 (N_15671,N_13588,N_14089);
nand U15672 (N_15672,N_14590,N_14572);
xor U15673 (N_15673,N_14100,N_13604);
nor U15674 (N_15674,N_14515,N_14870);
nand U15675 (N_15675,N_14255,N_14306);
and U15676 (N_15676,N_14232,N_12724);
xnor U15677 (N_15677,N_14695,N_13967);
nor U15678 (N_15678,N_14462,N_13362);
nand U15679 (N_15679,N_12501,N_14879);
xnor U15680 (N_15680,N_13749,N_12659);
and U15681 (N_15681,N_13262,N_14557);
and U15682 (N_15682,N_13117,N_14946);
xor U15683 (N_15683,N_14444,N_12797);
xnor U15684 (N_15684,N_14955,N_13272);
xnor U15685 (N_15685,N_13217,N_12813);
or U15686 (N_15686,N_14155,N_13717);
nor U15687 (N_15687,N_13475,N_14452);
xnor U15688 (N_15688,N_13916,N_13878);
nor U15689 (N_15689,N_12535,N_12514);
nor U15690 (N_15690,N_12896,N_12746);
nand U15691 (N_15691,N_14213,N_13247);
and U15692 (N_15692,N_14760,N_13509);
nand U15693 (N_15693,N_14033,N_12816);
and U15694 (N_15694,N_13690,N_12718);
and U15695 (N_15695,N_13380,N_14219);
or U15696 (N_15696,N_13805,N_13642);
xor U15697 (N_15697,N_13033,N_14271);
xor U15698 (N_15698,N_13985,N_14191);
and U15699 (N_15699,N_14900,N_13219);
or U15700 (N_15700,N_13615,N_12942);
nand U15701 (N_15701,N_14775,N_13778);
or U15702 (N_15702,N_13883,N_13444);
xor U15703 (N_15703,N_12688,N_13474);
nor U15704 (N_15704,N_14733,N_13572);
nor U15705 (N_15705,N_13635,N_14708);
nor U15706 (N_15706,N_12935,N_12936);
and U15707 (N_15707,N_13511,N_13791);
xor U15708 (N_15708,N_13309,N_13672);
and U15709 (N_15709,N_12564,N_13625);
xor U15710 (N_15710,N_13733,N_13552);
nor U15711 (N_15711,N_14372,N_13743);
xnor U15712 (N_15712,N_14613,N_14526);
xor U15713 (N_15713,N_14934,N_13970);
and U15714 (N_15714,N_12836,N_14596);
xnor U15715 (N_15715,N_13101,N_14980);
xnor U15716 (N_15716,N_14361,N_14968);
or U15717 (N_15717,N_12753,N_14652);
or U15718 (N_15718,N_13015,N_12851);
or U15719 (N_15719,N_13086,N_13612);
or U15720 (N_15720,N_12789,N_14984);
nor U15721 (N_15721,N_12977,N_12796);
xor U15722 (N_15722,N_14091,N_12887);
xnor U15723 (N_15723,N_13193,N_14086);
xor U15724 (N_15724,N_12573,N_13406);
or U15725 (N_15725,N_14537,N_13311);
xor U15726 (N_15726,N_14251,N_12744);
xor U15727 (N_15727,N_13500,N_14015);
and U15728 (N_15728,N_14087,N_13423);
or U15729 (N_15729,N_14865,N_14747);
nor U15730 (N_15730,N_13554,N_13416);
nand U15731 (N_15731,N_12690,N_14662);
xnor U15732 (N_15732,N_13266,N_13530);
nor U15733 (N_15733,N_13023,N_14534);
nand U15734 (N_15734,N_13936,N_14811);
or U15735 (N_15735,N_14038,N_12503);
and U15736 (N_15736,N_14224,N_14410);
or U15737 (N_15737,N_12963,N_13460);
nor U15738 (N_15738,N_13921,N_14389);
or U15739 (N_15739,N_12839,N_13986);
nand U15740 (N_15740,N_14650,N_13303);
xor U15741 (N_15741,N_14396,N_13284);
nand U15742 (N_15742,N_14516,N_14512);
nand U15743 (N_15743,N_13961,N_14297);
and U15744 (N_15744,N_12722,N_14110);
xor U15745 (N_15745,N_13673,N_12922);
or U15746 (N_15746,N_13996,N_12515);
nand U15747 (N_15747,N_14044,N_13637);
and U15748 (N_15748,N_14200,N_12629);
or U15749 (N_15749,N_14348,N_14058);
nand U15750 (N_15750,N_14688,N_14838);
nand U15751 (N_15751,N_13387,N_14851);
nand U15752 (N_15752,N_13232,N_13348);
or U15753 (N_15753,N_14333,N_13292);
nor U15754 (N_15754,N_13394,N_13037);
or U15755 (N_15755,N_12731,N_14962);
and U15756 (N_15756,N_13727,N_12908);
and U15757 (N_15757,N_13770,N_12888);
nor U15758 (N_15758,N_13294,N_14346);
or U15759 (N_15759,N_14083,N_14761);
and U15760 (N_15760,N_12747,N_14717);
and U15761 (N_15761,N_13600,N_13374);
nor U15762 (N_15762,N_13815,N_12567);
xnor U15763 (N_15763,N_14736,N_13410);
and U15764 (N_15764,N_14425,N_13343);
or U15765 (N_15765,N_13976,N_13535);
nor U15766 (N_15766,N_14935,N_13620);
nand U15767 (N_15767,N_13098,N_12687);
xnor U15768 (N_15768,N_13550,N_12679);
xor U15769 (N_15769,N_14052,N_13933);
nor U15770 (N_15770,N_14867,N_13065);
and U15771 (N_15771,N_13302,N_14175);
xnor U15772 (N_15772,N_13505,N_13336);
xor U15773 (N_15773,N_14053,N_13762);
nand U15774 (N_15774,N_13667,N_14975);
and U15775 (N_15775,N_14620,N_13070);
xnor U15776 (N_15776,N_12642,N_13595);
xor U15777 (N_15777,N_13162,N_12974);
xnor U15778 (N_15778,N_14204,N_14809);
and U15779 (N_15779,N_14243,N_13268);
nor U15780 (N_15780,N_13492,N_13662);
nand U15781 (N_15781,N_14587,N_13893);
nor U15782 (N_15782,N_14810,N_13368);
or U15783 (N_15783,N_14216,N_14170);
or U15784 (N_15784,N_14982,N_12803);
and U15785 (N_15785,N_14438,N_14981);
nor U15786 (N_15786,N_13992,N_14345);
nor U15787 (N_15787,N_14032,N_13187);
xnor U15788 (N_15788,N_12513,N_13578);
nand U15789 (N_15789,N_12548,N_12765);
xnor U15790 (N_15790,N_14491,N_13077);
nand U15791 (N_15791,N_13845,N_14218);
xor U15792 (N_15792,N_13745,N_14719);
or U15793 (N_15793,N_13719,N_14621);
or U15794 (N_15794,N_13591,N_14234);
or U15795 (N_15795,N_12907,N_12506);
nand U15796 (N_15796,N_13518,N_12972);
and U15797 (N_15797,N_13503,N_14334);
and U15798 (N_15798,N_12900,N_12686);
and U15799 (N_15799,N_13089,N_12950);
nor U15800 (N_15800,N_13092,N_14769);
nor U15801 (N_15801,N_13709,N_14525);
or U15802 (N_15802,N_14321,N_13983);
and U15803 (N_15803,N_14375,N_12998);
nand U15804 (N_15804,N_12899,N_13418);
nor U15805 (N_15805,N_14883,N_13932);
or U15806 (N_15806,N_13759,N_13099);
nor U15807 (N_15807,N_14611,N_13288);
or U15808 (N_15808,N_13477,N_13927);
or U15809 (N_15809,N_12820,N_13014);
nand U15810 (N_15810,N_12948,N_14046);
nand U15811 (N_15811,N_13544,N_13737);
nand U15812 (N_15812,N_13695,N_14950);
and U15813 (N_15813,N_14672,N_12670);
and U15814 (N_15814,N_14392,N_14095);
or U15815 (N_15815,N_13044,N_14727);
or U15816 (N_15816,N_13397,N_13000);
nand U15817 (N_15817,N_13445,N_13821);
and U15818 (N_15818,N_14336,N_13529);
and U15819 (N_15819,N_14614,N_12611);
nand U15820 (N_15820,N_13021,N_12656);
nand U15821 (N_15821,N_13804,N_12590);
xor U15822 (N_15822,N_12852,N_14993);
or U15823 (N_15823,N_13526,N_12616);
or U15824 (N_15824,N_12555,N_13938);
nor U15825 (N_15825,N_13906,N_12666);
xnor U15826 (N_15826,N_14402,N_13324);
xor U15827 (N_15827,N_14625,N_14654);
and U15828 (N_15828,N_13577,N_13559);
or U15829 (N_15829,N_13856,N_12647);
nor U15830 (N_15830,N_13885,N_14203);
nand U15831 (N_15831,N_13827,N_12559);
nand U15832 (N_15832,N_14543,N_12605);
xnor U15833 (N_15833,N_12602,N_14715);
and U15834 (N_15834,N_13443,N_13347);
nand U15835 (N_15835,N_13811,N_13345);
nand U15836 (N_15836,N_13006,N_12840);
xnor U15837 (N_15837,N_13276,N_13880);
nor U15838 (N_15838,N_14765,N_13713);
nand U15839 (N_15839,N_13981,N_13621);
xor U15840 (N_15840,N_14368,N_12560);
nand U15841 (N_15841,N_13102,N_14668);
and U15842 (N_15842,N_14173,N_14197);
and U15843 (N_15843,N_14064,N_14312);
nand U15844 (N_15844,N_14927,N_14818);
nand U15845 (N_15845,N_14545,N_14400);
and U15846 (N_15846,N_12707,N_14495);
and U15847 (N_15847,N_14407,N_14469);
xnor U15848 (N_15848,N_13446,N_14365);
nor U15849 (N_15849,N_13586,N_14233);
nor U15850 (N_15850,N_14248,N_14168);
nand U15851 (N_15851,N_14437,N_13833);
or U15852 (N_15852,N_14116,N_13792);
nand U15853 (N_15853,N_14122,N_14371);
nor U15854 (N_15854,N_13009,N_14693);
nand U15855 (N_15855,N_14475,N_14029);
and U15856 (N_15856,N_13539,N_13902);
xnor U15857 (N_15857,N_13052,N_14541);
or U15858 (N_15858,N_13229,N_14532);
xor U15859 (N_15859,N_13843,N_12575);
nand U15860 (N_15860,N_13614,N_13116);
nand U15861 (N_15861,N_14762,N_13049);
nor U15862 (N_15862,N_14136,N_13285);
xor U15863 (N_15863,N_13126,N_14580);
xor U15864 (N_15864,N_14284,N_13876);
or U15865 (N_15865,N_14059,N_13279);
and U15866 (N_15866,N_14957,N_14565);
or U15867 (N_15867,N_13293,N_13855);
xnor U15868 (N_15868,N_13386,N_14536);
xnor U15869 (N_15869,N_14553,N_12999);
nand U15870 (N_15870,N_12626,N_12697);
or U15871 (N_15871,N_12520,N_12967);
nand U15872 (N_15872,N_14182,N_13886);
and U15873 (N_15873,N_14129,N_12870);
xnor U15874 (N_15874,N_13143,N_14659);
nor U15875 (N_15875,N_14583,N_12916);
nor U15876 (N_15876,N_14691,N_14651);
and U15877 (N_15877,N_13735,N_13968);
xor U15878 (N_15878,N_13684,N_13708);
and U15879 (N_15879,N_13982,N_14222);
or U15880 (N_15880,N_13150,N_14006);
nand U15881 (N_15881,N_12952,N_13298);
or U15882 (N_15882,N_14344,N_12672);
nor U15883 (N_15883,N_14549,N_12929);
nand U15884 (N_15884,N_14897,N_13390);
nand U15885 (N_15885,N_12549,N_13541);
or U15886 (N_15886,N_13074,N_12644);
xor U15887 (N_15887,N_14877,N_14995);
and U15888 (N_15888,N_14324,N_13835);
nand U15889 (N_15889,N_13439,N_13356);
nor U15890 (N_15890,N_13013,N_14473);
and U15891 (N_15891,N_13257,N_14521);
xor U15892 (N_15892,N_14937,N_13178);
and U15893 (N_15893,N_14970,N_14686);
and U15894 (N_15894,N_13283,N_14359);
or U15895 (N_15895,N_14739,N_14463);
nor U15896 (N_15896,N_14286,N_12720);
xnor U15897 (N_15897,N_13388,N_13816);
and U15898 (N_15898,N_12785,N_14704);
nor U15899 (N_15899,N_14734,N_12895);
nand U15900 (N_15900,N_14960,N_14753);
nor U15901 (N_15901,N_12581,N_12830);
xnor U15902 (N_15902,N_12973,N_12988);
xor U15903 (N_15903,N_13944,N_13534);
and U15904 (N_15904,N_14489,N_13571);
xor U15905 (N_15905,N_14841,N_13105);
or U15906 (N_15906,N_14507,N_12828);
nand U15907 (N_15907,N_13771,N_13171);
and U15908 (N_15908,N_13763,N_13199);
nand U15909 (N_15909,N_13874,N_14568);
xor U15910 (N_15910,N_14758,N_13844);
or U15911 (N_15911,N_12691,N_14556);
or U15912 (N_15912,N_13928,N_12953);
or U15913 (N_15913,N_14102,N_13566);
and U15914 (N_15914,N_13402,N_13971);
and U15915 (N_15915,N_12673,N_14247);
nand U15916 (N_15916,N_14524,N_13147);
xor U15917 (N_15917,N_12829,N_12776);
xnor U15918 (N_15918,N_13253,N_14320);
nand U15919 (N_15919,N_14221,N_14813);
xnor U15920 (N_15920,N_14330,N_12958);
and U15921 (N_15921,N_12805,N_13834);
and U15922 (N_15922,N_12853,N_13447);
and U15923 (N_15923,N_14069,N_13159);
nand U15924 (N_15924,N_14158,N_12767);
and U15925 (N_15925,N_14156,N_13546);
nand U15926 (N_15926,N_13587,N_13924);
or U15927 (N_15927,N_14595,N_14144);
nor U15928 (N_15928,N_14644,N_13598);
and U15929 (N_15929,N_12792,N_13250);
and U15930 (N_15930,N_13382,N_14899);
xnor U15931 (N_15931,N_12678,N_14369);
nor U15932 (N_15932,N_12834,N_13470);
nor U15933 (N_15933,N_13123,N_14020);
or U15934 (N_15934,N_13055,N_13664);
or U15935 (N_15935,N_13129,N_14205);
xor U15936 (N_15936,N_12651,N_12654);
or U15937 (N_15937,N_14848,N_12565);
and U15938 (N_15938,N_13525,N_13028);
nand U15939 (N_15939,N_14135,N_14669);
or U15940 (N_15940,N_14687,N_12517);
and U15941 (N_15941,N_13753,N_13373);
or U15942 (N_15942,N_14097,N_13010);
nand U15943 (N_15943,N_13910,N_13221);
and U15944 (N_15944,N_14784,N_14656);
xnor U15945 (N_15945,N_12650,N_14414);
xnor U15946 (N_15946,N_13549,N_12729);
or U15947 (N_15947,N_14492,N_14983);
nor U15948 (N_15948,N_14752,N_12956);
nor U15949 (N_15949,N_14658,N_13087);
and U15950 (N_15950,N_14280,N_13548);
or U15951 (N_15951,N_14898,N_13202);
and U15952 (N_15952,N_12730,N_14681);
nor U15953 (N_15953,N_13256,N_14670);
nand U15954 (N_15954,N_14386,N_14910);
or U15955 (N_15955,N_14745,N_12597);
xor U15956 (N_15956,N_13602,N_13032);
nor U15957 (N_15957,N_14742,N_14105);
or U15958 (N_15958,N_12553,N_12582);
nand U15959 (N_15959,N_14710,N_13357);
nor U15960 (N_15960,N_13411,N_13502);
nor U15961 (N_15961,N_14314,N_14586);
xor U15962 (N_15962,N_13496,N_12749);
or U15963 (N_15963,N_14264,N_13497);
nor U15964 (N_15964,N_13464,N_14494);
or U15965 (N_15965,N_14133,N_14262);
or U15966 (N_15966,N_13056,N_14915);
or U15967 (N_15967,N_13780,N_14731);
xnor U15968 (N_15968,N_13106,N_14241);
xnor U15969 (N_15969,N_13801,N_14430);
and U15970 (N_15970,N_12770,N_14062);
or U15971 (N_15971,N_14188,N_14546);
nor U15972 (N_15972,N_14774,N_13093);
nand U15973 (N_15973,N_12596,N_14555);
nor U15974 (N_15974,N_13954,N_12962);
nand U15975 (N_15975,N_13700,N_13121);
xor U15976 (N_15976,N_12665,N_13941);
and U15977 (N_15977,N_14830,N_13214);
xor U15978 (N_15978,N_13677,N_13723);
or U15979 (N_15979,N_13741,N_14876);
nor U15980 (N_15980,N_14878,N_13515);
or U15981 (N_15981,N_13547,N_12512);
xor U15982 (N_15982,N_14435,N_12843);
nand U15983 (N_15983,N_14018,N_14913);
nand U15984 (N_15984,N_13919,N_14940);
and U15985 (N_15985,N_14192,N_14804);
xnor U15986 (N_15986,N_13148,N_14570);
nand U15987 (N_15987,N_14433,N_14275);
nand U15988 (N_15988,N_13487,N_13707);
nor U15989 (N_15989,N_14888,N_13824);
xnor U15990 (N_15990,N_13678,N_12723);
nand U15991 (N_15991,N_14788,N_13558);
and U15992 (N_15992,N_12986,N_14834);
nor U15993 (N_15993,N_12736,N_13775);
and U15994 (N_15994,N_13950,N_14441);
nand U15995 (N_15995,N_13641,N_13645);
or U15996 (N_15996,N_12874,N_13391);
nand U15997 (N_15997,N_12913,N_12585);
xnor U15998 (N_15998,N_14618,N_14464);
and U15999 (N_15999,N_14778,N_14858);
nor U16000 (N_16000,N_13375,N_13661);
nor U16001 (N_16001,N_12622,N_13601);
or U16002 (N_16002,N_12809,N_13030);
nand U16003 (N_16003,N_14961,N_13689);
xor U16004 (N_16004,N_13104,N_14178);
or U16005 (N_16005,N_13570,N_14641);
nor U16006 (N_16006,N_13603,N_14199);
or U16007 (N_16007,N_12808,N_13863);
or U16008 (N_16008,N_14638,N_14705);
or U16009 (N_16009,N_14226,N_14331);
nor U16010 (N_16010,N_13764,N_12579);
xor U16011 (N_16011,N_13458,N_12994);
xnor U16012 (N_16012,N_14012,N_12620);
or U16013 (N_16013,N_13583,N_13194);
nand U16014 (N_16014,N_13297,N_14124);
nand U16015 (N_16015,N_12802,N_12880);
xnor U16016 (N_16016,N_14721,N_12975);
and U16017 (N_16017,N_14355,N_14240);
nor U16018 (N_16018,N_14290,N_14081);
xor U16019 (N_16019,N_12519,N_14399);
nand U16020 (N_16020,N_14082,N_14501);
xnor U16021 (N_16021,N_13892,N_13877);
nor U16022 (N_16022,N_14859,N_13889);
nand U16023 (N_16023,N_14328,N_13660);
and U16024 (N_16024,N_14645,N_12521);
xnor U16025 (N_16025,N_13838,N_12648);
nand U16026 (N_16026,N_12636,N_14049);
and U16027 (N_16027,N_13188,N_13304);
or U16028 (N_16028,N_14889,N_12586);
xnor U16029 (N_16029,N_13125,N_13799);
nor U16030 (N_16030,N_13668,N_12621);
or U16031 (N_16031,N_14847,N_12835);
and U16032 (N_16032,N_13861,N_14907);
or U16033 (N_16033,N_14563,N_13640);
nor U16034 (N_16034,N_14996,N_13459);
nand U16035 (N_16035,N_13482,N_14840);
or U16036 (N_16036,N_13870,N_14412);
xor U16037 (N_16037,N_13699,N_13145);
xor U16038 (N_16038,N_13146,N_14931);
nand U16039 (N_16039,N_13420,N_12970);
and U16040 (N_16040,N_13860,N_13584);
nand U16041 (N_16041,N_14431,N_13896);
nor U16042 (N_16042,N_12638,N_12733);
nor U16043 (N_16043,N_13163,N_14707);
xor U16044 (N_16044,N_14268,N_13705);
nor U16045 (N_16045,N_14257,N_14930);
nor U16046 (N_16046,N_14636,N_14857);
nand U16047 (N_16047,N_14157,N_14387);
nor U16048 (N_16048,N_12745,N_14237);
nor U16049 (N_16049,N_14367,N_14394);
nor U16050 (N_16050,N_12798,N_13829);
and U16051 (N_16051,N_13524,N_13617);
xor U16052 (N_16052,N_12764,N_14265);
and U16053 (N_16053,N_13926,N_12677);
and U16054 (N_16054,N_12804,N_13355);
and U16055 (N_16055,N_14319,N_12740);
and U16056 (N_16056,N_13132,N_13180);
nor U16057 (N_16057,N_13593,N_12925);
and U16058 (N_16058,N_14619,N_14160);
xor U16059 (N_16059,N_13003,N_14880);
or U16060 (N_16060,N_14209,N_13112);
nand U16061 (N_16061,N_13494,N_13038);
nor U16062 (N_16062,N_14703,N_12795);
xor U16063 (N_16063,N_14517,N_12947);
nor U16064 (N_16064,N_13431,N_14341);
xnor U16065 (N_16065,N_13734,N_13372);
or U16066 (N_16066,N_13561,N_14964);
nand U16067 (N_16067,N_14242,N_14165);
xor U16068 (N_16068,N_13555,N_13235);
nor U16069 (N_16069,N_14947,N_13035);
and U16070 (N_16070,N_12819,N_13739);
and U16071 (N_16071,N_13430,N_14624);
and U16072 (N_16072,N_12671,N_14844);
and U16073 (N_16073,N_14831,N_13173);
and U16074 (N_16074,N_14814,N_12681);
nand U16075 (N_16075,N_13852,N_12826);
or U16076 (N_16076,N_14522,N_12793);
and U16077 (N_16077,N_12976,N_13008);
or U16078 (N_16078,N_14130,N_13005);
xor U16079 (N_16079,N_13964,N_13175);
nor U16080 (N_16080,N_12618,N_13131);
or U16081 (N_16081,N_13331,N_13124);
nand U16082 (N_16082,N_14193,N_14918);
nor U16083 (N_16083,N_12537,N_13802);
and U16084 (N_16084,N_12979,N_14607);
xnor U16085 (N_16085,N_13231,N_12572);
or U16086 (N_16086,N_14920,N_13360);
nand U16087 (N_16087,N_13978,N_14685);
nand U16088 (N_16088,N_14047,N_13264);
and U16089 (N_16089,N_14732,N_12949);
nand U16090 (N_16090,N_12600,N_14694);
nor U16091 (N_16091,N_13278,N_12505);
xor U16092 (N_16092,N_13563,N_14254);
nor U16093 (N_16093,N_14383,N_14706);
xor U16094 (N_16094,N_13107,N_13830);
or U16095 (N_16095,N_14126,N_13879);
xor U16096 (N_16096,N_12944,N_12685);
nor U16097 (N_16097,N_14612,N_14352);
or U16098 (N_16098,N_13404,N_12983);
nor U16099 (N_16099,N_13114,N_12661);
and U16100 (N_16100,N_12837,N_13862);
xnor U16101 (N_16101,N_13773,N_14630);
nand U16102 (N_16102,N_13096,N_14712);
nor U16103 (N_16103,N_14045,N_14528);
xnor U16104 (N_16104,N_13428,N_13020);
xor U16105 (N_16105,N_14245,N_14567);
nor U16106 (N_16106,N_13160,N_12669);
or U16107 (N_16107,N_12771,N_13205);
nand U16108 (N_16108,N_13498,N_14349);
or U16109 (N_16109,N_14142,N_14373);
nor U16110 (N_16110,N_13308,N_14770);
xnor U16111 (N_16111,N_14952,N_13341);
xor U16112 (N_16112,N_12588,N_14702);
and U16113 (N_16113,N_12660,N_13674);
xnor U16114 (N_16114,N_13945,N_13784);
xnor U16115 (N_16115,N_13965,N_14887);
xor U16116 (N_16116,N_14585,N_14866);
and U16117 (N_16117,N_13218,N_13342);
and U16118 (N_16118,N_14342,N_13710);
nor U16119 (N_16119,N_13623,N_14994);
and U16120 (N_16120,N_14322,N_14904);
and U16121 (N_16121,N_14725,N_14533);
nor U16122 (N_16122,N_13400,N_12762);
or U16123 (N_16123,N_13891,N_13321);
and U16124 (N_16124,N_14017,N_13467);
nor U16125 (N_16125,N_13436,N_13622);
nor U16126 (N_16126,N_14600,N_14294);
nor U16127 (N_16127,N_13899,N_14266);
xor U16128 (N_16128,N_14415,N_12606);
nor U16129 (N_16129,N_12645,N_12844);
and U16130 (N_16130,N_12577,N_13783);
nand U16131 (N_16131,N_12668,N_12867);
or U16132 (N_16132,N_12886,N_14606);
nor U16133 (N_16133,N_12783,N_13490);
nand U16134 (N_16134,N_14701,N_14358);
or U16135 (N_16135,N_12788,N_13789);
nor U16136 (N_16136,N_13853,N_13873);
nor U16137 (N_16137,N_13004,N_14832);
or U16138 (N_16138,N_14115,N_12566);
and U16139 (N_16139,N_13370,N_12824);
nand U16140 (N_16140,N_14944,N_13553);
xnor U16141 (N_16141,N_13628,N_14181);
or U16142 (N_16142,N_14364,N_13337);
nand U16143 (N_16143,N_14554,N_12751);
nor U16144 (N_16144,N_14339,N_14647);
nor U16145 (N_16145,N_14206,N_14189);
nand U16146 (N_16146,N_13018,N_14149);
xnor U16147 (N_16147,N_13940,N_13557);
nor U16148 (N_16148,N_14789,N_13966);
nand U16149 (N_16149,N_14754,N_12875);
or U16150 (N_16150,N_13407,N_14458);
and U16151 (N_16151,N_14413,N_13513);
nand U16152 (N_16152,N_13670,N_14172);
and U16153 (N_16153,N_13249,N_14093);
or U16154 (N_16154,N_12646,N_12704);
nand U16155 (N_16155,N_12984,N_12934);
or U16156 (N_16156,N_14305,N_13141);
nand U16157 (N_16157,N_14252,N_14959);
nor U16158 (N_16158,N_14043,N_14397);
nor U16159 (N_16159,N_14936,N_12735);
or U16160 (N_16160,N_13327,N_13334);
or U16161 (N_16161,N_14723,N_13585);
or U16162 (N_16162,N_12845,N_13017);
xor U16163 (N_16163,N_13481,N_12831);
and U16164 (N_16164,N_14627,N_14928);
and U16165 (N_16165,N_13463,N_14776);
and U16166 (N_16166,N_14176,N_13814);
and U16167 (N_16167,N_13624,N_12946);
xnor U16168 (N_16168,N_14653,N_12610);
nand U16169 (N_16169,N_13618,N_12541);
or U16170 (N_16170,N_12719,N_14118);
and U16171 (N_16171,N_14690,N_14643);
or U16172 (N_16172,N_14420,N_13951);
or U16173 (N_16173,N_12905,N_14311);
nor U16174 (N_16174,N_13195,N_14042);
nand U16175 (N_16175,N_13412,N_14843);
nand U16176 (N_16176,N_12700,N_13888);
and U16177 (N_16177,N_13471,N_13504);
nand U16178 (N_16178,N_13972,N_12760);
and U16179 (N_16179,N_12526,N_13508);
or U16180 (N_16180,N_13953,N_12921);
nand U16181 (N_16181,N_12617,N_13270);
and U16182 (N_16182,N_13488,N_14238);
nand U16183 (N_16183,N_14487,N_14000);
xor U16184 (N_16184,N_13722,N_12698);
and U16185 (N_16185,N_13060,N_14153);
xor U16186 (N_16186,N_14488,N_13120);
nand U16187 (N_16187,N_14125,N_14111);
or U16188 (N_16188,N_14187,N_13275);
nand U16189 (N_16189,N_13864,N_13115);
and U16190 (N_16190,N_13452,N_14718);
xor U16191 (N_16191,N_13937,N_14561);
nand U16192 (N_16192,N_13686,N_13434);
xor U16193 (N_16193,N_14360,N_12664);
nor U16194 (N_16194,N_14604,N_13682);
or U16195 (N_16195,N_14002,N_13413);
and U16196 (N_16196,N_14301,N_14634);
nand U16197 (N_16197,N_13865,N_13952);
nand U16198 (N_16198,N_14663,N_14343);
nor U16199 (N_16199,N_14958,N_14833);
or U16200 (N_16200,N_13903,N_14404);
nor U16201 (N_16201,N_14976,N_13142);
xor U16202 (N_16202,N_14550,N_14966);
xor U16203 (N_16203,N_14267,N_14744);
nor U16204 (N_16204,N_14773,N_13963);
xnor U16205 (N_16205,N_12547,N_14626);
xnor U16206 (N_16206,N_14479,N_13027);
and U16207 (N_16207,N_14917,N_13704);
or U16208 (N_16208,N_14798,N_13568);
nand U16209 (N_16209,N_14429,N_14239);
xnor U16210 (N_16210,N_14674,N_13626);
and U16211 (N_16211,N_13489,N_13619);
or U16212 (N_16212,N_14011,N_12981);
nand U16213 (N_16213,N_12755,N_14513);
and U16214 (N_16214,N_13371,N_14037);
xnor U16215 (N_16215,N_13738,N_12643);
and U16216 (N_16216,N_14610,N_13758);
nand U16217 (N_16217,N_12904,N_13468);
nand U16218 (N_16218,N_14325,N_13239);
and U16219 (N_16219,N_12750,N_13211);
and U16220 (N_16220,N_14198,N_14285);
nor U16221 (N_16221,N_13091,N_12710);
nor U16222 (N_16222,N_14519,N_12591);
xnor U16223 (N_16223,N_14787,N_13904);
and U16224 (N_16224,N_12833,N_14177);
nand U16225 (N_16225,N_13118,N_13236);
nand U16226 (N_16226,N_14292,N_13057);
nand U16227 (N_16227,N_13108,N_13698);
nor U16228 (N_16228,N_14746,N_13313);
or U16229 (N_16229,N_13772,N_13800);
or U16230 (N_16230,N_14529,N_14531);
nor U16231 (N_16231,N_13947,N_14295);
and U16232 (N_16232,N_12915,N_12693);
xor U16233 (N_16233,N_14860,N_14003);
or U16234 (N_16234,N_13109,N_14195);
or U16235 (N_16235,N_13681,N_13307);
or U16236 (N_16236,N_14577,N_13828);
xnor U16237 (N_16237,N_14309,N_13989);
nor U16238 (N_16238,N_14578,N_14104);
xor U16239 (N_16239,N_12966,N_13133);
or U16240 (N_16240,N_12625,N_13979);
or U16241 (N_16241,N_13797,N_13486);
nor U16242 (N_16242,N_14291,N_14977);
nor U16243 (N_16243,N_12933,N_12878);
nand U16244 (N_16244,N_12576,N_14048);
xor U16245 (N_16245,N_14609,N_12545);
and U16246 (N_16246,N_14796,N_14617);
nor U16247 (N_16247,N_13222,N_14985);
nor U16248 (N_16248,N_13848,N_13401);
nand U16249 (N_16249,N_13720,N_14031);
nand U16250 (N_16250,N_13041,N_14788);
nor U16251 (N_16251,N_13228,N_14081);
nor U16252 (N_16252,N_13692,N_12816);
nand U16253 (N_16253,N_14412,N_14404);
nand U16254 (N_16254,N_13555,N_14354);
xnor U16255 (N_16255,N_13741,N_14339);
or U16256 (N_16256,N_13618,N_14687);
and U16257 (N_16257,N_14798,N_14337);
and U16258 (N_16258,N_13639,N_14424);
or U16259 (N_16259,N_14013,N_14901);
or U16260 (N_16260,N_14608,N_14992);
nand U16261 (N_16261,N_14892,N_13229);
or U16262 (N_16262,N_14346,N_14421);
and U16263 (N_16263,N_14486,N_13003);
xnor U16264 (N_16264,N_12926,N_13516);
nand U16265 (N_16265,N_13258,N_13125);
and U16266 (N_16266,N_13457,N_13741);
and U16267 (N_16267,N_14055,N_14862);
xor U16268 (N_16268,N_13067,N_12902);
nand U16269 (N_16269,N_14915,N_14835);
and U16270 (N_16270,N_13733,N_13918);
or U16271 (N_16271,N_12641,N_13356);
and U16272 (N_16272,N_14422,N_14961);
or U16273 (N_16273,N_14834,N_14977);
or U16274 (N_16274,N_14908,N_13235);
nor U16275 (N_16275,N_13847,N_12638);
and U16276 (N_16276,N_14128,N_13182);
nand U16277 (N_16277,N_14080,N_13117);
and U16278 (N_16278,N_12588,N_14578);
nand U16279 (N_16279,N_13047,N_14390);
xor U16280 (N_16280,N_12726,N_13325);
nor U16281 (N_16281,N_13987,N_14055);
nor U16282 (N_16282,N_14902,N_14038);
and U16283 (N_16283,N_14880,N_12847);
nor U16284 (N_16284,N_13323,N_13126);
nor U16285 (N_16285,N_14657,N_14055);
nor U16286 (N_16286,N_12925,N_13137);
nor U16287 (N_16287,N_14392,N_12539);
nor U16288 (N_16288,N_13925,N_12901);
and U16289 (N_16289,N_13275,N_13711);
xor U16290 (N_16290,N_13852,N_12782);
or U16291 (N_16291,N_14846,N_14082);
and U16292 (N_16292,N_14305,N_14528);
xnor U16293 (N_16293,N_14870,N_14789);
nor U16294 (N_16294,N_13072,N_14194);
xnor U16295 (N_16295,N_14011,N_13517);
nor U16296 (N_16296,N_14989,N_14843);
nand U16297 (N_16297,N_14318,N_13286);
nand U16298 (N_16298,N_14500,N_13410);
or U16299 (N_16299,N_13210,N_13449);
or U16300 (N_16300,N_13505,N_14760);
or U16301 (N_16301,N_13346,N_13806);
nand U16302 (N_16302,N_14781,N_13187);
nor U16303 (N_16303,N_14500,N_12600);
nor U16304 (N_16304,N_13724,N_13003);
nor U16305 (N_16305,N_13394,N_14942);
xor U16306 (N_16306,N_13392,N_12705);
nand U16307 (N_16307,N_14651,N_14987);
nand U16308 (N_16308,N_12710,N_13917);
nor U16309 (N_16309,N_14004,N_12548);
xnor U16310 (N_16310,N_12586,N_12717);
xnor U16311 (N_16311,N_12711,N_14091);
and U16312 (N_16312,N_13573,N_13418);
or U16313 (N_16313,N_14515,N_14541);
nor U16314 (N_16314,N_12602,N_12603);
xor U16315 (N_16315,N_13941,N_13406);
and U16316 (N_16316,N_14814,N_13970);
nand U16317 (N_16317,N_12665,N_14630);
nand U16318 (N_16318,N_13447,N_12990);
xor U16319 (N_16319,N_14576,N_13306);
nor U16320 (N_16320,N_14642,N_12784);
xnor U16321 (N_16321,N_13499,N_13110);
nand U16322 (N_16322,N_12821,N_14461);
nand U16323 (N_16323,N_13638,N_14168);
nand U16324 (N_16324,N_12924,N_12689);
or U16325 (N_16325,N_14051,N_12984);
or U16326 (N_16326,N_12928,N_12854);
xnor U16327 (N_16327,N_13122,N_13147);
and U16328 (N_16328,N_14075,N_12501);
or U16329 (N_16329,N_13116,N_14984);
nand U16330 (N_16330,N_14926,N_14739);
nand U16331 (N_16331,N_14040,N_14395);
nand U16332 (N_16332,N_14474,N_12519);
nor U16333 (N_16333,N_14711,N_14394);
xnor U16334 (N_16334,N_13682,N_14320);
xnor U16335 (N_16335,N_14758,N_12927);
nand U16336 (N_16336,N_13951,N_14238);
and U16337 (N_16337,N_14274,N_12899);
nor U16338 (N_16338,N_13863,N_14700);
or U16339 (N_16339,N_13973,N_14959);
and U16340 (N_16340,N_14660,N_12977);
and U16341 (N_16341,N_13679,N_14712);
or U16342 (N_16342,N_13387,N_12868);
nand U16343 (N_16343,N_14603,N_12641);
nor U16344 (N_16344,N_13620,N_14911);
xor U16345 (N_16345,N_13277,N_14144);
nand U16346 (N_16346,N_12979,N_13259);
or U16347 (N_16347,N_13590,N_13738);
xnor U16348 (N_16348,N_13615,N_14540);
xor U16349 (N_16349,N_13244,N_14499);
xor U16350 (N_16350,N_13593,N_14840);
nand U16351 (N_16351,N_14165,N_14556);
nand U16352 (N_16352,N_13060,N_14750);
or U16353 (N_16353,N_14253,N_14283);
nand U16354 (N_16354,N_13497,N_13293);
xnor U16355 (N_16355,N_14638,N_13212);
xor U16356 (N_16356,N_12960,N_12746);
or U16357 (N_16357,N_14942,N_14473);
nor U16358 (N_16358,N_13571,N_13989);
nor U16359 (N_16359,N_14763,N_14707);
and U16360 (N_16360,N_14432,N_14777);
nor U16361 (N_16361,N_14904,N_13094);
nand U16362 (N_16362,N_13247,N_13440);
nor U16363 (N_16363,N_13645,N_14398);
and U16364 (N_16364,N_12601,N_12790);
nor U16365 (N_16365,N_13434,N_12817);
xor U16366 (N_16366,N_13057,N_14854);
xor U16367 (N_16367,N_13851,N_13537);
nand U16368 (N_16368,N_13183,N_13129);
or U16369 (N_16369,N_13999,N_13437);
nand U16370 (N_16370,N_13937,N_14747);
and U16371 (N_16371,N_13123,N_14578);
nand U16372 (N_16372,N_13386,N_14643);
or U16373 (N_16373,N_12932,N_14194);
and U16374 (N_16374,N_13167,N_13921);
nor U16375 (N_16375,N_14892,N_13860);
xnor U16376 (N_16376,N_14722,N_12568);
nor U16377 (N_16377,N_14538,N_14049);
nand U16378 (N_16378,N_13833,N_13652);
xnor U16379 (N_16379,N_14662,N_14133);
and U16380 (N_16380,N_14500,N_13720);
and U16381 (N_16381,N_13260,N_14980);
nor U16382 (N_16382,N_13846,N_14368);
nand U16383 (N_16383,N_14553,N_14875);
nor U16384 (N_16384,N_14102,N_14056);
nand U16385 (N_16385,N_13838,N_12985);
or U16386 (N_16386,N_12816,N_12822);
or U16387 (N_16387,N_12567,N_12873);
and U16388 (N_16388,N_14854,N_13178);
or U16389 (N_16389,N_12837,N_12765);
or U16390 (N_16390,N_13996,N_13968);
and U16391 (N_16391,N_12881,N_13184);
or U16392 (N_16392,N_12850,N_13236);
nor U16393 (N_16393,N_13358,N_14573);
and U16394 (N_16394,N_13666,N_13137);
or U16395 (N_16395,N_13948,N_13059);
or U16396 (N_16396,N_12514,N_14477);
or U16397 (N_16397,N_14411,N_14069);
nand U16398 (N_16398,N_13065,N_13058);
xor U16399 (N_16399,N_13791,N_12961);
or U16400 (N_16400,N_14225,N_13855);
nand U16401 (N_16401,N_12873,N_13640);
nand U16402 (N_16402,N_13500,N_13003);
nand U16403 (N_16403,N_13899,N_14785);
or U16404 (N_16404,N_13372,N_14193);
and U16405 (N_16405,N_13246,N_13505);
nor U16406 (N_16406,N_14359,N_13002);
or U16407 (N_16407,N_13368,N_13036);
and U16408 (N_16408,N_12900,N_14413);
and U16409 (N_16409,N_14140,N_12756);
or U16410 (N_16410,N_13981,N_13457);
nor U16411 (N_16411,N_14698,N_12847);
nor U16412 (N_16412,N_14715,N_12828);
or U16413 (N_16413,N_12715,N_13168);
or U16414 (N_16414,N_13023,N_13534);
nor U16415 (N_16415,N_13173,N_13537);
and U16416 (N_16416,N_12608,N_14005);
nor U16417 (N_16417,N_13739,N_14862);
xnor U16418 (N_16418,N_13802,N_13339);
or U16419 (N_16419,N_13756,N_14515);
and U16420 (N_16420,N_12624,N_13845);
nand U16421 (N_16421,N_12536,N_12836);
or U16422 (N_16422,N_14364,N_12894);
and U16423 (N_16423,N_14425,N_13577);
or U16424 (N_16424,N_12857,N_13791);
nor U16425 (N_16425,N_13957,N_14021);
and U16426 (N_16426,N_12719,N_13367);
and U16427 (N_16427,N_13767,N_14225);
or U16428 (N_16428,N_14673,N_13137);
or U16429 (N_16429,N_13333,N_14290);
and U16430 (N_16430,N_14152,N_12744);
and U16431 (N_16431,N_13097,N_13745);
xor U16432 (N_16432,N_13327,N_13079);
nor U16433 (N_16433,N_12945,N_14745);
or U16434 (N_16434,N_14805,N_13728);
or U16435 (N_16435,N_13503,N_13074);
xnor U16436 (N_16436,N_12767,N_14955);
nor U16437 (N_16437,N_13790,N_12583);
nand U16438 (N_16438,N_14828,N_12669);
nor U16439 (N_16439,N_13450,N_14531);
nor U16440 (N_16440,N_14653,N_13672);
nand U16441 (N_16441,N_13805,N_12949);
and U16442 (N_16442,N_13712,N_14849);
nor U16443 (N_16443,N_14239,N_13377);
or U16444 (N_16444,N_14319,N_14118);
nor U16445 (N_16445,N_14834,N_12955);
nand U16446 (N_16446,N_12620,N_14390);
nand U16447 (N_16447,N_14991,N_13369);
nand U16448 (N_16448,N_14678,N_14291);
and U16449 (N_16449,N_12517,N_14128);
or U16450 (N_16450,N_13247,N_13356);
and U16451 (N_16451,N_13276,N_13275);
xnor U16452 (N_16452,N_12838,N_13991);
xor U16453 (N_16453,N_13171,N_13098);
and U16454 (N_16454,N_14750,N_13441);
and U16455 (N_16455,N_13711,N_13674);
or U16456 (N_16456,N_13472,N_13131);
and U16457 (N_16457,N_14174,N_14539);
nand U16458 (N_16458,N_12979,N_14830);
or U16459 (N_16459,N_14259,N_14121);
xor U16460 (N_16460,N_13727,N_14126);
nand U16461 (N_16461,N_13114,N_12903);
nor U16462 (N_16462,N_12581,N_13059);
xor U16463 (N_16463,N_13967,N_12780);
nor U16464 (N_16464,N_13775,N_12822);
nand U16465 (N_16465,N_14263,N_14200);
nor U16466 (N_16466,N_12855,N_14658);
or U16467 (N_16467,N_14165,N_13142);
and U16468 (N_16468,N_14632,N_14993);
nor U16469 (N_16469,N_13828,N_13986);
or U16470 (N_16470,N_13350,N_13364);
nor U16471 (N_16471,N_12920,N_13819);
nor U16472 (N_16472,N_12588,N_13897);
nor U16473 (N_16473,N_13377,N_14223);
and U16474 (N_16474,N_12714,N_12957);
and U16475 (N_16475,N_13334,N_12593);
nand U16476 (N_16476,N_14832,N_14784);
nand U16477 (N_16477,N_12645,N_14877);
and U16478 (N_16478,N_12958,N_12973);
nor U16479 (N_16479,N_13666,N_14761);
nor U16480 (N_16480,N_14533,N_13147);
nor U16481 (N_16481,N_13542,N_12967);
or U16482 (N_16482,N_12768,N_13470);
or U16483 (N_16483,N_14628,N_13514);
xor U16484 (N_16484,N_14904,N_13839);
or U16485 (N_16485,N_13441,N_13229);
nor U16486 (N_16486,N_14873,N_13796);
xnor U16487 (N_16487,N_13155,N_14177);
and U16488 (N_16488,N_14152,N_14870);
xor U16489 (N_16489,N_13800,N_14389);
nor U16490 (N_16490,N_12509,N_13558);
nand U16491 (N_16491,N_14135,N_13554);
and U16492 (N_16492,N_13895,N_14555);
nor U16493 (N_16493,N_14127,N_12505);
xor U16494 (N_16494,N_13212,N_12769);
nand U16495 (N_16495,N_13282,N_13677);
xor U16496 (N_16496,N_12517,N_14941);
xor U16497 (N_16497,N_13338,N_14297);
xor U16498 (N_16498,N_14406,N_13370);
or U16499 (N_16499,N_13926,N_14567);
and U16500 (N_16500,N_14610,N_14537);
nand U16501 (N_16501,N_13307,N_14420);
xnor U16502 (N_16502,N_12795,N_13482);
nand U16503 (N_16503,N_13630,N_14915);
and U16504 (N_16504,N_13965,N_14855);
and U16505 (N_16505,N_14020,N_14205);
nand U16506 (N_16506,N_14053,N_13510);
or U16507 (N_16507,N_12605,N_13232);
nor U16508 (N_16508,N_13990,N_12686);
nand U16509 (N_16509,N_12621,N_14613);
or U16510 (N_16510,N_14385,N_12845);
or U16511 (N_16511,N_14549,N_13113);
or U16512 (N_16512,N_14114,N_14017);
and U16513 (N_16513,N_13767,N_13915);
and U16514 (N_16514,N_14877,N_14641);
nor U16515 (N_16515,N_12896,N_13620);
and U16516 (N_16516,N_13931,N_13674);
nor U16517 (N_16517,N_13140,N_12502);
nor U16518 (N_16518,N_14050,N_13965);
xnor U16519 (N_16519,N_14951,N_14755);
xor U16520 (N_16520,N_14820,N_14828);
nor U16521 (N_16521,N_12587,N_14453);
nand U16522 (N_16522,N_13346,N_14361);
xor U16523 (N_16523,N_13508,N_13947);
xor U16524 (N_16524,N_13951,N_14822);
xnor U16525 (N_16525,N_14862,N_14942);
or U16526 (N_16526,N_13853,N_14276);
nor U16527 (N_16527,N_12631,N_13486);
nor U16528 (N_16528,N_13414,N_14120);
or U16529 (N_16529,N_12720,N_14746);
nor U16530 (N_16530,N_14447,N_13173);
and U16531 (N_16531,N_12727,N_13695);
nand U16532 (N_16532,N_13441,N_14796);
nor U16533 (N_16533,N_13885,N_14262);
nand U16534 (N_16534,N_12784,N_12878);
and U16535 (N_16535,N_14407,N_12664);
or U16536 (N_16536,N_13702,N_13617);
nand U16537 (N_16537,N_12663,N_14693);
or U16538 (N_16538,N_13496,N_12803);
xor U16539 (N_16539,N_13510,N_13760);
nor U16540 (N_16540,N_12959,N_14818);
or U16541 (N_16541,N_14912,N_13401);
and U16542 (N_16542,N_14516,N_14513);
nand U16543 (N_16543,N_12743,N_13896);
nor U16544 (N_16544,N_13368,N_13254);
nand U16545 (N_16545,N_12861,N_13957);
nor U16546 (N_16546,N_12663,N_14186);
xnor U16547 (N_16547,N_14188,N_13968);
nor U16548 (N_16548,N_14901,N_13172);
and U16549 (N_16549,N_14109,N_13938);
and U16550 (N_16550,N_13767,N_14954);
or U16551 (N_16551,N_14664,N_12963);
and U16552 (N_16552,N_13791,N_13036);
or U16553 (N_16553,N_13205,N_13669);
nor U16554 (N_16554,N_13535,N_14592);
nand U16555 (N_16555,N_14903,N_14075);
or U16556 (N_16556,N_14588,N_13868);
xnor U16557 (N_16557,N_12957,N_13905);
or U16558 (N_16558,N_12985,N_14128);
xor U16559 (N_16559,N_12582,N_14586);
nand U16560 (N_16560,N_12695,N_13577);
or U16561 (N_16561,N_14127,N_13401);
and U16562 (N_16562,N_12596,N_13944);
and U16563 (N_16563,N_13082,N_14681);
and U16564 (N_16564,N_14468,N_14008);
xor U16565 (N_16565,N_12934,N_14722);
nor U16566 (N_16566,N_14802,N_12940);
xnor U16567 (N_16567,N_14750,N_12879);
xor U16568 (N_16568,N_13229,N_13633);
or U16569 (N_16569,N_12683,N_13874);
xor U16570 (N_16570,N_13053,N_13286);
xnor U16571 (N_16571,N_13027,N_12644);
xnor U16572 (N_16572,N_12663,N_13173);
nand U16573 (N_16573,N_13139,N_14537);
nand U16574 (N_16574,N_13004,N_13466);
xor U16575 (N_16575,N_13746,N_13568);
nand U16576 (N_16576,N_13032,N_13895);
nor U16577 (N_16577,N_14728,N_12696);
nand U16578 (N_16578,N_12838,N_14919);
and U16579 (N_16579,N_13221,N_13012);
xor U16580 (N_16580,N_14799,N_14428);
and U16581 (N_16581,N_14658,N_12648);
xor U16582 (N_16582,N_14620,N_12779);
and U16583 (N_16583,N_13550,N_13167);
and U16584 (N_16584,N_14878,N_13714);
and U16585 (N_16585,N_13600,N_13725);
xnor U16586 (N_16586,N_13787,N_12620);
nor U16587 (N_16587,N_12924,N_14211);
xor U16588 (N_16588,N_13184,N_14586);
xnor U16589 (N_16589,N_12795,N_13166);
nand U16590 (N_16590,N_13309,N_13001);
xnor U16591 (N_16591,N_12943,N_13308);
nand U16592 (N_16592,N_12897,N_13573);
nand U16593 (N_16593,N_14272,N_14944);
xnor U16594 (N_16594,N_13852,N_13797);
and U16595 (N_16595,N_12698,N_14565);
xor U16596 (N_16596,N_13641,N_13026);
or U16597 (N_16597,N_13123,N_12533);
xor U16598 (N_16598,N_14230,N_13291);
or U16599 (N_16599,N_13991,N_14427);
nand U16600 (N_16600,N_14257,N_14904);
or U16601 (N_16601,N_14131,N_14380);
nand U16602 (N_16602,N_14673,N_12522);
nor U16603 (N_16603,N_13593,N_14241);
and U16604 (N_16604,N_14899,N_14011);
nand U16605 (N_16605,N_14431,N_13379);
or U16606 (N_16606,N_13856,N_14357);
and U16607 (N_16607,N_13166,N_14136);
xnor U16608 (N_16608,N_14647,N_13548);
nand U16609 (N_16609,N_14879,N_13676);
nor U16610 (N_16610,N_12565,N_13095);
nor U16611 (N_16611,N_13483,N_13132);
nor U16612 (N_16612,N_12985,N_12876);
nand U16613 (N_16613,N_14406,N_14151);
and U16614 (N_16614,N_13285,N_14115);
xor U16615 (N_16615,N_14566,N_14688);
or U16616 (N_16616,N_13258,N_13590);
and U16617 (N_16617,N_13673,N_13711);
and U16618 (N_16618,N_14404,N_13495);
xor U16619 (N_16619,N_12631,N_12558);
and U16620 (N_16620,N_14020,N_13237);
nor U16621 (N_16621,N_13981,N_13877);
or U16622 (N_16622,N_14811,N_12669);
nor U16623 (N_16623,N_12667,N_13413);
and U16624 (N_16624,N_13622,N_13013);
and U16625 (N_16625,N_12680,N_13872);
nand U16626 (N_16626,N_13084,N_13831);
or U16627 (N_16627,N_14659,N_14741);
xnor U16628 (N_16628,N_12552,N_14081);
nor U16629 (N_16629,N_14771,N_13755);
or U16630 (N_16630,N_13621,N_13670);
and U16631 (N_16631,N_13251,N_14765);
and U16632 (N_16632,N_14739,N_12672);
nand U16633 (N_16633,N_13010,N_14182);
nand U16634 (N_16634,N_14328,N_13091);
xnor U16635 (N_16635,N_14202,N_14806);
nand U16636 (N_16636,N_13864,N_13372);
nor U16637 (N_16637,N_12904,N_14959);
nor U16638 (N_16638,N_12682,N_13124);
xnor U16639 (N_16639,N_12587,N_14323);
and U16640 (N_16640,N_12840,N_13628);
nor U16641 (N_16641,N_14933,N_12893);
xnor U16642 (N_16642,N_13327,N_14186);
and U16643 (N_16643,N_13493,N_12830);
or U16644 (N_16644,N_13492,N_14207);
nand U16645 (N_16645,N_13507,N_12588);
nand U16646 (N_16646,N_14963,N_13481);
and U16647 (N_16647,N_12710,N_14806);
xor U16648 (N_16648,N_14579,N_12933);
or U16649 (N_16649,N_14458,N_14337);
nand U16650 (N_16650,N_14830,N_13258);
nor U16651 (N_16651,N_12745,N_13269);
nor U16652 (N_16652,N_13012,N_12941);
xor U16653 (N_16653,N_14094,N_12603);
nand U16654 (N_16654,N_14330,N_14121);
and U16655 (N_16655,N_14977,N_13657);
nor U16656 (N_16656,N_13228,N_13235);
xnor U16657 (N_16657,N_13366,N_14020);
nor U16658 (N_16658,N_12811,N_14633);
and U16659 (N_16659,N_13793,N_14369);
nand U16660 (N_16660,N_12967,N_13031);
xnor U16661 (N_16661,N_13225,N_14330);
nand U16662 (N_16662,N_14454,N_13047);
nor U16663 (N_16663,N_13702,N_13051);
nand U16664 (N_16664,N_13074,N_14903);
nand U16665 (N_16665,N_14921,N_14289);
nor U16666 (N_16666,N_13309,N_13104);
xnor U16667 (N_16667,N_13969,N_12592);
or U16668 (N_16668,N_13433,N_14801);
xor U16669 (N_16669,N_14536,N_12522);
nor U16670 (N_16670,N_14362,N_13267);
xor U16671 (N_16671,N_12962,N_14550);
nor U16672 (N_16672,N_14198,N_14811);
xnor U16673 (N_16673,N_13584,N_14471);
or U16674 (N_16674,N_13258,N_14272);
nor U16675 (N_16675,N_14082,N_14629);
xor U16676 (N_16676,N_13453,N_13954);
nor U16677 (N_16677,N_14480,N_12676);
and U16678 (N_16678,N_12527,N_14316);
xnor U16679 (N_16679,N_14865,N_13183);
or U16680 (N_16680,N_14054,N_14165);
and U16681 (N_16681,N_13064,N_14912);
and U16682 (N_16682,N_14326,N_13264);
xor U16683 (N_16683,N_14615,N_12837);
or U16684 (N_16684,N_13176,N_12589);
nor U16685 (N_16685,N_14479,N_14409);
or U16686 (N_16686,N_13367,N_12708);
and U16687 (N_16687,N_14073,N_14023);
nor U16688 (N_16688,N_13697,N_14245);
or U16689 (N_16689,N_13813,N_12706);
and U16690 (N_16690,N_13368,N_13387);
or U16691 (N_16691,N_12661,N_12570);
nand U16692 (N_16692,N_13048,N_12555);
nor U16693 (N_16693,N_13920,N_13808);
or U16694 (N_16694,N_14502,N_14756);
xor U16695 (N_16695,N_13046,N_14517);
xor U16696 (N_16696,N_13905,N_14069);
nand U16697 (N_16697,N_14739,N_14340);
nor U16698 (N_16698,N_12880,N_12920);
or U16699 (N_16699,N_14797,N_13047);
nand U16700 (N_16700,N_14269,N_14499);
nand U16701 (N_16701,N_14324,N_14802);
xor U16702 (N_16702,N_14329,N_13820);
nand U16703 (N_16703,N_14953,N_14151);
nor U16704 (N_16704,N_14075,N_14599);
or U16705 (N_16705,N_14633,N_12861);
xor U16706 (N_16706,N_14884,N_12887);
nand U16707 (N_16707,N_14597,N_14989);
xor U16708 (N_16708,N_13273,N_14815);
nand U16709 (N_16709,N_14698,N_14974);
or U16710 (N_16710,N_13264,N_13469);
xnor U16711 (N_16711,N_14436,N_13834);
nor U16712 (N_16712,N_14381,N_13772);
nand U16713 (N_16713,N_13629,N_12575);
nor U16714 (N_16714,N_12873,N_13552);
nand U16715 (N_16715,N_14643,N_14513);
or U16716 (N_16716,N_12754,N_14129);
xor U16717 (N_16717,N_13983,N_14924);
xor U16718 (N_16718,N_14397,N_12778);
nand U16719 (N_16719,N_13317,N_14530);
or U16720 (N_16720,N_12871,N_14058);
nor U16721 (N_16721,N_12699,N_13106);
nand U16722 (N_16722,N_13959,N_14999);
xnor U16723 (N_16723,N_12716,N_14550);
nor U16724 (N_16724,N_13879,N_13913);
and U16725 (N_16725,N_14438,N_14107);
and U16726 (N_16726,N_13513,N_13247);
xor U16727 (N_16727,N_14913,N_13553);
and U16728 (N_16728,N_14521,N_13321);
xor U16729 (N_16729,N_13560,N_13455);
or U16730 (N_16730,N_12746,N_13613);
or U16731 (N_16731,N_13858,N_14147);
nor U16732 (N_16732,N_14546,N_12720);
and U16733 (N_16733,N_14005,N_14995);
and U16734 (N_16734,N_14811,N_14755);
nand U16735 (N_16735,N_13895,N_14281);
nor U16736 (N_16736,N_13800,N_13071);
and U16737 (N_16737,N_14854,N_13593);
xor U16738 (N_16738,N_14285,N_14224);
nand U16739 (N_16739,N_13331,N_14533);
nand U16740 (N_16740,N_13954,N_12668);
nor U16741 (N_16741,N_13126,N_14438);
xor U16742 (N_16742,N_14522,N_13265);
and U16743 (N_16743,N_12552,N_12777);
or U16744 (N_16744,N_14451,N_14933);
nand U16745 (N_16745,N_13412,N_14259);
or U16746 (N_16746,N_14006,N_13765);
nor U16747 (N_16747,N_12648,N_14619);
nor U16748 (N_16748,N_13308,N_13046);
and U16749 (N_16749,N_14360,N_13293);
nor U16750 (N_16750,N_14980,N_13306);
and U16751 (N_16751,N_14470,N_13619);
nand U16752 (N_16752,N_13148,N_14426);
nand U16753 (N_16753,N_13094,N_12896);
or U16754 (N_16754,N_13734,N_13663);
nand U16755 (N_16755,N_14268,N_12576);
nand U16756 (N_16756,N_12787,N_13883);
or U16757 (N_16757,N_13268,N_13063);
nand U16758 (N_16758,N_14117,N_14770);
xor U16759 (N_16759,N_12865,N_12919);
xnor U16760 (N_16760,N_14547,N_14277);
nor U16761 (N_16761,N_14637,N_13876);
nand U16762 (N_16762,N_13113,N_13087);
nand U16763 (N_16763,N_14190,N_14205);
nand U16764 (N_16764,N_14298,N_12768);
or U16765 (N_16765,N_13155,N_12864);
nor U16766 (N_16766,N_13683,N_13132);
nand U16767 (N_16767,N_13388,N_12509);
and U16768 (N_16768,N_13717,N_14741);
nand U16769 (N_16769,N_14316,N_13608);
nor U16770 (N_16770,N_12673,N_14666);
xnor U16771 (N_16771,N_12861,N_13458);
and U16772 (N_16772,N_13192,N_14052);
xnor U16773 (N_16773,N_13835,N_13823);
xor U16774 (N_16774,N_14304,N_12720);
nor U16775 (N_16775,N_13783,N_13062);
and U16776 (N_16776,N_14714,N_13719);
or U16777 (N_16777,N_13803,N_12950);
nand U16778 (N_16778,N_13550,N_13918);
nand U16779 (N_16779,N_14016,N_12599);
nor U16780 (N_16780,N_14092,N_12944);
and U16781 (N_16781,N_14704,N_12569);
nand U16782 (N_16782,N_14528,N_13271);
and U16783 (N_16783,N_13534,N_13389);
nor U16784 (N_16784,N_14934,N_13347);
or U16785 (N_16785,N_13308,N_14472);
or U16786 (N_16786,N_13754,N_13808);
and U16787 (N_16787,N_14644,N_12913);
xnor U16788 (N_16788,N_13175,N_12946);
and U16789 (N_16789,N_14966,N_14650);
nand U16790 (N_16790,N_14006,N_13038);
nor U16791 (N_16791,N_14744,N_14503);
nor U16792 (N_16792,N_14256,N_14558);
and U16793 (N_16793,N_13603,N_14286);
xor U16794 (N_16794,N_14510,N_12962);
and U16795 (N_16795,N_13217,N_14911);
xor U16796 (N_16796,N_12842,N_13387);
and U16797 (N_16797,N_12657,N_13612);
xnor U16798 (N_16798,N_13014,N_13042);
nand U16799 (N_16799,N_14202,N_14526);
or U16800 (N_16800,N_13555,N_14864);
or U16801 (N_16801,N_12854,N_13257);
and U16802 (N_16802,N_14242,N_14412);
nand U16803 (N_16803,N_12652,N_13822);
and U16804 (N_16804,N_13754,N_12885);
nor U16805 (N_16805,N_14707,N_14033);
nor U16806 (N_16806,N_13524,N_13045);
xor U16807 (N_16807,N_13648,N_14809);
nor U16808 (N_16808,N_14962,N_12726);
nor U16809 (N_16809,N_14486,N_14910);
xnor U16810 (N_16810,N_14331,N_12630);
or U16811 (N_16811,N_14073,N_13270);
nand U16812 (N_16812,N_13065,N_12760);
and U16813 (N_16813,N_14323,N_14458);
and U16814 (N_16814,N_13934,N_14282);
xor U16815 (N_16815,N_14456,N_14871);
or U16816 (N_16816,N_13279,N_14987);
nor U16817 (N_16817,N_13771,N_12608);
or U16818 (N_16818,N_13370,N_12979);
nand U16819 (N_16819,N_13719,N_14978);
nor U16820 (N_16820,N_14738,N_14950);
xor U16821 (N_16821,N_13408,N_14866);
and U16822 (N_16822,N_14692,N_13750);
and U16823 (N_16823,N_13780,N_14974);
nor U16824 (N_16824,N_14901,N_13505);
nor U16825 (N_16825,N_13807,N_13907);
xnor U16826 (N_16826,N_14471,N_14545);
xnor U16827 (N_16827,N_14788,N_13798);
or U16828 (N_16828,N_14552,N_13898);
nor U16829 (N_16829,N_14058,N_12536);
and U16830 (N_16830,N_14210,N_13413);
nor U16831 (N_16831,N_14366,N_14615);
nor U16832 (N_16832,N_12848,N_14581);
or U16833 (N_16833,N_13050,N_13651);
and U16834 (N_16834,N_13015,N_13638);
and U16835 (N_16835,N_12549,N_14018);
nand U16836 (N_16836,N_14541,N_13607);
nand U16837 (N_16837,N_14899,N_13865);
or U16838 (N_16838,N_14177,N_13286);
nand U16839 (N_16839,N_14588,N_14571);
and U16840 (N_16840,N_14489,N_13110);
nor U16841 (N_16841,N_12516,N_12535);
and U16842 (N_16842,N_14040,N_13386);
and U16843 (N_16843,N_12874,N_14559);
or U16844 (N_16844,N_14789,N_14818);
and U16845 (N_16845,N_14328,N_14573);
or U16846 (N_16846,N_12728,N_13423);
and U16847 (N_16847,N_13055,N_12594);
and U16848 (N_16848,N_14606,N_12524);
xnor U16849 (N_16849,N_14370,N_14421);
nor U16850 (N_16850,N_12646,N_12679);
and U16851 (N_16851,N_12504,N_14072);
xnor U16852 (N_16852,N_13369,N_13671);
or U16853 (N_16853,N_13122,N_14464);
and U16854 (N_16854,N_14811,N_14554);
or U16855 (N_16855,N_12811,N_14120);
xnor U16856 (N_16856,N_13513,N_12921);
xor U16857 (N_16857,N_14912,N_13049);
nor U16858 (N_16858,N_12983,N_14172);
xnor U16859 (N_16859,N_12615,N_12767);
nor U16860 (N_16860,N_13568,N_13865);
and U16861 (N_16861,N_12942,N_14169);
nor U16862 (N_16862,N_13422,N_13531);
nand U16863 (N_16863,N_12678,N_13794);
nor U16864 (N_16864,N_13513,N_13721);
xor U16865 (N_16865,N_12564,N_12744);
or U16866 (N_16866,N_14496,N_13930);
and U16867 (N_16867,N_14960,N_13714);
nor U16868 (N_16868,N_14994,N_12970);
and U16869 (N_16869,N_14258,N_13252);
xor U16870 (N_16870,N_12767,N_14494);
xor U16871 (N_16871,N_12833,N_14721);
nor U16872 (N_16872,N_12537,N_13848);
and U16873 (N_16873,N_12703,N_12937);
and U16874 (N_16874,N_14571,N_12759);
nand U16875 (N_16875,N_14368,N_13109);
nand U16876 (N_16876,N_12953,N_14644);
nor U16877 (N_16877,N_14502,N_14298);
xnor U16878 (N_16878,N_13859,N_12772);
nand U16879 (N_16879,N_13538,N_14210);
xnor U16880 (N_16880,N_13031,N_14183);
nand U16881 (N_16881,N_14080,N_12600);
nand U16882 (N_16882,N_12801,N_13195);
or U16883 (N_16883,N_14266,N_13604);
nand U16884 (N_16884,N_13020,N_14969);
xnor U16885 (N_16885,N_13777,N_14501);
or U16886 (N_16886,N_13334,N_14897);
nand U16887 (N_16887,N_14786,N_14267);
or U16888 (N_16888,N_12978,N_12993);
and U16889 (N_16889,N_14195,N_12824);
and U16890 (N_16890,N_13363,N_14427);
and U16891 (N_16891,N_14975,N_12582);
xnor U16892 (N_16892,N_12769,N_12723);
xor U16893 (N_16893,N_14143,N_13090);
xnor U16894 (N_16894,N_13741,N_14571);
and U16895 (N_16895,N_14253,N_13176);
nor U16896 (N_16896,N_14484,N_14203);
nand U16897 (N_16897,N_12562,N_14932);
nor U16898 (N_16898,N_13750,N_12594);
xnor U16899 (N_16899,N_14995,N_14461);
xor U16900 (N_16900,N_14899,N_13973);
and U16901 (N_16901,N_13649,N_13723);
and U16902 (N_16902,N_12874,N_13009);
xor U16903 (N_16903,N_12908,N_14312);
xor U16904 (N_16904,N_14925,N_12672);
or U16905 (N_16905,N_13899,N_13415);
xnor U16906 (N_16906,N_14053,N_14236);
xnor U16907 (N_16907,N_12728,N_14045);
and U16908 (N_16908,N_12914,N_13892);
xor U16909 (N_16909,N_14870,N_12600);
nor U16910 (N_16910,N_14175,N_12888);
xor U16911 (N_16911,N_13321,N_13346);
nand U16912 (N_16912,N_12616,N_14375);
or U16913 (N_16913,N_14497,N_14070);
and U16914 (N_16914,N_14903,N_14353);
nand U16915 (N_16915,N_12737,N_14617);
nor U16916 (N_16916,N_13610,N_13892);
nand U16917 (N_16917,N_13239,N_12877);
nand U16918 (N_16918,N_14402,N_13716);
or U16919 (N_16919,N_14878,N_13853);
and U16920 (N_16920,N_13005,N_12827);
nand U16921 (N_16921,N_13485,N_13079);
nand U16922 (N_16922,N_14576,N_14114);
xor U16923 (N_16923,N_12755,N_14804);
and U16924 (N_16924,N_13179,N_14492);
xor U16925 (N_16925,N_14758,N_12921);
nor U16926 (N_16926,N_13323,N_14887);
and U16927 (N_16927,N_13093,N_12703);
and U16928 (N_16928,N_14421,N_14653);
xnor U16929 (N_16929,N_13307,N_14076);
nor U16930 (N_16930,N_14386,N_13507);
nor U16931 (N_16931,N_14207,N_14905);
or U16932 (N_16932,N_14611,N_13708);
nor U16933 (N_16933,N_14374,N_12993);
and U16934 (N_16934,N_12834,N_12687);
nor U16935 (N_16935,N_12986,N_13660);
nand U16936 (N_16936,N_14718,N_13143);
xor U16937 (N_16937,N_13972,N_14012);
or U16938 (N_16938,N_14677,N_13020);
and U16939 (N_16939,N_14842,N_12970);
nor U16940 (N_16940,N_12616,N_13597);
xor U16941 (N_16941,N_14839,N_13870);
and U16942 (N_16942,N_12665,N_13477);
or U16943 (N_16943,N_13540,N_12857);
or U16944 (N_16944,N_14738,N_13366);
or U16945 (N_16945,N_13692,N_13303);
and U16946 (N_16946,N_13042,N_13961);
nand U16947 (N_16947,N_13896,N_12525);
nand U16948 (N_16948,N_13752,N_14690);
nand U16949 (N_16949,N_13590,N_13730);
xnor U16950 (N_16950,N_14545,N_14985);
xor U16951 (N_16951,N_14993,N_12736);
and U16952 (N_16952,N_14462,N_14600);
xnor U16953 (N_16953,N_14689,N_12569);
nand U16954 (N_16954,N_14136,N_13392);
nand U16955 (N_16955,N_14995,N_14257);
nand U16956 (N_16956,N_14510,N_13999);
xnor U16957 (N_16957,N_14343,N_13128);
nor U16958 (N_16958,N_13161,N_13430);
xnor U16959 (N_16959,N_13300,N_14407);
or U16960 (N_16960,N_14336,N_14381);
xor U16961 (N_16961,N_13224,N_12792);
xnor U16962 (N_16962,N_12862,N_14025);
or U16963 (N_16963,N_13332,N_13877);
xnor U16964 (N_16964,N_13833,N_12764);
or U16965 (N_16965,N_13238,N_12564);
xor U16966 (N_16966,N_12731,N_14307);
or U16967 (N_16967,N_14743,N_12918);
and U16968 (N_16968,N_12861,N_12696);
or U16969 (N_16969,N_12635,N_13157);
and U16970 (N_16970,N_14269,N_12825);
xor U16971 (N_16971,N_13946,N_13937);
xnor U16972 (N_16972,N_12611,N_13735);
nand U16973 (N_16973,N_13724,N_12837);
xnor U16974 (N_16974,N_12713,N_13305);
xnor U16975 (N_16975,N_14296,N_14952);
and U16976 (N_16976,N_13277,N_13127);
and U16977 (N_16977,N_14094,N_12788);
or U16978 (N_16978,N_14034,N_14371);
nand U16979 (N_16979,N_14772,N_13531);
or U16980 (N_16980,N_14918,N_14382);
or U16981 (N_16981,N_14217,N_13407);
nor U16982 (N_16982,N_13047,N_14826);
xor U16983 (N_16983,N_13579,N_13410);
or U16984 (N_16984,N_13297,N_13125);
nand U16985 (N_16985,N_14590,N_14827);
nand U16986 (N_16986,N_14051,N_13400);
or U16987 (N_16987,N_13620,N_14941);
nand U16988 (N_16988,N_13809,N_14503);
xnor U16989 (N_16989,N_13191,N_13774);
xnor U16990 (N_16990,N_14047,N_13321);
nor U16991 (N_16991,N_13296,N_12995);
xor U16992 (N_16992,N_12973,N_14663);
or U16993 (N_16993,N_13455,N_14350);
nand U16994 (N_16994,N_12949,N_14175);
nor U16995 (N_16995,N_13351,N_14520);
nand U16996 (N_16996,N_12969,N_14977);
nor U16997 (N_16997,N_14588,N_14774);
xor U16998 (N_16998,N_12833,N_13009);
nor U16999 (N_16999,N_13140,N_14982);
and U17000 (N_17000,N_14992,N_13439);
nor U17001 (N_17001,N_14823,N_13567);
or U17002 (N_17002,N_14605,N_13226);
nand U17003 (N_17003,N_14204,N_14599);
nand U17004 (N_17004,N_13844,N_14097);
or U17005 (N_17005,N_13105,N_14999);
xnor U17006 (N_17006,N_13436,N_12935);
or U17007 (N_17007,N_13489,N_14760);
nor U17008 (N_17008,N_13300,N_13651);
and U17009 (N_17009,N_14729,N_12608);
nor U17010 (N_17010,N_14507,N_13040);
nor U17011 (N_17011,N_12679,N_14889);
or U17012 (N_17012,N_13978,N_13599);
xnor U17013 (N_17013,N_12533,N_14285);
and U17014 (N_17014,N_14759,N_14624);
nand U17015 (N_17015,N_13613,N_14945);
nor U17016 (N_17016,N_14868,N_14286);
and U17017 (N_17017,N_12869,N_14027);
nor U17018 (N_17018,N_14399,N_14085);
or U17019 (N_17019,N_12614,N_14513);
or U17020 (N_17020,N_12923,N_13638);
or U17021 (N_17021,N_12942,N_13996);
xnor U17022 (N_17022,N_13982,N_14525);
nor U17023 (N_17023,N_14654,N_13572);
or U17024 (N_17024,N_13798,N_14289);
or U17025 (N_17025,N_14438,N_13284);
xnor U17026 (N_17026,N_14005,N_12597);
nand U17027 (N_17027,N_14271,N_13386);
nand U17028 (N_17028,N_14890,N_14880);
and U17029 (N_17029,N_13336,N_13493);
nor U17030 (N_17030,N_12970,N_14453);
and U17031 (N_17031,N_13876,N_12933);
and U17032 (N_17032,N_13858,N_13096);
nand U17033 (N_17033,N_12996,N_14258);
and U17034 (N_17034,N_14494,N_14937);
nor U17035 (N_17035,N_14971,N_13230);
and U17036 (N_17036,N_14513,N_12790);
xnor U17037 (N_17037,N_12707,N_12680);
or U17038 (N_17038,N_12853,N_14995);
and U17039 (N_17039,N_13793,N_13097);
xnor U17040 (N_17040,N_13630,N_13175);
nand U17041 (N_17041,N_13392,N_12525);
and U17042 (N_17042,N_13106,N_13262);
nor U17043 (N_17043,N_13455,N_14284);
xnor U17044 (N_17044,N_13421,N_14521);
or U17045 (N_17045,N_12764,N_12740);
xor U17046 (N_17046,N_13151,N_13535);
or U17047 (N_17047,N_14703,N_12868);
or U17048 (N_17048,N_12604,N_12526);
xor U17049 (N_17049,N_13106,N_14324);
and U17050 (N_17050,N_12671,N_13900);
nor U17051 (N_17051,N_13695,N_14942);
nor U17052 (N_17052,N_14571,N_13446);
xnor U17053 (N_17053,N_13370,N_13914);
and U17054 (N_17054,N_12683,N_12728);
xor U17055 (N_17055,N_13980,N_14063);
nor U17056 (N_17056,N_13478,N_12816);
or U17057 (N_17057,N_14218,N_13472);
or U17058 (N_17058,N_12918,N_13605);
nand U17059 (N_17059,N_13694,N_14727);
nor U17060 (N_17060,N_13125,N_12588);
and U17061 (N_17061,N_14688,N_14699);
nand U17062 (N_17062,N_13104,N_14307);
nor U17063 (N_17063,N_13542,N_13782);
or U17064 (N_17064,N_14054,N_13632);
and U17065 (N_17065,N_13521,N_13049);
nor U17066 (N_17066,N_14932,N_13901);
or U17067 (N_17067,N_13020,N_14360);
nor U17068 (N_17068,N_13186,N_13075);
nand U17069 (N_17069,N_14960,N_14779);
and U17070 (N_17070,N_13893,N_14591);
or U17071 (N_17071,N_12999,N_14435);
nor U17072 (N_17072,N_12575,N_12935);
and U17073 (N_17073,N_13416,N_14797);
xnor U17074 (N_17074,N_14681,N_13008);
or U17075 (N_17075,N_14838,N_12596);
and U17076 (N_17076,N_12864,N_14271);
xnor U17077 (N_17077,N_14611,N_13788);
nand U17078 (N_17078,N_14381,N_14091);
and U17079 (N_17079,N_13643,N_12835);
xor U17080 (N_17080,N_12713,N_13201);
xor U17081 (N_17081,N_13305,N_13182);
xor U17082 (N_17082,N_13773,N_14492);
nand U17083 (N_17083,N_13307,N_13024);
and U17084 (N_17084,N_12939,N_14264);
nor U17085 (N_17085,N_14788,N_14951);
xor U17086 (N_17086,N_13698,N_13807);
or U17087 (N_17087,N_14925,N_14044);
xor U17088 (N_17088,N_14904,N_13144);
nor U17089 (N_17089,N_12930,N_14884);
and U17090 (N_17090,N_14168,N_14568);
and U17091 (N_17091,N_13337,N_13811);
and U17092 (N_17092,N_13860,N_12900);
or U17093 (N_17093,N_13870,N_13738);
nor U17094 (N_17094,N_14991,N_14560);
nand U17095 (N_17095,N_13146,N_12663);
xor U17096 (N_17096,N_12835,N_13694);
xnor U17097 (N_17097,N_14340,N_12876);
nor U17098 (N_17098,N_13101,N_12698);
nor U17099 (N_17099,N_13326,N_14949);
or U17100 (N_17100,N_14044,N_14165);
and U17101 (N_17101,N_14287,N_13309);
nor U17102 (N_17102,N_13358,N_14089);
nand U17103 (N_17103,N_13191,N_14446);
nor U17104 (N_17104,N_13351,N_14779);
or U17105 (N_17105,N_14110,N_13586);
nand U17106 (N_17106,N_14011,N_14130);
or U17107 (N_17107,N_12508,N_13884);
nand U17108 (N_17108,N_13011,N_13211);
or U17109 (N_17109,N_13785,N_13199);
or U17110 (N_17110,N_13556,N_12904);
and U17111 (N_17111,N_14232,N_14021);
nor U17112 (N_17112,N_14070,N_12979);
nand U17113 (N_17113,N_14782,N_13353);
nand U17114 (N_17114,N_13329,N_13160);
nor U17115 (N_17115,N_13472,N_12681);
or U17116 (N_17116,N_13146,N_13035);
xnor U17117 (N_17117,N_13293,N_13678);
nand U17118 (N_17118,N_14046,N_12937);
xor U17119 (N_17119,N_14008,N_13196);
xor U17120 (N_17120,N_14320,N_13877);
nor U17121 (N_17121,N_13610,N_13367);
nand U17122 (N_17122,N_13291,N_14083);
nand U17123 (N_17123,N_13416,N_14331);
nor U17124 (N_17124,N_14378,N_12669);
nand U17125 (N_17125,N_14275,N_13991);
and U17126 (N_17126,N_13385,N_13611);
nand U17127 (N_17127,N_12884,N_12850);
or U17128 (N_17128,N_14180,N_14530);
nand U17129 (N_17129,N_12825,N_12635);
nor U17130 (N_17130,N_14685,N_13783);
and U17131 (N_17131,N_13564,N_13022);
xor U17132 (N_17132,N_12944,N_12714);
xor U17133 (N_17133,N_12805,N_14652);
xor U17134 (N_17134,N_12962,N_13096);
nor U17135 (N_17135,N_13570,N_13992);
or U17136 (N_17136,N_12783,N_12709);
or U17137 (N_17137,N_14817,N_14935);
nand U17138 (N_17138,N_13788,N_14136);
and U17139 (N_17139,N_14155,N_14704);
nor U17140 (N_17140,N_14403,N_12624);
xor U17141 (N_17141,N_13350,N_13284);
nor U17142 (N_17142,N_14409,N_13020);
xnor U17143 (N_17143,N_13135,N_12536);
or U17144 (N_17144,N_13801,N_13722);
or U17145 (N_17145,N_13758,N_13807);
or U17146 (N_17146,N_13868,N_13747);
and U17147 (N_17147,N_13956,N_14043);
nand U17148 (N_17148,N_14622,N_14787);
nand U17149 (N_17149,N_13781,N_14897);
or U17150 (N_17150,N_12829,N_13799);
and U17151 (N_17151,N_14639,N_13052);
or U17152 (N_17152,N_13190,N_13551);
xor U17153 (N_17153,N_13513,N_12552);
nand U17154 (N_17154,N_13829,N_14668);
xor U17155 (N_17155,N_14612,N_12994);
xor U17156 (N_17156,N_13205,N_12601);
nor U17157 (N_17157,N_14220,N_13404);
xor U17158 (N_17158,N_13640,N_13162);
or U17159 (N_17159,N_12530,N_14207);
nand U17160 (N_17160,N_14989,N_14352);
and U17161 (N_17161,N_13756,N_13522);
or U17162 (N_17162,N_14436,N_13048);
and U17163 (N_17163,N_13203,N_13409);
or U17164 (N_17164,N_13231,N_13788);
and U17165 (N_17165,N_12949,N_13990);
xor U17166 (N_17166,N_13164,N_12938);
or U17167 (N_17167,N_12834,N_14876);
and U17168 (N_17168,N_12799,N_13431);
nor U17169 (N_17169,N_14660,N_13040);
and U17170 (N_17170,N_14621,N_13626);
and U17171 (N_17171,N_12680,N_13147);
xnor U17172 (N_17172,N_13491,N_13455);
nor U17173 (N_17173,N_13061,N_12816);
or U17174 (N_17174,N_13840,N_13697);
and U17175 (N_17175,N_14909,N_13692);
nand U17176 (N_17176,N_12500,N_14461);
nor U17177 (N_17177,N_12897,N_13234);
nand U17178 (N_17178,N_13122,N_14012);
and U17179 (N_17179,N_12714,N_14227);
and U17180 (N_17180,N_13289,N_14963);
nand U17181 (N_17181,N_14089,N_14244);
or U17182 (N_17182,N_12841,N_13984);
and U17183 (N_17183,N_13394,N_12799);
nand U17184 (N_17184,N_14581,N_13020);
nor U17185 (N_17185,N_13195,N_13383);
or U17186 (N_17186,N_13765,N_13827);
nor U17187 (N_17187,N_14254,N_13181);
nand U17188 (N_17188,N_14030,N_13805);
nand U17189 (N_17189,N_13051,N_13081);
nor U17190 (N_17190,N_13960,N_12700);
or U17191 (N_17191,N_13349,N_12546);
nand U17192 (N_17192,N_14302,N_13823);
or U17193 (N_17193,N_13657,N_14252);
xor U17194 (N_17194,N_14418,N_14987);
nand U17195 (N_17195,N_14743,N_12572);
nand U17196 (N_17196,N_12941,N_13185);
nand U17197 (N_17197,N_13849,N_14717);
and U17198 (N_17198,N_12825,N_13411);
and U17199 (N_17199,N_13932,N_12605);
nor U17200 (N_17200,N_12692,N_14270);
and U17201 (N_17201,N_14391,N_14476);
and U17202 (N_17202,N_13381,N_14755);
nor U17203 (N_17203,N_12557,N_12731);
nand U17204 (N_17204,N_14440,N_13345);
xnor U17205 (N_17205,N_13397,N_13939);
and U17206 (N_17206,N_12610,N_14398);
or U17207 (N_17207,N_13309,N_12663);
nand U17208 (N_17208,N_14403,N_14922);
and U17209 (N_17209,N_13549,N_13468);
and U17210 (N_17210,N_13243,N_14544);
and U17211 (N_17211,N_14219,N_13425);
nor U17212 (N_17212,N_14062,N_14469);
xnor U17213 (N_17213,N_13649,N_12605);
nand U17214 (N_17214,N_14237,N_14941);
xor U17215 (N_17215,N_13749,N_14976);
or U17216 (N_17216,N_13519,N_14697);
nand U17217 (N_17217,N_14477,N_14755);
nor U17218 (N_17218,N_13028,N_14989);
xor U17219 (N_17219,N_14473,N_14426);
nor U17220 (N_17220,N_13206,N_12521);
or U17221 (N_17221,N_14782,N_14268);
nand U17222 (N_17222,N_13769,N_13944);
nand U17223 (N_17223,N_13516,N_14397);
nor U17224 (N_17224,N_13360,N_14179);
nand U17225 (N_17225,N_14727,N_14582);
or U17226 (N_17226,N_12658,N_13470);
nand U17227 (N_17227,N_14484,N_13749);
xor U17228 (N_17228,N_12858,N_13868);
or U17229 (N_17229,N_13582,N_12698);
xor U17230 (N_17230,N_13713,N_14919);
xor U17231 (N_17231,N_14673,N_13539);
or U17232 (N_17232,N_14275,N_13424);
nor U17233 (N_17233,N_14284,N_13078);
nand U17234 (N_17234,N_14635,N_14763);
nor U17235 (N_17235,N_13359,N_14112);
or U17236 (N_17236,N_13351,N_14214);
nand U17237 (N_17237,N_12682,N_12511);
nor U17238 (N_17238,N_13645,N_14518);
and U17239 (N_17239,N_13540,N_14506);
or U17240 (N_17240,N_13216,N_14451);
nor U17241 (N_17241,N_14977,N_12992);
nand U17242 (N_17242,N_14756,N_13862);
nor U17243 (N_17243,N_14897,N_13265);
nand U17244 (N_17244,N_13611,N_13233);
and U17245 (N_17245,N_12647,N_14821);
and U17246 (N_17246,N_14206,N_13835);
xnor U17247 (N_17247,N_13067,N_13182);
nand U17248 (N_17248,N_12756,N_13998);
or U17249 (N_17249,N_13573,N_13464);
nand U17250 (N_17250,N_13843,N_14969);
nand U17251 (N_17251,N_13806,N_13639);
nor U17252 (N_17252,N_13142,N_14368);
nor U17253 (N_17253,N_12793,N_12729);
xnor U17254 (N_17254,N_14400,N_13671);
or U17255 (N_17255,N_12643,N_13170);
xnor U17256 (N_17256,N_12500,N_13690);
nor U17257 (N_17257,N_14272,N_14960);
nor U17258 (N_17258,N_14251,N_13497);
nor U17259 (N_17259,N_13216,N_12673);
nand U17260 (N_17260,N_14869,N_12946);
and U17261 (N_17261,N_13221,N_13603);
or U17262 (N_17262,N_12704,N_12821);
nand U17263 (N_17263,N_13096,N_12958);
or U17264 (N_17264,N_14673,N_13368);
xnor U17265 (N_17265,N_12559,N_13276);
xnor U17266 (N_17266,N_13259,N_12506);
and U17267 (N_17267,N_14290,N_14125);
nor U17268 (N_17268,N_13875,N_14342);
nand U17269 (N_17269,N_13717,N_14291);
nor U17270 (N_17270,N_13845,N_13940);
nand U17271 (N_17271,N_12880,N_13892);
and U17272 (N_17272,N_12937,N_12825);
xnor U17273 (N_17273,N_14158,N_12819);
and U17274 (N_17274,N_12924,N_14772);
xnor U17275 (N_17275,N_12688,N_13838);
nor U17276 (N_17276,N_14931,N_12548);
nor U17277 (N_17277,N_13813,N_13963);
or U17278 (N_17278,N_13909,N_14516);
or U17279 (N_17279,N_13100,N_13304);
xor U17280 (N_17280,N_13009,N_14847);
or U17281 (N_17281,N_14614,N_13836);
xnor U17282 (N_17282,N_14803,N_13482);
or U17283 (N_17283,N_14714,N_14395);
nand U17284 (N_17284,N_14839,N_14064);
nand U17285 (N_17285,N_13298,N_14370);
xor U17286 (N_17286,N_14538,N_14048);
xnor U17287 (N_17287,N_12909,N_13465);
or U17288 (N_17288,N_12849,N_13138);
or U17289 (N_17289,N_14494,N_13427);
xnor U17290 (N_17290,N_13668,N_13919);
nand U17291 (N_17291,N_13131,N_14158);
or U17292 (N_17292,N_13864,N_12546);
nand U17293 (N_17293,N_12892,N_13662);
or U17294 (N_17294,N_13336,N_13828);
or U17295 (N_17295,N_12966,N_13984);
xor U17296 (N_17296,N_14717,N_13738);
or U17297 (N_17297,N_13295,N_13285);
xor U17298 (N_17298,N_14174,N_13875);
nor U17299 (N_17299,N_14489,N_14946);
nor U17300 (N_17300,N_12651,N_14469);
nand U17301 (N_17301,N_13451,N_12792);
nand U17302 (N_17302,N_14781,N_13096);
xor U17303 (N_17303,N_12802,N_14050);
nor U17304 (N_17304,N_13138,N_12816);
xor U17305 (N_17305,N_12554,N_13614);
xor U17306 (N_17306,N_12607,N_14961);
and U17307 (N_17307,N_14596,N_14327);
xnor U17308 (N_17308,N_13865,N_13637);
nor U17309 (N_17309,N_12942,N_13451);
nor U17310 (N_17310,N_14472,N_13809);
nor U17311 (N_17311,N_13809,N_13854);
nand U17312 (N_17312,N_14522,N_12772);
xor U17313 (N_17313,N_13798,N_14699);
and U17314 (N_17314,N_13452,N_14948);
nor U17315 (N_17315,N_13760,N_14118);
nand U17316 (N_17316,N_14386,N_14418);
nor U17317 (N_17317,N_12528,N_14642);
and U17318 (N_17318,N_13117,N_14417);
nor U17319 (N_17319,N_14029,N_12640);
nor U17320 (N_17320,N_14519,N_13293);
and U17321 (N_17321,N_14313,N_13125);
or U17322 (N_17322,N_13727,N_13237);
nor U17323 (N_17323,N_13993,N_13074);
nor U17324 (N_17324,N_12844,N_12557);
or U17325 (N_17325,N_14053,N_13991);
nor U17326 (N_17326,N_13829,N_12809);
and U17327 (N_17327,N_13905,N_13399);
or U17328 (N_17328,N_13346,N_14592);
and U17329 (N_17329,N_13524,N_13599);
or U17330 (N_17330,N_13416,N_12833);
and U17331 (N_17331,N_13991,N_12741);
or U17332 (N_17332,N_12956,N_13358);
or U17333 (N_17333,N_13590,N_12610);
or U17334 (N_17334,N_13704,N_13829);
nand U17335 (N_17335,N_13581,N_12691);
and U17336 (N_17336,N_14427,N_13583);
nor U17337 (N_17337,N_14960,N_14365);
xor U17338 (N_17338,N_12868,N_13366);
nand U17339 (N_17339,N_14356,N_14484);
nand U17340 (N_17340,N_14193,N_12502);
nand U17341 (N_17341,N_13676,N_14093);
and U17342 (N_17342,N_14760,N_14117);
and U17343 (N_17343,N_14509,N_14751);
or U17344 (N_17344,N_14934,N_14136);
or U17345 (N_17345,N_14032,N_14730);
xnor U17346 (N_17346,N_12763,N_13303);
xnor U17347 (N_17347,N_12949,N_14407);
and U17348 (N_17348,N_14739,N_13650);
xnor U17349 (N_17349,N_13208,N_14634);
nor U17350 (N_17350,N_13938,N_13151);
xnor U17351 (N_17351,N_13830,N_14653);
xnor U17352 (N_17352,N_13515,N_13933);
nand U17353 (N_17353,N_13001,N_14525);
nor U17354 (N_17354,N_13698,N_13902);
or U17355 (N_17355,N_14688,N_13443);
xor U17356 (N_17356,N_14736,N_12647);
nor U17357 (N_17357,N_13279,N_12814);
and U17358 (N_17358,N_14425,N_13497);
xnor U17359 (N_17359,N_13087,N_14511);
nand U17360 (N_17360,N_12837,N_13058);
nor U17361 (N_17361,N_13009,N_12920);
nand U17362 (N_17362,N_13606,N_14279);
nand U17363 (N_17363,N_13817,N_12827);
or U17364 (N_17364,N_14072,N_14117);
and U17365 (N_17365,N_13048,N_14952);
and U17366 (N_17366,N_13804,N_14805);
nor U17367 (N_17367,N_14402,N_13487);
xnor U17368 (N_17368,N_14884,N_13148);
xor U17369 (N_17369,N_13054,N_12654);
nand U17370 (N_17370,N_13925,N_12920);
nand U17371 (N_17371,N_12516,N_12538);
xnor U17372 (N_17372,N_14244,N_14722);
nor U17373 (N_17373,N_12827,N_13585);
xor U17374 (N_17374,N_12841,N_14337);
nor U17375 (N_17375,N_14834,N_12959);
or U17376 (N_17376,N_13961,N_14020);
xnor U17377 (N_17377,N_13923,N_14143);
xor U17378 (N_17378,N_14341,N_14851);
nand U17379 (N_17379,N_13222,N_14347);
xnor U17380 (N_17380,N_14994,N_14835);
nand U17381 (N_17381,N_13226,N_12656);
and U17382 (N_17382,N_14416,N_13069);
and U17383 (N_17383,N_14654,N_13731);
or U17384 (N_17384,N_12970,N_13688);
nand U17385 (N_17385,N_13720,N_14419);
nand U17386 (N_17386,N_14141,N_12754);
or U17387 (N_17387,N_13327,N_13789);
nand U17388 (N_17388,N_14105,N_14431);
nand U17389 (N_17389,N_12922,N_12766);
or U17390 (N_17390,N_14993,N_14884);
xnor U17391 (N_17391,N_14686,N_14626);
nor U17392 (N_17392,N_13689,N_13661);
and U17393 (N_17393,N_12608,N_12509);
nand U17394 (N_17394,N_12517,N_14992);
or U17395 (N_17395,N_14100,N_14913);
xor U17396 (N_17396,N_14599,N_14975);
and U17397 (N_17397,N_13411,N_13561);
xnor U17398 (N_17398,N_13503,N_13363);
and U17399 (N_17399,N_13295,N_13406);
or U17400 (N_17400,N_14981,N_14103);
nor U17401 (N_17401,N_12737,N_14183);
or U17402 (N_17402,N_14306,N_13988);
nor U17403 (N_17403,N_14906,N_13491);
nor U17404 (N_17404,N_12757,N_14931);
nand U17405 (N_17405,N_12768,N_14820);
or U17406 (N_17406,N_13985,N_14859);
nand U17407 (N_17407,N_13441,N_12946);
nand U17408 (N_17408,N_13440,N_14202);
nand U17409 (N_17409,N_13695,N_14939);
nor U17410 (N_17410,N_13027,N_13191);
nor U17411 (N_17411,N_13061,N_13471);
nor U17412 (N_17412,N_14335,N_14171);
and U17413 (N_17413,N_14764,N_14899);
or U17414 (N_17414,N_14380,N_13791);
nor U17415 (N_17415,N_13175,N_13300);
nand U17416 (N_17416,N_14951,N_14272);
nor U17417 (N_17417,N_14833,N_13137);
and U17418 (N_17418,N_12700,N_13001);
nand U17419 (N_17419,N_13419,N_13189);
nand U17420 (N_17420,N_13973,N_13925);
xor U17421 (N_17421,N_12870,N_12781);
or U17422 (N_17422,N_14328,N_14615);
or U17423 (N_17423,N_13510,N_13929);
nand U17424 (N_17424,N_12623,N_13136);
or U17425 (N_17425,N_12554,N_13369);
and U17426 (N_17426,N_14751,N_14813);
and U17427 (N_17427,N_14182,N_13957);
or U17428 (N_17428,N_12890,N_13891);
xnor U17429 (N_17429,N_13204,N_12814);
nor U17430 (N_17430,N_13479,N_13900);
xnor U17431 (N_17431,N_12566,N_12717);
nor U17432 (N_17432,N_12737,N_13006);
nor U17433 (N_17433,N_14631,N_13240);
xnor U17434 (N_17434,N_13367,N_13059);
nand U17435 (N_17435,N_13295,N_14331);
or U17436 (N_17436,N_13702,N_13880);
nor U17437 (N_17437,N_12623,N_13113);
nand U17438 (N_17438,N_12515,N_12986);
nor U17439 (N_17439,N_12550,N_13137);
nand U17440 (N_17440,N_13327,N_13874);
and U17441 (N_17441,N_13033,N_13818);
xnor U17442 (N_17442,N_12917,N_14823);
nor U17443 (N_17443,N_13524,N_13090);
or U17444 (N_17444,N_14669,N_13606);
nor U17445 (N_17445,N_14073,N_14292);
xnor U17446 (N_17446,N_14051,N_13041);
xor U17447 (N_17447,N_14366,N_12500);
xor U17448 (N_17448,N_13943,N_12659);
xor U17449 (N_17449,N_14202,N_13735);
nand U17450 (N_17450,N_13971,N_13594);
nand U17451 (N_17451,N_14493,N_12820);
nand U17452 (N_17452,N_14065,N_13403);
or U17453 (N_17453,N_12947,N_14911);
and U17454 (N_17454,N_14347,N_13863);
xnor U17455 (N_17455,N_13978,N_13355);
nor U17456 (N_17456,N_14698,N_14116);
nor U17457 (N_17457,N_13439,N_14232);
and U17458 (N_17458,N_12556,N_13683);
or U17459 (N_17459,N_14094,N_13483);
xnor U17460 (N_17460,N_13820,N_14674);
or U17461 (N_17461,N_14787,N_14408);
or U17462 (N_17462,N_14668,N_12639);
and U17463 (N_17463,N_12985,N_13725);
or U17464 (N_17464,N_14046,N_13470);
nand U17465 (N_17465,N_14082,N_14990);
nor U17466 (N_17466,N_14839,N_12861);
xnor U17467 (N_17467,N_13746,N_13911);
nor U17468 (N_17468,N_13196,N_14530);
nor U17469 (N_17469,N_13091,N_13055);
nor U17470 (N_17470,N_13567,N_14275);
nor U17471 (N_17471,N_13687,N_12716);
nor U17472 (N_17472,N_14186,N_13975);
and U17473 (N_17473,N_14136,N_14320);
or U17474 (N_17474,N_14344,N_13299);
nand U17475 (N_17475,N_12502,N_13511);
and U17476 (N_17476,N_12913,N_12894);
or U17477 (N_17477,N_14308,N_12524);
and U17478 (N_17478,N_14046,N_14127);
xnor U17479 (N_17479,N_13863,N_14497);
nor U17480 (N_17480,N_13658,N_13789);
xor U17481 (N_17481,N_14456,N_13979);
nor U17482 (N_17482,N_12549,N_14742);
xor U17483 (N_17483,N_12779,N_14861);
or U17484 (N_17484,N_13673,N_14160);
nor U17485 (N_17485,N_13015,N_12551);
nor U17486 (N_17486,N_13099,N_13281);
nor U17487 (N_17487,N_14133,N_13120);
and U17488 (N_17488,N_14674,N_12807);
nand U17489 (N_17489,N_14503,N_14920);
nand U17490 (N_17490,N_13121,N_12738);
nor U17491 (N_17491,N_14568,N_14648);
xor U17492 (N_17492,N_14403,N_12618);
or U17493 (N_17493,N_14575,N_12615);
or U17494 (N_17494,N_13512,N_14063);
nor U17495 (N_17495,N_12807,N_13624);
nand U17496 (N_17496,N_12866,N_13489);
xor U17497 (N_17497,N_14877,N_14888);
or U17498 (N_17498,N_13014,N_12615);
and U17499 (N_17499,N_13021,N_14281);
and U17500 (N_17500,N_15405,N_15429);
or U17501 (N_17501,N_15617,N_15391);
xnor U17502 (N_17502,N_16306,N_17265);
nor U17503 (N_17503,N_16979,N_17462);
and U17504 (N_17504,N_16585,N_15921);
nor U17505 (N_17505,N_17176,N_15265);
or U17506 (N_17506,N_17436,N_15852);
or U17507 (N_17507,N_15061,N_16770);
xnor U17508 (N_17508,N_16495,N_15817);
xnor U17509 (N_17509,N_16628,N_16052);
or U17510 (N_17510,N_16838,N_16635);
or U17511 (N_17511,N_16938,N_16487);
or U17512 (N_17512,N_17215,N_17303);
xnor U17513 (N_17513,N_17131,N_16912);
nor U17514 (N_17514,N_15945,N_16638);
and U17515 (N_17515,N_15428,N_15362);
xnor U17516 (N_17516,N_15084,N_17214);
nand U17517 (N_17517,N_16172,N_15583);
nand U17518 (N_17518,N_17494,N_15651);
and U17519 (N_17519,N_17413,N_15437);
and U17520 (N_17520,N_15769,N_17498);
nor U17521 (N_17521,N_16985,N_15110);
and U17522 (N_17522,N_15373,N_15984);
xor U17523 (N_17523,N_16233,N_15560);
nand U17524 (N_17524,N_16299,N_15038);
or U17525 (N_17525,N_16824,N_15126);
xor U17526 (N_17526,N_15460,N_16618);
xnor U17527 (N_17527,N_15714,N_16751);
nand U17528 (N_17528,N_17477,N_16232);
or U17529 (N_17529,N_16520,N_16948);
nand U17530 (N_17530,N_16396,N_15305);
xnor U17531 (N_17531,N_16900,N_15466);
nand U17532 (N_17532,N_16101,N_15514);
and U17533 (N_17533,N_17103,N_15462);
or U17534 (N_17534,N_16493,N_15726);
or U17535 (N_17535,N_16178,N_17314);
or U17536 (N_17536,N_16273,N_15117);
and U17537 (N_17537,N_17467,N_16524);
and U17538 (N_17538,N_15897,N_17197);
nand U17539 (N_17539,N_15159,N_17016);
nand U17540 (N_17540,N_17461,N_17340);
or U17541 (N_17541,N_15418,N_15006);
nand U17542 (N_17542,N_15664,N_17024);
and U17543 (N_17543,N_15350,N_17043);
nand U17544 (N_17544,N_16866,N_17470);
and U17545 (N_17545,N_15215,N_15051);
nand U17546 (N_17546,N_15426,N_15436);
or U17547 (N_17547,N_16566,N_16183);
xnor U17548 (N_17548,N_17159,N_16793);
nor U17549 (N_17549,N_15548,N_17006);
and U17550 (N_17550,N_15446,N_15231);
xnor U17551 (N_17551,N_17239,N_15316);
xnor U17552 (N_17552,N_16718,N_15195);
or U17553 (N_17553,N_15160,N_17089);
or U17554 (N_17554,N_15997,N_16880);
xor U17555 (N_17555,N_17489,N_17129);
xnor U17556 (N_17556,N_15237,N_16081);
xnor U17557 (N_17557,N_15191,N_15810);
nand U17558 (N_17558,N_15926,N_17000);
nand U17559 (N_17559,N_15590,N_15470);
and U17560 (N_17560,N_17308,N_15893);
nand U17561 (N_17561,N_15844,N_16499);
xnor U17562 (N_17562,N_16723,N_16312);
or U17563 (N_17563,N_15201,N_17408);
or U17564 (N_17564,N_15752,N_15993);
nor U17565 (N_17565,N_16182,N_17328);
nor U17566 (N_17566,N_16730,N_16486);
xnor U17567 (N_17567,N_15184,N_16674);
xnor U17568 (N_17568,N_15625,N_15613);
and U17569 (N_17569,N_16247,N_15511);
and U17570 (N_17570,N_16407,N_15455);
or U17571 (N_17571,N_17305,N_15032);
or U17572 (N_17572,N_17035,N_16847);
xnor U17573 (N_17573,N_15182,N_15659);
xor U17574 (N_17574,N_15318,N_15802);
xnor U17575 (N_17575,N_15230,N_17262);
xor U17576 (N_17576,N_17011,N_16672);
xnor U17577 (N_17577,N_16019,N_16889);
nor U17578 (N_17578,N_16909,N_15312);
and U17579 (N_17579,N_16675,N_16353);
xnor U17580 (N_17580,N_15414,N_15020);
nand U17581 (N_17581,N_16102,N_17237);
nor U17582 (N_17582,N_16141,N_17345);
and U17583 (N_17583,N_15857,N_16235);
or U17584 (N_17584,N_15435,N_15452);
and U17585 (N_17585,N_16630,N_15588);
xnor U17586 (N_17586,N_16278,N_16238);
nor U17587 (N_17587,N_17200,N_17032);
nand U17588 (N_17588,N_16657,N_15706);
xnor U17589 (N_17589,N_16735,N_15822);
or U17590 (N_17590,N_16901,N_17042);
nor U17591 (N_17591,N_16876,N_17376);
and U17592 (N_17592,N_15443,N_16171);
nor U17593 (N_17593,N_16083,N_16689);
and U17594 (N_17594,N_16927,N_15656);
nor U17595 (N_17595,N_16041,N_17435);
xor U17596 (N_17596,N_15695,N_15901);
nor U17597 (N_17597,N_15584,N_17329);
xnor U17598 (N_17598,N_16349,N_16040);
xor U17599 (N_17599,N_16255,N_16950);
nor U17600 (N_17600,N_15339,N_16414);
nor U17601 (N_17601,N_15207,N_17423);
and U17602 (N_17602,N_15448,N_16620);
nor U17603 (N_17603,N_15276,N_17317);
xnor U17604 (N_17604,N_17492,N_17458);
or U17605 (N_17605,N_16167,N_16127);
and U17606 (N_17606,N_16869,N_17058);
nand U17607 (N_17607,N_17065,N_16951);
or U17608 (N_17608,N_17087,N_16724);
nand U17609 (N_17609,N_17069,N_15570);
nand U17610 (N_17610,N_15727,N_17033);
nor U17611 (N_17611,N_15334,N_17247);
and U17612 (N_17612,N_16069,N_15853);
xnor U17613 (N_17613,N_16739,N_17294);
nand U17614 (N_17614,N_16429,N_17410);
or U17615 (N_17615,N_17420,N_16625);
xor U17616 (N_17616,N_16589,N_15874);
or U17617 (N_17617,N_15603,N_16882);
nand U17618 (N_17618,N_16545,N_15212);
and U17619 (N_17619,N_15325,N_15366);
nor U17620 (N_17620,N_15211,N_15925);
nor U17621 (N_17621,N_15115,N_16842);
and U17622 (N_17622,N_16116,N_16421);
nor U17623 (N_17623,N_16251,N_16667);
nand U17624 (N_17624,N_16700,N_16096);
and U17625 (N_17625,N_16305,N_15698);
and U17626 (N_17626,N_16248,N_15592);
nand U17627 (N_17627,N_15113,N_17459);
xor U17628 (N_17628,N_16276,N_15206);
nand U17629 (N_17629,N_17147,N_15492);
nand U17630 (N_17630,N_15392,N_16982);
nor U17631 (N_17631,N_15326,N_16764);
xnor U17632 (N_17632,N_15055,N_15454);
or U17633 (N_17633,N_15021,N_15292);
nor U17634 (N_17634,N_15861,N_16720);
nor U17635 (N_17635,N_15137,N_16448);
or U17636 (N_17636,N_16702,N_15682);
and U17637 (N_17637,N_16765,N_17037);
or U17638 (N_17638,N_16351,N_15124);
nor U17639 (N_17639,N_16343,N_15487);
nor U17640 (N_17640,N_15322,N_16144);
or U17641 (N_17641,N_16896,N_16510);
nand U17642 (N_17642,N_15968,N_17401);
xor U17643 (N_17643,N_15258,N_15840);
nand U17644 (N_17644,N_17402,N_16840);
nand U17645 (N_17645,N_15829,N_17444);
and U17646 (N_17646,N_15344,N_15071);
nor U17647 (N_17647,N_16825,N_17191);
and U17648 (N_17648,N_15858,N_15732);
nand U17649 (N_17649,N_17351,N_16898);
xor U17650 (N_17650,N_15547,N_16509);
nand U17651 (N_17651,N_17003,N_16086);
nor U17652 (N_17652,N_15631,N_16374);
nor U17653 (N_17653,N_17230,N_15027);
nor U17654 (N_17654,N_15776,N_15205);
nand U17655 (N_17655,N_15157,N_15639);
nor U17656 (N_17656,N_16789,N_16090);
and U17657 (N_17657,N_17210,N_16229);
nand U17658 (N_17658,N_15860,N_17448);
or U17659 (N_17659,N_16342,N_17479);
xnor U17660 (N_17660,N_15904,N_15304);
or U17661 (N_17661,N_16356,N_16669);
and U17662 (N_17662,N_15193,N_16465);
and U17663 (N_17663,N_15194,N_16892);
nor U17664 (N_17664,N_16389,N_16123);
or U17665 (N_17665,N_17460,N_15513);
and U17666 (N_17666,N_15715,N_16302);
nor U17667 (N_17667,N_16915,N_16234);
nor U17668 (N_17668,N_15379,N_16591);
and U17669 (N_17669,N_16957,N_15681);
and U17670 (N_17670,N_15210,N_15793);
and U17671 (N_17671,N_17365,N_16540);
nand U17672 (N_17672,N_15691,N_17219);
nor U17673 (N_17673,N_16942,N_16966);
or U17674 (N_17674,N_17140,N_16417);
xor U17675 (N_17675,N_16470,N_17051);
xor U17676 (N_17676,N_17300,N_16878);
and U17677 (N_17677,N_16451,N_16176);
xor U17678 (N_17678,N_16858,N_17185);
or U17679 (N_17679,N_17354,N_15250);
nand U17680 (N_17680,N_16188,N_15747);
or U17681 (N_17681,N_16446,N_15399);
nand U17682 (N_17682,N_17269,N_16679);
and U17683 (N_17683,N_16508,N_16968);
nor U17684 (N_17684,N_15125,N_15985);
xnor U17685 (N_17685,N_16798,N_15834);
xor U17686 (N_17686,N_17160,N_15891);
or U17687 (N_17687,N_16792,N_15828);
nor U17688 (N_17688,N_16129,N_15778);
xnor U17689 (N_17689,N_16627,N_16574);
xnor U17690 (N_17690,N_15256,N_17106);
or U17691 (N_17691,N_17403,N_16472);
and U17692 (N_17692,N_17199,N_15739);
xnor U17693 (N_17693,N_16920,N_15090);
and U17694 (N_17694,N_16242,N_15106);
nor U17695 (N_17695,N_16386,N_15842);
nor U17696 (N_17696,N_15238,N_15219);
and U17697 (N_17697,N_16652,N_16085);
xor U17698 (N_17698,N_17442,N_15257);
nand U17699 (N_17699,N_16523,N_15099);
nand U17700 (N_17700,N_17409,N_16130);
nand U17701 (N_17701,N_16485,N_17495);
nor U17702 (N_17702,N_16001,N_15552);
nor U17703 (N_17703,N_15242,N_17273);
xnor U17704 (N_17704,N_16296,N_15384);
nor U17705 (N_17705,N_16187,N_16425);
and U17706 (N_17706,N_17079,N_15712);
nor U17707 (N_17707,N_16837,N_16134);
nand U17708 (N_17708,N_16959,N_16411);
xnor U17709 (N_17709,N_16933,N_15886);
nand U17710 (N_17710,N_16157,N_15424);
or U17711 (N_17711,N_17184,N_17430);
xor U17712 (N_17712,N_16984,N_16831);
or U17713 (N_17713,N_17418,N_17235);
nand U17714 (N_17714,N_15836,N_16954);
xor U17715 (N_17715,N_16801,N_17233);
nor U17716 (N_17716,N_16681,N_16095);
xnor U17717 (N_17717,N_15505,N_15515);
or U17718 (N_17718,N_15410,N_15407);
nand U17719 (N_17719,N_17443,N_15542);
nand U17720 (N_17720,N_15493,N_15927);
nor U17721 (N_17721,N_17007,N_15811);
nor U17722 (N_17722,N_15598,N_15756);
xnor U17723 (N_17723,N_16070,N_15546);
xor U17724 (N_17724,N_17312,N_15266);
xor U17725 (N_17725,N_15202,N_15471);
nor U17726 (N_17726,N_16339,N_16026);
nand U17727 (N_17727,N_17204,N_16817);
nor U17728 (N_17728,N_16059,N_15672);
nand U17729 (N_17729,N_15315,N_15890);
xnor U17730 (N_17730,N_16094,N_15504);
and U17731 (N_17731,N_16453,N_16111);
nand U17732 (N_17732,N_17195,N_15233);
nor U17733 (N_17733,N_15724,N_15200);
xnor U17734 (N_17734,N_15610,N_15331);
xor U17735 (N_17735,N_15850,N_16197);
xor U17736 (N_17736,N_17277,N_15228);
and U17737 (N_17737,N_16303,N_17258);
nor U17738 (N_17738,N_16693,N_16500);
nor U17739 (N_17739,N_16972,N_17366);
xnor U17740 (N_17740,N_15516,N_15576);
nor U17741 (N_17741,N_16177,N_15889);
and U17742 (N_17742,N_16768,N_16164);
and U17743 (N_17743,N_15025,N_16314);
nor U17744 (N_17744,N_15544,N_16103);
xor U17745 (N_17745,N_15635,N_15794);
and U17746 (N_17746,N_17407,N_15742);
nor U17747 (N_17747,N_15088,N_15780);
and U17748 (N_17748,N_17092,N_15569);
nand U17749 (N_17749,N_16989,N_16553);
or U17750 (N_17750,N_15932,N_15924);
nor U17751 (N_17751,N_16281,N_16592);
nand U17752 (N_17752,N_17389,N_15571);
or U17753 (N_17753,N_17380,N_15019);
and U17754 (N_17754,N_16209,N_17446);
or U17755 (N_17755,N_15014,N_17055);
nor U17756 (N_17756,N_16051,N_15749);
nor U17757 (N_17757,N_17186,N_15039);
and U17758 (N_17758,N_15615,N_16511);
nand U17759 (N_17759,N_15243,N_15320);
and U17760 (N_17760,N_16269,N_15779);
or U17761 (N_17761,N_15523,N_16043);
and U17762 (N_17762,N_17093,N_16431);
nand U17763 (N_17763,N_15114,N_16267);
xor U17764 (N_17764,N_16551,N_16816);
and U17765 (N_17765,N_15646,N_17177);
or U17766 (N_17766,N_15575,N_16575);
nand U17767 (N_17767,N_16222,N_15653);
nor U17768 (N_17768,N_15758,N_15477);
or U17769 (N_17769,N_15234,N_16692);
or U17770 (N_17770,N_15181,N_15004);
nand U17771 (N_17771,N_15996,N_15536);
or U17772 (N_17772,N_15666,N_15813);
xor U17773 (N_17773,N_15060,N_15474);
and U17774 (N_17774,N_17068,N_15345);
or U17775 (N_17775,N_17468,N_15626);
or U17776 (N_17776,N_15442,N_16796);
xor U17777 (N_17777,N_15785,N_15669);
or U17778 (N_17778,N_15438,N_16594);
nand U17779 (N_17779,N_17124,N_16089);
and U17780 (N_17780,N_17449,N_15415);
nand U17781 (N_17781,N_15555,N_17137);
xnor U17782 (N_17782,N_16622,N_15746);
and U17783 (N_17783,N_15037,N_16297);
nand U17784 (N_17784,N_15464,N_15909);
xor U17785 (N_17785,N_16310,N_16328);
or U17786 (N_17786,N_15941,N_17179);
nor U17787 (N_17787,N_15644,N_16010);
or U17788 (N_17788,N_16120,N_15382);
nor U17789 (N_17789,N_15824,N_16512);
nor U17790 (N_17790,N_15713,N_15808);
or U17791 (N_17791,N_17346,N_16437);
and U17792 (N_17792,N_15358,N_15168);
nor U17793 (N_17793,N_15467,N_16680);
xor U17794 (N_17794,N_15658,N_15290);
nand U17795 (N_17795,N_16460,N_16136);
or U17796 (N_17796,N_15112,N_15629);
nor U17797 (N_17797,N_16691,N_15468);
nor U17798 (N_17798,N_15553,N_15872);
and U17799 (N_17799,N_16619,N_15971);
nand U17800 (N_17800,N_16639,N_16394);
and U17801 (N_17801,N_15688,N_15433);
nand U17802 (N_17802,N_15678,N_15273);
nor U17803 (N_17803,N_17450,N_16811);
or U17804 (N_17804,N_16150,N_15719);
nor U17805 (N_17805,N_16350,N_15223);
and U17806 (N_17806,N_15502,N_16686);
nor U17807 (N_17807,N_16533,N_15649);
or U17808 (N_17808,N_15476,N_16624);
xnor U17809 (N_17809,N_16109,N_17152);
nand U17810 (N_17810,N_16080,N_16936);
nor U17811 (N_17811,N_15611,N_17388);
xnor U17812 (N_17812,N_16827,N_15067);
or U17813 (N_17813,N_16941,N_17022);
nand U17814 (N_17814,N_16744,N_15692);
nor U17815 (N_17815,N_16206,N_16264);
nand U17816 (N_17816,N_15496,N_16370);
nor U17817 (N_17817,N_16364,N_16387);
and U17818 (N_17818,N_16148,N_15141);
or U17819 (N_17819,N_17132,N_15057);
nand U17820 (N_17820,N_16332,N_15915);
nor U17821 (N_17821,N_15917,N_16643);
nor U17822 (N_17822,N_17213,N_15143);
nor U17823 (N_17823,N_16623,N_16978);
xor U17824 (N_17824,N_16986,N_17339);
and U17825 (N_17825,N_15185,N_15637);
or U17826 (N_17826,N_15591,N_16252);
xnor U17827 (N_17827,N_16061,N_16721);
nand U17828 (N_17828,N_16929,N_15657);
and U17829 (N_17829,N_16087,N_16391);
xnor U17830 (N_17830,N_15532,N_15871);
or U17831 (N_17831,N_16039,N_16767);
nand U17832 (N_17832,N_16774,N_16772);
nand U17833 (N_17833,N_17284,N_17153);
and U17834 (N_17834,N_15260,N_15068);
and U17835 (N_17835,N_16308,N_15158);
xor U17836 (N_17836,N_15047,N_15307);
nand U17837 (N_17837,N_17382,N_16246);
xnor U17838 (N_17838,N_16947,N_15970);
nor U17839 (N_17839,N_15134,N_16382);
nor U17840 (N_17840,N_16658,N_16179);
and U17841 (N_17841,N_15285,N_15413);
xor U17842 (N_17842,N_16473,N_15512);
nand U17843 (N_17843,N_17078,N_15671);
or U17844 (N_17844,N_16044,N_15878);
nand U17845 (N_17845,N_16676,N_15680);
or U17846 (N_17846,N_15796,N_16218);
or U17847 (N_17847,N_16458,N_16018);
or U17848 (N_17848,N_16719,N_16397);
or U17849 (N_17849,N_16863,N_15267);
or U17850 (N_17850,N_17066,N_16993);
and U17851 (N_17851,N_16160,N_15192);
nor U17852 (N_17852,N_16185,N_16418);
nor U17853 (N_17853,N_16363,N_16703);
or U17854 (N_17854,N_16746,N_15275);
nand U17855 (N_17855,N_17421,N_17090);
nor U17856 (N_17856,N_16445,N_15109);
nor U17857 (N_17857,N_15558,N_17027);
or U17858 (N_17858,N_17263,N_16139);
and U17859 (N_17859,N_16734,N_15936);
xor U17860 (N_17860,N_16687,N_15495);
nand U17861 (N_17861,N_16262,N_16126);
nor U17862 (N_17862,N_17451,N_16226);
nor U17863 (N_17863,N_16047,N_16290);
and U17864 (N_17864,N_15648,N_17264);
or U17865 (N_17865,N_16385,N_16049);
nor U17866 (N_17866,N_16074,N_16527);
or U17867 (N_17867,N_17342,N_15819);
or U17868 (N_17868,N_16748,N_16257);
xor U17869 (N_17869,N_16315,N_15902);
and U17870 (N_17870,N_15684,N_16230);
xnor U17871 (N_17871,N_15076,N_15923);
and U17872 (N_17872,N_16549,N_17373);
or U17873 (N_17873,N_16991,N_15123);
or U17874 (N_17874,N_16464,N_15096);
nand U17875 (N_17875,N_17378,N_15518);
nand U17876 (N_17876,N_16336,N_17133);
nand U17877 (N_17877,N_16502,N_17161);
and U17878 (N_17878,N_15480,N_16728);
nand U17879 (N_17879,N_17381,N_15764);
and U17880 (N_17880,N_15083,N_15162);
or U17881 (N_17881,N_15792,N_16240);
or U17882 (N_17882,N_16921,N_17375);
xnor U17883 (N_17883,N_16999,N_17142);
or U17884 (N_17884,N_16964,N_16731);
xnor U17885 (N_17885,N_17225,N_16104);
nand U17886 (N_17886,N_16685,N_16565);
xor U17887 (N_17887,N_15204,N_15335);
nand U17888 (N_17888,N_16879,N_15333);
and U17889 (N_17889,N_15034,N_15948);
nor U17890 (N_17890,N_16195,N_15670);
nand U17891 (N_17891,N_15313,N_15577);
or U17892 (N_17892,N_17319,N_15255);
or U17893 (N_17893,N_16253,N_15760);
or U17894 (N_17894,N_16717,N_15735);
or U17895 (N_17895,N_16295,N_16958);
nor U17896 (N_17896,N_15655,N_17156);
nand U17897 (N_17897,N_17036,N_17119);
xor U17898 (N_17898,N_16987,N_16839);
and U17899 (N_17899,N_15284,N_17357);
nor U17900 (N_17900,N_15665,N_16355);
and U17901 (N_17901,N_17188,N_16268);
nor U17902 (N_17902,N_15221,N_17208);
and U17903 (N_17903,N_15865,N_16322);
and U17904 (N_17904,N_15489,N_17302);
or U17905 (N_17905,N_17292,N_16806);
nand U17906 (N_17906,N_16651,N_15832);
xnor U17907 (N_17907,N_17487,N_17044);
nor U17908 (N_17908,N_16304,N_16344);
or U17909 (N_17909,N_16482,N_15486);
and U17910 (N_17910,N_15906,N_16142);
xor U17911 (N_17911,N_16535,N_16563);
or U17912 (N_17912,N_15951,N_16057);
nor U17913 (N_17913,N_15403,N_17217);
or U17914 (N_17914,N_16128,N_17229);
and U17915 (N_17915,N_16406,N_16335);
and U17916 (N_17916,N_16404,N_15716);
nand U17917 (N_17917,N_16537,N_15703);
xor U17918 (N_17918,N_16440,N_17072);
nor U17919 (N_17919,N_17118,N_15314);
or U17920 (N_17920,N_16821,N_15485);
or U17921 (N_17921,N_15624,N_16568);
or U17922 (N_17922,N_17144,N_17018);
nand U17923 (N_17923,N_15013,N_16106);
xor U17924 (N_17924,N_16555,N_15950);
and U17925 (N_17925,N_16169,N_16376);
and U17926 (N_17926,N_15161,N_15643);
and U17927 (N_17927,N_17267,N_17395);
xor U17928 (N_17928,N_16983,N_16992);
nor U17929 (N_17929,N_16653,N_17041);
nand U17930 (N_17930,N_16097,N_17405);
or U17931 (N_17931,N_17431,N_15427);
nor U17932 (N_17932,N_15565,N_17295);
nand U17933 (N_17933,N_17231,N_17205);
nor U17934 (N_17934,N_16949,N_17253);
and U17935 (N_17935,N_17012,N_16547);
or U17936 (N_17936,N_16525,N_16832);
xor U17937 (N_17937,N_15245,N_15434);
nor U17938 (N_17938,N_16707,N_17100);
xor U17939 (N_17939,N_15774,N_16450);
and U17940 (N_17940,N_16249,N_15557);
nor U17941 (N_17941,N_17157,N_16347);
and U17942 (N_17942,N_15636,N_16601);
and U17943 (N_17943,N_16602,N_16153);
or U17944 (N_17944,N_15341,N_16334);
and U17945 (N_17945,N_16773,N_15676);
nand U17946 (N_17946,N_16053,N_15606);
nor U17947 (N_17947,N_15797,N_15801);
nand U17948 (N_17948,N_15864,N_15056);
nand U17949 (N_17949,N_16000,N_17399);
nand U17950 (N_17950,N_15701,N_15296);
and U17951 (N_17951,N_15826,N_15723);
or U17952 (N_17952,N_15431,N_16515);
nand U17953 (N_17953,N_17228,N_16497);
xor U17954 (N_17954,N_15073,N_17163);
or U17955 (N_17955,N_16256,N_15139);
nand U17956 (N_17956,N_15674,N_17464);
and U17957 (N_17957,N_16162,N_15298);
nand U17958 (N_17958,N_15116,N_16615);
nor U17959 (N_17959,N_16034,N_17173);
and U17960 (N_17960,N_16277,N_16196);
nand U17961 (N_17961,N_15481,N_16926);
xor U17962 (N_17962,N_16961,N_17138);
nor U17963 (N_17963,N_17488,N_15991);
and U17964 (N_17964,N_15609,N_16935);
and U17965 (N_17965,N_17146,N_16003);
or U17966 (N_17966,N_15738,N_16759);
xnor U17967 (N_17967,N_16704,N_17251);
xnor U17968 (N_17968,N_16813,N_16189);
and U17969 (N_17969,N_16517,N_16147);
nor U17970 (N_17970,N_15062,N_16902);
or U17971 (N_17971,N_16874,N_16705);
nand U17972 (N_17972,N_17048,N_15026);
or U17973 (N_17973,N_16002,N_16245);
nand U17974 (N_17974,N_16757,N_15277);
nor U17975 (N_17975,N_15521,N_16329);
nand U17976 (N_17976,N_15154,N_15987);
nand U17977 (N_17977,N_16763,N_16154);
or U17978 (N_17978,N_15937,N_16403);
xor U17979 (N_17979,N_15308,N_15705);
xor U17980 (N_17980,N_17491,N_15028);
nand U17981 (N_17981,N_15899,N_15227);
xnor U17982 (N_17982,N_16320,N_16513);
xnor U17983 (N_17983,N_15444,N_17088);
or U17984 (N_17984,N_15805,N_17271);
xor U17985 (N_17985,N_15843,N_15554);
nor U17986 (N_17986,N_17370,N_17166);
nor U17987 (N_17987,N_16844,N_15217);
nand U17988 (N_17988,N_16193,N_16932);
and U17989 (N_17989,N_15999,N_15001);
nor U17990 (N_17990,N_15710,N_15064);
nor U17991 (N_17991,N_17080,N_15751);
xnor U17992 (N_17992,N_15122,N_15599);
nor U17993 (N_17993,N_17178,N_16885);
xnor U17994 (N_17994,N_16841,N_17226);
and U17995 (N_17995,N_15053,N_16223);
nand U17996 (N_17996,N_16632,N_15709);
xor U17997 (N_17997,N_17322,N_15526);
nand U17998 (N_17998,N_17371,N_16780);
nor U17999 (N_17999,N_16014,N_15337);
nor U18000 (N_18000,N_16498,N_17394);
nor U18001 (N_18001,N_17260,N_16662);
xor U18002 (N_18002,N_16521,N_15142);
nor U18003 (N_18003,N_17256,N_15111);
nand U18004 (N_18004,N_16861,N_16970);
and U18005 (N_18005,N_16469,N_16969);
nor U18006 (N_18006,N_16413,N_15947);
xor U18007 (N_18007,N_16904,N_15809);
nor U18008 (N_18008,N_16456,N_15589);
xor U18009 (N_18009,N_15531,N_17279);
or U18010 (N_18010,N_16514,N_15903);
and U18011 (N_18011,N_17236,N_16997);
nand U18012 (N_18012,N_15965,N_16865);
xor U18013 (N_18013,N_15679,N_15015);
nand U18014 (N_18014,N_16576,N_16755);
or U18015 (N_18015,N_15069,N_17272);
and U18016 (N_18016,N_16597,N_17158);
nand U18017 (N_18017,N_16648,N_16800);
nor U18018 (N_18018,N_15767,N_17384);
nand U18019 (N_18019,N_16088,N_16205);
or U18020 (N_18020,N_16587,N_15994);
and U18021 (N_18021,N_15650,N_16042);
or U18022 (N_18022,N_16412,N_16626);
or U18023 (N_18023,N_16829,N_16113);
nor U18024 (N_18024,N_15880,N_15980);
xor U18025 (N_18025,N_15638,N_15788);
or U18026 (N_18026,N_16805,N_16378);
or U18027 (N_18027,N_17261,N_15484);
and U18028 (N_18028,N_15440,N_15740);
and U18029 (N_18029,N_16771,N_16531);
xnor U18030 (N_18030,N_16631,N_15128);
or U18031 (N_18031,N_15058,N_16833);
nand U18032 (N_18032,N_15827,N_15600);
and U18033 (N_18033,N_16608,N_17385);
nand U18034 (N_18034,N_16967,N_16005);
nor U18035 (N_18035,N_16732,N_15023);
nand U18036 (N_18036,N_16856,N_17296);
nor U18037 (N_18037,N_17454,N_15469);
and U18038 (N_18038,N_15416,N_17398);
nand U18039 (N_18039,N_16393,N_15866);
nor U18040 (N_18040,N_16855,N_16586);
and U18041 (N_18041,N_15841,N_16489);
xor U18042 (N_18042,N_17363,N_17324);
or U18043 (N_18043,N_15604,N_15354);
xor U18044 (N_18044,N_15849,N_17108);
nor U18045 (N_18045,N_16870,N_15317);
nor U18046 (N_18046,N_17490,N_16073);
or U18047 (N_18047,N_15929,N_16873);
nor U18048 (N_18048,N_15602,N_16518);
nor U18049 (N_18049,N_17134,N_16301);
xnor U18050 (N_18050,N_16490,N_17120);
nor U18051 (N_18051,N_16937,N_17143);
xor U18052 (N_18052,N_15800,N_15986);
or U18053 (N_18053,N_15961,N_16542);
and U18054 (N_18054,N_17220,N_16712);
or U18055 (N_18055,N_15582,N_16548);
and U18056 (N_18056,N_16809,N_15848);
nor U18057 (N_18057,N_16117,N_15208);
nor U18058 (N_18058,N_15170,N_15972);
xnor U18059 (N_18059,N_15506,N_17091);
and U18060 (N_18060,N_15197,N_16331);
and U18061 (N_18061,N_17139,N_17049);
and U18062 (N_18062,N_15640,N_15311);
nor U18063 (N_18063,N_16466,N_15080);
or U18064 (N_18064,N_15045,N_16250);
nand U18065 (N_18065,N_15867,N_16121);
nand U18066 (N_18066,N_15005,N_15831);
xnor U18067 (N_18067,N_16590,N_17001);
nand U18068 (N_18068,N_15838,N_15933);
or U18069 (N_18069,N_15072,N_15585);
xnor U18070 (N_18070,N_16782,N_15186);
xor U18071 (N_18071,N_17485,N_17334);
nor U18072 (N_18072,N_17417,N_15905);
nor U18073 (N_18073,N_16504,N_15895);
and U18074 (N_18074,N_15673,N_16522);
xor U18075 (N_18075,N_16236,N_16379);
nor U18076 (N_18076,N_16072,N_15456);
nor U18077 (N_18077,N_15699,N_16736);
nor U18078 (N_18078,N_17238,N_16955);
nand U18079 (N_18079,N_16893,N_15395);
xnor U18080 (N_18080,N_15174,N_15359);
nand U18081 (N_18081,N_17293,N_15851);
and U18082 (N_18082,N_16588,N_15995);
or U18083 (N_18083,N_17447,N_15882);
nand U18084 (N_18084,N_16559,N_15633);
and U18085 (N_18085,N_16606,N_17434);
nand U18086 (N_18086,N_16899,N_15291);
nor U18087 (N_18087,N_16327,N_16665);
or U18088 (N_18088,N_17023,N_16860);
xnor U18089 (N_18089,N_15420,N_16528);
and U18090 (N_18090,N_15616,N_17209);
nand U18091 (N_18091,N_15862,N_16836);
and U18092 (N_18092,N_17203,N_15783);
and U18093 (N_18093,N_15295,N_17175);
and U18094 (N_18094,N_17306,N_17466);
xor U18095 (N_18095,N_16914,N_16038);
xor U18096 (N_18096,N_16505,N_17171);
nand U18097 (N_18097,N_16420,N_16190);
and U18098 (N_18098,N_17170,N_15241);
nand U18099 (N_18099,N_17084,N_16371);
xor U18100 (N_18100,N_17481,N_16802);
or U18101 (N_18101,N_16380,N_17193);
or U18102 (N_18102,N_15095,N_16877);
or U18103 (N_18103,N_15900,N_15441);
nor U18104 (N_18104,N_17165,N_17113);
and U18105 (N_18105,N_15133,N_17073);
nor U18106 (N_18106,N_15940,N_15017);
xnor U18107 (N_18107,N_16220,N_17369);
nand U18108 (N_18108,N_17440,N_15654);
xor U18109 (N_18109,N_16062,N_15708);
xnor U18110 (N_18110,N_17327,N_17076);
nor U18111 (N_18111,N_15765,N_15240);
or U18112 (N_18112,N_16155,N_16733);
nand U18113 (N_18113,N_15118,N_16962);
xnor U18114 (N_18114,N_15928,N_17476);
and U18115 (N_18115,N_15030,N_16888);
or U18116 (N_18116,N_15002,N_16775);
or U18117 (N_18117,N_15302,N_15148);
and U18118 (N_18118,N_15772,N_15355);
nand U18119 (N_18119,N_16581,N_16677);
or U18120 (N_18120,N_17034,N_17309);
nand U18121 (N_18121,N_16633,N_17005);
xnor U18122 (N_18122,N_16384,N_16905);
and U18123 (N_18123,N_16781,N_15294);
or U18124 (N_18124,N_15562,N_15263);
and U18125 (N_18125,N_15007,N_16025);
xnor U18126 (N_18126,N_16434,N_15356);
nand U18127 (N_18127,N_15846,N_15696);
nand U18128 (N_18128,N_15031,N_15879);
xnor U18129 (N_18129,N_16670,N_15044);
or U18130 (N_18130,N_16060,N_16562);
or U18131 (N_18131,N_16359,N_16835);
and U18132 (N_18132,N_16028,N_17301);
and U18133 (N_18133,N_15310,N_16170);
nand U18134 (N_18134,N_17130,N_16207);
and U18135 (N_18135,N_16956,N_15264);
xnor U18136 (N_18136,N_16447,N_16145);
or U18137 (N_18137,N_16795,N_16480);
or U18138 (N_18138,N_16048,N_17116);
nor U18139 (N_18139,N_16820,N_16854);
nor U18140 (N_18140,N_15868,N_15898);
and U18141 (N_18141,N_16727,N_17297);
nor U18142 (N_18142,N_15482,N_16184);
nand U18143 (N_18143,N_16930,N_17248);
xor U18144 (N_18144,N_15040,N_16114);
nand U18145 (N_18145,N_17040,N_15188);
or U18146 (N_18146,N_15164,N_16595);
or U18147 (N_18147,N_17393,N_15102);
xor U18148 (N_18148,N_15942,N_15119);
nor U18149 (N_18149,N_16125,N_16713);
nand U18150 (N_18150,N_15324,N_16475);
or U18151 (N_18151,N_15402,N_15529);
nand U18152 (N_18152,N_15647,N_16641);
nand U18153 (N_18153,N_16138,N_15086);
and U18154 (N_18154,N_15966,N_16582);
nor U18155 (N_18155,N_16484,N_16851);
and U18156 (N_18156,N_15270,N_15894);
or U18157 (N_18157,N_17111,N_15097);
nand U18158 (N_18158,N_16872,N_17338);
nor U18159 (N_18159,N_15869,N_17315);
nor U18160 (N_18160,N_15149,N_16099);
nor U18161 (N_18161,N_16373,N_16289);
and U18162 (N_18162,N_16611,N_17141);
and U18163 (N_18163,N_16814,N_16390);
nand U18164 (N_18164,N_15417,N_15144);
nand U18165 (N_18165,N_15737,N_17455);
nand U18166 (N_18166,N_16375,N_15409);
nand U18167 (N_18167,N_15132,N_17274);
and U18168 (N_18168,N_15180,N_15579);
nand U18169 (N_18169,N_16092,N_17218);
and U18170 (N_18170,N_15107,N_16292);
and U18171 (N_18171,N_16023,N_16100);
xnor U18172 (N_18172,N_15042,N_15981);
or U18173 (N_18173,N_15763,N_15306);
xnor U18174 (N_18174,N_16180,N_16191);
nand U18175 (N_18175,N_15136,N_15203);
nand U18176 (N_18176,N_17198,N_16282);
xnor U18177 (N_18177,N_17017,N_17053);
nand U18178 (N_18178,N_15214,N_17059);
nor U18179 (N_18179,N_17275,N_15839);
xor U18180 (N_18180,N_16894,N_15820);
and U18181 (N_18181,N_17335,N_15368);
and U18182 (N_18182,N_16918,N_15235);
or U18183 (N_18183,N_17015,N_16076);
nor U18184 (N_18184,N_17187,N_16492);
or U18185 (N_18185,N_15010,N_16683);
or U18186 (N_18186,N_16293,N_15912);
and U18187 (N_18187,N_17333,N_16647);
nor U18188 (N_18188,N_16859,N_15008);
nand U18189 (N_18189,N_17360,N_15697);
nand U18190 (N_18190,N_15685,N_15108);
and U18191 (N_18191,N_16976,N_16006);
and U18192 (N_18192,N_16903,N_16640);
and U18193 (N_18193,N_16810,N_15074);
nor U18194 (N_18194,N_15367,N_17095);
nor U18195 (N_18195,N_15939,N_16055);
or U18196 (N_18196,N_16973,N_15394);
xor U18197 (N_18197,N_16365,N_15799);
nand U18198 (N_18198,N_15958,N_17484);
xor U18199 (N_18199,N_15973,N_16283);
and U18200 (N_18200,N_16165,N_17266);
and U18201 (N_18201,N_16455,N_15351);
xnor U18202 (N_18202,N_17452,N_15357);
nor U18203 (N_18203,N_15854,N_17350);
xor U18204 (N_18204,N_17270,N_15618);
and U18205 (N_18205,N_15525,N_15388);
xnor U18206 (N_18206,N_16036,N_17361);
nor U18207 (N_18207,N_15179,N_16093);
and U18208 (N_18208,N_15450,N_16922);
and U18209 (N_18209,N_15372,N_15533);
nand U18210 (N_18210,N_16311,N_16649);
nor U18211 (N_18211,N_16395,N_16785);
nor U18212 (N_18212,N_15381,N_17222);
and U18213 (N_18213,N_16210,N_15390);
nor U18214 (N_18214,N_15009,N_15375);
and U18215 (N_18215,N_15537,N_16593);
nand U18216 (N_18216,N_15596,N_15459);
or U18217 (N_18217,N_16091,N_16600);
and U18218 (N_18218,N_16368,N_17441);
or U18219 (N_18219,N_16298,N_15396);
nand U18220 (N_18220,N_17189,N_17362);
nor U18221 (N_18221,N_16199,N_16998);
xor U18222 (N_18222,N_16655,N_15750);
xnor U18223 (N_18223,N_15011,N_15540);
or U18224 (N_18224,N_15259,N_15363);
xnor U18225 (N_18225,N_16307,N_15608);
nand U18226 (N_18226,N_16266,N_15048);
and U18227 (N_18227,N_16318,N_15421);
and U18228 (N_18228,N_15627,N_16560);
nand U18229 (N_18229,N_17323,N_17259);
nand U18230 (N_18230,N_17474,N_15268);
or U18231 (N_18231,N_15172,N_15220);
nor U18232 (N_18232,N_16749,N_16786);
or U18233 (N_18233,N_15370,N_16064);
nor U18234 (N_18234,N_16607,N_16875);
nor U18235 (N_18235,N_15954,N_16452);
and U18236 (N_18236,N_17471,N_15667);
xor U18237 (N_18237,N_16803,N_17283);
nor U18238 (N_18238,N_15791,N_16629);
nand U18239 (N_18239,N_16925,N_16684);
nand U18240 (N_18240,N_15775,N_16584);
or U18241 (N_18241,N_15105,N_15248);
nor U18242 (N_18242,N_17321,N_17063);
xnor U18243 (N_18243,N_17221,N_17336);
nor U18244 (N_18244,N_15807,N_16642);
xnor U18245 (N_18245,N_15677,N_15377);
xnor U18246 (N_18246,N_15510,N_16690);
nand U18247 (N_18247,N_16225,N_15962);
nor U18248 (N_18248,N_15353,N_15524);
nor U18249 (N_18249,N_16324,N_15982);
or U18250 (N_18250,N_15527,N_16459);
and U18251 (N_18251,N_17422,N_17290);
or U18252 (N_18252,N_16503,N_16468);
nor U18253 (N_18253,N_16752,N_17353);
xnor U18254 (N_18254,N_16678,N_16695);
and U18255 (N_18255,N_16604,N_16202);
or U18256 (N_18256,N_15816,N_16995);
and U18257 (N_18257,N_15847,N_16402);
nand U18258 (N_18258,N_15408,N_15342);
nand U18259 (N_18259,N_15085,N_15156);
and U18260 (N_18260,N_17427,N_16037);
xnor U18261 (N_18261,N_16791,N_16501);
nand U18262 (N_18262,N_16068,N_16697);
nor U18263 (N_18263,N_15488,N_16573);
or U18264 (N_18264,N_16570,N_16952);
and U18265 (N_18265,N_17060,N_16291);
and U18266 (N_18266,N_17070,N_17453);
or U18267 (N_18267,N_16398,N_17250);
nand U18268 (N_18268,N_15559,N_16428);
and U18269 (N_18269,N_15120,N_15938);
nand U18270 (N_18270,N_16462,N_16423);
and U18271 (N_18271,N_15153,N_15328);
nor U18272 (N_18272,N_15722,N_15479);
or U18273 (N_18273,N_15041,N_16078);
or U18274 (N_18274,N_15759,N_17482);
nor U18275 (N_18275,N_15918,N_15361);
nor U18276 (N_18276,N_15593,N_15387);
xnor U18277 (N_18277,N_16476,N_16664);
and U18278 (N_18278,N_15877,N_15835);
nand U18279 (N_18279,N_16022,N_17010);
xnor U18280 (N_18280,N_16660,N_15823);
nor U18281 (N_18281,N_15404,N_15478);
and U18282 (N_18282,N_16325,N_15736);
xnor U18283 (N_18283,N_17437,N_16742);
nor U18284 (N_18284,N_17102,N_15165);
and U18285 (N_18285,N_15789,N_16722);
or U18286 (N_18286,N_16030,N_16654);
nand U18287 (N_18287,N_16797,N_15082);
nand U18288 (N_18288,N_17330,N_15702);
or U18289 (N_18289,N_15911,N_15497);
nand U18290 (N_18290,N_16330,N_15668);
or U18291 (N_18291,N_16323,N_17304);
nand U18292 (N_18292,N_16467,N_15449);
nor U18293 (N_18293,N_16988,N_16338);
or U18294 (N_18294,N_15630,N_17190);
xnor U18295 (N_18295,N_17276,N_15439);
or U18296 (N_18296,N_16016,N_17122);
nor U18297 (N_18297,N_15500,N_16449);
xor U18298 (N_18298,N_16158,N_17013);
nor U18299 (N_18299,N_15365,N_17245);
and U18300 (N_18300,N_17169,N_16745);
nor U18301 (N_18301,N_17383,N_15694);
xnor U18302 (N_18302,N_17117,N_16557);
and U18303 (N_18303,N_17288,N_15374);
nand U18304 (N_18304,N_15956,N_15930);
nor U18305 (N_18305,N_16477,N_16433);
xnor U18306 (N_18306,N_16945,N_16137);
nor U18307 (N_18307,N_15607,N_16284);
or U18308 (N_18308,N_16432,N_16804);
nor U18309 (N_18309,N_16636,N_16663);
xor U18310 (N_18310,N_15946,N_15121);
xnor U18311 (N_18311,N_16940,N_17182);
nor U18312 (N_18312,N_17234,N_17057);
nand U18313 (N_18313,N_16166,N_16131);
nand U18314 (N_18314,N_15196,N_17145);
or U18315 (N_18315,N_16392,N_15003);
nand U18316 (N_18316,N_15043,N_16911);
and U18317 (N_18317,N_15620,N_16819);
or U18318 (N_18318,N_16410,N_17252);
and U18319 (N_18319,N_16300,N_15229);
nand U18320 (N_18320,N_16761,N_17391);
or U18321 (N_18321,N_15884,N_17061);
and U18322 (N_18322,N_16424,N_15964);
xnor U18323 (N_18323,N_15327,N_17254);
nor U18324 (N_18324,N_15943,N_17240);
or U18325 (N_18325,N_17085,N_15472);
xnor U18326 (N_18326,N_16033,N_16066);
or U18327 (N_18327,N_16031,N_15271);
nand U18328 (N_18328,N_17356,N_16443);
or U18329 (N_18329,N_15171,N_15534);
or U18330 (N_18330,N_16071,N_16011);
xnor U18331 (N_18331,N_15189,N_16726);
nor U18332 (N_18332,N_15175,N_15978);
nor U18333 (N_18333,N_17404,N_16345);
xor U18334 (N_18334,N_17316,N_16481);
xor U18335 (N_18335,N_16494,N_15859);
and U18336 (N_18336,N_15837,N_15530);
nand U18337 (N_18337,N_15567,N_17298);
or U18338 (N_18338,N_17009,N_15745);
nand U18339 (N_18339,N_16203,N_17167);
nor U18340 (N_18340,N_15272,N_16556);
xor U18341 (N_18341,N_15499,N_17062);
xor U18342 (N_18342,N_17114,N_16341);
nor U18343 (N_18343,N_16754,N_16317);
or U18344 (N_18344,N_15281,N_15319);
and U18345 (N_18345,N_15689,N_16219);
nor U18346 (N_18346,N_16725,N_15718);
and U18347 (N_18347,N_16541,N_15873);
nor U18348 (N_18348,N_15130,N_17039);
nand U18349 (N_18349,N_16784,N_16706);
or U18350 (N_18350,N_16881,N_16644);
xor U18351 (N_18351,N_15049,N_15955);
nand U18352 (N_18352,N_15018,N_15422);
and U18353 (N_18353,N_17416,N_15795);
and U18354 (N_18354,N_17196,N_15297);
nand U18355 (N_18355,N_16286,N_15790);
or U18356 (N_18356,N_16572,N_15663);
nor U18357 (N_18357,N_15338,N_16173);
or U18358 (N_18358,N_15979,N_15908);
nand U18359 (N_18359,N_16561,N_16696);
nand U18360 (N_18360,N_16599,N_16035);
xor U18361 (N_18361,N_16079,N_15348);
or U18362 (N_18362,N_16974,N_17396);
nor U18363 (N_18363,N_17098,N_16007);
and U18364 (N_18364,N_15104,N_15528);
or U18365 (N_18365,N_16211,N_16483);
or U18366 (N_18366,N_15385,N_16288);
or U18367 (N_18367,N_16156,N_16361);
and U18368 (N_18368,N_15952,N_16146);
or U18369 (N_18369,N_16753,N_15881);
nand U18370 (N_18370,N_16471,N_15711);
nand U18371 (N_18371,N_16694,N_16354);
nor U18372 (N_18372,N_17101,N_16818);
and U18373 (N_18373,N_15458,N_16610);
nand U18374 (N_18374,N_16743,N_15743);
nor U18375 (N_18375,N_16923,N_15675);
xnor U18376 (N_18376,N_15825,N_15581);
or U18377 (N_18377,N_15717,N_17493);
or U18378 (N_18378,N_16309,N_15748);
and U18379 (N_18379,N_16671,N_16110);
xor U18380 (N_18380,N_17332,N_15568);
and U18381 (N_18381,N_16822,N_16826);
or U18382 (N_18382,N_15163,N_15914);
and U18383 (N_18383,N_16058,N_16758);
or U18384 (N_18384,N_16214,N_15239);
nand U18385 (N_18385,N_15587,N_15771);
nand U18386 (N_18386,N_15244,N_16263);
or U18387 (N_18387,N_15508,N_15700);
or U18388 (N_18388,N_16815,N_17211);
nand U18389 (N_18389,N_17285,N_15087);
nor U18390 (N_18390,N_17232,N_15731);
xor U18391 (N_18391,N_15509,N_16027);
and U18392 (N_18392,N_16848,N_15254);
and U18393 (N_18393,N_16279,N_17019);
or U18394 (N_18394,N_16917,N_16224);
nor U18395 (N_18395,N_16883,N_17473);
nor U18396 (N_18396,N_16163,N_16388);
nor U18397 (N_18397,N_15398,N_15803);
xor U18398 (N_18398,N_15236,N_16161);
xor U18399 (N_18399,N_16237,N_15815);
or U18400 (N_18400,N_16294,N_15463);
xnor U18401 (N_18401,N_16174,N_17439);
or U18402 (N_18402,N_16977,N_15693);
nor U18403 (N_18403,N_16666,N_16943);
nand U18404 (N_18404,N_15347,N_16788);
or U18405 (N_18405,N_16994,N_16944);
and U18406 (N_18406,N_16906,N_17415);
nor U18407 (N_18407,N_16701,N_15151);
nand U18408 (N_18408,N_15075,N_16488);
xnor U18409 (N_18409,N_16799,N_17168);
nor U18410 (N_18410,N_16215,N_16133);
or U18411 (N_18411,N_16032,N_17280);
and U18412 (N_18412,N_17419,N_17475);
nand U18413 (N_18413,N_15406,N_15580);
or U18414 (N_18414,N_16063,N_16009);
or U18415 (N_18415,N_16507,N_17326);
xnor U18416 (N_18416,N_16616,N_16422);
nor U18417 (N_18417,N_16864,N_16609);
and U18418 (N_18418,N_16769,N_16834);
xor U18419 (N_18419,N_15888,N_16122);
nand U18420 (N_18420,N_16119,N_15597);
xnor U18421 (N_18421,N_16200,N_15992);
nor U18422 (N_18422,N_16360,N_15960);
nand U18423 (N_18423,N_17224,N_16598);
nor U18424 (N_18424,N_16577,N_16435);
xor U18425 (N_18425,N_15491,N_15522);
or U18426 (N_18426,N_16454,N_15293);
nand U18427 (N_18427,N_15561,N_17465);
nand U18428 (N_18428,N_16274,N_15378);
or U18429 (N_18429,N_16550,N_15556);
nor U18430 (N_18430,N_16118,N_15863);
nor U18431 (N_18431,N_17151,N_16012);
or U18432 (N_18432,N_16852,N_15821);
and U18433 (N_18433,N_15289,N_15261);
or U18434 (N_18434,N_15262,N_15147);
nor U18435 (N_18435,N_17125,N_15475);
xor U18436 (N_18436,N_15094,N_15773);
nand U18437 (N_18437,N_16614,N_16020);
nand U18438 (N_18438,N_15786,N_16244);
nor U18439 (N_18439,N_15550,N_16316);
or U18440 (N_18440,N_16151,N_17480);
nand U18441 (N_18441,N_17377,N_17083);
nand U18442 (N_18442,N_16634,N_16673);
xnor U18443 (N_18443,N_15393,N_15551);
nor U18444 (N_18444,N_16939,N_16216);
and U18445 (N_18445,N_15252,N_15566);
nor U18446 (N_18446,N_16438,N_16149);
nor U18447 (N_18447,N_17094,N_17028);
and U18448 (N_18448,N_16213,N_16580);
nand U18449 (N_18449,N_16441,N_17425);
nand U18450 (N_18450,N_16897,N_15875);
nor U18451 (N_18451,N_16807,N_16479);
nand U18452 (N_18452,N_16461,N_15369);
and U18453 (N_18453,N_16546,N_17110);
or U18454 (N_18454,N_17064,N_16132);
and U18455 (N_18455,N_17463,N_16143);
and U18456 (N_18456,N_15451,N_16975);
nand U18457 (N_18457,N_15976,N_16583);
and U18458 (N_18458,N_16740,N_17379);
nor U18459 (N_18459,N_16221,N_17483);
nor U18460 (N_18460,N_17029,N_16212);
and U18461 (N_18461,N_16711,N_16098);
xnor U18462 (N_18462,N_16008,N_17020);
and U18463 (N_18463,N_15046,N_15628);
or U18464 (N_18464,N_16928,N_15279);
or U18465 (N_18465,N_15622,N_15349);
xnor U18466 (N_18466,N_17115,N_15150);
nor U18467 (N_18467,N_15412,N_16140);
nand U18468 (N_18468,N_16056,N_16275);
nand U18469 (N_18469,N_17496,N_15024);
nand U18470 (N_18470,N_15687,N_16168);
or U18471 (N_18471,N_15401,N_15352);
or U18472 (N_18472,N_17127,N_16208);
and U18473 (N_18473,N_15507,N_16787);
nor U18474 (N_18474,N_16346,N_15473);
nor U18475 (N_18475,N_16965,N_15360);
nand U18476 (N_18476,N_15761,N_16931);
nand U18477 (N_18477,N_17172,N_17355);
or U18478 (N_18478,N_17244,N_17246);
or U18479 (N_18479,N_15910,N_15101);
nor U18480 (N_18480,N_17359,N_16578);
or U18481 (N_18481,N_16013,N_16400);
nand U18482 (N_18482,N_16401,N_16077);
xnor U18483 (N_18483,N_16916,N_15078);
and U18484 (N_18484,N_15623,N_17112);
nor U18485 (N_18485,N_15050,N_17148);
xnor U18486 (N_18486,N_17438,N_16192);
nand U18487 (N_18487,N_15535,N_16175);
xor U18488 (N_18488,N_16613,N_16457);
or U18489 (N_18489,N_17255,N_15247);
or U18490 (N_18490,N_16075,N_16845);
xor U18491 (N_18491,N_16362,N_15818);
xnor U18492 (N_18492,N_15707,N_16741);
xor U18493 (N_18493,N_15806,N_17162);
and U18494 (N_18494,N_17386,N_16369);
nor U18495 (N_18495,N_17469,N_16710);
nand U18496 (N_18496,N_15321,N_16217);
and U18497 (N_18497,N_16688,N_16004);
nor U18498 (N_18498,N_15876,N_15586);
and U18499 (N_18499,N_16790,N_15812);
xor U18500 (N_18500,N_15246,N_16895);
xnor U18501 (N_18501,N_16427,N_15990);
xor U18502 (N_18502,N_17128,N_16405);
nand U18503 (N_18503,N_16564,N_16439);
nor U18504 (N_18504,N_16348,N_15892);
or U18505 (N_18505,N_17067,N_15187);
or U18506 (N_18506,N_17344,N_15103);
and U18507 (N_18507,N_16659,N_17406);
or U18508 (N_18508,N_15323,N_17286);
nor U18509 (N_18509,N_17047,N_16105);
nand U18510 (N_18510,N_16980,N_15066);
and U18511 (N_18511,N_15762,N_15766);
nand U18512 (N_18512,N_16934,N_17364);
xor U18513 (N_18513,N_15397,N_15453);
xnor U18514 (N_18514,N_15447,N_16029);
xor U18515 (N_18515,N_16054,N_16516);
and U18516 (N_18516,N_16709,N_17126);
nor U18517 (N_18517,N_15092,N_15957);
or U18518 (N_18518,N_17358,N_15782);
or U18519 (N_18519,N_16536,N_15364);
nor U18520 (N_18520,N_17347,N_15135);
and U18521 (N_18521,N_17086,N_16124);
nor U18522 (N_18522,N_16194,N_16021);
nand U18523 (N_18523,N_16871,N_16646);
xor U18524 (N_18524,N_17121,N_17282);
nand U18525 (N_18525,N_15690,N_16756);
xnor U18526 (N_18526,N_17105,N_16270);
nand U18527 (N_18527,N_15059,N_16538);
or U18528 (N_18528,N_15093,N_17216);
xor U18529 (N_18529,N_15016,N_15730);
and U18530 (N_18530,N_16645,N_17038);
nand U18531 (N_18531,N_16280,N_15178);
nor U18532 (N_18532,N_15376,N_15919);
and U18533 (N_18533,N_15621,N_16908);
nand U18534 (N_18534,N_16729,N_16239);
nand U18535 (N_18535,N_15140,N_16259);
nor U18536 (N_18536,N_16333,N_16924);
nor U18537 (N_18537,N_16271,N_17428);
xor U18538 (N_18538,N_16319,N_17002);
and U18539 (N_18539,N_15520,N_17374);
nor U18540 (N_18540,N_16907,N_17397);
nor U18541 (N_18541,N_15423,N_17291);
xor U18542 (N_18542,N_15983,N_15967);
nand U18543 (N_18543,N_15425,N_17432);
nand U18544 (N_18544,N_15216,N_15885);
or U18545 (N_18545,N_15077,N_15686);
xnor U18546 (N_18546,N_15605,N_17201);
xnor U18547 (N_18547,N_17325,N_17149);
and U18548 (N_18548,N_15798,N_16981);
nor U18549 (N_18549,N_16747,N_17313);
nor U18550 (N_18550,N_15035,N_17014);
nand U18551 (N_18551,N_15935,N_17241);
nor U18552 (N_18552,N_15169,N_15371);
nand U18553 (N_18553,N_17331,N_16884);
xor U18554 (N_18554,N_17054,N_17307);
nand U18555 (N_18555,N_15400,N_15232);
and U18556 (N_18556,N_15959,N_17206);
xnor U18557 (N_18557,N_15977,N_16946);
xnor U18558 (N_18558,N_16612,N_17123);
xor U18559 (N_18559,N_17107,N_15907);
or U18560 (N_18560,N_17183,N_16668);
nand U18561 (N_18561,N_16890,N_16015);
nor U18562 (N_18562,N_17456,N_17372);
or U18563 (N_18563,N_16372,N_17445);
nand U18564 (N_18564,N_16430,N_15249);
xor U18565 (N_18565,N_16971,N_16321);
nand U18566 (N_18566,N_15330,N_16603);
nor U18567 (N_18567,N_17278,N_15033);
nor U18568 (N_18568,N_15734,N_16357);
and U18569 (N_18569,N_15922,N_15494);
or U18570 (N_18570,N_15340,N_15855);
or U18571 (N_18571,N_16065,N_16808);
or U18572 (N_18572,N_15029,N_17457);
and U18573 (N_18573,N_15070,N_16963);
nand U18574 (N_18574,N_15222,N_15998);
or U18575 (N_18575,N_17368,N_15755);
or U18576 (N_18576,N_15517,N_17414);
nor U18577 (N_18577,N_15720,N_17497);
or U18578 (N_18578,N_16491,N_15601);
and U18579 (N_18579,N_15974,N_16868);
or U18580 (N_18580,N_15619,N_16135);
or U18581 (N_18581,N_17227,N_16415);
nand U18582 (N_18582,N_15595,N_16656);
xnor U18583 (N_18583,N_16830,N_16381);
nand U18584 (N_18584,N_15753,N_15000);
nor U18585 (N_18585,N_16714,N_15280);
and U18586 (N_18586,N_16285,N_15989);
or U18587 (N_18587,N_17242,N_15190);
nand U18588 (N_18588,N_15283,N_17310);
or U18589 (N_18589,N_16340,N_16779);
nor U18590 (N_18590,N_16539,N_16534);
nand U18591 (N_18591,N_15054,N_15641);
and U18592 (N_18592,N_16661,N_16474);
nand U18593 (N_18593,N_15089,N_15887);
or U18594 (N_18594,N_15642,N_15127);
and U18595 (N_18595,N_15419,N_15498);
and U18596 (N_18596,N_16426,N_15332);
nand U18597 (N_18597,N_17135,N_15411);
nand U18598 (N_18598,N_17164,N_15564);
nor U18599 (N_18599,N_17400,N_16867);
and U18600 (N_18600,N_15683,N_15614);
and U18601 (N_18601,N_16108,N_15660);
nand U18602 (N_18602,N_16496,N_15545);
xnor U18603 (N_18603,N_17387,N_16828);
nand U18604 (N_18604,N_17096,N_16107);
nor U18605 (N_18605,N_17026,N_15269);
xnor U18606 (N_18606,N_15022,N_16650);
nand U18607 (N_18607,N_17050,N_16254);
or U18608 (N_18608,N_15541,N_15777);
and U18609 (N_18609,N_15953,N_16258);
nor U18610 (N_18610,N_15274,N_15218);
or U18611 (N_18611,N_17008,N_15300);
or U18612 (N_18612,N_16352,N_17311);
nor U18613 (N_18613,N_16543,N_17154);
or U18614 (N_18614,N_16358,N_16919);
and U18615 (N_18615,N_16794,N_15091);
nor U18616 (N_18616,N_17202,N_17181);
and U18617 (N_18617,N_16778,N_15573);
xnor U18618 (N_18618,N_15634,N_15969);
nand U18619 (N_18619,N_15198,N_16409);
or U18620 (N_18620,N_17077,N_15152);
or U18621 (N_18621,N_15612,N_16084);
or U18622 (N_18622,N_15213,N_17411);
and U18623 (N_18623,N_17281,N_16699);
and U18624 (N_18624,N_16436,N_15733);
nand U18625 (N_18625,N_16596,N_16737);
and U18626 (N_18626,N_16846,N_15539);
nor U18627 (N_18627,N_16326,N_17341);
and U18628 (N_18628,N_16408,N_15975);
nand U18629 (N_18629,N_15870,N_17337);
or U18630 (N_18630,N_16272,N_15146);
xnor U18631 (N_18631,N_15225,N_15383);
or U18632 (N_18632,N_15100,N_17046);
and U18633 (N_18633,N_15949,N_16159);
nand U18634 (N_18634,N_15253,N_16617);
nand U18635 (N_18635,N_15944,N_15578);
nor U18636 (N_18636,N_16367,N_15503);
and U18637 (N_18637,N_17472,N_17150);
xnor U18638 (N_18638,N_15173,N_17174);
or U18639 (N_18639,N_15728,N_15065);
nand U18640 (N_18640,N_15288,N_16046);
nand U18641 (N_18641,N_17343,N_15704);
nor U18642 (N_18642,N_16530,N_17257);
and U18643 (N_18643,N_17348,N_17486);
xnor U18644 (N_18644,N_17136,N_16261);
nand U18645 (N_18645,N_16383,N_15224);
nand U18646 (N_18646,N_17352,N_17207);
nor U18647 (N_18647,N_17056,N_15052);
xor U18648 (N_18648,N_16024,N_15652);
xor U18649 (N_18649,N_15549,N_15770);
and U18650 (N_18650,N_15299,N_17025);
and U18651 (N_18651,N_17392,N_15916);
and U18652 (N_18652,N_16544,N_16843);
nor U18653 (N_18653,N_16529,N_16857);
nor U18654 (N_18654,N_17243,N_17299);
and U18655 (N_18655,N_17180,N_16783);
and U18656 (N_18656,N_15830,N_17004);
xnor U18657 (N_18657,N_16571,N_16198);
and U18658 (N_18658,N_15934,N_17030);
nand U18659 (N_18659,N_17071,N_17499);
or U18660 (N_18660,N_17075,N_15931);
and U18661 (N_18661,N_15177,N_17390);
nand U18662 (N_18662,N_15012,N_15432);
nand U18663 (N_18663,N_16243,N_16181);
nand U18664 (N_18664,N_16605,N_16766);
or U18665 (N_18665,N_17109,N_16777);
nand U18666 (N_18666,N_16738,N_15781);
and U18667 (N_18667,N_16853,N_16862);
xnor U18668 (N_18668,N_17052,N_15833);
or U18669 (N_18669,N_16891,N_15741);
and U18670 (N_18670,N_17249,N_16241);
nand U18671 (N_18671,N_16558,N_15336);
nand U18672 (N_18672,N_15166,N_16913);
and U18673 (N_18673,N_16050,N_16399);
and U18674 (N_18674,N_15572,N_17031);
xor U18675 (N_18675,N_16067,N_16569);
nor U18676 (N_18676,N_17320,N_15303);
nor U18677 (N_18677,N_15538,N_15784);
xor U18678 (N_18678,N_15519,N_17097);
or U18679 (N_18679,N_17426,N_16017);
and U18680 (N_18680,N_16716,N_15389);
or U18681 (N_18681,N_15063,N_17268);
nand U18682 (N_18682,N_16201,N_17192);
and U18683 (N_18683,N_16762,N_15145);
xor U18684 (N_18684,N_15036,N_17289);
xnor U18685 (N_18685,N_16442,N_15343);
xnor U18686 (N_18686,N_16526,N_15490);
and U18687 (N_18687,N_16579,N_17433);
and U18688 (N_18688,N_16313,N_15787);
xor U18689 (N_18689,N_15329,N_16478);
and U18690 (N_18690,N_15729,N_17074);
nor U18691 (N_18691,N_17412,N_16377);
or U18692 (N_18692,N_15098,N_16506);
and U18693 (N_18693,N_15430,N_16996);
nor U18694 (N_18694,N_15209,N_15963);
and U18695 (N_18695,N_16554,N_16760);
or U18696 (N_18696,N_16750,N_15883);
or U18697 (N_18697,N_15856,N_15804);
nor U18698 (N_18698,N_16204,N_16910);
nand U18699 (N_18699,N_15645,N_16228);
and U18700 (N_18700,N_17478,N_15725);
and U18701 (N_18701,N_16265,N_15845);
xnor U18702 (N_18702,N_16637,N_15386);
xnor U18703 (N_18703,N_16682,N_15131);
or U18704 (N_18704,N_15757,N_16186);
xnor U18705 (N_18705,N_16621,N_16886);
nor U18706 (N_18706,N_15988,N_17021);
nor U18707 (N_18707,N_15079,N_15662);
or U18708 (N_18708,N_16287,N_15594);
xnor U18709 (N_18709,N_15501,N_17082);
and U18710 (N_18710,N_16115,N_15754);
and U18711 (N_18711,N_16887,N_16519);
xor U18712 (N_18712,N_17424,N_15226);
nor U18713 (N_18713,N_16708,N_15563);
xor U18714 (N_18714,N_17318,N_15632);
and U18715 (N_18715,N_15483,N_15380);
xor U18716 (N_18716,N_17099,N_15457);
xnor U18717 (N_18717,N_16990,N_16231);
xnor U18718 (N_18718,N_16227,N_17212);
or U18719 (N_18719,N_15744,N_17429);
xnor U18720 (N_18720,N_15661,N_15278);
nand U18721 (N_18721,N_16419,N_15286);
xor U18722 (N_18722,N_16812,N_16715);
or U18723 (N_18723,N_15138,N_15081);
xnor U18724 (N_18724,N_15768,N_15155);
or U18725 (N_18725,N_16463,N_15129);
nand U18726 (N_18726,N_15574,N_17045);
nor U18727 (N_18727,N_17155,N_16045);
nor U18728 (N_18728,N_16552,N_15199);
and U18729 (N_18729,N_16953,N_16960);
nor U18730 (N_18730,N_15287,N_15913);
and U18731 (N_18731,N_15543,N_16112);
nand U18732 (N_18732,N_16337,N_15301);
nand U18733 (N_18733,N_16416,N_16444);
nand U18734 (N_18734,N_15282,N_15721);
or U18735 (N_18735,N_17287,N_17349);
xor U18736 (N_18736,N_15445,N_16152);
and U18737 (N_18737,N_16082,N_15309);
and U18738 (N_18738,N_16532,N_15346);
or U18739 (N_18739,N_15896,N_15251);
or U18740 (N_18740,N_16260,N_16776);
and U18741 (N_18741,N_15465,N_16366);
nand U18742 (N_18742,N_17194,N_15183);
xor U18743 (N_18743,N_17367,N_15814);
or U18744 (N_18744,N_17223,N_17104);
or U18745 (N_18745,N_17081,N_16850);
xor U18746 (N_18746,N_16698,N_15920);
and U18747 (N_18747,N_16849,N_15167);
nor U18748 (N_18748,N_15461,N_16567);
xor U18749 (N_18749,N_15176,N_16823);
or U18750 (N_18750,N_15009,N_16118);
and U18751 (N_18751,N_15429,N_15334);
nand U18752 (N_18752,N_17388,N_15237);
and U18753 (N_18753,N_15880,N_16215);
or U18754 (N_18754,N_16874,N_16217);
nand U18755 (N_18755,N_16434,N_15018);
nand U18756 (N_18756,N_15446,N_16653);
and U18757 (N_18757,N_16734,N_16230);
nor U18758 (N_18758,N_17161,N_15092);
and U18759 (N_18759,N_15316,N_17190);
or U18760 (N_18760,N_16678,N_17155);
and U18761 (N_18761,N_16581,N_15333);
nor U18762 (N_18762,N_15392,N_15402);
nand U18763 (N_18763,N_16151,N_16157);
nand U18764 (N_18764,N_15824,N_15713);
and U18765 (N_18765,N_16724,N_15639);
nand U18766 (N_18766,N_16608,N_15310);
nor U18767 (N_18767,N_17041,N_16582);
and U18768 (N_18768,N_16093,N_15646);
and U18769 (N_18769,N_15992,N_15460);
or U18770 (N_18770,N_16586,N_15342);
and U18771 (N_18771,N_15967,N_16396);
nor U18772 (N_18772,N_16543,N_17192);
or U18773 (N_18773,N_17280,N_16222);
nand U18774 (N_18774,N_16646,N_16111);
nand U18775 (N_18775,N_16836,N_17322);
xor U18776 (N_18776,N_16155,N_16222);
or U18777 (N_18777,N_15160,N_15597);
and U18778 (N_18778,N_15191,N_16176);
xor U18779 (N_18779,N_17290,N_15882);
xnor U18780 (N_18780,N_16516,N_15331);
nor U18781 (N_18781,N_15461,N_15552);
and U18782 (N_18782,N_17218,N_16395);
nor U18783 (N_18783,N_15929,N_15098);
and U18784 (N_18784,N_17022,N_15807);
or U18785 (N_18785,N_16127,N_15446);
or U18786 (N_18786,N_16724,N_15927);
nand U18787 (N_18787,N_15303,N_15819);
nor U18788 (N_18788,N_16453,N_16816);
nor U18789 (N_18789,N_15727,N_16308);
nand U18790 (N_18790,N_16159,N_16539);
or U18791 (N_18791,N_16130,N_15146);
nand U18792 (N_18792,N_17240,N_16541);
nor U18793 (N_18793,N_15089,N_16750);
nor U18794 (N_18794,N_15972,N_15696);
or U18795 (N_18795,N_15443,N_15067);
and U18796 (N_18796,N_16524,N_16886);
or U18797 (N_18797,N_16558,N_15282);
nand U18798 (N_18798,N_15725,N_15258);
and U18799 (N_18799,N_15172,N_16458);
and U18800 (N_18800,N_17049,N_17194);
or U18801 (N_18801,N_16154,N_15952);
and U18802 (N_18802,N_16762,N_16132);
nor U18803 (N_18803,N_16963,N_15377);
nor U18804 (N_18804,N_16184,N_16516);
or U18805 (N_18805,N_16389,N_16434);
nor U18806 (N_18806,N_15760,N_17139);
xnor U18807 (N_18807,N_15960,N_16664);
or U18808 (N_18808,N_16522,N_17061);
nand U18809 (N_18809,N_17296,N_15246);
xnor U18810 (N_18810,N_15187,N_16167);
or U18811 (N_18811,N_15205,N_15753);
or U18812 (N_18812,N_17048,N_16077);
nor U18813 (N_18813,N_15011,N_15968);
or U18814 (N_18814,N_15840,N_17304);
nand U18815 (N_18815,N_15722,N_15001);
xor U18816 (N_18816,N_16202,N_16990);
nand U18817 (N_18817,N_15776,N_17327);
xor U18818 (N_18818,N_15075,N_16707);
or U18819 (N_18819,N_17353,N_15605);
and U18820 (N_18820,N_15715,N_16760);
and U18821 (N_18821,N_16096,N_17015);
xnor U18822 (N_18822,N_15680,N_16508);
nand U18823 (N_18823,N_16990,N_17391);
or U18824 (N_18824,N_17446,N_15819);
nand U18825 (N_18825,N_16865,N_16179);
nor U18826 (N_18826,N_16600,N_15040);
or U18827 (N_18827,N_17283,N_16578);
and U18828 (N_18828,N_16590,N_15845);
nor U18829 (N_18829,N_16329,N_15419);
nor U18830 (N_18830,N_16441,N_16898);
xnor U18831 (N_18831,N_16969,N_16248);
nor U18832 (N_18832,N_16932,N_16862);
nor U18833 (N_18833,N_16695,N_15369);
and U18834 (N_18834,N_17326,N_17124);
and U18835 (N_18835,N_15980,N_15996);
nand U18836 (N_18836,N_16129,N_17125);
nand U18837 (N_18837,N_15290,N_17420);
and U18838 (N_18838,N_15993,N_15164);
and U18839 (N_18839,N_16130,N_17494);
nor U18840 (N_18840,N_15220,N_16060);
or U18841 (N_18841,N_15824,N_15002);
and U18842 (N_18842,N_17277,N_16442);
nand U18843 (N_18843,N_16963,N_16037);
nor U18844 (N_18844,N_17171,N_17306);
or U18845 (N_18845,N_15133,N_16251);
nand U18846 (N_18846,N_16049,N_16656);
nor U18847 (N_18847,N_16497,N_16487);
nor U18848 (N_18848,N_15492,N_16955);
nand U18849 (N_18849,N_15576,N_15482);
xor U18850 (N_18850,N_17282,N_15818);
or U18851 (N_18851,N_15785,N_16103);
xor U18852 (N_18852,N_15020,N_15198);
nor U18853 (N_18853,N_17233,N_15766);
or U18854 (N_18854,N_16330,N_17182);
nand U18855 (N_18855,N_16471,N_17493);
nand U18856 (N_18856,N_15301,N_15834);
nand U18857 (N_18857,N_16689,N_16137);
and U18858 (N_18858,N_15677,N_17354);
nand U18859 (N_18859,N_16717,N_16390);
nor U18860 (N_18860,N_16163,N_15074);
and U18861 (N_18861,N_15083,N_17152);
and U18862 (N_18862,N_15437,N_17469);
or U18863 (N_18863,N_15803,N_16634);
or U18864 (N_18864,N_15401,N_15486);
nand U18865 (N_18865,N_15440,N_15995);
nor U18866 (N_18866,N_15092,N_17188);
or U18867 (N_18867,N_17263,N_15152);
nand U18868 (N_18868,N_16207,N_15461);
or U18869 (N_18869,N_15173,N_16801);
nor U18870 (N_18870,N_15555,N_15064);
nand U18871 (N_18871,N_17175,N_16786);
nor U18872 (N_18872,N_16374,N_17309);
xnor U18873 (N_18873,N_15874,N_15918);
and U18874 (N_18874,N_15626,N_15016);
xnor U18875 (N_18875,N_17232,N_16789);
and U18876 (N_18876,N_16947,N_16231);
xnor U18877 (N_18877,N_17428,N_15586);
nand U18878 (N_18878,N_16593,N_17475);
nand U18879 (N_18879,N_16060,N_17113);
nand U18880 (N_18880,N_15724,N_16872);
xnor U18881 (N_18881,N_15927,N_17209);
nand U18882 (N_18882,N_16141,N_15262);
and U18883 (N_18883,N_16995,N_16911);
nand U18884 (N_18884,N_16556,N_16725);
xnor U18885 (N_18885,N_16224,N_16804);
nor U18886 (N_18886,N_16735,N_17154);
and U18887 (N_18887,N_16001,N_15002);
xnor U18888 (N_18888,N_15170,N_15025);
or U18889 (N_18889,N_15525,N_17273);
nand U18890 (N_18890,N_16475,N_15958);
nor U18891 (N_18891,N_15309,N_16394);
or U18892 (N_18892,N_16155,N_16482);
nor U18893 (N_18893,N_17106,N_16167);
nand U18894 (N_18894,N_15697,N_16887);
xor U18895 (N_18895,N_15066,N_17189);
nor U18896 (N_18896,N_16050,N_17400);
xnor U18897 (N_18897,N_15180,N_16121);
and U18898 (N_18898,N_16079,N_15037);
nand U18899 (N_18899,N_16095,N_15022);
nand U18900 (N_18900,N_16311,N_15255);
nand U18901 (N_18901,N_16092,N_16129);
xnor U18902 (N_18902,N_16641,N_15981);
and U18903 (N_18903,N_17316,N_17408);
and U18904 (N_18904,N_15621,N_17241);
nor U18905 (N_18905,N_16116,N_17114);
xor U18906 (N_18906,N_17293,N_16735);
or U18907 (N_18907,N_16655,N_16030);
nor U18908 (N_18908,N_16001,N_15724);
nand U18909 (N_18909,N_17316,N_16288);
or U18910 (N_18910,N_15683,N_15324);
xor U18911 (N_18911,N_15237,N_16487);
and U18912 (N_18912,N_15831,N_17071);
xnor U18913 (N_18913,N_16659,N_16617);
xor U18914 (N_18914,N_16047,N_15168);
or U18915 (N_18915,N_16750,N_15830);
xor U18916 (N_18916,N_15199,N_15164);
xnor U18917 (N_18917,N_17286,N_17100);
and U18918 (N_18918,N_15600,N_16699);
or U18919 (N_18919,N_17332,N_15200);
nor U18920 (N_18920,N_15348,N_15651);
xor U18921 (N_18921,N_16625,N_16093);
xnor U18922 (N_18922,N_17453,N_15175);
and U18923 (N_18923,N_16444,N_16196);
nor U18924 (N_18924,N_16674,N_16108);
or U18925 (N_18925,N_15429,N_16321);
or U18926 (N_18926,N_16784,N_17168);
or U18927 (N_18927,N_15990,N_15739);
nor U18928 (N_18928,N_15399,N_15001);
xnor U18929 (N_18929,N_16004,N_16234);
xnor U18930 (N_18930,N_15734,N_15253);
or U18931 (N_18931,N_16203,N_15496);
or U18932 (N_18932,N_16434,N_15833);
and U18933 (N_18933,N_15497,N_16487);
or U18934 (N_18934,N_17147,N_16285);
and U18935 (N_18935,N_15045,N_15370);
or U18936 (N_18936,N_15233,N_15221);
xor U18937 (N_18937,N_15750,N_16770);
or U18938 (N_18938,N_17013,N_16713);
nor U18939 (N_18939,N_17387,N_15431);
nor U18940 (N_18940,N_16166,N_16417);
xor U18941 (N_18941,N_17238,N_16077);
and U18942 (N_18942,N_15986,N_17075);
and U18943 (N_18943,N_15482,N_16330);
xnor U18944 (N_18944,N_17145,N_15372);
and U18945 (N_18945,N_16910,N_16807);
and U18946 (N_18946,N_16102,N_16699);
nand U18947 (N_18947,N_16809,N_15920);
nor U18948 (N_18948,N_16482,N_16078);
or U18949 (N_18949,N_16731,N_15386);
nand U18950 (N_18950,N_16263,N_16052);
nand U18951 (N_18951,N_15208,N_17208);
or U18952 (N_18952,N_16160,N_16528);
xor U18953 (N_18953,N_16812,N_17492);
xor U18954 (N_18954,N_15428,N_17185);
nor U18955 (N_18955,N_16322,N_15138);
and U18956 (N_18956,N_15440,N_16615);
xor U18957 (N_18957,N_17115,N_15669);
xnor U18958 (N_18958,N_15332,N_15966);
nor U18959 (N_18959,N_17116,N_17131);
nor U18960 (N_18960,N_16822,N_16322);
xnor U18961 (N_18961,N_16332,N_16590);
and U18962 (N_18962,N_16010,N_17312);
nor U18963 (N_18963,N_17179,N_16481);
nand U18964 (N_18964,N_15693,N_15804);
nor U18965 (N_18965,N_17293,N_17112);
or U18966 (N_18966,N_16669,N_17050);
nor U18967 (N_18967,N_15843,N_15739);
nand U18968 (N_18968,N_15869,N_15420);
xnor U18969 (N_18969,N_16715,N_15562);
xor U18970 (N_18970,N_15972,N_16949);
nand U18971 (N_18971,N_15336,N_15158);
xor U18972 (N_18972,N_15431,N_16219);
nand U18973 (N_18973,N_15845,N_16667);
xnor U18974 (N_18974,N_17305,N_16646);
xnor U18975 (N_18975,N_17294,N_15403);
and U18976 (N_18976,N_17439,N_17485);
xor U18977 (N_18977,N_15802,N_16502);
nor U18978 (N_18978,N_17357,N_15258);
xnor U18979 (N_18979,N_15559,N_15842);
nor U18980 (N_18980,N_16834,N_17499);
nor U18981 (N_18981,N_16750,N_16396);
xor U18982 (N_18982,N_15861,N_16201);
nand U18983 (N_18983,N_16319,N_15980);
or U18984 (N_18984,N_15576,N_15651);
nor U18985 (N_18985,N_17058,N_16761);
nor U18986 (N_18986,N_15953,N_15733);
or U18987 (N_18987,N_16246,N_15607);
or U18988 (N_18988,N_15301,N_15918);
xnor U18989 (N_18989,N_15078,N_15158);
xnor U18990 (N_18990,N_16164,N_15038);
nor U18991 (N_18991,N_16791,N_15649);
and U18992 (N_18992,N_15457,N_17281);
or U18993 (N_18993,N_16959,N_16974);
nor U18994 (N_18994,N_16094,N_15284);
or U18995 (N_18995,N_17260,N_17107);
nor U18996 (N_18996,N_15844,N_16360);
nand U18997 (N_18997,N_17241,N_17080);
nand U18998 (N_18998,N_16587,N_15708);
nand U18999 (N_18999,N_16444,N_15815);
and U19000 (N_19000,N_17302,N_16741);
and U19001 (N_19001,N_15376,N_17371);
and U19002 (N_19002,N_17330,N_16088);
or U19003 (N_19003,N_15456,N_17160);
or U19004 (N_19004,N_17151,N_17184);
xor U19005 (N_19005,N_15510,N_17188);
and U19006 (N_19006,N_15866,N_15276);
or U19007 (N_19007,N_16690,N_15320);
or U19008 (N_19008,N_16883,N_16631);
nor U19009 (N_19009,N_16098,N_15366);
or U19010 (N_19010,N_15036,N_16207);
nand U19011 (N_19011,N_16890,N_15794);
and U19012 (N_19012,N_15959,N_15337);
nand U19013 (N_19013,N_15702,N_15706);
and U19014 (N_19014,N_17256,N_16655);
or U19015 (N_19015,N_17263,N_15391);
nor U19016 (N_19016,N_16334,N_16663);
xor U19017 (N_19017,N_15719,N_17337);
nor U19018 (N_19018,N_17019,N_17347);
nor U19019 (N_19019,N_16532,N_16952);
or U19020 (N_19020,N_17163,N_17385);
nand U19021 (N_19021,N_16149,N_16537);
or U19022 (N_19022,N_15403,N_16197);
xor U19023 (N_19023,N_17315,N_15966);
or U19024 (N_19024,N_16035,N_16179);
and U19025 (N_19025,N_15005,N_16045);
and U19026 (N_19026,N_17420,N_16628);
and U19027 (N_19027,N_16770,N_15968);
and U19028 (N_19028,N_16248,N_16067);
nand U19029 (N_19029,N_15107,N_15266);
nand U19030 (N_19030,N_15561,N_15382);
nand U19031 (N_19031,N_16265,N_16526);
and U19032 (N_19032,N_15448,N_17345);
and U19033 (N_19033,N_17161,N_15069);
or U19034 (N_19034,N_15182,N_15082);
or U19035 (N_19035,N_16908,N_17107);
nand U19036 (N_19036,N_17141,N_17152);
or U19037 (N_19037,N_16157,N_17095);
or U19038 (N_19038,N_15777,N_17195);
nand U19039 (N_19039,N_16239,N_15093);
nor U19040 (N_19040,N_16333,N_17224);
and U19041 (N_19041,N_17341,N_15207);
nand U19042 (N_19042,N_16472,N_16248);
nand U19043 (N_19043,N_17253,N_15435);
xor U19044 (N_19044,N_15120,N_15926);
nor U19045 (N_19045,N_15149,N_17354);
nand U19046 (N_19046,N_15234,N_15820);
nor U19047 (N_19047,N_15561,N_16029);
and U19048 (N_19048,N_17269,N_17260);
and U19049 (N_19049,N_15840,N_16211);
nand U19050 (N_19050,N_16265,N_17016);
nand U19051 (N_19051,N_15034,N_16505);
and U19052 (N_19052,N_17472,N_15966);
nand U19053 (N_19053,N_17323,N_16573);
or U19054 (N_19054,N_16512,N_15003);
and U19055 (N_19055,N_16507,N_16627);
nand U19056 (N_19056,N_15421,N_15791);
xnor U19057 (N_19057,N_15227,N_15757);
or U19058 (N_19058,N_16946,N_17215);
nand U19059 (N_19059,N_16257,N_16253);
nor U19060 (N_19060,N_17110,N_17068);
nand U19061 (N_19061,N_16852,N_17018);
nand U19062 (N_19062,N_15880,N_16528);
and U19063 (N_19063,N_15946,N_16782);
nand U19064 (N_19064,N_15267,N_16543);
nor U19065 (N_19065,N_16514,N_16540);
or U19066 (N_19066,N_15094,N_15068);
or U19067 (N_19067,N_16743,N_16927);
or U19068 (N_19068,N_17458,N_17406);
nand U19069 (N_19069,N_15368,N_15806);
nor U19070 (N_19070,N_17261,N_16719);
or U19071 (N_19071,N_15617,N_15642);
or U19072 (N_19072,N_15489,N_15754);
nand U19073 (N_19073,N_15852,N_17384);
xnor U19074 (N_19074,N_17156,N_15012);
nor U19075 (N_19075,N_16878,N_17158);
nand U19076 (N_19076,N_17383,N_15715);
nand U19077 (N_19077,N_17282,N_17348);
xnor U19078 (N_19078,N_15029,N_16518);
nand U19079 (N_19079,N_15307,N_15682);
nor U19080 (N_19080,N_15591,N_15717);
nor U19081 (N_19081,N_15220,N_16547);
nor U19082 (N_19082,N_15246,N_16962);
nand U19083 (N_19083,N_17218,N_15696);
nor U19084 (N_19084,N_17337,N_17024);
and U19085 (N_19085,N_16368,N_15447);
nand U19086 (N_19086,N_16686,N_15501);
and U19087 (N_19087,N_16476,N_15135);
nor U19088 (N_19088,N_16153,N_15979);
xor U19089 (N_19089,N_15498,N_17404);
or U19090 (N_19090,N_15042,N_15945);
xor U19091 (N_19091,N_15783,N_16770);
nor U19092 (N_19092,N_15257,N_15810);
or U19093 (N_19093,N_17301,N_17268);
nor U19094 (N_19094,N_16110,N_15022);
nand U19095 (N_19095,N_15370,N_15586);
and U19096 (N_19096,N_16894,N_17134);
xor U19097 (N_19097,N_15291,N_16010);
or U19098 (N_19098,N_16850,N_16186);
xor U19099 (N_19099,N_15313,N_16515);
nor U19100 (N_19100,N_15126,N_15063);
or U19101 (N_19101,N_17049,N_17281);
or U19102 (N_19102,N_16942,N_15629);
nor U19103 (N_19103,N_17423,N_16828);
nand U19104 (N_19104,N_16000,N_15184);
or U19105 (N_19105,N_16750,N_16156);
xnor U19106 (N_19106,N_15760,N_16953);
or U19107 (N_19107,N_16998,N_16938);
and U19108 (N_19108,N_16466,N_15946);
and U19109 (N_19109,N_15300,N_15836);
nand U19110 (N_19110,N_15725,N_15582);
xnor U19111 (N_19111,N_15637,N_15028);
nand U19112 (N_19112,N_17107,N_15710);
or U19113 (N_19113,N_16212,N_15813);
xor U19114 (N_19114,N_15549,N_16562);
xnor U19115 (N_19115,N_16073,N_16696);
nor U19116 (N_19116,N_15290,N_16181);
nand U19117 (N_19117,N_15954,N_16830);
and U19118 (N_19118,N_17170,N_16680);
nand U19119 (N_19119,N_16346,N_16524);
nand U19120 (N_19120,N_16442,N_17370);
nor U19121 (N_19121,N_17424,N_16869);
and U19122 (N_19122,N_15966,N_15916);
nand U19123 (N_19123,N_17051,N_16343);
xnor U19124 (N_19124,N_15943,N_16276);
xor U19125 (N_19125,N_15794,N_15983);
and U19126 (N_19126,N_15512,N_15597);
or U19127 (N_19127,N_16841,N_16090);
or U19128 (N_19128,N_17109,N_16627);
nor U19129 (N_19129,N_15558,N_15093);
nor U19130 (N_19130,N_15816,N_16630);
nand U19131 (N_19131,N_15272,N_16202);
nor U19132 (N_19132,N_17172,N_16913);
nor U19133 (N_19133,N_16615,N_16864);
and U19134 (N_19134,N_16374,N_15079);
nor U19135 (N_19135,N_15503,N_17297);
xnor U19136 (N_19136,N_15229,N_16419);
and U19137 (N_19137,N_16901,N_16306);
nor U19138 (N_19138,N_17154,N_15108);
nor U19139 (N_19139,N_16373,N_15147);
nor U19140 (N_19140,N_16325,N_15363);
xnor U19141 (N_19141,N_17153,N_15082);
nand U19142 (N_19142,N_15506,N_17078);
nand U19143 (N_19143,N_15742,N_16327);
nand U19144 (N_19144,N_15865,N_16301);
nand U19145 (N_19145,N_17337,N_16492);
nor U19146 (N_19146,N_17379,N_16540);
or U19147 (N_19147,N_16166,N_16737);
nor U19148 (N_19148,N_15959,N_15339);
nand U19149 (N_19149,N_15561,N_16293);
or U19150 (N_19150,N_16798,N_16933);
or U19151 (N_19151,N_15114,N_17477);
nor U19152 (N_19152,N_17428,N_15310);
xnor U19153 (N_19153,N_16533,N_17456);
and U19154 (N_19154,N_16755,N_15329);
and U19155 (N_19155,N_15918,N_16524);
and U19156 (N_19156,N_15772,N_16634);
or U19157 (N_19157,N_16885,N_15468);
or U19158 (N_19158,N_16132,N_17479);
nor U19159 (N_19159,N_15081,N_15801);
nor U19160 (N_19160,N_16392,N_15499);
nand U19161 (N_19161,N_16852,N_15527);
and U19162 (N_19162,N_16162,N_16722);
or U19163 (N_19163,N_15239,N_17470);
and U19164 (N_19164,N_17053,N_17448);
and U19165 (N_19165,N_15177,N_16255);
or U19166 (N_19166,N_15434,N_16571);
and U19167 (N_19167,N_15707,N_16509);
nor U19168 (N_19168,N_15527,N_17243);
nand U19169 (N_19169,N_17482,N_15272);
nor U19170 (N_19170,N_16282,N_16475);
and U19171 (N_19171,N_15940,N_16243);
nand U19172 (N_19172,N_15069,N_16443);
nand U19173 (N_19173,N_16746,N_16503);
nand U19174 (N_19174,N_15034,N_16291);
or U19175 (N_19175,N_15719,N_17233);
nor U19176 (N_19176,N_16018,N_17359);
and U19177 (N_19177,N_15290,N_15089);
and U19178 (N_19178,N_15219,N_15234);
and U19179 (N_19179,N_15964,N_16184);
nand U19180 (N_19180,N_16755,N_15652);
and U19181 (N_19181,N_15840,N_16831);
nor U19182 (N_19182,N_16721,N_16904);
and U19183 (N_19183,N_16536,N_16113);
nor U19184 (N_19184,N_15579,N_17177);
and U19185 (N_19185,N_15326,N_15143);
nand U19186 (N_19186,N_16714,N_16839);
and U19187 (N_19187,N_16792,N_16140);
nor U19188 (N_19188,N_16436,N_16389);
or U19189 (N_19189,N_17045,N_16606);
or U19190 (N_19190,N_15588,N_16545);
xor U19191 (N_19191,N_17232,N_16116);
and U19192 (N_19192,N_17116,N_16862);
nand U19193 (N_19193,N_15864,N_17202);
nor U19194 (N_19194,N_17413,N_16354);
and U19195 (N_19195,N_16335,N_16097);
or U19196 (N_19196,N_15882,N_16813);
xnor U19197 (N_19197,N_15129,N_15694);
xor U19198 (N_19198,N_16442,N_15171);
nor U19199 (N_19199,N_15857,N_16545);
xor U19200 (N_19200,N_17141,N_15695);
or U19201 (N_19201,N_15881,N_17269);
and U19202 (N_19202,N_15724,N_15299);
and U19203 (N_19203,N_16296,N_17389);
xnor U19204 (N_19204,N_15873,N_17091);
nor U19205 (N_19205,N_15828,N_15532);
nor U19206 (N_19206,N_15800,N_16981);
or U19207 (N_19207,N_15716,N_16896);
nand U19208 (N_19208,N_16198,N_15255);
or U19209 (N_19209,N_16010,N_15562);
xor U19210 (N_19210,N_16454,N_17339);
nand U19211 (N_19211,N_17438,N_15362);
and U19212 (N_19212,N_15463,N_17300);
nor U19213 (N_19213,N_16561,N_16436);
and U19214 (N_19214,N_17263,N_16082);
nand U19215 (N_19215,N_16461,N_15340);
and U19216 (N_19216,N_16024,N_16972);
or U19217 (N_19217,N_16204,N_16814);
nand U19218 (N_19218,N_15038,N_16217);
nand U19219 (N_19219,N_15137,N_15477);
nand U19220 (N_19220,N_16916,N_15578);
and U19221 (N_19221,N_16865,N_15783);
or U19222 (N_19222,N_16776,N_15844);
nor U19223 (N_19223,N_15399,N_17361);
xnor U19224 (N_19224,N_17102,N_15037);
xnor U19225 (N_19225,N_16908,N_15152);
nor U19226 (N_19226,N_17213,N_17012);
nor U19227 (N_19227,N_17050,N_17468);
xnor U19228 (N_19228,N_16581,N_15418);
or U19229 (N_19229,N_15624,N_15083);
or U19230 (N_19230,N_15485,N_16994);
and U19231 (N_19231,N_17195,N_15692);
nor U19232 (N_19232,N_15870,N_16106);
or U19233 (N_19233,N_17196,N_16628);
xnor U19234 (N_19234,N_15063,N_16217);
or U19235 (N_19235,N_17490,N_17055);
and U19236 (N_19236,N_15697,N_15474);
or U19237 (N_19237,N_16196,N_15089);
xor U19238 (N_19238,N_15196,N_16414);
and U19239 (N_19239,N_16632,N_17054);
xor U19240 (N_19240,N_16249,N_15552);
nand U19241 (N_19241,N_16235,N_16622);
xor U19242 (N_19242,N_17178,N_16985);
nor U19243 (N_19243,N_16067,N_16836);
or U19244 (N_19244,N_15024,N_16023);
nand U19245 (N_19245,N_17342,N_16031);
and U19246 (N_19246,N_16764,N_15297);
nand U19247 (N_19247,N_15887,N_15786);
or U19248 (N_19248,N_15929,N_17327);
xnor U19249 (N_19249,N_16875,N_16146);
nand U19250 (N_19250,N_16689,N_16477);
and U19251 (N_19251,N_16059,N_16908);
nand U19252 (N_19252,N_17056,N_16392);
xor U19253 (N_19253,N_16684,N_15673);
nor U19254 (N_19254,N_16145,N_15413);
xnor U19255 (N_19255,N_16554,N_16694);
nor U19256 (N_19256,N_15269,N_15322);
nor U19257 (N_19257,N_16191,N_15411);
nor U19258 (N_19258,N_16811,N_17223);
xnor U19259 (N_19259,N_15740,N_15615);
nand U19260 (N_19260,N_16906,N_15866);
xor U19261 (N_19261,N_16194,N_15291);
nor U19262 (N_19262,N_16397,N_16429);
xor U19263 (N_19263,N_17418,N_15326);
xor U19264 (N_19264,N_15669,N_16218);
nor U19265 (N_19265,N_16434,N_16148);
nor U19266 (N_19266,N_15027,N_16279);
nor U19267 (N_19267,N_16149,N_16232);
nor U19268 (N_19268,N_16472,N_17203);
nor U19269 (N_19269,N_15433,N_15101);
xnor U19270 (N_19270,N_17400,N_15713);
xnor U19271 (N_19271,N_17151,N_15111);
or U19272 (N_19272,N_16213,N_15676);
and U19273 (N_19273,N_15698,N_16463);
nand U19274 (N_19274,N_16741,N_17146);
and U19275 (N_19275,N_17177,N_15403);
and U19276 (N_19276,N_15571,N_15783);
or U19277 (N_19277,N_15400,N_16999);
nand U19278 (N_19278,N_15752,N_17021);
nand U19279 (N_19279,N_16538,N_15370);
nand U19280 (N_19280,N_15292,N_15142);
and U19281 (N_19281,N_16217,N_16678);
nor U19282 (N_19282,N_16514,N_16833);
nor U19283 (N_19283,N_16244,N_17041);
nor U19284 (N_19284,N_16045,N_16532);
or U19285 (N_19285,N_16457,N_15267);
xor U19286 (N_19286,N_15858,N_16871);
xnor U19287 (N_19287,N_16256,N_15694);
or U19288 (N_19288,N_17400,N_16277);
and U19289 (N_19289,N_16380,N_16262);
or U19290 (N_19290,N_17197,N_16601);
and U19291 (N_19291,N_15175,N_16156);
nand U19292 (N_19292,N_15985,N_16057);
nor U19293 (N_19293,N_16825,N_17225);
nor U19294 (N_19294,N_16658,N_15765);
nand U19295 (N_19295,N_15478,N_17471);
and U19296 (N_19296,N_16756,N_15261);
nand U19297 (N_19297,N_16354,N_15318);
and U19298 (N_19298,N_17086,N_17032);
xor U19299 (N_19299,N_15483,N_15325);
nand U19300 (N_19300,N_16986,N_16334);
or U19301 (N_19301,N_17276,N_16009);
nor U19302 (N_19302,N_15773,N_15492);
nor U19303 (N_19303,N_16280,N_17133);
or U19304 (N_19304,N_15925,N_17215);
or U19305 (N_19305,N_16297,N_15517);
xnor U19306 (N_19306,N_16626,N_16514);
nor U19307 (N_19307,N_16585,N_16400);
or U19308 (N_19308,N_15759,N_16609);
and U19309 (N_19309,N_16946,N_16710);
and U19310 (N_19310,N_16489,N_16297);
nor U19311 (N_19311,N_15437,N_15503);
and U19312 (N_19312,N_17325,N_15240);
or U19313 (N_19313,N_17415,N_17051);
xor U19314 (N_19314,N_15401,N_15347);
nor U19315 (N_19315,N_15187,N_16435);
xnor U19316 (N_19316,N_17224,N_15513);
nor U19317 (N_19317,N_17282,N_15343);
xnor U19318 (N_19318,N_16918,N_15644);
xor U19319 (N_19319,N_15511,N_17462);
xor U19320 (N_19320,N_16350,N_17438);
and U19321 (N_19321,N_17087,N_17234);
and U19322 (N_19322,N_15608,N_16289);
nand U19323 (N_19323,N_15975,N_16055);
nor U19324 (N_19324,N_16987,N_16807);
xnor U19325 (N_19325,N_15992,N_16400);
or U19326 (N_19326,N_15439,N_15591);
nor U19327 (N_19327,N_17305,N_16217);
nand U19328 (N_19328,N_17479,N_16148);
and U19329 (N_19329,N_16457,N_16317);
nor U19330 (N_19330,N_16920,N_16980);
nor U19331 (N_19331,N_16918,N_15175);
and U19332 (N_19332,N_15067,N_17187);
nor U19333 (N_19333,N_15341,N_16151);
xor U19334 (N_19334,N_15554,N_17174);
nand U19335 (N_19335,N_17467,N_16307);
nor U19336 (N_19336,N_15098,N_15808);
nand U19337 (N_19337,N_15997,N_15327);
nand U19338 (N_19338,N_16379,N_15598);
or U19339 (N_19339,N_16828,N_15817);
or U19340 (N_19340,N_16739,N_15083);
and U19341 (N_19341,N_17106,N_15678);
nor U19342 (N_19342,N_15191,N_15636);
nand U19343 (N_19343,N_16527,N_15273);
and U19344 (N_19344,N_15754,N_15901);
xor U19345 (N_19345,N_15552,N_15785);
or U19346 (N_19346,N_15502,N_17137);
nand U19347 (N_19347,N_16723,N_15063);
and U19348 (N_19348,N_17028,N_17202);
and U19349 (N_19349,N_17260,N_16193);
and U19350 (N_19350,N_15039,N_17025);
and U19351 (N_19351,N_15875,N_15637);
xnor U19352 (N_19352,N_16773,N_16518);
nand U19353 (N_19353,N_17458,N_15746);
or U19354 (N_19354,N_15265,N_16326);
and U19355 (N_19355,N_16976,N_17168);
nand U19356 (N_19356,N_15995,N_15492);
and U19357 (N_19357,N_16048,N_15788);
or U19358 (N_19358,N_17212,N_16357);
nand U19359 (N_19359,N_15466,N_16164);
and U19360 (N_19360,N_16091,N_16880);
and U19361 (N_19361,N_15354,N_15460);
or U19362 (N_19362,N_16948,N_15576);
xor U19363 (N_19363,N_16277,N_15880);
nand U19364 (N_19364,N_15896,N_16210);
nand U19365 (N_19365,N_15461,N_16630);
and U19366 (N_19366,N_15127,N_17056);
and U19367 (N_19367,N_16602,N_15088);
and U19368 (N_19368,N_16864,N_15797);
xnor U19369 (N_19369,N_15217,N_17011);
nand U19370 (N_19370,N_15090,N_15325);
nor U19371 (N_19371,N_15513,N_15277);
or U19372 (N_19372,N_16086,N_15112);
xor U19373 (N_19373,N_17156,N_15399);
xor U19374 (N_19374,N_15963,N_15199);
xnor U19375 (N_19375,N_15962,N_16511);
and U19376 (N_19376,N_15399,N_15192);
nor U19377 (N_19377,N_15422,N_15627);
and U19378 (N_19378,N_15587,N_15888);
nor U19379 (N_19379,N_15677,N_17326);
nand U19380 (N_19380,N_17100,N_15049);
nand U19381 (N_19381,N_16759,N_15437);
nand U19382 (N_19382,N_15357,N_16148);
or U19383 (N_19383,N_15490,N_17496);
nand U19384 (N_19384,N_15249,N_17046);
and U19385 (N_19385,N_17021,N_16178);
nor U19386 (N_19386,N_17379,N_15082);
nor U19387 (N_19387,N_15433,N_15693);
xnor U19388 (N_19388,N_17208,N_16673);
or U19389 (N_19389,N_16568,N_16257);
nand U19390 (N_19390,N_16196,N_16911);
xnor U19391 (N_19391,N_15513,N_15605);
nand U19392 (N_19392,N_15496,N_16807);
nor U19393 (N_19393,N_17170,N_15539);
xnor U19394 (N_19394,N_17369,N_16413);
or U19395 (N_19395,N_15769,N_15410);
and U19396 (N_19396,N_15113,N_17209);
and U19397 (N_19397,N_16418,N_15762);
nand U19398 (N_19398,N_16345,N_15931);
or U19399 (N_19399,N_17384,N_17239);
nand U19400 (N_19400,N_15675,N_15276);
and U19401 (N_19401,N_15385,N_16653);
xnor U19402 (N_19402,N_16039,N_15190);
or U19403 (N_19403,N_16550,N_15818);
xnor U19404 (N_19404,N_17006,N_17186);
nand U19405 (N_19405,N_15694,N_15667);
xor U19406 (N_19406,N_16802,N_15629);
xor U19407 (N_19407,N_15978,N_17035);
nand U19408 (N_19408,N_15077,N_16079);
and U19409 (N_19409,N_15710,N_17367);
nor U19410 (N_19410,N_15519,N_16170);
or U19411 (N_19411,N_15844,N_15982);
xor U19412 (N_19412,N_17482,N_15204);
or U19413 (N_19413,N_17055,N_16942);
xor U19414 (N_19414,N_16775,N_16276);
and U19415 (N_19415,N_15973,N_16049);
xnor U19416 (N_19416,N_16504,N_16396);
or U19417 (N_19417,N_15630,N_16795);
or U19418 (N_19418,N_16501,N_15858);
or U19419 (N_19419,N_16193,N_16004);
or U19420 (N_19420,N_17073,N_15080);
nand U19421 (N_19421,N_16050,N_16842);
or U19422 (N_19422,N_17452,N_17279);
and U19423 (N_19423,N_16920,N_17353);
nand U19424 (N_19424,N_15847,N_16914);
xnor U19425 (N_19425,N_15775,N_15295);
and U19426 (N_19426,N_15210,N_15173);
xor U19427 (N_19427,N_17111,N_17166);
and U19428 (N_19428,N_17378,N_16445);
or U19429 (N_19429,N_15884,N_17092);
nor U19430 (N_19430,N_16138,N_17162);
and U19431 (N_19431,N_15221,N_17136);
or U19432 (N_19432,N_15910,N_16202);
nor U19433 (N_19433,N_15831,N_15649);
nor U19434 (N_19434,N_15421,N_15075);
or U19435 (N_19435,N_17232,N_16511);
and U19436 (N_19436,N_17046,N_16464);
xor U19437 (N_19437,N_17214,N_16174);
xnor U19438 (N_19438,N_16645,N_17403);
nor U19439 (N_19439,N_16748,N_15523);
or U19440 (N_19440,N_17379,N_16939);
nand U19441 (N_19441,N_16527,N_15338);
nor U19442 (N_19442,N_15105,N_16690);
xor U19443 (N_19443,N_15427,N_15466);
nor U19444 (N_19444,N_15588,N_17006);
and U19445 (N_19445,N_16299,N_17055);
or U19446 (N_19446,N_15116,N_15274);
nand U19447 (N_19447,N_16723,N_15205);
and U19448 (N_19448,N_16192,N_17004);
nand U19449 (N_19449,N_15360,N_17162);
or U19450 (N_19450,N_15323,N_16262);
nor U19451 (N_19451,N_15363,N_17349);
nand U19452 (N_19452,N_16831,N_15800);
or U19453 (N_19453,N_17166,N_15421);
xor U19454 (N_19454,N_17390,N_17265);
or U19455 (N_19455,N_15614,N_15184);
nand U19456 (N_19456,N_16056,N_15350);
nor U19457 (N_19457,N_15708,N_15456);
and U19458 (N_19458,N_15463,N_16884);
nand U19459 (N_19459,N_16201,N_17117);
and U19460 (N_19460,N_16762,N_15091);
or U19461 (N_19461,N_16357,N_16758);
nor U19462 (N_19462,N_15857,N_16736);
nor U19463 (N_19463,N_15022,N_16551);
nand U19464 (N_19464,N_15867,N_17351);
nor U19465 (N_19465,N_16414,N_16130);
and U19466 (N_19466,N_16857,N_16702);
nand U19467 (N_19467,N_17169,N_16716);
nor U19468 (N_19468,N_15477,N_16713);
xor U19469 (N_19469,N_16051,N_17339);
nand U19470 (N_19470,N_16640,N_15566);
nand U19471 (N_19471,N_17488,N_16428);
nand U19472 (N_19472,N_15570,N_15637);
nor U19473 (N_19473,N_15129,N_15273);
nor U19474 (N_19474,N_17497,N_17367);
xor U19475 (N_19475,N_15420,N_15913);
nand U19476 (N_19476,N_15087,N_15414);
xnor U19477 (N_19477,N_16578,N_17022);
nand U19478 (N_19478,N_16737,N_15293);
or U19479 (N_19479,N_16873,N_15614);
nor U19480 (N_19480,N_15616,N_16843);
xnor U19481 (N_19481,N_16664,N_17436);
nor U19482 (N_19482,N_15498,N_16008);
nand U19483 (N_19483,N_17291,N_15921);
or U19484 (N_19484,N_16320,N_15233);
nand U19485 (N_19485,N_17034,N_16160);
and U19486 (N_19486,N_17370,N_15321);
nor U19487 (N_19487,N_17218,N_15774);
and U19488 (N_19488,N_15366,N_16824);
nand U19489 (N_19489,N_17455,N_15300);
and U19490 (N_19490,N_15193,N_15811);
nand U19491 (N_19491,N_15732,N_15778);
nor U19492 (N_19492,N_17409,N_16363);
nor U19493 (N_19493,N_15699,N_15558);
nand U19494 (N_19494,N_16616,N_16026);
xnor U19495 (N_19495,N_15200,N_15277);
nand U19496 (N_19496,N_17048,N_16892);
xor U19497 (N_19497,N_16371,N_16794);
or U19498 (N_19498,N_16612,N_15468);
nor U19499 (N_19499,N_15217,N_16604);
nor U19500 (N_19500,N_16322,N_16320);
nor U19501 (N_19501,N_16188,N_15350);
nor U19502 (N_19502,N_15478,N_17198);
or U19503 (N_19503,N_16928,N_16321);
nor U19504 (N_19504,N_15158,N_15371);
nor U19505 (N_19505,N_15243,N_15827);
or U19506 (N_19506,N_15144,N_15985);
xnor U19507 (N_19507,N_17200,N_15250);
xor U19508 (N_19508,N_17388,N_15636);
and U19509 (N_19509,N_16536,N_15896);
nor U19510 (N_19510,N_15325,N_15950);
xnor U19511 (N_19511,N_15998,N_17384);
nor U19512 (N_19512,N_16098,N_15473);
nor U19513 (N_19513,N_17118,N_15645);
and U19514 (N_19514,N_17438,N_15779);
nor U19515 (N_19515,N_16915,N_15074);
nand U19516 (N_19516,N_16438,N_15936);
nor U19517 (N_19517,N_15631,N_15348);
nor U19518 (N_19518,N_17169,N_17322);
and U19519 (N_19519,N_15978,N_15466);
or U19520 (N_19520,N_16752,N_17086);
nor U19521 (N_19521,N_15541,N_16319);
xor U19522 (N_19522,N_15656,N_16420);
or U19523 (N_19523,N_15563,N_16213);
and U19524 (N_19524,N_15952,N_16728);
or U19525 (N_19525,N_16559,N_17161);
nor U19526 (N_19526,N_16976,N_16621);
nor U19527 (N_19527,N_15950,N_15672);
nor U19528 (N_19528,N_15126,N_17025);
nand U19529 (N_19529,N_16591,N_15444);
nor U19530 (N_19530,N_15689,N_15277);
and U19531 (N_19531,N_16903,N_15145);
xnor U19532 (N_19532,N_15695,N_15985);
nand U19533 (N_19533,N_16843,N_17061);
nand U19534 (N_19534,N_16286,N_16083);
xnor U19535 (N_19535,N_15171,N_15712);
xnor U19536 (N_19536,N_16811,N_17257);
xnor U19537 (N_19537,N_17496,N_15384);
xnor U19538 (N_19538,N_17242,N_15404);
or U19539 (N_19539,N_15999,N_17149);
xor U19540 (N_19540,N_17154,N_16383);
and U19541 (N_19541,N_15251,N_17293);
or U19542 (N_19542,N_16772,N_15545);
or U19543 (N_19543,N_17440,N_16720);
xnor U19544 (N_19544,N_17037,N_17213);
nor U19545 (N_19545,N_15051,N_15248);
nand U19546 (N_19546,N_16972,N_15766);
xor U19547 (N_19547,N_15824,N_15065);
nand U19548 (N_19548,N_16967,N_16096);
nor U19549 (N_19549,N_16126,N_15846);
or U19550 (N_19550,N_15229,N_16296);
nand U19551 (N_19551,N_17131,N_16085);
and U19552 (N_19552,N_15173,N_15030);
xnor U19553 (N_19553,N_16386,N_16950);
and U19554 (N_19554,N_16036,N_17294);
or U19555 (N_19555,N_16374,N_16147);
xor U19556 (N_19556,N_17258,N_17286);
xnor U19557 (N_19557,N_16125,N_15017);
nand U19558 (N_19558,N_16046,N_15795);
nor U19559 (N_19559,N_16563,N_15693);
xnor U19560 (N_19560,N_17390,N_16512);
nand U19561 (N_19561,N_17239,N_16595);
or U19562 (N_19562,N_15346,N_15588);
or U19563 (N_19563,N_16364,N_15001);
nand U19564 (N_19564,N_15177,N_16464);
nor U19565 (N_19565,N_16401,N_15947);
or U19566 (N_19566,N_15797,N_16513);
or U19567 (N_19567,N_16714,N_16221);
nor U19568 (N_19568,N_17036,N_16614);
xnor U19569 (N_19569,N_17444,N_15379);
nor U19570 (N_19570,N_17034,N_15217);
xor U19571 (N_19571,N_16103,N_16996);
nor U19572 (N_19572,N_15240,N_16487);
nor U19573 (N_19573,N_15539,N_16609);
nor U19574 (N_19574,N_17063,N_15403);
or U19575 (N_19575,N_16522,N_15578);
nor U19576 (N_19576,N_15990,N_16834);
xor U19577 (N_19577,N_15387,N_17032);
nor U19578 (N_19578,N_17384,N_17038);
or U19579 (N_19579,N_16452,N_15903);
nand U19580 (N_19580,N_16402,N_15641);
xnor U19581 (N_19581,N_16694,N_15670);
and U19582 (N_19582,N_15887,N_15344);
and U19583 (N_19583,N_15672,N_16959);
nand U19584 (N_19584,N_16421,N_17267);
or U19585 (N_19585,N_16536,N_15913);
and U19586 (N_19586,N_16200,N_15423);
nor U19587 (N_19587,N_16349,N_15637);
nor U19588 (N_19588,N_16634,N_15512);
or U19589 (N_19589,N_15206,N_15619);
and U19590 (N_19590,N_15751,N_16016);
and U19591 (N_19591,N_16881,N_15816);
and U19592 (N_19592,N_15337,N_15649);
nor U19593 (N_19593,N_17044,N_16679);
or U19594 (N_19594,N_15382,N_15805);
nand U19595 (N_19595,N_15127,N_15767);
nand U19596 (N_19596,N_15939,N_15954);
nor U19597 (N_19597,N_15223,N_16932);
and U19598 (N_19598,N_15449,N_15095);
nor U19599 (N_19599,N_16510,N_16599);
xor U19600 (N_19600,N_15748,N_15876);
nand U19601 (N_19601,N_17355,N_16921);
and U19602 (N_19602,N_15971,N_16298);
nor U19603 (N_19603,N_17076,N_16429);
and U19604 (N_19604,N_15030,N_16916);
nor U19605 (N_19605,N_17452,N_17180);
nor U19606 (N_19606,N_17377,N_15283);
nor U19607 (N_19607,N_15606,N_15812);
and U19608 (N_19608,N_16407,N_17353);
nor U19609 (N_19609,N_17461,N_16825);
xnor U19610 (N_19610,N_15972,N_17385);
xor U19611 (N_19611,N_17146,N_15188);
and U19612 (N_19612,N_16586,N_15148);
nand U19613 (N_19613,N_15770,N_16576);
xnor U19614 (N_19614,N_16548,N_15578);
and U19615 (N_19615,N_16779,N_15849);
nor U19616 (N_19616,N_16146,N_16697);
or U19617 (N_19617,N_17160,N_17323);
xor U19618 (N_19618,N_15660,N_16050);
nor U19619 (N_19619,N_17361,N_16793);
and U19620 (N_19620,N_15171,N_16405);
xnor U19621 (N_19621,N_16603,N_16968);
xnor U19622 (N_19622,N_16511,N_16196);
or U19623 (N_19623,N_16506,N_16400);
nor U19624 (N_19624,N_15219,N_17284);
nand U19625 (N_19625,N_15162,N_16788);
nor U19626 (N_19626,N_15480,N_16124);
or U19627 (N_19627,N_15158,N_16805);
or U19628 (N_19628,N_16806,N_16683);
xnor U19629 (N_19629,N_17475,N_17265);
nand U19630 (N_19630,N_15429,N_16850);
and U19631 (N_19631,N_15468,N_15333);
or U19632 (N_19632,N_15830,N_17105);
xor U19633 (N_19633,N_16630,N_17478);
and U19634 (N_19634,N_17144,N_17299);
xor U19635 (N_19635,N_17406,N_16312);
nor U19636 (N_19636,N_15244,N_17365);
xnor U19637 (N_19637,N_17489,N_17121);
or U19638 (N_19638,N_16262,N_15539);
nor U19639 (N_19639,N_16122,N_15964);
nand U19640 (N_19640,N_16472,N_16241);
nor U19641 (N_19641,N_16522,N_15944);
nand U19642 (N_19642,N_15372,N_15438);
xnor U19643 (N_19643,N_16308,N_15003);
xor U19644 (N_19644,N_16330,N_15059);
or U19645 (N_19645,N_17450,N_16164);
xor U19646 (N_19646,N_15368,N_15478);
and U19647 (N_19647,N_16768,N_16087);
nand U19648 (N_19648,N_15150,N_16959);
nand U19649 (N_19649,N_17312,N_16562);
and U19650 (N_19650,N_16564,N_15428);
and U19651 (N_19651,N_17301,N_16618);
nor U19652 (N_19652,N_15318,N_15976);
or U19653 (N_19653,N_15442,N_15957);
nand U19654 (N_19654,N_16832,N_15036);
nor U19655 (N_19655,N_16178,N_16998);
or U19656 (N_19656,N_15399,N_16643);
or U19657 (N_19657,N_17264,N_15333);
nand U19658 (N_19658,N_17174,N_15237);
nand U19659 (N_19659,N_15313,N_16119);
nand U19660 (N_19660,N_17214,N_16500);
nand U19661 (N_19661,N_16476,N_16059);
and U19662 (N_19662,N_16508,N_16709);
or U19663 (N_19663,N_15021,N_16373);
or U19664 (N_19664,N_15460,N_15772);
or U19665 (N_19665,N_17314,N_17092);
xnor U19666 (N_19666,N_16578,N_16582);
and U19667 (N_19667,N_16170,N_17482);
xor U19668 (N_19668,N_17187,N_17040);
and U19669 (N_19669,N_16813,N_15260);
xor U19670 (N_19670,N_15994,N_16002);
or U19671 (N_19671,N_16918,N_15196);
or U19672 (N_19672,N_17225,N_15448);
nand U19673 (N_19673,N_15688,N_15186);
nand U19674 (N_19674,N_15877,N_15435);
or U19675 (N_19675,N_15908,N_17151);
xor U19676 (N_19676,N_16240,N_15932);
or U19677 (N_19677,N_16643,N_17412);
xnor U19678 (N_19678,N_16799,N_16814);
or U19679 (N_19679,N_16991,N_15949);
nor U19680 (N_19680,N_16938,N_16358);
nand U19681 (N_19681,N_16220,N_16879);
nor U19682 (N_19682,N_17183,N_15819);
xnor U19683 (N_19683,N_15149,N_15711);
and U19684 (N_19684,N_15153,N_16350);
nor U19685 (N_19685,N_16219,N_16622);
xor U19686 (N_19686,N_16118,N_15626);
xnor U19687 (N_19687,N_16118,N_15343);
xor U19688 (N_19688,N_16199,N_15390);
nand U19689 (N_19689,N_15578,N_16427);
nor U19690 (N_19690,N_15504,N_15836);
nand U19691 (N_19691,N_15857,N_17459);
nor U19692 (N_19692,N_17494,N_16193);
nand U19693 (N_19693,N_17045,N_16416);
or U19694 (N_19694,N_16223,N_16603);
and U19695 (N_19695,N_16498,N_15966);
nor U19696 (N_19696,N_17366,N_16665);
nand U19697 (N_19697,N_15341,N_15793);
or U19698 (N_19698,N_17344,N_16812);
or U19699 (N_19699,N_16502,N_15574);
or U19700 (N_19700,N_17102,N_15775);
xnor U19701 (N_19701,N_15680,N_16823);
or U19702 (N_19702,N_16670,N_17202);
xor U19703 (N_19703,N_17167,N_15694);
and U19704 (N_19704,N_16587,N_17454);
nand U19705 (N_19705,N_16786,N_16112);
nand U19706 (N_19706,N_15542,N_17352);
nand U19707 (N_19707,N_17124,N_16506);
or U19708 (N_19708,N_15948,N_17251);
and U19709 (N_19709,N_16403,N_17113);
xor U19710 (N_19710,N_15793,N_16658);
nor U19711 (N_19711,N_17337,N_17464);
and U19712 (N_19712,N_17202,N_15228);
and U19713 (N_19713,N_16639,N_15887);
and U19714 (N_19714,N_15693,N_15453);
or U19715 (N_19715,N_16007,N_16089);
xor U19716 (N_19716,N_16007,N_16638);
nor U19717 (N_19717,N_15124,N_15028);
xor U19718 (N_19718,N_17451,N_15583);
or U19719 (N_19719,N_15275,N_15029);
or U19720 (N_19720,N_15272,N_16234);
or U19721 (N_19721,N_15676,N_17314);
nand U19722 (N_19722,N_17227,N_15943);
nor U19723 (N_19723,N_16917,N_15043);
nor U19724 (N_19724,N_15933,N_15643);
and U19725 (N_19725,N_15884,N_15146);
or U19726 (N_19726,N_17459,N_17164);
or U19727 (N_19727,N_15868,N_16432);
nand U19728 (N_19728,N_16089,N_16998);
nor U19729 (N_19729,N_15939,N_15203);
nor U19730 (N_19730,N_16036,N_16220);
or U19731 (N_19731,N_15828,N_17257);
or U19732 (N_19732,N_16988,N_17094);
or U19733 (N_19733,N_15658,N_16895);
and U19734 (N_19734,N_16164,N_16132);
nand U19735 (N_19735,N_15907,N_15084);
xor U19736 (N_19736,N_16755,N_15354);
xnor U19737 (N_19737,N_16461,N_16724);
or U19738 (N_19738,N_15418,N_15618);
or U19739 (N_19739,N_15411,N_15199);
and U19740 (N_19740,N_16906,N_15947);
nor U19741 (N_19741,N_16934,N_16805);
xnor U19742 (N_19742,N_15854,N_17080);
and U19743 (N_19743,N_16060,N_16272);
or U19744 (N_19744,N_17005,N_15576);
xnor U19745 (N_19745,N_17492,N_16494);
or U19746 (N_19746,N_15998,N_16348);
and U19747 (N_19747,N_16183,N_16516);
nor U19748 (N_19748,N_17047,N_15273);
or U19749 (N_19749,N_15331,N_15542);
nand U19750 (N_19750,N_15791,N_17438);
and U19751 (N_19751,N_15881,N_16545);
or U19752 (N_19752,N_15594,N_16748);
or U19753 (N_19753,N_17320,N_16175);
xor U19754 (N_19754,N_16133,N_15109);
nor U19755 (N_19755,N_17223,N_15502);
nor U19756 (N_19756,N_16645,N_16467);
nand U19757 (N_19757,N_15519,N_15299);
xor U19758 (N_19758,N_15019,N_16065);
and U19759 (N_19759,N_16416,N_17245);
and U19760 (N_19760,N_15492,N_15338);
nand U19761 (N_19761,N_15384,N_17168);
or U19762 (N_19762,N_16602,N_17317);
nand U19763 (N_19763,N_15299,N_16433);
nor U19764 (N_19764,N_15809,N_16708);
nand U19765 (N_19765,N_17267,N_16797);
nand U19766 (N_19766,N_17448,N_16040);
or U19767 (N_19767,N_17455,N_17116);
nor U19768 (N_19768,N_17447,N_16265);
nor U19769 (N_19769,N_15625,N_16829);
nand U19770 (N_19770,N_15473,N_16322);
nand U19771 (N_19771,N_15994,N_17109);
and U19772 (N_19772,N_16504,N_17176);
nor U19773 (N_19773,N_15545,N_17259);
xor U19774 (N_19774,N_15600,N_16348);
and U19775 (N_19775,N_15559,N_15358);
or U19776 (N_19776,N_17075,N_17341);
xor U19777 (N_19777,N_16277,N_15423);
nor U19778 (N_19778,N_16879,N_16503);
nand U19779 (N_19779,N_16852,N_15860);
xor U19780 (N_19780,N_15590,N_16145);
xor U19781 (N_19781,N_15510,N_17225);
and U19782 (N_19782,N_16238,N_15573);
or U19783 (N_19783,N_16169,N_15601);
nor U19784 (N_19784,N_16792,N_15943);
nor U19785 (N_19785,N_15153,N_15902);
or U19786 (N_19786,N_15107,N_16541);
and U19787 (N_19787,N_16197,N_15050);
nor U19788 (N_19788,N_15220,N_15307);
and U19789 (N_19789,N_15129,N_15825);
or U19790 (N_19790,N_16107,N_15612);
or U19791 (N_19791,N_15052,N_16451);
nor U19792 (N_19792,N_15037,N_16352);
xnor U19793 (N_19793,N_16955,N_17379);
nand U19794 (N_19794,N_15042,N_16092);
nand U19795 (N_19795,N_16780,N_17281);
and U19796 (N_19796,N_16606,N_17217);
or U19797 (N_19797,N_16703,N_15922);
nor U19798 (N_19798,N_17334,N_16089);
nor U19799 (N_19799,N_15682,N_15823);
and U19800 (N_19800,N_15075,N_15949);
nor U19801 (N_19801,N_16617,N_17462);
or U19802 (N_19802,N_15760,N_17036);
nand U19803 (N_19803,N_17020,N_16891);
xnor U19804 (N_19804,N_16085,N_16039);
xnor U19805 (N_19805,N_15368,N_15064);
nand U19806 (N_19806,N_17327,N_16672);
nor U19807 (N_19807,N_15996,N_17154);
xnor U19808 (N_19808,N_16244,N_15776);
xnor U19809 (N_19809,N_15924,N_16507);
or U19810 (N_19810,N_16000,N_15531);
nand U19811 (N_19811,N_17373,N_17053);
or U19812 (N_19812,N_15065,N_17392);
nand U19813 (N_19813,N_16838,N_15172);
or U19814 (N_19814,N_15482,N_16802);
xor U19815 (N_19815,N_16512,N_17415);
nor U19816 (N_19816,N_16561,N_15143);
or U19817 (N_19817,N_15338,N_16827);
or U19818 (N_19818,N_15283,N_17295);
and U19819 (N_19819,N_17396,N_15604);
or U19820 (N_19820,N_15282,N_17027);
xor U19821 (N_19821,N_17225,N_16493);
or U19822 (N_19822,N_15817,N_15447);
or U19823 (N_19823,N_15539,N_15832);
nand U19824 (N_19824,N_16834,N_16250);
xor U19825 (N_19825,N_16172,N_16378);
or U19826 (N_19826,N_16420,N_15886);
nand U19827 (N_19827,N_15178,N_15047);
nand U19828 (N_19828,N_15626,N_16998);
and U19829 (N_19829,N_16358,N_16235);
or U19830 (N_19830,N_16480,N_16513);
xor U19831 (N_19831,N_15488,N_16785);
xor U19832 (N_19832,N_15877,N_15409);
xor U19833 (N_19833,N_16317,N_17195);
xor U19834 (N_19834,N_17381,N_15106);
and U19835 (N_19835,N_15835,N_16813);
xor U19836 (N_19836,N_15068,N_17389);
and U19837 (N_19837,N_16773,N_15739);
xor U19838 (N_19838,N_17258,N_16213);
or U19839 (N_19839,N_16756,N_16056);
or U19840 (N_19840,N_16663,N_16707);
xnor U19841 (N_19841,N_15441,N_17374);
or U19842 (N_19842,N_15724,N_16530);
or U19843 (N_19843,N_16842,N_15580);
xor U19844 (N_19844,N_17022,N_17321);
nand U19845 (N_19845,N_16792,N_16673);
xnor U19846 (N_19846,N_15643,N_15368);
and U19847 (N_19847,N_17086,N_15216);
and U19848 (N_19848,N_15883,N_15863);
and U19849 (N_19849,N_16174,N_15562);
nor U19850 (N_19850,N_16705,N_17372);
nor U19851 (N_19851,N_16561,N_15539);
nor U19852 (N_19852,N_15347,N_15308);
nand U19853 (N_19853,N_17281,N_16309);
nor U19854 (N_19854,N_15171,N_16814);
or U19855 (N_19855,N_16341,N_17323);
nand U19856 (N_19856,N_15980,N_16036);
and U19857 (N_19857,N_16509,N_17411);
nand U19858 (N_19858,N_15792,N_16136);
xor U19859 (N_19859,N_15130,N_16316);
nor U19860 (N_19860,N_15242,N_15441);
and U19861 (N_19861,N_16214,N_15718);
and U19862 (N_19862,N_16844,N_16666);
xor U19863 (N_19863,N_15066,N_16208);
nor U19864 (N_19864,N_16654,N_16868);
xor U19865 (N_19865,N_15004,N_17227);
nand U19866 (N_19866,N_16657,N_15742);
or U19867 (N_19867,N_15025,N_16709);
xnor U19868 (N_19868,N_15807,N_16233);
and U19869 (N_19869,N_16998,N_16131);
nand U19870 (N_19870,N_15619,N_16800);
or U19871 (N_19871,N_17284,N_17057);
xnor U19872 (N_19872,N_15070,N_15208);
xnor U19873 (N_19873,N_16750,N_15310);
or U19874 (N_19874,N_16678,N_16794);
xnor U19875 (N_19875,N_16874,N_16363);
xor U19876 (N_19876,N_17465,N_15463);
or U19877 (N_19877,N_15664,N_16054);
and U19878 (N_19878,N_17377,N_15272);
or U19879 (N_19879,N_15022,N_16228);
nor U19880 (N_19880,N_17356,N_17183);
nor U19881 (N_19881,N_16640,N_16394);
nor U19882 (N_19882,N_17068,N_15507);
xor U19883 (N_19883,N_15520,N_15473);
or U19884 (N_19884,N_15187,N_17395);
or U19885 (N_19885,N_15070,N_16869);
nand U19886 (N_19886,N_15755,N_15743);
nand U19887 (N_19887,N_16018,N_17420);
xor U19888 (N_19888,N_16271,N_16407);
or U19889 (N_19889,N_15057,N_15164);
and U19890 (N_19890,N_16035,N_15702);
nor U19891 (N_19891,N_15418,N_15840);
nand U19892 (N_19892,N_15172,N_15361);
nand U19893 (N_19893,N_17369,N_15687);
nor U19894 (N_19894,N_15154,N_15242);
and U19895 (N_19895,N_16809,N_16663);
nand U19896 (N_19896,N_15698,N_15818);
nand U19897 (N_19897,N_16807,N_15837);
or U19898 (N_19898,N_16301,N_15395);
nor U19899 (N_19899,N_17391,N_16107);
xor U19900 (N_19900,N_17169,N_16971);
or U19901 (N_19901,N_15695,N_15391);
or U19902 (N_19902,N_17209,N_15019);
nor U19903 (N_19903,N_15818,N_17448);
xnor U19904 (N_19904,N_15915,N_15707);
nor U19905 (N_19905,N_15200,N_15926);
xor U19906 (N_19906,N_16142,N_16463);
xor U19907 (N_19907,N_17080,N_16734);
xor U19908 (N_19908,N_15784,N_16489);
nand U19909 (N_19909,N_15326,N_16561);
or U19910 (N_19910,N_17380,N_15850);
xor U19911 (N_19911,N_15740,N_16485);
and U19912 (N_19912,N_16055,N_16670);
nand U19913 (N_19913,N_16971,N_16410);
xnor U19914 (N_19914,N_16589,N_16982);
nor U19915 (N_19915,N_15782,N_17233);
nor U19916 (N_19916,N_16743,N_15774);
and U19917 (N_19917,N_16770,N_15586);
and U19918 (N_19918,N_15457,N_16506);
nand U19919 (N_19919,N_16166,N_15525);
nand U19920 (N_19920,N_16278,N_15225);
nand U19921 (N_19921,N_17266,N_15738);
nor U19922 (N_19922,N_16784,N_16150);
and U19923 (N_19923,N_16400,N_15509);
nand U19924 (N_19924,N_15890,N_16833);
or U19925 (N_19925,N_15806,N_15623);
and U19926 (N_19926,N_16412,N_15812);
or U19927 (N_19927,N_17392,N_16127);
nor U19928 (N_19928,N_16239,N_17379);
and U19929 (N_19929,N_16190,N_16680);
and U19930 (N_19930,N_15356,N_16612);
or U19931 (N_19931,N_15964,N_16489);
nor U19932 (N_19932,N_16162,N_17164);
or U19933 (N_19933,N_17014,N_16552);
nor U19934 (N_19934,N_15200,N_15747);
nor U19935 (N_19935,N_16601,N_17124);
xor U19936 (N_19936,N_15635,N_16765);
nand U19937 (N_19937,N_15321,N_17299);
nor U19938 (N_19938,N_16336,N_15024);
and U19939 (N_19939,N_17094,N_16946);
nand U19940 (N_19940,N_16043,N_17297);
and U19941 (N_19941,N_15327,N_16376);
xnor U19942 (N_19942,N_15559,N_16120);
nand U19943 (N_19943,N_15696,N_15949);
nand U19944 (N_19944,N_16558,N_17132);
nor U19945 (N_19945,N_15218,N_17047);
xnor U19946 (N_19946,N_15908,N_15888);
xor U19947 (N_19947,N_16484,N_15469);
or U19948 (N_19948,N_17061,N_16601);
nor U19949 (N_19949,N_16264,N_15369);
xnor U19950 (N_19950,N_16438,N_17326);
xor U19951 (N_19951,N_16276,N_15547);
and U19952 (N_19952,N_16738,N_15028);
nand U19953 (N_19953,N_15263,N_16101);
or U19954 (N_19954,N_16561,N_15694);
xor U19955 (N_19955,N_15981,N_15664);
and U19956 (N_19956,N_15781,N_17200);
or U19957 (N_19957,N_15067,N_15962);
nor U19958 (N_19958,N_15252,N_16935);
and U19959 (N_19959,N_15264,N_17179);
or U19960 (N_19960,N_16547,N_15637);
and U19961 (N_19961,N_16756,N_15229);
and U19962 (N_19962,N_16315,N_15332);
nor U19963 (N_19963,N_17073,N_15633);
and U19964 (N_19964,N_16139,N_16020);
xnor U19965 (N_19965,N_15799,N_17359);
nand U19966 (N_19966,N_17417,N_15897);
nand U19967 (N_19967,N_16498,N_15391);
nor U19968 (N_19968,N_16202,N_17319);
nand U19969 (N_19969,N_16519,N_16960);
or U19970 (N_19970,N_17270,N_15487);
nor U19971 (N_19971,N_17121,N_17244);
nor U19972 (N_19972,N_15849,N_17344);
or U19973 (N_19973,N_17277,N_17124);
or U19974 (N_19974,N_17455,N_15805);
nor U19975 (N_19975,N_16948,N_15429);
and U19976 (N_19976,N_15393,N_17481);
nor U19977 (N_19977,N_15781,N_16590);
and U19978 (N_19978,N_17204,N_16562);
nor U19979 (N_19979,N_16183,N_17236);
or U19980 (N_19980,N_17212,N_17337);
nand U19981 (N_19981,N_15950,N_16237);
or U19982 (N_19982,N_15942,N_15100);
and U19983 (N_19983,N_15450,N_16313);
or U19984 (N_19984,N_16048,N_17049);
nand U19985 (N_19985,N_15992,N_17074);
xnor U19986 (N_19986,N_16784,N_15350);
xor U19987 (N_19987,N_15157,N_16557);
nand U19988 (N_19988,N_16487,N_17174);
and U19989 (N_19989,N_15473,N_16507);
and U19990 (N_19990,N_15550,N_17185);
and U19991 (N_19991,N_16249,N_15800);
and U19992 (N_19992,N_15109,N_16046);
or U19993 (N_19993,N_17468,N_16629);
or U19994 (N_19994,N_15885,N_17248);
nand U19995 (N_19995,N_16951,N_15153);
nor U19996 (N_19996,N_16959,N_17036);
xnor U19997 (N_19997,N_16619,N_16187);
and U19998 (N_19998,N_16515,N_17158);
xnor U19999 (N_19999,N_15775,N_16932);
and U20000 (N_20000,N_17973,N_17591);
and U20001 (N_20001,N_18465,N_18849);
or U20002 (N_20002,N_19719,N_18612);
and U20003 (N_20003,N_17898,N_18911);
nand U20004 (N_20004,N_19276,N_19056);
nor U20005 (N_20005,N_17570,N_19922);
or U20006 (N_20006,N_19173,N_17517);
nor U20007 (N_20007,N_19963,N_19254);
xor U20008 (N_20008,N_19815,N_18402);
nand U20009 (N_20009,N_19337,N_18014);
nor U20010 (N_20010,N_18069,N_17752);
xnor U20011 (N_20011,N_18793,N_18901);
nor U20012 (N_20012,N_19491,N_18144);
or U20013 (N_20013,N_19722,N_18086);
or U20014 (N_20014,N_19425,N_17860);
or U20015 (N_20015,N_19852,N_18420);
and U20016 (N_20016,N_18288,N_17644);
or U20017 (N_20017,N_17954,N_18246);
xnor U20018 (N_20018,N_18076,N_19779);
nand U20019 (N_20019,N_19148,N_19451);
xor U20020 (N_20020,N_19913,N_18233);
and U20021 (N_20021,N_18831,N_19324);
or U20022 (N_20022,N_18674,N_19532);
nand U20023 (N_20023,N_19345,N_18422);
nor U20024 (N_20024,N_17607,N_18371);
nor U20025 (N_20025,N_17845,N_18613);
or U20026 (N_20026,N_17925,N_18324);
xor U20027 (N_20027,N_19608,N_17771);
and U20028 (N_20028,N_19320,N_19936);
xnor U20029 (N_20029,N_18467,N_18273);
and U20030 (N_20030,N_19756,N_19674);
nand U20031 (N_20031,N_19507,N_18515);
and U20032 (N_20032,N_19250,N_19831);
nor U20033 (N_20033,N_19099,N_19067);
nor U20034 (N_20034,N_18878,N_18764);
or U20035 (N_20035,N_19773,N_17783);
xnor U20036 (N_20036,N_17579,N_18451);
and U20037 (N_20037,N_18653,N_18463);
or U20038 (N_20038,N_18149,N_18815);
xnor U20039 (N_20039,N_19465,N_19906);
and U20040 (N_20040,N_19477,N_19270);
xnor U20041 (N_20041,N_19377,N_18956);
xor U20042 (N_20042,N_18182,N_19143);
nand U20043 (N_20043,N_18358,N_19241);
and U20044 (N_20044,N_18987,N_17541);
nor U20045 (N_20045,N_18944,N_19302);
nor U20046 (N_20046,N_17611,N_19058);
and U20047 (N_20047,N_19720,N_18430);
or U20048 (N_20048,N_18326,N_19182);
nor U20049 (N_20049,N_18130,N_18258);
nand U20050 (N_20050,N_18267,N_18279);
xnor U20051 (N_20051,N_19445,N_19764);
xor U20052 (N_20052,N_19338,N_18058);
nand U20053 (N_20053,N_18670,N_18100);
or U20054 (N_20054,N_19401,N_17618);
nor U20055 (N_20055,N_19725,N_18732);
or U20056 (N_20056,N_19277,N_19590);
or U20057 (N_20057,N_18973,N_19105);
or U20058 (N_20058,N_18360,N_18780);
or U20059 (N_20059,N_18364,N_19999);
and U20060 (N_20060,N_18209,N_18262);
nand U20061 (N_20061,N_18873,N_19778);
and U20062 (N_20062,N_19801,N_17828);
or U20063 (N_20063,N_17807,N_18630);
or U20064 (N_20064,N_18826,N_19861);
xor U20065 (N_20065,N_19935,N_18084);
xnor U20066 (N_20066,N_18984,N_18850);
and U20067 (N_20067,N_19592,N_19019);
or U20068 (N_20068,N_18458,N_18116);
nor U20069 (N_20069,N_18043,N_18204);
nand U20070 (N_20070,N_18718,N_18509);
and U20071 (N_20071,N_19979,N_17654);
or U20072 (N_20072,N_19329,N_18142);
or U20073 (N_20073,N_18589,N_19209);
and U20074 (N_20074,N_17521,N_18742);
and U20075 (N_20075,N_18398,N_18190);
nor U20076 (N_20076,N_18278,N_18841);
xnor U20077 (N_20077,N_17791,N_18401);
xor U20078 (N_20078,N_19095,N_18407);
or U20079 (N_20079,N_19600,N_18997);
xor U20080 (N_20080,N_19654,N_18047);
xor U20081 (N_20081,N_19718,N_18829);
and U20082 (N_20082,N_19761,N_19622);
and U20083 (N_20083,N_19016,N_18303);
and U20084 (N_20084,N_17645,N_19566);
and U20085 (N_20085,N_17887,N_18180);
or U20086 (N_20086,N_17581,N_18242);
xor U20087 (N_20087,N_18799,N_19141);
nand U20088 (N_20088,N_19111,N_18561);
and U20089 (N_20089,N_17946,N_19447);
and U20090 (N_20090,N_18853,N_19023);
or U20091 (N_20091,N_17933,N_19891);
or U20092 (N_20092,N_17693,N_18176);
and U20093 (N_20093,N_19998,N_19118);
nand U20094 (N_20094,N_18082,N_18281);
nand U20095 (N_20095,N_18221,N_19004);
nand U20096 (N_20096,N_17595,N_17503);
and U20097 (N_20097,N_19244,N_17883);
and U20098 (N_20098,N_18474,N_19269);
xor U20099 (N_20099,N_17533,N_17598);
xnor U20100 (N_20100,N_17605,N_19076);
nand U20101 (N_20101,N_19576,N_17620);
nor U20102 (N_20102,N_19112,N_18656);
and U20103 (N_20103,N_18934,N_19926);
xor U20104 (N_20104,N_19703,N_19154);
or U20105 (N_20105,N_18835,N_17586);
nor U20106 (N_20106,N_19029,N_19360);
and U20107 (N_20107,N_18601,N_17858);
nand U20108 (N_20108,N_19605,N_18717);
xnor U20109 (N_20109,N_18571,N_18808);
xnor U20110 (N_20110,N_19175,N_19835);
nor U20111 (N_20111,N_17934,N_19724);
or U20112 (N_20112,N_17944,N_18075);
and U20113 (N_20113,N_19033,N_18024);
nor U20114 (N_20114,N_19575,N_19663);
nand U20115 (N_20115,N_19267,N_19658);
nand U20116 (N_20116,N_19614,N_18498);
xor U20117 (N_20117,N_19496,N_19364);
nor U20118 (N_20118,N_19550,N_18165);
nand U20119 (N_20119,N_19647,N_19356);
nand U20120 (N_20120,N_18447,N_19129);
xnor U20121 (N_20121,N_17842,N_19909);
nor U20122 (N_20122,N_19069,N_19690);
nand U20123 (N_20123,N_18638,N_17950);
nor U20124 (N_20124,N_18170,N_18316);
nand U20125 (N_20125,N_18067,N_19051);
xor U20126 (N_20126,N_18197,N_17901);
xor U20127 (N_20127,N_17852,N_17646);
nand U20128 (N_20128,N_17709,N_18089);
nor U20129 (N_20129,N_18955,N_18198);
nand U20130 (N_20130,N_17781,N_18622);
nor U20131 (N_20131,N_19342,N_19196);
nand U20132 (N_20132,N_17970,N_19731);
nand U20133 (N_20133,N_18504,N_18148);
nor U20134 (N_20134,N_17879,N_18903);
xnor U20135 (N_20135,N_18918,N_17674);
or U20136 (N_20136,N_17544,N_18335);
nor U20137 (N_20137,N_19675,N_19730);
nand U20138 (N_20138,N_18887,N_19390);
nor U20139 (N_20139,N_18724,N_19279);
nand U20140 (N_20140,N_18369,N_19841);
and U20141 (N_20141,N_19140,N_19607);
and U20142 (N_20142,N_18833,N_18195);
or U20143 (N_20143,N_18909,N_18602);
nor U20144 (N_20144,N_18877,N_19085);
or U20145 (N_20145,N_19503,N_18529);
nand U20146 (N_20146,N_18794,N_19882);
nand U20147 (N_20147,N_18454,N_18244);
or U20148 (N_20148,N_17768,N_18660);
or U20149 (N_20149,N_17672,N_18415);
nor U20150 (N_20150,N_19316,N_19931);
nand U20151 (N_20151,N_18556,N_19122);
and U20152 (N_20152,N_17566,N_17535);
xnor U20153 (N_20153,N_19974,N_18658);
or U20154 (N_20154,N_18442,N_19977);
nand U20155 (N_20155,N_19744,N_19468);
or U20156 (N_20156,N_19948,N_19752);
and U20157 (N_20157,N_19312,N_18315);
nand U20158 (N_20158,N_18239,N_19704);
or U20159 (N_20159,N_19966,N_19934);
or U20160 (N_20160,N_19387,N_18910);
or U20161 (N_20161,N_18310,N_18203);
nand U20162 (N_20162,N_19262,N_19824);
nor U20163 (N_20163,N_18957,N_18605);
and U20164 (N_20164,N_18942,N_19010);
nor U20165 (N_20165,N_18517,N_19397);
and U20166 (N_20166,N_19457,N_19616);
nor U20167 (N_20167,N_18559,N_17732);
or U20168 (N_20168,N_18340,N_18889);
nand U20169 (N_20169,N_19746,N_19097);
xnor U20170 (N_20170,N_19484,N_18090);
nor U20171 (N_20171,N_19395,N_18205);
or U20172 (N_20172,N_18308,N_19827);
nor U20173 (N_20173,N_17710,N_19313);
or U20174 (N_20174,N_19193,N_18795);
nand U20175 (N_20175,N_19596,N_18830);
and U20176 (N_20176,N_19046,N_19449);
or U20177 (N_20177,N_17737,N_17751);
or U20178 (N_20178,N_18497,N_17715);
nor U20179 (N_20179,N_18035,N_18131);
or U20180 (N_20180,N_19783,N_18595);
nor U20181 (N_20181,N_19134,N_18277);
nor U20182 (N_20182,N_17866,N_18680);
nand U20183 (N_20183,N_19119,N_19346);
nor U20184 (N_20184,N_17941,N_17815);
xnor U20185 (N_20185,N_19200,N_18105);
xor U20186 (N_20186,N_18132,N_17844);
or U20187 (N_20187,N_19114,N_18744);
nor U20188 (N_20188,N_17801,N_18464);
nand U20189 (N_20189,N_19100,N_18749);
and U20190 (N_20190,N_17509,N_19971);
or U20191 (N_20191,N_18563,N_17692);
and U20192 (N_20192,N_18543,N_18624);
xnor U20193 (N_20193,N_17778,N_19167);
or U20194 (N_20194,N_19548,N_19866);
nand U20195 (N_20195,N_17892,N_17524);
nand U20196 (N_20196,N_18599,N_19867);
nor U20197 (N_20197,N_19836,N_18520);
nand U20198 (N_20198,N_19839,N_19304);
nor U20199 (N_20199,N_18557,N_19363);
or U20200 (N_20200,N_17758,N_19495);
and U20201 (N_20201,N_18140,N_19327);
or U20202 (N_20202,N_19463,N_18590);
or U20203 (N_20203,N_18238,N_18843);
or U20204 (N_20204,N_18542,N_19347);
nor U20205 (N_20205,N_19151,N_18797);
or U20206 (N_20206,N_17785,N_19003);
and U20207 (N_20207,N_19299,N_17580);
xnor U20208 (N_20208,N_18738,N_18922);
or U20209 (N_20209,N_17926,N_18490);
xnor U20210 (N_20210,N_19641,N_18582);
xor U20211 (N_20211,N_19450,N_19128);
nor U20212 (N_20212,N_18848,N_17914);
xnor U20213 (N_20213,N_18970,N_18023);
xnor U20214 (N_20214,N_19152,N_18450);
nor U20215 (N_20215,N_18354,N_18154);
nand U20216 (N_20216,N_19471,N_19405);
nor U20217 (N_20217,N_17929,N_18291);
and U20218 (N_20218,N_18917,N_18966);
and U20219 (N_20219,N_17540,N_19009);
nor U20220 (N_20220,N_19139,N_17742);
and U20221 (N_20221,N_17897,N_19514);
xor U20222 (N_20222,N_18857,N_19453);
nand U20223 (N_20223,N_18068,N_19384);
nor U20224 (N_20224,N_18899,N_19240);
nor U20225 (N_20225,N_18019,N_18768);
nand U20226 (N_20226,N_17585,N_19740);
or U20227 (N_20227,N_17964,N_19013);
and U20228 (N_20228,N_18696,N_18378);
nand U20229 (N_20229,N_18770,N_18048);
xnor U20230 (N_20230,N_18636,N_18339);
nand U20231 (N_20231,N_17673,N_19885);
xnor U20232 (N_20232,N_18269,N_18020);
or U20233 (N_20233,N_19753,N_19786);
or U20234 (N_20234,N_18568,N_18640);
or U20235 (N_20235,N_17888,N_18213);
and U20236 (N_20236,N_18760,N_19001);
nand U20237 (N_20237,N_17703,N_19766);
and U20238 (N_20238,N_19767,N_19245);
and U20239 (N_20239,N_19512,N_19020);
nor U20240 (N_20240,N_19452,N_18158);
and U20241 (N_20241,N_18964,N_17873);
nor U20242 (N_20242,N_18959,N_17655);
and U20243 (N_20243,N_17853,N_18384);
or U20244 (N_20244,N_17953,N_17619);
nor U20245 (N_20245,N_19082,N_17730);
or U20246 (N_20246,N_19919,N_19103);
nor U20247 (N_20247,N_17761,N_19601);
nand U20248 (N_20248,N_18778,N_18645);
nor U20249 (N_20249,N_19310,N_19775);
nand U20250 (N_20250,N_18336,N_19521);
and U20251 (N_20251,N_19127,N_18093);
nand U20252 (N_20252,N_19442,N_19096);
xor U20253 (N_20253,N_18280,N_18344);
or U20254 (N_20254,N_17664,N_19055);
nand U20255 (N_20255,N_17981,N_18210);
nor U20256 (N_20256,N_19043,N_18977);
nor U20257 (N_20257,N_17725,N_17832);
and U20258 (N_20258,N_19402,N_19696);
nand U20259 (N_20259,N_18684,N_18006);
xnor U20260 (N_20260,N_19899,N_19997);
xor U20261 (N_20261,N_19317,N_18252);
xnor U20262 (N_20262,N_19109,N_17938);
xor U20263 (N_20263,N_19933,N_19564);
nor U20264 (N_20264,N_18224,N_19093);
nor U20265 (N_20265,N_19849,N_19747);
nor U20266 (N_20266,N_18866,N_19281);
or U20267 (N_20267,N_17995,N_17958);
xnor U20268 (N_20268,N_19970,N_19102);
nor U20269 (N_20269,N_19263,N_19203);
nor U20270 (N_20270,N_19567,N_17916);
or U20271 (N_20271,N_19190,N_18828);
or U20272 (N_20272,N_19014,N_19782);
and U20273 (N_20273,N_19290,N_17790);
nor U20274 (N_20274,N_18581,N_18186);
nor U20275 (N_20275,N_18423,N_19079);
and U20276 (N_20276,N_18153,N_19274);
and U20277 (N_20277,N_18431,N_18033);
and U20278 (N_20278,N_18274,N_19878);
xnor U20279 (N_20279,N_19692,N_19407);
or U20280 (N_20280,N_17979,N_18791);
or U20281 (N_20281,N_19892,N_19462);
and U20282 (N_20282,N_17831,N_18410);
xor U20283 (N_20283,N_18177,N_19758);
or U20284 (N_20284,N_19220,N_19213);
xor U20285 (N_20285,N_17596,N_19264);
nand U20286 (N_20286,N_19538,N_17723);
xor U20287 (N_20287,N_18940,N_19392);
nor U20288 (N_20288,N_19958,N_19777);
xor U20289 (N_20289,N_18635,N_19678);
nor U20290 (N_20290,N_19309,N_19632);
and U20291 (N_20291,N_19502,N_18649);
nand U20292 (N_20292,N_18713,N_19604);
nor U20293 (N_20293,N_19186,N_19319);
or U20294 (N_20294,N_19938,N_18353);
or U20295 (N_20295,N_18160,N_18792);
nand U20296 (N_20296,N_18979,N_19519);
and U20297 (N_20297,N_18113,N_18604);
nand U20298 (N_20298,N_18372,N_17697);
nor U20299 (N_20299,N_19816,N_19625);
nor U20300 (N_20300,N_19195,N_18672);
nor U20301 (N_20301,N_19049,N_19711);
or U20302 (N_20302,N_18703,N_18508);
nor U20303 (N_20303,N_18620,N_18625);
xnor U20304 (N_20304,N_19523,N_19917);
nand U20305 (N_20305,N_19968,N_19957);
xnor U20306 (N_20306,N_18101,N_17635);
xnor U20307 (N_20307,N_19908,N_18477);
nand U20308 (N_20308,N_19757,N_17727);
nor U20309 (N_20309,N_17690,N_18247);
nor U20310 (N_20310,N_19661,N_17762);
or U20311 (N_20311,N_18096,N_18001);
xnor U20312 (N_20312,N_19559,N_19686);
and U20313 (N_20313,N_19833,N_19606);
xor U20314 (N_20314,N_19557,N_19573);
and U20315 (N_20315,N_19306,N_19236);
or U20316 (N_20316,N_17564,N_19094);
xor U20317 (N_20317,N_18173,N_18000);
nand U20318 (N_20318,N_19609,N_19699);
or U20319 (N_20319,N_18337,N_18462);
or U20320 (N_20320,N_17625,N_19469);
nand U20321 (N_20321,N_19965,N_18388);
and U20322 (N_20322,N_17743,N_17547);
nand U20323 (N_20323,N_17512,N_18054);
or U20324 (N_20324,N_19388,N_19296);
or U20325 (N_20325,N_19246,N_19930);
or U20326 (N_20326,N_18211,N_17658);
nand U20327 (N_20327,N_19983,N_18920);
nor U20328 (N_20328,N_19321,N_17928);
nand U20329 (N_20329,N_18623,N_19212);
xnor U20330 (N_20330,N_18255,N_19886);
nor U20331 (N_20331,N_19669,N_18057);
or U20332 (N_20332,N_19399,N_18259);
nor U20333 (N_20333,N_19283,N_19501);
nor U20334 (N_20334,N_17660,N_18208);
xor U20335 (N_20335,N_19499,N_18538);
or U20336 (N_20336,N_17532,N_19391);
and U20337 (N_20337,N_19727,N_18356);
nand U20338 (N_20338,N_19893,N_18932);
or U20339 (N_20339,N_19572,N_17889);
nor U20340 (N_20340,N_19166,N_17574);
xnor U20341 (N_20341,N_19701,N_18473);
or U20342 (N_20342,N_18924,N_18257);
nand U20343 (N_20343,N_19041,N_17683);
or U20344 (N_20344,N_19334,N_18106);
or U20345 (N_20345,N_19147,N_19640);
nor U20346 (N_20346,N_18567,N_18236);
xnor U20347 (N_20347,N_18135,N_17717);
nand U20348 (N_20348,N_19565,N_19047);
nand U20349 (N_20349,N_17506,N_18745);
or U20350 (N_20350,N_19207,N_17975);
xnor U20351 (N_20351,N_19822,N_17582);
nand U20352 (N_20352,N_19171,N_19184);
or U20353 (N_20353,N_18013,N_17840);
xnor U20354 (N_20354,N_18320,N_19634);
xnor U20355 (N_20355,N_17679,N_19707);
or U20356 (N_20356,N_17945,N_18689);
xor U20357 (N_20357,N_19921,N_19482);
xnor U20358 (N_20358,N_17738,N_19811);
xor U20359 (N_20359,N_19684,N_19568);
and U20360 (N_20360,N_18628,N_18097);
xnor U20361 (N_20361,N_19693,N_18010);
nand U20362 (N_20362,N_19403,N_19772);
or U20363 (N_20363,N_17553,N_19506);
or U20364 (N_20364,N_19860,N_18845);
nor U20365 (N_20365,N_18028,N_19064);
and U20366 (N_20366,N_19612,N_19574);
nor U20367 (N_20367,N_17802,N_18796);
and U20368 (N_20368,N_19736,N_19648);
nand U20369 (N_20369,N_19291,N_18935);
or U20370 (N_20370,N_17829,N_18521);
nor U20371 (N_20371,N_19856,N_19642);
nor U20372 (N_20372,N_18562,N_18731);
xnor U20373 (N_20373,N_19509,N_18648);
or U20374 (N_20374,N_18094,N_19176);
xor U20375 (N_20375,N_18382,N_19876);
or U20376 (N_20376,N_18725,N_19473);
and U20377 (N_20377,N_17707,N_17626);
and U20378 (N_20378,N_18588,N_18767);
nand U20379 (N_20379,N_19904,N_18884);
or U20380 (N_20380,N_19888,N_18968);
nand U20381 (N_20381,N_19526,N_19956);
or U20382 (N_20382,N_19052,N_19426);
nor U20383 (N_20383,N_19115,N_19982);
nor U20384 (N_20384,N_18237,N_18304);
xor U20385 (N_20385,N_18710,N_18234);
xor U20386 (N_20386,N_18699,N_18669);
and U20387 (N_20387,N_18871,N_18123);
and U20388 (N_20388,N_18004,N_19583);
or U20389 (N_20389,N_18061,N_19628);
nand U20390 (N_20390,N_17991,N_18307);
and U20391 (N_20391,N_19459,N_19946);
and U20392 (N_20392,N_18468,N_19687);
and U20393 (N_20393,N_17774,N_19163);
xor U20394 (N_20394,N_18074,N_19416);
nand U20395 (N_20395,N_19905,N_18800);
xor U20396 (N_20396,N_18720,N_19961);
or U20397 (N_20397,N_19895,N_19230);
nor U20398 (N_20398,N_19820,N_18129);
and U20399 (N_20399,N_17622,N_18389);
nand U20400 (N_20400,N_18188,N_19709);
or U20401 (N_20401,N_19768,N_19335);
or U20402 (N_20402,N_18298,N_18941);
xnor U20403 (N_20403,N_18548,N_18928);
and U20404 (N_20404,N_18663,N_19472);
xor U20405 (N_20405,N_18885,N_18958);
and U20406 (N_20406,N_19515,N_19884);
or U20407 (N_20407,N_19497,N_19536);
and U20408 (N_20408,N_19635,N_19443);
nand U20409 (N_20409,N_19900,N_18902);
nand U20410 (N_20410,N_19763,N_18930);
or U20411 (N_20411,N_17911,N_17731);
nor U20412 (N_20412,N_17992,N_18491);
and U20413 (N_20413,N_18499,N_18923);
nand U20414 (N_20414,N_19090,N_17859);
or U20415 (N_20415,N_18583,N_19098);
nor U20416 (N_20416,N_18708,N_18345);
or U20417 (N_20417,N_17968,N_19868);
or U20418 (N_20418,N_19551,N_18782);
nor U20419 (N_20419,N_18456,N_18719);
xor U20420 (N_20420,N_17977,N_18390);
or U20421 (N_20421,N_17657,N_18784);
or U20422 (N_20422,N_19932,N_19923);
nor U20423 (N_20423,N_18428,N_18781);
and U20424 (N_20424,N_17947,N_18592);
nor U20425 (N_20425,N_17969,N_17775);
and U20426 (N_20426,N_17675,N_18293);
and U20427 (N_20427,N_18925,N_18219);
or U20428 (N_20428,N_18801,N_18572);
or U20429 (N_20429,N_19570,N_19875);
xnor U20430 (N_20430,N_17538,N_19089);
nor U20431 (N_20431,N_18264,N_18155);
xor U20432 (N_20432,N_18042,N_19670);
nand U20433 (N_20433,N_18996,N_18394);
or U20434 (N_20434,N_17630,N_17502);
nand U20435 (N_20435,N_18951,N_17634);
or U20436 (N_20436,N_18120,N_18297);
xnor U20437 (N_20437,N_19879,N_19275);
and U20438 (N_20438,N_18697,N_17718);
and U20439 (N_20439,N_18196,N_19790);
xnor U20440 (N_20440,N_17716,N_19159);
xnor U20441 (N_20441,N_19417,N_19734);
nand U20442 (N_20442,N_17617,N_17592);
and U20443 (N_20443,N_18891,N_18493);
nor U20444 (N_20444,N_19863,N_17905);
nor U20445 (N_20445,N_17959,N_19649);
nand U20446 (N_20446,N_19234,N_18639);
nor U20447 (N_20447,N_19978,N_17702);
xnor U20448 (N_20448,N_19581,N_17680);
or U20449 (N_20449,N_19104,N_18145);
and U20450 (N_20450,N_19404,N_17767);
or U20451 (N_20451,N_18414,N_18416);
or U20452 (N_20452,N_19231,N_19000);
xnor U20453 (N_20453,N_17811,N_19537);
and U20454 (N_20454,N_19912,N_19819);
nor U20455 (N_20455,N_18365,N_18655);
nand U20456 (N_20456,N_17633,N_18954);
nand U20457 (N_20457,N_17554,N_17637);
or U20458 (N_20458,N_19042,N_18945);
nand U20459 (N_20459,N_18818,N_19421);
nand U20460 (N_20460,N_18174,N_19599);
nor U20461 (N_20461,N_18193,N_19698);
nor U20462 (N_20462,N_18164,N_18323);
xnor U20463 (N_20463,N_18051,N_19474);
and U20464 (N_20464,N_19695,N_17530);
nand U20465 (N_20465,N_17748,N_19774);
and U20466 (N_20466,N_19624,N_19610);
nor U20467 (N_20467,N_18694,N_18913);
nand U20468 (N_20468,N_19796,N_19406);
nand U20469 (N_20469,N_19708,N_18988);
or U20470 (N_20470,N_17960,N_18485);
nand U20471 (N_20471,N_19989,N_18466);
and U20472 (N_20472,N_19035,N_18788);
or U20473 (N_20473,N_18432,N_18730);
xor U20474 (N_20474,N_19528,N_18551);
xnor U20475 (N_20475,N_19880,N_17841);
nor U20476 (N_20476,N_18472,N_17906);
and U20477 (N_20477,N_19466,N_18633);
and U20478 (N_20478,N_19181,N_19224);
or U20479 (N_20479,N_18062,N_18534);
nor U20480 (N_20480,N_19222,N_18124);
nor U20481 (N_20481,N_19251,N_19427);
or U20482 (N_20482,N_17797,N_18265);
and U20483 (N_20483,N_18783,N_18434);
xnor U20484 (N_20484,N_19821,N_18757);
and U20485 (N_20485,N_18109,N_18540);
or U20486 (N_20486,N_18775,N_19508);
nor U20487 (N_20487,N_18117,N_18832);
nor U20488 (N_20488,N_19697,N_17756);
and U20489 (N_20489,N_19136,N_17627);
nand U20490 (N_20490,N_17910,N_18405);
nand U20491 (N_20491,N_17686,N_17563);
xnor U20492 (N_20492,N_19348,N_19994);
or U20493 (N_20493,N_18296,N_19343);
and U20494 (N_20494,N_18929,N_18514);
or U20495 (N_20495,N_17759,N_18199);
nand U20496 (N_20496,N_18050,N_18844);
nand U20497 (N_20497,N_18457,N_18285);
xor U20498 (N_20498,N_18448,N_18125);
nor U20499 (N_20499,N_18671,N_18693);
nor U20500 (N_20500,N_19541,N_19794);
or U20501 (N_20501,N_18009,N_18686);
or U20502 (N_20502,N_19024,N_18192);
nor U20503 (N_20503,N_19771,N_18126);
or U20504 (N_20504,N_17824,N_18867);
xnor U20505 (N_20505,N_18810,N_19848);
nor U20506 (N_20506,N_19705,N_18897);
nor U20507 (N_20507,N_17636,N_19619);
and U20508 (N_20508,N_17682,N_17653);
or U20509 (N_20509,N_18368,N_19394);
nor U20510 (N_20510,N_19784,N_18276);
nand U20511 (N_20511,N_18021,N_18709);
nand U20512 (N_20512,N_17862,N_19188);
and U20513 (N_20513,N_18552,N_19331);
xor U20514 (N_20514,N_19120,N_17561);
nor U20515 (N_20515,N_18723,N_18059);
nor U20516 (N_20516,N_19002,N_19239);
nor U20517 (N_20517,N_19988,N_19485);
or U20518 (N_20518,N_17921,N_19631);
and U20519 (N_20519,N_19877,N_19028);
xor U20520 (N_20520,N_17885,N_19301);
and U20521 (N_20521,N_19990,N_17770);
nor U20522 (N_20522,N_19488,N_17949);
nand U20523 (N_20523,N_19531,N_19265);
xor U20524 (N_20524,N_19543,N_18163);
and U20525 (N_20525,N_19735,N_17773);
xnor U20526 (N_20526,N_18769,N_18459);
and U20527 (N_20527,N_19637,N_18827);
and U20528 (N_20528,N_18282,N_19007);
nand U20529 (N_20529,N_18642,N_19925);
nor U20530 (N_20530,N_19106,N_17504);
xor U20531 (N_20531,N_17613,N_19621);
and U20532 (N_20532,N_18706,N_19791);
and U20533 (N_20533,N_18355,N_17780);
nor U20534 (N_20534,N_18044,N_18426);
and U20535 (N_20535,N_17578,N_18593);
nor U20536 (N_20536,N_17665,N_17576);
and U20537 (N_20537,N_18017,N_18321);
or U20538 (N_20538,N_18379,N_19257);
or U20539 (N_20539,N_19510,N_17930);
nor U20540 (N_20540,N_18519,N_18070);
nand U20541 (N_20541,N_19826,N_18138);
nor U20542 (N_20542,N_18095,N_17572);
and U20543 (N_20543,N_18151,N_18546);
xor U20544 (N_20544,N_17850,N_19578);
and U20545 (N_20545,N_19582,N_19593);
nand U20546 (N_20546,N_17684,N_19218);
nand U20547 (N_20547,N_19544,N_19890);
nor U20548 (N_20548,N_19470,N_19598);
xnor U20549 (N_20549,N_18251,N_17955);
xnor U20550 (N_20550,N_18361,N_17511);
xor U20551 (N_20551,N_18737,N_19738);
nor U20552 (N_20552,N_19591,N_18888);
nand U20553 (N_20553,N_19980,N_19872);
and U20554 (N_20554,N_18876,N_17837);
and U20555 (N_20555,N_18785,N_18092);
or U20556 (N_20556,N_18743,N_19185);
nand U20557 (N_20557,N_18518,N_18870);
nand U20558 (N_20558,N_17594,N_19396);
xnor U20559 (N_20559,N_18346,N_19202);
nor U20560 (N_20560,N_18270,N_17875);
nand U20561 (N_20561,N_19149,N_19288);
nand U20562 (N_20562,N_17940,N_19759);
and U20563 (N_20563,N_18982,N_18175);
nor U20564 (N_20564,N_19535,N_19483);
and U20565 (N_20565,N_18882,N_19344);
nor U20566 (N_20566,N_18185,N_17918);
nand U20567 (N_20567,N_17724,N_18501);
xnor U20568 (N_20568,N_19243,N_19145);
xor U20569 (N_20569,N_17868,N_19955);
or U20570 (N_20570,N_19993,N_17500);
nor U20571 (N_20571,N_19393,N_18650);
or U20572 (N_20572,N_19242,N_17990);
nor U20573 (N_20573,N_17501,N_18161);
nand U20574 (N_20574,N_18409,N_19553);
nor U20575 (N_20575,N_17830,N_18895);
nand U20576 (N_20576,N_18541,N_19737);
and U20577 (N_20577,N_18741,N_19838);
nor U20578 (N_20578,N_18790,N_19339);
nand U20579 (N_20579,N_18606,N_19065);
xor U20580 (N_20580,N_18046,N_17784);
and U20581 (N_20581,N_17652,N_18936);
xor U20582 (N_20582,N_17722,N_17825);
xnor U20583 (N_20583,N_18535,N_19691);
and U20584 (N_20584,N_17777,N_19563);
or U20585 (N_20585,N_18350,N_17745);
nor U20586 (N_20586,N_17719,N_19305);
xnor U20587 (N_20587,N_17855,N_19694);
nor U20588 (N_20588,N_19681,N_17839);
nor U20589 (N_20589,N_17843,N_18607);
xor U20590 (N_20590,N_18981,N_18055);
nor U20591 (N_20591,N_18322,N_17912);
xor U20592 (N_20592,N_19739,N_19336);
xnor U20593 (N_20593,N_18927,N_19742);
or U20594 (N_20594,N_19813,N_18376);
or U20595 (N_20595,N_19375,N_18726);
or U20596 (N_20596,N_19386,N_18565);
and U20597 (N_20597,N_18805,N_19529);
and U20598 (N_20598,N_18367,N_19741);
and U20599 (N_20599,N_19797,N_18272);
or U20600 (N_20600,N_19927,N_19048);
nand U20601 (N_20601,N_17820,N_18091);
and U20602 (N_20602,N_19062,N_17608);
or U20603 (N_20603,N_18370,N_18494);
and U20604 (N_20604,N_18578,N_19333);
nor U20605 (N_20605,N_18391,N_19898);
xor U20606 (N_20606,N_18617,N_18399);
and U20607 (N_20607,N_18716,N_17913);
and U20608 (N_20608,N_19644,N_18860);
and U20609 (N_20609,N_18919,N_17817);
nor U20610 (N_20610,N_19116,N_18654);
and U20611 (N_20611,N_18879,N_19793);
or U20612 (N_20612,N_19754,N_18122);
nor U20613 (N_20613,N_17942,N_19645);
or U20614 (N_20614,N_19776,N_18143);
or U20615 (N_20615,N_19969,N_18965);
xnor U20616 (N_20616,N_17863,N_19135);
or U20617 (N_20617,N_18359,N_19562);
nor U20618 (N_20618,N_18381,N_18812);
xor U20619 (N_20619,N_17746,N_17629);
and U20620 (N_20620,N_18937,N_19383);
and U20621 (N_20621,N_17939,N_18216);
nand U20622 (N_20622,N_19897,N_19133);
xor U20623 (N_20623,N_17896,N_18816);
and U20624 (N_20624,N_18331,N_17721);
or U20625 (N_20625,N_18228,N_18445);
or U20626 (N_20626,N_18644,N_18861);
nor U20627 (N_20627,N_18947,N_17798);
and U20628 (N_20628,N_19716,N_18475);
and U20629 (N_20629,N_17516,N_17537);
nor U20630 (N_20630,N_17776,N_18994);
or U20631 (N_20631,N_19018,N_18207);
nor U20632 (N_20632,N_19733,N_18286);
xnor U20633 (N_20633,N_17808,N_17836);
and U20634 (N_20634,N_19174,N_19762);
nand U20635 (N_20635,N_18438,N_18496);
nor U20636 (N_20636,N_18102,N_17861);
nor U20637 (N_20637,N_19683,N_18217);
and U20638 (N_20638,N_18201,N_19032);
xnor U20639 (N_20639,N_19547,N_17809);
and U20640 (N_20640,N_18727,N_18524);
and U20641 (N_20641,N_19676,N_18118);
nor U20642 (N_20642,N_17668,N_19289);
xor U20643 (N_20643,N_18411,N_19361);
or U20644 (N_20644,N_18275,N_18036);
nand U20645 (N_20645,N_17505,N_19286);
or U20646 (N_20646,N_17662,N_18516);
or U20647 (N_20647,N_17834,N_18698);
and U20648 (N_20648,N_18972,N_19237);
nor U20649 (N_20649,N_19430,N_19353);
xnor U20650 (N_20650,N_17602,N_18787);
or U20651 (N_20651,N_18759,N_18191);
xnor U20652 (N_20652,N_17584,N_19155);
and U20653 (N_20653,N_19354,N_19297);
or U20654 (N_20654,N_18931,N_18375);
nor U20655 (N_20655,N_19370,N_18235);
and U20656 (N_20656,N_19198,N_19549);
nand U20657 (N_20657,N_18063,N_18439);
nor U20658 (N_20658,N_19984,N_17667);
and U20659 (N_20659,N_18597,N_19380);
or U20660 (N_20660,N_17599,N_19210);
nand U20661 (N_20661,N_18011,N_19688);
nand U20662 (N_20662,N_19178,N_19987);
nor U20663 (N_20663,N_17542,N_17971);
and U20664 (N_20664,N_18777,N_18962);
nor U20665 (N_20665,N_17548,N_19814);
nor U20666 (N_20666,N_19072,N_19996);
or U20667 (N_20667,N_18218,N_18482);
nor U20668 (N_20668,N_18290,N_17565);
nor U20669 (N_20669,N_19788,N_18253);
nand U20670 (N_20670,N_18488,N_18002);
or U20671 (N_20671,N_19755,N_18666);
nor U20672 (N_20672,N_17757,N_18026);
xnor U20673 (N_20673,N_19124,N_18967);
xnor U20674 (N_20674,N_19962,N_18121);
or U20675 (N_20675,N_19428,N_18025);
nand U20676 (N_20676,N_17508,N_19086);
nor U20677 (N_20677,N_18157,N_18045);
xnor U20678 (N_20678,N_17936,N_17543);
or U20679 (N_20679,N_17531,N_19039);
nand U20680 (N_20680,N_19480,N_19187);
xor U20681 (N_20681,N_19271,N_18798);
or U20682 (N_20682,N_18421,N_17823);
nor U20683 (N_20683,N_19197,N_19308);
nand U20684 (N_20684,N_18834,N_19942);
xnor U20685 (N_20685,N_19054,N_17706);
nand U20686 (N_20686,N_18038,N_19597);
nand U20687 (N_20687,N_18260,N_18362);
xnor U20688 (N_20688,N_19323,N_19138);
and U20689 (N_20689,N_17688,N_18858);
xnor U20690 (N_20690,N_18225,N_19802);
xor U20691 (N_20691,N_18111,N_18373);
xnor U20692 (N_20692,N_19318,N_18859);
nand U20693 (N_20693,N_17567,N_19545);
nor U20694 (N_20694,N_19374,N_18240);
nor U20695 (N_20695,N_19579,N_17904);
xnor U20696 (N_20696,N_18425,N_18141);
nand U20697 (N_20697,N_17670,N_18975);
and U20698 (N_20698,N_19038,N_18007);
nand U20699 (N_20699,N_17812,N_19432);
xor U20700 (N_20700,N_17974,N_19087);
xnor U20701 (N_20701,N_17650,N_19940);
nand U20702 (N_20702,N_19855,N_17604);
nor U20703 (N_20703,N_19221,N_18429);
or U20704 (N_20704,N_18933,N_18687);
and U20705 (N_20705,N_19179,N_18729);
or U20706 (N_20706,N_19225,N_19907);
xnor U20707 (N_20707,N_18080,N_18573);
and U20708 (N_20708,N_17803,N_19525);
nand U20709 (N_20709,N_19303,N_17849);
xnor U20710 (N_20710,N_18609,N_18295);
and U20711 (N_20711,N_17838,N_18479);
or U20712 (N_20712,N_19369,N_19022);
and U20713 (N_20713,N_19494,N_17513);
and U20714 (N_20714,N_19729,N_18591);
or U20715 (N_20715,N_18854,N_19527);
and U20716 (N_20716,N_18580,N_18079);
nand U20717 (N_20717,N_17978,N_19721);
nand U20718 (N_20718,N_19967,N_17639);
nor U20719 (N_20719,N_18668,N_18313);
xnor U20720 (N_20720,N_18169,N_17787);
nor U20721 (N_20721,N_17821,N_19618);
and U20722 (N_20722,N_18053,N_17782);
xnor U20723 (N_20723,N_19493,N_18309);
nand U20724 (N_20724,N_18608,N_19216);
xor U20725 (N_20725,N_17691,N_18115);
or U20726 (N_20726,N_19662,N_18107);
nand U20727 (N_20727,N_18081,N_17569);
nor U20728 (N_20728,N_19467,N_18470);
and U20729 (N_20729,N_18245,N_18736);
or U20730 (N_20730,N_19362,N_19850);
xor U20731 (N_20731,N_18946,N_17744);
nand U20732 (N_20732,N_17902,N_19858);
nand U20733 (N_20733,N_19518,N_17813);
and U20734 (N_20734,N_17624,N_18446);
nand U20735 (N_20735,N_17518,N_18898);
nand U20736 (N_20736,N_18950,N_17612);
xnor U20737 (N_20737,N_17534,N_19659);
xnor U20738 (N_20738,N_19533,N_19194);
nor U20739 (N_20739,N_19229,N_19411);
nand U20740 (N_20740,N_19728,N_18487);
xnor U20741 (N_20741,N_19585,N_19172);
xnor U20742 (N_20742,N_19828,N_18461);
nor U20743 (N_20743,N_19400,N_18953);
and U20744 (N_20744,N_17962,N_19439);
nand U20745 (N_20745,N_18998,N_19456);
nand U20746 (N_20746,N_18611,N_18500);
and U20747 (N_20747,N_19045,N_17671);
nor U20748 (N_20748,N_17590,N_19434);
or U20749 (N_20749,N_19382,N_17510);
or U20750 (N_20750,N_18223,N_17891);
and U20751 (N_20751,N_19520,N_17708);
and U20752 (N_20752,N_19939,N_17677);
nor U20753 (N_20753,N_17577,N_17822);
and U20754 (N_20754,N_17733,N_18301);
and U20755 (N_20755,N_17994,N_19253);
and U20756 (N_20756,N_19615,N_18318);
or U20757 (N_20757,N_19078,N_19280);
and U20758 (N_20758,N_19044,N_18881);
or U20759 (N_20759,N_19611,N_19580);
xnor U20760 (N_20760,N_18673,N_19180);
xor U20761 (N_20761,N_17967,N_17552);
xor U20762 (N_20762,N_18249,N_18271);
nor U20763 (N_20763,N_18809,N_18078);
nor U20764 (N_20764,N_18691,N_19441);
or U20765 (N_20765,N_19673,N_19256);
nand U20766 (N_20766,N_17701,N_17632);
or U20767 (N_20767,N_18403,N_17689);
and U20768 (N_20768,N_17800,N_17870);
nor U20769 (N_20769,N_19025,N_18427);
nand U20770 (N_20770,N_19712,N_18900);
and U20771 (N_20771,N_17874,N_19745);
or U20772 (N_20772,N_18547,N_19057);
or U20773 (N_20773,N_17847,N_18762);
or U20774 (N_20774,N_19806,N_19646);
and U20775 (N_20775,N_19871,N_19255);
xnor U20776 (N_20776,N_18453,N_17519);
xnor U20777 (N_20777,N_18299,N_18733);
or U20778 (N_20778,N_18495,N_18661);
xnor U20779 (N_20779,N_19804,N_19170);
and U20780 (N_20780,N_19571,N_17545);
xor U20781 (N_20781,N_17982,N_18016);
and U20782 (N_20782,N_17884,N_17961);
xnor U20783 (N_20783,N_19322,N_18851);
nand U20784 (N_20784,N_17614,N_19371);
nor U20785 (N_20785,N_18452,N_18735);
nand U20786 (N_20786,N_18380,N_18734);
xor U20787 (N_20787,N_17997,N_18814);
and U20788 (N_20788,N_19546,N_19889);
nand U20789 (N_20789,N_17818,N_19666);
nor U20790 (N_20790,N_18437,N_18227);
nand U20791 (N_20791,N_17877,N_19588);
nor U20792 (N_20792,N_19260,N_19415);
xnor U20793 (N_20793,N_19294,N_18916);
nor U20794 (N_20794,N_17907,N_19944);
nor U20795 (N_20795,N_19132,N_19300);
xnor U20796 (N_20796,N_19702,N_19613);
and U20797 (N_20797,N_18863,N_19126);
and U20798 (N_20798,N_17694,N_19760);
nand U20799 (N_20799,N_19706,N_19081);
and U20800 (N_20800,N_18072,N_19870);
xnor U20801 (N_20801,N_18419,N_17589);
and U20802 (N_20802,N_17766,N_18560);
nor U20803 (N_20803,N_17999,N_19513);
or U20804 (N_20804,N_19315,N_19843);
nor U20805 (N_20805,N_19682,N_17765);
nand U20806 (N_20806,N_18266,N_19036);
nand U20807 (N_20807,N_18400,N_18688);
nand U20808 (N_20808,N_18893,N_17747);
or U20809 (N_20809,N_18821,N_18677);
xnor U20810 (N_20810,N_19558,N_17856);
nor U20811 (N_20811,N_18596,N_18136);
nand U20812 (N_20812,N_19227,N_19656);
nor U20813 (N_20813,N_18652,N_18890);
and U20814 (N_20814,N_18449,N_19005);
or U20815 (N_20815,N_17551,N_17687);
or U20816 (N_20816,N_19602,N_19498);
and U20817 (N_20817,N_18682,N_19249);
and U20818 (N_20818,N_18317,N_19351);
nand U20819 (N_20819,N_17980,N_18119);
or U20820 (N_20820,N_18338,N_18779);
nor U20821 (N_20821,N_18531,N_19995);
xor U20822 (N_20822,N_17583,N_18087);
xnor U20823 (N_20823,N_19101,N_18341);
or U20824 (N_20824,N_17867,N_19652);
and U20825 (N_20825,N_18505,N_19372);
and U20826 (N_20826,N_19454,N_17539);
xnor U20827 (N_20827,N_19832,N_19063);
nor U20828 (N_20828,N_17638,N_19478);
nor U20829 (N_20829,N_19689,N_19807);
nand U20830 (N_20830,N_19710,N_18681);
nand U20831 (N_20831,N_18484,N_18554);
nand U20832 (N_20832,N_19985,N_19438);
xnor U20833 (N_20833,N_18085,N_18511);
nor U20834 (N_20834,N_19358,N_19812);
or U20835 (N_20835,N_19869,N_18864);
or U20836 (N_20836,N_19413,N_18202);
xor U20837 (N_20837,N_18980,N_18527);
nor U20838 (N_20838,N_18753,N_19053);
nor U20839 (N_20839,N_18222,N_19715);
xor U20840 (N_20840,N_18184,N_19205);
or U20841 (N_20841,N_17894,N_18108);
nor U20842 (N_20842,N_19084,N_19770);
nor U20843 (N_20843,N_18305,N_18049);
or U20844 (N_20844,N_19340,N_17741);
or U20845 (N_20845,N_18386,N_18314);
nor U20846 (N_20846,N_19113,N_18865);
nand U20847 (N_20847,N_19153,N_19424);
xnor U20848 (N_20848,N_17895,N_19412);
or U20849 (N_20849,N_17550,N_18478);
nor U20850 (N_20850,N_18395,N_19887);
and U20851 (N_20851,N_19359,N_18231);
or U20852 (N_20852,N_19298,N_17819);
nand U20853 (N_20853,N_18088,N_18528);
or U20854 (N_20854,N_17750,N_18906);
nor U20855 (N_20855,N_19522,N_17786);
and U20856 (N_20856,N_19556,N_17763);
and U20857 (N_20857,N_17698,N_19748);
and U20858 (N_20858,N_19408,N_18990);
xor U20859 (N_20859,N_19458,N_19379);
xor U20860 (N_20860,N_18545,N_17857);
and U20861 (N_20861,N_17659,N_17527);
or U20862 (N_20862,N_18667,N_17736);
or U20863 (N_20863,N_19829,N_18214);
nor U20864 (N_20864,N_19924,N_17616);
and U20865 (N_20865,N_18243,N_19121);
nand U20866 (N_20866,N_17899,N_17963);
and U20867 (N_20867,N_18664,N_18683);
and U20868 (N_20868,N_18992,N_18641);
nand U20869 (N_20869,N_19123,N_17526);
and U20870 (N_20870,N_18526,N_18896);
and U20871 (N_20871,N_17601,N_17643);
and U20872 (N_20872,N_19131,N_18908);
nand U20873 (N_20873,N_17755,N_18302);
xor U20874 (N_20874,N_19341,N_19552);
nand U20875 (N_20875,N_18347,N_18676);
and U20876 (N_20876,N_19431,N_18030);
or U20877 (N_20877,N_19295,N_19750);
or U20878 (N_20878,N_19325,N_18629);
xor U20879 (N_20879,N_17536,N_18436);
or U20880 (N_20880,N_18241,N_17796);
nor U20881 (N_20881,N_19077,N_18110);
xnor U20882 (N_20882,N_18418,N_18230);
or U20883 (N_20883,N_17794,N_19945);
nor U20884 (N_20884,N_19307,N_18146);
or U20885 (N_20885,N_18993,N_19943);
nand U20886 (N_20886,N_19381,N_18083);
nor U20887 (N_20887,N_19328,N_18585);
nand U20888 (N_20888,N_18481,N_17986);
xor U20889 (N_20889,N_19830,N_17876);
nor U20890 (N_20890,N_18200,N_17587);
or U20891 (N_20891,N_18763,N_18575);
xor U20892 (N_20892,N_19660,N_18530);
nor U20893 (N_20893,N_19991,N_17835);
nor U20894 (N_20894,N_17799,N_17700);
and U20895 (N_20895,N_19657,N_19883);
xor U20896 (N_20896,N_17764,N_17972);
nor U20897 (N_20897,N_18804,N_17558);
xnor U20898 (N_20898,N_18943,N_18598);
and U20899 (N_20899,N_18306,N_18952);
nand U20900 (N_20900,N_18071,N_17965);
nor U20901 (N_20901,N_17720,N_18705);
xnor U20902 (N_20902,N_17681,N_19158);
and U20903 (N_20903,N_18536,N_17656);
nor U20904 (N_20904,N_19017,N_19150);
or U20905 (N_20905,N_19500,N_19714);
and U20906 (N_20906,N_18675,N_19070);
nand U20907 (N_20907,N_17923,N_19840);
xnor U20908 (N_20908,N_17920,N_18015);
nand U20909 (N_20909,N_18512,N_18150);
or U20910 (N_20910,N_19700,N_18766);
nand U20911 (N_20911,N_18976,N_18077);
and U20912 (N_20912,N_19617,N_19080);
xnor U20913 (N_20913,N_19420,N_17562);
xnor U20914 (N_20914,N_18872,N_19075);
nand U20915 (N_20915,N_18312,N_18393);
and U20916 (N_20916,N_19765,N_18647);
and U20917 (N_20917,N_17871,N_18690);
or U20918 (N_20918,N_18969,N_18751);
nand U20919 (N_20919,N_18949,N_17666);
xor U20920 (N_20920,N_19589,N_18406);
and U20921 (N_20921,N_19517,N_18254);
and U20922 (N_20922,N_17983,N_17931);
xnor U20923 (N_20923,N_18147,N_18029);
nand U20924 (N_20924,N_19422,N_19037);
and U20925 (N_20925,N_17712,N_18250);
and U20926 (N_20926,N_18978,N_19959);
and U20927 (N_20927,N_19929,N_19629);
and U20928 (N_20928,N_18875,N_19183);
nand U20929 (N_20929,N_17623,N_17989);
xor U20930 (N_20930,N_19894,N_17575);
xnor U20931 (N_20931,N_18342,N_17878);
nand U20932 (N_20932,N_18363,N_18172);
nor U20933 (N_20933,N_19146,N_18506);
nand U20934 (N_20934,N_18983,N_18614);
or U20935 (N_20935,N_19650,N_18824);
nand U20936 (N_20936,N_19685,N_18619);
nand U20937 (N_20937,N_18892,N_18584);
or U20938 (N_20938,N_18776,N_19620);
and U20939 (N_20939,N_18558,N_19789);
and U20940 (N_20940,N_19357,N_19259);
xnor U20941 (N_20941,N_19258,N_19554);
and U20942 (N_20942,N_18907,N_19460);
nand U20943 (N_20943,N_19160,N_18349);
nand U20944 (N_20944,N_18471,N_18586);
xor U20945 (N_20945,N_17754,N_19847);
xor U20946 (N_20946,N_19061,N_19108);
and U20947 (N_20947,N_19355,N_19092);
or U20948 (N_20948,N_19235,N_17886);
and U20949 (N_20949,N_18651,N_17640);
nor U20950 (N_20950,N_17810,N_19800);
and U20951 (N_20951,N_17932,N_17909);
nor U20952 (N_20952,N_17869,N_19584);
nand U20953 (N_20953,N_17779,N_18179);
nor U20954 (N_20954,N_19516,N_19168);
xnor U20955 (N_20955,N_19248,N_17520);
and U20956 (N_20956,N_19352,N_19368);
and U20957 (N_20957,N_18803,N_18333);
nor U20958 (N_20958,N_17846,N_18039);
and U20959 (N_20959,N_19284,N_18948);
or U20960 (N_20960,N_17711,N_18678);
nand U20961 (N_20961,N_19034,N_18289);
nor U20962 (N_20962,N_18099,N_17848);
and U20963 (N_20963,N_19015,N_19423);
nand U20964 (N_20964,N_17924,N_17556);
nand U20965 (N_20965,N_19803,N_19293);
nor U20966 (N_20966,N_18991,N_18746);
and U20967 (N_20967,N_19577,N_19144);
and U20968 (N_20968,N_19916,N_18041);
nand U20969 (N_20969,N_19542,N_19976);
nand U20970 (N_20970,N_18631,N_18921);
and U20971 (N_20971,N_18040,N_18037);
or U20972 (N_20972,N_18707,N_18334);
or U20973 (N_20973,N_19446,N_18162);
nand U20974 (N_20974,N_18183,N_19671);
xnor U20975 (N_20975,N_17814,N_19951);
nand U20976 (N_20976,N_18460,N_19915);
and U20977 (N_20977,N_17704,N_19914);
and U20978 (N_20978,N_18351,N_18692);
xnor U20979 (N_20979,N_19199,N_18840);
nand U20980 (N_20980,N_18722,N_17663);
xnor U20981 (N_20981,N_19638,N_19252);
nand U20982 (N_20982,N_18229,N_19461);
nand U20983 (N_20983,N_18774,N_19074);
nand U20984 (N_20984,N_19366,N_18300);
nor U20985 (N_20985,N_18206,N_18133);
nand U20986 (N_20986,N_18712,N_19950);
or U20987 (N_20987,N_19651,N_18539);
xor U20988 (N_20988,N_17864,N_19021);
and U20989 (N_20989,N_17795,N_18995);
xnor U20990 (N_20990,N_18440,N_19639);
or U20991 (N_20991,N_19844,N_17793);
nor U20992 (N_20992,N_19960,N_17573);
nor U20993 (N_20993,N_19540,N_18985);
and U20994 (N_20994,N_18615,N_19088);
and U20995 (N_20995,N_19083,N_19873);
nor U20996 (N_20996,N_18152,N_19211);
nand U20997 (N_20997,N_19292,N_17522);
nand U20998 (N_20998,N_19769,N_19492);
nand U20999 (N_20999,N_19233,N_19068);
nand U21000 (N_21000,N_18665,N_19376);
xor U21001 (N_21001,N_18846,N_19918);
nor U21002 (N_21002,N_18632,N_17993);
xnor U21003 (N_21003,N_18989,N_19191);
xor U21004 (N_21004,N_17678,N_18444);
or U21005 (N_21005,N_19031,N_18564);
nor U21006 (N_21006,N_19282,N_18820);
nor U21007 (N_21007,N_17523,N_19479);
and U21008 (N_21008,N_18027,N_19809);
nor U21009 (N_21009,N_19834,N_19219);
and U21010 (N_21010,N_18646,N_18594);
and U21011 (N_21011,N_18537,N_19903);
and U21012 (N_21012,N_19272,N_19595);
or U21013 (N_21013,N_19874,N_19278);
or U21014 (N_21014,N_17651,N_18603);
nand U21015 (N_21015,N_19157,N_17826);
nand U21016 (N_21016,N_18714,N_19818);
nand U21017 (N_21017,N_19845,N_18685);
or U21018 (N_21018,N_18616,N_18397);
nor U21019 (N_21019,N_17649,N_19953);
xnor U21020 (N_21020,N_19524,N_17789);
nor U21021 (N_21021,N_18139,N_19949);
nor U21022 (N_21022,N_17984,N_19862);
and U21023 (N_21023,N_19378,N_19189);
xor U21024 (N_21024,N_17956,N_18926);
xnor U21025 (N_21025,N_17966,N_19973);
nand U21026 (N_21026,N_19433,N_18443);
or U21027 (N_21027,N_19217,N_19448);
or U21028 (N_21028,N_18555,N_17903);
and U21029 (N_21029,N_19726,N_18034);
and U21030 (N_21030,N_19854,N_18503);
or U21031 (N_21031,N_18181,N_19798);
nand U21032 (N_21032,N_19215,N_18662);
nand U21033 (N_21033,N_19952,N_17805);
nor U21034 (N_21034,N_19437,N_17772);
or U21035 (N_21035,N_19534,N_18008);
or U21036 (N_21036,N_19365,N_19911);
and U21037 (N_21037,N_18343,N_18413);
and U21038 (N_21038,N_18761,N_18166);
xnor U21039 (N_21039,N_18311,N_19385);
nand U21040 (N_21040,N_19414,N_17753);
and U21041 (N_21041,N_19986,N_17515);
nand U21042 (N_21042,N_19668,N_17560);
and U21043 (N_21043,N_17557,N_18700);
nor U21044 (N_21044,N_19091,N_17606);
or U21045 (N_21045,N_18065,N_18837);
nand U21046 (N_21046,N_18412,N_18822);
or U21047 (N_21047,N_19232,N_18618);
xor U21048 (N_21048,N_18750,N_19273);
or U21049 (N_21049,N_17890,N_19743);
xor U21050 (N_21050,N_19169,N_18765);
and U21051 (N_21051,N_17792,N_19125);
xnor U21052 (N_21052,N_18711,N_18657);
or U21053 (N_21053,N_19992,N_19781);
nand U21054 (N_21054,N_18963,N_18748);
xor U21055 (N_21055,N_18550,N_19504);
and U21056 (N_21056,N_19142,N_18868);
xor U21057 (N_21057,N_19680,N_18492);
nor U21058 (N_21058,N_18938,N_18404);
nor U21059 (N_21059,N_19130,N_17647);
nand U21060 (N_21060,N_19655,N_19040);
or U21061 (N_21061,N_18212,N_18167);
xnor U21062 (N_21062,N_18838,N_19603);
and U21063 (N_21063,N_18839,N_18507);
and U21064 (N_21064,N_18914,N_19732);
and U21065 (N_21065,N_17705,N_17988);
and U21066 (N_21066,N_18525,N_19677);
or U21067 (N_21067,N_17600,N_17740);
nand U21068 (N_21068,N_18469,N_18357);
and U21069 (N_21069,N_19201,N_17865);
xor U21070 (N_21070,N_18283,N_19511);
and U21071 (N_21071,N_19865,N_19429);
or U21072 (N_21072,N_18752,N_18480);
xnor U21073 (N_21073,N_18032,N_19857);
or U21074 (N_21074,N_18187,N_18634);
xor U21075 (N_21075,N_18773,N_19464);
or U21076 (N_21076,N_18194,N_17816);
and U21077 (N_21077,N_17603,N_19825);
nand U21078 (N_21078,N_17915,N_19560);
or U21079 (N_21079,N_18579,N_19947);
nor U21080 (N_21080,N_17882,N_18012);
and U21081 (N_21081,N_17726,N_19837);
and U21082 (N_21082,N_17648,N_18855);
and U21083 (N_21083,N_18292,N_18823);
xor U21084 (N_21084,N_18566,N_18721);
and U21085 (N_21085,N_19008,N_18103);
nor U21086 (N_21086,N_19717,N_17729);
and U21087 (N_21087,N_19785,N_19192);
nor U21088 (N_21088,N_19012,N_18171);
nand U21089 (N_21089,N_18544,N_17827);
nor U21090 (N_21090,N_18377,N_19350);
nand U21091 (N_21091,N_19481,N_19410);
xor U21092 (N_21092,N_18220,N_18248);
and U21093 (N_21093,N_17806,N_19972);
nor U21094 (N_21094,N_17615,N_18533);
nand U21095 (N_21095,N_19030,N_18383);
xnor U21096 (N_21096,N_17976,N_17880);
xnor U21097 (N_21097,N_18570,N_18847);
nand U21098 (N_21098,N_18433,N_19653);
nand U21099 (N_21099,N_17900,N_19633);
and U21100 (N_21100,N_19864,N_17769);
nand U21101 (N_21101,N_18701,N_19489);
or U21102 (N_21102,N_19975,N_18695);
nand U21103 (N_21103,N_18366,N_18758);
and U21104 (N_21104,N_18754,N_17943);
or U21105 (N_21105,N_18348,N_19247);
nand U21106 (N_21106,N_18127,N_18073);
nand U21107 (N_21107,N_19920,N_18747);
and U21108 (N_21108,N_19846,N_19011);
nor U21109 (N_21109,N_17685,N_17919);
nor U21110 (N_21110,N_18114,N_18156);
and U21111 (N_21111,N_17952,N_19204);
nand U21112 (N_21112,N_18005,N_19373);
xnor U21113 (N_21113,N_19156,N_19026);
nand U21114 (N_21114,N_18031,N_17528);
xor U21115 (N_21115,N_19261,N_19853);
nor U21116 (N_21116,N_18325,N_18659);
and U21117 (N_21117,N_18999,N_18886);
and U21118 (N_21118,N_17728,N_18510);
or U21119 (N_21119,N_18704,N_18168);
xnor U21120 (N_21120,N_18553,N_18806);
nor U21121 (N_21121,N_18486,N_18905);
or U21122 (N_21122,N_18532,N_17996);
nor U21123 (N_21123,N_18786,N_18621);
and U21124 (N_21124,N_19059,N_19367);
nand U21125 (N_21125,N_19436,N_19206);
nand U21126 (N_21126,N_17699,N_18587);
nand U21127 (N_21127,N_18268,N_19117);
and U21128 (N_21128,N_18387,N_18417);
nand U21129 (N_21129,N_19314,N_19799);
xor U21130 (N_21130,N_17937,N_18263);
xnor U21131 (N_21131,N_17735,N_17893);
nor U21132 (N_21132,N_18728,N_19228);
or U21133 (N_21133,N_19851,N_17948);
or U21134 (N_21134,N_19586,N_19902);
nor U21135 (N_21135,N_17571,N_18374);
nand U21136 (N_21136,N_19630,N_18842);
and U21137 (N_21137,N_18066,N_18003);
xnor U21138 (N_21138,N_18287,N_19901);
xnor U21139 (N_21139,N_17788,N_18294);
nand U21140 (N_21140,N_19349,N_19214);
and U21141 (N_21141,N_19643,N_17669);
or U21142 (N_21142,N_19810,N_19419);
nand U21143 (N_21143,N_18522,N_18332);
or U21144 (N_21144,N_17927,N_18134);
and U21145 (N_21145,N_19311,N_19954);
and U21146 (N_21146,N_18637,N_17621);
xnor U21147 (N_21147,N_19285,N_19110);
and U21148 (N_21148,N_19505,N_19723);
xnor U21149 (N_21149,N_19006,N_17696);
or U21150 (N_21150,N_19418,N_18960);
or U21151 (N_21151,N_18912,N_17610);
nand U21152 (N_21152,N_17985,N_17525);
nor U21153 (N_21153,N_19941,N_17951);
and U21154 (N_21154,N_17908,N_19896);
or U21155 (N_21155,N_18408,N_17568);
xnor U21156 (N_21156,N_18064,N_18256);
and U21157 (N_21157,N_17609,N_17734);
or U21158 (N_21158,N_19667,N_18771);
and U21159 (N_21159,N_19409,N_18856);
xor U21160 (N_21160,N_17555,N_19842);
and U21161 (N_21161,N_19487,N_18915);
xnor U21162 (N_21162,N_19440,N_17546);
or U21163 (N_21163,N_18600,N_19594);
nor U21164 (N_21164,N_19050,N_18862);
nor U21165 (N_21165,N_19164,N_18883);
and U21166 (N_21166,N_19444,N_19665);
xor U21167 (N_21167,N_19664,N_18319);
and U21168 (N_21168,N_19569,N_18836);
nor U21169 (N_21169,N_19208,N_17661);
nand U21170 (N_21170,N_18894,N_18128);
and U21171 (N_21171,N_17987,N_18137);
xnor U21172 (N_21172,N_18874,N_17713);
and U21173 (N_21173,N_18329,N_17631);
or U21174 (N_21174,N_18825,N_17676);
nand U21175 (N_21175,N_17851,N_17935);
nand U21176 (N_21176,N_17593,N_19486);
nor U21177 (N_21177,N_17833,N_18441);
nand U21178 (N_21178,N_19587,N_18986);
nor U21179 (N_21179,N_19287,N_19672);
nand U21180 (N_21180,N_18018,N_18971);
nand U21181 (N_21181,N_19679,N_19626);
nor U21182 (N_21182,N_18435,N_18232);
nor U21183 (N_21183,N_18880,N_17872);
nand U21184 (N_21184,N_17597,N_18052);
or U21185 (N_21185,N_17760,N_18702);
nand U21186 (N_21186,N_18756,N_18483);
nand U21187 (N_21187,N_18098,N_19326);
and U21188 (N_21188,N_19792,N_19268);
or U21189 (N_21189,N_17695,N_19981);
or U21190 (N_21190,N_18424,N_19937);
and U21191 (N_21191,N_19780,N_18577);
and U21192 (N_21192,N_19332,N_19060);
nand U21193 (N_21193,N_19266,N_19636);
xnor U21194 (N_21194,N_19389,N_18626);
xnor U21195 (N_21195,N_18226,N_19910);
xnor U21196 (N_21196,N_18056,N_18523);
or U21197 (N_21197,N_19561,N_18813);
or U21198 (N_21198,N_17642,N_19964);
or U21199 (N_21199,N_19928,N_18869);
or U21200 (N_21200,N_18610,N_18627);
or U21201 (N_21201,N_19161,N_19066);
and U21202 (N_21202,N_19177,N_17549);
nand U21203 (N_21203,N_17922,N_18455);
nor U21204 (N_21204,N_18817,N_18476);
nor U21205 (N_21205,N_18739,N_18549);
and U21206 (N_21206,N_18740,N_18261);
xnor U21207 (N_21207,N_19859,N_18807);
or U21208 (N_21208,N_18502,N_19749);
and U21209 (N_21209,N_17749,N_18772);
xnor U21210 (N_21210,N_18802,N_18352);
nand U21211 (N_21211,N_19490,N_19530);
xor U21212 (N_21212,N_17881,N_19805);
nand U21213 (N_21213,N_18330,N_19137);
xnor U21214 (N_21214,N_19223,N_19787);
nand U21215 (N_21215,N_18904,N_17588);
and U21216 (N_21216,N_19435,N_19330);
and U21217 (N_21217,N_18392,N_18939);
nor U21218 (N_21218,N_19165,N_18819);
or U21219 (N_21219,N_19823,N_19226);
xnor U21220 (N_21220,N_18022,N_18215);
and U21221 (N_21221,N_19162,N_19539);
xor U21222 (N_21222,N_17739,N_18104);
and U21223 (N_21223,N_18489,N_18189);
or U21224 (N_21224,N_18643,N_18159);
or U21225 (N_21225,N_17628,N_18961);
nor U21226 (N_21226,N_17854,N_17714);
nand U21227 (N_21227,N_19073,N_18328);
and U21228 (N_21228,N_18974,N_19398);
nor U21229 (N_21229,N_18811,N_17507);
or U21230 (N_21230,N_19808,N_18178);
or U21231 (N_21231,N_18385,N_17998);
nand U21232 (N_21232,N_17529,N_17957);
and U21233 (N_21233,N_19238,N_18112);
nand U21234 (N_21234,N_18789,N_17917);
nor U21235 (N_21235,N_18755,N_19555);
xor U21236 (N_21236,N_19475,N_19476);
nor U21237 (N_21237,N_19881,N_18679);
or U21238 (N_21238,N_19455,N_17641);
nand U21239 (N_21239,N_18852,N_17804);
nand U21240 (N_21240,N_17514,N_18574);
and U21241 (N_21241,N_17559,N_18060);
nor U21242 (N_21242,N_18513,N_18569);
nand U21243 (N_21243,N_18327,N_18284);
nor U21244 (N_21244,N_19751,N_19107);
or U21245 (N_21245,N_18396,N_19027);
and U21246 (N_21246,N_19623,N_19817);
or U21247 (N_21247,N_18715,N_19713);
nand U21248 (N_21248,N_19795,N_19071);
xnor U21249 (N_21249,N_18576,N_19627);
nor U21250 (N_21250,N_18283,N_18895);
nor U21251 (N_21251,N_18006,N_17550);
or U21252 (N_21252,N_19489,N_19063);
nand U21253 (N_21253,N_18495,N_18857);
and U21254 (N_21254,N_18343,N_17878);
or U21255 (N_21255,N_18621,N_19117);
or U21256 (N_21256,N_17725,N_18304);
or U21257 (N_21257,N_19522,N_18062);
nand U21258 (N_21258,N_18630,N_17705);
or U21259 (N_21259,N_17718,N_18159);
and U21260 (N_21260,N_19768,N_17973);
nand U21261 (N_21261,N_18187,N_18997);
or U21262 (N_21262,N_18973,N_17906);
nand U21263 (N_21263,N_18656,N_19970);
and U21264 (N_21264,N_19634,N_18446);
nand U21265 (N_21265,N_18683,N_18318);
or U21266 (N_21266,N_19891,N_18881);
and U21267 (N_21267,N_18800,N_18409);
nand U21268 (N_21268,N_18996,N_19236);
and U21269 (N_21269,N_19042,N_19611);
or U21270 (N_21270,N_19824,N_19251);
nand U21271 (N_21271,N_18565,N_17686);
xnor U21272 (N_21272,N_19553,N_17683);
nor U21273 (N_21273,N_19441,N_18849);
or U21274 (N_21274,N_18063,N_19980);
nand U21275 (N_21275,N_18161,N_18208);
and U21276 (N_21276,N_18752,N_19802);
nand U21277 (N_21277,N_18458,N_17619);
nor U21278 (N_21278,N_19086,N_19907);
and U21279 (N_21279,N_19833,N_19249);
nor U21280 (N_21280,N_18374,N_19359);
or U21281 (N_21281,N_19077,N_18143);
xnor U21282 (N_21282,N_18117,N_19326);
or U21283 (N_21283,N_17697,N_19488);
and U21284 (N_21284,N_17776,N_19059);
and U21285 (N_21285,N_19280,N_19773);
and U21286 (N_21286,N_18383,N_19437);
nor U21287 (N_21287,N_18864,N_17962);
nor U21288 (N_21288,N_18772,N_17773);
nor U21289 (N_21289,N_19382,N_18575);
xnor U21290 (N_21290,N_17982,N_18526);
nand U21291 (N_21291,N_19596,N_18312);
and U21292 (N_21292,N_19183,N_17851);
xnor U21293 (N_21293,N_19894,N_19793);
nor U21294 (N_21294,N_18633,N_19049);
nand U21295 (N_21295,N_19415,N_19739);
xor U21296 (N_21296,N_17964,N_17547);
xor U21297 (N_21297,N_18305,N_18680);
and U21298 (N_21298,N_17766,N_17799);
xor U21299 (N_21299,N_17552,N_17612);
or U21300 (N_21300,N_17894,N_19695);
nand U21301 (N_21301,N_18988,N_19465);
and U21302 (N_21302,N_19510,N_19994);
xor U21303 (N_21303,N_18418,N_19265);
or U21304 (N_21304,N_19408,N_19142);
nand U21305 (N_21305,N_19732,N_19165);
nand U21306 (N_21306,N_19935,N_18836);
xor U21307 (N_21307,N_19027,N_19009);
or U21308 (N_21308,N_19933,N_17717);
and U21309 (N_21309,N_18687,N_18590);
nand U21310 (N_21310,N_19540,N_18458);
nor U21311 (N_21311,N_18492,N_17756);
xnor U21312 (N_21312,N_19825,N_18336);
nand U21313 (N_21313,N_18438,N_19383);
and U21314 (N_21314,N_18751,N_19647);
and U21315 (N_21315,N_18632,N_18514);
and U21316 (N_21316,N_19752,N_19984);
and U21317 (N_21317,N_19006,N_19255);
or U21318 (N_21318,N_18924,N_19832);
xor U21319 (N_21319,N_18543,N_17675);
xnor U21320 (N_21320,N_19606,N_19584);
or U21321 (N_21321,N_18192,N_18773);
or U21322 (N_21322,N_19324,N_18337);
or U21323 (N_21323,N_18332,N_19276);
nand U21324 (N_21324,N_18738,N_18847);
or U21325 (N_21325,N_19181,N_19685);
xnor U21326 (N_21326,N_19720,N_17937);
and U21327 (N_21327,N_17902,N_19053);
and U21328 (N_21328,N_19414,N_18795);
xnor U21329 (N_21329,N_19323,N_17596);
nand U21330 (N_21330,N_18755,N_17760);
xor U21331 (N_21331,N_19103,N_19996);
and U21332 (N_21332,N_17922,N_18256);
and U21333 (N_21333,N_17925,N_19859);
or U21334 (N_21334,N_18411,N_19859);
nand U21335 (N_21335,N_18622,N_17678);
and U21336 (N_21336,N_18055,N_17835);
and U21337 (N_21337,N_18463,N_19277);
nor U21338 (N_21338,N_19746,N_18863);
and U21339 (N_21339,N_19691,N_19696);
xnor U21340 (N_21340,N_19976,N_17514);
nor U21341 (N_21341,N_17641,N_19972);
nor U21342 (N_21342,N_18949,N_18552);
or U21343 (N_21343,N_18503,N_17823);
xnor U21344 (N_21344,N_19237,N_17851);
or U21345 (N_21345,N_18031,N_19767);
nand U21346 (N_21346,N_18731,N_17926);
nand U21347 (N_21347,N_17914,N_18671);
nor U21348 (N_21348,N_18915,N_18561);
and U21349 (N_21349,N_19299,N_19464);
nor U21350 (N_21350,N_18540,N_18684);
xor U21351 (N_21351,N_17534,N_19853);
and U21352 (N_21352,N_17731,N_17988);
or U21353 (N_21353,N_17762,N_17816);
or U21354 (N_21354,N_19308,N_19402);
and U21355 (N_21355,N_19708,N_19256);
xnor U21356 (N_21356,N_19325,N_19280);
and U21357 (N_21357,N_18252,N_19112);
and U21358 (N_21358,N_18464,N_17789);
nor U21359 (N_21359,N_18384,N_18303);
xnor U21360 (N_21360,N_18242,N_18421);
nor U21361 (N_21361,N_18278,N_17639);
and U21362 (N_21362,N_18123,N_18907);
and U21363 (N_21363,N_18144,N_19224);
nor U21364 (N_21364,N_19865,N_17519);
nor U21365 (N_21365,N_18438,N_19793);
nand U21366 (N_21366,N_17576,N_18494);
xor U21367 (N_21367,N_17832,N_18525);
and U21368 (N_21368,N_17876,N_17829);
nor U21369 (N_21369,N_18296,N_19330);
and U21370 (N_21370,N_18303,N_19188);
nand U21371 (N_21371,N_19334,N_19205);
xor U21372 (N_21372,N_19411,N_18110);
nand U21373 (N_21373,N_19427,N_17984);
nand U21374 (N_21374,N_17541,N_17921);
and U21375 (N_21375,N_19278,N_17776);
xor U21376 (N_21376,N_18077,N_19003);
xnor U21377 (N_21377,N_17907,N_19393);
nand U21378 (N_21378,N_18239,N_18689);
nand U21379 (N_21379,N_17662,N_18231);
and U21380 (N_21380,N_18543,N_19916);
xor U21381 (N_21381,N_19693,N_18274);
xor U21382 (N_21382,N_19053,N_18204);
nor U21383 (N_21383,N_18873,N_18609);
and U21384 (N_21384,N_17664,N_18982);
nand U21385 (N_21385,N_18408,N_19721);
and U21386 (N_21386,N_18300,N_19974);
nand U21387 (N_21387,N_18498,N_17577);
nor U21388 (N_21388,N_19896,N_18285);
xnor U21389 (N_21389,N_19198,N_19333);
and U21390 (N_21390,N_19192,N_19866);
or U21391 (N_21391,N_19199,N_19067);
nand U21392 (N_21392,N_18479,N_17902);
xor U21393 (N_21393,N_18181,N_18941);
nand U21394 (N_21394,N_17597,N_19437);
xnor U21395 (N_21395,N_19435,N_19847);
nor U21396 (N_21396,N_19154,N_19790);
nand U21397 (N_21397,N_19520,N_17691);
nor U21398 (N_21398,N_19626,N_19147);
or U21399 (N_21399,N_19746,N_19325);
or U21400 (N_21400,N_18290,N_19398);
xnor U21401 (N_21401,N_18268,N_17705);
nand U21402 (N_21402,N_18109,N_18574);
xnor U21403 (N_21403,N_17978,N_19988);
xor U21404 (N_21404,N_18602,N_18943);
and U21405 (N_21405,N_18143,N_18048);
or U21406 (N_21406,N_17589,N_19260);
nand U21407 (N_21407,N_17809,N_17621);
nand U21408 (N_21408,N_19983,N_17689);
or U21409 (N_21409,N_19493,N_18772);
or U21410 (N_21410,N_17757,N_18303);
nor U21411 (N_21411,N_17580,N_19539);
nor U21412 (N_21412,N_19978,N_19086);
or U21413 (N_21413,N_17677,N_19102);
nand U21414 (N_21414,N_19738,N_19532);
and U21415 (N_21415,N_18077,N_19611);
nor U21416 (N_21416,N_19243,N_19297);
xnor U21417 (N_21417,N_17533,N_19684);
xnor U21418 (N_21418,N_18854,N_18772);
and U21419 (N_21419,N_19574,N_19316);
or U21420 (N_21420,N_19868,N_18366);
or U21421 (N_21421,N_19462,N_18281);
and U21422 (N_21422,N_18733,N_17730);
nor U21423 (N_21423,N_18605,N_19872);
nor U21424 (N_21424,N_18937,N_17595);
nand U21425 (N_21425,N_18690,N_17915);
xor U21426 (N_21426,N_19256,N_19439);
or U21427 (N_21427,N_19769,N_18859);
or U21428 (N_21428,N_18603,N_18070);
nor U21429 (N_21429,N_17888,N_19527);
and U21430 (N_21430,N_19163,N_19475);
and U21431 (N_21431,N_19816,N_17561);
nand U21432 (N_21432,N_19950,N_18761);
nand U21433 (N_21433,N_18338,N_17542);
or U21434 (N_21434,N_18566,N_19040);
or U21435 (N_21435,N_19345,N_18093);
or U21436 (N_21436,N_19759,N_19640);
or U21437 (N_21437,N_19912,N_19400);
xor U21438 (N_21438,N_19037,N_19181);
and U21439 (N_21439,N_19776,N_18653);
or U21440 (N_21440,N_18300,N_19819);
and U21441 (N_21441,N_18718,N_19574);
or U21442 (N_21442,N_19402,N_18090);
and U21443 (N_21443,N_18705,N_17503);
xor U21444 (N_21444,N_19225,N_19429);
xnor U21445 (N_21445,N_19357,N_17579);
or U21446 (N_21446,N_19909,N_19792);
xnor U21447 (N_21447,N_17653,N_18162);
nand U21448 (N_21448,N_18314,N_17965);
and U21449 (N_21449,N_18540,N_17997);
nor U21450 (N_21450,N_17789,N_19985);
nor U21451 (N_21451,N_19218,N_18875);
nand U21452 (N_21452,N_18007,N_17832);
nor U21453 (N_21453,N_18567,N_18793);
xnor U21454 (N_21454,N_19243,N_19683);
nor U21455 (N_21455,N_19000,N_19286);
nor U21456 (N_21456,N_18890,N_17715);
nor U21457 (N_21457,N_19479,N_17565);
nand U21458 (N_21458,N_19422,N_17876);
and U21459 (N_21459,N_19439,N_18961);
and U21460 (N_21460,N_18215,N_17741);
and U21461 (N_21461,N_18979,N_17822);
xnor U21462 (N_21462,N_17985,N_17543);
or U21463 (N_21463,N_19707,N_18567);
or U21464 (N_21464,N_17854,N_18554);
or U21465 (N_21465,N_18887,N_19121);
or U21466 (N_21466,N_19417,N_17911);
and U21467 (N_21467,N_19017,N_19908);
nand U21468 (N_21468,N_19536,N_17652);
or U21469 (N_21469,N_18346,N_18870);
nand U21470 (N_21470,N_19298,N_19626);
nand U21471 (N_21471,N_19906,N_19411);
xnor U21472 (N_21472,N_18499,N_17718);
and U21473 (N_21473,N_18683,N_19226);
nor U21474 (N_21474,N_19692,N_17912);
and U21475 (N_21475,N_19382,N_19973);
or U21476 (N_21476,N_17707,N_19587);
and U21477 (N_21477,N_19602,N_18686);
xor U21478 (N_21478,N_18058,N_17656);
or U21479 (N_21479,N_19656,N_18709);
nor U21480 (N_21480,N_18982,N_18341);
or U21481 (N_21481,N_18900,N_18115);
and U21482 (N_21482,N_19952,N_17670);
xnor U21483 (N_21483,N_19897,N_19582);
nor U21484 (N_21484,N_18566,N_19411);
or U21485 (N_21485,N_18686,N_19556);
nor U21486 (N_21486,N_17587,N_19189);
and U21487 (N_21487,N_19616,N_19871);
and U21488 (N_21488,N_17928,N_18112);
nor U21489 (N_21489,N_19282,N_17506);
nor U21490 (N_21490,N_19181,N_17889);
and U21491 (N_21491,N_17678,N_18180);
nand U21492 (N_21492,N_19362,N_18529);
nor U21493 (N_21493,N_19259,N_19608);
xor U21494 (N_21494,N_19535,N_17722);
nand U21495 (N_21495,N_18656,N_18032);
nor U21496 (N_21496,N_19773,N_17839);
nor U21497 (N_21497,N_19225,N_17511);
xor U21498 (N_21498,N_19752,N_18368);
xnor U21499 (N_21499,N_18069,N_17756);
xnor U21500 (N_21500,N_18542,N_18086);
and U21501 (N_21501,N_19969,N_18017);
nand U21502 (N_21502,N_18043,N_19527);
and U21503 (N_21503,N_19866,N_19579);
xnor U21504 (N_21504,N_19376,N_19844);
nor U21505 (N_21505,N_18312,N_19829);
and U21506 (N_21506,N_19397,N_18150);
nor U21507 (N_21507,N_17544,N_17944);
and U21508 (N_21508,N_19126,N_19932);
and U21509 (N_21509,N_18187,N_19249);
xor U21510 (N_21510,N_17606,N_18095);
and U21511 (N_21511,N_18040,N_17832);
xor U21512 (N_21512,N_19366,N_17851);
xnor U21513 (N_21513,N_19315,N_19084);
xnor U21514 (N_21514,N_18153,N_19327);
or U21515 (N_21515,N_18764,N_17899);
nor U21516 (N_21516,N_19851,N_17619);
nor U21517 (N_21517,N_19792,N_19196);
nand U21518 (N_21518,N_18964,N_18498);
xnor U21519 (N_21519,N_18275,N_17579);
nand U21520 (N_21520,N_18971,N_18178);
and U21521 (N_21521,N_19157,N_17846);
nand U21522 (N_21522,N_19597,N_17564);
and U21523 (N_21523,N_18639,N_18817);
nand U21524 (N_21524,N_17987,N_17724);
nand U21525 (N_21525,N_18948,N_18156);
nand U21526 (N_21526,N_18852,N_17645);
or U21527 (N_21527,N_18172,N_18830);
or U21528 (N_21528,N_17878,N_19969);
and U21529 (N_21529,N_18478,N_18513);
or U21530 (N_21530,N_17692,N_17602);
and U21531 (N_21531,N_18544,N_19733);
and U21532 (N_21532,N_18214,N_17542);
xnor U21533 (N_21533,N_19713,N_19169);
xnor U21534 (N_21534,N_18891,N_18304);
xor U21535 (N_21535,N_19543,N_18900);
nor U21536 (N_21536,N_18899,N_19620);
or U21537 (N_21537,N_19987,N_18802);
xnor U21538 (N_21538,N_19961,N_17561);
nor U21539 (N_21539,N_19962,N_18838);
nor U21540 (N_21540,N_17519,N_18786);
and U21541 (N_21541,N_18021,N_18965);
xnor U21542 (N_21542,N_18911,N_17942);
nor U21543 (N_21543,N_17677,N_19415);
and U21544 (N_21544,N_18031,N_19248);
and U21545 (N_21545,N_19458,N_18290);
nor U21546 (N_21546,N_18259,N_17665);
or U21547 (N_21547,N_17785,N_19185);
or U21548 (N_21548,N_18669,N_17522);
or U21549 (N_21549,N_18577,N_19898);
nor U21550 (N_21550,N_18569,N_17736);
nand U21551 (N_21551,N_18208,N_17926);
or U21552 (N_21552,N_19510,N_17748);
or U21553 (N_21553,N_18830,N_17548);
and U21554 (N_21554,N_18284,N_17912);
nand U21555 (N_21555,N_19403,N_18212);
xor U21556 (N_21556,N_18835,N_17707);
nand U21557 (N_21557,N_18564,N_18257);
nor U21558 (N_21558,N_18320,N_18249);
nand U21559 (N_21559,N_19904,N_19725);
xnor U21560 (N_21560,N_18328,N_18492);
and U21561 (N_21561,N_17580,N_18585);
nand U21562 (N_21562,N_19615,N_19449);
nor U21563 (N_21563,N_17550,N_18504);
xnor U21564 (N_21564,N_19538,N_17638);
nor U21565 (N_21565,N_17638,N_18166);
xnor U21566 (N_21566,N_18602,N_19110);
and U21567 (N_21567,N_19503,N_19935);
and U21568 (N_21568,N_19227,N_18181);
xnor U21569 (N_21569,N_18551,N_17661);
or U21570 (N_21570,N_17890,N_18567);
and U21571 (N_21571,N_19481,N_17918);
or U21572 (N_21572,N_18490,N_19453);
xor U21573 (N_21573,N_19961,N_18335);
xnor U21574 (N_21574,N_17948,N_19625);
nor U21575 (N_21575,N_18947,N_18681);
xnor U21576 (N_21576,N_19958,N_19765);
xnor U21577 (N_21577,N_18234,N_18610);
nor U21578 (N_21578,N_18887,N_18449);
nand U21579 (N_21579,N_18037,N_19114);
and U21580 (N_21580,N_18494,N_19518);
nand U21581 (N_21581,N_18751,N_19765);
or U21582 (N_21582,N_18706,N_18349);
or U21583 (N_21583,N_18177,N_18361);
and U21584 (N_21584,N_18027,N_18057);
xor U21585 (N_21585,N_19627,N_19069);
or U21586 (N_21586,N_18517,N_19068);
xor U21587 (N_21587,N_19928,N_19175);
and U21588 (N_21588,N_19628,N_18793);
nand U21589 (N_21589,N_19369,N_19052);
xnor U21590 (N_21590,N_19838,N_19114);
nor U21591 (N_21591,N_18147,N_19219);
or U21592 (N_21592,N_18343,N_18840);
nand U21593 (N_21593,N_19032,N_19609);
or U21594 (N_21594,N_18152,N_18810);
nor U21595 (N_21595,N_19280,N_19924);
or U21596 (N_21596,N_19618,N_18182);
and U21597 (N_21597,N_18705,N_18267);
nand U21598 (N_21598,N_19976,N_19709);
nand U21599 (N_21599,N_17802,N_18281);
xor U21600 (N_21600,N_19683,N_19066);
nand U21601 (N_21601,N_17997,N_19165);
or U21602 (N_21602,N_19116,N_18510);
nand U21603 (N_21603,N_19349,N_18839);
or U21604 (N_21604,N_19357,N_18446);
or U21605 (N_21605,N_18595,N_19904);
nand U21606 (N_21606,N_19808,N_19935);
nor U21607 (N_21607,N_18814,N_19832);
and U21608 (N_21608,N_18716,N_19579);
xnor U21609 (N_21609,N_17952,N_19334);
nand U21610 (N_21610,N_18346,N_17801);
xor U21611 (N_21611,N_19501,N_18962);
nor U21612 (N_21612,N_19050,N_18244);
nor U21613 (N_21613,N_18120,N_19116);
xor U21614 (N_21614,N_18855,N_17501);
nand U21615 (N_21615,N_18427,N_19440);
nand U21616 (N_21616,N_18487,N_19940);
xor U21617 (N_21617,N_19487,N_18059);
nor U21618 (N_21618,N_18028,N_19925);
and U21619 (N_21619,N_19606,N_17806);
xor U21620 (N_21620,N_19697,N_17936);
nor U21621 (N_21621,N_18174,N_19344);
nand U21622 (N_21622,N_17956,N_19778);
nand U21623 (N_21623,N_18286,N_19058);
nor U21624 (N_21624,N_19623,N_18820);
nand U21625 (N_21625,N_18238,N_17869);
or U21626 (N_21626,N_18669,N_18133);
and U21627 (N_21627,N_18981,N_17948);
or U21628 (N_21628,N_19484,N_19319);
nand U21629 (N_21629,N_17785,N_19417);
or U21630 (N_21630,N_18768,N_19675);
and U21631 (N_21631,N_17827,N_17596);
xnor U21632 (N_21632,N_18917,N_19113);
and U21633 (N_21633,N_17738,N_18000);
nand U21634 (N_21634,N_17503,N_18806);
xnor U21635 (N_21635,N_19321,N_19016);
and U21636 (N_21636,N_18959,N_18544);
xor U21637 (N_21637,N_19783,N_19355);
xor U21638 (N_21638,N_17509,N_17539);
nor U21639 (N_21639,N_19970,N_19369);
and U21640 (N_21640,N_17524,N_17761);
nand U21641 (N_21641,N_19760,N_18111);
or U21642 (N_21642,N_18988,N_17818);
nor U21643 (N_21643,N_19200,N_19772);
and U21644 (N_21644,N_19539,N_19854);
and U21645 (N_21645,N_19052,N_18110);
xnor U21646 (N_21646,N_18503,N_19744);
xnor U21647 (N_21647,N_18370,N_18508);
or U21648 (N_21648,N_17575,N_18388);
and U21649 (N_21649,N_18055,N_18537);
or U21650 (N_21650,N_17683,N_19172);
nand U21651 (N_21651,N_17830,N_18927);
xnor U21652 (N_21652,N_18920,N_18164);
and U21653 (N_21653,N_18276,N_18678);
and U21654 (N_21654,N_19604,N_19164);
nand U21655 (N_21655,N_19201,N_17594);
and U21656 (N_21656,N_19119,N_19408);
nor U21657 (N_21657,N_19751,N_19271);
and U21658 (N_21658,N_18341,N_18787);
xnor U21659 (N_21659,N_19262,N_19032);
xnor U21660 (N_21660,N_18884,N_19463);
and U21661 (N_21661,N_17900,N_18697);
nor U21662 (N_21662,N_17852,N_18633);
xor U21663 (N_21663,N_19752,N_19542);
or U21664 (N_21664,N_18072,N_19062);
or U21665 (N_21665,N_19464,N_18085);
and U21666 (N_21666,N_18670,N_17787);
xnor U21667 (N_21667,N_18716,N_17974);
nor U21668 (N_21668,N_19005,N_19490);
nor U21669 (N_21669,N_17850,N_19586);
nand U21670 (N_21670,N_18428,N_18616);
and U21671 (N_21671,N_19158,N_18429);
or U21672 (N_21672,N_19393,N_18761);
nand U21673 (N_21673,N_18107,N_17965);
xnor U21674 (N_21674,N_18181,N_18474);
or U21675 (N_21675,N_18282,N_18246);
nand U21676 (N_21676,N_18989,N_18618);
nor U21677 (N_21677,N_19361,N_19777);
nor U21678 (N_21678,N_18734,N_18049);
nand U21679 (N_21679,N_18428,N_18929);
or U21680 (N_21680,N_18643,N_19626);
nor U21681 (N_21681,N_18371,N_18135);
or U21682 (N_21682,N_17885,N_18551);
and U21683 (N_21683,N_17803,N_19951);
nand U21684 (N_21684,N_19895,N_17842);
and U21685 (N_21685,N_18509,N_19237);
nand U21686 (N_21686,N_18351,N_18496);
nor U21687 (N_21687,N_19769,N_17877);
xnor U21688 (N_21688,N_19101,N_19393);
xnor U21689 (N_21689,N_19939,N_18559);
xnor U21690 (N_21690,N_17930,N_18307);
xor U21691 (N_21691,N_17997,N_19475);
and U21692 (N_21692,N_18612,N_17573);
nor U21693 (N_21693,N_18372,N_19837);
nand U21694 (N_21694,N_19987,N_18108);
nand U21695 (N_21695,N_17622,N_19885);
nand U21696 (N_21696,N_18493,N_19978);
and U21697 (N_21697,N_19577,N_17853);
nand U21698 (N_21698,N_19592,N_18345);
and U21699 (N_21699,N_19444,N_19930);
nand U21700 (N_21700,N_18816,N_17711);
and U21701 (N_21701,N_19852,N_18271);
nand U21702 (N_21702,N_18341,N_17657);
nor U21703 (N_21703,N_19338,N_19784);
or U21704 (N_21704,N_18295,N_18836);
nand U21705 (N_21705,N_19470,N_17976);
and U21706 (N_21706,N_19546,N_19013);
nand U21707 (N_21707,N_18274,N_19626);
xor U21708 (N_21708,N_19953,N_19223);
xor U21709 (N_21709,N_19872,N_17844);
or U21710 (N_21710,N_18049,N_19438);
nand U21711 (N_21711,N_18714,N_19826);
and U21712 (N_21712,N_19612,N_17916);
and U21713 (N_21713,N_19686,N_17765);
and U21714 (N_21714,N_19038,N_18987);
xnor U21715 (N_21715,N_18777,N_19616);
nor U21716 (N_21716,N_18446,N_19574);
and U21717 (N_21717,N_19788,N_18421);
xnor U21718 (N_21718,N_19631,N_19576);
and U21719 (N_21719,N_18063,N_18682);
xor U21720 (N_21720,N_19676,N_18962);
nand U21721 (N_21721,N_19634,N_18708);
xnor U21722 (N_21722,N_18994,N_18410);
and U21723 (N_21723,N_19435,N_18009);
nand U21724 (N_21724,N_18884,N_19446);
nor U21725 (N_21725,N_17859,N_18421);
nand U21726 (N_21726,N_18348,N_19185);
or U21727 (N_21727,N_19800,N_18946);
and U21728 (N_21728,N_17801,N_19868);
and U21729 (N_21729,N_18612,N_19957);
nand U21730 (N_21730,N_19737,N_18872);
or U21731 (N_21731,N_18808,N_19956);
nand U21732 (N_21732,N_19666,N_19518);
xor U21733 (N_21733,N_18127,N_17746);
and U21734 (N_21734,N_18766,N_19196);
or U21735 (N_21735,N_19817,N_17521);
or U21736 (N_21736,N_19609,N_18640);
and U21737 (N_21737,N_18810,N_19599);
nor U21738 (N_21738,N_19691,N_19755);
nor U21739 (N_21739,N_18502,N_19914);
xnor U21740 (N_21740,N_19645,N_19766);
nand U21741 (N_21741,N_17523,N_19133);
and U21742 (N_21742,N_18560,N_19908);
and U21743 (N_21743,N_18331,N_19679);
or U21744 (N_21744,N_18768,N_19723);
nor U21745 (N_21745,N_19532,N_19758);
or U21746 (N_21746,N_19485,N_17927);
and U21747 (N_21747,N_19230,N_18032);
nand U21748 (N_21748,N_18421,N_18369);
nor U21749 (N_21749,N_17655,N_19701);
or U21750 (N_21750,N_17571,N_19165);
nand U21751 (N_21751,N_18587,N_17555);
or U21752 (N_21752,N_17824,N_19274);
nor U21753 (N_21753,N_18647,N_18566);
xor U21754 (N_21754,N_18384,N_19737);
xnor U21755 (N_21755,N_18157,N_19504);
or U21756 (N_21756,N_18023,N_18671);
or U21757 (N_21757,N_19295,N_18184);
xnor U21758 (N_21758,N_18418,N_19876);
nor U21759 (N_21759,N_18297,N_19590);
nand U21760 (N_21760,N_18778,N_17571);
nor U21761 (N_21761,N_18684,N_19717);
nor U21762 (N_21762,N_19926,N_18592);
nand U21763 (N_21763,N_19655,N_18339);
nor U21764 (N_21764,N_18585,N_18319);
nor U21765 (N_21765,N_18608,N_18235);
and U21766 (N_21766,N_19744,N_19913);
and U21767 (N_21767,N_17624,N_18286);
nor U21768 (N_21768,N_18632,N_19098);
and U21769 (N_21769,N_18767,N_17893);
xor U21770 (N_21770,N_17972,N_18623);
xnor U21771 (N_21771,N_19210,N_18427);
and U21772 (N_21772,N_18798,N_19863);
nand U21773 (N_21773,N_19485,N_19280);
nor U21774 (N_21774,N_18896,N_18207);
nand U21775 (N_21775,N_18741,N_18517);
and U21776 (N_21776,N_17716,N_18613);
nor U21777 (N_21777,N_18841,N_19684);
and U21778 (N_21778,N_18886,N_18522);
xnor U21779 (N_21779,N_18022,N_18635);
and U21780 (N_21780,N_19021,N_19305);
nand U21781 (N_21781,N_19397,N_19381);
nor U21782 (N_21782,N_18275,N_18204);
nor U21783 (N_21783,N_17810,N_19189);
and U21784 (N_21784,N_18067,N_19848);
or U21785 (N_21785,N_18070,N_18580);
and U21786 (N_21786,N_19266,N_18253);
nand U21787 (N_21787,N_19102,N_17753);
and U21788 (N_21788,N_19614,N_19899);
xnor U21789 (N_21789,N_19488,N_18318);
nor U21790 (N_21790,N_19866,N_18429);
or U21791 (N_21791,N_19739,N_19803);
or U21792 (N_21792,N_19963,N_18613);
and U21793 (N_21793,N_19079,N_17842);
and U21794 (N_21794,N_19670,N_18299);
nand U21795 (N_21795,N_17866,N_18956);
nand U21796 (N_21796,N_17653,N_18715);
xor U21797 (N_21797,N_18284,N_17954);
nand U21798 (N_21798,N_18912,N_17965);
nand U21799 (N_21799,N_19689,N_18971);
nand U21800 (N_21800,N_18218,N_17904);
or U21801 (N_21801,N_18446,N_19148);
or U21802 (N_21802,N_18414,N_19235);
and U21803 (N_21803,N_19018,N_18869);
and U21804 (N_21804,N_19210,N_18696);
nor U21805 (N_21805,N_19845,N_17500);
and U21806 (N_21806,N_17864,N_19953);
or U21807 (N_21807,N_18165,N_19564);
and U21808 (N_21808,N_17518,N_19586);
nand U21809 (N_21809,N_19912,N_19541);
nand U21810 (N_21810,N_18573,N_18024);
and U21811 (N_21811,N_17573,N_19557);
and U21812 (N_21812,N_19861,N_19519);
nand U21813 (N_21813,N_19652,N_19717);
xor U21814 (N_21814,N_17627,N_19718);
nor U21815 (N_21815,N_19475,N_18960);
xnor U21816 (N_21816,N_18423,N_18072);
nand U21817 (N_21817,N_19391,N_19796);
nor U21818 (N_21818,N_17545,N_18782);
xnor U21819 (N_21819,N_19859,N_17642);
and U21820 (N_21820,N_18466,N_18988);
and U21821 (N_21821,N_17758,N_19967);
nor U21822 (N_21822,N_19643,N_18274);
nor U21823 (N_21823,N_18471,N_19230);
xor U21824 (N_21824,N_17919,N_18187);
nand U21825 (N_21825,N_19103,N_18449);
or U21826 (N_21826,N_19187,N_19804);
and U21827 (N_21827,N_19685,N_19320);
nor U21828 (N_21828,N_18305,N_17951);
nor U21829 (N_21829,N_19936,N_17711);
or U21830 (N_21830,N_18793,N_18324);
and U21831 (N_21831,N_19933,N_19423);
xnor U21832 (N_21832,N_18225,N_19106);
nand U21833 (N_21833,N_17816,N_19188);
xor U21834 (N_21834,N_18153,N_19208);
xor U21835 (N_21835,N_19996,N_18170);
and U21836 (N_21836,N_19052,N_18612);
xnor U21837 (N_21837,N_19928,N_17850);
nand U21838 (N_21838,N_18039,N_18693);
nor U21839 (N_21839,N_19375,N_19208);
nand U21840 (N_21840,N_19931,N_18538);
nand U21841 (N_21841,N_19441,N_19297);
or U21842 (N_21842,N_19139,N_19731);
and U21843 (N_21843,N_17756,N_18258);
nand U21844 (N_21844,N_18672,N_17745);
nand U21845 (N_21845,N_18189,N_17907);
nor U21846 (N_21846,N_17794,N_18774);
nand U21847 (N_21847,N_17975,N_18991);
or U21848 (N_21848,N_18232,N_18871);
nor U21849 (N_21849,N_18259,N_19349);
nand U21850 (N_21850,N_19300,N_18741);
or U21851 (N_21851,N_19908,N_18380);
nor U21852 (N_21852,N_18310,N_18887);
xnor U21853 (N_21853,N_19041,N_18881);
or U21854 (N_21854,N_19938,N_18365);
or U21855 (N_21855,N_19876,N_18717);
and U21856 (N_21856,N_18552,N_19010);
and U21857 (N_21857,N_19718,N_19781);
nand U21858 (N_21858,N_18464,N_17897);
nand U21859 (N_21859,N_19450,N_19309);
nor U21860 (N_21860,N_19988,N_19287);
nor U21861 (N_21861,N_17723,N_18990);
nand U21862 (N_21862,N_17562,N_18504);
or U21863 (N_21863,N_18758,N_19184);
and U21864 (N_21864,N_19985,N_18359);
and U21865 (N_21865,N_18986,N_18845);
or U21866 (N_21866,N_18080,N_19671);
nor U21867 (N_21867,N_18263,N_18574);
xor U21868 (N_21868,N_18271,N_17509);
nor U21869 (N_21869,N_19323,N_19157);
and U21870 (N_21870,N_18132,N_17881);
and U21871 (N_21871,N_18400,N_19081);
nor U21872 (N_21872,N_19529,N_19240);
and U21873 (N_21873,N_19832,N_17954);
or U21874 (N_21874,N_19017,N_19658);
nand U21875 (N_21875,N_19368,N_18220);
or U21876 (N_21876,N_18490,N_18647);
nor U21877 (N_21877,N_18497,N_19091);
or U21878 (N_21878,N_19871,N_19313);
and U21879 (N_21879,N_17811,N_18816);
or U21880 (N_21880,N_19694,N_18024);
nor U21881 (N_21881,N_18139,N_18014);
and U21882 (N_21882,N_17680,N_18044);
and U21883 (N_21883,N_19889,N_19093);
nor U21884 (N_21884,N_18475,N_17970);
and U21885 (N_21885,N_19628,N_18115);
xnor U21886 (N_21886,N_17821,N_17597);
and U21887 (N_21887,N_17538,N_18924);
or U21888 (N_21888,N_17718,N_17641);
and U21889 (N_21889,N_17951,N_18465);
nand U21890 (N_21890,N_19610,N_18541);
or U21891 (N_21891,N_17810,N_19140);
nor U21892 (N_21892,N_19955,N_18030);
xnor U21893 (N_21893,N_17541,N_17591);
nor U21894 (N_21894,N_18753,N_18963);
and U21895 (N_21895,N_17547,N_17597);
and U21896 (N_21896,N_19821,N_17983);
nand U21897 (N_21897,N_19368,N_19238);
xor U21898 (N_21898,N_19373,N_19273);
nor U21899 (N_21899,N_17646,N_19687);
nor U21900 (N_21900,N_18102,N_18346);
or U21901 (N_21901,N_18976,N_18646);
or U21902 (N_21902,N_19465,N_18994);
or U21903 (N_21903,N_19358,N_19491);
nand U21904 (N_21904,N_19220,N_19688);
or U21905 (N_21905,N_18644,N_18391);
xor U21906 (N_21906,N_18715,N_18959);
or U21907 (N_21907,N_18294,N_19170);
nor U21908 (N_21908,N_19537,N_19770);
and U21909 (N_21909,N_19743,N_18570);
nor U21910 (N_21910,N_18492,N_18236);
xnor U21911 (N_21911,N_18936,N_19386);
xor U21912 (N_21912,N_18268,N_17855);
nor U21913 (N_21913,N_18008,N_19143);
or U21914 (N_21914,N_19141,N_18566);
and U21915 (N_21915,N_17975,N_18824);
or U21916 (N_21916,N_18216,N_19519);
xnor U21917 (N_21917,N_18585,N_19890);
and U21918 (N_21918,N_18205,N_17600);
xnor U21919 (N_21919,N_17805,N_18529);
nor U21920 (N_21920,N_18420,N_18613);
nor U21921 (N_21921,N_19255,N_18027);
xnor U21922 (N_21922,N_19502,N_18758);
xnor U21923 (N_21923,N_19821,N_17518);
and U21924 (N_21924,N_19357,N_17973);
xnor U21925 (N_21925,N_18969,N_18177);
xor U21926 (N_21926,N_18961,N_18394);
xnor U21927 (N_21927,N_18472,N_17627);
and U21928 (N_21928,N_18844,N_18093);
and U21929 (N_21929,N_18333,N_19623);
or U21930 (N_21930,N_18455,N_19981);
nor U21931 (N_21931,N_18714,N_17506);
xnor U21932 (N_21932,N_18995,N_17871);
xnor U21933 (N_21933,N_18996,N_18975);
nand U21934 (N_21934,N_19894,N_19534);
nand U21935 (N_21935,N_19252,N_18972);
and U21936 (N_21936,N_18416,N_18349);
nand U21937 (N_21937,N_19803,N_18961);
or U21938 (N_21938,N_18709,N_18939);
and U21939 (N_21939,N_18804,N_17572);
nand U21940 (N_21940,N_19870,N_19110);
nor U21941 (N_21941,N_18695,N_18520);
xnor U21942 (N_21942,N_19521,N_17770);
and U21943 (N_21943,N_19327,N_17971);
nor U21944 (N_21944,N_18088,N_19030);
nor U21945 (N_21945,N_19729,N_19927);
nand U21946 (N_21946,N_19474,N_18633);
or U21947 (N_21947,N_18679,N_18680);
xor U21948 (N_21948,N_18833,N_19317);
xor U21949 (N_21949,N_19858,N_17634);
nor U21950 (N_21950,N_19030,N_17771);
and U21951 (N_21951,N_19183,N_19871);
xnor U21952 (N_21952,N_19640,N_17697);
xnor U21953 (N_21953,N_19735,N_19789);
nor U21954 (N_21954,N_17679,N_18922);
and U21955 (N_21955,N_19242,N_19909);
or U21956 (N_21956,N_19800,N_18137);
or U21957 (N_21957,N_17820,N_19937);
and U21958 (N_21958,N_19925,N_19446);
or U21959 (N_21959,N_18769,N_19839);
and U21960 (N_21960,N_18229,N_19389);
xor U21961 (N_21961,N_17577,N_19724);
nand U21962 (N_21962,N_17996,N_19848);
nor U21963 (N_21963,N_19580,N_19491);
and U21964 (N_21964,N_19252,N_18039);
nor U21965 (N_21965,N_19599,N_17968);
and U21966 (N_21966,N_17555,N_18204);
xor U21967 (N_21967,N_17723,N_18940);
nor U21968 (N_21968,N_19180,N_17954);
nor U21969 (N_21969,N_17649,N_19661);
nand U21970 (N_21970,N_19616,N_18350);
xor U21971 (N_21971,N_18834,N_19861);
nand U21972 (N_21972,N_19492,N_18230);
and U21973 (N_21973,N_18388,N_18266);
nand U21974 (N_21974,N_18328,N_19284);
and U21975 (N_21975,N_19044,N_18797);
nor U21976 (N_21976,N_19734,N_19542);
xnor U21977 (N_21977,N_19948,N_18999);
xor U21978 (N_21978,N_19814,N_19684);
nand U21979 (N_21979,N_18281,N_19712);
nor U21980 (N_21980,N_18795,N_18183);
xnor U21981 (N_21981,N_19519,N_19200);
xor U21982 (N_21982,N_18453,N_19051);
nand U21983 (N_21983,N_19007,N_19547);
nand U21984 (N_21984,N_18152,N_17927);
nor U21985 (N_21985,N_18902,N_18500);
and U21986 (N_21986,N_19174,N_17829);
xnor U21987 (N_21987,N_19464,N_18764);
nand U21988 (N_21988,N_19979,N_19125);
nor U21989 (N_21989,N_18664,N_18825);
xor U21990 (N_21990,N_18628,N_17755);
and U21991 (N_21991,N_17623,N_17740);
nand U21992 (N_21992,N_19882,N_18170);
and U21993 (N_21993,N_19008,N_17947);
nor U21994 (N_21994,N_17971,N_19044);
nor U21995 (N_21995,N_17774,N_19515);
and U21996 (N_21996,N_18363,N_18525);
and U21997 (N_21997,N_19273,N_18360);
nand U21998 (N_21998,N_19519,N_18699);
nor U21999 (N_21999,N_18450,N_18252);
or U22000 (N_22000,N_17850,N_18267);
nand U22001 (N_22001,N_19835,N_18093);
or U22002 (N_22002,N_17508,N_18598);
nand U22003 (N_22003,N_19536,N_17739);
nand U22004 (N_22004,N_18794,N_18443);
and U22005 (N_22005,N_19054,N_17653);
nor U22006 (N_22006,N_19062,N_18442);
or U22007 (N_22007,N_18467,N_17555);
nor U22008 (N_22008,N_19351,N_19910);
nand U22009 (N_22009,N_17766,N_19335);
and U22010 (N_22010,N_17625,N_19151);
nand U22011 (N_22011,N_18088,N_19162);
or U22012 (N_22012,N_19217,N_18231);
xor U22013 (N_22013,N_18551,N_19535);
nor U22014 (N_22014,N_17949,N_18548);
nor U22015 (N_22015,N_18418,N_17624);
nand U22016 (N_22016,N_19681,N_17758);
or U22017 (N_22017,N_19336,N_18796);
nand U22018 (N_22018,N_19008,N_19756);
xnor U22019 (N_22019,N_19745,N_19026);
or U22020 (N_22020,N_19122,N_19347);
nand U22021 (N_22021,N_19868,N_18565);
or U22022 (N_22022,N_18319,N_18274);
and U22023 (N_22023,N_18211,N_18378);
or U22024 (N_22024,N_18368,N_19683);
nand U22025 (N_22025,N_19615,N_18178);
xnor U22026 (N_22026,N_18575,N_17544);
or U22027 (N_22027,N_19586,N_18175);
or U22028 (N_22028,N_19644,N_19151);
nand U22029 (N_22029,N_17657,N_18565);
and U22030 (N_22030,N_18194,N_19689);
and U22031 (N_22031,N_19301,N_17655);
nor U22032 (N_22032,N_18208,N_18044);
and U22033 (N_22033,N_19631,N_19447);
xnor U22034 (N_22034,N_19617,N_18307);
xnor U22035 (N_22035,N_18435,N_18158);
or U22036 (N_22036,N_19914,N_18231);
and U22037 (N_22037,N_19896,N_17718);
or U22038 (N_22038,N_18379,N_19781);
or U22039 (N_22039,N_19290,N_18674);
or U22040 (N_22040,N_18513,N_18749);
or U22041 (N_22041,N_19252,N_18904);
nand U22042 (N_22042,N_19386,N_19381);
xnor U22043 (N_22043,N_18879,N_18722);
nand U22044 (N_22044,N_17792,N_19049);
or U22045 (N_22045,N_18383,N_18478);
or U22046 (N_22046,N_18986,N_19531);
nor U22047 (N_22047,N_18236,N_17990);
or U22048 (N_22048,N_17950,N_18796);
and U22049 (N_22049,N_18024,N_19072);
or U22050 (N_22050,N_18633,N_19838);
nand U22051 (N_22051,N_17501,N_17778);
xnor U22052 (N_22052,N_17881,N_18766);
or U22053 (N_22053,N_17949,N_18424);
nand U22054 (N_22054,N_19037,N_18020);
nand U22055 (N_22055,N_17940,N_17572);
nand U22056 (N_22056,N_19258,N_19539);
and U22057 (N_22057,N_18173,N_17653);
xor U22058 (N_22058,N_19162,N_17724);
nand U22059 (N_22059,N_19208,N_18758);
xor U22060 (N_22060,N_18263,N_18980);
and U22061 (N_22061,N_17605,N_19136);
nand U22062 (N_22062,N_18013,N_17652);
and U22063 (N_22063,N_18980,N_19196);
nand U22064 (N_22064,N_17525,N_18336);
nand U22065 (N_22065,N_18049,N_18192);
nor U22066 (N_22066,N_19283,N_18904);
xor U22067 (N_22067,N_18170,N_19233);
or U22068 (N_22068,N_18553,N_18516);
or U22069 (N_22069,N_19787,N_18240);
or U22070 (N_22070,N_18589,N_18827);
nand U22071 (N_22071,N_18410,N_17568);
nor U22072 (N_22072,N_18482,N_18441);
nand U22073 (N_22073,N_17600,N_18819);
or U22074 (N_22074,N_18738,N_18333);
nor U22075 (N_22075,N_17679,N_18887);
nor U22076 (N_22076,N_19825,N_18485);
or U22077 (N_22077,N_19302,N_18055);
nand U22078 (N_22078,N_19085,N_19481);
nand U22079 (N_22079,N_19368,N_18624);
and U22080 (N_22080,N_18308,N_19377);
nand U22081 (N_22081,N_18135,N_18131);
xor U22082 (N_22082,N_19269,N_18520);
and U22083 (N_22083,N_18866,N_19153);
xor U22084 (N_22084,N_18104,N_18603);
and U22085 (N_22085,N_19555,N_17658);
or U22086 (N_22086,N_19852,N_18443);
nor U22087 (N_22087,N_19438,N_17874);
nor U22088 (N_22088,N_18006,N_19424);
and U22089 (N_22089,N_19878,N_19301);
and U22090 (N_22090,N_19523,N_19110);
and U22091 (N_22091,N_19048,N_19749);
nor U22092 (N_22092,N_19990,N_19269);
or U22093 (N_22093,N_18671,N_19585);
nand U22094 (N_22094,N_17662,N_19579);
nor U22095 (N_22095,N_17560,N_17648);
or U22096 (N_22096,N_18812,N_19710);
nor U22097 (N_22097,N_18422,N_18642);
or U22098 (N_22098,N_19086,N_18111);
nor U22099 (N_22099,N_19195,N_18851);
xor U22100 (N_22100,N_19594,N_18521);
and U22101 (N_22101,N_18931,N_18219);
xor U22102 (N_22102,N_19189,N_17646);
and U22103 (N_22103,N_19806,N_19323);
or U22104 (N_22104,N_17934,N_18986);
and U22105 (N_22105,N_18962,N_18695);
xnor U22106 (N_22106,N_18171,N_18094);
xnor U22107 (N_22107,N_17579,N_19426);
nor U22108 (N_22108,N_18038,N_19321);
xor U22109 (N_22109,N_18205,N_19267);
and U22110 (N_22110,N_19829,N_18649);
xnor U22111 (N_22111,N_17951,N_19188);
nor U22112 (N_22112,N_19369,N_19539);
nand U22113 (N_22113,N_19543,N_19337);
xnor U22114 (N_22114,N_18416,N_18327);
or U22115 (N_22115,N_18687,N_19022);
and U22116 (N_22116,N_17788,N_19249);
nand U22117 (N_22117,N_19956,N_17866);
and U22118 (N_22118,N_19729,N_19733);
nand U22119 (N_22119,N_19381,N_18118);
or U22120 (N_22120,N_17509,N_19118);
nor U22121 (N_22121,N_19878,N_19051);
or U22122 (N_22122,N_19491,N_18659);
nand U22123 (N_22123,N_18012,N_18634);
nor U22124 (N_22124,N_18161,N_19274);
nand U22125 (N_22125,N_19088,N_17560);
nor U22126 (N_22126,N_19478,N_18000);
or U22127 (N_22127,N_18072,N_19602);
nand U22128 (N_22128,N_19805,N_18824);
nor U22129 (N_22129,N_18065,N_19648);
or U22130 (N_22130,N_19475,N_17823);
and U22131 (N_22131,N_18068,N_19556);
xnor U22132 (N_22132,N_19142,N_19238);
and U22133 (N_22133,N_18078,N_17882);
nor U22134 (N_22134,N_18367,N_19049);
nand U22135 (N_22135,N_18693,N_18146);
and U22136 (N_22136,N_18912,N_17816);
or U22137 (N_22137,N_19143,N_18029);
nand U22138 (N_22138,N_19013,N_18855);
nor U22139 (N_22139,N_17517,N_19848);
xnor U22140 (N_22140,N_17800,N_17755);
xor U22141 (N_22141,N_18719,N_18988);
xor U22142 (N_22142,N_18154,N_18650);
nand U22143 (N_22143,N_18799,N_17626);
nand U22144 (N_22144,N_19983,N_18143);
and U22145 (N_22145,N_19659,N_18536);
and U22146 (N_22146,N_18295,N_17846);
or U22147 (N_22147,N_17613,N_17959);
nor U22148 (N_22148,N_19688,N_19308);
xor U22149 (N_22149,N_19594,N_19103);
xnor U22150 (N_22150,N_18758,N_18679);
nand U22151 (N_22151,N_18297,N_18554);
nor U22152 (N_22152,N_18654,N_19668);
nand U22153 (N_22153,N_17874,N_18932);
xor U22154 (N_22154,N_17549,N_18376);
xnor U22155 (N_22155,N_18040,N_18652);
and U22156 (N_22156,N_17572,N_19939);
nand U22157 (N_22157,N_19554,N_17826);
nand U22158 (N_22158,N_18762,N_19110);
nand U22159 (N_22159,N_18569,N_18643);
and U22160 (N_22160,N_18194,N_19906);
nand U22161 (N_22161,N_17703,N_19476);
and U22162 (N_22162,N_18798,N_18270);
nand U22163 (N_22163,N_18013,N_19412);
xor U22164 (N_22164,N_17876,N_18573);
nor U22165 (N_22165,N_19175,N_18140);
xnor U22166 (N_22166,N_18250,N_17840);
xor U22167 (N_22167,N_19577,N_19831);
or U22168 (N_22168,N_19385,N_18426);
xnor U22169 (N_22169,N_18103,N_19455);
nand U22170 (N_22170,N_18301,N_18175);
or U22171 (N_22171,N_19218,N_18003);
or U22172 (N_22172,N_17831,N_19574);
and U22173 (N_22173,N_19440,N_19574);
nand U22174 (N_22174,N_19168,N_18728);
nor U22175 (N_22175,N_19550,N_19458);
nor U22176 (N_22176,N_19599,N_18251);
nor U22177 (N_22177,N_17656,N_18465);
nor U22178 (N_22178,N_18006,N_19397);
nand U22179 (N_22179,N_18295,N_18516);
xor U22180 (N_22180,N_18131,N_17905);
xnor U22181 (N_22181,N_18838,N_18822);
or U22182 (N_22182,N_18092,N_18964);
nand U22183 (N_22183,N_18376,N_18706);
xnor U22184 (N_22184,N_18000,N_19556);
nor U22185 (N_22185,N_19718,N_18175);
nor U22186 (N_22186,N_17932,N_19122);
xor U22187 (N_22187,N_18229,N_18006);
and U22188 (N_22188,N_19208,N_18419);
or U22189 (N_22189,N_17713,N_19527);
nor U22190 (N_22190,N_18898,N_18654);
xor U22191 (N_22191,N_18074,N_19406);
nand U22192 (N_22192,N_17805,N_19870);
and U22193 (N_22193,N_18570,N_19616);
xnor U22194 (N_22194,N_18311,N_18394);
nor U22195 (N_22195,N_19474,N_19676);
and U22196 (N_22196,N_18831,N_19368);
or U22197 (N_22197,N_18116,N_18967);
or U22198 (N_22198,N_18599,N_19206);
and U22199 (N_22199,N_17540,N_19535);
nor U22200 (N_22200,N_17792,N_19357);
or U22201 (N_22201,N_18291,N_18049);
xnor U22202 (N_22202,N_17974,N_18206);
nand U22203 (N_22203,N_19643,N_17785);
xor U22204 (N_22204,N_19108,N_18267);
xor U22205 (N_22205,N_18627,N_18445);
xor U22206 (N_22206,N_19994,N_19611);
xor U22207 (N_22207,N_18666,N_17582);
or U22208 (N_22208,N_19145,N_19551);
and U22209 (N_22209,N_18098,N_18259);
nor U22210 (N_22210,N_18504,N_17749);
or U22211 (N_22211,N_18540,N_17662);
or U22212 (N_22212,N_19231,N_18065);
or U22213 (N_22213,N_19459,N_18309);
nand U22214 (N_22214,N_18122,N_18806);
nand U22215 (N_22215,N_19052,N_18539);
and U22216 (N_22216,N_18921,N_19603);
nand U22217 (N_22217,N_18196,N_18864);
nand U22218 (N_22218,N_19060,N_18366);
xnor U22219 (N_22219,N_18483,N_18733);
nand U22220 (N_22220,N_17545,N_18781);
and U22221 (N_22221,N_18787,N_19726);
xor U22222 (N_22222,N_18862,N_17871);
xor U22223 (N_22223,N_19111,N_17587);
or U22224 (N_22224,N_17516,N_18082);
and U22225 (N_22225,N_17982,N_19460);
xor U22226 (N_22226,N_18169,N_18771);
nor U22227 (N_22227,N_18899,N_19233);
nand U22228 (N_22228,N_17832,N_19686);
xor U22229 (N_22229,N_19235,N_19142);
and U22230 (N_22230,N_19737,N_18924);
nor U22231 (N_22231,N_19905,N_19207);
nand U22232 (N_22232,N_18388,N_18357);
xnor U22233 (N_22233,N_18277,N_19563);
or U22234 (N_22234,N_18587,N_19345);
xnor U22235 (N_22235,N_19271,N_19510);
nand U22236 (N_22236,N_17735,N_18618);
nor U22237 (N_22237,N_18801,N_19153);
nand U22238 (N_22238,N_18050,N_19426);
nand U22239 (N_22239,N_18578,N_18353);
nand U22240 (N_22240,N_19082,N_19097);
nor U22241 (N_22241,N_19811,N_19989);
or U22242 (N_22242,N_18031,N_17774);
nand U22243 (N_22243,N_19514,N_19053);
nor U22244 (N_22244,N_17585,N_19097);
and U22245 (N_22245,N_19428,N_19867);
nor U22246 (N_22246,N_19035,N_19389);
nand U22247 (N_22247,N_18942,N_18556);
and U22248 (N_22248,N_19073,N_19504);
or U22249 (N_22249,N_17764,N_17879);
xnor U22250 (N_22250,N_19261,N_18653);
xnor U22251 (N_22251,N_18888,N_18140);
nand U22252 (N_22252,N_19215,N_18637);
nor U22253 (N_22253,N_19340,N_19282);
nor U22254 (N_22254,N_17855,N_18760);
nor U22255 (N_22255,N_19192,N_19303);
xnor U22256 (N_22256,N_18753,N_17722);
xor U22257 (N_22257,N_17676,N_18882);
xnor U22258 (N_22258,N_19610,N_19184);
xor U22259 (N_22259,N_19563,N_19719);
nor U22260 (N_22260,N_17703,N_19710);
and U22261 (N_22261,N_17615,N_18218);
or U22262 (N_22262,N_19083,N_18836);
nand U22263 (N_22263,N_18593,N_19065);
nor U22264 (N_22264,N_19126,N_19129);
or U22265 (N_22265,N_17762,N_19019);
nand U22266 (N_22266,N_18008,N_18405);
nor U22267 (N_22267,N_17695,N_19335);
nand U22268 (N_22268,N_19912,N_18841);
nand U22269 (N_22269,N_19532,N_19380);
nand U22270 (N_22270,N_18183,N_17981);
xnor U22271 (N_22271,N_19530,N_19246);
xnor U22272 (N_22272,N_19984,N_19614);
and U22273 (N_22273,N_19234,N_19341);
xor U22274 (N_22274,N_19300,N_17790);
or U22275 (N_22275,N_18881,N_18448);
nor U22276 (N_22276,N_18061,N_19073);
or U22277 (N_22277,N_19912,N_18899);
and U22278 (N_22278,N_17854,N_17716);
xnor U22279 (N_22279,N_17574,N_19963);
and U22280 (N_22280,N_19284,N_19306);
xnor U22281 (N_22281,N_19942,N_19607);
xor U22282 (N_22282,N_17972,N_17845);
nand U22283 (N_22283,N_19551,N_18712);
nor U22284 (N_22284,N_19383,N_18153);
nor U22285 (N_22285,N_18152,N_17978);
nand U22286 (N_22286,N_17838,N_18667);
xnor U22287 (N_22287,N_19797,N_19891);
or U22288 (N_22288,N_17674,N_17974);
and U22289 (N_22289,N_18711,N_18160);
and U22290 (N_22290,N_17505,N_18637);
or U22291 (N_22291,N_19642,N_19812);
xnor U22292 (N_22292,N_19805,N_19673);
or U22293 (N_22293,N_19013,N_18610);
and U22294 (N_22294,N_19427,N_19797);
xnor U22295 (N_22295,N_19327,N_17512);
nand U22296 (N_22296,N_19610,N_17521);
nand U22297 (N_22297,N_18844,N_19338);
nor U22298 (N_22298,N_19249,N_18485);
and U22299 (N_22299,N_19388,N_19104);
nand U22300 (N_22300,N_19017,N_18875);
and U22301 (N_22301,N_18084,N_18939);
or U22302 (N_22302,N_18027,N_19103);
or U22303 (N_22303,N_17926,N_19031);
and U22304 (N_22304,N_19307,N_18676);
xnor U22305 (N_22305,N_18973,N_17574);
nor U22306 (N_22306,N_17986,N_19462);
and U22307 (N_22307,N_17830,N_18257);
and U22308 (N_22308,N_17763,N_18593);
and U22309 (N_22309,N_19203,N_19050);
nand U22310 (N_22310,N_17962,N_17842);
nor U22311 (N_22311,N_18264,N_17876);
nor U22312 (N_22312,N_18261,N_19947);
nand U22313 (N_22313,N_19758,N_18301);
or U22314 (N_22314,N_18000,N_18459);
or U22315 (N_22315,N_18495,N_18775);
nor U22316 (N_22316,N_19659,N_18376);
nand U22317 (N_22317,N_18806,N_19804);
xnor U22318 (N_22318,N_18095,N_18885);
nand U22319 (N_22319,N_19586,N_18133);
and U22320 (N_22320,N_19281,N_18621);
nand U22321 (N_22321,N_19657,N_18823);
and U22322 (N_22322,N_19445,N_17725);
or U22323 (N_22323,N_18020,N_18138);
and U22324 (N_22324,N_18182,N_18791);
nand U22325 (N_22325,N_19003,N_19502);
nor U22326 (N_22326,N_18887,N_19989);
nand U22327 (N_22327,N_18512,N_18029);
nand U22328 (N_22328,N_18765,N_18779);
xor U22329 (N_22329,N_17595,N_18655);
or U22330 (N_22330,N_19321,N_18149);
xnor U22331 (N_22331,N_18654,N_17772);
or U22332 (N_22332,N_19775,N_18353);
or U22333 (N_22333,N_18396,N_17608);
nor U22334 (N_22334,N_19921,N_17757);
nand U22335 (N_22335,N_19836,N_18679);
nor U22336 (N_22336,N_18470,N_19522);
and U22337 (N_22337,N_18515,N_18338);
nor U22338 (N_22338,N_19507,N_18833);
and U22339 (N_22339,N_18859,N_19089);
nand U22340 (N_22340,N_19628,N_19995);
and U22341 (N_22341,N_18317,N_19430);
xnor U22342 (N_22342,N_19052,N_19228);
and U22343 (N_22343,N_19789,N_17739);
or U22344 (N_22344,N_18177,N_19311);
or U22345 (N_22345,N_17742,N_19824);
nor U22346 (N_22346,N_18902,N_17577);
nor U22347 (N_22347,N_19446,N_18594);
and U22348 (N_22348,N_18542,N_17973);
xnor U22349 (N_22349,N_18481,N_17955);
xor U22350 (N_22350,N_18134,N_17537);
and U22351 (N_22351,N_17548,N_19552);
nor U22352 (N_22352,N_18666,N_19736);
xor U22353 (N_22353,N_17808,N_18695);
or U22354 (N_22354,N_18647,N_19647);
or U22355 (N_22355,N_19117,N_17700);
and U22356 (N_22356,N_19674,N_19387);
and U22357 (N_22357,N_18270,N_19601);
and U22358 (N_22358,N_17915,N_19753);
or U22359 (N_22359,N_19992,N_19460);
nor U22360 (N_22360,N_18613,N_19103);
and U22361 (N_22361,N_17930,N_18432);
nor U22362 (N_22362,N_18414,N_18290);
or U22363 (N_22363,N_19854,N_17543);
and U22364 (N_22364,N_18378,N_19359);
nand U22365 (N_22365,N_18709,N_17686);
or U22366 (N_22366,N_18037,N_18914);
nand U22367 (N_22367,N_18994,N_19881);
or U22368 (N_22368,N_18552,N_18791);
or U22369 (N_22369,N_18097,N_18872);
or U22370 (N_22370,N_18855,N_18800);
nor U22371 (N_22371,N_17720,N_19794);
nand U22372 (N_22372,N_19158,N_18634);
or U22373 (N_22373,N_19327,N_18346);
xnor U22374 (N_22374,N_17971,N_18424);
nor U22375 (N_22375,N_18791,N_17508);
or U22376 (N_22376,N_19172,N_19572);
and U22377 (N_22377,N_19635,N_19906);
or U22378 (N_22378,N_18347,N_19436);
and U22379 (N_22379,N_19966,N_17849);
or U22380 (N_22380,N_19461,N_17771);
nand U22381 (N_22381,N_19023,N_19334);
and U22382 (N_22382,N_18294,N_19333);
or U22383 (N_22383,N_18341,N_17543);
nand U22384 (N_22384,N_18765,N_17628);
and U22385 (N_22385,N_19118,N_18727);
nand U22386 (N_22386,N_17719,N_19215);
or U22387 (N_22387,N_18591,N_18460);
nor U22388 (N_22388,N_17881,N_19579);
xnor U22389 (N_22389,N_19342,N_18542);
nand U22390 (N_22390,N_18455,N_18601);
or U22391 (N_22391,N_18743,N_18474);
or U22392 (N_22392,N_19511,N_18982);
nand U22393 (N_22393,N_19379,N_18703);
or U22394 (N_22394,N_18423,N_19561);
and U22395 (N_22395,N_18541,N_19054);
nand U22396 (N_22396,N_18085,N_18334);
xnor U22397 (N_22397,N_17777,N_19961);
xor U22398 (N_22398,N_18442,N_18202);
or U22399 (N_22399,N_17821,N_19109);
nor U22400 (N_22400,N_17560,N_19815);
nand U22401 (N_22401,N_17524,N_18865);
nand U22402 (N_22402,N_17634,N_19234);
nand U22403 (N_22403,N_18191,N_18453);
nand U22404 (N_22404,N_19787,N_18950);
and U22405 (N_22405,N_17744,N_19879);
nor U22406 (N_22406,N_19235,N_17912);
and U22407 (N_22407,N_19239,N_19906);
and U22408 (N_22408,N_19219,N_19972);
nor U22409 (N_22409,N_19223,N_19346);
nor U22410 (N_22410,N_17776,N_18966);
or U22411 (N_22411,N_18498,N_18827);
nand U22412 (N_22412,N_18210,N_18691);
nor U22413 (N_22413,N_19254,N_19044);
or U22414 (N_22414,N_19920,N_18486);
or U22415 (N_22415,N_17510,N_18737);
nand U22416 (N_22416,N_17716,N_17793);
nor U22417 (N_22417,N_18509,N_17758);
and U22418 (N_22418,N_19045,N_18773);
or U22419 (N_22419,N_17648,N_18555);
or U22420 (N_22420,N_18881,N_18308);
nand U22421 (N_22421,N_18151,N_18033);
or U22422 (N_22422,N_18789,N_18466);
nand U22423 (N_22423,N_17808,N_18857);
nand U22424 (N_22424,N_18973,N_19123);
xnor U22425 (N_22425,N_18475,N_17869);
nand U22426 (N_22426,N_19771,N_18342);
nor U22427 (N_22427,N_19921,N_17962);
and U22428 (N_22428,N_19367,N_18076);
or U22429 (N_22429,N_19343,N_18931);
nand U22430 (N_22430,N_19400,N_19332);
nor U22431 (N_22431,N_17640,N_18783);
nor U22432 (N_22432,N_17598,N_19831);
nor U22433 (N_22433,N_18621,N_17864);
nand U22434 (N_22434,N_17779,N_19483);
xor U22435 (N_22435,N_18325,N_19979);
and U22436 (N_22436,N_17581,N_18318);
and U22437 (N_22437,N_19742,N_18336);
xnor U22438 (N_22438,N_19866,N_18660);
and U22439 (N_22439,N_18494,N_19726);
nor U22440 (N_22440,N_18345,N_19051);
nor U22441 (N_22441,N_18153,N_19175);
xnor U22442 (N_22442,N_19135,N_19742);
and U22443 (N_22443,N_19823,N_19490);
or U22444 (N_22444,N_19946,N_18963);
or U22445 (N_22445,N_19944,N_18659);
xnor U22446 (N_22446,N_18771,N_17639);
and U22447 (N_22447,N_17825,N_17636);
and U22448 (N_22448,N_18286,N_19435);
and U22449 (N_22449,N_18747,N_19997);
or U22450 (N_22450,N_18658,N_19549);
nor U22451 (N_22451,N_18915,N_18849);
nor U22452 (N_22452,N_19675,N_18366);
or U22453 (N_22453,N_19109,N_18209);
nor U22454 (N_22454,N_18611,N_18836);
and U22455 (N_22455,N_17849,N_18926);
xor U22456 (N_22456,N_18249,N_17843);
and U22457 (N_22457,N_18132,N_19912);
and U22458 (N_22458,N_19425,N_17855);
nand U22459 (N_22459,N_19144,N_18773);
and U22460 (N_22460,N_18902,N_17702);
nand U22461 (N_22461,N_17597,N_18414);
or U22462 (N_22462,N_18880,N_18021);
or U22463 (N_22463,N_19098,N_18160);
and U22464 (N_22464,N_18201,N_17922);
nand U22465 (N_22465,N_18103,N_17914);
nand U22466 (N_22466,N_18816,N_19127);
or U22467 (N_22467,N_18445,N_19270);
nand U22468 (N_22468,N_18568,N_18057);
nand U22469 (N_22469,N_18460,N_19531);
and U22470 (N_22470,N_19520,N_19414);
or U22471 (N_22471,N_18245,N_19176);
nand U22472 (N_22472,N_18159,N_17697);
xnor U22473 (N_22473,N_18034,N_18004);
nor U22474 (N_22474,N_19282,N_17551);
nor U22475 (N_22475,N_18826,N_19313);
xor U22476 (N_22476,N_18681,N_19117);
nor U22477 (N_22477,N_19039,N_19859);
and U22478 (N_22478,N_19641,N_18380);
or U22479 (N_22479,N_19777,N_18293);
and U22480 (N_22480,N_17694,N_19015);
and U22481 (N_22481,N_19117,N_18690);
or U22482 (N_22482,N_17826,N_18792);
and U22483 (N_22483,N_19583,N_17762);
or U22484 (N_22484,N_19233,N_18671);
xor U22485 (N_22485,N_18235,N_17514);
and U22486 (N_22486,N_18260,N_19269);
nor U22487 (N_22487,N_18356,N_19659);
xnor U22488 (N_22488,N_18011,N_19971);
or U22489 (N_22489,N_19049,N_17637);
or U22490 (N_22490,N_17880,N_18157);
nor U22491 (N_22491,N_19133,N_18913);
and U22492 (N_22492,N_18793,N_19917);
and U22493 (N_22493,N_18447,N_18736);
nor U22494 (N_22494,N_19477,N_19318);
or U22495 (N_22495,N_18055,N_18508);
nor U22496 (N_22496,N_19557,N_19545);
nor U22497 (N_22497,N_19987,N_18456);
and U22498 (N_22498,N_19021,N_17616);
nand U22499 (N_22499,N_19276,N_18945);
xor U22500 (N_22500,N_21375,N_21663);
nor U22501 (N_22501,N_20722,N_20995);
nor U22502 (N_22502,N_20864,N_21606);
or U22503 (N_22503,N_22351,N_22231);
nand U22504 (N_22504,N_20752,N_21153);
or U22505 (N_22505,N_20213,N_21665);
xnor U22506 (N_22506,N_22263,N_21285);
or U22507 (N_22507,N_21897,N_22009);
nand U22508 (N_22508,N_20252,N_22473);
and U22509 (N_22509,N_21392,N_22395);
xnor U22510 (N_22510,N_22301,N_22293);
and U22511 (N_22511,N_22305,N_21998);
nor U22512 (N_22512,N_22219,N_20781);
nor U22513 (N_22513,N_21825,N_21910);
nand U22514 (N_22514,N_20868,N_20943);
xnor U22515 (N_22515,N_21247,N_20518);
and U22516 (N_22516,N_20225,N_21455);
xor U22517 (N_22517,N_21556,N_20556);
or U22518 (N_22518,N_21369,N_20942);
or U22519 (N_22519,N_22382,N_20650);
or U22520 (N_22520,N_20396,N_20885);
xnor U22521 (N_22521,N_22255,N_22157);
and U22522 (N_22522,N_22410,N_20585);
xor U22523 (N_22523,N_20709,N_22215);
nor U22524 (N_22524,N_20140,N_22398);
and U22525 (N_22525,N_22432,N_21016);
nand U22526 (N_22526,N_20229,N_20680);
nand U22527 (N_22527,N_21751,N_22026);
xnor U22528 (N_22528,N_20924,N_21077);
xor U22529 (N_22529,N_21393,N_20121);
nand U22530 (N_22530,N_21734,N_21299);
nand U22531 (N_22531,N_20696,N_20871);
nand U22532 (N_22532,N_21927,N_21164);
nand U22533 (N_22533,N_21633,N_20976);
xor U22534 (N_22534,N_22133,N_20228);
xor U22535 (N_22535,N_20199,N_20082);
nand U22536 (N_22536,N_21487,N_22274);
nor U22537 (N_22537,N_22162,N_20936);
xnor U22538 (N_22538,N_21173,N_20381);
and U22539 (N_22539,N_22191,N_20421);
and U22540 (N_22540,N_21997,N_20046);
nand U22541 (N_22541,N_20376,N_21205);
xnor U22542 (N_22542,N_21182,N_20548);
nand U22543 (N_22543,N_22006,N_22053);
and U22544 (N_22544,N_20125,N_21593);
or U22545 (N_22545,N_21072,N_22275);
xnor U22546 (N_22546,N_21968,N_21097);
and U22547 (N_22547,N_21867,N_21919);
or U22548 (N_22548,N_21730,N_20947);
and U22549 (N_22549,N_20610,N_20857);
nor U22550 (N_22550,N_21436,N_20542);
nor U22551 (N_22551,N_20867,N_22063);
or U22552 (N_22552,N_21690,N_21559);
xnor U22553 (N_22553,N_20915,N_20134);
nand U22554 (N_22554,N_21971,N_20427);
xor U22555 (N_22555,N_21201,N_20766);
nor U22556 (N_22556,N_21470,N_21132);
xor U22557 (N_22557,N_21461,N_21847);
xor U22558 (N_22558,N_20838,N_21157);
nand U22559 (N_22559,N_20579,N_22295);
xor U22560 (N_22560,N_21036,N_20767);
nor U22561 (N_22561,N_20703,N_20632);
nand U22562 (N_22562,N_22059,N_21188);
and U22563 (N_22563,N_20623,N_20794);
nor U22564 (N_22564,N_21994,N_22159);
xnor U22565 (N_22565,N_20517,N_22490);
and U22566 (N_22566,N_20330,N_20823);
nor U22567 (N_22567,N_20979,N_22400);
and U22568 (N_22568,N_21141,N_21579);
nand U22569 (N_22569,N_20394,N_22271);
and U22570 (N_22570,N_21151,N_22047);
nand U22571 (N_22571,N_20844,N_21404);
nor U22572 (N_22572,N_21604,N_21992);
or U22573 (N_22573,N_22298,N_21373);
and U22574 (N_22574,N_22206,N_22299);
nand U22575 (N_22575,N_22349,N_22423);
nand U22576 (N_22576,N_20592,N_21017);
nor U22577 (N_22577,N_21826,N_21475);
or U22578 (N_22578,N_20404,N_22156);
and U22579 (N_22579,N_22233,N_21671);
nor U22580 (N_22580,N_22463,N_22135);
and U22581 (N_22581,N_20360,N_20522);
xnor U22582 (N_22582,N_21526,N_21323);
and U22583 (N_22583,N_22336,N_22049);
and U22584 (N_22584,N_22377,N_20222);
or U22585 (N_22585,N_21331,N_20303);
xnor U22586 (N_22586,N_22213,N_20185);
nand U22587 (N_22587,N_21830,N_22358);
xor U22588 (N_22588,N_21869,N_20711);
nand U22589 (N_22589,N_22252,N_21066);
and U22590 (N_22590,N_21549,N_20744);
and U22591 (N_22591,N_20695,N_22128);
xor U22592 (N_22592,N_22268,N_20965);
xnor U22593 (N_22593,N_20032,N_20092);
nand U22594 (N_22594,N_21854,N_22048);
xnor U22595 (N_22595,N_20903,N_21314);
or U22596 (N_22596,N_20710,N_20606);
nand U22597 (N_22597,N_20021,N_20999);
and U22598 (N_22598,N_21150,N_22331);
nand U22599 (N_22599,N_21948,N_20932);
or U22600 (N_22600,N_20079,N_22112);
nand U22601 (N_22601,N_21598,N_20509);
xnor U22602 (N_22602,N_20175,N_22467);
or U22603 (N_22603,N_22344,N_22326);
nor U22604 (N_22604,N_20118,N_20814);
xor U22605 (N_22605,N_21868,N_20900);
nand U22606 (N_22606,N_21144,N_20403);
xnor U22607 (N_22607,N_21935,N_20897);
xnor U22608 (N_22608,N_21602,N_21889);
and U22609 (N_22609,N_21000,N_20624);
or U22610 (N_22610,N_20042,N_21685);
nor U22611 (N_22611,N_21410,N_22454);
or U22612 (N_22612,N_21725,N_20786);
and U22613 (N_22613,N_20086,N_21710);
xor U22614 (N_22614,N_20634,N_22227);
nand U22615 (N_22615,N_20797,N_21506);
xnor U22616 (N_22616,N_20597,N_22054);
and U22617 (N_22617,N_21135,N_20078);
nor U22618 (N_22618,N_21381,N_20350);
nor U22619 (N_22619,N_20813,N_20869);
and U22620 (N_22620,N_20075,N_20436);
xor U22621 (N_22621,N_20973,N_22003);
and U22622 (N_22622,N_21440,N_20720);
or U22623 (N_22623,N_21419,N_20574);
nor U22624 (N_22624,N_21585,N_21763);
or U22625 (N_22625,N_20070,N_21528);
and U22626 (N_22626,N_21858,N_22038);
nand U22627 (N_22627,N_21672,N_21791);
or U22628 (N_22628,N_20980,N_21040);
xor U22629 (N_22629,N_20646,N_22447);
xor U22630 (N_22630,N_21399,N_21222);
and U22631 (N_22631,N_21566,N_22125);
nand U22632 (N_22632,N_20519,N_21319);
or U22633 (N_22633,N_20895,N_21865);
and U22634 (N_22634,N_21257,N_20790);
and U22635 (N_22635,N_21387,N_21864);
xnor U22636 (N_22636,N_22126,N_21228);
nand U22637 (N_22637,N_20656,N_20176);
and U22638 (N_22638,N_20017,N_21978);
and U22639 (N_22639,N_21263,N_20635);
nand U22640 (N_22640,N_21425,N_22105);
or U22641 (N_22641,N_21238,N_21025);
xor U22642 (N_22642,N_20174,N_20273);
or U22643 (N_22643,N_21915,N_20978);
nor U22644 (N_22644,N_22015,N_22402);
xor U22645 (N_22645,N_22070,N_20398);
xnor U22646 (N_22646,N_20494,N_20644);
nand U22647 (N_22647,N_22315,N_20798);
or U22648 (N_22648,N_21167,N_22401);
or U22649 (N_22649,N_20605,N_20254);
and U22650 (N_22650,N_21619,N_20312);
and U22651 (N_22651,N_21874,N_22118);
or U22652 (N_22652,N_20311,N_20777);
xor U22653 (N_22653,N_21177,N_22267);
nor U22654 (N_22654,N_22272,N_21286);
xnor U22655 (N_22655,N_22165,N_20670);
or U22656 (N_22656,N_20948,N_20365);
nor U22657 (N_22657,N_20166,N_22117);
or U22658 (N_22658,N_21248,N_21474);
nand U22659 (N_22659,N_22373,N_21824);
and U22660 (N_22660,N_20505,N_21415);
nand U22661 (N_22661,N_20609,N_20637);
nor U22662 (N_22662,N_21525,N_21533);
nor U22663 (N_22663,N_22071,N_21755);
nand U22664 (N_22664,N_22376,N_21091);
nand U22665 (N_22665,N_20926,N_22102);
xor U22666 (N_22666,N_21693,N_21784);
or U22667 (N_22667,N_20682,N_20158);
or U22668 (N_22668,N_21667,N_20690);
nor U22669 (N_22669,N_20861,N_22458);
nor U22670 (N_22670,N_20791,N_22142);
nor U22671 (N_22671,N_20465,N_21045);
nor U22672 (N_22672,N_21877,N_20458);
nand U22673 (N_22673,N_22014,N_22166);
and U22674 (N_22674,N_21115,N_22039);
xnor U22675 (N_22675,N_21575,N_20054);
and U22676 (N_22676,N_21493,N_21796);
xnor U22677 (N_22677,N_21850,N_21291);
nor U22678 (N_22678,N_21655,N_20387);
and U22679 (N_22679,N_21908,N_21152);
or U22680 (N_22680,N_20661,N_21512);
xnor U22681 (N_22681,N_21303,N_21804);
or U22682 (N_22682,N_20717,N_21609);
or U22683 (N_22683,N_21316,N_22290);
or U22684 (N_22684,N_20432,N_20329);
or U22685 (N_22685,N_20507,N_21273);
nand U22686 (N_22686,N_21518,N_22066);
nand U22687 (N_22687,N_22188,N_22235);
or U22688 (N_22688,N_20619,N_20383);
and U22689 (N_22689,N_21787,N_20860);
nor U22690 (N_22690,N_21843,N_20059);
nand U22691 (N_22691,N_21959,N_20968);
nor U22692 (N_22692,N_20570,N_20859);
nor U22693 (N_22693,N_22438,N_20004);
or U22694 (N_22694,N_20233,N_22228);
and U22695 (N_22695,N_21673,N_22388);
and U22696 (N_22696,N_20386,N_21428);
and U22697 (N_22697,N_20761,N_20916);
or U22698 (N_22698,N_20810,N_20935);
and U22699 (N_22699,N_21960,N_22197);
or U22700 (N_22700,N_21355,N_20099);
nor U22701 (N_22701,N_20490,N_22332);
nor U22702 (N_22702,N_21180,N_22248);
and U22703 (N_22703,N_20291,N_20066);
or U22704 (N_22704,N_20593,N_20776);
nand U22705 (N_22705,N_20728,N_20259);
or U22706 (N_22706,N_22346,N_21189);
xor U22707 (N_22707,N_20002,N_22359);
and U22708 (N_22708,N_20547,N_22074);
and U22709 (N_22709,N_21862,N_21210);
and U22710 (N_22710,N_20561,N_20789);
or U22711 (N_22711,N_21603,N_21343);
xnor U22712 (N_22712,N_20120,N_20706);
nand U22713 (N_22713,N_21922,N_20313);
nor U22714 (N_22714,N_20461,N_20622);
and U22715 (N_22715,N_20788,N_20697);
and U22716 (N_22716,N_21417,N_22010);
nand U22717 (N_22717,N_20039,N_20799);
nor U22718 (N_22718,N_21028,N_20256);
and U22719 (N_22719,N_21571,N_21772);
or U22720 (N_22720,N_21005,N_20994);
and U22721 (N_22721,N_21237,N_20841);
and U22722 (N_22722,N_21010,N_20468);
nand U22723 (N_22723,N_22236,N_22282);
or U22724 (N_22724,N_21274,N_22444);
xnor U22725 (N_22725,N_21148,N_21236);
nand U22726 (N_22726,N_22040,N_20364);
xor U22727 (N_22727,N_22325,N_20663);
or U22728 (N_22728,N_22285,N_22453);
and U22729 (N_22729,N_22088,N_21112);
or U22730 (N_22730,N_20564,N_21006);
and U22731 (N_22731,N_20485,N_21536);
nand U22732 (N_22732,N_20544,N_21795);
xor U22733 (N_22733,N_20827,N_20148);
and U22734 (N_22734,N_20025,N_21296);
nor U22735 (N_22735,N_21870,N_20455);
and U22736 (N_22736,N_22189,N_21437);
nor U22737 (N_22737,N_20685,N_21271);
nand U22738 (N_22738,N_20630,N_20563);
nand U22739 (N_22739,N_20629,N_20305);
or U22740 (N_22740,N_21995,N_21743);
or U22741 (N_22741,N_20482,N_20715);
nand U22742 (N_22742,N_22499,N_22451);
nor U22743 (N_22743,N_20076,N_22161);
nor U22744 (N_22744,N_20642,N_21562);
nand U22745 (N_22745,N_20253,N_21906);
xor U22746 (N_22746,N_21880,N_20601);
and U22747 (N_22747,N_21371,N_22435);
xor U22748 (N_22748,N_21856,N_20940);
xor U22749 (N_22749,N_20850,N_20196);
and U22750 (N_22750,N_21614,N_20114);
nor U22751 (N_22751,N_21714,N_20189);
nand U22752 (N_22752,N_21485,N_20912);
or U22753 (N_22753,N_20130,N_20904);
nor U22754 (N_22754,N_21996,N_20055);
nor U22755 (N_22755,N_21365,N_22424);
nor U22756 (N_22756,N_21557,N_21389);
nand U22757 (N_22757,N_21642,N_20603);
nor U22758 (N_22758,N_21241,N_21447);
and U22759 (N_22759,N_21081,N_21432);
or U22760 (N_22760,N_20090,N_21678);
nor U22761 (N_22761,N_21814,N_21591);
xnor U22762 (N_22762,N_21914,N_21810);
or U22763 (N_22763,N_22439,N_20466);
nand U22764 (N_22764,N_21165,N_21523);
nand U22765 (N_22765,N_21484,N_22368);
and U22766 (N_22766,N_22429,N_21728);
or U22767 (N_22767,N_21191,N_20881);
nand U22768 (N_22768,N_21260,N_20746);
nand U22769 (N_22769,N_20049,N_21721);
and U22770 (N_22770,N_20657,N_21508);
nor U22771 (N_22771,N_21053,N_22449);
nand U22772 (N_22772,N_20373,N_20489);
nand U22773 (N_22773,N_21888,N_21022);
xnor U22774 (N_22774,N_21354,N_22044);
nor U22775 (N_22775,N_21283,N_21762);
nor U22776 (N_22776,N_20280,N_21169);
nor U22777 (N_22777,N_21125,N_21809);
or U22778 (N_22778,N_20257,N_22442);
nand U22779 (N_22779,N_21021,N_22122);
and U22780 (N_22780,N_21050,N_22391);
xor U22781 (N_22781,N_20782,N_21403);
nor U22782 (N_22782,N_20156,N_20111);
and U22783 (N_22783,N_20566,N_21894);
nand U22784 (N_22784,N_20285,N_21278);
and U22785 (N_22785,N_22232,N_22276);
and U22786 (N_22786,N_22193,N_21746);
xor U22787 (N_22787,N_22115,N_21264);
nand U22788 (N_22788,N_21925,N_20986);
nand U22789 (N_22789,N_20759,N_20845);
nand U22790 (N_22790,N_21044,N_21815);
nand U22791 (N_22791,N_20545,N_22075);
xor U22792 (N_22792,N_22278,N_22329);
nand U22793 (N_22793,N_22257,N_21401);
nor U22794 (N_22794,N_20414,N_21033);
and U22795 (N_22795,N_21938,N_21058);
xnor U22796 (N_22796,N_21570,N_21691);
or U22797 (N_22797,N_22093,N_21659);
xnor U22798 (N_22798,N_20428,N_22001);
nand U22799 (N_22799,N_21962,N_20179);
or U22800 (N_22800,N_20723,N_20824);
xor U22801 (N_22801,N_21345,N_20358);
or U22802 (N_22802,N_20307,N_22243);
or U22803 (N_22803,N_21226,N_20407);
nor U22804 (N_22804,N_22050,N_20647);
xor U22805 (N_22805,N_21563,N_20769);
xnor U22806 (N_22806,N_22201,N_21510);
xnor U22807 (N_22807,N_20219,N_22472);
or U22808 (N_22808,N_20793,N_21406);
nor U22809 (N_22809,N_22216,N_20377);
and U22810 (N_22810,N_21356,N_20586);
and U22811 (N_22811,N_21262,N_20437);
xnor U22812 (N_22812,N_22330,N_22405);
or U22813 (N_22813,N_21706,N_20319);
and U22814 (N_22814,N_20502,N_20535);
xnor U22815 (N_22815,N_21550,N_20701);
or U22816 (N_22816,N_21459,N_20523);
or U22817 (N_22817,N_20462,N_22393);
nand U22818 (N_22818,N_20380,N_20829);
nand U22819 (N_22819,N_20512,N_21729);
and U22820 (N_22820,N_21414,N_20872);
or U22821 (N_22821,N_22296,N_21634);
nor U22822 (N_22822,N_20626,N_22154);
and U22823 (N_22823,N_22462,N_20530);
and U22824 (N_22824,N_20478,N_21653);
and U22825 (N_22825,N_21358,N_22364);
xnor U22826 (N_22826,N_21620,N_20992);
and U22827 (N_22827,N_20119,N_22341);
and U22828 (N_22828,N_20721,N_20889);
xor U22829 (N_22829,N_21680,N_21229);
or U22830 (N_22830,N_22323,N_21501);
nor U22831 (N_22831,N_20266,N_21084);
xnor U22832 (N_22832,N_20031,N_20007);
nor U22833 (N_22833,N_20539,N_22264);
nor U22834 (N_22834,N_22011,N_22194);
nand U22835 (N_22835,N_21713,N_20678);
xor U22836 (N_22836,N_20138,N_21255);
nand U22837 (N_22837,N_22476,N_20297);
and U22838 (N_22838,N_20045,N_20809);
xnor U22839 (N_22839,N_21329,N_20552);
and U22840 (N_22840,N_22459,N_21715);
nand U22841 (N_22841,N_22083,N_20057);
nand U22842 (N_22842,N_21617,N_22306);
nand U22843 (N_22843,N_22404,N_21088);
xor U22844 (N_22844,N_21096,N_21564);
nand U22845 (N_22845,N_22277,N_20348);
and U22846 (N_22846,N_20754,N_22307);
or U22847 (N_22847,N_22247,N_20424);
xnor U22848 (N_22848,N_21986,N_21702);
nand U22849 (N_22849,N_20843,N_21515);
or U22850 (N_22850,N_21532,N_21011);
nor U22851 (N_22851,N_20464,N_22378);
xor U22852 (N_22852,N_20359,N_21970);
nor U22853 (N_22853,N_21382,N_21929);
and U22854 (N_22854,N_20371,N_20426);
or U22855 (N_22855,N_21932,N_22149);
xor U22856 (N_22856,N_20875,N_20040);
nor U22857 (N_22857,N_21792,N_20499);
nor U22858 (N_22858,N_20191,N_22024);
nand U22859 (N_22859,N_21244,N_20802);
and U22860 (N_22860,N_20141,N_20217);
or U22861 (N_22861,N_20338,N_22132);
or U22862 (N_22862,N_21463,N_22036);
nand U22863 (N_22863,N_21321,N_20200);
and U22864 (N_22864,N_21396,N_22080);
xnor U22865 (N_22865,N_22407,N_21174);
and U22866 (N_22866,N_22057,N_21085);
or U22867 (N_22867,N_20016,N_22428);
or U22868 (N_22868,N_21335,N_20699);
xor U22869 (N_22869,N_20378,N_20083);
xor U22870 (N_22870,N_22374,N_21435);
nor U22871 (N_22871,N_21947,N_20308);
nand U22872 (N_22872,N_22324,N_20971);
xnor U22873 (N_22873,N_20149,N_20975);
nor U22874 (N_22874,N_20352,N_22079);
or U22875 (N_22875,N_21126,N_21307);
xor U22876 (N_22876,N_20208,N_22109);
or U22877 (N_22877,N_21531,N_20483);
nor U22878 (N_22878,N_20135,N_20104);
and U22879 (N_22879,N_20557,N_21430);
xor U22880 (N_22880,N_22062,N_20608);
nor U22881 (N_22881,N_20132,N_22380);
and U22882 (N_22882,N_20639,N_20631);
and U22883 (N_22883,N_21042,N_20613);
xnor U22884 (N_22884,N_20729,N_20908);
or U22885 (N_22885,N_21488,N_20206);
or U22886 (N_22886,N_20892,N_20438);
nor U22887 (N_22887,N_21350,N_20209);
or U22888 (N_22888,N_22350,N_20345);
and U22889 (N_22889,N_22212,N_21583);
or U22890 (N_22890,N_22217,N_20649);
xor U22891 (N_22891,N_20488,N_21985);
xnor U22892 (N_22892,N_20249,N_21819);
or U22893 (N_22893,N_21254,N_22465);
nor U22894 (N_22894,N_22460,N_21993);
nor U22895 (N_22895,N_21124,N_20361);
xor U22896 (N_22896,N_21320,N_20727);
or U22897 (N_22897,N_22244,N_21544);
or U22898 (N_22898,N_21103,N_22027);
or U22899 (N_22899,N_22089,N_20621);
or U22900 (N_22900,N_20451,N_21920);
xnor U22901 (N_22901,N_22229,N_21094);
nor U22902 (N_22902,N_20261,N_21905);
xnor U22903 (N_22903,N_21213,N_20470);
and U22904 (N_22904,N_21267,N_21773);
or U22905 (N_22905,N_22077,N_22167);
xnor U22906 (N_22906,N_21046,N_22005);
nand U22907 (N_22907,N_21800,N_20238);
nor U22908 (N_22908,N_21626,N_22218);
and U22909 (N_22909,N_21266,N_21225);
and U22910 (N_22910,N_22384,N_22238);
or U22911 (N_22911,N_20851,N_20340);
xnor U22912 (N_22912,N_22372,N_21958);
and U22913 (N_22913,N_21344,N_21361);
nand U22914 (N_22914,N_20375,N_20389);
nor U22915 (N_22915,N_20058,N_20846);
nand U22916 (N_22916,N_21421,N_21251);
and U22917 (N_22917,N_22196,N_20453);
and U22918 (N_22918,N_20237,N_20471);
xor U22919 (N_22919,N_22094,N_20452);
nor U22920 (N_22920,N_22099,N_21982);
xnor U22921 (N_22921,N_21901,N_20107);
xor U22922 (N_22922,N_21163,N_22058);
nor U22923 (N_22923,N_22023,N_21457);
and U22924 (N_22924,N_21902,N_21963);
nor U22925 (N_22925,N_20234,N_21765);
nand U22926 (N_22926,N_21298,N_21217);
xor U22927 (N_22927,N_20318,N_20572);
nor U22928 (N_22928,N_22396,N_22414);
nor U22929 (N_22929,N_21269,N_21941);
or U22930 (N_22930,N_22427,N_20704);
nor U22931 (N_22931,N_21194,N_21704);
nand U22932 (N_22932,N_20840,N_21293);
nor U22933 (N_22933,N_22035,N_20714);
or U22934 (N_22934,N_21121,N_20966);
or U22935 (N_22935,N_20773,N_20410);
nand U22936 (N_22936,N_22390,N_21065);
or U22937 (N_22937,N_22443,N_22098);
and U22938 (N_22938,N_22185,N_22113);
and U22939 (N_22939,N_22137,N_21138);
nor U22940 (N_22940,N_20677,N_22448);
nand U22941 (N_22941,N_22420,N_22004);
nor U22942 (N_22942,N_21711,N_22202);
or U22943 (N_22943,N_21179,N_21822);
nand U22944 (N_22944,N_20289,N_22261);
or U22945 (N_22945,N_20446,N_20416);
or U22946 (N_22946,N_20949,N_21412);
nand U22947 (N_22947,N_20290,N_21047);
nand U22948 (N_22948,N_20898,N_21756);
xor U22949 (N_22949,N_20641,N_22087);
and U22950 (N_22950,N_22345,N_22184);
and U22951 (N_22951,N_20477,N_21422);
and U22952 (N_22952,N_20423,N_20355);
nand U22953 (N_22953,N_21964,N_22221);
nand U22954 (N_22954,N_21080,N_20521);
and U22955 (N_22955,N_21913,N_21162);
and U22956 (N_22956,N_20441,N_21836);
and U22957 (N_22957,N_20137,N_21268);
nor U22958 (N_22958,N_20469,N_20300);
nor U22959 (N_22959,N_20988,N_22356);
xor U22960 (N_22960,N_21990,N_21280);
nand U22961 (N_22961,N_21108,N_20106);
xnor U22962 (N_22962,N_20963,N_21505);
xnor U22963 (N_22963,N_21168,N_22265);
xnor U22964 (N_22964,N_21043,N_22352);
or U22965 (N_22965,N_20894,N_20983);
nand U22966 (N_22966,N_20192,N_20506);
and U22967 (N_22967,N_20805,N_22179);
xnor U22968 (N_22968,N_21580,N_21524);
nor U22969 (N_22969,N_22020,N_21154);
and U22970 (N_22970,N_22170,N_21584);
or U22971 (N_22971,N_22480,N_21117);
nor U22972 (N_22972,N_22226,N_21279);
nor U22973 (N_22973,N_20336,N_21879);
nor U22974 (N_22974,N_20084,N_20958);
nor U22975 (N_22975,N_22171,N_20939);
nand U22976 (N_22976,N_21397,N_21209);
nor U22977 (N_22977,N_20591,N_22129);
nor U22978 (N_22978,N_21852,N_20351);
nand U22979 (N_22979,N_21778,N_20113);
xor U22980 (N_22980,N_20147,N_20491);
or U22981 (N_22981,N_22241,N_21362);
nor U22982 (N_22982,N_21774,N_21082);
nand U22983 (N_22983,N_21724,N_22338);
nor U22984 (N_22984,N_21338,N_20064);
or U22985 (N_22985,N_22239,N_21666);
and U22986 (N_22986,N_21402,N_21857);
nor U22987 (N_22987,N_20529,N_20891);
or U22988 (N_22988,N_20770,N_21893);
and U22989 (N_22989,N_21187,N_21480);
nand U22990 (N_22990,N_21712,N_20751);
nand U22991 (N_22991,N_22160,N_20420);
or U22992 (N_22992,N_20184,N_20740);
nand U22993 (N_22993,N_20476,N_22280);
nand U22994 (N_22994,N_20785,N_20836);
xnor U22995 (N_22995,N_21923,N_20652);
nand U22996 (N_22996,N_20034,N_21789);
nand U22997 (N_22997,N_22457,N_20905);
and U22998 (N_22998,N_21987,N_21829);
xnor U22999 (N_22999,N_21689,N_20671);
or U23000 (N_23000,N_20731,N_21038);
or U23001 (N_23001,N_21186,N_21977);
or U23002 (N_23002,N_21788,N_21409);
or U23003 (N_23003,N_22445,N_21383);
nor U23004 (N_23004,N_20930,N_21687);
or U23005 (N_23005,N_20304,N_21473);
and U23006 (N_23006,N_21211,N_20339);
and U23007 (N_23007,N_21311,N_21966);
nor U23008 (N_23008,N_20538,N_22123);
xnor U23009 (N_23009,N_22131,N_20600);
and U23010 (N_23010,N_20473,N_22335);
nand U23011 (N_23011,N_21546,N_21003);
or U23012 (N_23012,N_21051,N_22343);
nor U23013 (N_23013,N_22486,N_21675);
and U23014 (N_23014,N_21243,N_22141);
xor U23015 (N_23015,N_20664,N_21129);
or U23016 (N_23016,N_20286,N_20931);
or U23017 (N_23017,N_21739,N_21265);
or U23018 (N_23018,N_20161,N_20172);
or U23019 (N_23019,N_20808,N_21939);
nand U23020 (N_23020,N_22164,N_20203);
and U23021 (N_23021,N_22190,N_21426);
or U23022 (N_23022,N_22311,N_21511);
and U23023 (N_23023,N_20676,N_20748);
or U23024 (N_23024,N_21592,N_22353);
nor U23025 (N_23025,N_21844,N_21246);
xnor U23026 (N_23026,N_21221,N_22091);
or U23027 (N_23027,N_21936,N_20879);
xor U23028 (N_23028,N_22455,N_21808);
nand U23029 (N_23029,N_22032,N_21628);
xnor U23030 (N_23030,N_21543,N_22153);
or U23031 (N_23031,N_22294,N_20833);
nand U23032 (N_23032,N_20000,N_21871);
or U23033 (N_23033,N_20571,N_21090);
xnor U23034 (N_23034,N_22333,N_21067);
or U23035 (N_23035,N_20094,N_20370);
or U23036 (N_23036,N_21860,N_21954);
nand U23037 (N_23037,N_21853,N_20077);
or U23038 (N_23038,N_20753,N_21832);
xor U23039 (N_23039,N_21542,N_20990);
xnor U23040 (N_23040,N_21450,N_22081);
or U23041 (N_23041,N_21337,N_21757);
nor U23042 (N_23042,N_22288,N_21695);
nor U23043 (N_23043,N_21821,N_20887);
and U23044 (N_23044,N_21288,N_20018);
nand U23045 (N_23045,N_21438,N_22195);
or U23046 (N_23046,N_20126,N_20614);
or U23047 (N_23047,N_20100,N_21109);
xnor U23048 (N_23048,N_20449,N_20194);
xnor U23049 (N_23049,N_20354,N_21890);
and U23050 (N_23050,N_21520,N_21818);
xnor U23051 (N_23051,N_21032,N_22092);
xor U23052 (N_23052,N_21882,N_21351);
and U23053 (N_23053,N_22078,N_22479);
xor U23054 (N_23054,N_22357,N_21813);
or U23055 (N_23055,N_20982,N_20514);
nor U23056 (N_23056,N_21921,N_21917);
nor U23057 (N_23057,N_21594,N_20153);
xor U23058 (N_23058,N_20231,N_21453);
nand U23059 (N_23059,N_21411,N_20131);
nor U23060 (N_23060,N_22406,N_21621);
xor U23061 (N_23061,N_21181,N_21468);
and U23062 (N_23062,N_22273,N_21753);
nor U23063 (N_23063,N_21486,N_20041);
nand U23064 (N_23064,N_22104,N_21202);
or U23065 (N_23065,N_20594,N_20665);
or U23066 (N_23066,N_20640,N_20101);
and U23067 (N_23067,N_20133,N_21433);
xor U23068 (N_23068,N_20232,N_21553);
nand U23069 (N_23069,N_20325,N_20362);
and U23070 (N_23070,N_20533,N_21806);
or U23071 (N_23071,N_20242,N_20448);
nand U23072 (N_23072,N_22174,N_20177);
nand U23073 (N_23073,N_20328,N_21176);
xnor U23074 (N_23074,N_20136,N_20248);
or U23075 (N_23075,N_20143,N_22158);
and U23076 (N_23076,N_21837,N_20950);
and U23077 (N_23077,N_22469,N_20822);
and U23078 (N_23078,N_20015,N_22130);
or U23079 (N_23079,N_20109,N_21582);
and U23080 (N_23080,N_22019,N_22220);
and U23081 (N_23081,N_22456,N_20651);
xor U23082 (N_23082,N_20792,N_21374);
nor U23083 (N_23083,N_22143,N_20265);
xnor U23084 (N_23084,N_20828,N_21200);
and U23085 (N_23085,N_20275,N_20739);
nand U23086 (N_23086,N_21114,N_21215);
or U23087 (N_23087,N_21008,N_20484);
nor U23088 (N_23088,N_21545,N_20413);
nand U23089 (N_23089,N_20804,N_21903);
or U23090 (N_23090,N_21647,N_21799);
and U23091 (N_23091,N_21083,N_21976);
nor U23092 (N_23092,N_20719,N_22370);
nor U23093 (N_23093,N_20024,N_21731);
nand U23094 (N_23094,N_20050,N_22251);
nand U23095 (N_23095,N_22322,N_21366);
xnor U23096 (N_23096,N_22101,N_20115);
xnor U23097 (N_23097,N_21353,N_22371);
xnor U23098 (N_23098,N_21887,N_22334);
nor U23099 (N_23099,N_20124,N_22292);
nand U23100 (N_23100,N_20803,N_22145);
nand U23101 (N_23101,N_20977,N_20178);
or U23102 (N_23102,N_21002,N_22139);
and U23103 (N_23103,N_21708,N_20620);
nand U23104 (N_23104,N_22286,N_21846);
or U23105 (N_23105,N_21700,N_20246);
nor U23106 (N_23106,N_21390,N_21881);
nand U23107 (N_23107,N_20784,N_21380);
nand U23108 (N_23108,N_20314,N_20648);
and U23109 (N_23109,N_20800,N_20281);
or U23110 (N_23110,N_21400,N_20095);
xnor U23111 (N_23111,N_21497,N_21649);
nor U23112 (N_23112,N_20165,N_21489);
or U23113 (N_23113,N_21195,N_21481);
nor U23114 (N_23114,N_20399,N_21054);
xor U23115 (N_23115,N_21817,N_22316);
xnor U23116 (N_23116,N_22249,N_21456);
nor U23117 (N_23117,N_21287,N_21336);
and U23118 (N_23118,N_20888,N_20730);
nand U23119 (N_23119,N_20555,N_21347);
nor U23120 (N_23120,N_21979,N_21328);
or U23121 (N_23121,N_22279,N_21441);
or U23122 (N_23122,N_21597,N_21926);
nor U23123 (N_23123,N_20862,N_20302);
or U23124 (N_23124,N_20689,N_21692);
xor U23125 (N_23125,N_20741,N_20612);
nor U23126 (N_23126,N_20551,N_22169);
nor U23127 (N_23127,N_22433,N_20734);
nand U23128 (N_23128,N_20097,N_20224);
nor U23129 (N_23129,N_22007,N_20144);
nor U23130 (N_23130,N_20890,N_22055);
xnor U23131 (N_23131,N_21965,N_21716);
or U23132 (N_23132,N_20599,N_20938);
or U23133 (N_23133,N_20516,N_21242);
or U23134 (N_23134,N_21681,N_20392);
and U23135 (N_23135,N_21113,N_21218);
nand U23136 (N_23136,N_21504,N_20959);
nand U23137 (N_23137,N_21555,N_21220);
nand U23138 (N_23138,N_21041,N_20666);
nor U23139 (N_23139,N_21062,N_21136);
and U23140 (N_23140,N_20356,N_21276);
nand U23141 (N_23141,N_21950,N_21644);
nor U23142 (N_23142,N_22319,N_21172);
nand U23143 (N_23143,N_21698,N_21931);
or U23144 (N_23144,N_21749,N_20486);
and U23145 (N_23145,N_22022,N_20953);
nor U23146 (N_23146,N_21648,N_20183);
nor U23147 (N_23147,N_22441,N_20998);
xnor U23148 (N_23148,N_22086,N_22199);
and U23149 (N_23149,N_20504,N_21030);
nand U23150 (N_23150,N_20067,N_22041);
nand U23151 (N_23151,N_21750,N_21878);
xor U23152 (N_23152,N_20896,N_20615);
nor U23153 (N_23153,N_21376,N_21143);
nor U23154 (N_23154,N_21631,N_20287);
and U23155 (N_23155,N_21308,N_21640);
xor U23156 (N_23156,N_20433,N_21657);
nand U23157 (N_23157,N_22042,N_20964);
nand U23158 (N_23158,N_20725,N_21781);
nand U23159 (N_23159,N_21037,N_22367);
xor U23160 (N_23160,N_21984,N_20029);
and U23161 (N_23161,N_20241,N_21975);
nand U23162 (N_23162,N_21029,N_21378);
or U23163 (N_23163,N_21462,N_20960);
nor U23164 (N_23164,N_20481,N_21305);
xnor U23165 (N_23165,N_21107,N_21733);
xor U23166 (N_23166,N_22461,N_22491);
nand U23167 (N_23167,N_20700,N_21233);
nor U23168 (N_23168,N_22254,N_20524);
xor U23169 (N_23169,N_20341,N_20487);
nand U23170 (N_23170,N_20282,N_20945);
nor U23171 (N_23171,N_21100,N_20532);
nor U23172 (N_23172,N_20479,N_20684);
or U23173 (N_23173,N_20750,N_20215);
or U23174 (N_23174,N_20913,N_20764);
or U23175 (N_23175,N_21281,N_20235);
xnor U23176 (N_23176,N_21178,N_20408);
nand U23177 (N_23177,N_20151,N_20014);
nand U23178 (N_23178,N_22234,N_20815);
nand U23179 (N_23179,N_21284,N_20668);
or U23180 (N_23180,N_21969,N_21074);
and U23181 (N_23181,N_21637,N_20272);
xnor U23182 (N_23182,N_20274,N_20157);
nand U23183 (N_23183,N_21304,N_22494);
and U23184 (N_23184,N_21061,N_22379);
xnor U23185 (N_23185,N_20756,N_20775);
and U23186 (N_23186,N_20139,N_22237);
xnor U23187 (N_23187,N_20712,N_20858);
nand U23188 (N_23188,N_22016,N_20013);
and U23189 (N_23189,N_20779,N_21391);
xor U23190 (N_23190,N_21261,N_22262);
nor U23191 (N_23191,N_21554,N_21367);
and U23192 (N_23192,N_21718,N_20353);
or U23193 (N_23193,N_21290,N_20211);
and U23194 (N_23194,N_21630,N_21875);
xor U23195 (N_23195,N_21945,N_21767);
nor U23196 (N_23196,N_21654,N_21636);
or U23197 (N_23197,N_20293,N_21024);
nor U23198 (N_23198,N_20117,N_21764);
nand U23199 (N_23199,N_21034,N_22147);
xnor U23200 (N_23200,N_20985,N_21703);
or U23201 (N_23201,N_21498,N_20655);
nor U23202 (N_23202,N_21615,N_22152);
and U23203 (N_23203,N_20240,N_21439);
nor U23204 (N_23204,N_21547,N_20023);
and U23205 (N_23205,N_20401,N_21670);
nor U23206 (N_23206,N_22375,N_22284);
nor U23207 (N_23207,N_20443,N_22387);
nand U23208 (N_23208,N_20033,N_21701);
nand U23209 (N_23209,N_21629,N_22310);
or U23210 (N_23210,N_22096,N_20991);
xnor U23211 (N_23211,N_20724,N_21048);
nand U23212 (N_23212,N_21495,N_21424);
nand U23213 (N_23213,N_21023,N_22100);
and U23214 (N_23214,N_21310,N_21790);
or U23215 (N_23215,N_21601,N_21558);
xnor U23216 (N_23216,N_21794,N_20758);
xor U23217 (N_23217,N_20877,N_21004);
xor U23218 (N_23218,N_21540,N_21651);
and U23219 (N_23219,N_20220,N_22363);
nor U23220 (N_23220,N_21610,N_21300);
xnor U23221 (N_23221,N_21529,N_20439);
and U23222 (N_23222,N_22222,N_21184);
or U23223 (N_23223,N_21622,N_21249);
nand U23224 (N_23224,N_20283,N_20037);
xor U23225 (N_23225,N_21616,N_20425);
nand U23226 (N_23226,N_21087,N_20718);
xor U23227 (N_23227,N_20170,N_22250);
and U23228 (N_23228,N_21900,N_21981);
and U23229 (N_23229,N_22090,N_20434);
nor U23230 (N_23230,N_20961,N_20645);
xnor U23231 (N_23231,N_20497,N_20849);
or U23232 (N_23232,N_22450,N_20088);
nor U23233 (N_23233,N_22116,N_20474);
nor U23234 (N_23234,N_20587,N_20698);
or U23235 (N_23235,N_20839,N_21232);
xnor U23236 (N_23236,N_20911,N_21227);
and U23237 (N_23237,N_20418,N_21793);
or U23238 (N_23238,N_21899,N_20636);
nand U23239 (N_23239,N_22205,N_22186);
and U23240 (N_23240,N_21330,N_22269);
nor U23241 (N_23241,N_21196,N_20541);
nand U23242 (N_23242,N_20129,N_20576);
or U23243 (N_23243,N_20030,N_20028);
or U23244 (N_23244,N_21686,N_21206);
nand U23245 (N_23245,N_22211,N_21957);
nor U23246 (N_23246,N_20195,N_20659);
xnor U23247 (N_23247,N_22484,N_22033);
and U23248 (N_23248,N_21185,N_21127);
nand U23249 (N_23249,N_20589,N_21443);
and U23250 (N_23250,N_20331,N_20142);
or U23251 (N_23251,N_22134,N_21577);
or U23252 (N_23252,N_21384,N_20301);
nor U23253 (N_23253,N_20391,N_22386);
and U23254 (N_23254,N_20537,N_21859);
xnor U23255 (N_23255,N_20022,N_22493);
xor U23256 (N_23256,N_21527,N_21472);
xor U23257 (N_23257,N_22259,N_21190);
and U23258 (N_23258,N_21193,N_20295);
nand U23259 (N_23259,N_20182,N_20933);
nand U23260 (N_23260,N_21953,N_21595);
and U23261 (N_23261,N_21203,N_21776);
nor U23262 (N_23262,N_21145,N_20581);
nand U23263 (N_23263,N_21886,N_20667);
and U23264 (N_23264,N_22127,N_21420);
nand U23265 (N_23265,N_22495,N_22421);
and U23266 (N_23266,N_21918,N_20288);
or U23267 (N_23267,N_21538,N_20440);
nor U23268 (N_23268,N_22031,N_21253);
nand U23269 (N_23269,N_20653,N_21624);
xor U23270 (N_23270,N_20673,N_21797);
or U23271 (N_23271,N_20006,N_20052);
or U23272 (N_23272,N_20638,N_20853);
xnor U23273 (N_23273,N_21798,N_20880);
and U23274 (N_23274,N_21160,N_20929);
or U23275 (N_23275,N_21245,N_20883);
and U23276 (N_23276,N_22366,N_20654);
nand U23277 (N_23277,N_21635,N_21357);
xnor U23278 (N_23278,N_22355,N_21643);
or U23279 (N_23279,N_21568,N_21198);
nor U23280 (N_23280,N_21892,N_21705);
xnor U23281 (N_23281,N_20197,N_20061);
and U23282 (N_23282,N_20691,N_20848);
nor U23283 (N_23283,N_21578,N_20707);
nor U23284 (N_23284,N_22478,N_20527);
or U23285 (N_23285,N_21052,N_20921);
xnor U23286 (N_23286,N_21709,N_20674);
nor U23287 (N_23287,N_22069,N_21407);
nand U23288 (N_23288,N_20292,N_21095);
and U23289 (N_23289,N_20508,N_21552);
or U23290 (N_23290,N_20063,N_21590);
nor U23291 (N_23291,N_22204,N_21086);
or U23292 (N_23292,N_21551,N_21650);
or U23293 (N_23293,N_21891,N_22245);
nor U23294 (N_23294,N_21294,N_21388);
and U23295 (N_23295,N_20768,N_22317);
nor U23296 (N_23296,N_20327,N_21664);
nor U23297 (N_23297,N_21360,N_22291);
nand U23298 (N_23298,N_21801,N_20442);
and U23299 (N_23299,N_21842,N_22208);
and U23300 (N_23300,N_21183,N_22392);
xnor U23301 (N_23301,N_20837,N_20204);
nor U23302 (N_23302,N_21156,N_21098);
nand U23303 (N_23303,N_21988,N_20069);
nor U23304 (N_23304,N_21333,N_20498);
or U23305 (N_23305,N_20510,N_20834);
nand U23306 (N_23306,N_21073,N_21502);
or U23307 (N_23307,N_22385,N_20616);
xnor U23308 (N_23308,N_20447,N_21216);
or U23309 (N_23309,N_20925,N_21394);
nor U23310 (N_23310,N_20584,N_22389);
nand U23311 (N_23311,N_21668,N_21079);
xor U23312 (N_23312,N_22013,N_20745);
nor U23313 (N_23313,N_20951,N_21446);
nand U23314 (N_23314,N_22309,N_22413);
and U23315 (N_23315,N_21039,N_21717);
xnor U23316 (N_23316,N_21754,N_20430);
and U23317 (N_23317,N_22436,N_20914);
nor U23318 (N_23318,N_20244,N_20239);
and U23319 (N_23319,N_21170,N_22246);
xor U23320 (N_23320,N_20081,N_20444);
or U23321 (N_23321,N_20012,N_20760);
or U23322 (N_23322,N_20379,N_20186);
and U23323 (N_23323,N_20956,N_21779);
and U23324 (N_23324,N_22103,N_21758);
nor U23325 (N_23325,N_21214,N_20733);
nand U23326 (N_23326,N_21834,N_20475);
or U23327 (N_23327,N_21155,N_21352);
nor U23328 (N_23328,N_21605,N_21139);
nand U23329 (N_23329,N_20520,N_21372);
and U23330 (N_23330,N_20787,N_22489);
xnor U23331 (N_23331,N_21576,N_21761);
nor U23332 (N_23332,N_20575,N_20952);
nor U23333 (N_23333,N_22312,N_20847);
nor U23334 (N_23334,N_21452,N_21334);
nand U23335 (N_23335,N_22108,N_21197);
nand U23336 (N_23336,N_20618,N_20780);
xnor U23337 (N_23337,N_21060,N_20159);
nor U23338 (N_23338,N_21745,N_20495);
nor U23339 (N_23339,N_21159,N_22155);
nand U23340 (N_23340,N_21063,N_20087);
or U23341 (N_23341,N_20854,N_21748);
and U23342 (N_23342,N_20335,N_20954);
or U23343 (N_23343,N_21503,N_21377);
nand U23344 (N_23344,N_21600,N_22416);
nand U23345 (N_23345,N_21980,N_21466);
and U23346 (N_23346,N_21332,N_21478);
or U23347 (N_23347,N_21561,N_21683);
nand U23348 (N_23348,N_20216,N_20974);
nor U23349 (N_23349,N_22409,N_21530);
and U23350 (N_23350,N_22209,N_21427);
xor U23351 (N_23351,N_20906,N_22342);
or U23352 (N_23352,N_21031,N_20765);
or U23353 (N_23353,N_22302,N_22422);
and U23354 (N_23354,N_21588,N_21092);
nand U23355 (N_23355,N_20909,N_20450);
nand U23356 (N_23356,N_20511,N_20672);
or U23357 (N_23357,N_22181,N_22474);
nand U23358 (N_23358,N_21317,N_22176);
or U23359 (N_23359,N_20560,N_22419);
nor U23360 (N_23360,N_20236,N_20419);
xnor U23361 (N_23361,N_20053,N_22107);
nor U23362 (N_23362,N_20578,N_21611);
nand U23363 (N_23363,N_21099,N_20346);
nor U23364 (N_23364,N_21519,N_20269);
nor U23365 (N_23365,N_21937,N_21009);
or U23366 (N_23366,N_20927,N_21315);
and U23367 (N_23367,N_20611,N_20969);
xnor U23368 (N_23368,N_21398,N_21952);
nand U23369 (N_23369,N_20749,N_20243);
xnor U23370 (N_23370,N_22097,N_20382);
nor U23371 (N_23371,N_22111,N_21483);
and U23372 (N_23372,N_21102,N_21252);
and U23373 (N_23373,N_21123,N_21479);
xor U23374 (N_23374,N_20214,N_21339);
xnor U23375 (N_23375,N_20922,N_22417);
and U23376 (N_23376,N_21370,N_21223);
and U23377 (N_23377,N_20073,N_22084);
nand U23378 (N_23378,N_21110,N_20918);
and U23379 (N_23379,N_20317,N_21494);
nand U23380 (N_23380,N_20011,N_21924);
nand U23381 (N_23381,N_21760,N_21688);
or U23382 (N_23382,N_21104,N_22477);
or U23383 (N_23383,N_21140,N_21574);
or U23384 (N_23384,N_21707,N_21318);
xnor U23385 (N_23385,N_21840,N_21499);
nand U23386 (N_23386,N_20878,N_22327);
nand U23387 (N_23387,N_21885,N_20366);
xnor U23388 (N_23388,N_20628,N_21207);
xor U23389 (N_23389,N_20093,N_20020);
and U23390 (N_23390,N_22198,N_21161);
xnor U23391 (N_23391,N_21855,N_21956);
nor U23392 (N_23392,N_20155,N_22082);
nand U23393 (N_23393,N_22483,N_21027);
xnor U23394 (N_23394,N_21934,N_21131);
nand U23395 (N_23395,N_20492,N_20227);
nand U23396 (N_23396,N_21608,N_22328);
nand U23397 (N_23397,N_20169,N_21146);
and U23398 (N_23398,N_22002,N_21055);
nor U23399 (N_23399,N_21641,N_22183);
xor U23400 (N_23400,N_22182,N_21312);
nor U23401 (N_23401,N_21147,N_21780);
xnor U23402 (N_23402,N_20526,N_20549);
xor U23403 (N_23403,N_21258,N_20876);
xnor U23404 (N_23404,N_21514,N_20686);
or U23405 (N_23405,N_22440,N_20893);
nand U23406 (N_23406,N_22397,N_21967);
or U23407 (N_23407,N_21295,N_22256);
xnor U23408 (N_23408,N_21572,N_20515);
nand U23409 (N_23409,N_21625,N_22138);
nor U23410 (N_23410,N_21727,N_21560);
nand U23411 (N_23411,N_20842,N_20112);
nor U23412 (N_23412,N_22136,N_20198);
and U23413 (N_23413,N_21064,N_21158);
nor U23414 (N_23414,N_20503,N_20207);
nor U23415 (N_23415,N_20981,N_21828);
or U23416 (N_23416,N_21607,N_21416);
or U23417 (N_23417,N_21912,N_22313);
and U23418 (N_23418,N_21827,N_20818);
nand U23419 (N_23419,N_20262,N_21904);
or U23420 (N_23420,N_21884,N_21142);
nand U23421 (N_23421,N_20901,N_21522);
nand U23422 (N_23422,N_21297,N_20415);
nor U23423 (N_23423,N_21674,N_22072);
nor U23424 (N_23424,N_21581,N_21219);
or U23425 (N_23425,N_21057,N_20467);
nor U23426 (N_23426,N_20831,N_20310);
xor U23427 (N_23427,N_20188,N_22052);
nor U23428 (N_23428,N_20043,N_21049);
nand U23429 (N_23429,N_20278,N_21035);
nor U23430 (N_23430,N_20435,N_22287);
nor U23431 (N_23431,N_20732,N_20811);
or U23432 (N_23432,N_21509,N_20688);
nand U23433 (N_23433,N_21224,N_21662);
and U23434 (N_23434,N_20298,N_20160);
nand U23435 (N_23435,N_22060,N_21723);
nand U23436 (N_23436,N_21876,N_21944);
nor U23437 (N_23437,N_21282,N_21661);
xnor U23438 (N_23438,N_21833,N_20996);
xor U23439 (N_23439,N_21972,N_21272);
xor U23440 (N_23440,N_21943,N_21839);
nand U23441 (N_23441,N_22289,N_21240);
nor U23442 (N_23442,N_22418,N_21777);
nor U23443 (N_23443,N_22177,N_20145);
and U23444 (N_23444,N_21676,N_22148);
or U23445 (N_23445,N_22144,N_21078);
xnor U23446 (N_23446,N_22119,N_21658);
or U23447 (N_23447,N_20886,N_22361);
or U23448 (N_23448,N_21596,N_21093);
or U23449 (N_23449,N_20816,N_20604);
or U23450 (N_23450,N_20367,N_22394);
or U23451 (N_23451,N_21348,N_21786);
nor U23452 (N_23452,N_20596,N_22043);
xnor U23453 (N_23453,N_20173,N_22068);
and U23454 (N_23454,N_21449,N_22431);
nor U23455 (N_23455,N_20390,N_22304);
and U23456 (N_23456,N_21012,N_22308);
and U23457 (N_23457,N_22321,N_22253);
nand U23458 (N_23458,N_20743,N_20536);
or U23459 (N_23459,N_21363,N_21565);
xor U23460 (N_23460,N_20801,N_20819);
or U23461 (N_23461,N_20633,N_21270);
xnor U23462 (N_23462,N_20683,N_20460);
xor U23463 (N_23463,N_21171,N_21231);
xnor U23464 (N_23464,N_22408,N_20008);
or U23465 (N_23465,N_22021,N_22240);
nor U23466 (N_23466,N_21259,N_20060);
nor U23467 (N_23467,N_20694,N_20493);
xor U23468 (N_23468,N_20500,N_21639);
and U23469 (N_23469,N_21632,N_22283);
and U23470 (N_23470,N_20910,N_20003);
or U23471 (N_23471,N_22497,N_20919);
nor U23472 (N_23472,N_21386,N_22120);
and U23473 (N_23473,N_20102,N_20902);
or U23474 (N_23474,N_20316,N_21464);
xnor U23475 (N_23475,N_21492,N_21638);
and U23476 (N_23476,N_21646,N_20681);
xor U23477 (N_23477,N_22200,N_21118);
nor U23478 (N_23478,N_21623,N_20588);
xor U23479 (N_23479,N_22266,N_20202);
and U23480 (N_23480,N_21292,N_20250);
xor U23481 (N_23481,N_20068,N_20820);
nand U23482 (N_23482,N_20937,N_20795);
and U23483 (N_23483,N_22073,N_20344);
nand U23484 (N_23484,N_20127,N_21250);
nand U23485 (N_23485,N_20736,N_20309);
nand U23486 (N_23486,N_21679,N_21068);
nand U23487 (N_23487,N_20337,N_20096);
and U23488 (N_23488,N_21521,N_21346);
or U23489 (N_23489,N_21469,N_22121);
nor U23490 (N_23490,N_21500,N_21627);
nand U23491 (N_23491,N_20944,N_20409);
and U23492 (N_23492,N_21771,N_20675);
nor U23493 (N_23493,N_20429,N_21669);
nor U23494 (N_23494,N_22168,N_22481);
nor U23495 (N_23495,N_20221,N_21326);
nor U23496 (N_23496,N_20554,N_21645);
or U23497 (N_23497,N_20957,N_22260);
xor U23498 (N_23498,N_21302,N_21105);
nand U23499 (N_23499,N_20110,N_20762);
xnor U23500 (N_23500,N_22485,N_20832);
and U23501 (N_23501,N_22415,N_22488);
nor U23502 (N_23502,N_21482,N_21014);
or U23503 (N_23503,N_21408,N_21434);
nor U23504 (N_23504,N_21465,N_20830);
nor U23505 (N_23505,N_20187,N_20627);
and U23506 (N_23506,N_20368,N_20417);
or U23507 (N_23507,N_20255,N_20163);
nand U23508 (N_23508,N_22178,N_22106);
nand U23509 (N_23509,N_21418,N_21119);
xnor U23510 (N_23510,N_22175,N_20569);
xnor U23511 (N_23511,N_21946,N_20412);
nand U23512 (N_23512,N_21122,N_21327);
nor U23513 (N_23513,N_21866,N_22223);
and U23514 (N_23514,N_20687,N_21467);
or U23515 (N_23515,N_22225,N_20454);
xnor U23516 (N_23516,N_20267,N_20573);
or U23517 (N_23517,N_20755,N_21340);
nand U23518 (N_23518,N_20726,N_21277);
xnor U23519 (N_23519,N_21783,N_21744);
nor U23520 (N_23520,N_21026,N_20874);
nand U23521 (N_23521,N_21015,N_20546);
xnor U23522 (N_23522,N_21541,N_21071);
and U23523 (N_23523,N_22000,N_21694);
xor U23524 (N_23524,N_21831,N_21120);
or U23525 (N_23525,N_20277,N_22399);
nand U23526 (N_23526,N_21275,N_20038);
xor U23527 (N_23527,N_20056,N_22124);
and U23528 (N_23528,N_20321,N_20263);
xnor U23529 (N_23529,N_20372,N_21134);
and U23530 (N_23530,N_20071,N_20128);
or U23531 (N_23531,N_22018,N_21820);
nor U23532 (N_23532,N_21239,N_22339);
nand U23533 (N_23533,N_20993,N_20577);
nor U23534 (N_23534,N_20374,N_22452);
nand U23535 (N_23535,N_20009,N_20669);
nor U23536 (N_23536,N_20154,N_20284);
and U23537 (N_23537,N_21851,N_22347);
and U23538 (N_23538,N_20783,N_21873);
xor U23539 (N_23539,N_20513,N_20384);
xor U23540 (N_23540,N_22114,N_20738);
and U23541 (N_23541,N_21537,N_20251);
xnor U23542 (N_23542,N_20643,N_20852);
and U23543 (N_23543,N_20294,N_21423);
nand U23544 (N_23544,N_21306,N_20602);
and U23545 (N_23545,N_20496,N_22207);
and U23546 (N_23546,N_21454,N_20065);
or U23547 (N_23547,N_20946,N_21368);
nor U23548 (N_23548,N_20658,N_21444);
nand U23549 (N_23549,N_20342,N_20821);
nor U23550 (N_23550,N_20230,N_20472);
nor U23551 (N_23551,N_22037,N_20431);
and U23552 (N_23552,N_20402,N_21802);
nor U23553 (N_23553,N_21013,N_22303);
xnor U23554 (N_23554,N_20019,N_20268);
xnor U23555 (N_23555,N_20873,N_20558);
nand U23556 (N_23556,N_21192,N_20713);
nand U23557 (N_23557,N_20422,N_22224);
and U23558 (N_23558,N_20917,N_21137);
xor U23559 (N_23559,N_20072,N_22140);
and U23560 (N_23560,N_20972,N_21895);
xnor U23561 (N_23561,N_21732,N_21741);
nand U23562 (N_23562,N_22151,N_22065);
nor U23563 (N_23563,N_21752,N_20772);
xnor U23564 (N_23564,N_21613,N_20595);
or U23565 (N_23565,N_21737,N_20817);
xor U23566 (N_23566,N_21872,N_20559);
and U23567 (N_23567,N_21911,N_20270);
xnor U23568 (N_23568,N_20567,N_22426);
xor U23569 (N_23569,N_21069,N_21149);
or U23570 (N_23570,N_21587,N_20363);
nand U23571 (N_23571,N_21696,N_22297);
or U23572 (N_23572,N_22300,N_20343);
nand U23573 (N_23573,N_21199,N_20299);
xor U23574 (N_23574,N_20705,N_22067);
xor U23575 (N_23575,N_20984,N_21983);
xor U23576 (N_23576,N_21807,N_21111);
nor U23577 (N_23577,N_21289,N_21697);
nor U23578 (N_23578,N_22061,N_20774);
or U23579 (N_23579,N_20598,N_22173);
nor U23580 (N_23580,N_20036,N_20181);
nor U23581 (N_23581,N_20865,N_20322);
nor U23582 (N_23582,N_22163,N_20035);
and U23583 (N_23583,N_20866,N_22028);
nor U23584 (N_23584,N_20349,N_20369);
nand U23585 (N_23585,N_20796,N_21916);
nand U23586 (N_23586,N_20742,N_20702);
xor U23587 (N_23587,N_21007,N_22430);
or U23588 (N_23588,N_20044,N_21999);
xor U23589 (N_23589,N_20967,N_20226);
or U23590 (N_23590,N_20085,N_21618);
nor U23591 (N_23591,N_22365,N_20607);
nor U23592 (N_23592,N_20306,N_21883);
nor U23593 (N_23593,N_22214,N_20562);
or U23594 (N_23594,N_22437,N_20091);
nor U23595 (N_23595,N_21586,N_21720);
xnor U23596 (N_23596,N_20190,N_20899);
and U23597 (N_23597,N_21534,N_20164);
or U23598 (N_23598,N_21429,N_21766);
nand U23599 (N_23599,N_21089,N_20480);
xor U23600 (N_23600,N_21458,N_20010);
or U23601 (N_23601,N_21722,N_22381);
or U23602 (N_23602,N_20323,N_22482);
or U23603 (N_23603,N_20201,N_22146);
nand U23604 (N_23604,N_22362,N_20385);
xor U23605 (N_23605,N_21612,N_21861);
or U23606 (N_23606,N_21823,N_21841);
xnor U23607 (N_23607,N_21324,N_21059);
and U23608 (N_23608,N_22464,N_21548);
nor U23609 (N_23609,N_20357,N_22180);
nand U23610 (N_23610,N_20395,N_20276);
nand U23611 (N_23611,N_20205,N_20757);
xnor U23612 (N_23612,N_21848,N_20411);
or U23613 (N_23613,N_21325,N_20716);
or U23614 (N_23614,N_22203,N_20150);
xnor U23615 (N_23615,N_21413,N_20884);
nor U23616 (N_23616,N_20806,N_22492);
and U23617 (N_23617,N_20393,N_21128);
nand U23618 (N_23618,N_22369,N_22475);
nor U23619 (N_23619,N_20970,N_20333);
xnor U23620 (N_23620,N_22242,N_21166);
and U23621 (N_23621,N_22320,N_22064);
nor U23622 (N_23622,N_20074,N_21942);
nand U23623 (N_23623,N_21451,N_20051);
nand U23624 (N_23624,N_22281,N_20320);
nor U23625 (N_23625,N_21395,N_20388);
and U23626 (N_23626,N_21507,N_21496);
or U23627 (N_23627,N_22056,N_20692);
xnor U23628 (N_23628,N_20162,N_20347);
or U23629 (N_23629,N_21516,N_21735);
or U23630 (N_23630,N_22192,N_22470);
nor U23631 (N_23631,N_21656,N_21020);
nand U23632 (N_23632,N_20271,N_20617);
nor U23633 (N_23633,N_22412,N_21477);
and U23634 (N_23634,N_20027,N_20907);
and U23635 (N_23635,N_22466,N_20326);
xor U23636 (N_23636,N_20332,N_20540);
xnor U23637 (N_23637,N_20456,N_20920);
or U23638 (N_23638,N_20457,N_21907);
and U23639 (N_23639,N_22425,N_21208);
nand U23640 (N_23640,N_21928,N_20997);
and U23641 (N_23641,N_20583,N_21539);
nand U23642 (N_23642,N_20406,N_20928);
nor U23643 (N_23643,N_20582,N_21973);
xnor U23644 (N_23644,N_20080,N_22230);
xor U23645 (N_23645,N_20315,N_20264);
xnor U23646 (N_23646,N_22187,N_20870);
nor U23647 (N_23647,N_20693,N_20098);
or U23648 (N_23648,N_22012,N_21364);
xnor U23649 (N_23649,N_21018,N_20400);
and U23650 (N_23650,N_22487,N_21379);
and U23651 (N_23651,N_20625,N_21234);
and U23652 (N_23652,N_21204,N_21385);
or U23653 (N_23653,N_22270,N_20807);
nand U23654 (N_23654,N_21940,N_21769);
nand U23655 (N_23655,N_20501,N_20763);
nand U23656 (N_23656,N_21898,N_22150);
and U23657 (N_23657,N_20825,N_20989);
and U23658 (N_23658,N_20459,N_21684);
nor U23659 (N_23659,N_22085,N_22258);
xor U23660 (N_23660,N_21974,N_22318);
nand U23661 (N_23661,N_21736,N_21256);
nor U23662 (N_23662,N_22095,N_21768);
xor U23663 (N_23663,N_21838,N_22046);
nand U23664 (N_23664,N_22434,N_21445);
and U23665 (N_23665,N_20048,N_20212);
and U23666 (N_23666,N_21431,N_21341);
or U23667 (N_23667,N_21811,N_20463);
or U23668 (N_23668,N_21235,N_20005);
nor U23669 (N_23669,N_20955,N_21726);
or U23670 (N_23670,N_21019,N_20882);
nand U23671 (N_23671,N_21738,N_22468);
or U23672 (N_23672,N_22030,N_20590);
and U23673 (N_23673,N_20826,N_20122);
xor U23674 (N_23674,N_20260,N_21909);
nand U23675 (N_23675,N_22498,N_21476);
nor U23676 (N_23676,N_21442,N_21513);
nand U23677 (N_23677,N_20001,N_22340);
xnor U23678 (N_23678,N_21567,N_22360);
nor U23679 (N_23679,N_21933,N_20735);
and U23680 (N_23680,N_20923,N_21056);
or U23681 (N_23681,N_20218,N_22034);
and U23682 (N_23682,N_20152,N_21812);
and U23683 (N_23683,N_20123,N_20531);
and U23684 (N_23684,N_21896,N_21816);
nand U23685 (N_23685,N_21471,N_20580);
and U23686 (N_23686,N_20534,N_21742);
and U23687 (N_23687,N_20047,N_20835);
or U23688 (N_23688,N_21991,N_21845);
or U23689 (N_23689,N_20210,N_21460);
nor U23690 (N_23690,N_20771,N_20863);
nor U23691 (N_23691,N_20778,N_20812);
nand U23692 (N_23692,N_20941,N_22017);
xnor U23693 (N_23693,N_21133,N_22314);
and U23694 (N_23694,N_21342,N_21930);
xor U23695 (N_23695,N_20167,N_21803);
or U23696 (N_23696,N_20171,N_21770);
or U23697 (N_23697,N_21989,N_20550);
and U23698 (N_23698,N_22354,N_22029);
xnor U23699 (N_23699,N_21313,N_20108);
xnor U23700 (N_23700,N_22045,N_20747);
nand U23701 (N_23701,N_21652,N_22076);
or U23702 (N_23702,N_21517,N_22446);
nand U23703 (N_23703,N_21785,N_21448);
and U23704 (N_23704,N_21949,N_22210);
xnor U23705 (N_23705,N_21740,N_20405);
nor U23706 (N_23706,N_20247,N_20168);
and U23707 (N_23707,N_20258,N_21535);
nor U23708 (N_23708,N_21001,N_21747);
xnor U23709 (N_23709,N_21849,N_20855);
and U23710 (N_23710,N_21212,N_22471);
nand U23711 (N_23711,N_21682,N_20223);
or U23712 (N_23712,N_20528,N_20662);
and U23713 (N_23713,N_21699,N_20987);
nor U23714 (N_23714,N_22383,N_20296);
and U23715 (N_23715,N_21719,N_20856);
and U23716 (N_23716,N_21835,N_21660);
nor U23717 (N_23717,N_21573,N_20934);
and U23718 (N_23718,N_20543,N_20279);
nor U23719 (N_23719,N_20026,N_20062);
nor U23720 (N_23720,N_20679,N_21075);
or U23721 (N_23721,N_21175,N_21405);
and U23722 (N_23722,N_21116,N_21349);
and U23723 (N_23723,N_21759,N_20962);
nor U23724 (N_23724,N_21491,N_20146);
nand U23725 (N_23725,N_21359,N_20660);
or U23726 (N_23726,N_21309,N_22110);
or U23727 (N_23727,N_21569,N_21805);
xor U23728 (N_23728,N_20397,N_20245);
nand U23729 (N_23729,N_20737,N_20334);
and U23730 (N_23730,N_22008,N_20553);
or U23731 (N_23731,N_21782,N_22403);
and U23732 (N_23732,N_20525,N_20116);
nand U23733 (N_23733,N_21599,N_20568);
nor U23734 (N_23734,N_20565,N_21677);
or U23735 (N_23735,N_22025,N_20103);
xor U23736 (N_23736,N_21589,N_21775);
nor U23737 (N_23737,N_21130,N_20708);
nand U23738 (N_23738,N_21076,N_21951);
xnor U23739 (N_23739,N_21301,N_20105);
nor U23740 (N_23740,N_21955,N_22172);
and U23741 (N_23741,N_22337,N_21230);
nor U23742 (N_23742,N_21961,N_21070);
nor U23743 (N_23743,N_20324,N_20089);
nand U23744 (N_23744,N_22496,N_21101);
or U23745 (N_23745,N_22051,N_21863);
xor U23746 (N_23746,N_21322,N_20445);
or U23747 (N_23747,N_21490,N_20193);
or U23748 (N_23748,N_20180,N_21106);
and U23749 (N_23749,N_22348,N_22411);
xnor U23750 (N_23750,N_20108,N_21475);
nand U23751 (N_23751,N_21362,N_22256);
and U23752 (N_23752,N_21932,N_22184);
or U23753 (N_23753,N_21624,N_20555);
nand U23754 (N_23754,N_21385,N_20426);
and U23755 (N_23755,N_20448,N_21184);
xnor U23756 (N_23756,N_21758,N_21803);
xnor U23757 (N_23757,N_20848,N_21666);
and U23758 (N_23758,N_22088,N_20465);
or U23759 (N_23759,N_22292,N_20964);
nor U23760 (N_23760,N_20906,N_20258);
or U23761 (N_23761,N_20828,N_20140);
xnor U23762 (N_23762,N_22123,N_20446);
nor U23763 (N_23763,N_21986,N_21480);
or U23764 (N_23764,N_20415,N_21460);
xor U23765 (N_23765,N_20997,N_21072);
xor U23766 (N_23766,N_20213,N_22214);
nand U23767 (N_23767,N_20013,N_21594);
nand U23768 (N_23768,N_21209,N_20321);
xnor U23769 (N_23769,N_21902,N_21290);
xnor U23770 (N_23770,N_20357,N_22236);
nand U23771 (N_23771,N_21411,N_20288);
xnor U23772 (N_23772,N_21386,N_20478);
or U23773 (N_23773,N_20298,N_20171);
xor U23774 (N_23774,N_20516,N_21686);
nand U23775 (N_23775,N_21647,N_22427);
nand U23776 (N_23776,N_20090,N_22226);
and U23777 (N_23777,N_21464,N_20758);
xnor U23778 (N_23778,N_21441,N_21654);
nor U23779 (N_23779,N_20286,N_20934);
nand U23780 (N_23780,N_20737,N_20982);
and U23781 (N_23781,N_21679,N_22454);
or U23782 (N_23782,N_21387,N_22251);
nor U23783 (N_23783,N_21343,N_20876);
nand U23784 (N_23784,N_21070,N_20008);
nor U23785 (N_23785,N_21494,N_22203);
xor U23786 (N_23786,N_21436,N_21692);
or U23787 (N_23787,N_22061,N_21514);
nand U23788 (N_23788,N_21070,N_21020);
and U23789 (N_23789,N_20581,N_20372);
nand U23790 (N_23790,N_21746,N_22241);
xor U23791 (N_23791,N_21239,N_20521);
or U23792 (N_23792,N_20609,N_20908);
xnor U23793 (N_23793,N_21419,N_20809);
or U23794 (N_23794,N_22216,N_20000);
or U23795 (N_23795,N_20999,N_20928);
nor U23796 (N_23796,N_20966,N_22210);
nor U23797 (N_23797,N_20523,N_20057);
nand U23798 (N_23798,N_21590,N_22379);
or U23799 (N_23799,N_20884,N_20882);
and U23800 (N_23800,N_21722,N_22314);
xor U23801 (N_23801,N_22174,N_21887);
nor U23802 (N_23802,N_20063,N_21866);
nor U23803 (N_23803,N_21081,N_21784);
nor U23804 (N_23804,N_22454,N_20386);
and U23805 (N_23805,N_21376,N_22388);
or U23806 (N_23806,N_20278,N_21304);
nor U23807 (N_23807,N_20153,N_21641);
nand U23808 (N_23808,N_20834,N_21029);
or U23809 (N_23809,N_21850,N_20661);
nor U23810 (N_23810,N_22262,N_20121);
nor U23811 (N_23811,N_20719,N_21034);
nor U23812 (N_23812,N_20124,N_20770);
and U23813 (N_23813,N_20445,N_21876);
nand U23814 (N_23814,N_21340,N_21835);
or U23815 (N_23815,N_22298,N_21266);
or U23816 (N_23816,N_21822,N_20994);
nor U23817 (N_23817,N_21567,N_22049);
or U23818 (N_23818,N_21529,N_22376);
or U23819 (N_23819,N_22471,N_21585);
and U23820 (N_23820,N_22320,N_20540);
and U23821 (N_23821,N_21045,N_20012);
nand U23822 (N_23822,N_22237,N_21962);
xor U23823 (N_23823,N_20857,N_20882);
and U23824 (N_23824,N_20857,N_20312);
and U23825 (N_23825,N_21743,N_20006);
xor U23826 (N_23826,N_21702,N_20232);
nand U23827 (N_23827,N_22338,N_20903);
nand U23828 (N_23828,N_20181,N_20737);
xor U23829 (N_23829,N_22458,N_20237);
xor U23830 (N_23830,N_20660,N_20978);
nand U23831 (N_23831,N_20376,N_22245);
nor U23832 (N_23832,N_20732,N_20135);
or U23833 (N_23833,N_20366,N_20399);
and U23834 (N_23834,N_21130,N_21975);
or U23835 (N_23835,N_20519,N_21265);
xnor U23836 (N_23836,N_20860,N_21039);
and U23837 (N_23837,N_21566,N_22108);
nor U23838 (N_23838,N_22394,N_21011);
and U23839 (N_23839,N_20855,N_20242);
and U23840 (N_23840,N_21387,N_22157);
nor U23841 (N_23841,N_21082,N_20786);
nor U23842 (N_23842,N_20787,N_20356);
or U23843 (N_23843,N_21358,N_20142);
nand U23844 (N_23844,N_21246,N_21559);
and U23845 (N_23845,N_21220,N_20965);
nand U23846 (N_23846,N_22433,N_21167);
nand U23847 (N_23847,N_22475,N_20331);
nand U23848 (N_23848,N_22197,N_21848);
nand U23849 (N_23849,N_21260,N_20340);
nand U23850 (N_23850,N_20516,N_21571);
nor U23851 (N_23851,N_20409,N_21460);
or U23852 (N_23852,N_20810,N_21696);
nand U23853 (N_23853,N_21334,N_22451);
and U23854 (N_23854,N_20300,N_22352);
nor U23855 (N_23855,N_21935,N_21050);
xor U23856 (N_23856,N_20663,N_21864);
nand U23857 (N_23857,N_22355,N_20485);
or U23858 (N_23858,N_21775,N_21058);
or U23859 (N_23859,N_22250,N_21109);
and U23860 (N_23860,N_20184,N_20148);
nor U23861 (N_23861,N_22105,N_20531);
xnor U23862 (N_23862,N_21661,N_20137);
nand U23863 (N_23863,N_20033,N_20685);
xor U23864 (N_23864,N_21459,N_20010);
and U23865 (N_23865,N_21063,N_21181);
or U23866 (N_23866,N_21363,N_21861);
xnor U23867 (N_23867,N_21021,N_21146);
nor U23868 (N_23868,N_21257,N_22262);
nor U23869 (N_23869,N_21505,N_21356);
or U23870 (N_23870,N_21267,N_20456);
or U23871 (N_23871,N_21947,N_21191);
nand U23872 (N_23872,N_21764,N_20250);
or U23873 (N_23873,N_21832,N_20689);
nand U23874 (N_23874,N_22075,N_20119);
nand U23875 (N_23875,N_21873,N_22460);
nand U23876 (N_23876,N_22055,N_20978);
or U23877 (N_23877,N_20499,N_21909);
and U23878 (N_23878,N_22171,N_20037);
nand U23879 (N_23879,N_22104,N_20028);
and U23880 (N_23880,N_21066,N_20714);
or U23881 (N_23881,N_22330,N_22033);
xor U23882 (N_23882,N_21685,N_20401);
xor U23883 (N_23883,N_21855,N_20932);
and U23884 (N_23884,N_20937,N_20391);
nor U23885 (N_23885,N_21656,N_20422);
xor U23886 (N_23886,N_20521,N_21312);
xor U23887 (N_23887,N_20174,N_20255);
nor U23888 (N_23888,N_21367,N_21173);
and U23889 (N_23889,N_21754,N_20104);
nand U23890 (N_23890,N_20292,N_21685);
nor U23891 (N_23891,N_20738,N_22314);
nor U23892 (N_23892,N_21137,N_21797);
nor U23893 (N_23893,N_20527,N_21798);
xnor U23894 (N_23894,N_21598,N_21188);
or U23895 (N_23895,N_21778,N_21285);
or U23896 (N_23896,N_21200,N_21288);
nand U23897 (N_23897,N_22212,N_22203);
nand U23898 (N_23898,N_20201,N_21655);
and U23899 (N_23899,N_22095,N_21855);
xnor U23900 (N_23900,N_20060,N_21659);
nand U23901 (N_23901,N_21112,N_20597);
or U23902 (N_23902,N_20383,N_20327);
nor U23903 (N_23903,N_22109,N_22263);
xor U23904 (N_23904,N_21578,N_20676);
nor U23905 (N_23905,N_22426,N_20574);
xnor U23906 (N_23906,N_21312,N_21177);
nor U23907 (N_23907,N_21124,N_21389);
and U23908 (N_23908,N_20781,N_20188);
or U23909 (N_23909,N_21435,N_21930);
or U23910 (N_23910,N_21580,N_22289);
xnor U23911 (N_23911,N_20283,N_20228);
or U23912 (N_23912,N_20737,N_21973);
nor U23913 (N_23913,N_20030,N_20993);
or U23914 (N_23914,N_20235,N_21169);
nand U23915 (N_23915,N_22070,N_21876);
and U23916 (N_23916,N_20347,N_20047);
or U23917 (N_23917,N_21585,N_21354);
nor U23918 (N_23918,N_21297,N_21560);
nand U23919 (N_23919,N_20479,N_22101);
xor U23920 (N_23920,N_21527,N_21652);
nand U23921 (N_23921,N_20680,N_22179);
or U23922 (N_23922,N_20854,N_21193);
xnor U23923 (N_23923,N_21993,N_20954);
xor U23924 (N_23924,N_21674,N_20807);
nand U23925 (N_23925,N_22398,N_22444);
nor U23926 (N_23926,N_20113,N_20692);
and U23927 (N_23927,N_22019,N_20505);
or U23928 (N_23928,N_21793,N_20370);
nand U23929 (N_23929,N_21424,N_21897);
and U23930 (N_23930,N_21994,N_22332);
xnor U23931 (N_23931,N_21345,N_22362);
xor U23932 (N_23932,N_20170,N_21142);
or U23933 (N_23933,N_21486,N_22060);
xnor U23934 (N_23934,N_22166,N_22486);
nor U23935 (N_23935,N_22421,N_20986);
and U23936 (N_23936,N_20799,N_21788);
nand U23937 (N_23937,N_20860,N_22233);
or U23938 (N_23938,N_20903,N_20639);
xnor U23939 (N_23939,N_22377,N_20587);
or U23940 (N_23940,N_20623,N_22164);
xnor U23941 (N_23941,N_21809,N_20556);
nand U23942 (N_23942,N_21712,N_20602);
nor U23943 (N_23943,N_22314,N_20619);
nand U23944 (N_23944,N_20653,N_20798);
or U23945 (N_23945,N_21006,N_21120);
nor U23946 (N_23946,N_22332,N_21149);
xnor U23947 (N_23947,N_20672,N_21353);
nor U23948 (N_23948,N_22356,N_21587);
or U23949 (N_23949,N_22177,N_21460);
and U23950 (N_23950,N_22351,N_21715);
nor U23951 (N_23951,N_22045,N_22146);
and U23952 (N_23952,N_21931,N_20170);
and U23953 (N_23953,N_20663,N_20928);
xor U23954 (N_23954,N_21852,N_21927);
nor U23955 (N_23955,N_20733,N_21049);
nand U23956 (N_23956,N_20379,N_22192);
nand U23957 (N_23957,N_21677,N_21933);
or U23958 (N_23958,N_20439,N_21274);
and U23959 (N_23959,N_20559,N_20091);
nand U23960 (N_23960,N_20045,N_20875);
xor U23961 (N_23961,N_21919,N_22499);
and U23962 (N_23962,N_21434,N_21405);
or U23963 (N_23963,N_22109,N_22264);
and U23964 (N_23964,N_21688,N_20586);
xor U23965 (N_23965,N_21072,N_22074);
nand U23966 (N_23966,N_20651,N_20256);
or U23967 (N_23967,N_20745,N_22349);
nand U23968 (N_23968,N_20898,N_20058);
nand U23969 (N_23969,N_20034,N_21555);
xor U23970 (N_23970,N_21483,N_20502);
xor U23971 (N_23971,N_20432,N_20045);
nand U23972 (N_23972,N_22069,N_21192);
or U23973 (N_23973,N_20310,N_20545);
nand U23974 (N_23974,N_21863,N_20378);
xor U23975 (N_23975,N_22345,N_21789);
and U23976 (N_23976,N_20442,N_21938);
and U23977 (N_23977,N_21250,N_21676);
nand U23978 (N_23978,N_21667,N_20343);
xor U23979 (N_23979,N_22213,N_20007);
nor U23980 (N_23980,N_21817,N_20539);
xnor U23981 (N_23981,N_21753,N_20006);
nand U23982 (N_23982,N_20333,N_20073);
xor U23983 (N_23983,N_21064,N_21399);
xnor U23984 (N_23984,N_20395,N_21108);
and U23985 (N_23985,N_20297,N_20521);
or U23986 (N_23986,N_20333,N_21158);
or U23987 (N_23987,N_20370,N_20169);
nor U23988 (N_23988,N_21567,N_22035);
xor U23989 (N_23989,N_22289,N_21668);
nand U23990 (N_23990,N_21965,N_20189);
and U23991 (N_23991,N_20989,N_22135);
nand U23992 (N_23992,N_21401,N_20066);
nor U23993 (N_23993,N_21511,N_21784);
xnor U23994 (N_23994,N_20592,N_20938);
xor U23995 (N_23995,N_21629,N_21924);
nand U23996 (N_23996,N_22162,N_20686);
and U23997 (N_23997,N_20677,N_20282);
nand U23998 (N_23998,N_22145,N_21024);
or U23999 (N_23999,N_21488,N_21597);
and U24000 (N_24000,N_20731,N_20313);
and U24001 (N_24001,N_21092,N_22242);
and U24002 (N_24002,N_21480,N_20365);
nand U24003 (N_24003,N_20460,N_20372);
or U24004 (N_24004,N_21721,N_22463);
nor U24005 (N_24005,N_22111,N_21778);
xnor U24006 (N_24006,N_20440,N_22396);
and U24007 (N_24007,N_22068,N_21600);
xor U24008 (N_24008,N_22039,N_22021);
nand U24009 (N_24009,N_22483,N_20541);
nand U24010 (N_24010,N_20475,N_20946);
or U24011 (N_24011,N_20733,N_20256);
nor U24012 (N_24012,N_21268,N_20728);
and U24013 (N_24013,N_20612,N_22361);
or U24014 (N_24014,N_22061,N_21659);
xnor U24015 (N_24015,N_22295,N_20050);
nor U24016 (N_24016,N_22295,N_22487);
xnor U24017 (N_24017,N_21281,N_20147);
and U24018 (N_24018,N_20948,N_21059);
and U24019 (N_24019,N_21311,N_22089);
or U24020 (N_24020,N_21768,N_20986);
or U24021 (N_24021,N_22342,N_20833);
nand U24022 (N_24022,N_20434,N_20536);
xnor U24023 (N_24023,N_22408,N_22092);
or U24024 (N_24024,N_21444,N_21729);
nor U24025 (N_24025,N_20089,N_21350);
or U24026 (N_24026,N_22201,N_21341);
nand U24027 (N_24027,N_20692,N_20697);
nor U24028 (N_24028,N_21129,N_20523);
nand U24029 (N_24029,N_20443,N_21233);
and U24030 (N_24030,N_20152,N_20990);
nor U24031 (N_24031,N_22360,N_21942);
or U24032 (N_24032,N_21691,N_21496);
nand U24033 (N_24033,N_20108,N_20003);
or U24034 (N_24034,N_21010,N_20086);
nand U24035 (N_24035,N_20008,N_22002);
nor U24036 (N_24036,N_20937,N_21590);
nand U24037 (N_24037,N_22094,N_21819);
nor U24038 (N_24038,N_22264,N_22414);
nand U24039 (N_24039,N_20983,N_22370);
xor U24040 (N_24040,N_21609,N_20823);
nand U24041 (N_24041,N_22316,N_22027);
nand U24042 (N_24042,N_20547,N_21136);
nor U24043 (N_24043,N_22459,N_20615);
or U24044 (N_24044,N_22348,N_21956);
nand U24045 (N_24045,N_20736,N_20603);
xnor U24046 (N_24046,N_22094,N_20870);
nor U24047 (N_24047,N_21123,N_20271);
nor U24048 (N_24048,N_22479,N_21721);
and U24049 (N_24049,N_22478,N_20959);
nand U24050 (N_24050,N_21779,N_20100);
nor U24051 (N_24051,N_20313,N_20089);
nor U24052 (N_24052,N_20757,N_20004);
nor U24053 (N_24053,N_22384,N_20876);
and U24054 (N_24054,N_22166,N_20023);
and U24055 (N_24055,N_22226,N_20982);
nand U24056 (N_24056,N_22334,N_22415);
or U24057 (N_24057,N_21605,N_20068);
and U24058 (N_24058,N_20891,N_20507);
xor U24059 (N_24059,N_20507,N_22218);
nand U24060 (N_24060,N_22211,N_20103);
and U24061 (N_24061,N_22192,N_20622);
nand U24062 (N_24062,N_20744,N_21332);
nor U24063 (N_24063,N_21492,N_20119);
or U24064 (N_24064,N_20450,N_22142);
nor U24065 (N_24065,N_20213,N_20450);
nand U24066 (N_24066,N_21518,N_20218);
nor U24067 (N_24067,N_21230,N_22325);
nand U24068 (N_24068,N_20489,N_22112);
or U24069 (N_24069,N_20534,N_21668);
and U24070 (N_24070,N_21653,N_21851);
xor U24071 (N_24071,N_20830,N_20648);
and U24072 (N_24072,N_22071,N_21926);
and U24073 (N_24073,N_21554,N_20989);
or U24074 (N_24074,N_20444,N_20171);
and U24075 (N_24075,N_22238,N_22454);
nand U24076 (N_24076,N_22114,N_20638);
nor U24077 (N_24077,N_20005,N_21152);
nand U24078 (N_24078,N_20203,N_20810);
or U24079 (N_24079,N_20188,N_22401);
nand U24080 (N_24080,N_22324,N_21654);
nor U24081 (N_24081,N_21929,N_21503);
xor U24082 (N_24082,N_20529,N_21538);
or U24083 (N_24083,N_22237,N_21163);
or U24084 (N_24084,N_22139,N_21643);
or U24085 (N_24085,N_20722,N_20810);
nand U24086 (N_24086,N_21531,N_20593);
nand U24087 (N_24087,N_21796,N_21939);
xnor U24088 (N_24088,N_20476,N_22384);
nor U24089 (N_24089,N_20472,N_22301);
or U24090 (N_24090,N_20586,N_20765);
nor U24091 (N_24091,N_21611,N_22372);
and U24092 (N_24092,N_20981,N_20733);
xnor U24093 (N_24093,N_20763,N_20394);
or U24094 (N_24094,N_21717,N_22193);
or U24095 (N_24095,N_20740,N_21702);
nand U24096 (N_24096,N_21169,N_22283);
nor U24097 (N_24097,N_21974,N_20994);
or U24098 (N_24098,N_22272,N_21057);
nor U24099 (N_24099,N_20762,N_21152);
nand U24100 (N_24100,N_21795,N_20854);
and U24101 (N_24101,N_22070,N_20366);
nor U24102 (N_24102,N_20953,N_20129);
xnor U24103 (N_24103,N_20194,N_21380);
nor U24104 (N_24104,N_20000,N_21729);
xor U24105 (N_24105,N_20203,N_21695);
nor U24106 (N_24106,N_21949,N_21103);
nor U24107 (N_24107,N_21034,N_22121);
or U24108 (N_24108,N_20436,N_20040);
nor U24109 (N_24109,N_21288,N_22154);
or U24110 (N_24110,N_20613,N_22117);
or U24111 (N_24111,N_20669,N_21377);
nor U24112 (N_24112,N_22232,N_21878);
nor U24113 (N_24113,N_20796,N_20954);
xor U24114 (N_24114,N_21577,N_20513);
and U24115 (N_24115,N_21760,N_21423);
or U24116 (N_24116,N_22251,N_20189);
or U24117 (N_24117,N_20891,N_21027);
nand U24118 (N_24118,N_21410,N_20110);
or U24119 (N_24119,N_20174,N_21027);
nor U24120 (N_24120,N_21094,N_21407);
or U24121 (N_24121,N_20963,N_20090);
and U24122 (N_24122,N_21830,N_21302);
xnor U24123 (N_24123,N_21257,N_22295);
nand U24124 (N_24124,N_21592,N_21823);
nor U24125 (N_24125,N_20385,N_22136);
nand U24126 (N_24126,N_20950,N_21623);
xnor U24127 (N_24127,N_20020,N_20957);
and U24128 (N_24128,N_21284,N_21523);
or U24129 (N_24129,N_20508,N_20297);
or U24130 (N_24130,N_22474,N_20045);
xnor U24131 (N_24131,N_21353,N_21172);
and U24132 (N_24132,N_21909,N_20768);
nor U24133 (N_24133,N_20299,N_21202);
and U24134 (N_24134,N_22415,N_20556);
or U24135 (N_24135,N_21014,N_21510);
and U24136 (N_24136,N_21735,N_20421);
or U24137 (N_24137,N_20853,N_21187);
or U24138 (N_24138,N_22429,N_21532);
nor U24139 (N_24139,N_20218,N_20382);
xnor U24140 (N_24140,N_20956,N_21553);
or U24141 (N_24141,N_21613,N_22493);
nand U24142 (N_24142,N_20531,N_20270);
or U24143 (N_24143,N_20438,N_21289);
and U24144 (N_24144,N_20398,N_21187);
xor U24145 (N_24145,N_21298,N_21792);
or U24146 (N_24146,N_21059,N_20187);
xor U24147 (N_24147,N_20397,N_21519);
nand U24148 (N_24148,N_21593,N_20957);
nand U24149 (N_24149,N_20899,N_21706);
nand U24150 (N_24150,N_22060,N_21264);
or U24151 (N_24151,N_22372,N_20430);
xnor U24152 (N_24152,N_22496,N_20197);
nand U24153 (N_24153,N_20178,N_21231);
nor U24154 (N_24154,N_22426,N_20609);
or U24155 (N_24155,N_22029,N_21424);
and U24156 (N_24156,N_22364,N_21142);
nand U24157 (N_24157,N_20743,N_22405);
and U24158 (N_24158,N_22309,N_20937);
xnor U24159 (N_24159,N_22079,N_20737);
xor U24160 (N_24160,N_20513,N_20355);
nor U24161 (N_24161,N_22377,N_21511);
nand U24162 (N_24162,N_20304,N_21234);
xnor U24163 (N_24163,N_20146,N_21989);
xor U24164 (N_24164,N_22492,N_22102);
and U24165 (N_24165,N_21519,N_21794);
or U24166 (N_24166,N_21741,N_21632);
nor U24167 (N_24167,N_21295,N_21888);
or U24168 (N_24168,N_21135,N_20698);
nand U24169 (N_24169,N_20354,N_21466);
and U24170 (N_24170,N_22109,N_20654);
nand U24171 (N_24171,N_21787,N_20614);
and U24172 (N_24172,N_21597,N_21700);
nand U24173 (N_24173,N_22104,N_22410);
nor U24174 (N_24174,N_21132,N_21417);
nand U24175 (N_24175,N_20552,N_22055);
and U24176 (N_24176,N_21801,N_22041);
and U24177 (N_24177,N_22187,N_20469);
xor U24178 (N_24178,N_21223,N_20407);
or U24179 (N_24179,N_21688,N_21510);
nor U24180 (N_24180,N_20930,N_21977);
nor U24181 (N_24181,N_22380,N_21896);
nand U24182 (N_24182,N_21282,N_21366);
xnor U24183 (N_24183,N_21668,N_21161);
or U24184 (N_24184,N_20432,N_21307);
and U24185 (N_24185,N_21792,N_20341);
xor U24186 (N_24186,N_22167,N_20903);
nand U24187 (N_24187,N_21384,N_20983);
nand U24188 (N_24188,N_20721,N_20182);
or U24189 (N_24189,N_21813,N_22420);
nor U24190 (N_24190,N_20144,N_21412);
or U24191 (N_24191,N_21760,N_21525);
and U24192 (N_24192,N_21707,N_21652);
nand U24193 (N_24193,N_20334,N_21398);
xnor U24194 (N_24194,N_20925,N_22093);
xnor U24195 (N_24195,N_22382,N_20192);
and U24196 (N_24196,N_22269,N_20868);
nor U24197 (N_24197,N_21814,N_20417);
or U24198 (N_24198,N_22120,N_20861);
and U24199 (N_24199,N_21695,N_21388);
xnor U24200 (N_24200,N_20196,N_21980);
nor U24201 (N_24201,N_22242,N_20261);
xnor U24202 (N_24202,N_21499,N_21526);
nand U24203 (N_24203,N_20410,N_21712);
xnor U24204 (N_24204,N_21613,N_21885);
nor U24205 (N_24205,N_22284,N_21721);
and U24206 (N_24206,N_21579,N_20535);
nand U24207 (N_24207,N_21313,N_21996);
or U24208 (N_24208,N_20014,N_20119);
nand U24209 (N_24209,N_21274,N_22421);
nand U24210 (N_24210,N_22031,N_20379);
nor U24211 (N_24211,N_21891,N_22180);
nor U24212 (N_24212,N_21929,N_21756);
and U24213 (N_24213,N_21223,N_21340);
or U24214 (N_24214,N_22204,N_20549);
nand U24215 (N_24215,N_21275,N_21634);
xnor U24216 (N_24216,N_20179,N_22313);
or U24217 (N_24217,N_20889,N_22210);
and U24218 (N_24218,N_20743,N_21989);
nor U24219 (N_24219,N_20068,N_20171);
nor U24220 (N_24220,N_20198,N_21421);
nor U24221 (N_24221,N_22019,N_21731);
or U24222 (N_24222,N_21291,N_20470);
and U24223 (N_24223,N_21704,N_20113);
xor U24224 (N_24224,N_21049,N_20811);
or U24225 (N_24225,N_21576,N_20940);
nand U24226 (N_24226,N_20191,N_20765);
or U24227 (N_24227,N_21205,N_20358);
or U24228 (N_24228,N_20270,N_20789);
nor U24229 (N_24229,N_22330,N_20805);
nand U24230 (N_24230,N_21680,N_20834);
nand U24231 (N_24231,N_20136,N_22442);
xor U24232 (N_24232,N_21416,N_21746);
nand U24233 (N_24233,N_20265,N_21517);
xnor U24234 (N_24234,N_22077,N_21075);
xnor U24235 (N_24235,N_20397,N_22072);
nand U24236 (N_24236,N_20869,N_20714);
nand U24237 (N_24237,N_21980,N_21999);
xor U24238 (N_24238,N_20210,N_21242);
or U24239 (N_24239,N_21930,N_20833);
nand U24240 (N_24240,N_20444,N_20582);
nand U24241 (N_24241,N_21443,N_21985);
and U24242 (N_24242,N_21638,N_22047);
nor U24243 (N_24243,N_21934,N_22437);
nand U24244 (N_24244,N_21862,N_20899);
nor U24245 (N_24245,N_21543,N_20485);
or U24246 (N_24246,N_20105,N_20840);
and U24247 (N_24247,N_21948,N_21941);
and U24248 (N_24248,N_22416,N_21716);
xnor U24249 (N_24249,N_21001,N_21907);
or U24250 (N_24250,N_21977,N_21882);
xor U24251 (N_24251,N_21809,N_22328);
nand U24252 (N_24252,N_21135,N_22120);
and U24253 (N_24253,N_21275,N_21344);
nand U24254 (N_24254,N_22442,N_21136);
nand U24255 (N_24255,N_20803,N_21381);
or U24256 (N_24256,N_21541,N_22272);
or U24257 (N_24257,N_21243,N_20704);
xnor U24258 (N_24258,N_20294,N_20592);
or U24259 (N_24259,N_22455,N_22430);
or U24260 (N_24260,N_20886,N_22232);
and U24261 (N_24261,N_21499,N_21518);
or U24262 (N_24262,N_20093,N_21006);
xor U24263 (N_24263,N_20882,N_20984);
nand U24264 (N_24264,N_20720,N_22116);
or U24265 (N_24265,N_21049,N_22374);
and U24266 (N_24266,N_20903,N_21493);
nor U24267 (N_24267,N_21148,N_21364);
nand U24268 (N_24268,N_20391,N_20641);
and U24269 (N_24269,N_21796,N_21531);
xnor U24270 (N_24270,N_21570,N_20055);
and U24271 (N_24271,N_22218,N_20496);
nor U24272 (N_24272,N_21388,N_20133);
xnor U24273 (N_24273,N_20297,N_20540);
and U24274 (N_24274,N_21037,N_22136);
nand U24275 (N_24275,N_20314,N_21555);
nor U24276 (N_24276,N_22064,N_22229);
xnor U24277 (N_24277,N_21746,N_22156);
nor U24278 (N_24278,N_22116,N_20691);
nand U24279 (N_24279,N_21589,N_21104);
nor U24280 (N_24280,N_22223,N_20883);
xor U24281 (N_24281,N_21140,N_20975);
nor U24282 (N_24282,N_21965,N_20240);
or U24283 (N_24283,N_21877,N_21753);
or U24284 (N_24284,N_20516,N_22263);
or U24285 (N_24285,N_21521,N_21256);
or U24286 (N_24286,N_20532,N_22497);
or U24287 (N_24287,N_22361,N_22041);
nor U24288 (N_24288,N_20575,N_21632);
nor U24289 (N_24289,N_21543,N_21788);
and U24290 (N_24290,N_21348,N_20350);
and U24291 (N_24291,N_21749,N_20854);
and U24292 (N_24292,N_21317,N_22078);
or U24293 (N_24293,N_20548,N_20278);
nand U24294 (N_24294,N_21733,N_22323);
or U24295 (N_24295,N_20330,N_20021);
and U24296 (N_24296,N_21224,N_21537);
xor U24297 (N_24297,N_20999,N_22254);
or U24298 (N_24298,N_21967,N_21047);
and U24299 (N_24299,N_21284,N_21150);
and U24300 (N_24300,N_21517,N_21277);
and U24301 (N_24301,N_21463,N_20768);
nand U24302 (N_24302,N_21788,N_22167);
and U24303 (N_24303,N_21920,N_21532);
and U24304 (N_24304,N_20736,N_22335);
or U24305 (N_24305,N_20589,N_21276);
and U24306 (N_24306,N_22172,N_20103);
xnor U24307 (N_24307,N_22200,N_21710);
nand U24308 (N_24308,N_21815,N_20503);
or U24309 (N_24309,N_22124,N_20627);
nor U24310 (N_24310,N_21529,N_20945);
nand U24311 (N_24311,N_22283,N_20428);
xnor U24312 (N_24312,N_22437,N_20428);
or U24313 (N_24313,N_20154,N_22205);
nor U24314 (N_24314,N_20474,N_20331);
nand U24315 (N_24315,N_20290,N_21231);
xnor U24316 (N_24316,N_22277,N_20697);
or U24317 (N_24317,N_20436,N_22239);
or U24318 (N_24318,N_20304,N_22380);
nand U24319 (N_24319,N_21569,N_20767);
nor U24320 (N_24320,N_21378,N_21187);
or U24321 (N_24321,N_20881,N_21743);
xor U24322 (N_24322,N_21365,N_20421);
or U24323 (N_24323,N_20931,N_21882);
nand U24324 (N_24324,N_21434,N_22408);
xor U24325 (N_24325,N_20989,N_21605);
or U24326 (N_24326,N_21334,N_21398);
and U24327 (N_24327,N_21958,N_20546);
nor U24328 (N_24328,N_22438,N_22113);
or U24329 (N_24329,N_21272,N_21758);
or U24330 (N_24330,N_21214,N_21889);
and U24331 (N_24331,N_20206,N_20534);
and U24332 (N_24332,N_21821,N_20121);
or U24333 (N_24333,N_21048,N_21399);
xor U24334 (N_24334,N_21276,N_21849);
nor U24335 (N_24335,N_21000,N_21771);
nand U24336 (N_24336,N_22461,N_22289);
nor U24337 (N_24337,N_22436,N_22100);
or U24338 (N_24338,N_21401,N_21411);
nand U24339 (N_24339,N_20217,N_21182);
or U24340 (N_24340,N_20884,N_21049);
and U24341 (N_24341,N_21638,N_21423);
or U24342 (N_24342,N_20840,N_20419);
and U24343 (N_24343,N_20183,N_22339);
and U24344 (N_24344,N_21903,N_20176);
xor U24345 (N_24345,N_20991,N_22148);
xnor U24346 (N_24346,N_20663,N_20573);
or U24347 (N_24347,N_21770,N_21191);
and U24348 (N_24348,N_21878,N_22398);
and U24349 (N_24349,N_22021,N_21104);
nand U24350 (N_24350,N_21053,N_21390);
nor U24351 (N_24351,N_22119,N_21522);
xor U24352 (N_24352,N_20039,N_20670);
xor U24353 (N_24353,N_20379,N_20143);
nand U24354 (N_24354,N_20318,N_20892);
and U24355 (N_24355,N_20758,N_20994);
or U24356 (N_24356,N_20079,N_21616);
nand U24357 (N_24357,N_20537,N_20600);
nor U24358 (N_24358,N_22414,N_20996);
and U24359 (N_24359,N_21568,N_22238);
nand U24360 (N_24360,N_20207,N_21314);
nor U24361 (N_24361,N_21643,N_21135);
nor U24362 (N_24362,N_21352,N_21893);
nor U24363 (N_24363,N_22364,N_22267);
nor U24364 (N_24364,N_21267,N_20380);
xor U24365 (N_24365,N_22045,N_22413);
nor U24366 (N_24366,N_21292,N_20428);
and U24367 (N_24367,N_21858,N_22146);
or U24368 (N_24368,N_21527,N_21131);
xor U24369 (N_24369,N_21287,N_20522);
or U24370 (N_24370,N_21921,N_21581);
nor U24371 (N_24371,N_21597,N_20404);
and U24372 (N_24372,N_20828,N_21311);
xnor U24373 (N_24373,N_20650,N_22224);
or U24374 (N_24374,N_21668,N_22271);
and U24375 (N_24375,N_21384,N_21138);
and U24376 (N_24376,N_21629,N_21770);
nor U24377 (N_24377,N_21936,N_21216);
xnor U24378 (N_24378,N_20454,N_21321);
nor U24379 (N_24379,N_22172,N_21377);
nand U24380 (N_24380,N_20138,N_21213);
xor U24381 (N_24381,N_21528,N_22358);
nor U24382 (N_24382,N_21008,N_21516);
xnor U24383 (N_24383,N_20953,N_20761);
nand U24384 (N_24384,N_22242,N_20859);
or U24385 (N_24385,N_20673,N_22184);
xnor U24386 (N_24386,N_20361,N_21527);
xor U24387 (N_24387,N_22475,N_21505);
nor U24388 (N_24388,N_20612,N_20108);
and U24389 (N_24389,N_21228,N_20969);
or U24390 (N_24390,N_22401,N_22313);
or U24391 (N_24391,N_21540,N_22394);
nor U24392 (N_24392,N_22298,N_21215);
and U24393 (N_24393,N_20646,N_21541);
or U24394 (N_24394,N_22029,N_22475);
nor U24395 (N_24395,N_20947,N_20143);
xnor U24396 (N_24396,N_21301,N_20136);
and U24397 (N_24397,N_20300,N_20396);
or U24398 (N_24398,N_22033,N_20383);
nor U24399 (N_24399,N_20984,N_20488);
or U24400 (N_24400,N_21581,N_21028);
or U24401 (N_24401,N_20131,N_20693);
nor U24402 (N_24402,N_22222,N_22240);
xor U24403 (N_24403,N_21172,N_22243);
or U24404 (N_24404,N_20876,N_22404);
xor U24405 (N_24405,N_21265,N_21453);
nand U24406 (N_24406,N_21659,N_20714);
xor U24407 (N_24407,N_20222,N_20381);
or U24408 (N_24408,N_22454,N_21766);
and U24409 (N_24409,N_22205,N_20298);
nor U24410 (N_24410,N_21640,N_20914);
or U24411 (N_24411,N_20086,N_21535);
or U24412 (N_24412,N_20588,N_20785);
or U24413 (N_24413,N_20112,N_21195);
nor U24414 (N_24414,N_20703,N_21450);
or U24415 (N_24415,N_20792,N_21161);
and U24416 (N_24416,N_21458,N_20563);
or U24417 (N_24417,N_21503,N_20018);
or U24418 (N_24418,N_21443,N_21722);
or U24419 (N_24419,N_21628,N_21415);
or U24420 (N_24420,N_20140,N_22294);
or U24421 (N_24421,N_20315,N_21899);
nand U24422 (N_24422,N_20283,N_22083);
nand U24423 (N_24423,N_20470,N_21257);
nor U24424 (N_24424,N_22487,N_22384);
xor U24425 (N_24425,N_21869,N_20221);
and U24426 (N_24426,N_22195,N_21725);
xor U24427 (N_24427,N_20338,N_21204);
xor U24428 (N_24428,N_21067,N_21057);
xnor U24429 (N_24429,N_20809,N_21554);
nor U24430 (N_24430,N_20430,N_22231);
and U24431 (N_24431,N_20183,N_20991);
or U24432 (N_24432,N_20151,N_21697);
nand U24433 (N_24433,N_22317,N_22380);
or U24434 (N_24434,N_20003,N_22294);
xnor U24435 (N_24435,N_20372,N_21395);
nor U24436 (N_24436,N_21806,N_21644);
xor U24437 (N_24437,N_20827,N_20553);
or U24438 (N_24438,N_20339,N_21647);
nand U24439 (N_24439,N_20390,N_21663);
nand U24440 (N_24440,N_21963,N_20079);
or U24441 (N_24441,N_20422,N_21024);
xnor U24442 (N_24442,N_20221,N_20059);
nor U24443 (N_24443,N_20692,N_21347);
xnor U24444 (N_24444,N_22014,N_22398);
xnor U24445 (N_24445,N_20784,N_21382);
xor U24446 (N_24446,N_20901,N_20431);
or U24447 (N_24447,N_22496,N_21347);
nand U24448 (N_24448,N_22205,N_20226);
xnor U24449 (N_24449,N_22220,N_21665);
or U24450 (N_24450,N_21819,N_21633);
and U24451 (N_24451,N_21356,N_21531);
nand U24452 (N_24452,N_21674,N_21270);
xor U24453 (N_24453,N_20983,N_21836);
nor U24454 (N_24454,N_20882,N_21433);
nand U24455 (N_24455,N_22094,N_20803);
and U24456 (N_24456,N_21413,N_22287);
and U24457 (N_24457,N_20437,N_21010);
nand U24458 (N_24458,N_21061,N_20902);
xor U24459 (N_24459,N_21199,N_22403);
nor U24460 (N_24460,N_20840,N_20431);
nand U24461 (N_24461,N_22434,N_21045);
or U24462 (N_24462,N_21035,N_21176);
or U24463 (N_24463,N_21552,N_20217);
nand U24464 (N_24464,N_21101,N_21172);
or U24465 (N_24465,N_22497,N_20398);
nand U24466 (N_24466,N_22149,N_21891);
nor U24467 (N_24467,N_20435,N_21356);
or U24468 (N_24468,N_20452,N_20987);
xor U24469 (N_24469,N_20719,N_21525);
nand U24470 (N_24470,N_20475,N_20358);
nor U24471 (N_24471,N_21952,N_20273);
nand U24472 (N_24472,N_21928,N_21859);
nor U24473 (N_24473,N_21340,N_21654);
nand U24474 (N_24474,N_21371,N_20594);
nand U24475 (N_24475,N_20776,N_22439);
xnor U24476 (N_24476,N_21744,N_21040);
or U24477 (N_24477,N_20963,N_21107);
nor U24478 (N_24478,N_21402,N_22074);
xor U24479 (N_24479,N_20304,N_21054);
xor U24480 (N_24480,N_20351,N_22082);
or U24481 (N_24481,N_22442,N_20035);
nand U24482 (N_24482,N_20349,N_22060);
nor U24483 (N_24483,N_20360,N_20247);
and U24484 (N_24484,N_20718,N_20255);
xor U24485 (N_24485,N_21504,N_21073);
xor U24486 (N_24486,N_20268,N_20102);
nand U24487 (N_24487,N_22345,N_21159);
xnor U24488 (N_24488,N_20902,N_22337);
nand U24489 (N_24489,N_21860,N_21281);
nor U24490 (N_24490,N_21458,N_21732);
or U24491 (N_24491,N_20629,N_20136);
and U24492 (N_24492,N_22397,N_21666);
and U24493 (N_24493,N_21061,N_21368);
or U24494 (N_24494,N_21650,N_21519);
nand U24495 (N_24495,N_21903,N_21344);
and U24496 (N_24496,N_21962,N_20893);
xnor U24497 (N_24497,N_20107,N_20538);
xnor U24498 (N_24498,N_20604,N_20544);
and U24499 (N_24499,N_21656,N_21681);
xor U24500 (N_24500,N_20588,N_22319);
xnor U24501 (N_24501,N_20977,N_20180);
nor U24502 (N_24502,N_21738,N_21645);
xor U24503 (N_24503,N_21056,N_20901);
or U24504 (N_24504,N_22383,N_21163);
nand U24505 (N_24505,N_21125,N_20009);
or U24506 (N_24506,N_20681,N_20403);
nand U24507 (N_24507,N_21562,N_21340);
nand U24508 (N_24508,N_22467,N_21383);
and U24509 (N_24509,N_20920,N_21086);
xnor U24510 (N_24510,N_21640,N_22151);
nand U24511 (N_24511,N_21677,N_21028);
xor U24512 (N_24512,N_22330,N_21103);
nand U24513 (N_24513,N_21230,N_21634);
or U24514 (N_24514,N_22179,N_21045);
nor U24515 (N_24515,N_22355,N_20378);
nor U24516 (N_24516,N_21411,N_21521);
or U24517 (N_24517,N_21904,N_20238);
or U24518 (N_24518,N_22341,N_22404);
nor U24519 (N_24519,N_20185,N_20302);
nand U24520 (N_24520,N_20196,N_21871);
nor U24521 (N_24521,N_21427,N_20622);
nand U24522 (N_24522,N_21730,N_20183);
or U24523 (N_24523,N_21914,N_20200);
and U24524 (N_24524,N_20687,N_21715);
or U24525 (N_24525,N_20440,N_21565);
xnor U24526 (N_24526,N_22222,N_22414);
or U24527 (N_24527,N_22094,N_21070);
and U24528 (N_24528,N_22304,N_20791);
nand U24529 (N_24529,N_21294,N_20308);
nor U24530 (N_24530,N_21461,N_22143);
nor U24531 (N_24531,N_21601,N_22322);
or U24532 (N_24532,N_20524,N_22204);
and U24533 (N_24533,N_20286,N_21283);
nand U24534 (N_24534,N_22206,N_20743);
and U24535 (N_24535,N_21096,N_20616);
or U24536 (N_24536,N_22389,N_21395);
nor U24537 (N_24537,N_20513,N_21108);
or U24538 (N_24538,N_20021,N_20137);
nor U24539 (N_24539,N_22439,N_22469);
and U24540 (N_24540,N_20878,N_20443);
or U24541 (N_24541,N_22303,N_22454);
or U24542 (N_24542,N_21264,N_20963);
xnor U24543 (N_24543,N_21933,N_21005);
nand U24544 (N_24544,N_21279,N_22140);
nand U24545 (N_24545,N_21034,N_21721);
nor U24546 (N_24546,N_20297,N_20616);
or U24547 (N_24547,N_21133,N_20691);
nor U24548 (N_24548,N_21195,N_21739);
nor U24549 (N_24549,N_21830,N_21975);
or U24550 (N_24550,N_22440,N_21256);
or U24551 (N_24551,N_21260,N_20812);
or U24552 (N_24552,N_20890,N_22091);
and U24553 (N_24553,N_21960,N_20104);
nand U24554 (N_24554,N_21124,N_21257);
xor U24555 (N_24555,N_20516,N_22034);
xnor U24556 (N_24556,N_20079,N_21734);
or U24557 (N_24557,N_21817,N_21439);
xor U24558 (N_24558,N_21526,N_21544);
xor U24559 (N_24559,N_21359,N_20123);
nand U24560 (N_24560,N_21714,N_21589);
or U24561 (N_24561,N_21297,N_21804);
nand U24562 (N_24562,N_20534,N_20576);
nor U24563 (N_24563,N_21320,N_22152);
nor U24564 (N_24564,N_21752,N_20257);
nor U24565 (N_24565,N_22273,N_20501);
nor U24566 (N_24566,N_21310,N_21931);
and U24567 (N_24567,N_21796,N_21670);
xor U24568 (N_24568,N_21919,N_21476);
and U24569 (N_24569,N_21974,N_21978);
and U24570 (N_24570,N_22317,N_21734);
and U24571 (N_24571,N_20880,N_21479);
xor U24572 (N_24572,N_21190,N_21479);
and U24573 (N_24573,N_20644,N_22157);
nand U24574 (N_24574,N_21573,N_20431);
xnor U24575 (N_24575,N_22134,N_21559);
nand U24576 (N_24576,N_21590,N_20952);
nand U24577 (N_24577,N_21981,N_20078);
and U24578 (N_24578,N_21444,N_22278);
xnor U24579 (N_24579,N_20481,N_21321);
xor U24580 (N_24580,N_21873,N_21697);
and U24581 (N_24581,N_22272,N_21293);
or U24582 (N_24582,N_21678,N_22324);
xor U24583 (N_24583,N_20145,N_22404);
nand U24584 (N_24584,N_21969,N_22436);
and U24585 (N_24585,N_22296,N_20432);
or U24586 (N_24586,N_21882,N_21857);
or U24587 (N_24587,N_22260,N_21547);
or U24588 (N_24588,N_22013,N_21442);
and U24589 (N_24589,N_22458,N_20877);
nor U24590 (N_24590,N_21947,N_20630);
and U24591 (N_24591,N_21890,N_22258);
nand U24592 (N_24592,N_21075,N_22057);
or U24593 (N_24593,N_22293,N_21143);
xnor U24594 (N_24594,N_20113,N_22466);
nand U24595 (N_24595,N_22434,N_21530);
or U24596 (N_24596,N_22159,N_20058);
and U24597 (N_24597,N_22336,N_20905);
nor U24598 (N_24598,N_20873,N_20746);
xnor U24599 (N_24599,N_20505,N_20388);
or U24600 (N_24600,N_20462,N_22071);
xor U24601 (N_24601,N_22151,N_20249);
or U24602 (N_24602,N_20706,N_21315);
nor U24603 (N_24603,N_21091,N_22124);
and U24604 (N_24604,N_20590,N_21405);
and U24605 (N_24605,N_20680,N_20493);
or U24606 (N_24606,N_20720,N_20379);
xnor U24607 (N_24607,N_20164,N_20717);
nor U24608 (N_24608,N_21577,N_20049);
xnor U24609 (N_24609,N_21404,N_21127);
and U24610 (N_24610,N_21014,N_21101);
xor U24611 (N_24611,N_21898,N_21797);
or U24612 (N_24612,N_21311,N_20820);
and U24613 (N_24613,N_20821,N_20102);
xnor U24614 (N_24614,N_20143,N_20670);
xor U24615 (N_24615,N_22009,N_21717);
nor U24616 (N_24616,N_22031,N_20315);
or U24617 (N_24617,N_20559,N_21297);
nor U24618 (N_24618,N_20213,N_21755);
nand U24619 (N_24619,N_21794,N_21086);
or U24620 (N_24620,N_21880,N_20147);
xnor U24621 (N_24621,N_20462,N_22052);
xor U24622 (N_24622,N_20688,N_21804);
nand U24623 (N_24623,N_21842,N_20385);
or U24624 (N_24624,N_20906,N_21519);
nand U24625 (N_24625,N_21783,N_20651);
nor U24626 (N_24626,N_20627,N_22159);
or U24627 (N_24627,N_21798,N_21174);
nand U24628 (N_24628,N_20918,N_20273);
nand U24629 (N_24629,N_21380,N_21840);
nor U24630 (N_24630,N_22160,N_20815);
nor U24631 (N_24631,N_22211,N_21589);
nor U24632 (N_24632,N_21352,N_22002);
nor U24633 (N_24633,N_22322,N_20763);
or U24634 (N_24634,N_21145,N_20261);
nand U24635 (N_24635,N_22392,N_20693);
and U24636 (N_24636,N_20293,N_20529);
xnor U24637 (N_24637,N_21078,N_21924);
and U24638 (N_24638,N_22040,N_21460);
or U24639 (N_24639,N_21479,N_21578);
xor U24640 (N_24640,N_22164,N_20131);
nand U24641 (N_24641,N_21526,N_22301);
or U24642 (N_24642,N_20140,N_20573);
nor U24643 (N_24643,N_21957,N_21231);
or U24644 (N_24644,N_21895,N_21509);
or U24645 (N_24645,N_20269,N_21927);
nor U24646 (N_24646,N_21798,N_22251);
nor U24647 (N_24647,N_22156,N_20201);
xor U24648 (N_24648,N_21713,N_20218);
or U24649 (N_24649,N_20316,N_22233);
and U24650 (N_24650,N_22125,N_21983);
nor U24651 (N_24651,N_22318,N_21358);
xnor U24652 (N_24652,N_20969,N_20641);
or U24653 (N_24653,N_21336,N_22335);
and U24654 (N_24654,N_21899,N_21533);
xnor U24655 (N_24655,N_22412,N_20868);
xor U24656 (N_24656,N_22048,N_20387);
nor U24657 (N_24657,N_21093,N_21014);
and U24658 (N_24658,N_22026,N_21844);
nand U24659 (N_24659,N_22339,N_20253);
nand U24660 (N_24660,N_20376,N_21256);
xnor U24661 (N_24661,N_21958,N_22364);
or U24662 (N_24662,N_20772,N_21134);
or U24663 (N_24663,N_22170,N_21195);
or U24664 (N_24664,N_22432,N_21391);
or U24665 (N_24665,N_21356,N_21268);
or U24666 (N_24666,N_22033,N_20176);
or U24667 (N_24667,N_21519,N_21251);
or U24668 (N_24668,N_21883,N_21112);
nor U24669 (N_24669,N_21421,N_21135);
or U24670 (N_24670,N_20915,N_22419);
and U24671 (N_24671,N_21862,N_22436);
or U24672 (N_24672,N_20504,N_20958);
nor U24673 (N_24673,N_21641,N_22083);
or U24674 (N_24674,N_21467,N_20774);
nor U24675 (N_24675,N_21400,N_20471);
nand U24676 (N_24676,N_22445,N_22058);
and U24677 (N_24677,N_21725,N_20899);
or U24678 (N_24678,N_20362,N_20991);
and U24679 (N_24679,N_21208,N_22195);
nand U24680 (N_24680,N_20459,N_21608);
xnor U24681 (N_24681,N_22318,N_22408);
nor U24682 (N_24682,N_22043,N_20338);
and U24683 (N_24683,N_22476,N_21503);
or U24684 (N_24684,N_20155,N_20542);
nor U24685 (N_24685,N_21565,N_20728);
nand U24686 (N_24686,N_20061,N_21079);
nor U24687 (N_24687,N_20021,N_20796);
nor U24688 (N_24688,N_21300,N_20177);
nor U24689 (N_24689,N_20891,N_22207);
xor U24690 (N_24690,N_22180,N_21849);
nor U24691 (N_24691,N_22242,N_21161);
xnor U24692 (N_24692,N_21568,N_21282);
and U24693 (N_24693,N_20270,N_20294);
and U24694 (N_24694,N_22109,N_22259);
or U24695 (N_24695,N_20570,N_22384);
xor U24696 (N_24696,N_22364,N_22079);
xor U24697 (N_24697,N_20552,N_20893);
or U24698 (N_24698,N_21785,N_21337);
xor U24699 (N_24699,N_20860,N_20599);
and U24700 (N_24700,N_21485,N_22388);
xnor U24701 (N_24701,N_22127,N_20911);
xor U24702 (N_24702,N_22477,N_20934);
nor U24703 (N_24703,N_21586,N_21242);
or U24704 (N_24704,N_22355,N_22091);
or U24705 (N_24705,N_21045,N_20798);
nor U24706 (N_24706,N_20380,N_20349);
or U24707 (N_24707,N_20261,N_20504);
nor U24708 (N_24708,N_21566,N_22191);
nand U24709 (N_24709,N_22434,N_21875);
nor U24710 (N_24710,N_22287,N_21351);
nand U24711 (N_24711,N_22194,N_20981);
nor U24712 (N_24712,N_20875,N_21299);
nand U24713 (N_24713,N_20785,N_22339);
and U24714 (N_24714,N_20641,N_21873);
nand U24715 (N_24715,N_22284,N_21286);
nand U24716 (N_24716,N_20186,N_21432);
and U24717 (N_24717,N_22358,N_20898);
and U24718 (N_24718,N_20758,N_20813);
nand U24719 (N_24719,N_21853,N_20089);
or U24720 (N_24720,N_20581,N_22094);
nor U24721 (N_24721,N_20630,N_20013);
nor U24722 (N_24722,N_21120,N_22453);
nor U24723 (N_24723,N_20655,N_20538);
or U24724 (N_24724,N_22242,N_20689);
nor U24725 (N_24725,N_20571,N_20836);
xor U24726 (N_24726,N_20606,N_22026);
or U24727 (N_24727,N_21144,N_21863);
xor U24728 (N_24728,N_20890,N_20160);
nand U24729 (N_24729,N_22494,N_22004);
or U24730 (N_24730,N_20512,N_21294);
nand U24731 (N_24731,N_22179,N_21562);
nand U24732 (N_24732,N_20997,N_21212);
xor U24733 (N_24733,N_20230,N_21644);
and U24734 (N_24734,N_21573,N_21078);
nand U24735 (N_24735,N_20439,N_20414);
or U24736 (N_24736,N_20100,N_20086);
xnor U24737 (N_24737,N_22258,N_20339);
nand U24738 (N_24738,N_22392,N_20256);
or U24739 (N_24739,N_22495,N_20312);
and U24740 (N_24740,N_20639,N_22303);
or U24741 (N_24741,N_20407,N_20861);
nor U24742 (N_24742,N_20869,N_21503);
and U24743 (N_24743,N_22101,N_21901);
or U24744 (N_24744,N_21967,N_21257);
or U24745 (N_24745,N_21668,N_21727);
nor U24746 (N_24746,N_21053,N_20152);
and U24747 (N_24747,N_20219,N_21529);
nand U24748 (N_24748,N_21974,N_20889);
nand U24749 (N_24749,N_20271,N_22009);
or U24750 (N_24750,N_20480,N_21048);
nand U24751 (N_24751,N_21497,N_21340);
xor U24752 (N_24752,N_21946,N_21168);
nor U24753 (N_24753,N_22068,N_20188);
and U24754 (N_24754,N_20343,N_21493);
nand U24755 (N_24755,N_22044,N_21407);
nand U24756 (N_24756,N_22171,N_21235);
nand U24757 (N_24757,N_21397,N_20235);
and U24758 (N_24758,N_21952,N_20994);
and U24759 (N_24759,N_20211,N_20927);
nor U24760 (N_24760,N_22404,N_21406);
or U24761 (N_24761,N_20184,N_22214);
and U24762 (N_24762,N_21482,N_20669);
xnor U24763 (N_24763,N_21099,N_21918);
nand U24764 (N_24764,N_22095,N_22419);
nand U24765 (N_24765,N_21136,N_21962);
xnor U24766 (N_24766,N_21714,N_20583);
or U24767 (N_24767,N_20116,N_21445);
nor U24768 (N_24768,N_20427,N_20292);
nor U24769 (N_24769,N_21805,N_20137);
nand U24770 (N_24770,N_20159,N_21684);
or U24771 (N_24771,N_22435,N_22444);
nor U24772 (N_24772,N_20202,N_21137);
nand U24773 (N_24773,N_20386,N_20837);
nand U24774 (N_24774,N_21776,N_20167);
and U24775 (N_24775,N_21781,N_22261);
nand U24776 (N_24776,N_20521,N_22279);
xor U24777 (N_24777,N_21760,N_20494);
xor U24778 (N_24778,N_22350,N_20398);
or U24779 (N_24779,N_20873,N_21971);
xnor U24780 (N_24780,N_21875,N_20046);
or U24781 (N_24781,N_22102,N_21415);
nand U24782 (N_24782,N_21990,N_21797);
or U24783 (N_24783,N_22273,N_22256);
and U24784 (N_24784,N_20262,N_21011);
and U24785 (N_24785,N_21931,N_20795);
and U24786 (N_24786,N_20055,N_20312);
and U24787 (N_24787,N_20943,N_20719);
xnor U24788 (N_24788,N_21187,N_21037);
xnor U24789 (N_24789,N_20967,N_21755);
nor U24790 (N_24790,N_21647,N_21312);
xnor U24791 (N_24791,N_21187,N_21541);
or U24792 (N_24792,N_21264,N_20308);
or U24793 (N_24793,N_20143,N_22018);
xor U24794 (N_24794,N_22458,N_21875);
xnor U24795 (N_24795,N_20652,N_22276);
or U24796 (N_24796,N_21729,N_21897);
nor U24797 (N_24797,N_22388,N_20132);
nand U24798 (N_24798,N_20957,N_20983);
and U24799 (N_24799,N_21836,N_21215);
or U24800 (N_24800,N_21763,N_20900);
and U24801 (N_24801,N_20062,N_21753);
nand U24802 (N_24802,N_21942,N_21908);
nand U24803 (N_24803,N_22137,N_20309);
and U24804 (N_24804,N_20196,N_20798);
and U24805 (N_24805,N_20798,N_22465);
nor U24806 (N_24806,N_22498,N_21479);
xnor U24807 (N_24807,N_21177,N_20819);
and U24808 (N_24808,N_22368,N_21666);
xnor U24809 (N_24809,N_20671,N_20210);
xor U24810 (N_24810,N_20334,N_20536);
nand U24811 (N_24811,N_20016,N_21225);
nand U24812 (N_24812,N_21610,N_20664);
or U24813 (N_24813,N_21749,N_20721);
nor U24814 (N_24814,N_20742,N_20938);
and U24815 (N_24815,N_22252,N_20760);
xnor U24816 (N_24816,N_22190,N_20040);
xnor U24817 (N_24817,N_21350,N_21120);
xor U24818 (N_24818,N_21200,N_21095);
nor U24819 (N_24819,N_21870,N_20279);
or U24820 (N_24820,N_20143,N_20745);
or U24821 (N_24821,N_21278,N_21397);
or U24822 (N_24822,N_22435,N_21993);
xnor U24823 (N_24823,N_20690,N_20826);
nand U24824 (N_24824,N_21225,N_21044);
or U24825 (N_24825,N_21830,N_21161);
or U24826 (N_24826,N_22372,N_22198);
nor U24827 (N_24827,N_22482,N_22389);
and U24828 (N_24828,N_20764,N_21069);
or U24829 (N_24829,N_20606,N_20201);
or U24830 (N_24830,N_21062,N_20356);
and U24831 (N_24831,N_20846,N_20398);
nand U24832 (N_24832,N_22121,N_21447);
and U24833 (N_24833,N_21608,N_22293);
xor U24834 (N_24834,N_21527,N_22064);
nor U24835 (N_24835,N_20366,N_20902);
or U24836 (N_24836,N_22090,N_22373);
nand U24837 (N_24837,N_20156,N_20115);
nand U24838 (N_24838,N_21291,N_21748);
nor U24839 (N_24839,N_21675,N_21179);
and U24840 (N_24840,N_21124,N_21696);
and U24841 (N_24841,N_20091,N_20058);
or U24842 (N_24842,N_21023,N_20022);
or U24843 (N_24843,N_21712,N_21353);
nand U24844 (N_24844,N_22344,N_22378);
nor U24845 (N_24845,N_20044,N_22267);
or U24846 (N_24846,N_20530,N_22177);
nand U24847 (N_24847,N_20524,N_22341);
and U24848 (N_24848,N_20306,N_22358);
nor U24849 (N_24849,N_22390,N_21506);
nand U24850 (N_24850,N_21104,N_21818);
and U24851 (N_24851,N_21378,N_21175);
nand U24852 (N_24852,N_21124,N_22177);
or U24853 (N_24853,N_21946,N_21073);
and U24854 (N_24854,N_21150,N_20248);
xnor U24855 (N_24855,N_21695,N_20564);
nand U24856 (N_24856,N_21817,N_21931);
and U24857 (N_24857,N_20542,N_21408);
and U24858 (N_24858,N_21317,N_21860);
nor U24859 (N_24859,N_21257,N_22186);
xnor U24860 (N_24860,N_21792,N_22466);
nand U24861 (N_24861,N_20566,N_20838);
and U24862 (N_24862,N_21474,N_21282);
and U24863 (N_24863,N_20137,N_21424);
or U24864 (N_24864,N_20303,N_21586);
and U24865 (N_24865,N_22276,N_22198);
xor U24866 (N_24866,N_21303,N_21316);
nand U24867 (N_24867,N_21242,N_21909);
nand U24868 (N_24868,N_22123,N_20923);
nor U24869 (N_24869,N_20452,N_20640);
nor U24870 (N_24870,N_21495,N_21863);
xor U24871 (N_24871,N_20580,N_21317);
or U24872 (N_24872,N_21812,N_22335);
or U24873 (N_24873,N_20245,N_20085);
nand U24874 (N_24874,N_20151,N_22069);
and U24875 (N_24875,N_20579,N_20605);
or U24876 (N_24876,N_20067,N_21754);
xor U24877 (N_24877,N_22090,N_22274);
xor U24878 (N_24878,N_22046,N_20384);
nor U24879 (N_24879,N_21948,N_21357);
or U24880 (N_24880,N_21115,N_21347);
nor U24881 (N_24881,N_22191,N_21081);
or U24882 (N_24882,N_21040,N_20458);
nand U24883 (N_24883,N_21964,N_21240);
and U24884 (N_24884,N_20063,N_20900);
nand U24885 (N_24885,N_20155,N_20764);
or U24886 (N_24886,N_21431,N_21349);
or U24887 (N_24887,N_21881,N_20152);
or U24888 (N_24888,N_20911,N_21697);
or U24889 (N_24889,N_21684,N_20146);
and U24890 (N_24890,N_20533,N_20801);
nand U24891 (N_24891,N_21518,N_21164);
and U24892 (N_24892,N_21870,N_20633);
xnor U24893 (N_24893,N_22022,N_21076);
xor U24894 (N_24894,N_21606,N_21075);
nor U24895 (N_24895,N_22439,N_22427);
nor U24896 (N_24896,N_20551,N_21665);
nor U24897 (N_24897,N_20143,N_20338);
nand U24898 (N_24898,N_20131,N_20881);
and U24899 (N_24899,N_21585,N_20335);
nor U24900 (N_24900,N_20823,N_20273);
or U24901 (N_24901,N_21146,N_21895);
nor U24902 (N_24902,N_21492,N_20207);
or U24903 (N_24903,N_21104,N_20149);
or U24904 (N_24904,N_22405,N_21716);
nand U24905 (N_24905,N_20232,N_21613);
or U24906 (N_24906,N_21484,N_20382);
and U24907 (N_24907,N_21596,N_20160);
nand U24908 (N_24908,N_21324,N_20005);
or U24909 (N_24909,N_22437,N_21133);
nor U24910 (N_24910,N_20210,N_20988);
and U24911 (N_24911,N_20032,N_22450);
or U24912 (N_24912,N_21913,N_21580);
nand U24913 (N_24913,N_20510,N_20360);
or U24914 (N_24914,N_21286,N_21910);
and U24915 (N_24915,N_20910,N_20396);
or U24916 (N_24916,N_21240,N_22434);
nand U24917 (N_24917,N_20471,N_22048);
xor U24918 (N_24918,N_21552,N_22212);
and U24919 (N_24919,N_21377,N_22191);
nor U24920 (N_24920,N_21330,N_20642);
nand U24921 (N_24921,N_20714,N_22490);
nor U24922 (N_24922,N_21027,N_20869);
xnor U24923 (N_24923,N_21743,N_20364);
and U24924 (N_24924,N_21358,N_21089);
or U24925 (N_24925,N_20466,N_20877);
or U24926 (N_24926,N_20298,N_21710);
nand U24927 (N_24927,N_21289,N_20583);
or U24928 (N_24928,N_20719,N_22159);
and U24929 (N_24929,N_20938,N_20780);
or U24930 (N_24930,N_20610,N_20203);
nor U24931 (N_24931,N_21383,N_21528);
xor U24932 (N_24932,N_21799,N_21770);
and U24933 (N_24933,N_22381,N_21766);
and U24934 (N_24934,N_20289,N_20874);
or U24935 (N_24935,N_20533,N_22177);
xnor U24936 (N_24936,N_22441,N_21044);
and U24937 (N_24937,N_22135,N_21821);
and U24938 (N_24938,N_22122,N_20245);
nand U24939 (N_24939,N_21021,N_21194);
xor U24940 (N_24940,N_21270,N_20342);
and U24941 (N_24941,N_22208,N_20377);
nand U24942 (N_24942,N_22497,N_20332);
and U24943 (N_24943,N_21295,N_21566);
and U24944 (N_24944,N_21325,N_21423);
xnor U24945 (N_24945,N_21732,N_21901);
and U24946 (N_24946,N_21294,N_21762);
xor U24947 (N_24947,N_21747,N_21954);
and U24948 (N_24948,N_21643,N_22271);
xnor U24949 (N_24949,N_22317,N_22125);
and U24950 (N_24950,N_21720,N_22187);
and U24951 (N_24951,N_20709,N_21985);
and U24952 (N_24952,N_20931,N_21845);
nor U24953 (N_24953,N_21156,N_21518);
xor U24954 (N_24954,N_20600,N_20674);
nor U24955 (N_24955,N_21990,N_20973);
xor U24956 (N_24956,N_21441,N_21847);
xor U24957 (N_24957,N_21254,N_20964);
nor U24958 (N_24958,N_20014,N_22105);
or U24959 (N_24959,N_21435,N_21062);
nor U24960 (N_24960,N_22316,N_20817);
and U24961 (N_24961,N_22010,N_21330);
nand U24962 (N_24962,N_21385,N_21386);
nor U24963 (N_24963,N_20436,N_21482);
and U24964 (N_24964,N_20083,N_22084);
or U24965 (N_24965,N_20477,N_20918);
nor U24966 (N_24966,N_22151,N_21543);
nor U24967 (N_24967,N_21684,N_21879);
or U24968 (N_24968,N_22112,N_20787);
and U24969 (N_24969,N_20663,N_21190);
xnor U24970 (N_24970,N_22192,N_20923);
nor U24971 (N_24971,N_22206,N_21956);
xor U24972 (N_24972,N_20473,N_21058);
xnor U24973 (N_24973,N_21927,N_21556);
nor U24974 (N_24974,N_20257,N_22002);
nand U24975 (N_24975,N_22016,N_21317);
nand U24976 (N_24976,N_20906,N_20695);
nand U24977 (N_24977,N_22445,N_21507);
or U24978 (N_24978,N_21752,N_22366);
nand U24979 (N_24979,N_22399,N_20906);
nand U24980 (N_24980,N_21016,N_20459);
nor U24981 (N_24981,N_21749,N_21876);
nand U24982 (N_24982,N_21463,N_20845);
nor U24983 (N_24983,N_21394,N_20756);
and U24984 (N_24984,N_21736,N_22327);
nand U24985 (N_24985,N_20002,N_21973);
nand U24986 (N_24986,N_20576,N_21198);
nand U24987 (N_24987,N_21708,N_21866);
or U24988 (N_24988,N_20123,N_21752);
nor U24989 (N_24989,N_20409,N_21330);
xor U24990 (N_24990,N_20520,N_22296);
or U24991 (N_24991,N_22316,N_21136);
nor U24992 (N_24992,N_21652,N_22214);
xor U24993 (N_24993,N_20353,N_20847);
nor U24994 (N_24994,N_20966,N_20019);
nor U24995 (N_24995,N_21914,N_20290);
nor U24996 (N_24996,N_21088,N_21602);
nor U24997 (N_24997,N_21448,N_22056);
or U24998 (N_24998,N_21013,N_21196);
nor U24999 (N_24999,N_21882,N_21746);
or U25000 (N_25000,N_22861,N_24506);
xor U25001 (N_25001,N_23451,N_22663);
xnor U25002 (N_25002,N_24769,N_23220);
and U25003 (N_25003,N_23677,N_24205);
xnor U25004 (N_25004,N_23455,N_23438);
and U25005 (N_25005,N_23461,N_23803);
nand U25006 (N_25006,N_22649,N_22779);
or U25007 (N_25007,N_23727,N_24005);
nor U25008 (N_25008,N_22599,N_23067);
nand U25009 (N_25009,N_24496,N_22659);
nor U25010 (N_25010,N_22627,N_22672);
nor U25011 (N_25011,N_23215,N_22676);
nor U25012 (N_25012,N_23201,N_24728);
xnor U25013 (N_25013,N_24214,N_24000);
or U25014 (N_25014,N_22966,N_24433);
xor U25015 (N_25015,N_23753,N_24550);
or U25016 (N_25016,N_24579,N_23573);
or U25017 (N_25017,N_24782,N_23048);
xor U25018 (N_25018,N_23761,N_24501);
nor U25019 (N_25019,N_23975,N_23935);
xnor U25020 (N_25020,N_24658,N_24617);
xnor U25021 (N_25021,N_24291,N_23366);
nand U25022 (N_25022,N_22588,N_23113);
or U25023 (N_25023,N_22786,N_24230);
or U25024 (N_25024,N_22681,N_23069);
nor U25025 (N_25025,N_22541,N_24806);
and U25026 (N_25026,N_24355,N_23190);
xnor U25027 (N_25027,N_24905,N_23966);
xor U25028 (N_25028,N_23791,N_23183);
nand U25029 (N_25029,N_24545,N_24553);
and U25030 (N_25030,N_23167,N_24758);
xor U25031 (N_25031,N_24733,N_24389);
or U25032 (N_25032,N_22893,N_24079);
nor U25033 (N_25033,N_22742,N_23592);
nand U25034 (N_25034,N_24700,N_24390);
or U25035 (N_25035,N_22698,N_23572);
nand U25036 (N_25036,N_22558,N_23867);
nor U25037 (N_25037,N_23529,N_23468);
nand U25038 (N_25038,N_23619,N_24591);
nand U25039 (N_25039,N_24552,N_23017);
and U25040 (N_25040,N_24116,N_24138);
nor U25041 (N_25041,N_24858,N_23551);
nand U25042 (N_25042,N_23784,N_24075);
nor U25043 (N_25043,N_23528,N_24041);
nor U25044 (N_25044,N_24266,N_23777);
nor U25045 (N_25045,N_23846,N_22655);
nand U25046 (N_25046,N_22868,N_23748);
and U25047 (N_25047,N_22835,N_24683);
xor U25048 (N_25048,N_24687,N_23842);
xnor U25049 (N_25049,N_22890,N_23974);
nand U25050 (N_25050,N_22833,N_23755);
or U25051 (N_25051,N_24673,N_24292);
or U25052 (N_25052,N_24654,N_24734);
nand U25053 (N_25053,N_23499,N_23374);
or U25054 (N_25054,N_23238,N_23819);
nand U25055 (N_25055,N_22678,N_22842);
and U25056 (N_25056,N_23825,N_23298);
xor U25057 (N_25057,N_24463,N_24601);
and U25058 (N_25058,N_24935,N_24805);
nand U25059 (N_25059,N_22554,N_24678);
and U25060 (N_25060,N_23149,N_22756);
and U25061 (N_25061,N_23599,N_24690);
nand U25062 (N_25062,N_23684,N_24134);
nand U25063 (N_25063,N_23005,N_22725);
nor U25064 (N_25064,N_22917,N_24794);
nor U25065 (N_25065,N_23348,N_24454);
or U25066 (N_25066,N_24539,N_23914);
or U25067 (N_25067,N_22899,N_22507);
or U25068 (N_25068,N_23336,N_23603);
or U25069 (N_25069,N_23887,N_23273);
or U25070 (N_25070,N_24692,N_22533);
nand U25071 (N_25071,N_24816,N_23924);
and U25072 (N_25072,N_24367,N_24953);
xnor U25073 (N_25073,N_23085,N_23396);
nand U25074 (N_25074,N_23503,N_23895);
nand U25075 (N_25075,N_23504,N_24476);
xnor U25076 (N_25076,N_22812,N_23849);
nor U25077 (N_25077,N_24263,N_24333);
nor U25078 (N_25078,N_24376,N_23870);
or U25079 (N_25079,N_23088,N_23591);
nor U25080 (N_25080,N_24561,N_24066);
nand U25081 (N_25081,N_23200,N_22780);
and U25082 (N_25082,N_24373,N_22894);
nor U25083 (N_25083,N_24779,N_22668);
or U25084 (N_25084,N_24439,N_24098);
or U25085 (N_25085,N_23831,N_22568);
or U25086 (N_25086,N_24135,N_24767);
nor U25087 (N_25087,N_24440,N_24809);
and U25088 (N_25088,N_23590,N_24613);
or U25089 (N_25089,N_23737,N_24147);
nor U25090 (N_25090,N_22903,N_24069);
xor U25091 (N_25091,N_22956,N_22595);
nand U25092 (N_25092,N_22854,N_22777);
nor U25093 (N_25093,N_23342,N_22590);
nand U25094 (N_25094,N_22945,N_22845);
nor U25095 (N_25095,N_24954,N_23557);
or U25096 (N_25096,N_23163,N_24231);
nor U25097 (N_25097,N_23637,N_22712);
and U25098 (N_25098,N_22720,N_23743);
and U25099 (N_25099,N_22506,N_23493);
xor U25100 (N_25100,N_23520,N_23286);
or U25101 (N_25101,N_23968,N_22578);
or U25102 (N_25102,N_24896,N_23308);
and U25103 (N_25103,N_23302,N_24639);
nor U25104 (N_25104,N_22865,N_23064);
nand U25105 (N_25105,N_22788,N_23459);
and U25106 (N_25106,N_23317,N_23061);
or U25107 (N_25107,N_23478,N_23740);
and U25108 (N_25108,N_23577,N_24795);
xor U25109 (N_25109,N_24818,N_24270);
or U25110 (N_25110,N_24090,N_23567);
nor U25111 (N_25111,N_24691,N_23343);
or U25112 (N_25112,N_24260,N_24777);
nand U25113 (N_25113,N_23800,N_24973);
xor U25114 (N_25114,N_23664,N_24558);
nand U25115 (N_25115,N_23647,N_24473);
or U25116 (N_25116,N_23383,N_23741);
and U25117 (N_25117,N_24120,N_22616);
nor U25118 (N_25118,N_24479,N_24073);
nand U25119 (N_25119,N_24760,N_24108);
xor U25120 (N_25120,N_22792,N_24398);
and U25121 (N_25121,N_23834,N_24856);
nor U25122 (N_25122,N_23646,N_24505);
and U25123 (N_25123,N_23119,N_24036);
nor U25124 (N_25124,N_23414,N_23514);
or U25125 (N_25125,N_22796,N_24302);
nand U25126 (N_25126,N_23227,N_23291);
nor U25127 (N_25127,N_23062,N_22722);
nand U25128 (N_25128,N_22939,N_22948);
or U25129 (N_25129,N_23435,N_24308);
nor U25130 (N_25130,N_22751,N_22933);
or U25131 (N_25131,N_23845,N_24634);
nand U25132 (N_25132,N_24877,N_22697);
xnor U25133 (N_25133,N_22920,N_22888);
and U25134 (N_25134,N_23057,N_24406);
or U25135 (N_25135,N_23657,N_23415);
and U25136 (N_25136,N_24365,N_24277);
nand U25137 (N_25137,N_23594,N_24414);
xnor U25138 (N_25138,N_23222,N_22858);
nand U25139 (N_25139,N_22885,N_23606);
nor U25140 (N_25140,N_23103,N_23548);
xnor U25141 (N_25141,N_23159,N_24698);
or U25142 (N_25142,N_23033,N_24922);
nand U25143 (N_25143,N_22638,N_24722);
nand U25144 (N_25144,N_24282,N_22843);
xnor U25145 (N_25145,N_24768,N_24570);
nand U25146 (N_25146,N_22863,N_22636);
xor U25147 (N_25147,N_22944,N_22693);
nand U25148 (N_25148,N_23705,N_24290);
or U25149 (N_25149,N_24730,N_22852);
xnor U25150 (N_25150,N_24857,N_24085);
and U25151 (N_25151,N_24494,N_24220);
and U25152 (N_25152,N_23077,N_23002);
xnor U25153 (N_25153,N_24188,N_24315);
and U25154 (N_25154,N_24024,N_23367);
and U25155 (N_25155,N_24656,N_22776);
xnor U25156 (N_25156,N_22910,N_23984);
xnor U25157 (N_25157,N_22529,N_24737);
and U25158 (N_25158,N_24182,N_24747);
or U25159 (N_25159,N_23198,N_23771);
nand U25160 (N_25160,N_23875,N_24250);
and U25161 (N_25161,N_24206,N_23477);
xnor U25162 (N_25162,N_24055,N_23956);
and U25163 (N_25163,N_23563,N_23538);
nand U25164 (N_25164,N_23155,N_23495);
nand U25165 (N_25165,N_22979,N_22584);
xor U25166 (N_25166,N_24094,N_24299);
or U25167 (N_25167,N_23526,N_24169);
nor U25168 (N_25168,N_23187,N_22930);
nor U25169 (N_25169,N_24559,N_23651);
xor U25170 (N_25170,N_23392,N_22550);
or U25171 (N_25171,N_22935,N_24287);
nand U25172 (N_25172,N_23742,N_24099);
nand U25173 (N_25173,N_24364,N_24710);
xor U25174 (N_25174,N_23690,N_23643);
or U25175 (N_25175,N_23445,N_24172);
nor U25176 (N_25176,N_24585,N_23472);
nand U25177 (N_25177,N_23624,N_23991);
nor U25178 (N_25178,N_22700,N_23211);
xor U25179 (N_25179,N_24633,N_23213);
xnor U25180 (N_25180,N_22901,N_23282);
nand U25181 (N_25181,N_24604,N_22962);
or U25182 (N_25182,N_24838,N_23714);
or U25183 (N_25183,N_23506,N_23447);
xnor U25184 (N_25184,N_23158,N_24681);
nand U25185 (N_25185,N_24577,N_24101);
or U25186 (N_25186,N_23919,N_24859);
and U25187 (N_25187,N_23145,N_23874);
nor U25188 (N_25188,N_23066,N_24898);
xor U25189 (N_25189,N_23332,N_22977);
and U25190 (N_25190,N_22664,N_23857);
xnor U25191 (N_25191,N_24117,N_24648);
nand U25192 (N_25192,N_24983,N_23723);
and U25193 (N_25193,N_22582,N_24474);
nor U25194 (N_25194,N_23247,N_23494);
nand U25195 (N_25195,N_22932,N_24798);
and U25196 (N_25196,N_22696,N_24401);
nor U25197 (N_25197,N_22889,N_22791);
and U25198 (N_25198,N_24854,N_23010);
or U25199 (N_25199,N_22512,N_22784);
and U25200 (N_25200,N_22807,N_24142);
or U25201 (N_25201,N_23147,N_23071);
and U25202 (N_25202,N_24209,N_24426);
and U25203 (N_25203,N_24227,N_23667);
or U25204 (N_25204,N_23299,N_22973);
nand U25205 (N_25205,N_24104,N_23574);
and U25206 (N_25206,N_23822,N_22954);
and U25207 (N_25207,N_23231,N_24486);
or U25208 (N_25208,N_23878,N_23533);
or U25209 (N_25209,N_24490,N_22654);
and U25210 (N_25210,N_24933,N_23007);
and U25211 (N_25211,N_23688,N_23386);
nand U25212 (N_25212,N_23369,N_24669);
nor U25213 (N_25213,N_24920,N_23730);
or U25214 (N_25214,N_23865,N_23821);
nand U25215 (N_25215,N_24304,N_23703);
nor U25216 (N_25216,N_24504,N_23859);
xor U25217 (N_25217,N_24238,N_24014);
xnor U25218 (N_25218,N_24595,N_22774);
nor U25219 (N_25219,N_24129,N_24919);
xnor U25220 (N_25220,N_23123,N_24848);
xnor U25221 (N_25221,N_23818,N_23905);
and U25222 (N_25222,N_22574,N_23540);
nor U25223 (N_25223,N_22704,N_22591);
or U25224 (N_25224,N_24672,N_23259);
xnor U25225 (N_25225,N_24774,N_22794);
nand U25226 (N_25226,N_23549,N_24438);
nor U25227 (N_25227,N_22614,N_23118);
nand U25228 (N_25228,N_24589,N_23104);
and U25229 (N_25229,N_23823,N_24598);
xnor U25230 (N_25230,N_24314,N_22949);
nor U25231 (N_25231,N_24067,N_24403);
nor U25232 (N_25232,N_22543,N_24921);
and U25233 (N_25233,N_23334,N_23749);
or U25234 (N_25234,N_22740,N_23694);
nor U25235 (N_25235,N_24757,N_23604);
or U25236 (N_25236,N_22708,N_23294);
or U25237 (N_25237,N_24471,N_23902);
and U25238 (N_25238,N_23600,N_23125);
nand U25239 (N_25239,N_23307,N_23004);
xnor U25240 (N_25240,N_23138,N_22919);
or U25241 (N_25241,N_24432,N_24118);
or U25242 (N_25242,N_24624,N_22563);
nand U25243 (N_25243,N_22675,N_23735);
and U25244 (N_25244,N_24420,N_23691);
xor U25245 (N_25245,N_22832,N_24374);
or U25246 (N_25246,N_23841,N_24799);
xnor U25247 (N_25247,N_24849,N_23426);
nand U25248 (N_25248,N_23869,N_23612);
and U25249 (N_25249,N_22746,N_23750);
or U25250 (N_25250,N_22719,N_23253);
or U25251 (N_25251,N_23279,N_23744);
or U25252 (N_25252,N_23850,N_22866);
nor U25253 (N_25253,N_23847,N_22934);
nand U25254 (N_25254,N_24917,N_23450);
nand U25255 (N_25255,N_22647,N_24133);
nor U25256 (N_25256,N_24960,N_23745);
xor U25257 (N_25257,N_23958,N_24415);
and U25258 (N_25258,N_23693,N_23434);
nand U25259 (N_25259,N_24725,N_24833);
or U25260 (N_25260,N_22619,N_22749);
or U25261 (N_25261,N_24186,N_23997);
and U25262 (N_25262,N_22705,N_23801);
xnor U25263 (N_25263,N_22994,N_24430);
nand U25264 (N_25264,N_24939,N_23797);
xnor U25265 (N_25265,N_23285,N_24265);
and U25266 (N_25266,N_24045,N_24904);
or U25267 (N_25267,N_23006,N_23805);
nor U25268 (N_25268,N_22798,N_22823);
xnor U25269 (N_25269,N_24313,N_23030);
nor U25270 (N_25270,N_22646,N_23830);
nand U25271 (N_25271,N_22844,N_23661);
xor U25272 (N_25272,N_24622,N_24636);
and U25273 (N_25273,N_23152,N_23115);
nand U25274 (N_25274,N_24942,N_24663);
nor U25275 (N_25275,N_23542,N_24618);
xnor U25276 (N_25276,N_23385,N_24033);
xor U25277 (N_25277,N_24294,N_24827);
nor U25278 (N_25278,N_24808,N_24867);
xnor U25279 (N_25279,N_23794,N_24985);
nor U25280 (N_25280,N_24458,N_24635);
nor U25281 (N_25281,N_23787,N_24309);
nand U25282 (N_25282,N_23463,N_24732);
nor U25283 (N_25283,N_24358,N_24177);
nor U25284 (N_25284,N_24351,N_23656);
nand U25285 (N_25285,N_23880,N_22905);
nand U25286 (N_25286,N_23901,N_24223);
nand U25287 (N_25287,N_24168,N_22970);
and U25288 (N_25288,N_23150,N_23546);
nor U25289 (N_25289,N_23885,N_22955);
nand U25290 (N_25290,N_23981,N_23863);
nand U25291 (N_25291,N_23862,N_24517);
nor U25292 (N_25292,N_22797,N_23673);
and U25293 (N_25293,N_23252,N_24652);
and U25294 (N_25294,N_22817,N_24608);
nor U25295 (N_25295,N_24100,N_24512);
and U25296 (N_25296,N_23474,N_23733);
nor U25297 (N_25297,N_24707,N_23970);
and U25298 (N_25298,N_23233,N_23593);
nor U25299 (N_25299,N_24802,N_24864);
and U25300 (N_25300,N_24980,N_22617);
nand U25301 (N_25301,N_23934,N_22565);
xnor U25302 (N_25302,N_23040,N_24926);
xor U25303 (N_25303,N_22625,N_24123);
nand U25304 (N_25304,N_23918,N_24300);
nand U25305 (N_25305,N_22660,N_24880);
nand U25306 (N_25306,N_23012,N_22810);
and U25307 (N_25307,N_22583,N_23930);
nor U25308 (N_25308,N_22857,N_23925);
nand U25309 (N_25309,N_22562,N_22771);
nor U25310 (N_25310,N_24058,N_22897);
nor U25311 (N_25311,N_23602,N_22609);
nand U25312 (N_25312,N_24083,N_24044);
nand U25313 (N_25313,N_22764,N_24026);
or U25314 (N_25314,N_24199,N_23219);
or U25315 (N_25315,N_24019,N_24952);
xor U25316 (N_25316,N_24679,N_24711);
nor U25317 (N_25317,N_23676,N_24957);
or U25318 (N_25318,N_24784,N_24626);
or U25319 (N_25319,N_23711,N_23817);
xnor U25320 (N_25320,N_24137,N_23789);
xor U25321 (N_25321,N_24434,N_22605);
nor U25322 (N_25322,N_23462,N_24006);
xor U25323 (N_25323,N_23939,N_23700);
nor U25324 (N_25324,N_22772,N_23382);
nand U25325 (N_25325,N_22587,N_22753);
xor U25326 (N_25326,N_24200,N_23900);
or U25327 (N_25327,N_22913,N_23413);
xor U25328 (N_25328,N_23024,N_23621);
or U25329 (N_25329,N_24261,N_24824);
nor U25330 (N_25330,N_22846,N_23756);
and U25331 (N_25331,N_23195,N_23804);
nand U25332 (N_25332,N_24705,N_23370);
xor U25333 (N_25333,N_22701,N_22855);
xnor U25334 (N_25334,N_24551,N_23708);
nor U25335 (N_25335,N_23553,N_24825);
and U25336 (N_25336,N_24927,N_24885);
xor U25337 (N_25337,N_23028,N_24916);
and U25338 (N_25338,N_24071,N_23019);
nand U25339 (N_25339,N_23671,N_24457);
xnor U25340 (N_25340,N_24720,N_24978);
or U25341 (N_25341,N_23508,N_24152);
xor U25342 (N_25342,N_23047,N_24422);
nor U25343 (N_25343,N_23571,N_24937);
xor U25344 (N_25344,N_23390,N_23683);
nand U25345 (N_25345,N_23223,N_23160);
nand U25346 (N_25346,N_24107,N_24670);
or U25347 (N_25347,N_22514,N_22633);
and U25348 (N_25348,N_24323,N_24792);
xor U25349 (N_25349,N_22824,N_22853);
xor U25350 (N_25350,N_22782,N_23512);
xnor U25351 (N_25351,N_23449,N_23073);
nor U25352 (N_25352,N_24326,N_22989);
nor U25353 (N_25353,N_24031,N_23486);
xnor U25354 (N_25354,N_24240,N_24424);
nand U25355 (N_25355,N_24130,N_24567);
or U25356 (N_25356,N_23992,N_22508);
nor U25357 (N_25357,N_24832,N_23456);
nor U25358 (N_25358,N_23853,N_23217);
or U25359 (N_25359,N_23126,N_23908);
or U25360 (N_25360,N_23100,N_24187);
xor U25361 (N_25361,N_24537,N_22602);
nor U25362 (N_25362,N_23243,N_23613);
or U25363 (N_25363,N_23957,N_22809);
nand U25364 (N_25364,N_22570,N_23829);
xnor U25365 (N_25365,N_23584,N_24191);
xnor U25366 (N_25366,N_24081,N_24882);
and U25367 (N_25367,N_24763,N_23751);
and U25368 (N_25368,N_23096,N_24468);
or U25369 (N_25369,N_24103,N_23547);
nand U25370 (N_25370,N_24274,N_24462);
nor U25371 (N_25371,N_23060,N_23176);
nor U25372 (N_25372,N_24482,N_22735);
and U25373 (N_25373,N_23785,N_24571);
nor U25374 (N_25374,N_24455,N_23263);
and U25375 (N_25375,N_23099,N_24534);
xnor U25376 (N_25376,N_23162,N_24127);
nor U25377 (N_25377,N_24740,N_24106);
xnor U25378 (N_25378,N_22959,N_22790);
and U25379 (N_25379,N_22608,N_24331);
xor U25380 (N_25380,N_23178,N_23587);
and U25381 (N_25381,N_23431,N_24507);
xnor U25382 (N_25382,N_23632,N_22838);
xor U25383 (N_25383,N_24158,N_23618);
nand U25384 (N_25384,N_24350,N_23555);
or U25385 (N_25385,N_22527,N_24021);
and U25386 (N_25386,N_22581,N_24427);
nand U25387 (N_25387,N_24716,N_22811);
or U25388 (N_25388,N_22680,N_24979);
or U25389 (N_25389,N_24091,N_23649);
xnor U25390 (N_25390,N_22656,N_22523);
nand U25391 (N_25391,N_22569,N_22951);
and U25392 (N_25392,N_24377,N_23582);
and U25393 (N_25393,N_24157,N_24017);
and U25394 (N_25394,N_23543,N_23391);
or U25395 (N_25395,N_23454,N_22825);
and U25396 (N_25396,N_24050,N_24043);
nor U25397 (N_25397,N_24170,N_24337);
nor U25398 (N_25398,N_23325,N_22561);
xnor U25399 (N_25399,N_23835,N_23368);
or U25400 (N_25400,N_23436,N_23883);
or U25401 (N_25401,N_22500,N_23402);
or U25402 (N_25402,N_23045,N_24362);
nor U25403 (N_25403,N_23046,N_22830);
or U25404 (N_25404,N_23614,N_22585);
nand U25405 (N_25405,N_23311,N_23575);
or U25406 (N_25406,N_24185,N_23535);
xor U25407 (N_25407,N_24623,N_23026);
xnor U25408 (N_25408,N_23906,N_24801);
nor U25409 (N_25409,N_23009,N_22610);
or U25410 (N_25410,N_24475,N_24583);
nor U25411 (N_25411,N_22606,N_23722);
nand U25412 (N_25412,N_23907,N_24823);
nand U25413 (N_25413,N_24023,N_24759);
and U25414 (N_25414,N_24297,N_23168);
nor U25415 (N_25415,N_24460,N_22960);
nand U25416 (N_25416,N_24369,N_24602);
nor U25417 (N_25417,N_23469,N_23429);
or U25418 (N_25418,N_23692,N_24229);
or U25419 (N_25419,N_23892,N_23080);
nand U25420 (N_25420,N_22634,N_22626);
and U25421 (N_25421,N_22723,N_23419);
xor U25422 (N_25422,N_24176,N_24407);
or U25423 (N_25423,N_22566,N_23824);
nand U25424 (N_25424,N_23287,N_22537);
nand U25425 (N_25425,N_22938,N_22998);
nor U25426 (N_25426,N_23645,N_23278);
and U25427 (N_25427,N_23097,N_23458);
nor U25428 (N_25428,N_24655,N_22873);
and U25429 (N_25429,N_24755,N_23362);
or U25430 (N_25430,N_23716,N_24410);
nand U25431 (N_25431,N_23037,N_23866);
or U25432 (N_25432,N_24876,N_24568);
or U25433 (N_25433,N_24908,N_23254);
and U25434 (N_25434,N_23679,N_23623);
nand U25435 (N_25435,N_24616,N_23815);
nand U25436 (N_25436,N_23795,N_23265);
nand U25437 (N_25437,N_24975,N_23448);
and U25438 (N_25438,N_23164,N_24166);
and U25439 (N_25439,N_23654,N_24564);
nor U25440 (N_25440,N_24444,N_23399);
nand U25441 (N_25441,N_23739,N_24712);
xnor U25442 (N_25442,N_24531,N_23442);
and U25443 (N_25443,N_22971,N_22849);
nand U25444 (N_25444,N_24371,N_22926);
and U25445 (N_25445,N_24829,N_24888);
nor U25446 (N_25446,N_23305,N_24027);
nand U25447 (N_25447,N_22726,N_22769);
nor U25448 (N_25448,N_23359,N_24140);
nor U25449 (N_25449,N_24347,N_24521);
xor U25450 (N_25450,N_23562,N_24007);
nor U25451 (N_25451,N_24820,N_24442);
nor U25452 (N_25452,N_22884,N_23146);
and U25453 (N_25453,N_22921,N_23439);
nand U25454 (N_25454,N_24153,N_24605);
or U25455 (N_25455,N_22773,N_22652);
xnor U25456 (N_25456,N_23094,N_23515);
nor U25457 (N_25457,N_23773,N_23728);
and U25458 (N_25458,N_22691,N_24162);
or U25459 (N_25459,N_24491,N_23297);
or U25460 (N_25460,N_24503,N_22642);
and U25461 (N_25461,N_24217,N_23827);
nand U25462 (N_25462,N_22556,N_24252);
and U25463 (N_25463,N_22732,N_22848);
or U25464 (N_25464,N_23262,N_24974);
nand U25465 (N_25465,N_24180,N_24063);
and U25466 (N_25466,N_24630,N_23389);
and U25467 (N_25467,N_23052,N_23525);
and U25468 (N_25468,N_24074,N_22906);
or U25469 (N_25469,N_24837,N_24772);
nand U25470 (N_25470,N_24487,N_23709);
or U25471 (N_25471,N_24582,N_24020);
xnor U25472 (N_25472,N_24717,N_22631);
xnor U25473 (N_25473,N_24751,N_23086);
nand U25474 (N_25474,N_24542,N_23316);
xor U25475 (N_25475,N_24178,N_23492);
or U25476 (N_25476,N_23638,N_22997);
and U25477 (N_25477,N_24943,N_24596);
xnor U25478 (N_25478,N_23670,N_24619);
or U25479 (N_25479,N_22643,N_24388);
nand U25480 (N_25480,N_24597,N_24575);
or U25481 (N_25481,N_22763,N_23585);
or U25482 (N_25482,N_23102,N_23806);
nand U25483 (N_25483,N_23107,N_23781);
nor U25484 (N_25484,N_23281,N_23798);
nand U25485 (N_25485,N_24741,N_22531);
nand U25486 (N_25486,N_24171,N_23221);
nor U25487 (N_25487,N_22958,N_23877);
nand U25488 (N_25488,N_24516,N_23264);
xor U25489 (N_25489,N_24909,N_23633);
nor U25490 (N_25490,N_22628,N_23652);
xnor U25491 (N_25491,N_23020,N_24372);
xnor U25492 (N_25492,N_24453,N_24119);
or U25493 (N_25493,N_24184,N_23202);
nor U25494 (N_25494,N_24329,N_23078);
nand U25495 (N_25495,N_24883,N_23153);
or U25496 (N_25496,N_24286,N_23995);
nand U25497 (N_25497,N_24951,N_23425);
and U25498 (N_25498,N_22754,N_23736);
and U25499 (N_25499,N_24674,N_23199);
and U25500 (N_25500,N_22692,N_24399);
nor U25501 (N_25501,N_24251,N_23903);
xor U25502 (N_25502,N_24968,N_23489);
xor U25503 (N_25503,N_24914,N_23888);
nand U25504 (N_25504,N_23669,N_23464);
nor U25505 (N_25505,N_24533,N_23376);
nor U25506 (N_25506,N_24785,N_23860);
and U25507 (N_25507,N_23802,N_22645);
nor U25508 (N_25508,N_24895,N_22552);
nor U25509 (N_25509,N_23379,N_24484);
and U25510 (N_25510,N_22737,N_22503);
nor U25511 (N_25511,N_24148,N_22925);
or U25512 (N_25512,N_22657,N_24677);
and U25513 (N_25513,N_22878,N_22912);
and U25514 (N_25514,N_23081,N_23813);
nor U25515 (N_25515,N_22819,N_23851);
xnor U25516 (N_25516,N_24746,N_24621);
and U25517 (N_25517,N_24385,N_23566);
and U25518 (N_25518,N_23191,N_23890);
xnor U25519 (N_25519,N_24325,N_22651);
nand U25520 (N_25520,N_23365,N_23018);
and U25521 (N_25521,N_23128,N_22957);
or U25522 (N_25522,N_24843,N_24703);
and U25523 (N_25523,N_22761,N_24124);
xor U25524 (N_25524,N_23564,N_22621);
or U25525 (N_25525,N_23720,N_24901);
or U25526 (N_25526,N_23672,N_22721);
xor U25527 (N_25527,N_23290,N_23443);
nor U25528 (N_25528,N_23059,N_24042);
or U25529 (N_25529,N_23848,N_24940);
nor U25530 (N_25530,N_22891,N_23554);
or U25531 (N_25531,N_23837,N_23864);
nand U25532 (N_25532,N_24894,N_24029);
and U25533 (N_25533,N_23039,N_24773);
nand U25534 (N_25534,N_23154,N_23063);
and U25535 (N_25535,N_23023,N_24198);
nor U25536 (N_25536,N_24967,N_23886);
and U25537 (N_25537,N_24814,N_24334);
xnor U25538 (N_25538,N_24456,N_23142);
nand U25539 (N_25539,N_23569,N_22671);
nand U25540 (N_25540,N_23420,N_23397);
nand U25541 (N_25541,N_24999,N_22524);
nand U25542 (N_25542,N_24111,N_24844);
or U25543 (N_25543,N_23224,N_23036);
nand U25544 (N_25544,N_23350,N_24946);
nor U25545 (N_25545,N_23109,N_23891);
and U25546 (N_25546,N_23725,N_23707);
nor U25547 (N_25547,N_22923,N_24243);
nand U25548 (N_25548,N_24594,N_23375);
nand U25549 (N_25549,N_22694,N_23432);
and U25550 (N_25550,N_24990,N_24466);
or U25551 (N_25551,N_23347,N_24528);
nor U25552 (N_25552,N_22604,N_23774);
nand U25553 (N_25553,N_24899,N_23084);
and U25554 (N_25554,N_22673,N_22573);
nand U25555 (N_25555,N_23082,N_24037);
or U25556 (N_25556,N_24642,N_23595);
nand U25557 (N_25557,N_23457,N_22504);
or U25558 (N_25558,N_22870,N_22766);
xor U25559 (N_25559,N_23288,N_22978);
xnor U25560 (N_25560,N_24163,N_24327);
or U25561 (N_25561,N_23799,N_23648);
or U25562 (N_25562,N_23301,N_23516);
and U25563 (N_25563,N_23872,N_24721);
nor U25564 (N_25564,N_23346,N_23101);
nor U25565 (N_25565,N_24811,N_23986);
nor U25566 (N_25566,N_22516,N_24072);
or U25567 (N_25567,N_24102,N_22685);
and U25568 (N_25568,N_23793,N_22641);
nor U25569 (N_25569,N_24640,N_22778);
nor U25570 (N_25570,N_23556,N_24451);
nand U25571 (N_25571,N_24906,N_22632);
nor U25572 (N_25572,N_24324,N_23779);
nand U25573 (N_25573,N_23884,N_24524);
and U25574 (N_25574,N_23559,N_24813);
and U25575 (N_25575,N_23008,N_22887);
and U25576 (N_25576,N_24723,N_23129);
xnor U25577 (N_25577,N_24097,N_24393);
or U25578 (N_25578,N_24139,N_23873);
nor U25579 (N_25579,N_24514,N_24776);
nand U25580 (N_25580,N_23079,N_22898);
nor U25581 (N_25581,N_22501,N_22553);
and U25582 (N_25582,N_24408,N_22695);
nor U25583 (N_25583,N_23226,N_22505);
nand U25584 (N_25584,N_24413,N_23196);
nand U25585 (N_25585,N_22943,N_22598);
xor U25586 (N_25586,N_24646,N_23921);
or U25587 (N_25587,N_24500,N_22689);
xnor U25588 (N_25588,N_22867,N_22549);
and U25589 (N_25589,N_22580,N_23232);
or U25590 (N_25590,N_24082,N_23530);
xnor U25591 (N_25591,N_23240,N_24025);
or U25592 (N_25592,N_22814,N_23518);
nor U25593 (N_25593,N_22521,N_23214);
and U25594 (N_25594,N_24064,N_22759);
xor U25595 (N_25595,N_24345,N_24057);
or U25596 (N_25596,N_24208,N_24788);
xor U25597 (N_25597,N_23453,N_24167);
and U25598 (N_25598,N_24461,N_24929);
nor U25599 (N_25599,N_23678,N_22882);
nand U25600 (N_25600,N_24032,N_23858);
nor U25601 (N_25601,N_23732,N_23245);
and U25602 (N_25602,N_24949,N_24224);
nor U25603 (N_25603,N_22829,N_23446);
or U25604 (N_25604,N_24089,N_24497);
nand U25605 (N_25605,N_24984,N_23384);
xor U25606 (N_25606,N_22687,N_23193);
or U25607 (N_25607,N_24053,N_24892);
xor U25608 (N_25608,N_24095,N_24445);
nor U25609 (N_25609,N_24569,N_24890);
nor U25610 (N_25610,N_23625,N_24477);
xor U25611 (N_25611,N_23378,N_24532);
nand U25612 (N_25612,N_24870,N_24947);
xor U25613 (N_25613,N_23689,N_24836);
xor U25614 (N_25614,N_24271,N_24256);
and U25615 (N_25615,N_24873,N_23032);
xnor U25616 (N_25616,N_23973,N_23904);
nand U25617 (N_25617,N_23271,N_24643);
or U25618 (N_25618,N_24667,N_24418);
xor U25619 (N_25619,N_24826,N_24380);
or U25620 (N_25620,N_24012,N_23320);
or U25621 (N_25621,N_22667,N_24003);
xor U25622 (N_25622,N_23122,N_23581);
xor U25623 (N_25623,N_24803,N_24628);
nor U25624 (N_25624,N_23630,N_23854);
or U25625 (N_25625,N_23790,N_23373);
and U25626 (N_25626,N_23388,N_24241);
nor U25627 (N_25627,N_23424,N_23329);
or U25628 (N_25628,N_23717,N_23134);
and U25629 (N_25629,N_22999,N_22972);
and U25630 (N_25630,N_22679,N_23275);
or U25631 (N_25631,N_23133,N_23629);
and U25632 (N_25632,N_23879,N_24641);
nand U25633 (N_25633,N_24397,N_23626);
xor U25634 (N_25634,N_23117,N_23954);
xnor U25635 (N_25635,N_23042,N_22734);
and U25636 (N_25636,N_23210,N_24761);
or U25637 (N_25637,N_23184,N_24267);
nand U25638 (N_25638,N_23203,N_22575);
and U25639 (N_25639,N_23558,N_23016);
and U25640 (N_25640,N_24994,N_24499);
and U25641 (N_25641,N_22760,N_24666);
nand U25642 (N_25642,N_24987,N_24697);
xor U25643 (N_25643,N_24845,N_24540);
nor U25644 (N_25644,N_22744,N_22743);
and U25645 (N_25645,N_22927,N_23339);
nand U25646 (N_25646,N_24296,N_23565);
nand U25647 (N_25647,N_23927,N_24386);
xnor U25648 (N_25648,N_22834,N_22942);
nand U25649 (N_25649,N_23015,N_24659);
nand U25650 (N_25650,N_22787,N_23401);
or U25651 (N_25651,N_24931,N_22969);
xnor U25652 (N_25652,N_24684,N_24245);
and U25653 (N_25653,N_22594,N_23828);
or U25654 (N_25654,N_22800,N_24340);
nor U25655 (N_25655,N_24638,N_24047);
or U25656 (N_25656,N_23738,N_24748);
xnor U25657 (N_25657,N_24915,N_22991);
and U25658 (N_25658,N_24258,N_23072);
nand U25659 (N_25659,N_22896,N_24190);
nand U25660 (N_25660,N_23173,N_23121);
nand U25661 (N_25661,N_23055,N_23687);
and U25662 (N_25662,N_23928,N_23372);
nand U25663 (N_25663,N_24114,N_22674);
and U25664 (N_25664,N_22576,N_23810);
or U25665 (N_25665,N_23327,N_24912);
or U25666 (N_25666,N_22513,N_24918);
nor U25667 (N_25667,N_24611,N_23180);
xnor U25668 (N_25668,N_23112,N_24966);
xor U25669 (N_25669,N_24151,N_24498);
xnor U25670 (N_25670,N_23607,N_24196);
and U25671 (N_25671,N_24143,N_22789);
nand U25672 (N_25672,N_22929,N_23333);
nand U25673 (N_25673,N_24425,N_22551);
or U25674 (N_25674,N_24900,N_24657);
and U25675 (N_25675,N_23433,N_23519);
or U25676 (N_25676,N_22559,N_23729);
xor U25677 (N_25677,N_24587,N_24713);
or U25678 (N_25678,N_23760,N_23544);
and U25679 (N_25679,N_24213,N_22547);
or U25680 (N_25680,N_23274,N_23620);
xor U25681 (N_25681,N_23792,N_24964);
or U25682 (N_25682,N_23967,N_24753);
nand U25683 (N_25683,N_24273,N_24651);
nand U25684 (N_25684,N_23768,N_23759);
nand U25685 (N_25685,N_23955,N_23038);
and U25686 (N_25686,N_22711,N_23143);
nand U25687 (N_25687,N_23985,N_24714);
and U25688 (N_25688,N_22859,N_24727);
nor U25689 (N_25689,N_23812,N_23937);
nand U25690 (N_25690,N_24771,N_23951);
or U25691 (N_25691,N_24749,N_24972);
and U25692 (N_25692,N_24303,N_24828);
nor U25693 (N_25693,N_23165,N_23137);
and U25694 (N_25694,N_24417,N_23933);
xnor U25695 (N_25695,N_24936,N_23182);
nor U25696 (N_25696,N_24530,N_24841);
nor U25697 (N_25697,N_24804,N_23511);
and U25698 (N_25698,N_24335,N_23513);
or U25699 (N_25699,N_24378,N_23947);
nor U25700 (N_25700,N_24661,N_24357);
nand U25701 (N_25701,N_22729,N_24718);
nor U25702 (N_25702,N_24881,N_23898);
xnor U25703 (N_25703,N_22985,N_22546);
xnor U25704 (N_25704,N_22528,N_22532);
nand U25705 (N_25705,N_24520,N_24902);
nor U25706 (N_25706,N_24495,N_24481);
nand U25707 (N_25707,N_24402,N_22862);
and U25708 (N_25708,N_23502,N_23139);
nor U25709 (N_25709,N_23641,N_23277);
nor U25710 (N_25710,N_23931,N_24150);
and U25711 (N_25711,N_24181,N_23310);
and U25712 (N_25712,N_23208,N_23699);
or U25713 (N_25713,N_24056,N_22765);
and U25714 (N_25714,N_23653,N_23313);
or U25715 (N_25715,N_23280,N_24923);
xor U25716 (N_25716,N_23161,N_23982);
and U25717 (N_25717,N_24086,N_23093);
nor U25718 (N_25718,N_23911,N_23576);
nand U25719 (N_25719,N_24375,N_24179);
nor U25720 (N_25720,N_22597,N_22795);
nand U25721 (N_25721,N_22620,N_24578);
nor U25722 (N_25722,N_24736,N_24288);
xor U25723 (N_25723,N_22984,N_23229);
and U25724 (N_25724,N_22733,N_24996);
or U25725 (N_25725,N_22775,N_24204);
or U25726 (N_25726,N_22534,N_23539);
and U25727 (N_25727,N_23488,N_22850);
nor U25728 (N_25728,N_23460,N_24361);
xnor U25729 (N_25729,N_22511,N_23655);
or U25730 (N_25730,N_24600,N_24061);
xor U25731 (N_25731,N_24051,N_24631);
nand U25732 (N_25732,N_24059,N_23524);
or U25733 (N_25733,N_23719,N_23136);
xnor U25734 (N_25734,N_24671,N_22535);
or U25735 (N_25735,N_24281,N_22665);
and U25736 (N_25736,N_24660,N_22941);
xnor U25737 (N_25737,N_22987,N_24834);
and U25738 (N_25738,N_23505,N_23144);
or U25739 (N_25739,N_23437,N_23330);
nand U25740 (N_25740,N_24913,N_22702);
nor U25741 (N_25741,N_23003,N_24387);
and U25742 (N_25742,N_23141,N_22682);
and U25743 (N_25743,N_24603,N_24750);
nor U25744 (N_25744,N_24316,N_23349);
and U25745 (N_25745,N_23380,N_22618);
nor U25746 (N_25746,N_24510,N_23029);
nand U25747 (N_25747,N_24470,N_23423);
nand U25748 (N_25748,N_23068,N_24685);
xnor U25749 (N_25749,N_23767,N_22983);
or U25750 (N_25750,N_24336,N_22911);
or U25751 (N_25751,N_24096,N_23315);
and U25752 (N_25752,N_23151,N_24431);
nand U25753 (N_25753,N_24001,N_23065);
nand U25754 (N_25754,N_24956,N_24412);
nand U25755 (N_25755,N_23946,N_24348);
nand U25756 (N_25756,N_24192,N_24093);
or U25757 (N_25757,N_23545,N_23408);
and U25758 (N_25758,N_22988,N_23811);
nor U25759 (N_25759,N_22840,N_23731);
nor U25760 (N_25760,N_23074,N_24556);
or U25761 (N_25761,N_23027,N_24541);
or U25762 (N_25762,N_23283,N_23712);
xor U25763 (N_25763,N_23580,N_22630);
nor U25764 (N_25764,N_23156,N_23272);
and U25765 (N_25765,N_22847,N_24754);
and U25766 (N_25766,N_23352,N_22542);
or U25767 (N_25767,N_23361,N_23394);
nand U25768 (N_25768,N_23179,N_22706);
nor U25769 (N_25769,N_23605,N_23171);
nand U25770 (N_25770,N_23941,N_22860);
xor U25771 (N_25771,N_24429,N_23940);
and U25772 (N_25772,N_24203,N_23323);
xnor U25773 (N_25773,N_22530,N_22548);
or U25774 (N_25774,N_23570,N_24592);
and U25775 (N_25775,N_22869,N_24584);
or U25776 (N_25776,N_24159,N_23110);
or U25777 (N_25777,N_23255,N_23762);
nor U25778 (N_25778,N_24739,N_24318);
and U25779 (N_25779,N_23044,N_24305);
and U25780 (N_25780,N_24965,N_23132);
nand U25781 (N_25781,N_22816,N_23990);
nand U25782 (N_25782,N_24464,N_23763);
and U25783 (N_25783,N_24039,N_24268);
nor U25784 (N_25784,N_22781,N_24607);
and U25785 (N_25785,N_23411,N_24793);
nand U25786 (N_25786,N_23345,N_23788);
or U25787 (N_25787,N_24863,N_24790);
or U25788 (N_25788,N_23031,N_22982);
nand U25789 (N_25789,N_22874,N_24566);
xnor U25790 (N_25790,N_23328,N_23807);
xor U25791 (N_25791,N_24038,N_23013);
or U25792 (N_25792,N_23899,N_24306);
or U25793 (N_25793,N_23910,N_23943);
and U25794 (N_25794,N_22831,N_24565);
and U25795 (N_25795,N_24211,N_24903);
xor U25796 (N_25796,N_24536,N_24195);
and U25797 (N_25797,N_23251,N_24035);
xnor U25798 (N_25798,N_24786,N_23706);
nand U25799 (N_25799,N_23289,N_23754);
nor U25800 (N_25800,N_23076,N_24696);
or U25801 (N_25801,N_24391,N_24629);
nor U25802 (N_25802,N_24368,N_24787);
and U25803 (N_25803,N_24791,N_24557);
nand U25804 (N_25804,N_24886,N_24259);
and U25805 (N_25805,N_23228,N_24543);
and U25806 (N_25806,N_23197,N_23896);
xnor U25807 (N_25807,N_24855,N_23296);
or U25808 (N_25808,N_23106,N_22730);
xnor U25809 (N_25809,N_23665,N_23422);
xnor U25810 (N_25810,N_24349,N_23758);
or U25811 (N_25811,N_23249,N_24775);
nand U25812 (N_25812,N_24606,N_23070);
nand U25813 (N_25813,N_23523,N_22952);
nor U25814 (N_25814,N_23681,N_24110);
xnor U25815 (N_25815,N_24030,N_23043);
nor U25816 (N_25816,N_22806,N_24513);
and U25817 (N_25817,N_24928,N_22937);
nand U25818 (N_25818,N_24489,N_24706);
and U25819 (N_25819,N_22669,N_24982);
nor U25820 (N_25820,N_24022,N_24360);
or U25821 (N_25821,N_22699,N_24366);
nand U25822 (N_25822,N_22518,N_22895);
nor U25823 (N_25823,N_24962,N_24992);
and U25824 (N_25824,N_24465,N_23615);
nand U25825 (N_25825,N_22758,N_23353);
nand U25826 (N_25826,N_24969,N_23976);
xor U25827 (N_25827,N_22918,N_24976);
and U25828 (N_25828,N_24446,N_23809);
nand U25829 (N_25829,N_23983,N_22745);
and U25830 (N_25830,N_23335,N_22990);
and U25831 (N_25831,N_24588,N_22826);
or U25832 (N_25832,N_24709,N_23640);
and U25833 (N_25833,N_23541,N_23521);
xor U25834 (N_25834,N_23135,N_23098);
nand U25835 (N_25835,N_23111,N_24645);
or U25836 (N_25836,N_23701,N_22639);
nor U25837 (N_25837,N_24879,N_23778);
xor U25838 (N_25838,N_22623,N_24009);
and U25839 (N_25839,N_22572,N_23598);
or U25840 (N_25840,N_23148,N_24586);
nand U25841 (N_25841,N_22515,N_23490);
xor U25842 (N_25842,N_23838,N_22589);
and U25843 (N_25843,N_23988,N_24839);
or U25844 (N_25844,N_24756,N_23318);
nor U25845 (N_25845,N_24627,N_23644);
nand U25846 (N_25846,N_23936,N_24149);
and U25847 (N_25847,N_24715,N_23170);
or U25848 (N_25848,N_23400,N_24131);
and U25849 (N_25849,N_22755,N_23627);
nor U25850 (N_25850,N_23484,N_23025);
xor U25851 (N_25851,N_23882,N_23480);
xnor U25852 (N_25852,N_24394,N_22900);
nand U25853 (N_25853,N_23230,N_23212);
or U25854 (N_25854,N_22875,N_23969);
nand U25855 (N_25855,N_23826,N_24650);
and U25856 (N_25856,N_23909,N_23836);
nor U25857 (N_25857,N_24478,N_24342);
nor U25858 (N_25858,N_23014,N_22611);
or U25859 (N_25859,N_23485,N_23406);
or U25860 (N_25860,N_24860,N_23250);
nor U25861 (N_25861,N_24126,N_23476);
and U25862 (N_25862,N_22607,N_24239);
nor U25863 (N_25863,N_23978,N_23715);
xor U25864 (N_25864,N_23444,N_23635);
or U25865 (N_25865,N_23398,N_22710);
and U25866 (N_25866,N_23021,N_23686);
nand U25867 (N_25867,N_22593,N_23186);
or U25868 (N_25868,N_24459,N_22648);
nand U25869 (N_25869,N_24341,N_24469);
nand U25870 (N_25870,N_24544,N_23816);
and U25871 (N_25871,N_23218,N_23949);
xnor U25872 (N_25872,N_22613,N_24948);
xor U25873 (N_25873,N_24573,N_23300);
xor U25874 (N_25874,N_22635,N_23916);
xnor U25875 (N_25875,N_22714,N_24576);
nand U25876 (N_25876,N_24644,N_24526);
nor U25877 (N_25877,N_23236,N_24076);
xnor U25878 (N_25878,N_24052,N_23395);
nor U25879 (N_25879,N_23207,N_22544);
nor U25880 (N_25880,N_23579,N_24991);
or U25881 (N_25881,N_24742,N_23972);
xor U25882 (N_25882,N_24695,N_24745);
nand U25883 (N_25883,N_24136,N_23405);
nor U25884 (N_25884,N_24262,N_23696);
or U25885 (N_25885,N_23531,N_24702);
nand U25886 (N_25886,N_24411,N_22940);
xor U25887 (N_25887,N_22683,N_24002);
nand U25888 (N_25888,N_23948,N_24404);
nand U25889 (N_25889,N_22557,N_23358);
or U25890 (N_25890,N_22975,N_24236);
xor U25891 (N_25891,N_24924,N_22748);
nor U25892 (N_25892,N_24704,N_23256);
nor U25893 (N_25893,N_23239,N_24729);
and U25894 (N_25894,N_23188,N_23979);
nor U25895 (N_25895,N_24997,N_23075);
nand U25896 (N_25896,N_23839,N_24523);
and U25897 (N_25897,N_23241,N_23268);
nor U25898 (N_25898,N_22828,N_24048);
xnor U25899 (N_25899,N_24452,N_23861);
nor U25900 (N_25900,N_24272,N_24610);
nor U25901 (N_25901,N_24502,N_22931);
nand U25902 (N_25902,N_23832,N_23871);
xor U25903 (N_25903,N_23616,N_24765);
and U25904 (N_25904,N_22644,N_23536);
and U25905 (N_25905,N_24046,N_23479);
or U25906 (N_25906,N_22653,N_22802);
nand U25907 (N_25907,N_23270,N_23095);
or U25908 (N_25908,N_24384,N_24812);
nor U25909 (N_25909,N_24443,N_23276);
nor U25910 (N_25910,N_23953,N_22688);
and U25911 (N_25911,N_23769,N_24423);
and U25912 (N_25912,N_24932,N_24807);
nand U25913 (N_25913,N_23962,N_24878);
xor U25914 (N_25914,N_24155,N_22818);
xnor U25915 (N_25915,N_24738,N_24183);
nor U25916 (N_25916,N_24781,N_23876);
nor U25917 (N_25917,N_23552,N_24682);
or U25918 (N_25918,N_24861,N_24248);
xor U25919 (N_25919,N_24080,N_23089);
nor U25920 (N_25920,N_24437,N_24122);
and U25921 (N_25921,N_23295,N_22995);
nand U25922 (N_25922,N_24851,N_24647);
nor U25923 (N_25923,N_24590,N_24049);
or U25924 (N_25924,N_23430,N_23596);
nor U25925 (N_25925,N_24509,N_24219);
nor U25926 (N_25926,N_23244,N_24034);
nor U25927 (N_25927,N_23304,N_22992);
nor U25928 (N_25928,N_24554,N_23695);
xnor U25929 (N_25929,N_23660,N_23517);
nor U25930 (N_25930,N_22502,N_24938);
nor U25931 (N_25931,N_24889,N_23452);
or U25932 (N_25932,N_23814,N_22864);
nand U25933 (N_25933,N_22592,N_24279);
and U25934 (N_25934,N_24986,N_24538);
nor U25935 (N_25935,N_22837,N_24842);
nor U25936 (N_25936,N_23377,N_23852);
nor U25937 (N_25937,N_22953,N_24068);
nor U25938 (N_25938,N_24527,N_22827);
xor U25939 (N_25939,N_23412,N_24632);
xnor U25940 (N_25940,N_24210,N_24441);
and U25941 (N_25941,N_24593,N_24637);
and U25942 (N_25942,N_23284,N_24321);
nand U25943 (N_25943,N_22650,N_24708);
nand U25944 (N_25944,N_24354,N_23428);
and U25945 (N_25945,N_23124,N_23685);
and U25946 (N_25946,N_22841,N_24396);
xnor U25947 (N_25947,N_24092,N_23617);
and U25948 (N_25948,N_22658,N_22718);
nor U25949 (N_25949,N_24485,N_24925);
or U25950 (N_25950,N_23465,N_23786);
nor U25951 (N_25951,N_24911,N_24865);
xor U25952 (N_25952,N_23844,N_23680);
nand U25953 (N_25953,N_23977,N_22684);
nor U25954 (N_25954,N_23980,N_23091);
nor U25955 (N_25955,N_24549,N_23360);
nor U25956 (N_25956,N_24831,N_22964);
xor U25957 (N_25957,N_22724,N_22976);
nand U25958 (N_25958,N_23181,N_24293);
or U25959 (N_25959,N_24796,N_22709);
nand U25960 (N_25960,N_22876,N_24253);
nor U25961 (N_25961,N_22871,N_23820);
nor U25962 (N_25962,N_24247,N_23355);
or U25963 (N_25963,N_24662,N_23306);
nor U25964 (N_25964,N_24356,N_24338);
xnor U25965 (N_25965,N_22560,N_23726);
xnor U25966 (N_25966,N_24620,N_24233);
or U25967 (N_25967,N_23496,N_24298);
nand U25968 (N_25968,N_24435,N_23855);
and U25969 (N_25969,N_23475,N_24154);
or U25970 (N_25970,N_23000,N_24971);
nand U25971 (N_25971,N_24379,N_23421);
and U25972 (N_25972,N_22555,N_24289);
xor U25973 (N_25973,N_24174,N_24013);
nor U25974 (N_25974,N_24783,N_22522);
xor U25975 (N_25975,N_24546,N_23235);
or U25976 (N_25976,N_24599,N_24693);
nand U25977 (N_25977,N_22577,N_23527);
and U25978 (N_25978,N_24165,N_23237);
xnor U25979 (N_25979,N_22996,N_23331);
nand U25980 (N_25980,N_23209,N_22739);
nand U25981 (N_25981,N_23926,N_24649);
nand U25982 (N_25982,N_24065,N_24560);
nor U25983 (N_25983,N_22946,N_23467);
and U25984 (N_25984,N_23108,N_24472);
nand U25985 (N_25985,N_22596,N_22902);
and U25986 (N_25986,N_24830,N_24850);
and U25987 (N_25987,N_22851,N_24242);
and U25988 (N_25988,N_24295,N_24132);
nor U25989 (N_25989,N_23169,N_22713);
nor U25990 (N_25990,N_23491,N_23292);
or U25991 (N_25991,N_23772,N_24887);
nor U25992 (N_25992,N_22768,N_22993);
nor U25993 (N_25993,N_22803,N_24780);
xor U25994 (N_25994,N_24930,N_24852);
nor U25995 (N_25995,N_24207,N_24370);
nor U25996 (N_25996,N_23668,N_23952);
and U25997 (N_25997,N_24580,N_23364);
nand U25998 (N_25998,N_22579,N_23808);
and U25999 (N_25999,N_23482,N_24175);
or U26000 (N_26000,N_23628,N_24989);
or U26001 (N_26001,N_24615,N_24084);
or U26002 (N_26002,N_23698,N_24688);
xor U26003 (N_26003,N_22813,N_24254);
or U26004 (N_26004,N_24392,N_24893);
nor U26005 (N_26005,N_22677,N_22963);
and U26006 (N_26006,N_23611,N_23631);
and U26007 (N_26007,N_24810,N_22690);
nand U26008 (N_26008,N_24015,N_23441);
or U26009 (N_26009,N_23780,N_23601);
nand U26010 (N_26010,N_22793,N_22728);
or U26011 (N_26011,N_23257,N_24778);
xnor U26012 (N_26012,N_23034,N_23642);
nor U26013 (N_26013,N_23510,N_24945);
nand U26014 (N_26014,N_24492,N_22961);
nor U26015 (N_26015,N_22907,N_23713);
nor U26016 (N_26016,N_24955,N_22770);
nor U26017 (N_26017,N_23131,N_23945);
and U26018 (N_26018,N_23471,N_24981);
or U26019 (N_26019,N_23965,N_23560);
nand U26020 (N_26020,N_24574,N_24255);
xor U26021 (N_26021,N_22856,N_23022);
nand U26022 (N_26022,N_23260,N_23500);
nor U26023 (N_26023,N_24821,N_24221);
nand U26024 (N_26024,N_24891,N_23766);
nand U26025 (N_26025,N_22757,N_23993);
or U26026 (N_26026,N_24519,N_24866);
or U26027 (N_26027,N_24202,N_23796);
or U26028 (N_26028,N_24070,N_23610);
and U26029 (N_26029,N_24121,N_23783);
nand U26030 (N_26030,N_24535,N_24555);
or U26031 (N_26031,N_24872,N_23532);
xnor U26032 (N_26032,N_23987,N_24869);
nand U26033 (N_26033,N_23470,N_23185);
or U26034 (N_26034,N_24694,N_22715);
xor U26035 (N_26035,N_22600,N_24562);
and U26036 (N_26036,N_22526,N_24689);
or U26037 (N_26037,N_22879,N_23418);
nand U26038 (N_26038,N_23659,N_24330);
xor U26039 (N_26039,N_23609,N_24719);
nand U26040 (N_26040,N_23938,N_23204);
xnor U26041 (N_26041,N_23942,N_22804);
or U26042 (N_26042,N_23326,N_23371);
nor U26043 (N_26043,N_23588,N_23674);
or U26044 (N_26044,N_23312,N_24653);
and U26045 (N_26045,N_23409,N_23466);
and U26046 (N_26046,N_24246,N_24193);
and U26047 (N_26047,N_23724,N_24686);
or U26048 (N_26048,N_23293,N_24764);
nand U26049 (N_26049,N_24609,N_23913);
xnor U26050 (N_26050,N_24060,N_23056);
xnor U26051 (N_26051,N_23964,N_24874);
xor U26052 (N_26052,N_22540,N_23416);
nor U26053 (N_26053,N_23971,N_22520);
nor U26054 (N_26054,N_24105,N_23752);
xnor U26055 (N_26055,N_23054,N_24884);
and U26056 (N_26056,N_23897,N_24249);
nor U26057 (N_26057,N_23105,N_24450);
xor U26058 (N_26058,N_22839,N_24731);
nor U26059 (N_26059,N_23746,N_23639);
nor U26060 (N_26060,N_24483,N_24665);
xor U26061 (N_26061,N_22767,N_24197);
and U26062 (N_26062,N_23267,N_22967);
or U26063 (N_26063,N_24317,N_24160);
nor U26064 (N_26064,N_24815,N_23923);
xnor U26065 (N_26065,N_24343,N_23881);
xnor U26066 (N_26066,N_23550,N_24322);
and U26067 (N_26067,N_24382,N_23675);
xor U26068 (N_26068,N_23501,N_24113);
and U26069 (N_26069,N_22586,N_24115);
or U26070 (N_26070,N_22801,N_23206);
or U26071 (N_26071,N_23309,N_24161);
or U26072 (N_26072,N_22872,N_22603);
nand U26073 (N_26073,N_23950,N_24789);
or U26074 (N_26074,N_23765,N_23922);
or U26075 (N_26075,N_24934,N_24226);
nand U26076 (N_26076,N_24871,N_23522);
nor U26077 (N_26077,N_23734,N_24752);
and U26078 (N_26078,N_23998,N_24363);
xor U26079 (N_26079,N_22936,N_23770);
or U26080 (N_26080,N_23166,N_24383);
nand U26081 (N_26081,N_24419,N_23507);
or U26082 (N_26082,N_24156,N_22717);
xor U26083 (N_26083,N_23561,N_24743);
nand U26084 (N_26084,N_23087,N_23189);
and U26085 (N_26085,N_22716,N_24201);
nor U26086 (N_26086,N_22877,N_23840);
and U26087 (N_26087,N_24332,N_22703);
xnor U26088 (N_26088,N_22662,N_24770);
nor U26089 (N_26089,N_23242,N_24409);
nor U26090 (N_26090,N_23856,N_24194);
xnor U26091 (N_26091,N_23843,N_24278);
or U26092 (N_26092,N_24232,N_24998);
nand U26093 (N_26093,N_22968,N_24285);
nand U26094 (N_26094,N_24436,N_24675);
xnor U26095 (N_26095,N_22615,N_23944);
xor U26096 (N_26096,N_24008,N_24062);
or U26097 (N_26097,N_23001,N_24817);
nand U26098 (N_26098,N_24835,N_24146);
xnor U26099 (N_26099,N_22545,N_24144);
nor U26100 (N_26100,N_23959,N_23697);
xnor U26101 (N_26101,N_23035,N_23989);
or U26102 (N_26102,N_23049,N_24680);
xor U26103 (N_26103,N_23757,N_24488);
or U26104 (N_26104,N_23483,N_24237);
xnor U26105 (N_26105,N_23261,N_24941);
and U26106 (N_26106,N_23764,N_22670);
and U26107 (N_26107,N_23172,N_23589);
xor U26108 (N_26108,N_23351,N_24280);
nand U26109 (N_26109,N_24222,N_23120);
nand U26110 (N_26110,N_22881,N_23407);
xor U26111 (N_26111,N_23534,N_23622);
or U26112 (N_26112,N_24054,N_24958);
or U26113 (N_26113,N_23996,N_23586);
nor U26114 (N_26114,N_23417,N_24018);
nand U26115 (N_26115,N_24625,N_23354);
and U26116 (N_26116,N_24244,N_22519);
xnor U26117 (N_26117,N_23833,N_24612);
xor U26118 (N_26118,N_23234,N_23747);
xor U26119 (N_26119,N_24339,N_24448);
or U26120 (N_26120,N_23663,N_23393);
nor U26121 (N_26121,N_24218,N_23920);
or U26122 (N_26122,N_24301,N_24381);
nor U26123 (N_26123,N_24228,N_23083);
nor U26124 (N_26124,N_23090,N_22950);
nand U26125 (N_26125,N_24087,N_22525);
xor U26126 (N_26126,N_24563,N_24234);
nand U26127 (N_26127,N_24359,N_24346);
nand U26128 (N_26128,N_23404,N_24173);
nor U26129 (N_26129,N_23338,N_23868);
or U26130 (N_26130,N_23568,N_23889);
xnor U26131 (N_26131,N_23410,N_23440);
xor U26132 (N_26132,N_24897,N_23658);
xor U26133 (N_26133,N_22880,N_24993);
nor U26134 (N_26134,N_23363,N_23776);
and U26135 (N_26135,N_24312,N_24701);
or U26136 (N_26136,N_24311,N_24726);
or U26137 (N_26137,N_24212,N_22928);
nand U26138 (N_26138,N_22986,N_23782);
and U26139 (N_26139,N_24548,N_23319);
or U26140 (N_26140,N_24529,N_24040);
and U26141 (N_26141,N_23216,N_24447);
xnor U26142 (N_26142,N_22747,N_23915);
xnor U26143 (N_26143,N_22822,N_24868);
or U26144 (N_26144,N_23650,N_24011);
or U26145 (N_26145,N_22915,N_24819);
nand U26146 (N_26146,N_23963,N_24078);
or U26147 (N_26147,N_23710,N_22883);
and U26148 (N_26148,N_24235,N_23537);
nor U26149 (N_26149,N_22836,N_22510);
and U26150 (N_26150,N_23258,N_23058);
and U26151 (N_26151,N_23932,N_24164);
or U26152 (N_26152,N_24515,N_23498);
or U26153 (N_26153,N_24724,N_22892);
nor U26154 (N_26154,N_23175,N_23775);
nand U26155 (N_26155,N_23381,N_22571);
nor U26156 (N_26156,N_24766,N_24077);
and U26157 (N_26157,N_24699,N_24257);
and U26158 (N_26158,N_23509,N_23497);
or U26159 (N_26159,N_24216,N_22981);
nor U26160 (N_26160,N_22752,N_24988);
xor U26161 (N_26161,N_22612,N_24762);
nand U26162 (N_26162,N_23666,N_23357);
or U26163 (N_26163,N_24797,N_22820);
and U26164 (N_26164,N_23894,N_23704);
and U26165 (N_26165,N_24664,N_24480);
or U26166 (N_26166,N_23177,N_24511);
nand U26167 (N_26167,N_24352,N_23403);
nand U26168 (N_26168,N_23269,N_23205);
or U26169 (N_26169,N_24010,N_23961);
or U26170 (N_26170,N_24421,N_22509);
nor U26171 (N_26171,N_22914,N_23174);
xor U26172 (N_26172,N_24400,N_22916);
or U26173 (N_26173,N_23473,N_24109);
and U26174 (N_26174,N_23324,N_24328);
nor U26175 (N_26175,N_24189,N_22622);
and U26176 (N_26176,N_22909,N_23041);
or U26177 (N_26177,N_23718,N_22947);
and U26178 (N_26178,N_24353,N_22980);
and U26179 (N_26179,N_23246,N_24395);
and U26180 (N_26180,N_24944,N_23130);
xor U26181 (N_26181,N_24822,N_23929);
xnor U26182 (N_26182,N_22517,N_23702);
xor U26183 (N_26183,N_22624,N_22808);
or U26184 (N_26184,N_22539,N_22731);
nand U26185 (N_26185,N_24145,N_23999);
and U26186 (N_26186,N_24522,N_24264);
nand U26187 (N_26187,N_24307,N_24141);
and U26188 (N_26188,N_23053,N_23578);
and U26189 (N_26189,N_23427,N_22536);
and U26190 (N_26190,N_23387,N_22750);
and U26191 (N_26191,N_24581,N_24344);
nand U26192 (N_26192,N_22762,N_24128);
or U26193 (N_26193,N_24112,N_22904);
nand U26194 (N_26194,N_23340,N_23116);
or U26195 (N_26195,N_24961,N_24970);
or U26196 (N_26196,N_24004,N_24269);
xnor U26197 (N_26197,N_22805,N_22799);
xor U26198 (N_26198,N_22707,N_22538);
or U26199 (N_26199,N_23114,N_22629);
nor U26200 (N_26200,N_24416,N_22741);
and U26201 (N_26201,N_24676,N_22564);
nor U26202 (N_26202,N_23662,N_24275);
or U26203 (N_26203,N_24572,N_23051);
and U26204 (N_26204,N_22661,N_24088);
nand U26205 (N_26205,N_24405,N_23322);
nand U26206 (N_26206,N_22785,N_23356);
nor U26207 (N_26207,N_24125,N_23608);
xnor U26208 (N_26208,N_22821,N_23636);
nand U26209 (N_26209,N_23682,N_23303);
nand U26210 (N_26210,N_22686,N_22666);
nor U26211 (N_26211,N_22886,N_24547);
xnor U26212 (N_26212,N_23248,N_24614);
or U26213 (N_26213,N_23481,N_23597);
nand U26214 (N_26214,N_24668,N_23583);
or U26215 (N_26215,N_23092,N_24508);
and U26216 (N_26216,N_24963,N_23721);
nor U26217 (N_26217,N_24840,N_22640);
or U26218 (N_26218,N_22908,N_23321);
or U26219 (N_26219,N_24847,N_22974);
nand U26220 (N_26220,N_24518,N_23194);
or U26221 (N_26221,N_23912,N_23225);
nor U26222 (N_26222,N_23634,N_23266);
nand U26223 (N_26223,N_22601,N_24284);
xnor U26224 (N_26224,N_22924,N_24283);
nor U26225 (N_26225,N_23337,N_23050);
or U26226 (N_26226,N_24428,N_24977);
and U26227 (N_26227,N_24907,N_23487);
xnor U26228 (N_26228,N_23127,N_22815);
nand U26229 (N_26229,N_23341,N_24853);
nor U26230 (N_26230,N_23344,N_23192);
nor U26231 (N_26231,N_22637,N_24310);
xor U26232 (N_26232,N_22567,N_24016);
xnor U26233 (N_26233,N_24744,N_24276);
nand U26234 (N_26234,N_24862,N_24320);
xor U26235 (N_26235,N_23157,N_24910);
nand U26236 (N_26236,N_22727,N_23011);
nand U26237 (N_26237,N_22965,N_23140);
nand U26238 (N_26238,N_24846,N_24875);
nor U26239 (N_26239,N_22736,N_24735);
and U26240 (N_26240,N_24449,N_24225);
nand U26241 (N_26241,N_24525,N_23960);
xor U26242 (N_26242,N_24959,N_24215);
or U26243 (N_26243,N_22783,N_24493);
or U26244 (N_26244,N_23893,N_23994);
or U26245 (N_26245,N_22922,N_24319);
nand U26246 (N_26246,N_22738,N_24950);
nand U26247 (N_26247,N_24467,N_23917);
or U26248 (N_26248,N_24995,N_24028);
and U26249 (N_26249,N_23314,N_24800);
nand U26250 (N_26250,N_23880,N_22654);
nand U26251 (N_26251,N_24975,N_24148);
and U26252 (N_26252,N_22844,N_24628);
xnor U26253 (N_26253,N_24393,N_23944);
and U26254 (N_26254,N_22662,N_23258);
and U26255 (N_26255,N_23429,N_22723);
nor U26256 (N_26256,N_23975,N_22866);
and U26257 (N_26257,N_23483,N_23922);
or U26258 (N_26258,N_23530,N_24129);
and U26259 (N_26259,N_24575,N_24950);
or U26260 (N_26260,N_23693,N_24972);
nor U26261 (N_26261,N_22504,N_24329);
and U26262 (N_26262,N_23854,N_23596);
xnor U26263 (N_26263,N_24737,N_23075);
nor U26264 (N_26264,N_23719,N_24531);
xnor U26265 (N_26265,N_23319,N_23524);
xor U26266 (N_26266,N_24242,N_22680);
and U26267 (N_26267,N_23383,N_23666);
and U26268 (N_26268,N_24855,N_22508);
nor U26269 (N_26269,N_24785,N_23505);
nand U26270 (N_26270,N_23762,N_24021);
and U26271 (N_26271,N_24109,N_23884);
or U26272 (N_26272,N_23953,N_24079);
nor U26273 (N_26273,N_22952,N_23008);
and U26274 (N_26274,N_24964,N_24368);
nand U26275 (N_26275,N_22501,N_23275);
nand U26276 (N_26276,N_23482,N_24357);
nand U26277 (N_26277,N_23515,N_23428);
or U26278 (N_26278,N_24266,N_24456);
or U26279 (N_26279,N_22500,N_23575);
and U26280 (N_26280,N_24551,N_23997);
or U26281 (N_26281,N_23526,N_24258);
xnor U26282 (N_26282,N_24259,N_24871);
and U26283 (N_26283,N_23510,N_23005);
nor U26284 (N_26284,N_24129,N_23897);
or U26285 (N_26285,N_24720,N_22643);
nand U26286 (N_26286,N_23075,N_24075);
nor U26287 (N_26287,N_24788,N_22725);
xor U26288 (N_26288,N_22990,N_23522);
xnor U26289 (N_26289,N_23120,N_22724);
and U26290 (N_26290,N_24761,N_24791);
nor U26291 (N_26291,N_22777,N_24727);
and U26292 (N_26292,N_23125,N_22762);
or U26293 (N_26293,N_24734,N_24365);
and U26294 (N_26294,N_23445,N_24791);
nand U26295 (N_26295,N_23581,N_24548);
nor U26296 (N_26296,N_24453,N_23596);
nand U26297 (N_26297,N_24149,N_24965);
xnor U26298 (N_26298,N_24286,N_23557);
or U26299 (N_26299,N_23567,N_23606);
nor U26300 (N_26300,N_24398,N_23005);
nand U26301 (N_26301,N_23909,N_23953);
xnor U26302 (N_26302,N_23676,N_24897);
xor U26303 (N_26303,N_22626,N_23059);
and U26304 (N_26304,N_24620,N_22738);
nor U26305 (N_26305,N_23040,N_23479);
and U26306 (N_26306,N_24545,N_24338);
xnor U26307 (N_26307,N_24152,N_22789);
or U26308 (N_26308,N_22672,N_24127);
or U26309 (N_26309,N_24450,N_24052);
nor U26310 (N_26310,N_24913,N_24401);
nor U26311 (N_26311,N_24410,N_24343);
xnor U26312 (N_26312,N_23028,N_24180);
nand U26313 (N_26313,N_23417,N_24539);
nand U26314 (N_26314,N_24814,N_24193);
and U26315 (N_26315,N_24202,N_24639);
xnor U26316 (N_26316,N_24374,N_23237);
nor U26317 (N_26317,N_22541,N_23186);
nand U26318 (N_26318,N_23934,N_24080);
nor U26319 (N_26319,N_23931,N_24646);
nand U26320 (N_26320,N_23504,N_23124);
xnor U26321 (N_26321,N_24815,N_24674);
nand U26322 (N_26322,N_24915,N_23569);
xor U26323 (N_26323,N_23853,N_22834);
nor U26324 (N_26324,N_22510,N_23785);
or U26325 (N_26325,N_24944,N_23623);
xnor U26326 (N_26326,N_23382,N_22611);
or U26327 (N_26327,N_23818,N_23699);
xor U26328 (N_26328,N_23611,N_24815);
or U26329 (N_26329,N_23203,N_23692);
nand U26330 (N_26330,N_23065,N_24105);
nand U26331 (N_26331,N_23229,N_23596);
xnor U26332 (N_26332,N_24153,N_23359);
xnor U26333 (N_26333,N_24016,N_24786);
nor U26334 (N_26334,N_22966,N_24265);
xor U26335 (N_26335,N_23404,N_23509);
nor U26336 (N_26336,N_24384,N_22579);
nor U26337 (N_26337,N_22580,N_22719);
and U26338 (N_26338,N_23699,N_22962);
nor U26339 (N_26339,N_24516,N_23249);
nor U26340 (N_26340,N_24536,N_23609);
xnor U26341 (N_26341,N_24547,N_23858);
xor U26342 (N_26342,N_24288,N_24520);
and U26343 (N_26343,N_23000,N_23676);
and U26344 (N_26344,N_23627,N_23909);
nor U26345 (N_26345,N_24845,N_24458);
or U26346 (N_26346,N_23116,N_23660);
and U26347 (N_26347,N_23167,N_22819);
nand U26348 (N_26348,N_23682,N_24249);
nor U26349 (N_26349,N_23174,N_24147);
nand U26350 (N_26350,N_23822,N_22977);
nand U26351 (N_26351,N_24163,N_24362);
xor U26352 (N_26352,N_22599,N_22741);
and U26353 (N_26353,N_22930,N_24846);
xor U26354 (N_26354,N_22525,N_24325);
nor U26355 (N_26355,N_24968,N_24033);
xnor U26356 (N_26356,N_22871,N_23631);
or U26357 (N_26357,N_23623,N_24166);
nand U26358 (N_26358,N_23126,N_23603);
xor U26359 (N_26359,N_23352,N_23343);
or U26360 (N_26360,N_24246,N_23411);
or U26361 (N_26361,N_22864,N_23815);
and U26362 (N_26362,N_23002,N_22999);
or U26363 (N_26363,N_23288,N_23133);
nand U26364 (N_26364,N_24245,N_24586);
xnor U26365 (N_26365,N_24303,N_22786);
nand U26366 (N_26366,N_23162,N_23624);
nand U26367 (N_26367,N_23422,N_22594);
and U26368 (N_26368,N_23655,N_23054);
nor U26369 (N_26369,N_22770,N_23739);
or U26370 (N_26370,N_24134,N_24098);
and U26371 (N_26371,N_24496,N_24656);
nor U26372 (N_26372,N_24490,N_24841);
or U26373 (N_26373,N_24445,N_22999);
nor U26374 (N_26374,N_23231,N_24070);
nand U26375 (N_26375,N_22539,N_24209);
xnor U26376 (N_26376,N_22911,N_24866);
nor U26377 (N_26377,N_24550,N_23974);
xnor U26378 (N_26378,N_23626,N_22730);
nor U26379 (N_26379,N_23100,N_24519);
nand U26380 (N_26380,N_23665,N_24908);
and U26381 (N_26381,N_23410,N_23992);
nand U26382 (N_26382,N_23388,N_22677);
nor U26383 (N_26383,N_23160,N_23040);
and U26384 (N_26384,N_23706,N_23096);
and U26385 (N_26385,N_24079,N_23440);
and U26386 (N_26386,N_24425,N_23151);
or U26387 (N_26387,N_23639,N_24624);
nand U26388 (N_26388,N_23698,N_24064);
and U26389 (N_26389,N_22572,N_23753);
nor U26390 (N_26390,N_22538,N_23276);
nor U26391 (N_26391,N_24578,N_24974);
nor U26392 (N_26392,N_22816,N_22713);
nor U26393 (N_26393,N_24320,N_24148);
nor U26394 (N_26394,N_22504,N_24421);
or U26395 (N_26395,N_22806,N_24240);
and U26396 (N_26396,N_23010,N_23264);
nand U26397 (N_26397,N_24888,N_24525);
nor U26398 (N_26398,N_23950,N_24097);
xnor U26399 (N_26399,N_22989,N_22563);
nor U26400 (N_26400,N_23645,N_23850);
xnor U26401 (N_26401,N_24098,N_23750);
nor U26402 (N_26402,N_24937,N_24434);
xor U26403 (N_26403,N_23069,N_24727);
and U26404 (N_26404,N_22996,N_23093);
or U26405 (N_26405,N_24212,N_23305);
nand U26406 (N_26406,N_23478,N_23887);
or U26407 (N_26407,N_23535,N_23851);
nand U26408 (N_26408,N_23001,N_24081);
and U26409 (N_26409,N_23000,N_23576);
or U26410 (N_26410,N_23126,N_24742);
and U26411 (N_26411,N_23273,N_22708);
nand U26412 (N_26412,N_24350,N_23171);
and U26413 (N_26413,N_24711,N_23195);
nand U26414 (N_26414,N_24312,N_24669);
nor U26415 (N_26415,N_23398,N_22850);
nand U26416 (N_26416,N_22947,N_24545);
and U26417 (N_26417,N_24000,N_22684);
nand U26418 (N_26418,N_23678,N_22693);
or U26419 (N_26419,N_24005,N_22795);
nor U26420 (N_26420,N_22509,N_22793);
or U26421 (N_26421,N_22675,N_22715);
nand U26422 (N_26422,N_23836,N_23689);
or U26423 (N_26423,N_22522,N_22844);
nor U26424 (N_26424,N_24770,N_22709);
nand U26425 (N_26425,N_23015,N_23800);
nor U26426 (N_26426,N_23588,N_23397);
xnor U26427 (N_26427,N_23203,N_24049);
xor U26428 (N_26428,N_24115,N_22842);
or U26429 (N_26429,N_22776,N_24141);
or U26430 (N_26430,N_24692,N_22571);
nand U26431 (N_26431,N_22545,N_24789);
xnor U26432 (N_26432,N_24286,N_24466);
xor U26433 (N_26433,N_23295,N_24967);
xnor U26434 (N_26434,N_24457,N_23105);
nand U26435 (N_26435,N_23128,N_22922);
nor U26436 (N_26436,N_22732,N_23756);
or U26437 (N_26437,N_24280,N_22998);
nor U26438 (N_26438,N_24485,N_24738);
nor U26439 (N_26439,N_24405,N_24019);
and U26440 (N_26440,N_23882,N_23266);
and U26441 (N_26441,N_23316,N_23580);
or U26442 (N_26442,N_24611,N_24365);
nor U26443 (N_26443,N_23316,N_24956);
or U26444 (N_26444,N_24506,N_24595);
and U26445 (N_26445,N_24878,N_22753);
or U26446 (N_26446,N_22970,N_24298);
or U26447 (N_26447,N_23268,N_23670);
xor U26448 (N_26448,N_24561,N_24797);
and U26449 (N_26449,N_24227,N_22549);
xor U26450 (N_26450,N_22543,N_24806);
nand U26451 (N_26451,N_24213,N_23483);
or U26452 (N_26452,N_23491,N_23012);
nand U26453 (N_26453,N_22688,N_24474);
xnor U26454 (N_26454,N_22822,N_24728);
nor U26455 (N_26455,N_24358,N_22728);
xor U26456 (N_26456,N_23616,N_23913);
nand U26457 (N_26457,N_24535,N_24931);
nor U26458 (N_26458,N_24762,N_23358);
xor U26459 (N_26459,N_22913,N_22506);
nand U26460 (N_26460,N_23089,N_22828);
and U26461 (N_26461,N_22540,N_23628);
xnor U26462 (N_26462,N_24902,N_23605);
nand U26463 (N_26463,N_24762,N_24972);
nand U26464 (N_26464,N_23273,N_23583);
nand U26465 (N_26465,N_24777,N_23341);
or U26466 (N_26466,N_23092,N_22637);
xnor U26467 (N_26467,N_24988,N_22922);
xor U26468 (N_26468,N_24889,N_22501);
nand U26469 (N_26469,N_24671,N_24716);
or U26470 (N_26470,N_24589,N_23571);
and U26471 (N_26471,N_23391,N_22835);
and U26472 (N_26472,N_22542,N_22863);
nor U26473 (N_26473,N_22892,N_22866);
or U26474 (N_26474,N_24146,N_22941);
nor U26475 (N_26475,N_23543,N_23800);
xnor U26476 (N_26476,N_24685,N_22680);
xnor U26477 (N_26477,N_24852,N_23211);
and U26478 (N_26478,N_22681,N_22635);
or U26479 (N_26479,N_23752,N_23597);
nand U26480 (N_26480,N_24926,N_24991);
xor U26481 (N_26481,N_22978,N_23300);
or U26482 (N_26482,N_24644,N_24339);
and U26483 (N_26483,N_24368,N_24839);
or U26484 (N_26484,N_24313,N_22917);
or U26485 (N_26485,N_22815,N_24407);
nor U26486 (N_26486,N_24062,N_23419);
xor U26487 (N_26487,N_24684,N_24010);
nor U26488 (N_26488,N_23944,N_24766);
or U26489 (N_26489,N_24055,N_23492);
nor U26490 (N_26490,N_24212,N_24296);
nor U26491 (N_26491,N_22896,N_23277);
or U26492 (N_26492,N_23345,N_23000);
and U26493 (N_26493,N_23674,N_22726);
and U26494 (N_26494,N_24895,N_22929);
xor U26495 (N_26495,N_23726,N_22806);
or U26496 (N_26496,N_23014,N_23440);
nand U26497 (N_26497,N_22533,N_23367);
or U26498 (N_26498,N_23865,N_22622);
nand U26499 (N_26499,N_24601,N_24851);
nor U26500 (N_26500,N_24108,N_24472);
or U26501 (N_26501,N_23207,N_23735);
xor U26502 (N_26502,N_24004,N_22622);
nand U26503 (N_26503,N_23362,N_24642);
or U26504 (N_26504,N_23557,N_23967);
and U26505 (N_26505,N_23206,N_23766);
nand U26506 (N_26506,N_24448,N_22931);
nor U26507 (N_26507,N_23806,N_23088);
nand U26508 (N_26508,N_24449,N_24195);
or U26509 (N_26509,N_24136,N_24374);
nand U26510 (N_26510,N_24157,N_23800);
and U26511 (N_26511,N_22617,N_24339);
or U26512 (N_26512,N_24341,N_22834);
and U26513 (N_26513,N_23184,N_23293);
nor U26514 (N_26514,N_24155,N_23167);
or U26515 (N_26515,N_24263,N_23949);
and U26516 (N_26516,N_24502,N_24012);
and U26517 (N_26517,N_23985,N_24204);
nand U26518 (N_26518,N_22955,N_23594);
and U26519 (N_26519,N_23022,N_24944);
nor U26520 (N_26520,N_22988,N_23722);
nand U26521 (N_26521,N_23828,N_23243);
nor U26522 (N_26522,N_23385,N_22548);
xnor U26523 (N_26523,N_24119,N_23778);
or U26524 (N_26524,N_23383,N_23795);
and U26525 (N_26525,N_22804,N_24528);
nand U26526 (N_26526,N_24263,N_24423);
or U26527 (N_26527,N_22645,N_23473);
or U26528 (N_26528,N_23556,N_24342);
or U26529 (N_26529,N_23002,N_23179);
xnor U26530 (N_26530,N_24372,N_24792);
nand U26531 (N_26531,N_23913,N_23033);
or U26532 (N_26532,N_23241,N_23538);
nor U26533 (N_26533,N_24383,N_24376);
or U26534 (N_26534,N_24792,N_24654);
or U26535 (N_26535,N_24448,N_23040);
or U26536 (N_26536,N_23031,N_23936);
xor U26537 (N_26537,N_24406,N_24342);
or U26538 (N_26538,N_23188,N_23805);
or U26539 (N_26539,N_24041,N_23326);
nor U26540 (N_26540,N_24662,N_22847);
xor U26541 (N_26541,N_22533,N_23552);
nor U26542 (N_26542,N_22863,N_24949);
and U26543 (N_26543,N_23753,N_22868);
and U26544 (N_26544,N_24361,N_24658);
and U26545 (N_26545,N_24118,N_24632);
and U26546 (N_26546,N_22662,N_22522);
nor U26547 (N_26547,N_22506,N_24758);
nand U26548 (N_26548,N_23374,N_23852);
or U26549 (N_26549,N_24598,N_23504);
nand U26550 (N_26550,N_24134,N_23707);
nor U26551 (N_26551,N_22633,N_24459);
nor U26552 (N_26552,N_23787,N_23549);
or U26553 (N_26553,N_23677,N_23993);
and U26554 (N_26554,N_23894,N_24892);
and U26555 (N_26555,N_24715,N_23549);
nand U26556 (N_26556,N_24132,N_23192);
xor U26557 (N_26557,N_23695,N_23633);
xor U26558 (N_26558,N_22983,N_22621);
or U26559 (N_26559,N_24775,N_22688);
or U26560 (N_26560,N_24129,N_22964);
xor U26561 (N_26561,N_24167,N_24666);
or U26562 (N_26562,N_24075,N_24289);
or U26563 (N_26563,N_23481,N_23031);
and U26564 (N_26564,N_24567,N_22843);
or U26565 (N_26565,N_24803,N_22950);
xor U26566 (N_26566,N_23268,N_23563);
or U26567 (N_26567,N_24620,N_22583);
nand U26568 (N_26568,N_23141,N_23276);
and U26569 (N_26569,N_23628,N_23332);
nor U26570 (N_26570,N_24329,N_24312);
and U26571 (N_26571,N_23540,N_23880);
xnor U26572 (N_26572,N_23809,N_22911);
nor U26573 (N_26573,N_23114,N_22628);
nand U26574 (N_26574,N_23137,N_22536);
nor U26575 (N_26575,N_24423,N_23803);
and U26576 (N_26576,N_23803,N_23582);
and U26577 (N_26577,N_24052,N_24411);
nor U26578 (N_26578,N_23807,N_23636);
nor U26579 (N_26579,N_22883,N_24524);
nor U26580 (N_26580,N_24087,N_23671);
nor U26581 (N_26581,N_24844,N_24711);
nor U26582 (N_26582,N_23378,N_24749);
and U26583 (N_26583,N_23820,N_23147);
nor U26584 (N_26584,N_24684,N_24133);
xor U26585 (N_26585,N_23178,N_24414);
nor U26586 (N_26586,N_23634,N_22920);
or U26587 (N_26587,N_24262,N_24708);
or U26588 (N_26588,N_24701,N_24352);
xnor U26589 (N_26589,N_24184,N_22639);
or U26590 (N_26590,N_23892,N_23256);
xnor U26591 (N_26591,N_23183,N_24269);
nand U26592 (N_26592,N_24905,N_22729);
nand U26593 (N_26593,N_22920,N_24498);
and U26594 (N_26594,N_24605,N_24957);
nor U26595 (N_26595,N_24810,N_23465);
nand U26596 (N_26596,N_23725,N_23226);
and U26597 (N_26597,N_24331,N_24599);
nor U26598 (N_26598,N_23301,N_24313);
or U26599 (N_26599,N_23281,N_23244);
or U26600 (N_26600,N_23229,N_23754);
and U26601 (N_26601,N_24749,N_24611);
nand U26602 (N_26602,N_24609,N_24584);
nor U26603 (N_26603,N_23715,N_23194);
nor U26604 (N_26604,N_23504,N_24833);
and U26605 (N_26605,N_24575,N_23453);
or U26606 (N_26606,N_23211,N_22752);
nand U26607 (N_26607,N_23147,N_23727);
and U26608 (N_26608,N_24996,N_23262);
xor U26609 (N_26609,N_24022,N_23136);
or U26610 (N_26610,N_22920,N_23894);
and U26611 (N_26611,N_24936,N_24066);
nand U26612 (N_26612,N_22684,N_24835);
or U26613 (N_26613,N_24221,N_24282);
nand U26614 (N_26614,N_23172,N_24919);
or U26615 (N_26615,N_22886,N_24641);
nor U26616 (N_26616,N_22795,N_24795);
and U26617 (N_26617,N_23427,N_24930);
nand U26618 (N_26618,N_24389,N_24502);
nand U26619 (N_26619,N_23343,N_24377);
or U26620 (N_26620,N_22648,N_22617);
and U26621 (N_26621,N_23506,N_24017);
or U26622 (N_26622,N_24690,N_24830);
nor U26623 (N_26623,N_22555,N_23992);
and U26624 (N_26624,N_24277,N_23512);
nor U26625 (N_26625,N_23633,N_24321);
xnor U26626 (N_26626,N_23613,N_22720);
or U26627 (N_26627,N_23539,N_24131);
nor U26628 (N_26628,N_24871,N_22529);
and U26629 (N_26629,N_23775,N_23616);
nand U26630 (N_26630,N_24707,N_24311);
nor U26631 (N_26631,N_24591,N_23099);
and U26632 (N_26632,N_22889,N_23489);
xnor U26633 (N_26633,N_24950,N_23957);
nor U26634 (N_26634,N_24614,N_24152);
and U26635 (N_26635,N_24383,N_23904);
xnor U26636 (N_26636,N_22518,N_22568);
nor U26637 (N_26637,N_23332,N_24125);
xnor U26638 (N_26638,N_23103,N_22985);
xnor U26639 (N_26639,N_22987,N_22893);
nor U26640 (N_26640,N_23199,N_24881);
or U26641 (N_26641,N_24587,N_24302);
xnor U26642 (N_26642,N_23054,N_23366);
nor U26643 (N_26643,N_23229,N_23026);
xnor U26644 (N_26644,N_24218,N_23423);
and U26645 (N_26645,N_23239,N_23751);
nand U26646 (N_26646,N_23624,N_24988);
nand U26647 (N_26647,N_22897,N_23440);
nor U26648 (N_26648,N_23997,N_23117);
and U26649 (N_26649,N_24794,N_23144);
xor U26650 (N_26650,N_24443,N_23287);
nand U26651 (N_26651,N_22771,N_24477);
nor U26652 (N_26652,N_22949,N_22602);
and U26653 (N_26653,N_23132,N_24466);
or U26654 (N_26654,N_24298,N_24117);
nand U26655 (N_26655,N_23436,N_23250);
xnor U26656 (N_26656,N_23116,N_23589);
nand U26657 (N_26657,N_23942,N_22708);
nor U26658 (N_26658,N_23023,N_23415);
xnor U26659 (N_26659,N_24744,N_23631);
nand U26660 (N_26660,N_24148,N_23028);
nand U26661 (N_26661,N_23401,N_22658);
and U26662 (N_26662,N_24437,N_24416);
or U26663 (N_26663,N_23019,N_24905);
and U26664 (N_26664,N_23843,N_24565);
and U26665 (N_26665,N_23867,N_22906);
nand U26666 (N_26666,N_23999,N_24342);
or U26667 (N_26667,N_24031,N_24800);
and U26668 (N_26668,N_24069,N_24642);
nor U26669 (N_26669,N_23706,N_23936);
and U26670 (N_26670,N_23877,N_24359);
xnor U26671 (N_26671,N_24666,N_22791);
nor U26672 (N_26672,N_23399,N_24611);
nor U26673 (N_26673,N_22584,N_24403);
and U26674 (N_26674,N_23161,N_23979);
nand U26675 (N_26675,N_24198,N_23905);
nor U26676 (N_26676,N_24786,N_22822);
nor U26677 (N_26677,N_24930,N_23904);
nand U26678 (N_26678,N_23838,N_22661);
and U26679 (N_26679,N_24885,N_22591);
or U26680 (N_26680,N_22874,N_24767);
and U26681 (N_26681,N_23683,N_24913);
or U26682 (N_26682,N_22567,N_24315);
nor U26683 (N_26683,N_23621,N_24840);
and U26684 (N_26684,N_23684,N_22970);
or U26685 (N_26685,N_24638,N_23234);
or U26686 (N_26686,N_24108,N_24107);
nor U26687 (N_26687,N_22722,N_22882);
or U26688 (N_26688,N_23124,N_23417);
nor U26689 (N_26689,N_23871,N_23214);
and U26690 (N_26690,N_24764,N_24341);
nand U26691 (N_26691,N_24481,N_24287);
or U26692 (N_26692,N_24646,N_24343);
nand U26693 (N_26693,N_23032,N_23675);
nand U26694 (N_26694,N_23594,N_23042);
nand U26695 (N_26695,N_22641,N_24783);
xnor U26696 (N_26696,N_22514,N_24061);
nor U26697 (N_26697,N_23265,N_22662);
nand U26698 (N_26698,N_22594,N_23104);
or U26699 (N_26699,N_24280,N_24369);
xnor U26700 (N_26700,N_24287,N_23067);
nand U26701 (N_26701,N_23188,N_24177);
or U26702 (N_26702,N_23125,N_23962);
nand U26703 (N_26703,N_24520,N_24786);
nor U26704 (N_26704,N_23016,N_24291);
xnor U26705 (N_26705,N_23692,N_23885);
xnor U26706 (N_26706,N_24880,N_24617);
nand U26707 (N_26707,N_23839,N_23897);
xor U26708 (N_26708,N_23587,N_23398);
and U26709 (N_26709,N_24724,N_23462);
or U26710 (N_26710,N_22750,N_22769);
xor U26711 (N_26711,N_22972,N_22886);
and U26712 (N_26712,N_24383,N_22959);
nand U26713 (N_26713,N_24669,N_22999);
and U26714 (N_26714,N_24789,N_23497);
nand U26715 (N_26715,N_24215,N_22791);
and U26716 (N_26716,N_24009,N_23749);
nor U26717 (N_26717,N_22974,N_22928);
nand U26718 (N_26718,N_23774,N_24422);
nor U26719 (N_26719,N_22762,N_24305);
nand U26720 (N_26720,N_24191,N_23830);
xor U26721 (N_26721,N_24439,N_23796);
xnor U26722 (N_26722,N_23428,N_23102);
xor U26723 (N_26723,N_23219,N_22812);
xor U26724 (N_26724,N_24060,N_24214);
xor U26725 (N_26725,N_24623,N_23958);
and U26726 (N_26726,N_22837,N_24217);
nor U26727 (N_26727,N_23977,N_23398);
and U26728 (N_26728,N_24613,N_22718);
nand U26729 (N_26729,N_23834,N_23804);
xor U26730 (N_26730,N_24968,N_22982);
nand U26731 (N_26731,N_22861,N_23836);
and U26732 (N_26732,N_22938,N_22529);
xor U26733 (N_26733,N_23965,N_23148);
xnor U26734 (N_26734,N_24107,N_23621);
xor U26735 (N_26735,N_24698,N_23184);
or U26736 (N_26736,N_23179,N_23413);
and U26737 (N_26737,N_24504,N_22974);
nor U26738 (N_26738,N_22848,N_23189);
or U26739 (N_26739,N_23315,N_23534);
and U26740 (N_26740,N_24062,N_23303);
nand U26741 (N_26741,N_23760,N_22650);
and U26742 (N_26742,N_22566,N_22755);
and U26743 (N_26743,N_24608,N_23402);
and U26744 (N_26744,N_23381,N_23082);
nand U26745 (N_26745,N_24366,N_23081);
xnor U26746 (N_26746,N_24234,N_24678);
or U26747 (N_26747,N_24734,N_24744);
xnor U26748 (N_26748,N_23798,N_22695);
or U26749 (N_26749,N_24677,N_23306);
or U26750 (N_26750,N_24113,N_22575);
xor U26751 (N_26751,N_23018,N_23873);
or U26752 (N_26752,N_23417,N_23270);
nor U26753 (N_26753,N_22787,N_24560);
nand U26754 (N_26754,N_23520,N_23736);
xor U26755 (N_26755,N_23447,N_24749);
nor U26756 (N_26756,N_24078,N_24691);
xnor U26757 (N_26757,N_23347,N_22933);
and U26758 (N_26758,N_23780,N_24546);
or U26759 (N_26759,N_23170,N_22646);
nor U26760 (N_26760,N_22730,N_24065);
or U26761 (N_26761,N_23775,N_24389);
nand U26762 (N_26762,N_23839,N_24779);
and U26763 (N_26763,N_24502,N_24078);
or U26764 (N_26764,N_23291,N_24644);
nor U26765 (N_26765,N_24119,N_23492);
or U26766 (N_26766,N_24102,N_23974);
nor U26767 (N_26767,N_23452,N_24317);
nand U26768 (N_26768,N_23727,N_24396);
and U26769 (N_26769,N_23931,N_24315);
xnor U26770 (N_26770,N_23618,N_23254);
nand U26771 (N_26771,N_24986,N_24514);
xor U26772 (N_26772,N_22773,N_24069);
nand U26773 (N_26773,N_22661,N_23710);
and U26774 (N_26774,N_24344,N_24375);
xor U26775 (N_26775,N_24794,N_22512);
nand U26776 (N_26776,N_23304,N_24486);
nor U26777 (N_26777,N_22915,N_24608);
nand U26778 (N_26778,N_24049,N_24887);
or U26779 (N_26779,N_24291,N_22535);
xor U26780 (N_26780,N_23004,N_23636);
nor U26781 (N_26781,N_24458,N_23511);
or U26782 (N_26782,N_22754,N_23397);
or U26783 (N_26783,N_24940,N_22916);
xnor U26784 (N_26784,N_23451,N_24124);
and U26785 (N_26785,N_24986,N_23615);
xnor U26786 (N_26786,N_24653,N_22731);
nand U26787 (N_26787,N_22615,N_23374);
nand U26788 (N_26788,N_24184,N_22552);
and U26789 (N_26789,N_23272,N_23823);
and U26790 (N_26790,N_24608,N_24773);
and U26791 (N_26791,N_22981,N_22512);
nor U26792 (N_26792,N_23711,N_23561);
xnor U26793 (N_26793,N_23297,N_23052);
nand U26794 (N_26794,N_24936,N_23851);
xnor U26795 (N_26795,N_22957,N_23412);
xnor U26796 (N_26796,N_23498,N_22681);
nand U26797 (N_26797,N_23835,N_23064);
nand U26798 (N_26798,N_23344,N_24266);
nand U26799 (N_26799,N_23261,N_24889);
nand U26800 (N_26800,N_22836,N_22870);
nand U26801 (N_26801,N_22925,N_22624);
nor U26802 (N_26802,N_24442,N_24749);
xnor U26803 (N_26803,N_22632,N_24580);
nor U26804 (N_26804,N_22861,N_24923);
and U26805 (N_26805,N_24935,N_23914);
or U26806 (N_26806,N_23893,N_24876);
and U26807 (N_26807,N_22710,N_22603);
xnor U26808 (N_26808,N_22560,N_23683);
nand U26809 (N_26809,N_23587,N_23551);
and U26810 (N_26810,N_22687,N_23957);
nor U26811 (N_26811,N_24813,N_22659);
and U26812 (N_26812,N_23043,N_24326);
or U26813 (N_26813,N_23191,N_24599);
nand U26814 (N_26814,N_23184,N_22617);
or U26815 (N_26815,N_24450,N_22691);
or U26816 (N_26816,N_24096,N_24001);
nor U26817 (N_26817,N_24771,N_24793);
nand U26818 (N_26818,N_24345,N_22943);
and U26819 (N_26819,N_22935,N_22595);
nor U26820 (N_26820,N_23333,N_24688);
nor U26821 (N_26821,N_23633,N_23023);
nor U26822 (N_26822,N_24689,N_23453);
nand U26823 (N_26823,N_23392,N_23617);
xor U26824 (N_26824,N_23000,N_22718);
nor U26825 (N_26825,N_24853,N_23180);
or U26826 (N_26826,N_22643,N_22609);
or U26827 (N_26827,N_24264,N_24922);
nor U26828 (N_26828,N_24549,N_23156);
nor U26829 (N_26829,N_23197,N_22667);
xor U26830 (N_26830,N_22622,N_23400);
or U26831 (N_26831,N_23736,N_22905);
or U26832 (N_26832,N_24441,N_23135);
and U26833 (N_26833,N_23616,N_24332);
nand U26834 (N_26834,N_24098,N_24917);
xnor U26835 (N_26835,N_23199,N_22562);
nand U26836 (N_26836,N_23188,N_22673);
nand U26837 (N_26837,N_23895,N_23532);
or U26838 (N_26838,N_23586,N_23490);
or U26839 (N_26839,N_24020,N_24805);
or U26840 (N_26840,N_24289,N_22813);
xnor U26841 (N_26841,N_23575,N_24920);
and U26842 (N_26842,N_23425,N_22659);
xnor U26843 (N_26843,N_24197,N_22644);
xnor U26844 (N_26844,N_22696,N_24973);
and U26845 (N_26845,N_23372,N_24394);
and U26846 (N_26846,N_24369,N_23644);
and U26847 (N_26847,N_24651,N_24502);
and U26848 (N_26848,N_23252,N_24853);
nor U26849 (N_26849,N_24218,N_22754);
nor U26850 (N_26850,N_24024,N_22896);
and U26851 (N_26851,N_23758,N_23126);
or U26852 (N_26852,N_23107,N_23486);
nand U26853 (N_26853,N_23324,N_22543);
or U26854 (N_26854,N_24986,N_24563);
or U26855 (N_26855,N_23909,N_22678);
and U26856 (N_26856,N_24773,N_24801);
nand U26857 (N_26857,N_23521,N_23473);
or U26858 (N_26858,N_23193,N_22568);
xor U26859 (N_26859,N_23747,N_23041);
or U26860 (N_26860,N_23053,N_22979);
xor U26861 (N_26861,N_23676,N_24777);
nand U26862 (N_26862,N_22982,N_23698);
xnor U26863 (N_26863,N_22839,N_24693);
nor U26864 (N_26864,N_24645,N_24764);
and U26865 (N_26865,N_24138,N_24817);
xnor U26866 (N_26866,N_22894,N_23208);
and U26867 (N_26867,N_23486,N_23973);
or U26868 (N_26868,N_24694,N_22885);
or U26869 (N_26869,N_22931,N_24492);
xnor U26870 (N_26870,N_24436,N_24874);
or U26871 (N_26871,N_23673,N_24097);
or U26872 (N_26872,N_22881,N_24078);
nor U26873 (N_26873,N_22792,N_24335);
nand U26874 (N_26874,N_23831,N_24451);
and U26875 (N_26875,N_23005,N_24844);
or U26876 (N_26876,N_23300,N_23252);
nor U26877 (N_26877,N_24008,N_23280);
or U26878 (N_26878,N_23242,N_24563);
xor U26879 (N_26879,N_22897,N_24657);
and U26880 (N_26880,N_23906,N_23717);
nor U26881 (N_26881,N_23504,N_24512);
and U26882 (N_26882,N_24725,N_23614);
and U26883 (N_26883,N_22992,N_23864);
and U26884 (N_26884,N_22909,N_22974);
nor U26885 (N_26885,N_24420,N_24370);
and U26886 (N_26886,N_23417,N_23584);
and U26887 (N_26887,N_23787,N_22541);
xor U26888 (N_26888,N_23541,N_24253);
xor U26889 (N_26889,N_22662,N_24722);
xnor U26890 (N_26890,N_24828,N_24209);
or U26891 (N_26891,N_23236,N_24370);
nand U26892 (N_26892,N_22730,N_23160);
nor U26893 (N_26893,N_23760,N_23676);
xnor U26894 (N_26894,N_24263,N_23678);
nor U26895 (N_26895,N_23371,N_23455);
or U26896 (N_26896,N_22574,N_23289);
or U26897 (N_26897,N_23070,N_23699);
nor U26898 (N_26898,N_23409,N_23025);
xnor U26899 (N_26899,N_24957,N_24200);
and U26900 (N_26900,N_23426,N_23003);
nor U26901 (N_26901,N_22830,N_24404);
or U26902 (N_26902,N_24094,N_23373);
and U26903 (N_26903,N_24192,N_22943);
nand U26904 (N_26904,N_23854,N_24064);
xor U26905 (N_26905,N_23288,N_24925);
and U26906 (N_26906,N_23565,N_22702);
xor U26907 (N_26907,N_23993,N_23084);
nor U26908 (N_26908,N_23283,N_22639);
nand U26909 (N_26909,N_23722,N_23657);
nor U26910 (N_26910,N_23037,N_24431);
xor U26911 (N_26911,N_24275,N_23265);
nor U26912 (N_26912,N_24345,N_24294);
nand U26913 (N_26913,N_22644,N_24638);
xnor U26914 (N_26914,N_24519,N_24511);
and U26915 (N_26915,N_23339,N_23370);
nor U26916 (N_26916,N_24417,N_22935);
nor U26917 (N_26917,N_22969,N_23847);
or U26918 (N_26918,N_23747,N_24950);
or U26919 (N_26919,N_23974,N_24632);
nor U26920 (N_26920,N_23553,N_22785);
nor U26921 (N_26921,N_22824,N_22613);
or U26922 (N_26922,N_24253,N_23461);
or U26923 (N_26923,N_22935,N_23395);
or U26924 (N_26924,N_23641,N_24782);
xor U26925 (N_26925,N_23504,N_24080);
nor U26926 (N_26926,N_24647,N_24494);
nor U26927 (N_26927,N_22823,N_23424);
nor U26928 (N_26928,N_24075,N_24486);
xnor U26929 (N_26929,N_24175,N_23348);
or U26930 (N_26930,N_24007,N_24895);
and U26931 (N_26931,N_22643,N_22712);
or U26932 (N_26932,N_24085,N_24651);
nor U26933 (N_26933,N_23635,N_23766);
nor U26934 (N_26934,N_24685,N_23263);
and U26935 (N_26935,N_24638,N_23041);
nor U26936 (N_26936,N_23048,N_23878);
nor U26937 (N_26937,N_22716,N_23318);
nand U26938 (N_26938,N_24997,N_22515);
or U26939 (N_26939,N_23929,N_22613);
or U26940 (N_26940,N_23595,N_23071);
and U26941 (N_26941,N_23115,N_23128);
nor U26942 (N_26942,N_24666,N_24632);
xnor U26943 (N_26943,N_24843,N_24448);
nand U26944 (N_26944,N_22560,N_24431);
xor U26945 (N_26945,N_23359,N_23700);
or U26946 (N_26946,N_24911,N_22649);
nand U26947 (N_26947,N_24235,N_23453);
or U26948 (N_26948,N_23311,N_23033);
nor U26949 (N_26949,N_23574,N_24034);
or U26950 (N_26950,N_24922,N_24716);
xor U26951 (N_26951,N_24995,N_24810);
xor U26952 (N_26952,N_24457,N_22976);
nand U26953 (N_26953,N_24478,N_23130);
and U26954 (N_26954,N_23754,N_23471);
xnor U26955 (N_26955,N_24796,N_22630);
or U26956 (N_26956,N_24338,N_23670);
or U26957 (N_26957,N_23918,N_23360);
or U26958 (N_26958,N_23809,N_23384);
nand U26959 (N_26959,N_22709,N_24909);
or U26960 (N_26960,N_23358,N_22864);
and U26961 (N_26961,N_23894,N_24062);
xor U26962 (N_26962,N_23767,N_23353);
nor U26963 (N_26963,N_24623,N_23201);
xnor U26964 (N_26964,N_24473,N_22965);
and U26965 (N_26965,N_24003,N_23234);
nor U26966 (N_26966,N_24028,N_22803);
nor U26967 (N_26967,N_23745,N_24339);
nand U26968 (N_26968,N_24114,N_22965);
xnor U26969 (N_26969,N_23375,N_23055);
and U26970 (N_26970,N_23054,N_23602);
xnor U26971 (N_26971,N_23402,N_23280);
xor U26972 (N_26972,N_24913,N_23836);
and U26973 (N_26973,N_23382,N_24673);
and U26974 (N_26974,N_24850,N_24431);
xor U26975 (N_26975,N_24414,N_23754);
nand U26976 (N_26976,N_23416,N_23720);
nand U26977 (N_26977,N_22622,N_23955);
and U26978 (N_26978,N_24132,N_23646);
or U26979 (N_26979,N_24530,N_22848);
xor U26980 (N_26980,N_24396,N_23182);
nand U26981 (N_26981,N_23693,N_23547);
nand U26982 (N_26982,N_23370,N_23671);
xnor U26983 (N_26983,N_22520,N_24190);
nor U26984 (N_26984,N_24432,N_22745);
nand U26985 (N_26985,N_23529,N_22986);
xnor U26986 (N_26986,N_24847,N_24459);
or U26987 (N_26987,N_23845,N_24588);
and U26988 (N_26988,N_22769,N_23313);
and U26989 (N_26989,N_23698,N_22882);
xnor U26990 (N_26990,N_23518,N_24826);
and U26991 (N_26991,N_22846,N_23627);
nor U26992 (N_26992,N_24841,N_24094);
or U26993 (N_26993,N_23460,N_23216);
and U26994 (N_26994,N_22606,N_24919);
nor U26995 (N_26995,N_22885,N_22987);
or U26996 (N_26996,N_24581,N_23962);
nor U26997 (N_26997,N_24601,N_22784);
nand U26998 (N_26998,N_24275,N_23655);
nor U26999 (N_26999,N_23891,N_22640);
xor U27000 (N_27000,N_24966,N_22876);
nor U27001 (N_27001,N_23526,N_23089);
nand U27002 (N_27002,N_24274,N_24737);
or U27003 (N_27003,N_24261,N_23288);
nand U27004 (N_27004,N_23077,N_24025);
nand U27005 (N_27005,N_24458,N_23538);
nand U27006 (N_27006,N_23979,N_24933);
and U27007 (N_27007,N_22843,N_24913);
or U27008 (N_27008,N_24436,N_24730);
xor U27009 (N_27009,N_23935,N_22763);
xor U27010 (N_27010,N_23688,N_24375);
nor U27011 (N_27011,N_22844,N_22677);
nor U27012 (N_27012,N_23244,N_24322);
and U27013 (N_27013,N_24451,N_23855);
xnor U27014 (N_27014,N_23902,N_24657);
xnor U27015 (N_27015,N_24344,N_24226);
or U27016 (N_27016,N_23690,N_23168);
nor U27017 (N_27017,N_24782,N_23606);
or U27018 (N_27018,N_23039,N_24971);
nand U27019 (N_27019,N_23528,N_22687);
nand U27020 (N_27020,N_22676,N_24785);
nor U27021 (N_27021,N_24619,N_23707);
xnor U27022 (N_27022,N_22940,N_23518);
nand U27023 (N_27023,N_23597,N_23094);
or U27024 (N_27024,N_24257,N_23273);
and U27025 (N_27025,N_23911,N_23136);
nor U27026 (N_27026,N_23452,N_23648);
nand U27027 (N_27027,N_23327,N_23498);
or U27028 (N_27028,N_23951,N_22812);
or U27029 (N_27029,N_23529,N_23943);
nor U27030 (N_27030,N_24955,N_24856);
nand U27031 (N_27031,N_23305,N_22584);
and U27032 (N_27032,N_22984,N_24332);
and U27033 (N_27033,N_23518,N_24093);
xor U27034 (N_27034,N_24438,N_23287);
nor U27035 (N_27035,N_24886,N_24416);
nor U27036 (N_27036,N_24942,N_23858);
nor U27037 (N_27037,N_23916,N_23574);
nand U27038 (N_27038,N_23375,N_24854);
or U27039 (N_27039,N_24058,N_22921);
or U27040 (N_27040,N_22530,N_23815);
and U27041 (N_27041,N_22647,N_23093);
and U27042 (N_27042,N_23477,N_22735);
xor U27043 (N_27043,N_23986,N_24861);
and U27044 (N_27044,N_24480,N_24282);
and U27045 (N_27045,N_24505,N_24066);
nor U27046 (N_27046,N_23166,N_22659);
or U27047 (N_27047,N_24609,N_22680);
and U27048 (N_27048,N_24854,N_23675);
nand U27049 (N_27049,N_24209,N_24119);
nor U27050 (N_27050,N_23981,N_23609);
or U27051 (N_27051,N_23660,N_24444);
nand U27052 (N_27052,N_22941,N_23111);
xnor U27053 (N_27053,N_23099,N_22741);
or U27054 (N_27054,N_22876,N_23931);
and U27055 (N_27055,N_23085,N_23571);
nand U27056 (N_27056,N_24384,N_22984);
and U27057 (N_27057,N_24525,N_23085);
or U27058 (N_27058,N_24037,N_23132);
xnor U27059 (N_27059,N_24770,N_24971);
nand U27060 (N_27060,N_24115,N_24135);
and U27061 (N_27061,N_23784,N_23084);
nor U27062 (N_27062,N_22810,N_22851);
nand U27063 (N_27063,N_23312,N_23073);
nand U27064 (N_27064,N_23080,N_24659);
nor U27065 (N_27065,N_23923,N_23066);
xor U27066 (N_27066,N_23149,N_23191);
or U27067 (N_27067,N_24536,N_24690);
nand U27068 (N_27068,N_24206,N_24576);
and U27069 (N_27069,N_24274,N_23356);
xnor U27070 (N_27070,N_23632,N_22604);
and U27071 (N_27071,N_24849,N_23722);
and U27072 (N_27072,N_24691,N_24568);
or U27073 (N_27073,N_24383,N_22840);
nor U27074 (N_27074,N_24050,N_24218);
and U27075 (N_27075,N_24181,N_23733);
xor U27076 (N_27076,N_22637,N_24757);
or U27077 (N_27077,N_22976,N_23306);
nand U27078 (N_27078,N_22597,N_23478);
xor U27079 (N_27079,N_24947,N_24714);
xor U27080 (N_27080,N_23723,N_23631);
nand U27081 (N_27081,N_24733,N_23451);
nor U27082 (N_27082,N_23870,N_22823);
nor U27083 (N_27083,N_23918,N_23434);
nand U27084 (N_27084,N_24549,N_24283);
nor U27085 (N_27085,N_24116,N_24952);
xnor U27086 (N_27086,N_24495,N_23837);
xnor U27087 (N_27087,N_23458,N_24261);
xnor U27088 (N_27088,N_23678,N_23367);
and U27089 (N_27089,N_24892,N_22730);
nor U27090 (N_27090,N_23582,N_23415);
nor U27091 (N_27091,N_23532,N_23261);
nor U27092 (N_27092,N_23904,N_24588);
or U27093 (N_27093,N_22668,N_23321);
and U27094 (N_27094,N_22797,N_24732);
xor U27095 (N_27095,N_24922,N_24125);
nand U27096 (N_27096,N_23376,N_22925);
nand U27097 (N_27097,N_24782,N_22656);
xnor U27098 (N_27098,N_24309,N_24734);
nand U27099 (N_27099,N_23308,N_24963);
nor U27100 (N_27100,N_24795,N_24045);
xnor U27101 (N_27101,N_24867,N_22773);
xnor U27102 (N_27102,N_23773,N_24948);
nor U27103 (N_27103,N_24519,N_24145);
xnor U27104 (N_27104,N_24898,N_22872);
xor U27105 (N_27105,N_23112,N_23807);
or U27106 (N_27106,N_24283,N_23481);
nand U27107 (N_27107,N_24131,N_24257);
or U27108 (N_27108,N_22903,N_24710);
or U27109 (N_27109,N_24065,N_23416);
or U27110 (N_27110,N_23463,N_23736);
or U27111 (N_27111,N_24790,N_22682);
xor U27112 (N_27112,N_22891,N_24979);
xor U27113 (N_27113,N_24712,N_23397);
and U27114 (N_27114,N_24688,N_23762);
or U27115 (N_27115,N_24825,N_23886);
or U27116 (N_27116,N_24203,N_23404);
nand U27117 (N_27117,N_23026,N_23516);
nand U27118 (N_27118,N_24072,N_23955);
and U27119 (N_27119,N_22621,N_22874);
nor U27120 (N_27120,N_23628,N_22774);
nor U27121 (N_27121,N_23269,N_23195);
and U27122 (N_27122,N_23188,N_23984);
and U27123 (N_27123,N_24313,N_23736);
xnor U27124 (N_27124,N_24625,N_24726);
nor U27125 (N_27125,N_23900,N_23481);
and U27126 (N_27126,N_23334,N_23641);
and U27127 (N_27127,N_24513,N_23427);
xor U27128 (N_27128,N_24773,N_23494);
nand U27129 (N_27129,N_22645,N_22630);
nand U27130 (N_27130,N_23703,N_23028);
xnor U27131 (N_27131,N_23930,N_23102);
and U27132 (N_27132,N_23529,N_22597);
or U27133 (N_27133,N_23180,N_24585);
nand U27134 (N_27134,N_23379,N_23788);
nand U27135 (N_27135,N_23985,N_24862);
and U27136 (N_27136,N_23514,N_24733);
nand U27137 (N_27137,N_24807,N_22546);
and U27138 (N_27138,N_22598,N_23150);
or U27139 (N_27139,N_23912,N_24744);
nor U27140 (N_27140,N_24353,N_23450);
xnor U27141 (N_27141,N_23435,N_22538);
and U27142 (N_27142,N_24206,N_24679);
and U27143 (N_27143,N_23813,N_22848);
or U27144 (N_27144,N_24912,N_24563);
or U27145 (N_27145,N_23916,N_24579);
nand U27146 (N_27146,N_24192,N_22568);
xnor U27147 (N_27147,N_22937,N_24224);
nor U27148 (N_27148,N_22943,N_24504);
or U27149 (N_27149,N_23832,N_24151);
nor U27150 (N_27150,N_22852,N_23432);
or U27151 (N_27151,N_24137,N_22556);
nand U27152 (N_27152,N_23070,N_23183);
xor U27153 (N_27153,N_24325,N_24046);
xnor U27154 (N_27154,N_24863,N_23616);
nand U27155 (N_27155,N_23357,N_22588);
and U27156 (N_27156,N_23342,N_22708);
or U27157 (N_27157,N_23690,N_22913);
nand U27158 (N_27158,N_24756,N_23528);
nand U27159 (N_27159,N_22947,N_23565);
nand U27160 (N_27160,N_24290,N_23217);
nand U27161 (N_27161,N_24399,N_24658);
and U27162 (N_27162,N_23336,N_23506);
nand U27163 (N_27163,N_23469,N_23227);
nand U27164 (N_27164,N_23752,N_24400);
nand U27165 (N_27165,N_23922,N_24864);
nor U27166 (N_27166,N_22784,N_23189);
nor U27167 (N_27167,N_23897,N_23439);
or U27168 (N_27168,N_24245,N_24444);
nand U27169 (N_27169,N_23937,N_24094);
or U27170 (N_27170,N_24645,N_22500);
xnor U27171 (N_27171,N_24435,N_22943);
xor U27172 (N_27172,N_22826,N_23084);
or U27173 (N_27173,N_23029,N_23170);
and U27174 (N_27174,N_24639,N_22903);
nor U27175 (N_27175,N_23972,N_24697);
and U27176 (N_27176,N_22908,N_22990);
and U27177 (N_27177,N_22682,N_24167);
and U27178 (N_27178,N_24700,N_24645);
nor U27179 (N_27179,N_23167,N_24098);
xor U27180 (N_27180,N_24813,N_23321);
or U27181 (N_27181,N_24798,N_23784);
and U27182 (N_27182,N_22687,N_23050);
and U27183 (N_27183,N_23829,N_23764);
or U27184 (N_27184,N_24343,N_23464);
or U27185 (N_27185,N_24184,N_24933);
and U27186 (N_27186,N_22758,N_24487);
and U27187 (N_27187,N_24419,N_22877);
nand U27188 (N_27188,N_22779,N_22534);
and U27189 (N_27189,N_23493,N_24494);
or U27190 (N_27190,N_24377,N_23273);
xor U27191 (N_27191,N_24554,N_23041);
or U27192 (N_27192,N_24388,N_24084);
nand U27193 (N_27193,N_22566,N_22738);
or U27194 (N_27194,N_24708,N_24846);
or U27195 (N_27195,N_23345,N_24397);
nor U27196 (N_27196,N_22667,N_22720);
and U27197 (N_27197,N_22523,N_23546);
nand U27198 (N_27198,N_22979,N_23693);
xnor U27199 (N_27199,N_22554,N_23344);
and U27200 (N_27200,N_23528,N_22787);
and U27201 (N_27201,N_23841,N_24869);
nor U27202 (N_27202,N_22606,N_24844);
nor U27203 (N_27203,N_23222,N_23074);
and U27204 (N_27204,N_22852,N_23117);
and U27205 (N_27205,N_24202,N_22757);
nor U27206 (N_27206,N_23631,N_24598);
nand U27207 (N_27207,N_24546,N_24482);
xnor U27208 (N_27208,N_23850,N_23734);
or U27209 (N_27209,N_23881,N_22941);
nor U27210 (N_27210,N_24593,N_23628);
and U27211 (N_27211,N_22804,N_24675);
and U27212 (N_27212,N_22741,N_23035);
and U27213 (N_27213,N_24257,N_24559);
or U27214 (N_27214,N_23192,N_22586);
xor U27215 (N_27215,N_23998,N_24025);
xor U27216 (N_27216,N_24438,N_23542);
and U27217 (N_27217,N_22918,N_24500);
xor U27218 (N_27218,N_22824,N_22884);
or U27219 (N_27219,N_24905,N_23645);
nor U27220 (N_27220,N_23475,N_23492);
nand U27221 (N_27221,N_23345,N_24386);
or U27222 (N_27222,N_23434,N_24506);
nor U27223 (N_27223,N_23982,N_24203);
nand U27224 (N_27224,N_24468,N_22837);
or U27225 (N_27225,N_23813,N_23612);
nand U27226 (N_27226,N_23197,N_23465);
nand U27227 (N_27227,N_22563,N_24536);
xnor U27228 (N_27228,N_24841,N_23214);
xor U27229 (N_27229,N_24195,N_23759);
and U27230 (N_27230,N_24087,N_23306);
or U27231 (N_27231,N_23677,N_23340);
xnor U27232 (N_27232,N_24177,N_23516);
and U27233 (N_27233,N_23416,N_22585);
and U27234 (N_27234,N_24173,N_23128);
and U27235 (N_27235,N_23704,N_22586);
nand U27236 (N_27236,N_24614,N_23058);
or U27237 (N_27237,N_24812,N_22623);
nand U27238 (N_27238,N_23618,N_22563);
nor U27239 (N_27239,N_23376,N_24132);
xnor U27240 (N_27240,N_23934,N_23484);
or U27241 (N_27241,N_24898,N_22979);
nand U27242 (N_27242,N_23593,N_23337);
nand U27243 (N_27243,N_23724,N_23715);
and U27244 (N_27244,N_24695,N_24930);
nor U27245 (N_27245,N_24641,N_23368);
nand U27246 (N_27246,N_23282,N_22570);
nand U27247 (N_27247,N_23979,N_22691);
and U27248 (N_27248,N_24416,N_22758);
and U27249 (N_27249,N_24779,N_24851);
xor U27250 (N_27250,N_22814,N_23862);
and U27251 (N_27251,N_24088,N_22611);
and U27252 (N_27252,N_23908,N_23242);
and U27253 (N_27253,N_24663,N_22836);
xor U27254 (N_27254,N_23072,N_23493);
or U27255 (N_27255,N_22618,N_23717);
and U27256 (N_27256,N_22974,N_22957);
or U27257 (N_27257,N_24602,N_23794);
nor U27258 (N_27258,N_24074,N_23338);
nand U27259 (N_27259,N_23495,N_22859);
and U27260 (N_27260,N_22807,N_24534);
nor U27261 (N_27261,N_23582,N_23666);
or U27262 (N_27262,N_24920,N_23126);
xor U27263 (N_27263,N_24056,N_23831);
xnor U27264 (N_27264,N_22766,N_23608);
nor U27265 (N_27265,N_22732,N_24494);
xnor U27266 (N_27266,N_23025,N_23876);
xor U27267 (N_27267,N_24689,N_24678);
or U27268 (N_27268,N_23098,N_23322);
nand U27269 (N_27269,N_24313,N_24732);
xnor U27270 (N_27270,N_22700,N_23063);
and U27271 (N_27271,N_24381,N_24937);
nand U27272 (N_27272,N_24002,N_23386);
and U27273 (N_27273,N_23231,N_23075);
or U27274 (N_27274,N_22716,N_23730);
nor U27275 (N_27275,N_23946,N_23700);
nor U27276 (N_27276,N_24353,N_24462);
or U27277 (N_27277,N_24720,N_23770);
or U27278 (N_27278,N_23422,N_24369);
nand U27279 (N_27279,N_24058,N_23643);
nor U27280 (N_27280,N_23301,N_23487);
xor U27281 (N_27281,N_24946,N_24913);
nand U27282 (N_27282,N_24497,N_23952);
and U27283 (N_27283,N_24182,N_23376);
and U27284 (N_27284,N_22888,N_23987);
xnor U27285 (N_27285,N_23453,N_23521);
or U27286 (N_27286,N_23585,N_23675);
nand U27287 (N_27287,N_23001,N_23991);
xnor U27288 (N_27288,N_23727,N_23293);
nor U27289 (N_27289,N_23377,N_22785);
and U27290 (N_27290,N_23803,N_24600);
nand U27291 (N_27291,N_23295,N_23541);
nand U27292 (N_27292,N_24273,N_22886);
and U27293 (N_27293,N_24211,N_22565);
or U27294 (N_27294,N_23742,N_24755);
and U27295 (N_27295,N_24082,N_23604);
and U27296 (N_27296,N_24387,N_23931);
nand U27297 (N_27297,N_23878,N_24510);
xnor U27298 (N_27298,N_24587,N_22711);
nor U27299 (N_27299,N_23879,N_24627);
nor U27300 (N_27300,N_23530,N_23701);
nand U27301 (N_27301,N_23321,N_22965);
and U27302 (N_27302,N_22790,N_24092);
or U27303 (N_27303,N_22714,N_22567);
xnor U27304 (N_27304,N_24086,N_24521);
or U27305 (N_27305,N_24455,N_24247);
and U27306 (N_27306,N_24305,N_23808);
nand U27307 (N_27307,N_24962,N_22927);
or U27308 (N_27308,N_23338,N_24710);
xor U27309 (N_27309,N_24248,N_24606);
and U27310 (N_27310,N_22517,N_23230);
and U27311 (N_27311,N_23557,N_24883);
or U27312 (N_27312,N_22567,N_23947);
nand U27313 (N_27313,N_24046,N_23395);
or U27314 (N_27314,N_24288,N_23834);
nand U27315 (N_27315,N_23210,N_24078);
and U27316 (N_27316,N_23686,N_24164);
or U27317 (N_27317,N_23863,N_23493);
nand U27318 (N_27318,N_24846,N_24667);
or U27319 (N_27319,N_22666,N_23111);
nor U27320 (N_27320,N_24648,N_23272);
nor U27321 (N_27321,N_23827,N_23273);
nand U27322 (N_27322,N_23833,N_22893);
nor U27323 (N_27323,N_22803,N_24560);
or U27324 (N_27324,N_23369,N_24026);
xnor U27325 (N_27325,N_23219,N_23364);
nor U27326 (N_27326,N_24889,N_24216);
nor U27327 (N_27327,N_22896,N_24970);
and U27328 (N_27328,N_23376,N_24738);
or U27329 (N_27329,N_23491,N_23143);
xor U27330 (N_27330,N_23210,N_22628);
nor U27331 (N_27331,N_23831,N_22873);
or U27332 (N_27332,N_22656,N_23081);
nor U27333 (N_27333,N_23071,N_24612);
and U27334 (N_27334,N_24097,N_23786);
xnor U27335 (N_27335,N_23005,N_22853);
nor U27336 (N_27336,N_23858,N_23926);
xnor U27337 (N_27337,N_22688,N_24180);
nor U27338 (N_27338,N_24560,N_24355);
nor U27339 (N_27339,N_22861,N_22530);
nand U27340 (N_27340,N_24697,N_22907);
nor U27341 (N_27341,N_23055,N_24339);
xnor U27342 (N_27342,N_24151,N_24743);
and U27343 (N_27343,N_22646,N_23815);
nor U27344 (N_27344,N_24380,N_24542);
nor U27345 (N_27345,N_24987,N_24644);
nand U27346 (N_27346,N_23659,N_22994);
and U27347 (N_27347,N_22695,N_23614);
nor U27348 (N_27348,N_22712,N_24916);
or U27349 (N_27349,N_24951,N_24958);
or U27350 (N_27350,N_23407,N_23748);
nor U27351 (N_27351,N_24150,N_22810);
nor U27352 (N_27352,N_24574,N_23306);
nor U27353 (N_27353,N_23042,N_24719);
or U27354 (N_27354,N_23096,N_23149);
xnor U27355 (N_27355,N_23261,N_22581);
and U27356 (N_27356,N_24148,N_23550);
and U27357 (N_27357,N_24823,N_24459);
nand U27358 (N_27358,N_23169,N_23524);
and U27359 (N_27359,N_24574,N_22535);
and U27360 (N_27360,N_23990,N_23485);
nor U27361 (N_27361,N_23092,N_22864);
nor U27362 (N_27362,N_22933,N_23553);
and U27363 (N_27363,N_23684,N_23115);
nand U27364 (N_27364,N_24072,N_23905);
nor U27365 (N_27365,N_23633,N_24280);
nand U27366 (N_27366,N_23955,N_23931);
or U27367 (N_27367,N_23057,N_23214);
nor U27368 (N_27368,N_23916,N_24669);
nor U27369 (N_27369,N_22901,N_24781);
or U27370 (N_27370,N_23801,N_23090);
or U27371 (N_27371,N_22717,N_23596);
and U27372 (N_27372,N_24912,N_22965);
nand U27373 (N_27373,N_23679,N_23070);
nor U27374 (N_27374,N_24282,N_24088);
nor U27375 (N_27375,N_24973,N_24934);
or U27376 (N_27376,N_23841,N_22674);
nor U27377 (N_27377,N_22504,N_22909);
and U27378 (N_27378,N_24219,N_24511);
xnor U27379 (N_27379,N_24867,N_24271);
or U27380 (N_27380,N_24082,N_22668);
and U27381 (N_27381,N_24771,N_24479);
nand U27382 (N_27382,N_24928,N_23830);
nor U27383 (N_27383,N_24425,N_24352);
nand U27384 (N_27384,N_24318,N_23350);
nor U27385 (N_27385,N_23163,N_24904);
xnor U27386 (N_27386,N_24898,N_22576);
or U27387 (N_27387,N_24056,N_23607);
and U27388 (N_27388,N_24559,N_23218);
and U27389 (N_27389,N_23032,N_22949);
or U27390 (N_27390,N_24569,N_22508);
or U27391 (N_27391,N_22744,N_22971);
nand U27392 (N_27392,N_24232,N_22578);
or U27393 (N_27393,N_23731,N_23134);
or U27394 (N_27394,N_23991,N_23704);
and U27395 (N_27395,N_23341,N_23723);
nand U27396 (N_27396,N_23503,N_23432);
nor U27397 (N_27397,N_24471,N_23568);
nand U27398 (N_27398,N_24866,N_22862);
xor U27399 (N_27399,N_23462,N_24422);
nor U27400 (N_27400,N_22940,N_23861);
xor U27401 (N_27401,N_23416,N_23021);
and U27402 (N_27402,N_24148,N_23341);
or U27403 (N_27403,N_23430,N_24173);
nand U27404 (N_27404,N_24812,N_24037);
and U27405 (N_27405,N_22872,N_23327);
and U27406 (N_27406,N_22868,N_23754);
nand U27407 (N_27407,N_23748,N_23645);
nand U27408 (N_27408,N_23316,N_23145);
nand U27409 (N_27409,N_22970,N_23357);
xnor U27410 (N_27410,N_23372,N_23223);
nand U27411 (N_27411,N_24993,N_24531);
or U27412 (N_27412,N_24283,N_23678);
xor U27413 (N_27413,N_24102,N_23972);
and U27414 (N_27414,N_23931,N_23649);
nand U27415 (N_27415,N_23383,N_24029);
xor U27416 (N_27416,N_23130,N_24930);
nor U27417 (N_27417,N_23183,N_24608);
and U27418 (N_27418,N_24190,N_24406);
nor U27419 (N_27419,N_23445,N_24065);
and U27420 (N_27420,N_24440,N_22518);
nand U27421 (N_27421,N_24560,N_24229);
nand U27422 (N_27422,N_24875,N_23701);
and U27423 (N_27423,N_22922,N_24658);
or U27424 (N_27424,N_24098,N_24735);
and U27425 (N_27425,N_23109,N_22922);
and U27426 (N_27426,N_23874,N_23892);
nand U27427 (N_27427,N_24240,N_22684);
nor U27428 (N_27428,N_22747,N_23522);
nand U27429 (N_27429,N_23466,N_23664);
nor U27430 (N_27430,N_23902,N_24542);
and U27431 (N_27431,N_23630,N_23493);
xor U27432 (N_27432,N_22846,N_22841);
xor U27433 (N_27433,N_24808,N_24523);
xnor U27434 (N_27434,N_24436,N_22526);
nand U27435 (N_27435,N_24453,N_23886);
nor U27436 (N_27436,N_23786,N_24979);
xor U27437 (N_27437,N_23492,N_22733);
and U27438 (N_27438,N_24890,N_24626);
nor U27439 (N_27439,N_23799,N_24644);
nor U27440 (N_27440,N_22849,N_23204);
and U27441 (N_27441,N_23101,N_23515);
or U27442 (N_27442,N_23362,N_22922);
nand U27443 (N_27443,N_23471,N_24786);
xnor U27444 (N_27444,N_23193,N_23262);
nor U27445 (N_27445,N_23724,N_23484);
and U27446 (N_27446,N_22722,N_24583);
nand U27447 (N_27447,N_24898,N_24760);
xor U27448 (N_27448,N_24263,N_23171);
nor U27449 (N_27449,N_24578,N_24910);
nand U27450 (N_27450,N_24629,N_24720);
or U27451 (N_27451,N_22732,N_24728);
or U27452 (N_27452,N_23183,N_24323);
nor U27453 (N_27453,N_24201,N_24994);
and U27454 (N_27454,N_22630,N_24947);
nor U27455 (N_27455,N_24201,N_23306);
and U27456 (N_27456,N_23356,N_24993);
xor U27457 (N_27457,N_24211,N_23349);
and U27458 (N_27458,N_22891,N_23685);
nor U27459 (N_27459,N_24513,N_23315);
xnor U27460 (N_27460,N_24435,N_24971);
xnor U27461 (N_27461,N_23552,N_22634);
nor U27462 (N_27462,N_23944,N_23465);
xnor U27463 (N_27463,N_24150,N_24916);
xor U27464 (N_27464,N_23431,N_23487);
nor U27465 (N_27465,N_23690,N_23500);
xnor U27466 (N_27466,N_22842,N_24883);
nor U27467 (N_27467,N_23287,N_23095);
nand U27468 (N_27468,N_23671,N_23054);
xor U27469 (N_27469,N_24958,N_24681);
and U27470 (N_27470,N_23071,N_24901);
and U27471 (N_27471,N_24575,N_23590);
xor U27472 (N_27472,N_24015,N_23787);
nor U27473 (N_27473,N_23669,N_24500);
and U27474 (N_27474,N_23795,N_24286);
nor U27475 (N_27475,N_23534,N_23539);
and U27476 (N_27476,N_24290,N_24611);
nand U27477 (N_27477,N_24542,N_24872);
or U27478 (N_27478,N_23068,N_23735);
nand U27479 (N_27479,N_24469,N_23709);
or U27480 (N_27480,N_24910,N_23396);
or U27481 (N_27481,N_23725,N_23052);
and U27482 (N_27482,N_23120,N_23049);
and U27483 (N_27483,N_22749,N_23144);
xor U27484 (N_27484,N_24272,N_23379);
and U27485 (N_27485,N_24242,N_22958);
xor U27486 (N_27486,N_24438,N_24884);
nor U27487 (N_27487,N_24347,N_22631);
or U27488 (N_27488,N_22891,N_22794);
nand U27489 (N_27489,N_22855,N_24425);
nand U27490 (N_27490,N_22708,N_23070);
nor U27491 (N_27491,N_24109,N_22803);
or U27492 (N_27492,N_23185,N_23141);
nor U27493 (N_27493,N_23069,N_24970);
nor U27494 (N_27494,N_23642,N_23535);
xor U27495 (N_27495,N_24732,N_22537);
nand U27496 (N_27496,N_22847,N_24712);
nor U27497 (N_27497,N_24718,N_24906);
nand U27498 (N_27498,N_24611,N_23063);
xor U27499 (N_27499,N_23977,N_24591);
or U27500 (N_27500,N_25342,N_26004);
xnor U27501 (N_27501,N_27142,N_25121);
nand U27502 (N_27502,N_26904,N_25625);
xor U27503 (N_27503,N_25716,N_26268);
nand U27504 (N_27504,N_26378,N_25129);
or U27505 (N_27505,N_25918,N_26459);
nand U27506 (N_27506,N_25046,N_26149);
nor U27507 (N_27507,N_25854,N_26440);
xnor U27508 (N_27508,N_25627,N_27038);
nand U27509 (N_27509,N_26603,N_26607);
xor U27510 (N_27510,N_25325,N_25338);
or U27511 (N_27511,N_25025,N_26157);
xor U27512 (N_27512,N_25041,N_25305);
nand U27513 (N_27513,N_25717,N_27018);
nor U27514 (N_27514,N_27310,N_26439);
nor U27515 (N_27515,N_26698,N_25761);
xnor U27516 (N_27516,N_25950,N_27254);
nand U27517 (N_27517,N_25240,N_27364);
nand U27518 (N_27518,N_25150,N_27279);
nand U27519 (N_27519,N_25005,N_27218);
nand U27520 (N_27520,N_25275,N_25406);
xnor U27521 (N_27521,N_27007,N_25862);
and U27522 (N_27522,N_26708,N_26019);
xnor U27523 (N_27523,N_26688,N_25510);
nand U27524 (N_27524,N_26505,N_26065);
or U27525 (N_27525,N_26283,N_27098);
and U27526 (N_27526,N_25254,N_26976);
or U27527 (N_27527,N_25418,N_27325);
and U27528 (N_27528,N_26430,N_26160);
nor U27529 (N_27529,N_25927,N_26547);
nand U27530 (N_27530,N_27297,N_25459);
nand U27531 (N_27531,N_26108,N_27300);
and U27532 (N_27532,N_26363,N_27049);
or U27533 (N_27533,N_26189,N_25452);
and U27534 (N_27534,N_25273,N_27406);
xor U27535 (N_27535,N_25888,N_26828);
nand U27536 (N_27536,N_26248,N_25394);
and U27537 (N_27537,N_25614,N_26204);
nor U27538 (N_27538,N_25742,N_27008);
xnor U27539 (N_27539,N_25944,N_27308);
or U27540 (N_27540,N_25965,N_25955);
and U27541 (N_27541,N_25904,N_26826);
nor U27542 (N_27542,N_26765,N_27210);
xor U27543 (N_27543,N_26924,N_27052);
xor U27544 (N_27544,N_25568,N_25815);
or U27545 (N_27545,N_25086,N_25577);
nor U27546 (N_27546,N_27138,N_25163);
nor U27547 (N_27547,N_25045,N_25047);
xnor U27548 (N_27548,N_26866,N_25509);
nand U27549 (N_27549,N_25424,N_26062);
nand U27550 (N_27550,N_25177,N_27075);
nand U27551 (N_27551,N_26519,N_26344);
and U27552 (N_27552,N_26389,N_27477);
xor U27553 (N_27553,N_27175,N_25170);
nor U27554 (N_27554,N_25304,N_26721);
and U27555 (N_27555,N_25724,N_25668);
nor U27556 (N_27556,N_25503,N_26234);
or U27557 (N_27557,N_25658,N_26402);
nor U27558 (N_27558,N_26461,N_27078);
or U27559 (N_27559,N_25663,N_27436);
and U27560 (N_27560,N_26984,N_27013);
and U27561 (N_27561,N_27378,N_25286);
nor U27562 (N_27562,N_27022,N_26096);
xnor U27563 (N_27563,N_26627,N_26712);
and U27564 (N_27564,N_27041,N_25922);
and U27565 (N_27565,N_27226,N_26791);
nand U27566 (N_27566,N_27445,N_27459);
or U27567 (N_27567,N_26464,N_26396);
or U27568 (N_27568,N_27331,N_27021);
nand U27569 (N_27569,N_26507,N_25814);
nor U27570 (N_27570,N_25383,N_26905);
xnor U27571 (N_27571,N_27489,N_25091);
xor U27572 (N_27572,N_27404,N_25841);
nand U27573 (N_27573,N_26284,N_25554);
or U27574 (N_27574,N_25237,N_25136);
or U27575 (N_27575,N_26832,N_26111);
or U27576 (N_27576,N_26636,N_26939);
xor U27577 (N_27577,N_26117,N_26563);
nand U27578 (N_27578,N_25594,N_26576);
xnor U27579 (N_27579,N_26139,N_25068);
and U27580 (N_27580,N_26960,N_25032);
nand U27581 (N_27581,N_25592,N_26305);
nand U27582 (N_27582,N_25781,N_25793);
and U27583 (N_27583,N_26083,N_27464);
xnor U27584 (N_27584,N_25337,N_26035);
nand U27585 (N_27585,N_25680,N_26289);
nor U27586 (N_27586,N_25193,N_25480);
nor U27587 (N_27587,N_27143,N_25849);
nor U27588 (N_27588,N_26129,N_26333);
and U27589 (N_27589,N_25699,N_25312);
nand U27590 (N_27590,N_25514,N_25882);
nand U27591 (N_27591,N_25207,N_25903);
or U27592 (N_27592,N_25789,N_25948);
and U27593 (N_27593,N_25544,N_26038);
nand U27594 (N_27594,N_26392,N_26938);
and U27595 (N_27595,N_25479,N_25930);
nand U27596 (N_27596,N_25428,N_27133);
nor U27597 (N_27597,N_27189,N_26020);
nand U27598 (N_27598,N_25249,N_26867);
nor U27599 (N_27599,N_26114,N_26818);
or U27600 (N_27600,N_27322,N_25727);
xor U27601 (N_27601,N_25077,N_26612);
and U27602 (N_27602,N_26314,N_27330);
xnor U27603 (N_27603,N_25593,N_26123);
and U27604 (N_27604,N_25219,N_25106);
and U27605 (N_27605,N_25661,N_26957);
nand U27606 (N_27606,N_25471,N_25453);
or U27607 (N_27607,N_27301,N_26029);
and U27608 (N_27608,N_25739,N_25199);
nand U27609 (N_27609,N_25518,N_26266);
and U27610 (N_27610,N_25116,N_26777);
xor U27611 (N_27611,N_25547,N_25075);
xnor U27612 (N_27612,N_26794,N_25203);
xnor U27613 (N_27613,N_27357,N_26012);
and U27614 (N_27614,N_27213,N_26232);
xnor U27615 (N_27615,N_25819,N_25560);
or U27616 (N_27616,N_27263,N_26931);
nand U27617 (N_27617,N_27177,N_25691);
nand U27618 (N_27618,N_26571,N_26550);
or U27619 (N_27619,N_26328,N_26713);
nor U27620 (N_27620,N_25248,N_27043);
nor U27621 (N_27621,N_26608,N_27244);
xnor U27622 (N_27622,N_26492,N_25654);
or U27623 (N_27623,N_25111,N_25039);
xnor U27624 (N_27624,N_25519,N_26021);
or U27625 (N_27625,N_27173,N_26041);
and U27626 (N_27626,N_26558,N_25335);
and U27627 (N_27627,N_26143,N_25541);
or U27628 (N_27628,N_25468,N_26176);
nor U27629 (N_27629,N_25701,N_25404);
nand U27630 (N_27630,N_26733,N_26231);
nand U27631 (N_27631,N_26899,N_27207);
and U27632 (N_27632,N_26452,N_26512);
xor U27633 (N_27633,N_27024,N_25164);
nor U27634 (N_27634,N_25900,N_26748);
nor U27635 (N_27635,N_27487,N_27296);
or U27636 (N_27636,N_27382,N_25341);
nor U27637 (N_27637,N_25863,N_26634);
and U27638 (N_27638,N_25413,N_26797);
and U27639 (N_27639,N_26564,N_26103);
nand U27640 (N_27640,N_25787,N_25443);
xor U27641 (N_27641,N_26925,N_25396);
nor U27642 (N_27642,N_26953,N_25268);
or U27643 (N_27643,N_26187,N_26124);
xor U27644 (N_27644,N_27299,N_25125);
nand U27645 (N_27645,N_26584,N_26438);
and U27646 (N_27646,N_26730,N_25651);
nor U27647 (N_27647,N_25957,N_26329);
and U27648 (N_27648,N_25195,N_26516);
nand U27649 (N_27649,N_25392,N_27433);
nor U27650 (N_27650,N_26660,N_27232);
nand U27651 (N_27651,N_25719,N_26849);
xnor U27652 (N_27652,N_27336,N_26731);
or U27653 (N_27653,N_25079,N_27412);
xor U27654 (N_27654,N_27395,N_25867);
xnor U27655 (N_27655,N_25543,N_26705);
nor U27656 (N_27656,N_27202,N_25878);
and U27657 (N_27657,N_27221,N_25721);
nor U27658 (N_27658,N_27381,N_25178);
nand U27659 (N_27659,N_26127,N_26413);
or U27660 (N_27660,N_27397,N_25104);
xnor U27661 (N_27661,N_25036,N_25650);
and U27662 (N_27662,N_26914,N_27060);
nor U27663 (N_27663,N_25576,N_27039);
or U27664 (N_27664,N_26592,N_26493);
and U27665 (N_27665,N_25314,N_26681);
and U27666 (N_27666,N_25364,N_25843);
and U27667 (N_27667,N_26572,N_25081);
xnor U27668 (N_27668,N_25154,N_25209);
nor U27669 (N_27669,N_27063,N_25901);
and U27670 (N_27670,N_26495,N_27341);
or U27671 (N_27671,N_26435,N_26170);
or U27672 (N_27672,N_26784,N_25708);
or U27673 (N_27673,N_25945,N_25848);
nor U27674 (N_27674,N_26478,N_26741);
nor U27675 (N_27675,N_25282,N_26851);
and U27676 (N_27676,N_26726,N_25967);
nand U27677 (N_27677,N_27234,N_26319);
nand U27678 (N_27678,N_27214,N_26001);
nor U27679 (N_27679,N_27256,N_26715);
xor U27680 (N_27680,N_25968,N_26522);
nand U27681 (N_27681,N_25958,N_27014);
or U27682 (N_27682,N_26222,N_27485);
or U27683 (N_27683,N_26729,N_26624);
or U27684 (N_27684,N_27385,N_26936);
and U27685 (N_27685,N_26874,N_25504);
nor U27686 (N_27686,N_26207,N_27134);
xnor U27687 (N_27687,N_25052,N_26467);
nor U27688 (N_27688,N_26946,N_25498);
xnor U27689 (N_27689,N_26372,N_25629);
and U27690 (N_27690,N_26498,N_25871);
xnor U27691 (N_27691,N_25357,N_27276);
and U27692 (N_27692,N_25458,N_26227);
nor U27693 (N_27693,N_25756,N_26484);
nand U27694 (N_27694,N_27199,N_25358);
nand U27695 (N_27695,N_25261,N_25135);
xnor U27696 (N_27696,N_27118,N_26393);
or U27697 (N_27697,N_25931,N_26906);
nor U27698 (N_27698,N_25983,N_26552);
or U27699 (N_27699,N_25331,N_25709);
or U27700 (N_27700,N_25251,N_25346);
nand U27701 (N_27701,N_25360,N_25559);
and U27702 (N_27702,N_27344,N_27170);
nand U27703 (N_27703,N_25776,N_26412);
or U27704 (N_27704,N_26813,N_25430);
nand U27705 (N_27705,N_25907,N_26026);
nand U27706 (N_27706,N_26542,N_25890);
and U27707 (N_27707,N_27200,N_25087);
or U27708 (N_27708,N_25398,N_26643);
or U27709 (N_27709,N_26480,N_25235);
nand U27710 (N_27710,N_27291,N_27122);
nor U27711 (N_27711,N_25940,N_26320);
or U27712 (N_27712,N_26864,N_25711);
or U27713 (N_27713,N_25946,N_26738);
nor U27714 (N_27714,N_26064,N_26561);
xor U27715 (N_27715,N_26311,N_27069);
nand U27716 (N_27716,N_25905,N_25018);
nand U27717 (N_27717,N_25806,N_26959);
or U27718 (N_27718,N_25666,N_27027);
and U27719 (N_27719,N_27194,N_25085);
or U27720 (N_27720,N_27083,N_26089);
nor U27721 (N_27721,N_26782,N_27298);
nor U27722 (N_27722,N_26743,N_26657);
and U27723 (N_27723,N_27411,N_27313);
nand U27724 (N_27724,N_26274,N_25124);
and U27725 (N_27725,N_26555,N_27281);
xor U27726 (N_27726,N_26271,N_25466);
and U27727 (N_27727,N_25347,N_26210);
nor U27728 (N_27728,N_26678,N_25771);
nor U27729 (N_27729,N_26821,N_26302);
and U27730 (N_27730,N_25734,N_25454);
or U27731 (N_27731,N_27430,N_25645);
or U27732 (N_27732,N_25852,N_27429);
or U27733 (N_27733,N_26460,N_25168);
nor U27734 (N_27734,N_26406,N_25231);
or U27735 (N_27735,N_26940,N_27483);
and U27736 (N_27736,N_25403,N_25921);
nand U27737 (N_27737,N_25622,N_25444);
xnor U27738 (N_27738,N_25733,N_27283);
nand U27739 (N_27739,N_25484,N_25798);
xnor U27740 (N_27740,N_26500,N_26810);
and U27741 (N_27741,N_26308,N_26449);
and U27742 (N_27742,N_26072,N_26597);
nor U27743 (N_27743,N_25992,N_25677);
and U27744 (N_27744,N_26005,N_27285);
and U27745 (N_27745,N_25552,N_25746);
xor U27746 (N_27746,N_27498,N_27186);
and U27747 (N_27747,N_27348,N_26618);
xor U27748 (N_27748,N_26750,N_26888);
and U27749 (N_27749,N_25247,N_25832);
nor U27750 (N_27750,N_26093,N_26321);
or U27751 (N_27751,N_26186,N_25099);
and U27752 (N_27752,N_25065,N_25440);
nand U27753 (N_27753,N_25752,N_26795);
or U27754 (N_27754,N_26540,N_25555);
nand U27755 (N_27755,N_25427,N_26174);
nand U27756 (N_27756,N_26120,N_26628);
xor U27757 (N_27757,N_27439,N_25672);
nand U27758 (N_27758,N_25179,N_26808);
or U27759 (N_27759,N_26298,N_25865);
nor U27760 (N_27760,N_27440,N_25311);
nand U27761 (N_27761,N_26916,N_26796);
nor U27762 (N_27762,N_25082,N_25550);
xnor U27763 (N_27763,N_27103,N_25763);
or U27764 (N_27764,N_25595,N_26669);
xnor U27765 (N_27765,N_27204,N_27471);
nand U27766 (N_27766,N_25842,N_26704);
nor U27767 (N_27767,N_27111,N_26685);
or U27768 (N_27768,N_26476,N_26380);
or U27769 (N_27769,N_25876,N_27164);
xnor U27770 (N_27770,N_25605,N_26422);
nor U27771 (N_27771,N_26557,N_25587);
and U27772 (N_27772,N_25546,N_26690);
and U27773 (N_27773,N_25208,N_25571);
and U27774 (N_27774,N_27461,N_27094);
and U27775 (N_27775,N_25486,N_25840);
or U27776 (N_27776,N_25380,N_26399);
or U27777 (N_27777,N_27413,N_25644);
or U27778 (N_27778,N_26307,N_25103);
nand U27779 (N_27779,N_25094,N_26727);
and U27780 (N_27780,N_27087,N_25616);
nand U27781 (N_27781,N_26104,N_25391);
and U27782 (N_27782,N_25031,N_26691);
and U27783 (N_27783,N_26148,N_26518);
nand U27784 (N_27784,N_26194,N_27176);
and U27785 (N_27785,N_26742,N_25093);
xnor U27786 (N_27786,N_26679,N_26682);
and U27787 (N_27787,N_25212,N_27080);
xor U27788 (N_27788,N_27184,N_25202);
nand U27789 (N_27789,N_25575,N_26315);
xnor U27790 (N_27790,N_25875,N_26740);
nand U27791 (N_27791,N_25660,N_25230);
nor U27792 (N_27792,N_25336,N_26102);
or U27793 (N_27793,N_27437,N_25043);
and U27794 (N_27794,N_26028,N_26523);
xnor U27795 (N_27795,N_25063,N_25321);
nand U27796 (N_27796,N_26285,N_27141);
nor U27797 (N_27797,N_26774,N_26567);
nor U27798 (N_27798,N_25038,N_27153);
xor U27799 (N_27799,N_26985,N_26767);
xor U27800 (N_27800,N_26641,N_25790);
nand U27801 (N_27801,N_27262,N_26358);
and U27802 (N_27802,N_25161,N_26228);
or U27803 (N_27803,N_27419,N_26168);
nand U27804 (N_27804,N_25066,N_26840);
and U27805 (N_27805,N_26893,N_26884);
nand U27806 (N_27806,N_25143,N_26286);
nor U27807 (N_27807,N_25657,N_27320);
nand U27808 (N_27808,N_25461,N_26463);
nor U27809 (N_27809,N_26214,N_25131);
nor U27810 (N_27810,N_25956,N_25538);
nand U27811 (N_27811,N_26054,N_26580);
xor U27812 (N_27812,N_26684,N_25299);
and U27813 (N_27813,N_27252,N_26415);
nor U27814 (N_27814,N_25976,N_25123);
nand U27815 (N_27815,N_26544,N_27268);
xnor U27816 (N_27816,N_27315,N_26419);
nand U27817 (N_27817,N_25778,N_25457);
nor U27818 (N_27818,N_25590,N_25953);
and U27819 (N_27819,N_26366,N_26197);
nor U27820 (N_27820,N_27452,N_27114);
xor U27821 (N_27821,N_26002,N_25117);
nor U27822 (N_27822,N_26229,N_26489);
xor U27823 (N_27823,N_27386,N_27157);
xor U27824 (N_27824,N_25057,N_26462);
nand U27825 (N_27825,N_26639,N_26973);
or U27826 (N_27826,N_27280,N_25234);
xnor U27827 (N_27827,N_26839,N_26898);
or U27828 (N_27828,N_25869,N_26473);
nand U27829 (N_27829,N_25864,N_26428);
and U27830 (N_27830,N_25906,N_26923);
nand U27831 (N_27831,N_25088,N_27146);
nor U27832 (N_27832,N_25916,N_25700);
nor U27833 (N_27833,N_26891,N_25310);
xor U27834 (N_27834,N_27261,N_26133);
nand U27835 (N_27835,N_27212,N_26631);
nor U27836 (N_27836,N_26722,N_26070);
nor U27837 (N_27837,N_26847,N_25307);
or U27838 (N_27838,N_26574,N_25653);
nor U27839 (N_27839,N_27121,N_25167);
nand U27840 (N_27840,N_25426,N_26689);
and U27841 (N_27841,N_25954,N_26932);
and U27842 (N_27842,N_26340,N_26913);
nor U27843 (N_27843,N_26009,N_26693);
xor U27844 (N_27844,N_25994,N_25515);
nor U27845 (N_27845,N_26056,N_26115);
xnor U27846 (N_27846,N_25238,N_25301);
and U27847 (N_27847,N_27460,N_26746);
or U27848 (N_27848,N_26728,N_27323);
and U27849 (N_27849,N_25023,N_25786);
nand U27850 (N_27850,N_25608,N_26211);
nand U27851 (N_27851,N_25416,N_26881);
or U27852 (N_27852,N_26078,N_26646);
nand U27853 (N_27853,N_26977,N_26536);
nand U27854 (N_27854,N_26404,N_26894);
xor U27855 (N_27855,N_25157,N_26051);
nand U27856 (N_27856,N_27292,N_27425);
xor U27857 (N_27857,N_26342,N_26309);
xor U27858 (N_27858,N_26471,N_25603);
or U27859 (N_27859,N_26073,N_26303);
xor U27860 (N_27860,N_25825,N_26875);
nor U27861 (N_27861,N_25588,N_26766);
nor U27862 (N_27862,N_27484,N_26040);
or U27863 (N_27863,N_26861,N_27045);
xor U27864 (N_27864,N_25362,N_25937);
or U27865 (N_27865,N_27120,N_26582);
or U27866 (N_27866,N_27162,N_26249);
nor U27867 (N_27867,N_25977,N_27392);
or U27868 (N_27868,N_25521,N_27126);
and U27869 (N_27869,N_26836,N_26095);
nand U27870 (N_27870,N_26215,N_26508);
or U27871 (N_27871,N_27174,N_25799);
and U27872 (N_27872,N_25987,N_26956);
xnor U27873 (N_27873,N_27472,N_26658);
or U27874 (N_27874,N_27289,N_25715);
xnor U27875 (N_27875,N_27102,N_25780);
nor U27876 (N_27876,N_25562,N_26150);
nand U27877 (N_27877,N_27352,N_26998);
nand U27878 (N_27878,N_26562,N_26494);
nand U27879 (N_27879,N_26367,N_27286);
nand U27880 (N_27880,N_25545,N_27277);
xnor U27881 (N_27881,N_26395,N_25183);
nand U27882 (N_27882,N_26087,N_25279);
nor U27883 (N_27883,N_26725,N_25455);
nor U27884 (N_27884,N_26843,N_26573);
and U27885 (N_27885,N_25485,N_26496);
or U27886 (N_27886,N_26510,N_26757);
nand U27887 (N_27887,N_26699,N_26272);
and U27888 (N_27888,N_26092,N_26859);
nor U27889 (N_27889,N_26023,N_25000);
xnor U27890 (N_27890,N_27132,N_26779);
or U27891 (N_27891,N_26525,N_26619);
xor U27892 (N_27892,N_25422,N_26667);
xnor U27893 (N_27893,N_25511,N_26997);
and U27894 (N_27894,N_25643,N_25939);
and U27895 (N_27895,N_25271,N_25049);
nor U27896 (N_27896,N_26988,N_26933);
or U27897 (N_27897,N_25894,N_26887);
or U27898 (N_27898,N_26736,N_26252);
nand U27899 (N_27899,N_25765,N_26497);
nand U27900 (N_27900,N_27115,N_25565);
and U27901 (N_27901,N_27359,N_26506);
nor U27902 (N_27902,N_27407,N_25172);
and U27903 (N_27903,N_25563,N_25487);
and U27904 (N_27904,N_26981,N_26650);
and U27905 (N_27905,N_27044,N_26762);
and U27906 (N_27906,N_26674,N_26786);
or U27907 (N_27907,N_25263,N_25017);
or U27908 (N_27908,N_26820,N_25634);
and U27909 (N_27909,N_25762,N_26747);
nor U27910 (N_27910,N_26374,N_25813);
and U27911 (N_27911,N_26027,N_25012);
xor U27912 (N_27912,N_27019,N_26593);
nor U27913 (N_27913,N_26645,N_25612);
nand U27914 (N_27914,N_26436,N_26253);
nand U27915 (N_27915,N_26306,N_25943);
nor U27916 (N_27916,N_27034,N_25870);
and U27917 (N_27917,N_27227,N_26481);
xor U27918 (N_27918,N_26057,N_27067);
or U27919 (N_27919,N_26896,N_26091);
nor U27920 (N_27920,N_27274,N_26834);
nor U27921 (N_27921,N_25860,N_26015);
nor U27922 (N_27922,N_25624,N_26225);
and U27923 (N_27923,N_25205,N_26598);
and U27924 (N_27924,N_26236,N_26094);
and U27925 (N_27925,N_26457,N_26242);
xnor U27926 (N_27926,N_27092,N_26968);
nand U27927 (N_27927,N_26651,N_26131);
nand U27928 (N_27928,N_27343,N_25283);
nand U27929 (N_27929,N_25564,N_26668);
or U27930 (N_27930,N_26018,N_26433);
nand U27931 (N_27931,N_27077,N_25146);
nand U27932 (N_27932,N_25236,N_27420);
and U27933 (N_27933,N_27006,N_26672);
xnor U27934 (N_27934,N_27020,N_26902);
and U27935 (N_27935,N_26250,N_25028);
and U27936 (N_27936,N_27005,N_26318);
xor U27937 (N_27937,N_26310,N_26151);
or U27938 (N_27938,N_26400,N_25008);
or U27939 (N_27939,N_27042,N_26431);
and U27940 (N_27940,N_26798,N_27182);
and U27941 (N_27941,N_25072,N_25995);
nand U27942 (N_27942,N_27119,N_27444);
or U27943 (N_27943,N_26900,N_26857);
nor U27944 (N_27944,N_25759,N_27136);
nor U27945 (N_27945,N_25753,N_26987);
nor U27946 (N_27946,N_26080,N_25796);
nand U27947 (N_27947,N_25446,N_27128);
xnor U27948 (N_27948,N_26944,N_26856);
or U27949 (N_27949,N_27100,N_25874);
nand U27950 (N_27950,N_25489,N_27259);
nor U27951 (N_27951,N_26814,N_26206);
xnor U27952 (N_27952,N_25108,N_25229);
xor U27953 (N_27953,N_25144,N_25128);
or U27954 (N_27954,N_25908,N_26361);
nand U27955 (N_27955,N_25245,N_26384);
and U27956 (N_27956,N_25500,N_25419);
nor U27957 (N_27957,N_25879,N_27365);
or U27958 (N_27958,N_25553,N_27159);
nand U27959 (N_27959,N_26238,N_27187);
and U27960 (N_27960,N_26017,N_25365);
or U27961 (N_27961,N_26135,N_26753);
nand U27962 (N_27962,N_27394,N_27458);
or U27963 (N_27963,N_26130,N_27455);
and U27964 (N_27964,N_27282,N_25706);
xor U27965 (N_27965,N_25166,N_26291);
xnor U27966 (N_27966,N_26034,N_26613);
nand U27967 (N_27967,N_26756,N_26259);
nor U27968 (N_27968,N_25022,N_25986);
or U27969 (N_27969,N_25142,N_25175);
or U27970 (N_27970,N_26735,N_25070);
xor U27971 (N_27971,N_25496,N_26600);
xnor U27972 (N_27972,N_25926,N_26192);
and U27973 (N_27973,N_25421,N_27015);
or U27974 (N_27974,N_25626,N_26076);
or U27975 (N_27975,N_25784,N_27065);
nor U27976 (N_27976,N_26427,N_27393);
nor U27977 (N_27977,N_27306,N_25192);
nor U27978 (N_27978,N_26515,N_25100);
xnor U27979 (N_27979,N_26951,N_25258);
nand U27980 (N_27980,N_25291,N_25817);
nor U27981 (N_27981,N_27434,N_26890);
xor U27982 (N_27982,N_26749,N_25507);
nand U27983 (N_27983,N_25679,N_26853);
xor U27984 (N_27984,N_26443,N_27145);
xor U27985 (N_27985,N_27229,N_26845);
nand U27986 (N_27986,N_26219,N_27288);
nor U27987 (N_27987,N_26485,N_26181);
xnor U27988 (N_27988,N_26180,N_26348);
nor U27989 (N_27989,N_25159,N_26156);
nand U27990 (N_27990,N_25517,N_25829);
or U27991 (N_27991,N_25712,N_26455);
nand U27992 (N_27992,N_26616,N_27481);
or U27993 (N_27993,N_25631,N_25395);
xor U27994 (N_27994,N_26137,N_27081);
nand U27995 (N_27995,N_25589,N_27032);
nand U27996 (N_27996,N_25833,N_26324);
nand U27997 (N_27997,N_27368,N_27046);
xnor U27998 (N_27998,N_26972,N_25308);
xnor U27999 (N_27999,N_25348,N_27371);
nand U28000 (N_28000,N_27399,N_25714);
nor U28001 (N_28001,N_25736,N_26346);
nor U28002 (N_28002,N_27064,N_25206);
xor U28003 (N_28003,N_25689,N_26829);
nor U28004 (N_28004,N_26416,N_25738);
or U28005 (N_28005,N_25540,N_27294);
xor U28006 (N_28006,N_27169,N_26125);
or U28007 (N_28007,N_27462,N_25808);
nor U28008 (N_28008,N_27293,N_25145);
or U28009 (N_28009,N_25615,N_27197);
xnor U28010 (N_28010,N_25053,N_25647);
or U28011 (N_28011,N_25303,N_25477);
nor U28012 (N_28012,N_25010,N_25685);
nand U28013 (N_28013,N_25078,N_25429);
xnor U28014 (N_28014,N_25266,N_26869);
nor U28015 (N_28015,N_27108,N_25501);
xnor U28016 (N_28016,N_26470,N_26964);
and U28017 (N_28017,N_26244,N_25051);
and U28018 (N_28018,N_26714,N_27026);
and U28019 (N_28019,N_26633,N_26339);
xnor U28020 (N_28020,N_27470,N_25726);
xor U28021 (N_28021,N_27037,N_25020);
nor U28022 (N_28022,N_26293,N_26061);
nand U28023 (N_28023,N_25095,N_26989);
and U28024 (N_28024,N_25999,N_26016);
or U28025 (N_28025,N_25532,N_27245);
or U28026 (N_28026,N_27329,N_25913);
nand U28027 (N_28027,N_26524,N_25173);
nand U28028 (N_28028,N_27057,N_25343);
nand U28029 (N_28029,N_25030,N_26671);
nand U28030 (N_28030,N_27193,N_26110);
or U28031 (N_28031,N_25583,N_26644);
or U28032 (N_28032,N_25425,N_25407);
and U28033 (N_28033,N_25290,N_25872);
and U28034 (N_28034,N_26201,N_26490);
xor U28035 (N_28035,N_25339,N_25371);
xor U28036 (N_28036,N_26256,N_26982);
and U28037 (N_28037,N_25035,N_25324);
nand U28038 (N_28038,N_26364,N_25329);
nand U28039 (N_28039,N_26842,N_27486);
nor U28040 (N_28040,N_25558,N_26630);
or U28041 (N_28041,N_25188,N_25579);
and U28042 (N_28042,N_27260,N_26245);
nor U28043 (N_28043,N_26434,N_26136);
nor U28044 (N_28044,N_26203,N_27354);
xnor U28045 (N_28045,N_27168,N_27442);
nand U28046 (N_28046,N_25770,N_26615);
nor U28047 (N_28047,N_25936,N_25853);
xor U28048 (N_28048,N_25633,N_26677);
nand U28049 (N_28049,N_26218,N_26281);
or U28050 (N_28050,N_25621,N_26353);
and U28051 (N_28051,N_25274,N_25223);
nand U28052 (N_28052,N_25495,N_26037);
or U28053 (N_28053,N_27474,N_26383);
nor U28054 (N_28054,N_27055,N_25190);
and U28055 (N_28055,N_26806,N_26871);
xor U28056 (N_28056,N_26441,N_26701);
nor U28057 (N_28057,N_27383,N_26589);
and U28058 (N_28058,N_25899,N_27050);
nor U28059 (N_28059,N_25809,N_26267);
nand U28060 (N_28060,N_26610,N_25476);
and U28061 (N_28061,N_26408,N_26410);
or U28062 (N_28062,N_25265,N_26696);
nand U28063 (N_28063,N_25196,N_27305);
nor U28064 (N_28064,N_25332,N_26623);
and U28065 (N_28065,N_25990,N_25272);
xnor U28066 (N_28066,N_26474,N_26915);
or U28067 (N_28067,N_26442,N_26841);
and U28068 (N_28068,N_25749,N_27499);
nand U28069 (N_28069,N_25640,N_25949);
xnor U28070 (N_28070,N_26418,N_27195);
nand U28071 (N_28071,N_26152,N_27091);
nor U28072 (N_28072,N_25333,N_25988);
or U28073 (N_28073,N_25777,N_25417);
nand U28074 (N_28074,N_25855,N_26336);
and U28075 (N_28075,N_25508,N_25751);
xor U28076 (N_28076,N_25572,N_25334);
or U28077 (N_28077,N_27101,N_26179);
nor U28078 (N_28078,N_25233,N_25294);
or U28079 (N_28079,N_26835,N_26546);
or U28080 (N_28080,N_26119,N_26912);
or U28081 (N_28081,N_26118,N_27110);
and U28082 (N_28082,N_25635,N_26257);
nand U28083 (N_28083,N_25885,N_25408);
or U28084 (N_28084,N_26453,N_25978);
nor U28085 (N_28085,N_27248,N_27082);
xor U28086 (N_28086,N_27066,N_26526);
xor U28087 (N_28087,N_26069,N_25092);
or U28088 (N_28088,N_25409,N_26554);
and U28089 (N_28089,N_27328,N_27396);
and U28090 (N_28090,N_27109,N_26775);
nor U28091 (N_28091,N_25845,N_27265);
or U28092 (N_28092,N_26652,N_25973);
xnor U28093 (N_28093,N_26013,N_25002);
nand U28094 (N_28094,N_26886,N_26169);
nor U28095 (N_28095,N_26969,N_26343);
or U28096 (N_28096,N_26486,N_25319);
and U28097 (N_28097,N_26446,N_26105);
nand U28098 (N_28098,N_26885,N_26665);
nor U28099 (N_28099,N_25027,N_26648);
nor U28100 (N_28100,N_25122,N_25646);
and U28101 (N_28101,N_26659,N_25316);
and U28102 (N_28102,N_26548,N_25133);
and U28103 (N_28103,N_26263,N_25184);
and U28104 (N_28104,N_27191,N_27482);
nand U28105 (N_28105,N_26217,N_26469);
nand U28106 (N_28106,N_25152,N_25648);
xor U28107 (N_28107,N_25215,N_25102);
nor U28108 (N_28108,N_26421,N_26172);
nor U28109 (N_28109,N_26566,N_26647);
or U28110 (N_28110,N_25379,N_26527);
nor U28111 (N_28111,N_25984,N_25060);
nand U28112 (N_28112,N_26594,N_25016);
xor U28113 (N_28113,N_25084,N_27002);
xor U28114 (N_28114,N_26697,N_25456);
nor U28115 (N_28115,N_25449,N_25991);
nor U28116 (N_28116,N_26978,N_27269);
and U28117 (N_28117,N_27001,N_25354);
nor U28118 (N_28118,N_25367,N_26687);
or U28119 (N_28119,N_27070,N_25243);
xnor U28120 (N_28120,N_26590,N_26334);
or U28121 (N_28121,N_25998,N_25182);
or U28122 (N_28122,N_27158,N_26141);
nor U28123 (N_28123,N_26892,N_27116);
xnor U28124 (N_28124,N_26955,N_25839);
xnor U28125 (N_28125,N_26534,N_26394);
nand U28126 (N_28126,N_25582,N_25985);
xor U28127 (N_28127,N_25915,N_27417);
nor U28128 (N_28128,N_26246,N_27465);
xor U28129 (N_28129,N_26039,N_26388);
xnor U28130 (N_28130,N_26805,N_26780);
xnor U28131 (N_28131,N_25326,N_27373);
xor U28132 (N_28132,N_25493,N_25447);
and U28133 (N_28133,N_26723,N_26790);
and U28134 (N_28134,N_26055,N_26113);
or U28135 (N_28135,N_25216,N_26220);
xnor U28136 (N_28136,N_26530,N_25551);
nor U28137 (N_28137,N_26538,N_25080);
nand U28138 (N_28138,N_25004,N_26200);
xnor U28139 (N_28139,N_25747,N_25935);
or U28140 (N_28140,N_26583,N_27361);
nand U28141 (N_28141,N_25800,N_25069);
xnor U28142 (N_28142,N_27031,N_25067);
nor U28143 (N_28143,N_26241,N_25816);
and U28144 (N_28144,N_26850,N_25919);
nand U28145 (N_28145,N_26719,N_25887);
nor U28146 (N_28146,N_27339,N_26878);
nor U28147 (N_28147,N_26732,N_25704);
xor U28148 (N_28148,N_26049,N_26014);
xnor U28149 (N_28149,N_26895,N_25481);
xnor U28150 (N_28150,N_25652,N_26085);
nor U28151 (N_28151,N_27068,N_27161);
or U28152 (N_28152,N_25917,N_25090);
nand U28153 (N_28153,N_25420,N_27167);
xor U28154 (N_28154,N_26819,N_25527);
and U28155 (N_28155,N_25698,N_27448);
nor U28156 (N_28156,N_26031,N_27163);
nand U28157 (N_28157,N_26454,N_27362);
and U28158 (N_28158,N_27246,N_27071);
and U28159 (N_28159,N_26036,N_25934);
and U28160 (N_28160,N_26638,N_26811);
and U28161 (N_28161,N_27072,N_25941);
xnor U28162 (N_28162,N_26254,N_25101);
and U28163 (N_28163,N_25754,N_25598);
nand U28164 (N_28164,N_27056,N_25516);
xnor U28165 (N_28165,N_25021,N_25531);
and U28166 (N_28166,N_25232,N_25970);
and U28167 (N_28167,N_26067,N_25054);
or U28168 (N_28168,N_25764,N_25609);
and U28169 (N_28169,N_27030,N_27287);
or U28170 (N_28170,N_27228,N_25441);
nand U28171 (N_28171,N_27171,N_25381);
nand U28172 (N_28172,N_26661,N_27029);
nand U28173 (N_28173,N_26999,N_25656);
or U28174 (N_28174,N_27150,N_25774);
nor U28175 (N_28175,N_26331,N_25359);
and U28176 (N_28176,N_25376,N_27180);
nor U28177 (N_28177,N_25801,N_26273);
nand U28178 (N_28178,N_25886,N_25649);
nor U28179 (N_28179,N_26323,N_27196);
nor U28180 (N_28180,N_26042,N_27398);
xor U28181 (N_28181,N_26620,N_26287);
nand U28182 (N_28182,N_25826,N_26585);
nand U28183 (N_28183,N_25171,N_27370);
or U28184 (N_28184,N_27342,N_25533);
xor U28185 (N_28185,N_25641,N_25439);
nor U28186 (N_28186,N_26175,N_27401);
or U28187 (N_28187,N_26185,N_27205);
and U28188 (N_28188,N_25344,N_26581);
or U28189 (N_28189,N_27495,N_25828);
or U28190 (N_28190,N_25473,N_25601);
or U28191 (N_28191,N_25561,N_25891);
and U28192 (N_28192,N_27473,N_27000);
nand U28193 (N_28193,N_26709,N_26980);
or U28194 (N_28194,N_26673,N_27016);
and U28195 (N_28195,N_27243,N_25227);
nor U28196 (N_28196,N_27321,N_27048);
xor U28197 (N_28197,N_26437,N_26502);
and U28198 (N_28198,N_25580,N_27284);
and U28199 (N_28199,N_25389,N_26025);
and U28200 (N_28200,N_25393,N_26138);
nand U28201 (N_28201,N_26971,N_25410);
nor U28202 (N_28202,N_27079,N_25617);
nor U28203 (N_28203,N_27480,N_27233);
xnor U28204 (N_28204,N_26962,N_26377);
nor U28205 (N_28205,N_25156,N_25676);
and U28206 (N_28206,N_25802,N_25276);
nor U28207 (N_28207,N_27242,N_25925);
xnor U28208 (N_28208,N_26686,N_25019);
and U28209 (N_28209,N_25729,N_25024);
nor U28210 (N_28210,N_25064,N_25620);
nand U28211 (N_28211,N_26785,N_25837);
nor U28212 (N_28212,N_26199,N_26362);
nor U28213 (N_28213,N_25570,N_25474);
nor U28214 (N_28214,N_26341,N_27369);
xnor U28215 (N_28215,N_26086,N_27166);
or U28216 (N_28216,N_25370,N_27211);
xor U28217 (N_28217,N_26059,N_27496);
xor U28218 (N_28218,N_26047,N_27257);
nor U28219 (N_28219,N_27450,N_26804);
nand U28220 (N_28220,N_25896,N_26759);
or U28221 (N_28221,N_25897,N_25548);
and U28222 (N_28222,N_25297,N_26154);
and U28223 (N_28223,N_26935,N_27475);
or U28224 (N_28224,N_27340,N_26134);
and U28225 (N_28225,N_26033,N_26876);
nand U28226 (N_28226,N_26807,N_25827);
nor U28227 (N_28227,N_27453,N_27428);
nor U28228 (N_28228,N_25911,N_25289);
nor U28229 (N_28229,N_25194,N_25566);
xnor U28230 (N_28230,N_26863,N_27104);
xnor U28231 (N_28231,N_26365,N_26195);
and U28232 (N_28232,N_25013,N_26386);
or U28233 (N_28233,N_26226,N_27010);
nand U28234 (N_28234,N_25669,N_27208);
or U28235 (N_28235,N_25373,N_25963);
xor U28236 (N_28236,N_25692,N_26098);
and U28237 (N_28237,N_27181,N_27017);
or U28238 (N_28238,N_25745,N_25792);
or U28239 (N_28239,N_25382,N_25355);
xnor U28240 (N_28240,N_26163,N_26409);
xor U28241 (N_28241,N_25850,N_27009);
nor U28242 (N_28242,N_26071,N_26838);
or U28243 (N_28243,N_27238,N_26182);
and U28244 (N_28244,N_25529,N_26290);
xnor U28245 (N_28245,N_26514,N_26848);
or U28246 (N_28246,N_26251,N_25981);
nand U28247 (N_28247,N_25488,N_27432);
xnor U28248 (N_28248,N_25535,N_26282);
nor U28249 (N_28249,N_25225,N_25349);
and U28250 (N_28250,N_27028,N_26966);
or U28251 (N_28251,N_25866,N_27147);
or U28252 (N_28252,N_26769,N_26313);
xnor U28253 (N_28253,N_27384,N_27255);
or U28254 (N_28254,N_27236,N_26979);
nand U28255 (N_28255,N_25785,N_25137);
nor U28256 (N_28256,N_26487,N_26196);
nand U28257 (N_28257,N_26622,N_26060);
and U28258 (N_28258,N_26943,N_25450);
nand U28259 (N_28259,N_25637,N_26255);
nor U28260 (N_28260,N_25037,N_25805);
nand U28261 (N_28261,N_25881,N_25851);
xnor U28262 (N_28262,N_25285,N_25463);
and U28263 (N_28263,N_25390,N_25569);
nor U28264 (N_28264,N_26751,N_25375);
or U28265 (N_28265,N_26356,N_26707);
nand U28266 (N_28266,N_27040,N_25492);
and U28267 (N_28267,N_25942,N_25042);
nor U28268 (N_28268,N_27117,N_26146);
and U28269 (N_28269,N_25361,N_25134);
and U28270 (N_28270,N_25220,N_27353);
or U28271 (N_28271,N_25369,N_26209);
xor U28272 (N_28272,N_26737,N_25033);
xnor U28273 (N_28273,N_26854,N_26846);
or U28274 (N_28274,N_25769,N_27438);
or U28275 (N_28275,N_25412,N_25702);
and U28276 (N_28276,N_27250,N_26653);
or U28277 (N_28277,N_25639,N_26626);
or U28278 (N_28278,N_25750,N_25665);
or U28279 (N_28279,N_27224,N_27188);
and U28280 (N_28280,N_25821,N_27468);
or U28281 (N_28281,N_26755,N_26787);
nand U28282 (N_28282,N_26202,N_26862);
and U28283 (N_28283,N_27402,N_26405);
xnor U28284 (N_28284,N_26276,N_26304);
nor U28285 (N_28285,N_25001,N_26908);
nand U28286 (N_28286,N_26337,N_25824);
nor U28287 (N_28287,N_25214,N_27273);
xnor U28288 (N_28288,N_26077,N_26535);
nor U28289 (N_28289,N_25636,N_25252);
and U28290 (N_28290,N_27319,N_26279);
nand U28291 (N_28291,N_26666,N_26007);
xor U28292 (N_28292,N_25604,N_25722);
nor U28293 (N_28293,N_25744,N_25522);
nand U28294 (N_28294,N_25284,N_27140);
nand U28295 (N_28295,N_27151,N_25902);
nor U28296 (N_28296,N_26556,N_27059);
xor U28297 (N_28297,N_26983,N_27113);
and U28298 (N_28298,N_27219,N_26198);
and U28299 (N_28299,N_25269,N_25823);
nor U28300 (N_28300,N_25323,N_26407);
and U28301 (N_28301,N_26280,N_27388);
nor U28302 (N_28302,N_25924,N_27327);
and U28303 (N_28303,N_25317,N_26776);
or U28304 (N_28304,N_25313,N_25997);
and U28305 (N_28305,N_26444,N_25300);
and U28306 (N_28306,N_26359,N_26870);
xor U28307 (N_28307,N_25026,N_25822);
nor U28308 (N_28308,N_25255,N_25151);
or U28309 (N_28309,N_26531,N_27497);
or U28310 (N_28310,N_25695,N_25606);
nor U28311 (N_28311,N_26617,N_26802);
or U28312 (N_28312,N_25490,N_26447);
nand U28313 (N_28313,N_26360,N_26860);
nand U28314 (N_28314,N_26475,N_26664);
and U28315 (N_28315,N_27311,N_25278);
or U28316 (N_28316,N_25351,N_25898);
and U28317 (N_28317,N_25138,N_25844);
nand U28318 (N_28318,N_25932,N_25728);
and U28319 (N_28319,N_25707,N_26799);
xor U28320 (N_28320,N_26112,N_25556);
xor U28321 (N_28321,N_25345,N_25411);
nor U28322 (N_28322,N_26058,N_27247);
xor U28323 (N_28323,N_26216,N_25293);
or U28324 (N_28324,N_27156,N_27003);
nand U28325 (N_28325,N_25971,N_26006);
xor U28326 (N_28326,N_27215,N_25262);
nor U28327 (N_28327,N_26155,N_27165);
nor U28328 (N_28328,N_25920,N_26420);
xnor U28329 (N_28329,N_25098,N_25979);
and U28330 (N_28330,N_26397,N_26889);
xnor U28331 (N_28331,N_25847,N_26614);
and U28332 (N_28332,N_26052,N_25794);
xnor U28333 (N_28333,N_26178,N_26954);
xor U28334 (N_28334,N_27375,N_26164);
nand U28335 (N_28335,N_26165,N_25270);
or U28336 (N_28336,N_26852,N_27154);
xnor U28337 (N_28337,N_27446,N_26166);
and U28338 (N_28338,N_26167,N_25757);
or U28339 (N_28339,N_25868,N_26716);
xor U28340 (N_28340,N_26587,N_26398);
nor U28341 (N_28341,N_26926,N_26509);
xor U28342 (N_28342,N_27266,N_27467);
nor U28343 (N_28343,N_25014,N_25549);
or U28344 (N_28344,N_26929,N_26711);
nor U28345 (N_28345,N_27178,N_27424);
nand U28346 (N_28346,N_26937,N_26488);
and U28347 (N_28347,N_27272,N_25226);
xnor U28348 (N_28348,N_25584,N_26635);
nand U28349 (N_28349,N_27097,N_27391);
or U28350 (N_28350,N_27418,N_27372);
xnor U28351 (N_28351,N_25180,N_25048);
or U28352 (N_28352,N_26401,N_26517);
xor U28353 (N_28353,N_27222,N_27084);
and U28354 (N_28354,N_26423,N_25720);
xor U28355 (N_28355,N_26760,N_26240);
nor U28356 (N_28356,N_25228,N_25831);
nor U28357 (N_28357,N_26816,N_25464);
nor U28358 (N_28358,N_26144,N_25034);
xor U28359 (N_28359,N_25187,N_26683);
nor U28360 (N_28360,N_26761,N_26961);
or U28361 (N_28361,N_25530,N_25198);
nand U28362 (N_28362,N_26379,N_26521);
or U28363 (N_28363,N_26763,N_26043);
nand U28364 (N_28364,N_25893,N_25264);
nand U28365 (N_28365,N_26801,N_27139);
or U28366 (N_28366,N_27443,N_27304);
and U28367 (N_28367,N_25578,N_27400);
nor U28368 (N_28368,N_27479,N_25244);
xor U28369 (N_28369,N_25155,N_25993);
and U28370 (N_28370,N_26789,N_27235);
nand U28371 (N_28371,N_27374,N_26003);
xor U28372 (N_28372,N_27490,N_27012);
xnor U28373 (N_28373,N_27358,N_26354);
xor U28374 (N_28374,N_25119,N_26528);
xor U28375 (N_28375,N_27387,N_26670);
xor U28376 (N_28376,N_25483,N_27303);
nand U28377 (N_28377,N_25096,N_25682);
nor U28378 (N_28378,N_25961,N_25423);
nor U28379 (N_28379,N_25674,N_26317);
nor U28380 (N_28380,N_26800,N_25242);
xnor U28381 (N_28381,N_26773,N_25623);
and U28382 (N_28382,N_25740,N_25132);
nor U28383 (N_28383,N_26596,N_26296);
nor U28384 (N_28384,N_25011,N_26230);
nand U28385 (N_28385,N_27312,N_26588);
xor U28386 (N_28386,N_26865,N_27264);
and U28387 (N_28387,N_26606,N_27426);
or U28388 (N_28388,N_26483,N_26831);
or U28389 (N_28389,N_25309,N_25386);
xnor U28390 (N_28390,N_26312,N_27183);
nor U28391 (N_28391,N_27225,N_25952);
xor U28392 (N_28392,N_25951,N_26565);
xnor U28393 (N_28393,N_25528,N_25074);
xor U28394 (N_28394,N_26549,N_26700);
nor U28395 (N_28395,N_25830,N_25755);
and U28396 (N_28396,N_27249,N_25292);
or U28397 (N_28397,N_27333,N_26258);
nand U28398 (N_28398,N_27144,N_26472);
and U28399 (N_28399,N_25006,N_26918);
and U28400 (N_28400,N_26771,N_25114);
or U28401 (N_28401,N_27316,N_26261);
nor U28402 (N_28402,N_25573,N_27347);
nor U28403 (N_28403,N_25318,N_25241);
nand U28404 (N_28404,N_26390,N_25322);
nand U28405 (N_28405,N_27447,N_26642);
nor U28406 (N_28406,N_25460,N_25611);
xor U28407 (N_28407,N_27160,N_26879);
nor U28408 (N_28408,N_26792,N_25628);
or U28409 (N_28409,N_25073,N_25678);
or U28410 (N_28410,N_26903,N_25224);
nor U28411 (N_28411,N_27367,N_27493);
nand U28412 (N_28412,N_26662,N_26601);
xor U28413 (N_28413,N_25586,N_25856);
and U28414 (N_28414,N_26482,N_25737);
or U28415 (N_28415,N_25596,N_27457);
xnor U28416 (N_28416,N_25451,N_26996);
and U28417 (N_28417,N_25003,N_26823);
nor U28418 (N_28418,N_26010,N_27076);
nor U28419 (N_28419,N_26084,N_26883);
nor U28420 (N_28420,N_27423,N_26301);
or U28421 (N_28421,N_25857,N_25415);
nand U28422 (N_28422,N_26702,N_27270);
nor U28423 (N_28423,N_26269,N_25710);
or U28424 (N_28424,N_25007,N_25374);
or U28425 (N_28425,N_25914,N_27356);
xnor U28426 (N_28426,N_27454,N_26068);
nand U28427 (N_28427,N_25807,N_26676);
and U28428 (N_28428,N_26822,N_25526);
nand U28429 (N_28429,N_25858,N_26770);
nand U28430 (N_28430,N_26809,N_26595);
xnor U28431 (N_28431,N_26425,N_27427);
and U28432 (N_28432,N_27107,N_26833);
nand U28433 (N_28433,N_25494,N_26764);
and U28434 (N_28434,N_26075,N_25257);
xnor U28435 (N_28435,N_26191,N_25520);
xnor U28436 (N_28436,N_25210,N_27307);
or U28437 (N_28437,N_25378,N_25201);
xor U28438 (N_28438,N_25204,N_25512);
or U28439 (N_28439,N_26451,N_25141);
nor U28440 (N_28440,N_25475,N_27335);
and U28441 (N_28441,N_25873,N_26815);
nand U28442 (N_28442,N_25768,N_26458);
nor U28443 (N_28443,N_26551,N_25200);
and U28444 (N_28444,N_25662,N_25811);
or U28445 (N_28445,N_25502,N_25996);
nand U28446 (N_28446,N_25980,N_25295);
nand U28447 (N_28447,N_26994,N_27149);
or U28448 (N_28448,N_25281,N_25040);
nor U28449 (N_28449,N_25688,N_25909);
xor U28450 (N_28450,N_25810,N_26116);
nor U28451 (N_28451,N_26569,N_26872);
nand U28452 (N_28452,N_25705,N_26501);
nor U28453 (N_28453,N_25537,N_27223);
nor U28454 (N_28454,N_27127,N_27025);
nor U28455 (N_28455,N_26243,N_25933);
or U28456 (N_28456,N_27314,N_25015);
or U28457 (N_28457,N_25741,N_25445);
and U28458 (N_28458,N_25912,N_25433);
xnor U28459 (N_28459,N_26429,N_26739);
xnor U28460 (N_28460,N_27326,N_26147);
nand U28461 (N_28461,N_25260,N_26858);
nor U28462 (N_28462,N_25288,N_26239);
xnor U28463 (N_28463,N_26637,N_26625);
xnor U28464 (N_28464,N_25029,N_26873);
nand U28465 (N_28465,N_26193,N_25505);
nand U28466 (N_28466,N_25482,N_25923);
xor U28467 (N_28467,N_26327,N_25470);
or U28468 (N_28468,N_26132,N_25363);
and U28469 (N_28469,N_26024,N_26053);
xnor U28470 (N_28470,N_25638,N_26706);
or U28471 (N_28471,N_25684,N_26967);
nor U28472 (N_28472,N_26316,N_26663);
nor U28473 (N_28473,N_25139,N_25818);
xnor U28474 (N_28474,N_26781,N_26830);
or U28475 (N_28475,N_26591,N_25089);
and U28476 (N_28476,N_25169,N_26717);
and U28477 (N_28477,N_26223,N_26827);
nor U28478 (N_28478,N_26745,N_25671);
nand U28479 (N_28479,N_26000,N_26347);
nand U28480 (N_28480,N_25109,N_25055);
xnor U28481 (N_28481,N_25972,N_26351);
nand U28482 (N_28482,N_25696,N_27349);
or U28483 (N_28483,N_26907,N_25723);
xnor U28484 (N_28484,N_25165,N_25478);
nand U28485 (N_28485,N_26371,N_25766);
nand U28486 (N_28486,N_27036,N_26575);
xor U28487 (N_28487,N_25239,N_25525);
xnor U28488 (N_28488,N_27230,N_25735);
nand U28489 (N_28489,N_27390,N_25113);
nand U28490 (N_28490,N_26604,N_27058);
or U28491 (N_28491,N_26768,N_26734);
or U28492 (N_28492,N_26909,N_25536);
nand U28493 (N_28493,N_25846,N_26744);
and U28494 (N_28494,N_26090,N_25713);
xnor U28495 (N_28495,N_27451,N_25218);
nand U28496 (N_28496,N_26930,N_25694);
and U28497 (N_28497,N_26088,N_26101);
xnor U28498 (N_28498,N_26965,N_25384);
xor U28499 (N_28499,N_26710,N_27302);
or U28500 (N_28500,N_26897,N_26974);
nor U28501 (N_28501,N_27172,N_26553);
or U28502 (N_28502,N_27237,N_26654);
xnor U28503 (N_28503,N_25880,N_26529);
and U28504 (N_28504,N_25120,N_27201);
or U28505 (N_28505,N_25126,N_26975);
nor U28506 (N_28506,N_25889,N_26694);
and U28507 (N_28507,N_27130,N_26656);
or U28508 (N_28508,N_25591,N_26609);
nor U28509 (N_28509,N_25910,N_26158);
xnor U28510 (N_28510,N_26919,N_26126);
and U28511 (N_28511,N_26183,N_26511);
xor U28512 (N_28512,N_26373,N_26579);
nand U28513 (N_28513,N_27192,N_26602);
and U28514 (N_28514,N_27123,N_27035);
xor U28515 (N_28515,N_25506,N_26950);
or U28516 (N_28516,N_25610,N_26326);
nand U28517 (N_28517,N_25929,N_27152);
nand U28518 (N_28518,N_27488,N_25320);
xnor U28519 (N_28519,N_25105,N_27095);
or U28520 (N_28520,N_26855,N_26986);
xnor U28521 (N_28521,N_26928,N_25760);
or U28522 (N_28522,N_25697,N_26142);
xor U28523 (N_28523,N_26424,N_25328);
or U28524 (N_28524,N_26543,N_26533);
and U28525 (N_28525,N_25186,N_26171);
and U28526 (N_28526,N_27088,N_25581);
nand U28527 (N_28527,N_26948,N_26991);
or U28528 (N_28528,N_26491,N_27004);
nor U28529 (N_28529,N_27416,N_26288);
and U28530 (N_28530,N_25664,N_26958);
or U28531 (N_28531,N_26793,N_27135);
xnor U28532 (N_28532,N_26277,N_26921);
xor U28533 (N_28533,N_26778,N_27089);
nor U28534 (N_28534,N_26465,N_25217);
nor U28535 (N_28535,N_25574,N_26720);
nand U28536 (N_28536,N_26213,N_25602);
and U28537 (N_28537,N_26300,N_25725);
or U28538 (N_28538,N_26910,N_25221);
and U28539 (N_28539,N_26299,N_25795);
xor U28540 (N_28540,N_25397,N_27267);
nor U28541 (N_28541,N_26260,N_25767);
nor U28542 (N_28542,N_25197,N_26097);
or U28543 (N_28543,N_26330,N_27492);
nand U28544 (N_28544,N_25340,N_25189);
nor U28545 (N_28545,N_25797,N_27011);
or U28546 (N_28546,N_25982,N_25859);
or U28547 (N_28547,N_26880,N_26578);
and U28548 (N_28548,N_25056,N_26417);
or U28549 (N_28549,N_26559,N_25153);
xnor U28550 (N_28550,N_25585,N_27377);
nand U28551 (N_28551,N_25773,N_25250);
or U28552 (N_28552,N_25834,N_25959);
nand U28553 (N_28553,N_27033,N_26560);
nor U28554 (N_28554,N_26817,N_27053);
nor U28555 (N_28555,N_25071,N_25534);
xnor U28556 (N_28556,N_27403,N_27217);
nor U28557 (N_28557,N_25147,N_26153);
and U28558 (N_28558,N_27415,N_27360);
xor U28559 (N_28559,N_25772,N_26477);
or U28560 (N_28560,N_25687,N_25465);
nor U28561 (N_28561,N_26322,N_26403);
nor U28562 (N_28562,N_25352,N_26349);
nand U28563 (N_28563,N_26537,N_26161);
or U28564 (N_28564,N_27346,N_26901);
and U28565 (N_28565,N_26992,N_25600);
and U28566 (N_28566,N_26426,N_26503);
and U28567 (N_28567,N_25246,N_26173);
and U28568 (N_28568,N_27085,N_26122);
and U28569 (N_28569,N_25059,N_26100);
or U28570 (N_28570,N_26456,N_25989);
and U28571 (N_28571,N_25211,N_27441);
xnor U28572 (N_28572,N_26963,N_25812);
nor U28573 (N_28573,N_27309,N_25513);
or U28574 (N_28574,N_25112,N_27023);
nor U28575 (N_28575,N_26754,N_25174);
nand U28576 (N_28576,N_26381,N_25044);
xnor U28577 (N_28577,N_25366,N_25377);
or U28578 (N_28578,N_25287,N_25542);
nand U28579 (N_28579,N_26520,N_26278);
xor U28580 (N_28580,N_25435,N_27414);
or U28581 (N_28581,N_26675,N_25181);
nor U28582 (N_28582,N_25330,N_27216);
xor U28583 (N_28583,N_25703,N_26844);
or U28584 (N_28584,N_25524,N_27431);
nand U28585 (N_28585,N_27241,N_25659);
and U28586 (N_28586,N_26011,N_27405);
nand U28587 (N_28587,N_27240,N_26050);
or U28588 (N_28588,N_25353,N_26352);
xnor U28589 (N_28589,N_27350,N_27290);
and U28590 (N_28590,N_26695,N_27332);
nor U28591 (N_28591,N_25432,N_25966);
nor U28592 (N_28592,N_25405,N_26235);
nor U28593 (N_28593,N_26621,N_27275);
nor U28594 (N_28594,N_25803,N_26577);
xor U28595 (N_28595,N_26788,N_25356);
and U28596 (N_28596,N_27494,N_27190);
nor U28597 (N_28597,N_26008,N_26382);
xnor U28598 (N_28598,N_27054,N_26411);
xnor U28599 (N_28599,N_25130,N_26140);
nor U28600 (N_28600,N_25462,N_27073);
xor U28601 (N_28601,N_27148,N_26387);
or U28602 (N_28602,N_26945,N_26297);
or U28603 (N_28603,N_25491,N_27099);
xor U28604 (N_28604,N_25567,N_27408);
nor U28605 (N_28605,N_25058,N_25884);
and U28606 (N_28606,N_25836,N_26294);
nor U28607 (N_28607,N_25804,N_25400);
nand U28608 (N_28608,N_25306,N_25185);
and U28609 (N_28609,N_26332,N_25693);
and U28610 (N_28610,N_27129,N_25838);
xnor U28611 (N_28611,N_26450,N_26445);
nand U28612 (N_28612,N_26532,N_26629);
nand U28613 (N_28613,N_26825,N_26032);
or U28614 (N_28614,N_25061,N_26045);
xor U28615 (N_28615,N_25402,N_26048);
nor U28616 (N_28616,N_25681,N_27096);
nand U28617 (N_28617,N_25368,N_26837);
and U28618 (N_28618,N_26803,N_26990);
nor U28619 (N_28619,N_27258,N_27338);
and U28620 (N_28620,N_25437,N_26190);
nand U28621 (N_28621,N_26568,N_26649);
xor U28622 (N_28622,N_25748,N_25327);
xor U28623 (N_28623,N_26376,N_25783);
and U28624 (N_28624,N_25743,N_25731);
xnor U28625 (N_28625,N_26369,N_25670);
xnor U28626 (N_28626,N_26724,N_25118);
nand U28627 (N_28627,N_25467,N_27155);
nor U28628 (N_28628,N_25683,N_26128);
xor U28629 (N_28629,N_25642,N_25732);
nor U28630 (N_28630,N_26350,N_26335);
or U28631 (N_28631,N_25779,N_26391);
nor U28632 (N_28632,N_25176,N_25277);
nor U28633 (N_28633,N_25718,N_26692);
or U28634 (N_28634,N_26927,N_27410);
nand U28635 (N_28635,N_27317,N_26212);
or U28636 (N_28636,N_26824,N_26375);
and U28637 (N_28637,N_25619,N_26030);
nor U28638 (N_28638,N_25436,N_26338);
or U28639 (N_28639,N_26368,N_26275);
xor U28640 (N_28640,N_27062,N_25350);
nand U28641 (N_28641,N_27231,N_25267);
xor U28642 (N_28642,N_26264,N_27421);
or U28643 (N_28643,N_25673,N_27124);
xnor U28644 (N_28644,N_26758,N_25431);
xnor U28645 (N_28645,N_26325,N_25302);
nand U28646 (N_28646,N_26237,N_27074);
nor U28647 (N_28647,N_25613,N_25969);
xor U28648 (N_28648,N_26468,N_26941);
or U28649 (N_28649,N_26545,N_26022);
nand U28650 (N_28650,N_26718,N_25158);
nand U28651 (N_28651,N_26099,N_26177);
and U28652 (N_28652,N_25557,N_26145);
xnor U28653 (N_28653,N_25960,N_25599);
and U28654 (N_28654,N_25895,N_25730);
xnor U28655 (N_28655,N_26877,N_26947);
xor U28656 (N_28656,N_25974,N_27131);
and U28657 (N_28657,N_27422,N_26605);
and U28658 (N_28658,N_25497,N_25213);
or U28659 (N_28659,N_25861,N_25686);
and U28660 (N_28660,N_25788,N_26949);
nor U28661 (N_28661,N_26074,N_25076);
nor U28662 (N_28662,N_27179,N_27278);
or U28663 (N_28663,N_27206,N_27355);
and U28664 (N_28664,N_26106,N_25667);
nand U28665 (N_28665,N_27363,N_25298);
nand U28666 (N_28666,N_25975,N_26952);
nor U28667 (N_28667,N_25438,N_26934);
nor U28668 (N_28668,N_27251,N_27239);
xor U28669 (N_28669,N_25630,N_25191);
nand U28670 (N_28670,N_26355,N_25892);
and U28671 (N_28671,N_25962,N_26632);
and U28672 (N_28672,N_25097,N_26159);
and U28673 (N_28673,N_25675,N_26917);
or U28674 (N_28674,N_25782,N_25115);
and U28675 (N_28675,N_26247,N_26082);
xnor U28676 (N_28676,N_27351,N_25791);
xor U28677 (N_28677,N_26922,N_26262);
or U28678 (N_28678,N_27318,N_27106);
nand U28679 (N_28679,N_27466,N_27185);
nand U28680 (N_28680,N_27253,N_25928);
or U28681 (N_28681,N_27051,N_26184);
nand U28682 (N_28682,N_27090,N_25162);
nor U28683 (N_28683,N_26265,N_25775);
and U28684 (N_28684,N_26292,N_26205);
nor U28685 (N_28685,N_26611,N_26121);
and U28686 (N_28686,N_26570,N_27086);
and U28687 (N_28687,N_25442,N_26385);
nor U28688 (N_28688,N_26079,N_25607);
and U28689 (N_28689,N_25434,N_26270);
nand U28690 (N_28690,N_27478,N_27463);
and U28691 (N_28691,N_27198,N_27476);
nor U28692 (N_28692,N_27380,N_25296);
nand U28693 (N_28693,N_25414,N_27105);
xor U28694 (N_28694,N_26345,N_25539);
and U28695 (N_28695,N_25469,N_25009);
and U28696 (N_28696,N_27409,N_27209);
nand U28697 (N_28697,N_25280,N_26911);
or U28698 (N_28698,N_25399,N_26772);
nand U28699 (N_28699,N_27137,N_25964);
xnor U28700 (N_28700,N_25877,N_25523);
or U28701 (N_28701,N_25372,N_27093);
nand U28702 (N_28702,N_26370,N_26752);
xnor U28703 (N_28703,N_25110,N_26703);
or U28704 (N_28704,N_26466,N_26541);
nand U28705 (N_28705,N_25387,N_26295);
and U28706 (N_28706,N_27366,N_27491);
nor U28707 (N_28707,N_26233,N_25499);
nand U28708 (N_28708,N_26868,N_26107);
and U28709 (N_28709,N_27449,N_26942);
nor U28710 (N_28710,N_26221,N_26414);
or U28711 (N_28711,N_27324,N_26063);
and U28712 (N_28712,N_26655,N_26812);
nand U28713 (N_28713,N_25148,N_26046);
xnor U28714 (N_28714,N_27271,N_27334);
nor U28715 (N_28715,N_26783,N_25448);
nand U28716 (N_28716,N_25597,N_25947);
nand U28717 (N_28717,N_25690,N_26357);
or U28718 (N_28718,N_25385,N_26640);
or U28719 (N_28719,N_26599,N_27376);
or U28720 (N_28720,N_26970,N_27337);
or U28721 (N_28721,N_27220,N_26993);
nor U28722 (N_28722,N_27345,N_25632);
xor U28723 (N_28723,N_26109,N_26208);
nand U28724 (N_28724,N_26188,N_26499);
xnor U28725 (N_28725,N_25050,N_25472);
or U28726 (N_28726,N_26882,N_26448);
and U28727 (N_28727,N_25655,N_25618);
and U28728 (N_28728,N_25083,N_27469);
xor U28729 (N_28729,N_27389,N_25253);
and U28730 (N_28730,N_25835,N_27203);
xnor U28731 (N_28731,N_25160,N_26044);
nand U28732 (N_28732,N_27125,N_26995);
nand U28733 (N_28733,N_27047,N_27435);
nand U28734 (N_28734,N_25127,N_25388);
nand U28735 (N_28735,N_27295,N_26479);
xnor U28736 (N_28736,N_26504,N_25938);
and U28737 (N_28737,N_25062,N_26513);
or U28738 (N_28738,N_25401,N_25222);
nor U28739 (N_28739,N_26432,N_25140);
nand U28740 (N_28740,N_25315,N_26162);
or U28741 (N_28741,N_26081,N_27112);
nand U28742 (N_28742,N_25758,N_26920);
or U28743 (N_28743,N_26586,N_25820);
nor U28744 (N_28744,N_27379,N_26066);
nand U28745 (N_28745,N_26680,N_27456);
or U28746 (N_28746,N_27061,N_25883);
nor U28747 (N_28747,N_26539,N_26224);
xor U28748 (N_28748,N_25107,N_25256);
and U28749 (N_28749,N_25149,N_25259);
nor U28750 (N_28750,N_25108,N_25134);
xnor U28751 (N_28751,N_26320,N_26954);
or U28752 (N_28752,N_27375,N_25394);
and U28753 (N_28753,N_26354,N_25552);
xnor U28754 (N_28754,N_26034,N_25951);
nor U28755 (N_28755,N_26686,N_26127);
or U28756 (N_28756,N_25673,N_27455);
nand U28757 (N_28757,N_26134,N_27313);
nor U28758 (N_28758,N_27059,N_26382);
or U28759 (N_28759,N_25435,N_25385);
xor U28760 (N_28760,N_26139,N_26355);
nand U28761 (N_28761,N_26687,N_25678);
xor U28762 (N_28762,N_25876,N_27415);
or U28763 (N_28763,N_25815,N_25283);
or U28764 (N_28764,N_26679,N_26007);
nor U28765 (N_28765,N_25013,N_27401);
xnor U28766 (N_28766,N_26360,N_27166);
nand U28767 (N_28767,N_26746,N_26807);
nand U28768 (N_28768,N_26053,N_27144);
nor U28769 (N_28769,N_25426,N_26339);
nor U28770 (N_28770,N_27259,N_26342);
nand U28771 (N_28771,N_25073,N_27205);
and U28772 (N_28772,N_25288,N_25915);
xnor U28773 (N_28773,N_25414,N_27033);
nand U28774 (N_28774,N_26541,N_27063);
or U28775 (N_28775,N_26561,N_26170);
nor U28776 (N_28776,N_26578,N_25952);
nand U28777 (N_28777,N_27044,N_26016);
nor U28778 (N_28778,N_26581,N_26954);
nand U28779 (N_28779,N_26967,N_25376);
nor U28780 (N_28780,N_26788,N_26274);
xnor U28781 (N_28781,N_25910,N_25457);
nor U28782 (N_28782,N_26253,N_26211);
or U28783 (N_28783,N_26436,N_25276);
nand U28784 (N_28784,N_25479,N_25038);
nor U28785 (N_28785,N_26390,N_26353);
nor U28786 (N_28786,N_26456,N_27116);
xor U28787 (N_28787,N_25322,N_25349);
or U28788 (N_28788,N_26542,N_26425);
nand U28789 (N_28789,N_27218,N_26294);
or U28790 (N_28790,N_26767,N_26350);
xor U28791 (N_28791,N_26552,N_27117);
xnor U28792 (N_28792,N_25983,N_26371);
or U28793 (N_28793,N_25699,N_25015);
and U28794 (N_28794,N_25678,N_26072);
nand U28795 (N_28795,N_25655,N_25993);
nor U28796 (N_28796,N_26794,N_25164);
nand U28797 (N_28797,N_25565,N_27498);
xor U28798 (N_28798,N_25216,N_25774);
nor U28799 (N_28799,N_25008,N_25483);
or U28800 (N_28800,N_25527,N_26060);
and U28801 (N_28801,N_26483,N_25120);
nand U28802 (N_28802,N_26782,N_26645);
xor U28803 (N_28803,N_26614,N_25479);
nand U28804 (N_28804,N_27428,N_27031);
or U28805 (N_28805,N_27494,N_27042);
and U28806 (N_28806,N_26801,N_27145);
xnor U28807 (N_28807,N_26892,N_25375);
xnor U28808 (N_28808,N_25087,N_25950);
xnor U28809 (N_28809,N_25436,N_25778);
nand U28810 (N_28810,N_25104,N_27179);
nor U28811 (N_28811,N_26598,N_26080);
and U28812 (N_28812,N_26783,N_26773);
xor U28813 (N_28813,N_26560,N_25011);
nor U28814 (N_28814,N_25472,N_25879);
xor U28815 (N_28815,N_26779,N_25306);
or U28816 (N_28816,N_25919,N_26640);
nor U28817 (N_28817,N_27271,N_25398);
nand U28818 (N_28818,N_25909,N_25314);
and U28819 (N_28819,N_25934,N_27075);
xor U28820 (N_28820,N_25372,N_27483);
xnor U28821 (N_28821,N_25367,N_25138);
nor U28822 (N_28822,N_25839,N_25201);
or U28823 (N_28823,N_26639,N_26045);
nand U28824 (N_28824,N_26176,N_26610);
or U28825 (N_28825,N_27094,N_26829);
xor U28826 (N_28826,N_27084,N_27495);
nor U28827 (N_28827,N_26568,N_26085);
nand U28828 (N_28828,N_25595,N_26058);
xor U28829 (N_28829,N_25603,N_25253);
or U28830 (N_28830,N_27055,N_27012);
xor U28831 (N_28831,N_26592,N_25440);
nand U28832 (N_28832,N_26474,N_25475);
nor U28833 (N_28833,N_25081,N_26033);
and U28834 (N_28834,N_25386,N_26005);
xnor U28835 (N_28835,N_26000,N_25721);
xor U28836 (N_28836,N_27334,N_27342);
xnor U28837 (N_28837,N_27266,N_27454);
and U28838 (N_28838,N_25279,N_27153);
nand U28839 (N_28839,N_25067,N_25281);
xnor U28840 (N_28840,N_25172,N_25624);
and U28841 (N_28841,N_25263,N_26796);
nor U28842 (N_28842,N_26320,N_25782);
nor U28843 (N_28843,N_25537,N_25973);
nor U28844 (N_28844,N_26477,N_25253);
xnor U28845 (N_28845,N_25275,N_26092);
nand U28846 (N_28846,N_27123,N_26822);
and U28847 (N_28847,N_27171,N_25203);
xor U28848 (N_28848,N_27449,N_26300);
xnor U28849 (N_28849,N_26414,N_25401);
and U28850 (N_28850,N_26651,N_26309);
and U28851 (N_28851,N_27279,N_27299);
nand U28852 (N_28852,N_25920,N_26394);
or U28853 (N_28853,N_25626,N_27439);
xnor U28854 (N_28854,N_27435,N_25007);
and U28855 (N_28855,N_27144,N_26068);
and U28856 (N_28856,N_25921,N_26091);
or U28857 (N_28857,N_27213,N_26595);
nand U28858 (N_28858,N_25619,N_25418);
nor U28859 (N_28859,N_25559,N_26551);
nor U28860 (N_28860,N_27295,N_26586);
and U28861 (N_28861,N_25084,N_25923);
or U28862 (N_28862,N_25343,N_25267);
or U28863 (N_28863,N_27227,N_25766);
and U28864 (N_28864,N_25295,N_25415);
nor U28865 (N_28865,N_26738,N_25588);
and U28866 (N_28866,N_25909,N_26863);
nor U28867 (N_28867,N_25768,N_27293);
nor U28868 (N_28868,N_25500,N_26692);
or U28869 (N_28869,N_25221,N_26629);
or U28870 (N_28870,N_27323,N_26842);
nand U28871 (N_28871,N_26762,N_25648);
or U28872 (N_28872,N_25511,N_25111);
xnor U28873 (N_28873,N_26723,N_27453);
and U28874 (N_28874,N_25335,N_26867);
and U28875 (N_28875,N_25397,N_25759);
or U28876 (N_28876,N_26837,N_26158);
nand U28877 (N_28877,N_26693,N_25737);
nor U28878 (N_28878,N_26411,N_26919);
nand U28879 (N_28879,N_26609,N_26802);
nand U28880 (N_28880,N_27273,N_25211);
xor U28881 (N_28881,N_26330,N_25042);
or U28882 (N_28882,N_25277,N_25743);
nor U28883 (N_28883,N_27220,N_26711);
nand U28884 (N_28884,N_27491,N_25633);
and U28885 (N_28885,N_25828,N_25465);
and U28886 (N_28886,N_25618,N_25766);
xor U28887 (N_28887,N_26862,N_26871);
xor U28888 (N_28888,N_26503,N_25982);
nor U28889 (N_28889,N_25505,N_26679);
or U28890 (N_28890,N_27440,N_25663);
and U28891 (N_28891,N_26577,N_26372);
nand U28892 (N_28892,N_25015,N_27051);
or U28893 (N_28893,N_25757,N_25420);
nor U28894 (N_28894,N_25101,N_25304);
or U28895 (N_28895,N_26346,N_25055);
nor U28896 (N_28896,N_25825,N_25757);
xor U28897 (N_28897,N_26146,N_25846);
and U28898 (N_28898,N_25608,N_25863);
and U28899 (N_28899,N_25118,N_26893);
xor U28900 (N_28900,N_26014,N_26257);
or U28901 (N_28901,N_26580,N_26318);
nand U28902 (N_28902,N_26902,N_26216);
nor U28903 (N_28903,N_26357,N_26004);
or U28904 (N_28904,N_26665,N_25191);
and U28905 (N_28905,N_27049,N_26274);
or U28906 (N_28906,N_26837,N_26966);
and U28907 (N_28907,N_25845,N_26392);
xor U28908 (N_28908,N_27037,N_26077);
nand U28909 (N_28909,N_25013,N_26146);
xnor U28910 (N_28910,N_25972,N_26173);
and U28911 (N_28911,N_26959,N_25801);
nor U28912 (N_28912,N_26552,N_26835);
nand U28913 (N_28913,N_25350,N_25706);
nor U28914 (N_28914,N_27320,N_27213);
nor U28915 (N_28915,N_26622,N_26571);
nor U28916 (N_28916,N_27076,N_26110);
or U28917 (N_28917,N_26555,N_25456);
nor U28918 (N_28918,N_25651,N_25092);
or U28919 (N_28919,N_27455,N_27016);
xor U28920 (N_28920,N_27373,N_26576);
or U28921 (N_28921,N_26006,N_26667);
and U28922 (N_28922,N_25452,N_26955);
or U28923 (N_28923,N_25955,N_26329);
nor U28924 (N_28924,N_25721,N_26623);
xnor U28925 (N_28925,N_26403,N_27009);
nand U28926 (N_28926,N_25382,N_25768);
nor U28927 (N_28927,N_25990,N_27052);
nand U28928 (N_28928,N_27343,N_25585);
or U28929 (N_28929,N_27330,N_26414);
or U28930 (N_28930,N_25870,N_26715);
and U28931 (N_28931,N_27319,N_26510);
xor U28932 (N_28932,N_25757,N_25154);
nand U28933 (N_28933,N_26017,N_26771);
nand U28934 (N_28934,N_27021,N_26798);
or U28935 (N_28935,N_25508,N_25761);
nor U28936 (N_28936,N_25441,N_25067);
or U28937 (N_28937,N_25150,N_25551);
and U28938 (N_28938,N_26245,N_26292);
nor U28939 (N_28939,N_25225,N_27350);
and U28940 (N_28940,N_25548,N_25815);
or U28941 (N_28941,N_26821,N_25447);
or U28942 (N_28942,N_25770,N_25443);
xnor U28943 (N_28943,N_26905,N_27279);
nor U28944 (N_28944,N_26448,N_25823);
xor U28945 (N_28945,N_26968,N_25228);
and U28946 (N_28946,N_25979,N_25248);
xor U28947 (N_28947,N_26651,N_26004);
nor U28948 (N_28948,N_26620,N_26954);
or U28949 (N_28949,N_25932,N_26897);
or U28950 (N_28950,N_27054,N_26374);
and U28951 (N_28951,N_26840,N_26090);
or U28952 (N_28952,N_26925,N_25679);
or U28953 (N_28953,N_27036,N_26178);
nand U28954 (N_28954,N_26008,N_25518);
nand U28955 (N_28955,N_27207,N_26217);
nor U28956 (N_28956,N_25418,N_25469);
or U28957 (N_28957,N_25408,N_26242);
nand U28958 (N_28958,N_25249,N_26363);
or U28959 (N_28959,N_25418,N_27255);
or U28960 (N_28960,N_25706,N_26127);
nor U28961 (N_28961,N_27009,N_25007);
xnor U28962 (N_28962,N_25088,N_25257);
nand U28963 (N_28963,N_25197,N_25914);
nand U28964 (N_28964,N_27467,N_25398);
xor U28965 (N_28965,N_25549,N_25634);
nand U28966 (N_28966,N_26096,N_26938);
nand U28967 (N_28967,N_25074,N_27415);
and U28968 (N_28968,N_25236,N_25955);
or U28969 (N_28969,N_25897,N_27326);
nand U28970 (N_28970,N_25358,N_26645);
and U28971 (N_28971,N_25323,N_26342);
xor U28972 (N_28972,N_27080,N_27067);
and U28973 (N_28973,N_25467,N_26963);
xnor U28974 (N_28974,N_27288,N_26218);
and U28975 (N_28975,N_27244,N_27255);
nor U28976 (N_28976,N_26811,N_25021);
nand U28977 (N_28977,N_26866,N_26209);
or U28978 (N_28978,N_25699,N_27123);
xnor U28979 (N_28979,N_25785,N_26357);
or U28980 (N_28980,N_27499,N_26818);
or U28981 (N_28981,N_25440,N_25999);
xnor U28982 (N_28982,N_25763,N_25363);
nand U28983 (N_28983,N_27270,N_25338);
and U28984 (N_28984,N_26963,N_27116);
xnor U28985 (N_28985,N_27265,N_26249);
nand U28986 (N_28986,N_26824,N_26737);
nand U28987 (N_28987,N_26653,N_26618);
and U28988 (N_28988,N_25988,N_26776);
nor U28989 (N_28989,N_26340,N_26876);
nor U28990 (N_28990,N_26837,N_25523);
or U28991 (N_28991,N_25209,N_27259);
and U28992 (N_28992,N_26757,N_25381);
xnor U28993 (N_28993,N_26212,N_25234);
and U28994 (N_28994,N_26611,N_27108);
and U28995 (N_28995,N_25413,N_27400);
and U28996 (N_28996,N_25042,N_27370);
and U28997 (N_28997,N_26287,N_25931);
xnor U28998 (N_28998,N_25004,N_25958);
nor U28999 (N_28999,N_26312,N_25497);
or U29000 (N_29000,N_26311,N_26096);
nor U29001 (N_29001,N_27436,N_26443);
nand U29002 (N_29002,N_26339,N_27302);
and U29003 (N_29003,N_26256,N_25051);
and U29004 (N_29004,N_27260,N_27236);
nand U29005 (N_29005,N_25700,N_26119);
or U29006 (N_29006,N_25472,N_27411);
xor U29007 (N_29007,N_26307,N_26121);
nor U29008 (N_29008,N_26689,N_27096);
and U29009 (N_29009,N_26917,N_27122);
nor U29010 (N_29010,N_26822,N_25230);
xnor U29011 (N_29011,N_26170,N_26515);
nor U29012 (N_29012,N_27470,N_25250);
and U29013 (N_29013,N_25748,N_27331);
nand U29014 (N_29014,N_26740,N_26789);
and U29015 (N_29015,N_25799,N_26874);
nand U29016 (N_29016,N_25805,N_27326);
nand U29017 (N_29017,N_25395,N_25532);
nor U29018 (N_29018,N_26560,N_26621);
nor U29019 (N_29019,N_26318,N_26833);
nand U29020 (N_29020,N_25535,N_26602);
nand U29021 (N_29021,N_26736,N_26196);
and U29022 (N_29022,N_25022,N_25684);
xnor U29023 (N_29023,N_27262,N_25381);
xor U29024 (N_29024,N_25904,N_26353);
nand U29025 (N_29025,N_26567,N_25148);
or U29026 (N_29026,N_25971,N_27151);
and U29027 (N_29027,N_26812,N_25447);
nand U29028 (N_29028,N_27221,N_26442);
or U29029 (N_29029,N_26525,N_25088);
and U29030 (N_29030,N_26204,N_25813);
xnor U29031 (N_29031,N_25447,N_26844);
nand U29032 (N_29032,N_26102,N_26612);
and U29033 (N_29033,N_27480,N_26714);
or U29034 (N_29034,N_25181,N_25529);
or U29035 (N_29035,N_25101,N_25520);
nand U29036 (N_29036,N_27448,N_25928);
and U29037 (N_29037,N_26670,N_26537);
nand U29038 (N_29038,N_26324,N_25922);
xnor U29039 (N_29039,N_26672,N_26012);
xor U29040 (N_29040,N_26300,N_25174);
or U29041 (N_29041,N_25915,N_26615);
or U29042 (N_29042,N_26957,N_25172);
and U29043 (N_29043,N_25788,N_25308);
nand U29044 (N_29044,N_27444,N_27332);
nand U29045 (N_29045,N_27412,N_27282);
nor U29046 (N_29046,N_26847,N_27172);
nor U29047 (N_29047,N_27388,N_27297);
xnor U29048 (N_29048,N_25404,N_26646);
xnor U29049 (N_29049,N_26372,N_25175);
nor U29050 (N_29050,N_26509,N_26297);
xnor U29051 (N_29051,N_25159,N_26147);
xor U29052 (N_29052,N_26332,N_25169);
nor U29053 (N_29053,N_26787,N_27208);
nor U29054 (N_29054,N_26125,N_25026);
and U29055 (N_29055,N_25198,N_25283);
and U29056 (N_29056,N_26408,N_26039);
nand U29057 (N_29057,N_26034,N_26930);
xnor U29058 (N_29058,N_25136,N_26852);
and U29059 (N_29059,N_26949,N_26814);
nor U29060 (N_29060,N_26266,N_27429);
nand U29061 (N_29061,N_26169,N_26859);
nor U29062 (N_29062,N_27180,N_25473);
or U29063 (N_29063,N_26446,N_26594);
or U29064 (N_29064,N_26752,N_26923);
or U29065 (N_29065,N_25425,N_26628);
and U29066 (N_29066,N_26759,N_26933);
and U29067 (N_29067,N_26762,N_25014);
nor U29068 (N_29068,N_27465,N_26466);
xor U29069 (N_29069,N_25801,N_25256);
and U29070 (N_29070,N_27414,N_27177);
or U29071 (N_29071,N_25518,N_26199);
nor U29072 (N_29072,N_26137,N_25816);
and U29073 (N_29073,N_25872,N_26858);
and U29074 (N_29074,N_27001,N_25178);
or U29075 (N_29075,N_27076,N_26285);
or U29076 (N_29076,N_25126,N_25505);
nor U29077 (N_29077,N_26913,N_27177);
xnor U29078 (N_29078,N_25695,N_27069);
nor U29079 (N_29079,N_26387,N_25726);
nor U29080 (N_29080,N_26207,N_26314);
xnor U29081 (N_29081,N_26846,N_26866);
and U29082 (N_29082,N_27452,N_26113);
or U29083 (N_29083,N_25618,N_26821);
or U29084 (N_29084,N_25754,N_25623);
xor U29085 (N_29085,N_25116,N_25139);
nand U29086 (N_29086,N_26534,N_27487);
and U29087 (N_29087,N_25326,N_25024);
nor U29088 (N_29088,N_26913,N_27000);
or U29089 (N_29089,N_25721,N_25024);
nand U29090 (N_29090,N_25622,N_25117);
xnor U29091 (N_29091,N_26919,N_26062);
or U29092 (N_29092,N_26933,N_26452);
and U29093 (N_29093,N_25053,N_25115);
or U29094 (N_29094,N_26299,N_25890);
nor U29095 (N_29095,N_26507,N_25641);
or U29096 (N_29096,N_25828,N_26560);
xnor U29097 (N_29097,N_25201,N_26578);
nand U29098 (N_29098,N_25707,N_25144);
and U29099 (N_29099,N_25895,N_26686);
xnor U29100 (N_29100,N_26804,N_26981);
or U29101 (N_29101,N_26943,N_26667);
or U29102 (N_29102,N_25300,N_26560);
or U29103 (N_29103,N_26922,N_26301);
and U29104 (N_29104,N_25862,N_25199);
nand U29105 (N_29105,N_26055,N_26768);
xnor U29106 (N_29106,N_26555,N_25728);
xor U29107 (N_29107,N_25780,N_25162);
and U29108 (N_29108,N_26998,N_26301);
xnor U29109 (N_29109,N_26452,N_26396);
nand U29110 (N_29110,N_26452,N_27033);
or U29111 (N_29111,N_26108,N_27155);
or U29112 (N_29112,N_25397,N_25781);
nand U29113 (N_29113,N_25420,N_27273);
nor U29114 (N_29114,N_26020,N_25767);
or U29115 (N_29115,N_25300,N_27367);
or U29116 (N_29116,N_26093,N_26086);
and U29117 (N_29117,N_25190,N_25068);
and U29118 (N_29118,N_25495,N_25855);
nor U29119 (N_29119,N_27381,N_26885);
nor U29120 (N_29120,N_27261,N_25168);
nand U29121 (N_29121,N_25377,N_25650);
and U29122 (N_29122,N_26965,N_26991);
or U29123 (N_29123,N_25180,N_26646);
xor U29124 (N_29124,N_26000,N_26144);
or U29125 (N_29125,N_26192,N_25020);
or U29126 (N_29126,N_27200,N_27209);
or U29127 (N_29127,N_26312,N_25918);
nor U29128 (N_29128,N_25555,N_26368);
nor U29129 (N_29129,N_25223,N_26131);
xor U29130 (N_29130,N_26129,N_25051);
and U29131 (N_29131,N_26137,N_25834);
xor U29132 (N_29132,N_26478,N_25440);
and U29133 (N_29133,N_26613,N_25054);
or U29134 (N_29134,N_26056,N_25951);
xor U29135 (N_29135,N_26547,N_25621);
or U29136 (N_29136,N_26043,N_27120);
or U29137 (N_29137,N_26973,N_25536);
nand U29138 (N_29138,N_25781,N_25274);
xnor U29139 (N_29139,N_27368,N_26457);
or U29140 (N_29140,N_25843,N_25437);
xnor U29141 (N_29141,N_25799,N_26266);
xnor U29142 (N_29142,N_26878,N_25434);
and U29143 (N_29143,N_26952,N_27059);
and U29144 (N_29144,N_25218,N_25343);
and U29145 (N_29145,N_27335,N_25928);
or U29146 (N_29146,N_26222,N_27331);
nand U29147 (N_29147,N_25161,N_26021);
nand U29148 (N_29148,N_26634,N_25790);
nor U29149 (N_29149,N_25930,N_26404);
and U29150 (N_29150,N_25652,N_25883);
nand U29151 (N_29151,N_25429,N_25799);
nand U29152 (N_29152,N_25940,N_25846);
and U29153 (N_29153,N_25720,N_26765);
or U29154 (N_29154,N_26854,N_27449);
xor U29155 (N_29155,N_25200,N_26991);
and U29156 (N_29156,N_26833,N_25450);
nor U29157 (N_29157,N_26854,N_27058);
nor U29158 (N_29158,N_25704,N_27461);
xnor U29159 (N_29159,N_27245,N_26941);
nand U29160 (N_29160,N_25809,N_26543);
xnor U29161 (N_29161,N_25627,N_27218);
or U29162 (N_29162,N_26391,N_27184);
nor U29163 (N_29163,N_25114,N_26419);
or U29164 (N_29164,N_26117,N_26607);
nand U29165 (N_29165,N_25622,N_27064);
xor U29166 (N_29166,N_26937,N_27005);
nand U29167 (N_29167,N_27169,N_25048);
xor U29168 (N_29168,N_27226,N_26128);
xor U29169 (N_29169,N_25182,N_25245);
and U29170 (N_29170,N_26743,N_27457);
xor U29171 (N_29171,N_25074,N_25315);
nand U29172 (N_29172,N_25979,N_26063);
and U29173 (N_29173,N_26187,N_26680);
nor U29174 (N_29174,N_25624,N_25909);
xnor U29175 (N_29175,N_26325,N_25502);
xnor U29176 (N_29176,N_27389,N_27131);
nor U29177 (N_29177,N_25899,N_25821);
nor U29178 (N_29178,N_26984,N_27274);
and U29179 (N_29179,N_25770,N_26696);
and U29180 (N_29180,N_26311,N_25676);
and U29181 (N_29181,N_26397,N_27445);
nor U29182 (N_29182,N_25575,N_26833);
nand U29183 (N_29183,N_25587,N_27310);
nand U29184 (N_29184,N_25976,N_25817);
xnor U29185 (N_29185,N_25862,N_26707);
nor U29186 (N_29186,N_26237,N_25637);
or U29187 (N_29187,N_27004,N_26002);
or U29188 (N_29188,N_25896,N_26950);
or U29189 (N_29189,N_26318,N_25642);
or U29190 (N_29190,N_25772,N_26760);
nand U29191 (N_29191,N_26490,N_25627);
nand U29192 (N_29192,N_25500,N_25516);
and U29193 (N_29193,N_25759,N_26295);
and U29194 (N_29194,N_26421,N_25601);
nor U29195 (N_29195,N_25134,N_25847);
or U29196 (N_29196,N_25830,N_25632);
nand U29197 (N_29197,N_26890,N_26637);
and U29198 (N_29198,N_26342,N_25927);
and U29199 (N_29199,N_25592,N_25729);
or U29200 (N_29200,N_26000,N_26683);
nand U29201 (N_29201,N_26975,N_26026);
xor U29202 (N_29202,N_25771,N_27329);
nor U29203 (N_29203,N_27075,N_25864);
and U29204 (N_29204,N_25442,N_25964);
xor U29205 (N_29205,N_26799,N_27333);
and U29206 (N_29206,N_26739,N_26126);
nor U29207 (N_29207,N_27434,N_25167);
nand U29208 (N_29208,N_27366,N_25274);
nor U29209 (N_29209,N_26314,N_26829);
and U29210 (N_29210,N_26393,N_25234);
nand U29211 (N_29211,N_25359,N_26783);
nand U29212 (N_29212,N_27425,N_25567);
nor U29213 (N_29213,N_25578,N_25350);
xor U29214 (N_29214,N_25879,N_26422);
or U29215 (N_29215,N_25082,N_26376);
nor U29216 (N_29216,N_25027,N_25506);
xnor U29217 (N_29217,N_25206,N_25054);
nand U29218 (N_29218,N_25466,N_26666);
nand U29219 (N_29219,N_26091,N_26063);
and U29220 (N_29220,N_27143,N_26861);
xnor U29221 (N_29221,N_25299,N_26856);
and U29222 (N_29222,N_25355,N_25138);
nand U29223 (N_29223,N_25605,N_26510);
nor U29224 (N_29224,N_26899,N_26593);
xor U29225 (N_29225,N_25253,N_25504);
or U29226 (N_29226,N_27472,N_26298);
xnor U29227 (N_29227,N_26342,N_25597);
and U29228 (N_29228,N_27448,N_25367);
and U29229 (N_29229,N_26713,N_25672);
nor U29230 (N_29230,N_26287,N_25556);
nand U29231 (N_29231,N_27313,N_26779);
nand U29232 (N_29232,N_25732,N_25220);
nand U29233 (N_29233,N_27092,N_25458);
xor U29234 (N_29234,N_27334,N_25567);
or U29235 (N_29235,N_26271,N_25945);
xnor U29236 (N_29236,N_25003,N_25422);
and U29237 (N_29237,N_25262,N_27120);
nand U29238 (N_29238,N_26410,N_25999);
nor U29239 (N_29239,N_26730,N_26854);
or U29240 (N_29240,N_27406,N_27270);
or U29241 (N_29241,N_27465,N_27034);
nand U29242 (N_29242,N_25954,N_26744);
nor U29243 (N_29243,N_25532,N_25581);
xnor U29244 (N_29244,N_27299,N_25828);
nand U29245 (N_29245,N_25484,N_25420);
nor U29246 (N_29246,N_26337,N_27460);
xnor U29247 (N_29247,N_27097,N_26457);
or U29248 (N_29248,N_26189,N_26097);
or U29249 (N_29249,N_26732,N_25008);
nor U29250 (N_29250,N_26571,N_25208);
nor U29251 (N_29251,N_26530,N_25413);
xnor U29252 (N_29252,N_27258,N_25581);
nor U29253 (N_29253,N_27134,N_25860);
and U29254 (N_29254,N_27288,N_26609);
xnor U29255 (N_29255,N_25551,N_27108);
or U29256 (N_29256,N_27228,N_25678);
and U29257 (N_29257,N_25500,N_25208);
nor U29258 (N_29258,N_25687,N_25599);
xor U29259 (N_29259,N_25011,N_25272);
xnor U29260 (N_29260,N_25881,N_26317);
and U29261 (N_29261,N_27464,N_26827);
and U29262 (N_29262,N_25305,N_27031);
xor U29263 (N_29263,N_25181,N_25967);
and U29264 (N_29264,N_25251,N_25544);
or U29265 (N_29265,N_25145,N_25090);
nor U29266 (N_29266,N_26335,N_27425);
nand U29267 (N_29267,N_26510,N_25055);
xnor U29268 (N_29268,N_26488,N_27212);
xor U29269 (N_29269,N_26021,N_25890);
or U29270 (N_29270,N_26192,N_25065);
xor U29271 (N_29271,N_25574,N_26096);
nor U29272 (N_29272,N_25941,N_27320);
nand U29273 (N_29273,N_27497,N_25439);
and U29274 (N_29274,N_25493,N_25337);
and U29275 (N_29275,N_26472,N_26041);
nor U29276 (N_29276,N_25155,N_25471);
and U29277 (N_29277,N_27302,N_26014);
or U29278 (N_29278,N_26343,N_26070);
or U29279 (N_29279,N_25399,N_26136);
xnor U29280 (N_29280,N_25348,N_26948);
and U29281 (N_29281,N_27291,N_25378);
nor U29282 (N_29282,N_27210,N_25606);
xnor U29283 (N_29283,N_25420,N_27276);
or U29284 (N_29284,N_25517,N_26447);
nand U29285 (N_29285,N_27181,N_25794);
or U29286 (N_29286,N_25640,N_27419);
nor U29287 (N_29287,N_25635,N_25448);
nor U29288 (N_29288,N_25797,N_25973);
nor U29289 (N_29289,N_25275,N_26673);
nor U29290 (N_29290,N_25238,N_25044);
or U29291 (N_29291,N_25885,N_26397);
nor U29292 (N_29292,N_26034,N_27120);
and U29293 (N_29293,N_25667,N_26184);
nor U29294 (N_29294,N_25360,N_26657);
xnor U29295 (N_29295,N_26183,N_27309);
nor U29296 (N_29296,N_27068,N_26230);
or U29297 (N_29297,N_26710,N_25669);
nor U29298 (N_29298,N_27048,N_25345);
nand U29299 (N_29299,N_25110,N_25866);
nand U29300 (N_29300,N_26224,N_26045);
and U29301 (N_29301,N_27114,N_25046);
nor U29302 (N_29302,N_27483,N_27146);
nor U29303 (N_29303,N_26239,N_25648);
and U29304 (N_29304,N_25539,N_26294);
nand U29305 (N_29305,N_25202,N_25578);
nor U29306 (N_29306,N_25956,N_26348);
xor U29307 (N_29307,N_25385,N_27038);
nor U29308 (N_29308,N_26376,N_27138);
nor U29309 (N_29309,N_27043,N_26748);
and U29310 (N_29310,N_27208,N_25936);
nand U29311 (N_29311,N_26501,N_26566);
nand U29312 (N_29312,N_25333,N_26455);
nor U29313 (N_29313,N_26163,N_27030);
nor U29314 (N_29314,N_27056,N_25662);
nand U29315 (N_29315,N_26531,N_27228);
nand U29316 (N_29316,N_26387,N_26618);
or U29317 (N_29317,N_27153,N_26043);
xor U29318 (N_29318,N_26649,N_26730);
nor U29319 (N_29319,N_26692,N_26272);
xnor U29320 (N_29320,N_26627,N_25492);
or U29321 (N_29321,N_26599,N_25960);
xnor U29322 (N_29322,N_26684,N_25061);
and U29323 (N_29323,N_26695,N_26480);
nand U29324 (N_29324,N_27263,N_27453);
and U29325 (N_29325,N_25553,N_26832);
nand U29326 (N_29326,N_26593,N_25995);
and U29327 (N_29327,N_27308,N_26551);
and U29328 (N_29328,N_25234,N_25721);
or U29329 (N_29329,N_27475,N_26851);
and U29330 (N_29330,N_25277,N_26124);
and U29331 (N_29331,N_26214,N_25105);
xor U29332 (N_29332,N_25891,N_26741);
nor U29333 (N_29333,N_26951,N_26821);
and U29334 (N_29334,N_26511,N_27489);
xnor U29335 (N_29335,N_25565,N_25756);
nand U29336 (N_29336,N_27024,N_25482);
nand U29337 (N_29337,N_27439,N_26147);
nor U29338 (N_29338,N_25438,N_26238);
nand U29339 (N_29339,N_26920,N_27437);
nand U29340 (N_29340,N_26853,N_25833);
nand U29341 (N_29341,N_26783,N_26152);
nor U29342 (N_29342,N_26201,N_25463);
xor U29343 (N_29343,N_25614,N_27432);
nor U29344 (N_29344,N_27089,N_25167);
nand U29345 (N_29345,N_27078,N_27181);
xnor U29346 (N_29346,N_25409,N_27097);
or U29347 (N_29347,N_26391,N_26050);
xor U29348 (N_29348,N_26683,N_26301);
and U29349 (N_29349,N_26262,N_25506);
nor U29350 (N_29350,N_26871,N_26332);
nand U29351 (N_29351,N_26706,N_25491);
and U29352 (N_29352,N_27303,N_25169);
nor U29353 (N_29353,N_27499,N_27168);
or U29354 (N_29354,N_26211,N_26932);
and U29355 (N_29355,N_25138,N_26002);
nor U29356 (N_29356,N_25493,N_27498);
nand U29357 (N_29357,N_25058,N_27049);
nor U29358 (N_29358,N_26210,N_27157);
nand U29359 (N_29359,N_26201,N_25856);
and U29360 (N_29360,N_26767,N_27227);
and U29361 (N_29361,N_25857,N_25825);
or U29362 (N_29362,N_26743,N_25225);
or U29363 (N_29363,N_26652,N_26635);
or U29364 (N_29364,N_26034,N_26564);
and U29365 (N_29365,N_26629,N_25425);
or U29366 (N_29366,N_26449,N_27283);
nor U29367 (N_29367,N_26549,N_27259);
or U29368 (N_29368,N_27074,N_25746);
nor U29369 (N_29369,N_26894,N_25258);
xnor U29370 (N_29370,N_25916,N_25447);
nand U29371 (N_29371,N_26459,N_25864);
nor U29372 (N_29372,N_26358,N_25587);
and U29373 (N_29373,N_25487,N_27143);
xor U29374 (N_29374,N_25707,N_27011);
and U29375 (N_29375,N_26801,N_27117);
and U29376 (N_29376,N_26989,N_25050);
or U29377 (N_29377,N_27439,N_25969);
or U29378 (N_29378,N_26284,N_26387);
or U29379 (N_29379,N_25903,N_26784);
xor U29380 (N_29380,N_25500,N_25641);
nand U29381 (N_29381,N_26191,N_27395);
or U29382 (N_29382,N_27494,N_25227);
or U29383 (N_29383,N_25134,N_26825);
nand U29384 (N_29384,N_25418,N_25819);
nor U29385 (N_29385,N_26184,N_27046);
nor U29386 (N_29386,N_26005,N_26633);
nor U29387 (N_29387,N_25667,N_26946);
xnor U29388 (N_29388,N_26995,N_26910);
xnor U29389 (N_29389,N_27287,N_26613);
xnor U29390 (N_29390,N_25942,N_26934);
or U29391 (N_29391,N_26103,N_25851);
or U29392 (N_29392,N_26351,N_25598);
xnor U29393 (N_29393,N_25556,N_27077);
nand U29394 (N_29394,N_25234,N_26585);
xnor U29395 (N_29395,N_26575,N_25446);
and U29396 (N_29396,N_27311,N_26833);
and U29397 (N_29397,N_26038,N_26735);
and U29398 (N_29398,N_26929,N_26376);
nor U29399 (N_29399,N_27122,N_26354);
and U29400 (N_29400,N_26639,N_26615);
xnor U29401 (N_29401,N_25976,N_25511);
or U29402 (N_29402,N_25363,N_26402);
and U29403 (N_29403,N_25581,N_25823);
or U29404 (N_29404,N_27475,N_26214);
nor U29405 (N_29405,N_26512,N_26833);
nand U29406 (N_29406,N_26134,N_26075);
or U29407 (N_29407,N_26905,N_25726);
and U29408 (N_29408,N_25310,N_25608);
and U29409 (N_29409,N_25990,N_25078);
nand U29410 (N_29410,N_27186,N_25514);
nand U29411 (N_29411,N_26407,N_26831);
or U29412 (N_29412,N_26815,N_25036);
or U29413 (N_29413,N_26313,N_26446);
and U29414 (N_29414,N_26787,N_26544);
xor U29415 (N_29415,N_26072,N_26523);
xnor U29416 (N_29416,N_27405,N_27341);
xnor U29417 (N_29417,N_27179,N_25072);
or U29418 (N_29418,N_25608,N_26272);
xnor U29419 (N_29419,N_27141,N_25112);
xor U29420 (N_29420,N_26491,N_25989);
or U29421 (N_29421,N_27144,N_25180);
xor U29422 (N_29422,N_25368,N_25678);
xor U29423 (N_29423,N_26723,N_27157);
xnor U29424 (N_29424,N_25464,N_27483);
nand U29425 (N_29425,N_27219,N_26738);
and U29426 (N_29426,N_26277,N_27068);
and U29427 (N_29427,N_26180,N_25911);
xnor U29428 (N_29428,N_25549,N_27330);
xor U29429 (N_29429,N_26053,N_26189);
nor U29430 (N_29430,N_26579,N_25776);
and U29431 (N_29431,N_27350,N_25046);
nor U29432 (N_29432,N_25756,N_25050);
xnor U29433 (N_29433,N_26355,N_25582);
and U29434 (N_29434,N_26926,N_25746);
nor U29435 (N_29435,N_26300,N_25444);
and U29436 (N_29436,N_25046,N_25070);
nand U29437 (N_29437,N_25624,N_25130);
nor U29438 (N_29438,N_26720,N_26090);
and U29439 (N_29439,N_27086,N_27021);
and U29440 (N_29440,N_26211,N_25067);
xor U29441 (N_29441,N_25354,N_26064);
nor U29442 (N_29442,N_25363,N_26962);
and U29443 (N_29443,N_26141,N_25075);
and U29444 (N_29444,N_27134,N_25072);
nor U29445 (N_29445,N_26739,N_27097);
nand U29446 (N_29446,N_27069,N_26414);
and U29447 (N_29447,N_27289,N_27209);
and U29448 (N_29448,N_26373,N_26273);
nand U29449 (N_29449,N_26853,N_25175);
nand U29450 (N_29450,N_26654,N_26825);
or U29451 (N_29451,N_26019,N_25242);
nand U29452 (N_29452,N_25489,N_26568);
and U29453 (N_29453,N_26505,N_25070);
nor U29454 (N_29454,N_27246,N_26804);
xor U29455 (N_29455,N_27488,N_25832);
and U29456 (N_29456,N_27380,N_25407);
xor U29457 (N_29457,N_25087,N_25328);
nor U29458 (N_29458,N_25265,N_27274);
or U29459 (N_29459,N_27481,N_26101);
nor U29460 (N_29460,N_25945,N_25212);
and U29461 (N_29461,N_27291,N_26586);
nor U29462 (N_29462,N_26436,N_25722);
nor U29463 (N_29463,N_27276,N_25062);
nor U29464 (N_29464,N_25953,N_27201);
nor U29465 (N_29465,N_25598,N_27335);
nor U29466 (N_29466,N_26701,N_27449);
nand U29467 (N_29467,N_26707,N_25664);
and U29468 (N_29468,N_27442,N_25606);
nand U29469 (N_29469,N_26099,N_26404);
nor U29470 (N_29470,N_27409,N_26299);
nor U29471 (N_29471,N_25677,N_25569);
or U29472 (N_29472,N_27332,N_25573);
and U29473 (N_29473,N_26338,N_25645);
and U29474 (N_29474,N_26173,N_26236);
and U29475 (N_29475,N_27235,N_27006);
or U29476 (N_29476,N_25452,N_25601);
or U29477 (N_29477,N_25059,N_25812);
nand U29478 (N_29478,N_25165,N_26026);
xnor U29479 (N_29479,N_25233,N_27436);
nor U29480 (N_29480,N_25151,N_26636);
nand U29481 (N_29481,N_27342,N_25093);
or U29482 (N_29482,N_25618,N_27425);
or U29483 (N_29483,N_25919,N_26879);
or U29484 (N_29484,N_25038,N_26769);
and U29485 (N_29485,N_25559,N_26380);
and U29486 (N_29486,N_25652,N_25913);
xnor U29487 (N_29487,N_27032,N_25437);
nor U29488 (N_29488,N_25023,N_25134);
nor U29489 (N_29489,N_25353,N_25240);
or U29490 (N_29490,N_25752,N_25542);
and U29491 (N_29491,N_25788,N_27091);
and U29492 (N_29492,N_25651,N_26696);
nor U29493 (N_29493,N_26676,N_26371);
nand U29494 (N_29494,N_25183,N_26515);
nor U29495 (N_29495,N_27233,N_27244);
and U29496 (N_29496,N_26116,N_26589);
and U29497 (N_29497,N_27355,N_26542);
xor U29498 (N_29498,N_27002,N_27364);
nor U29499 (N_29499,N_26634,N_25690);
xnor U29500 (N_29500,N_26478,N_26063);
nand U29501 (N_29501,N_26191,N_27133);
nand U29502 (N_29502,N_26438,N_27029);
nor U29503 (N_29503,N_25509,N_27427);
nor U29504 (N_29504,N_25749,N_25514);
nand U29505 (N_29505,N_25688,N_25963);
or U29506 (N_29506,N_26470,N_27474);
or U29507 (N_29507,N_25705,N_26700);
nand U29508 (N_29508,N_26082,N_25921);
and U29509 (N_29509,N_25434,N_25969);
xnor U29510 (N_29510,N_26765,N_27203);
or U29511 (N_29511,N_27251,N_26760);
xor U29512 (N_29512,N_27101,N_26856);
xnor U29513 (N_29513,N_26890,N_26166);
xnor U29514 (N_29514,N_27151,N_27022);
xor U29515 (N_29515,N_25805,N_25234);
and U29516 (N_29516,N_25918,N_26205);
nand U29517 (N_29517,N_25383,N_25002);
and U29518 (N_29518,N_27285,N_26731);
nand U29519 (N_29519,N_27218,N_25028);
nor U29520 (N_29520,N_25580,N_25186);
nand U29521 (N_29521,N_25190,N_26721);
or U29522 (N_29522,N_26976,N_26797);
nand U29523 (N_29523,N_26901,N_26044);
and U29524 (N_29524,N_27314,N_27094);
nand U29525 (N_29525,N_26568,N_26084);
nor U29526 (N_29526,N_25364,N_26651);
xnor U29527 (N_29527,N_26758,N_25791);
nor U29528 (N_29528,N_26922,N_27242);
and U29529 (N_29529,N_26961,N_26136);
xnor U29530 (N_29530,N_26593,N_27469);
xor U29531 (N_29531,N_26849,N_25608);
and U29532 (N_29532,N_25071,N_27014);
nand U29533 (N_29533,N_26463,N_26119);
and U29534 (N_29534,N_26561,N_26968);
nand U29535 (N_29535,N_26224,N_25623);
and U29536 (N_29536,N_25332,N_25614);
nand U29537 (N_29537,N_25572,N_25831);
or U29538 (N_29538,N_27004,N_25024);
nand U29539 (N_29539,N_26237,N_26863);
nor U29540 (N_29540,N_25028,N_26344);
nand U29541 (N_29541,N_26473,N_25953);
and U29542 (N_29542,N_25292,N_26302);
or U29543 (N_29543,N_26027,N_27298);
and U29544 (N_29544,N_26488,N_25915);
nor U29545 (N_29545,N_25239,N_26493);
nand U29546 (N_29546,N_26820,N_25033);
nor U29547 (N_29547,N_27009,N_26480);
and U29548 (N_29548,N_26390,N_25600);
or U29549 (N_29549,N_27320,N_27386);
xor U29550 (N_29550,N_25629,N_25616);
or U29551 (N_29551,N_27023,N_25815);
nor U29552 (N_29552,N_26573,N_25633);
or U29553 (N_29553,N_26290,N_26074);
nand U29554 (N_29554,N_26666,N_25323);
xor U29555 (N_29555,N_26859,N_26301);
or U29556 (N_29556,N_27295,N_26496);
nand U29557 (N_29557,N_26506,N_25495);
or U29558 (N_29558,N_27462,N_26946);
nand U29559 (N_29559,N_26926,N_25102);
xor U29560 (N_29560,N_26728,N_26701);
or U29561 (N_29561,N_25496,N_25146);
or U29562 (N_29562,N_26901,N_26173);
nand U29563 (N_29563,N_26164,N_25119);
and U29564 (N_29564,N_25434,N_26292);
nand U29565 (N_29565,N_25649,N_26429);
or U29566 (N_29566,N_26895,N_25154);
xnor U29567 (N_29567,N_26733,N_25018);
xnor U29568 (N_29568,N_26013,N_27182);
xor U29569 (N_29569,N_27220,N_25816);
nor U29570 (N_29570,N_27392,N_26808);
or U29571 (N_29571,N_25451,N_26033);
nor U29572 (N_29572,N_25662,N_26588);
xor U29573 (N_29573,N_26174,N_25771);
xor U29574 (N_29574,N_25354,N_26452);
and U29575 (N_29575,N_25422,N_25157);
and U29576 (N_29576,N_25712,N_26085);
nand U29577 (N_29577,N_26424,N_27457);
or U29578 (N_29578,N_26513,N_27241);
and U29579 (N_29579,N_25009,N_25096);
nor U29580 (N_29580,N_26167,N_26934);
xor U29581 (N_29581,N_26044,N_25087);
xnor U29582 (N_29582,N_26509,N_27210);
or U29583 (N_29583,N_26675,N_27357);
xnor U29584 (N_29584,N_25081,N_26958);
nand U29585 (N_29585,N_26494,N_26552);
or U29586 (N_29586,N_25919,N_25991);
nor U29587 (N_29587,N_26404,N_25963);
nor U29588 (N_29588,N_25364,N_26283);
or U29589 (N_29589,N_25802,N_26612);
or U29590 (N_29590,N_25303,N_25707);
and U29591 (N_29591,N_27041,N_26998);
nor U29592 (N_29592,N_26914,N_26726);
xor U29593 (N_29593,N_26119,N_25505);
nor U29594 (N_29594,N_26304,N_25153);
xnor U29595 (N_29595,N_26577,N_26893);
or U29596 (N_29596,N_25188,N_25369);
nor U29597 (N_29597,N_26357,N_26388);
xor U29598 (N_29598,N_25665,N_27348);
xor U29599 (N_29599,N_26240,N_26008);
nand U29600 (N_29600,N_25332,N_25766);
nand U29601 (N_29601,N_26128,N_26133);
nor U29602 (N_29602,N_25745,N_26726);
nor U29603 (N_29603,N_26816,N_27359);
xnor U29604 (N_29604,N_26859,N_27299);
nor U29605 (N_29605,N_25652,N_26260);
and U29606 (N_29606,N_26283,N_25293);
nand U29607 (N_29607,N_25040,N_26954);
nand U29608 (N_29608,N_27328,N_25156);
xor U29609 (N_29609,N_25121,N_26033);
nand U29610 (N_29610,N_25217,N_27145);
nand U29611 (N_29611,N_25759,N_26554);
nand U29612 (N_29612,N_25323,N_26313);
or U29613 (N_29613,N_26771,N_27058);
and U29614 (N_29614,N_26436,N_26335);
xnor U29615 (N_29615,N_26465,N_25348);
nor U29616 (N_29616,N_26167,N_27321);
xor U29617 (N_29617,N_25353,N_26419);
or U29618 (N_29618,N_25287,N_25832);
nor U29619 (N_29619,N_25330,N_25769);
xnor U29620 (N_29620,N_26965,N_26043);
nand U29621 (N_29621,N_26581,N_26734);
nor U29622 (N_29622,N_26360,N_26361);
nand U29623 (N_29623,N_27072,N_26115);
nor U29624 (N_29624,N_27046,N_27280);
nor U29625 (N_29625,N_26670,N_25681);
nor U29626 (N_29626,N_26978,N_25065);
xnor U29627 (N_29627,N_25504,N_25261);
nand U29628 (N_29628,N_25924,N_27478);
nor U29629 (N_29629,N_25027,N_26365);
or U29630 (N_29630,N_26461,N_25336);
xnor U29631 (N_29631,N_25559,N_25975);
and U29632 (N_29632,N_26694,N_25071);
nor U29633 (N_29633,N_27323,N_25980);
nor U29634 (N_29634,N_25480,N_27066);
or U29635 (N_29635,N_25282,N_26465);
and U29636 (N_29636,N_26637,N_25563);
nand U29637 (N_29637,N_25619,N_25268);
nand U29638 (N_29638,N_26485,N_26237);
nor U29639 (N_29639,N_25523,N_25063);
xor U29640 (N_29640,N_25423,N_25863);
and U29641 (N_29641,N_27488,N_26974);
nand U29642 (N_29642,N_26050,N_26867);
xnor U29643 (N_29643,N_26176,N_25023);
and U29644 (N_29644,N_26459,N_25257);
xor U29645 (N_29645,N_26548,N_26087);
nor U29646 (N_29646,N_27012,N_26400);
xor U29647 (N_29647,N_26163,N_25968);
or U29648 (N_29648,N_26436,N_26338);
and U29649 (N_29649,N_26887,N_26488);
and U29650 (N_29650,N_25007,N_26558);
and U29651 (N_29651,N_25463,N_25648);
xor U29652 (N_29652,N_25975,N_25068);
or U29653 (N_29653,N_26619,N_26055);
xnor U29654 (N_29654,N_26765,N_26602);
and U29655 (N_29655,N_27144,N_26712);
nand U29656 (N_29656,N_27277,N_26041);
and U29657 (N_29657,N_26304,N_25247);
or U29658 (N_29658,N_25615,N_25692);
or U29659 (N_29659,N_25517,N_26495);
and U29660 (N_29660,N_25078,N_25969);
xnor U29661 (N_29661,N_26566,N_26947);
xnor U29662 (N_29662,N_27193,N_26206);
nor U29663 (N_29663,N_26210,N_25455);
nor U29664 (N_29664,N_27293,N_25041);
and U29665 (N_29665,N_25265,N_25461);
or U29666 (N_29666,N_26414,N_25808);
nor U29667 (N_29667,N_25451,N_27291);
nor U29668 (N_29668,N_26091,N_26650);
nor U29669 (N_29669,N_26724,N_27298);
and U29670 (N_29670,N_26682,N_26728);
or U29671 (N_29671,N_27146,N_25194);
nand U29672 (N_29672,N_27263,N_25712);
and U29673 (N_29673,N_26405,N_26407);
and U29674 (N_29674,N_26856,N_26528);
xor U29675 (N_29675,N_25521,N_27362);
or U29676 (N_29676,N_26908,N_25752);
nor U29677 (N_29677,N_26160,N_27213);
nor U29678 (N_29678,N_27352,N_25031);
nand U29679 (N_29679,N_25670,N_27425);
nand U29680 (N_29680,N_27420,N_25120);
nand U29681 (N_29681,N_27261,N_26044);
and U29682 (N_29682,N_25561,N_27323);
nor U29683 (N_29683,N_27098,N_27147);
or U29684 (N_29684,N_26446,N_26774);
nor U29685 (N_29685,N_26341,N_25303);
and U29686 (N_29686,N_26610,N_27386);
or U29687 (N_29687,N_26440,N_26846);
nor U29688 (N_29688,N_25074,N_27175);
and U29689 (N_29689,N_25644,N_25870);
xnor U29690 (N_29690,N_27123,N_25723);
and U29691 (N_29691,N_25636,N_26936);
nor U29692 (N_29692,N_26587,N_25564);
xor U29693 (N_29693,N_26871,N_25947);
nand U29694 (N_29694,N_27060,N_25494);
xor U29695 (N_29695,N_27272,N_25399);
and U29696 (N_29696,N_25285,N_27344);
and U29697 (N_29697,N_25569,N_27170);
nand U29698 (N_29698,N_25125,N_25329);
xor U29699 (N_29699,N_26816,N_25664);
xnor U29700 (N_29700,N_25944,N_25264);
or U29701 (N_29701,N_27063,N_26143);
and U29702 (N_29702,N_25235,N_25063);
nand U29703 (N_29703,N_25602,N_25842);
and U29704 (N_29704,N_27470,N_27192);
and U29705 (N_29705,N_26793,N_27148);
nand U29706 (N_29706,N_27476,N_25301);
and U29707 (N_29707,N_25544,N_25932);
nand U29708 (N_29708,N_25852,N_25193);
nor U29709 (N_29709,N_26596,N_26426);
or U29710 (N_29710,N_26742,N_25355);
or U29711 (N_29711,N_25701,N_27340);
nand U29712 (N_29712,N_26436,N_25132);
nand U29713 (N_29713,N_27190,N_26405);
nor U29714 (N_29714,N_26584,N_25820);
or U29715 (N_29715,N_26025,N_25792);
or U29716 (N_29716,N_26459,N_25113);
nor U29717 (N_29717,N_26408,N_26460);
nand U29718 (N_29718,N_26280,N_27232);
xor U29719 (N_29719,N_26606,N_26999);
or U29720 (N_29720,N_26628,N_27207);
nor U29721 (N_29721,N_26319,N_26627);
or U29722 (N_29722,N_26223,N_26138);
and U29723 (N_29723,N_27414,N_25211);
nand U29724 (N_29724,N_27314,N_26043);
xnor U29725 (N_29725,N_25663,N_25739);
and U29726 (N_29726,N_25060,N_25811);
or U29727 (N_29727,N_25617,N_26918);
nor U29728 (N_29728,N_25534,N_26570);
nand U29729 (N_29729,N_27388,N_25067);
nor U29730 (N_29730,N_25731,N_25529);
nor U29731 (N_29731,N_26624,N_26093);
and U29732 (N_29732,N_25691,N_27303);
or U29733 (N_29733,N_25706,N_26057);
nand U29734 (N_29734,N_26526,N_25293);
nor U29735 (N_29735,N_27178,N_25217);
nor U29736 (N_29736,N_26955,N_25228);
nand U29737 (N_29737,N_26596,N_25666);
nor U29738 (N_29738,N_25960,N_25534);
or U29739 (N_29739,N_26177,N_27118);
and U29740 (N_29740,N_25383,N_26843);
or U29741 (N_29741,N_26486,N_26247);
nand U29742 (N_29742,N_25269,N_25510);
and U29743 (N_29743,N_26947,N_27075);
or U29744 (N_29744,N_26984,N_25500);
or U29745 (N_29745,N_25944,N_26245);
and U29746 (N_29746,N_25963,N_27414);
nor U29747 (N_29747,N_27003,N_27357);
and U29748 (N_29748,N_26500,N_26425);
and U29749 (N_29749,N_25544,N_25572);
xnor U29750 (N_29750,N_25161,N_25379);
nor U29751 (N_29751,N_25995,N_25074);
nor U29752 (N_29752,N_25908,N_25455);
and U29753 (N_29753,N_27337,N_25585);
xnor U29754 (N_29754,N_25191,N_27418);
and U29755 (N_29755,N_26506,N_27288);
or U29756 (N_29756,N_26881,N_25679);
xnor U29757 (N_29757,N_25806,N_26510);
nor U29758 (N_29758,N_27026,N_26280);
xor U29759 (N_29759,N_27263,N_27052);
xor U29760 (N_29760,N_26875,N_26508);
and U29761 (N_29761,N_26695,N_25981);
and U29762 (N_29762,N_27304,N_25580);
xor U29763 (N_29763,N_25851,N_25765);
and U29764 (N_29764,N_26665,N_25208);
or U29765 (N_29765,N_26312,N_25574);
nand U29766 (N_29766,N_25687,N_26347);
nand U29767 (N_29767,N_27479,N_26678);
nor U29768 (N_29768,N_27097,N_25578);
and U29769 (N_29769,N_26431,N_26415);
and U29770 (N_29770,N_26985,N_25471);
or U29771 (N_29771,N_25337,N_25712);
nor U29772 (N_29772,N_25313,N_25522);
xnor U29773 (N_29773,N_26988,N_25694);
nand U29774 (N_29774,N_27334,N_25938);
and U29775 (N_29775,N_25968,N_25580);
nor U29776 (N_29776,N_26078,N_26324);
xnor U29777 (N_29777,N_25350,N_25387);
and U29778 (N_29778,N_25298,N_25789);
or U29779 (N_29779,N_26757,N_26783);
or U29780 (N_29780,N_25022,N_26501);
or U29781 (N_29781,N_25744,N_27048);
and U29782 (N_29782,N_26331,N_27373);
and U29783 (N_29783,N_26425,N_26989);
and U29784 (N_29784,N_27256,N_25441);
nor U29785 (N_29785,N_25401,N_26329);
nor U29786 (N_29786,N_25286,N_25555);
and U29787 (N_29787,N_27066,N_25674);
or U29788 (N_29788,N_25697,N_27444);
or U29789 (N_29789,N_25941,N_25693);
nand U29790 (N_29790,N_26382,N_25740);
xor U29791 (N_29791,N_26830,N_25880);
and U29792 (N_29792,N_26767,N_25167);
or U29793 (N_29793,N_25941,N_25982);
and U29794 (N_29794,N_25062,N_26480);
nand U29795 (N_29795,N_25425,N_26332);
nor U29796 (N_29796,N_26065,N_27008);
xor U29797 (N_29797,N_26975,N_26402);
or U29798 (N_29798,N_27366,N_25571);
xor U29799 (N_29799,N_25934,N_25290);
xnor U29800 (N_29800,N_26107,N_27238);
or U29801 (N_29801,N_26830,N_26663);
nor U29802 (N_29802,N_25430,N_25939);
and U29803 (N_29803,N_25667,N_25009);
nand U29804 (N_29804,N_25824,N_25517);
or U29805 (N_29805,N_26460,N_26961);
xor U29806 (N_29806,N_27099,N_26803);
nand U29807 (N_29807,N_25081,N_26971);
nor U29808 (N_29808,N_25838,N_25989);
or U29809 (N_29809,N_25432,N_27109);
xnor U29810 (N_29810,N_25712,N_26110);
nand U29811 (N_29811,N_27053,N_27387);
or U29812 (N_29812,N_26100,N_26612);
xnor U29813 (N_29813,N_26503,N_26383);
nor U29814 (N_29814,N_25262,N_27497);
and U29815 (N_29815,N_27471,N_25860);
and U29816 (N_29816,N_27255,N_25746);
xor U29817 (N_29817,N_26758,N_25191);
xor U29818 (N_29818,N_25379,N_25531);
and U29819 (N_29819,N_26579,N_25125);
and U29820 (N_29820,N_27392,N_25043);
nand U29821 (N_29821,N_25958,N_25926);
nand U29822 (N_29822,N_26056,N_26443);
nor U29823 (N_29823,N_25278,N_25789);
and U29824 (N_29824,N_25926,N_26517);
and U29825 (N_29825,N_25097,N_25887);
nand U29826 (N_29826,N_25092,N_27037);
nand U29827 (N_29827,N_27308,N_26337);
and U29828 (N_29828,N_27078,N_25768);
or U29829 (N_29829,N_26271,N_26415);
or U29830 (N_29830,N_26151,N_26447);
nand U29831 (N_29831,N_25242,N_26321);
nand U29832 (N_29832,N_25426,N_25557);
or U29833 (N_29833,N_25281,N_27268);
xor U29834 (N_29834,N_26449,N_27409);
nand U29835 (N_29835,N_25855,N_26203);
xor U29836 (N_29836,N_25408,N_27471);
xnor U29837 (N_29837,N_25276,N_27390);
or U29838 (N_29838,N_26096,N_27440);
nor U29839 (N_29839,N_25386,N_25376);
or U29840 (N_29840,N_26819,N_25781);
nand U29841 (N_29841,N_26814,N_26678);
nor U29842 (N_29842,N_25642,N_25731);
nor U29843 (N_29843,N_25182,N_26328);
xor U29844 (N_29844,N_26613,N_27073);
nor U29845 (N_29845,N_26694,N_27376);
nand U29846 (N_29846,N_27096,N_26727);
nand U29847 (N_29847,N_26829,N_26739);
and U29848 (N_29848,N_25620,N_25681);
or U29849 (N_29849,N_26472,N_25924);
nand U29850 (N_29850,N_25424,N_26273);
nor U29851 (N_29851,N_26915,N_26311);
and U29852 (N_29852,N_27264,N_25567);
xor U29853 (N_29853,N_25959,N_25475);
or U29854 (N_29854,N_26565,N_25610);
nor U29855 (N_29855,N_25981,N_25388);
nor U29856 (N_29856,N_27375,N_27089);
and U29857 (N_29857,N_27057,N_27058);
nor U29858 (N_29858,N_25168,N_27125);
xor U29859 (N_29859,N_25408,N_26525);
xor U29860 (N_29860,N_26376,N_25821);
nor U29861 (N_29861,N_26288,N_26449);
nor U29862 (N_29862,N_26356,N_25835);
and U29863 (N_29863,N_26942,N_26648);
nor U29864 (N_29864,N_25811,N_25149);
nand U29865 (N_29865,N_26959,N_25304);
or U29866 (N_29866,N_26612,N_25273);
nand U29867 (N_29867,N_25712,N_26960);
xor U29868 (N_29868,N_25514,N_25038);
nand U29869 (N_29869,N_27030,N_26316);
or U29870 (N_29870,N_25643,N_27225);
or U29871 (N_29871,N_25390,N_25398);
nor U29872 (N_29872,N_25212,N_26050);
or U29873 (N_29873,N_25477,N_25668);
nor U29874 (N_29874,N_25162,N_25019);
or U29875 (N_29875,N_27073,N_25172);
or U29876 (N_29876,N_25174,N_27457);
nor U29877 (N_29877,N_26550,N_26030);
and U29878 (N_29878,N_25307,N_27194);
nand U29879 (N_29879,N_25222,N_26104);
xnor U29880 (N_29880,N_25094,N_25590);
nor U29881 (N_29881,N_26208,N_26471);
nor U29882 (N_29882,N_27480,N_25867);
nor U29883 (N_29883,N_26521,N_26814);
xor U29884 (N_29884,N_25059,N_27413);
and U29885 (N_29885,N_27461,N_26324);
nor U29886 (N_29886,N_25991,N_26364);
nor U29887 (N_29887,N_27104,N_25601);
xor U29888 (N_29888,N_25019,N_26221);
or U29889 (N_29889,N_25450,N_26341);
xor U29890 (N_29890,N_26145,N_26335);
nand U29891 (N_29891,N_27180,N_25635);
xnor U29892 (N_29892,N_27163,N_27441);
nor U29893 (N_29893,N_26690,N_27181);
nand U29894 (N_29894,N_25208,N_26049);
and U29895 (N_29895,N_26847,N_27209);
nand U29896 (N_29896,N_27042,N_27432);
xnor U29897 (N_29897,N_26830,N_26913);
and U29898 (N_29898,N_27322,N_25178);
and U29899 (N_29899,N_27425,N_26176);
xor U29900 (N_29900,N_26015,N_26799);
nand U29901 (N_29901,N_26961,N_25713);
and U29902 (N_29902,N_25085,N_26769);
xnor U29903 (N_29903,N_26779,N_27078);
or U29904 (N_29904,N_27334,N_26987);
and U29905 (N_29905,N_25725,N_25180);
nor U29906 (N_29906,N_25262,N_26444);
nor U29907 (N_29907,N_25693,N_25107);
nor U29908 (N_29908,N_26486,N_26735);
and U29909 (N_29909,N_27392,N_26551);
and U29910 (N_29910,N_27100,N_27095);
xor U29911 (N_29911,N_25213,N_25698);
and U29912 (N_29912,N_26307,N_27314);
nor U29913 (N_29913,N_26514,N_26426);
and U29914 (N_29914,N_26942,N_26789);
and U29915 (N_29915,N_25654,N_25460);
nand U29916 (N_29916,N_25397,N_25112);
xnor U29917 (N_29917,N_26407,N_27145);
and U29918 (N_29918,N_26124,N_26449);
and U29919 (N_29919,N_26731,N_25930);
nand U29920 (N_29920,N_26712,N_26677);
or U29921 (N_29921,N_25066,N_27334);
and U29922 (N_29922,N_26885,N_26055);
nand U29923 (N_29923,N_27428,N_27253);
nand U29924 (N_29924,N_25855,N_25652);
nand U29925 (N_29925,N_26929,N_26152);
nand U29926 (N_29926,N_26838,N_26701);
nor U29927 (N_29927,N_25991,N_25010);
or U29928 (N_29928,N_26884,N_26208);
nor U29929 (N_29929,N_25216,N_25595);
or U29930 (N_29930,N_26221,N_26653);
nand U29931 (N_29931,N_25935,N_26521);
xor U29932 (N_29932,N_26933,N_26022);
or U29933 (N_29933,N_26478,N_26060);
and U29934 (N_29934,N_25367,N_25290);
nand U29935 (N_29935,N_26954,N_26400);
nand U29936 (N_29936,N_26286,N_25798);
and U29937 (N_29937,N_27326,N_26567);
nor U29938 (N_29938,N_27314,N_26079);
nand U29939 (N_29939,N_25825,N_26820);
xor U29940 (N_29940,N_26668,N_25344);
nand U29941 (N_29941,N_25184,N_26965);
or U29942 (N_29942,N_25900,N_25031);
nor U29943 (N_29943,N_26012,N_26990);
nand U29944 (N_29944,N_25708,N_25445);
nand U29945 (N_29945,N_26685,N_27340);
nor U29946 (N_29946,N_25281,N_27119);
nor U29947 (N_29947,N_26296,N_25011);
and U29948 (N_29948,N_25627,N_27321);
or U29949 (N_29949,N_26589,N_25408);
nand U29950 (N_29950,N_27206,N_26024);
or U29951 (N_29951,N_25522,N_26264);
xnor U29952 (N_29952,N_26213,N_25562);
or U29953 (N_29953,N_26344,N_25533);
and U29954 (N_29954,N_26727,N_26764);
and U29955 (N_29955,N_27121,N_25638);
nand U29956 (N_29956,N_27377,N_25842);
xnor U29957 (N_29957,N_25034,N_26635);
or U29958 (N_29958,N_26203,N_27184);
nand U29959 (N_29959,N_26713,N_26727);
xor U29960 (N_29960,N_25121,N_26324);
nand U29961 (N_29961,N_26767,N_26847);
nand U29962 (N_29962,N_26773,N_26057);
xor U29963 (N_29963,N_26127,N_26623);
nor U29964 (N_29964,N_27436,N_26590);
or U29965 (N_29965,N_26108,N_26452);
nor U29966 (N_29966,N_26363,N_25819);
or U29967 (N_29967,N_27230,N_25110);
xnor U29968 (N_29968,N_26626,N_25222);
and U29969 (N_29969,N_25739,N_26962);
xnor U29970 (N_29970,N_26599,N_25202);
nand U29971 (N_29971,N_27354,N_25517);
nor U29972 (N_29972,N_25125,N_25628);
xor U29973 (N_29973,N_25647,N_26331);
or U29974 (N_29974,N_25971,N_25590);
or U29975 (N_29975,N_27297,N_26623);
nor U29976 (N_29976,N_25390,N_25920);
and U29977 (N_29977,N_26569,N_26885);
nor U29978 (N_29978,N_25262,N_25002);
nor U29979 (N_29979,N_26087,N_27173);
and U29980 (N_29980,N_26557,N_25235);
or U29981 (N_29981,N_26511,N_25454);
xor U29982 (N_29982,N_27183,N_26719);
and U29983 (N_29983,N_26388,N_25717);
and U29984 (N_29984,N_25152,N_26101);
or U29985 (N_29985,N_25658,N_25639);
xnor U29986 (N_29986,N_27377,N_26676);
nand U29987 (N_29987,N_27069,N_26239);
nand U29988 (N_29988,N_25594,N_27273);
nor U29989 (N_29989,N_25755,N_26805);
nor U29990 (N_29990,N_25673,N_26714);
nand U29991 (N_29991,N_26892,N_26040);
and U29992 (N_29992,N_25563,N_25505);
xor U29993 (N_29993,N_26576,N_25429);
and U29994 (N_29994,N_26003,N_26727);
or U29995 (N_29995,N_26275,N_26578);
nor U29996 (N_29996,N_26472,N_27159);
xnor U29997 (N_29997,N_25541,N_26128);
nor U29998 (N_29998,N_26850,N_26947);
xor U29999 (N_29999,N_27102,N_25025);
nand U30000 (N_30000,N_29629,N_28470);
and U30001 (N_30001,N_29990,N_27911);
or U30002 (N_30002,N_29258,N_28831);
nor U30003 (N_30003,N_29577,N_28532);
nor U30004 (N_30004,N_28628,N_28841);
or U30005 (N_30005,N_29870,N_29017);
or U30006 (N_30006,N_29509,N_29021);
or U30007 (N_30007,N_28271,N_29063);
nor U30008 (N_30008,N_29222,N_28530);
nor U30009 (N_30009,N_28574,N_29574);
nor U30010 (N_30010,N_28169,N_27616);
or U30011 (N_30011,N_28144,N_28132);
nor U30012 (N_30012,N_27829,N_29849);
and U30013 (N_30013,N_28363,N_28160);
nand U30014 (N_30014,N_28550,N_29967);
or U30015 (N_30015,N_28100,N_29736);
nor U30016 (N_30016,N_28661,N_27681);
xnor U30017 (N_30017,N_29984,N_28340);
or U30018 (N_30018,N_29442,N_27672);
nor U30019 (N_30019,N_29330,N_29262);
nor U30020 (N_30020,N_29395,N_29275);
and U30021 (N_30021,N_29575,N_27569);
nand U30022 (N_30022,N_29050,N_28619);
and U30023 (N_30023,N_28905,N_28190);
and U30024 (N_30024,N_29435,N_29365);
or U30025 (N_30025,N_28672,N_29935);
xor U30026 (N_30026,N_28447,N_27804);
or U30027 (N_30027,N_28675,N_28255);
xnor U30028 (N_30028,N_29926,N_29093);
nor U30029 (N_30029,N_29468,N_29617);
nand U30030 (N_30030,N_27729,N_29476);
and U30031 (N_30031,N_28801,N_28591);
and U30032 (N_30032,N_28895,N_28967);
or U30033 (N_30033,N_29770,N_29631);
xor U30034 (N_30034,N_27834,N_29303);
xor U30035 (N_30035,N_29679,N_28156);
xor U30036 (N_30036,N_28108,N_28147);
nor U30037 (N_30037,N_29115,N_28388);
and U30038 (N_30038,N_28287,N_28537);
xnor U30039 (N_30039,N_28161,N_29372);
xnor U30040 (N_30040,N_29988,N_28982);
xnor U30041 (N_30041,N_28113,N_28378);
nand U30042 (N_30042,N_28561,N_28797);
and U30043 (N_30043,N_27667,N_28913);
xor U30044 (N_30044,N_29220,N_28579);
and U30045 (N_30045,N_29920,N_27972);
xnor U30046 (N_30046,N_29122,N_29046);
nor U30047 (N_30047,N_29841,N_28788);
nor U30048 (N_30048,N_28731,N_27590);
nand U30049 (N_30049,N_27784,N_29894);
nor U30050 (N_30050,N_28314,N_29380);
and U30051 (N_30051,N_27823,N_28868);
or U30052 (N_30052,N_29832,N_29661);
xor U30053 (N_30053,N_29359,N_29813);
and U30054 (N_30054,N_29453,N_29623);
nand U30055 (N_30055,N_28383,N_27604);
nor U30056 (N_30056,N_28010,N_28838);
nor U30057 (N_30057,N_28594,N_27579);
or U30058 (N_30058,N_29970,N_27827);
nand U30059 (N_30059,N_28517,N_27956);
nor U30060 (N_30060,N_29824,N_29100);
nand U30061 (N_30061,N_29178,N_28696);
or U30062 (N_30062,N_27927,N_29354);
nand U30063 (N_30063,N_28029,N_27586);
xor U30064 (N_30064,N_28624,N_29067);
nand U30065 (N_30065,N_27662,N_27753);
or U30066 (N_30066,N_27786,N_29202);
nor U30067 (N_30067,N_28541,N_29737);
nor U30068 (N_30068,N_28510,N_28299);
nand U30069 (N_30069,N_28700,N_28833);
or U30070 (N_30070,N_28695,N_29898);
xor U30071 (N_30071,N_28995,N_28865);
and U30072 (N_30072,N_29566,N_29759);
nor U30073 (N_30073,N_27635,N_28998);
nand U30074 (N_30074,N_28877,N_28024);
and U30075 (N_30075,N_29191,N_29855);
or U30076 (N_30076,N_28268,N_29217);
nor U30077 (N_30077,N_29627,N_28687);
and U30078 (N_30078,N_27844,N_29792);
and U30079 (N_30079,N_29428,N_27670);
or U30080 (N_30080,N_28544,N_29181);
nor U30081 (N_30081,N_29301,N_29868);
xnor U30082 (N_30082,N_29538,N_28957);
and U30083 (N_30083,N_29537,N_28577);
or U30084 (N_30084,N_27717,N_27840);
or U30085 (N_30085,N_29644,N_27895);
and U30086 (N_30086,N_29276,N_29865);
xnor U30087 (N_30087,N_28435,N_28637);
xor U30088 (N_30088,N_28630,N_29862);
nor U30089 (N_30089,N_28973,N_28805);
nor U30090 (N_30090,N_29867,N_28473);
xor U30091 (N_30091,N_29129,N_28273);
or U30092 (N_30092,N_27820,N_28732);
xnor U30093 (N_30093,N_29923,N_28937);
nor U30094 (N_30094,N_28475,N_27585);
or U30095 (N_30095,N_29700,N_28610);
nand U30096 (N_30096,N_28825,N_28744);
nor U30097 (N_30097,N_29422,N_29236);
or U30098 (N_30098,N_29244,N_28055);
or U30099 (N_30099,N_29170,N_29607);
or U30100 (N_30100,N_28275,N_28751);
xor U30101 (N_30101,N_29135,N_29155);
or U30102 (N_30102,N_28168,N_29601);
nor U30103 (N_30103,N_29916,N_27600);
nand U30104 (N_30104,N_29513,N_29444);
or U30105 (N_30105,N_28768,N_29801);
or U30106 (N_30106,N_29549,N_29141);
xnor U30107 (N_30107,N_29251,N_29750);
or U30108 (N_30108,N_29140,N_29766);
nor U30109 (N_30109,N_29972,N_28520);
nand U30110 (N_30110,N_28873,N_27899);
and U30111 (N_30111,N_28536,N_29676);
nand U30112 (N_30112,N_28699,N_27847);
or U30113 (N_30113,N_28439,N_29340);
nand U30114 (N_30114,N_29775,N_28240);
nor U30115 (N_30115,N_28880,N_28708);
nand U30116 (N_30116,N_28802,N_28143);
and U30117 (N_30117,N_28923,N_28760);
or U30118 (N_30118,N_29411,N_28897);
xnor U30119 (N_30119,N_28634,N_29197);
nand U30120 (N_30120,N_29794,N_27835);
nor U30121 (N_30121,N_27602,N_28674);
or U30122 (N_30122,N_28236,N_27733);
nand U30123 (N_30123,N_27738,N_28209);
nand U30124 (N_30124,N_28703,N_28824);
or U30125 (N_30125,N_27902,N_29126);
nor U30126 (N_30126,N_29002,N_28211);
and U30127 (N_30127,N_28583,N_29119);
nand U30128 (N_30128,N_27671,N_29522);
xnor U30129 (N_30129,N_29507,N_29596);
and U30130 (N_30130,N_28898,N_28627);
nand U30131 (N_30131,N_27760,N_27664);
nand U30132 (N_30132,N_28763,N_29568);
nor U30133 (N_30133,N_29738,N_29233);
xnor U30134 (N_30134,N_29001,N_28924);
xor U30135 (N_30135,N_29532,N_28774);
and U30136 (N_30136,N_29316,N_28582);
xor U30137 (N_30137,N_28789,N_27938);
or U30138 (N_30138,N_28887,N_27658);
xnor U30139 (N_30139,N_27526,N_28403);
xor U30140 (N_30140,N_29040,N_27969);
nand U30141 (N_30141,N_27767,N_29345);
and U30142 (N_30142,N_29449,N_27503);
nor U30143 (N_30143,N_28373,N_27621);
and U30144 (N_30144,N_29706,N_28064);
or U30145 (N_30145,N_29719,N_27841);
nor U30146 (N_30146,N_29284,N_28542);
and U30147 (N_30147,N_28538,N_29746);
nor U30148 (N_30148,N_28656,N_28045);
xor U30149 (N_30149,N_27543,N_27742);
xor U30150 (N_30150,N_28607,N_28975);
nand U30151 (N_30151,N_27513,N_29593);
nor U30152 (N_30152,N_27560,N_29803);
nand U30153 (N_30153,N_29866,N_28772);
and U30154 (N_30154,N_29863,N_27505);
nand U30155 (N_30155,N_28007,N_29246);
or U30156 (N_30156,N_28545,N_29039);
xnor U30157 (N_30157,N_29496,N_29368);
xnor U30158 (N_30158,N_29470,N_29090);
and U30159 (N_30159,N_29249,N_28092);
xnor U30160 (N_30160,N_27705,N_29618);
xor U30161 (N_30161,N_27863,N_27925);
nand U30162 (N_30162,N_28586,N_27553);
or U30163 (N_30163,N_27994,N_27606);
nor U30164 (N_30164,N_28256,N_28620);
and U30165 (N_30165,N_27855,N_29531);
nand U30166 (N_30166,N_27577,N_28552);
and U30167 (N_30167,N_28391,N_28228);
or U30168 (N_30168,N_29708,N_27960);
xor U30169 (N_30169,N_28643,N_27952);
xor U30170 (N_30170,N_28886,N_28401);
nor U30171 (N_30171,N_27741,N_28988);
nand U30172 (N_30172,N_29844,N_27620);
nand U30173 (N_30173,N_27548,N_28167);
or U30174 (N_30174,N_29225,N_29843);
or U30175 (N_30175,N_29536,N_28269);
xor U30176 (N_30176,N_29749,N_28863);
xor U30177 (N_30177,N_28931,N_28557);
nor U30178 (N_30178,N_29952,N_29314);
and U30179 (N_30179,N_29200,N_27625);
nor U30180 (N_30180,N_28300,N_27564);
nand U30181 (N_30181,N_27923,N_28008);
or U30182 (N_30182,N_29412,N_27985);
and U30183 (N_30183,N_29572,N_27688);
and U30184 (N_30184,N_28237,N_27580);
or U30185 (N_30185,N_27563,N_29296);
nand U30186 (N_30186,N_27836,N_29027);
and U30187 (N_30187,N_28953,N_28921);
or U30188 (N_30188,N_29059,N_28964);
nor U30189 (N_30189,N_28543,N_29207);
nand U30190 (N_30190,N_28040,N_29189);
or U30191 (N_30191,N_29374,N_29559);
nor U30192 (N_30192,N_27929,N_29208);
nor U30193 (N_30193,N_29034,N_27963);
nand U30194 (N_30194,N_28251,N_29118);
or U30195 (N_30195,N_29905,N_29701);
xnor U30196 (N_30196,N_29655,N_29148);
xor U30197 (N_30197,N_27856,N_27905);
and U30198 (N_30198,N_29430,N_29263);
nand U30199 (N_30199,N_28157,N_29633);
nand U30200 (N_30200,N_28837,N_29180);
nor U30201 (N_30201,N_28290,N_28413);
nand U30202 (N_30202,N_27850,N_28062);
and U30203 (N_30203,N_29343,N_29025);
nand U30204 (N_30204,N_28005,N_29804);
or U30205 (N_30205,N_28407,N_28899);
nor U30206 (N_30206,N_28963,N_28765);
or U30207 (N_30207,N_28486,N_29239);
or U30208 (N_30208,N_28996,N_28481);
and U30209 (N_30209,N_29165,N_28668);
nor U30210 (N_30210,N_27603,N_27608);
nand U30211 (N_30211,N_28793,N_27522);
nand U30212 (N_30212,N_29097,N_29931);
nor U30213 (N_30213,N_28662,N_29290);
nand U30214 (N_30214,N_27615,N_29709);
nand U30215 (N_30215,N_28710,N_28981);
xnor U30216 (N_30216,N_27737,N_29780);
nor U30217 (N_30217,N_29163,N_28685);
and U30218 (N_30218,N_29543,N_28468);
or U30219 (N_30219,N_28362,N_29198);
xnor U30220 (N_30220,N_27907,N_29871);
and U30221 (N_30221,N_27726,N_29159);
xor U30222 (N_30222,N_28239,N_27822);
nor U30223 (N_30223,N_29080,N_29688);
nand U30224 (N_30224,N_27818,N_28212);
or U30225 (N_30225,N_28930,N_28095);
and U30226 (N_30226,N_29283,N_28224);
and U30227 (N_30227,N_29669,N_29098);
nor U30228 (N_30228,N_28462,N_28641);
and U30229 (N_30229,N_28480,N_27695);
xnor U30230 (N_30230,N_27536,N_29014);
and U30231 (N_30231,N_28684,N_29425);
and U30232 (N_30232,N_29611,N_28432);
and U30233 (N_30233,N_28639,N_28799);
and U30234 (N_30234,N_28016,N_28234);
xor U30235 (N_30235,N_29230,N_29557);
xnor U30236 (N_30236,N_27533,N_28631);
nor U30237 (N_30237,N_29015,N_29973);
and U30238 (N_30238,N_27830,N_29819);
or U30239 (N_30239,N_27613,N_28770);
nor U30240 (N_30240,N_29667,N_27906);
or U30241 (N_30241,N_29143,N_29319);
xnor U30242 (N_30242,N_29592,N_29735);
and U30243 (N_30243,N_29854,N_29899);
nand U30244 (N_30244,N_27881,N_28644);
nand U30245 (N_30245,N_27649,N_29282);
xor U30246 (N_30246,N_29499,N_29114);
and U30247 (N_30247,N_29707,N_29448);
nand U30248 (N_30248,N_28404,N_29399);
or U30249 (N_30249,N_29698,N_27768);
and U30250 (N_30250,N_28111,N_28343);
nor U30251 (N_30251,N_27531,N_28215);
and U30252 (N_30252,N_29880,N_29771);
nand U30253 (N_30253,N_28783,N_29182);
nor U30254 (N_30254,N_27552,N_29045);
and U30255 (N_30255,N_28806,N_29711);
xnor U30256 (N_30256,N_29919,N_27675);
or U30257 (N_30257,N_27958,N_28935);
or U30258 (N_30258,N_28585,N_27566);
xnor U30259 (N_30259,N_29394,N_29542);
or U30260 (N_30260,N_28203,N_28498);
and U30261 (N_30261,N_28729,N_28068);
and U30262 (N_30262,N_29881,N_28118);
nor U30263 (N_30263,N_29765,N_27848);
and U30264 (N_30264,N_29602,N_29721);
xor U30265 (N_30265,N_28056,N_28356);
xor U30266 (N_30266,N_28743,N_29320);
xor U30267 (N_30267,N_28222,N_29304);
nand U30268 (N_30268,N_29030,N_28245);
and U30269 (N_30269,N_29156,N_29007);
nor U30270 (N_30270,N_29598,N_28735);
nor U30271 (N_30271,N_29949,N_29049);
xnor U30272 (N_30272,N_28341,N_27607);
and U30273 (N_30273,N_28775,N_28795);
nand U30274 (N_30274,N_29681,N_29190);
xor U30275 (N_30275,N_28028,N_29504);
or U30276 (N_30276,N_27731,N_27727);
nor U30277 (N_30277,N_28123,N_29578);
or U30278 (N_30278,N_29397,N_27891);
nand U30279 (N_30279,N_29875,N_29152);
nand U30280 (N_30280,N_27601,N_28929);
nor U30281 (N_30281,N_28546,N_29616);
xor U30282 (N_30282,N_28658,N_28102);
nor U30283 (N_30283,N_29295,N_29622);
xnor U30284 (N_30284,N_27720,N_29166);
nor U30285 (N_30285,N_29362,N_29396);
nor U30286 (N_30286,N_29584,N_27959);
and U30287 (N_30287,N_27546,N_27551);
xnor U30288 (N_30288,N_28089,N_29378);
xnor U30289 (N_30289,N_29512,N_29255);
and U30290 (N_30290,N_29619,N_29324);
or U30291 (N_30291,N_28612,N_28985);
or U30292 (N_30292,N_28676,N_28002);
or U30293 (N_30293,N_29101,N_28655);
xor U30294 (N_30294,N_28645,N_28214);
or U30295 (N_30295,N_27814,N_29036);
and U30296 (N_30296,N_27624,N_28515);
nor U30297 (N_30297,N_28578,N_27932);
xor U30298 (N_30298,N_27928,N_28826);
and U30299 (N_30299,N_28048,N_28712);
nand U30300 (N_30300,N_28592,N_29951);
nor U30301 (N_30301,N_28364,N_27641);
xor U30302 (N_30302,N_28246,N_29704);
nor U30303 (N_30303,N_27965,N_29267);
nand U30304 (N_30304,N_29408,N_29227);
nand U30305 (N_30305,N_29337,N_28085);
xnor U30306 (N_30306,N_28472,N_27523);
and U30307 (N_30307,N_28411,N_29254);
and U30308 (N_30308,N_28947,N_28130);
nor U30309 (N_30309,N_27696,N_29082);
xor U30310 (N_30310,N_29514,N_29966);
nand U30311 (N_30311,N_27584,N_28315);
nand U30312 (N_30312,N_28421,N_29223);
or U30313 (N_30313,N_28742,N_29414);
xor U30314 (N_30314,N_28459,N_28164);
and U30315 (N_30315,N_28600,N_29278);
or U30316 (N_30316,N_28001,N_28922);
nand U30317 (N_30317,N_29544,N_29778);
xnor U30318 (N_30318,N_29634,N_29248);
nor U30319 (N_30319,N_29398,N_27817);
nand U30320 (N_30320,N_29828,N_29686);
xor U30321 (N_30321,N_27721,N_29084);
nor U30322 (N_30322,N_28372,N_29665);
or U30323 (N_30323,N_28127,N_28116);
nand U30324 (N_30324,N_29471,N_29274);
xor U30325 (N_30325,N_27936,N_28183);
and U30326 (N_30326,N_29438,N_28054);
nor U30327 (N_30327,N_28835,N_28344);
xnor U30328 (N_30328,N_29840,N_28813);
xnor U30329 (N_30329,N_28397,N_29107);
or U30330 (N_30330,N_27622,N_27904);
or U30331 (N_30331,N_27796,N_29974);
or U30332 (N_30332,N_29964,N_28412);
or U30333 (N_30333,N_27964,N_28919);
nand U30334 (N_30334,N_29127,N_28115);
nand U30335 (N_30335,N_27659,N_29436);
or U30336 (N_30336,N_27833,N_28329);
or U30337 (N_30337,N_29710,N_28036);
nor U30338 (N_30338,N_29666,N_29418);
nand U30339 (N_30339,N_28306,N_28944);
nor U30340 (N_30340,N_28145,N_28023);
xnor U30341 (N_30341,N_28406,N_29297);
nor U30342 (N_30342,N_28253,N_29272);
or U30343 (N_30343,N_29954,N_27744);
nor U30344 (N_30344,N_27734,N_29877);
xnor U30345 (N_30345,N_28442,N_29130);
nor U30346 (N_30346,N_29961,N_29960);
or U30347 (N_30347,N_29035,N_27728);
xnor U30348 (N_30348,N_29104,N_28090);
nand U30349 (N_30349,N_29876,N_28954);
nor U30350 (N_30350,N_28946,N_29071);
or U30351 (N_30351,N_29091,N_27980);
nor U30352 (N_30352,N_28476,N_28261);
and U30353 (N_30353,N_29886,N_29756);
and U30354 (N_30354,N_29480,N_29102);
or U30355 (N_30355,N_28279,N_28501);
nand U30356 (N_30356,N_29802,N_28956);
or U30357 (N_30357,N_29564,N_29264);
nor U30358 (N_30358,N_27687,N_29016);
and U30359 (N_30359,N_28354,N_29762);
nor U30360 (N_30360,N_28918,N_27500);
and U30361 (N_30361,N_28017,N_28690);
xor U30362 (N_30362,N_28094,N_28844);
and U30363 (N_30363,N_28086,N_29358);
or U30364 (N_30364,N_28121,N_29705);
or U30365 (N_30365,N_28339,N_29790);
nand U30366 (N_30366,N_28018,N_29033);
and U30367 (N_30367,N_29740,N_27576);
nand U30368 (N_30368,N_28405,N_28642);
or U30369 (N_30369,N_27873,N_29313);
and U30370 (N_30370,N_29921,N_28664);
or U30371 (N_30371,N_29594,N_28888);
nor U30372 (N_30372,N_29702,N_29725);
xnor U30373 (N_30373,N_29475,N_29767);
nor U30374 (N_30374,N_29786,N_28444);
and U30375 (N_30375,N_29253,N_29569);
and U30376 (N_30376,N_27587,N_28349);
nand U30377 (N_30377,N_29585,N_28352);
and U30378 (N_30378,N_27668,N_29716);
xor U30379 (N_30379,N_27669,N_29603);
nand U30380 (N_30380,N_29493,N_29519);
nand U30381 (N_30381,N_28876,N_29257);
or U30382 (N_30382,N_27711,N_28249);
xnor U30383 (N_30383,N_27708,N_28911);
nand U30384 (N_30384,N_29461,N_29506);
xor U30385 (N_30385,N_29534,N_28387);
and U30386 (N_30386,N_27997,N_29987);
nor U30387 (N_30387,N_29630,N_28096);
and U30388 (N_30388,N_27866,N_28626);
xnor U30389 (N_30389,N_28969,N_29694);
nand U30390 (N_30390,N_28181,N_28746);
nand U30391 (N_30391,N_27754,N_29146);
nor U30392 (N_30392,N_28051,N_27698);
xor U30393 (N_30393,N_29347,N_29431);
and U30394 (N_30394,N_29454,N_28519);
or U30395 (N_30395,N_29250,N_29099);
and U30396 (N_30396,N_29648,N_29271);
nand U30397 (N_30397,N_29730,N_29927);
nor U30398 (N_30398,N_27745,N_29144);
xor U30399 (N_30399,N_27865,N_27699);
xnor U30400 (N_30400,N_28323,N_29419);
or U30401 (N_30401,N_29072,N_27795);
xnor U30402 (N_30402,N_28061,N_27530);
xor U30403 (N_30403,N_28031,N_28333);
or U30404 (N_30404,N_27521,N_29747);
and U30405 (N_30405,N_27593,N_27771);
nand U30406 (N_30406,N_29979,N_29901);
nor U30407 (N_30407,N_29367,N_27516);
nor U30408 (N_30408,N_28910,N_29911);
xnor U30409 (N_30409,N_28422,N_28248);
or U30410 (N_30410,N_28526,N_27640);
nor U30411 (N_30411,N_29168,N_28336);
nor U30412 (N_30412,N_27637,N_29020);
xor U30413 (N_30413,N_28595,N_29932);
nand U30414 (N_30414,N_27534,N_27802);
xnor U30415 (N_30415,N_27719,N_29680);
xor U30416 (N_30416,N_29579,N_27581);
nor U30417 (N_30417,N_28893,N_27639);
and U30418 (N_30418,N_28854,N_27686);
and U30419 (N_30419,N_28778,N_28948);
nand U30420 (N_30420,N_27950,N_29024);
nor U30421 (N_30421,N_28338,N_28223);
nor U30422 (N_30422,N_29851,N_28635);
nand U30423 (N_30423,N_29896,N_27931);
nor U30424 (N_30424,N_28894,N_28625);
nor U30425 (N_30425,N_29978,N_29560);
nand U30426 (N_30426,N_28283,N_27901);
nor U30427 (N_30427,N_28896,N_28436);
or U30428 (N_30428,N_28431,N_28026);
nor U30429 (N_30429,N_29293,N_29861);
or U30430 (N_30430,N_29462,N_29713);
nand U30431 (N_30431,N_28414,N_27713);
or U30432 (N_30432,N_27890,N_28129);
nand U30433 (N_30433,N_28126,N_29226);
nand U30434 (N_30434,N_28836,N_28265);
nor U30435 (N_30435,N_28093,N_28158);
and U30436 (N_30436,N_28736,N_28716);
and U30437 (N_30437,N_28153,N_29668);
xor U30438 (N_30438,N_27506,N_29369);
or U30439 (N_30439,N_27643,N_29975);
or U30440 (N_30440,N_28081,N_28616);
and U30441 (N_30441,N_27812,N_27588);
nor U30442 (N_30442,N_29799,N_29820);
and U30443 (N_30443,N_29580,N_28219);
or U30444 (N_30444,N_27599,N_28327);
nand U30445 (N_30445,N_28355,N_28705);
or U30446 (N_30446,N_29968,N_27511);
and U30447 (N_30447,N_27751,N_28989);
xor U30448 (N_30448,N_29077,N_29769);
and U30449 (N_30449,N_28434,N_29908);
xor U30450 (N_30450,N_27646,N_28599);
nand U30451 (N_30451,N_28613,N_29787);
and U30452 (N_30452,N_29069,N_29210);
nand U30453 (N_30453,N_28231,N_27790);
nand U30454 (N_30454,N_29692,N_27594);
or U30455 (N_30455,N_29848,N_29652);
xnor U30456 (N_30456,N_28791,N_27707);
and U30457 (N_30457,N_28322,N_27990);
nor U30458 (N_30458,N_27650,N_29204);
nand U30459 (N_30459,N_27633,N_28576);
nor U30460 (N_30460,N_28866,N_28451);
and U30461 (N_30461,N_29605,N_28313);
and U30462 (N_30462,N_29341,N_28021);
and U30463 (N_30463,N_29539,N_27981);
nand U30464 (N_30464,N_29467,N_27630);
and U30465 (N_30465,N_28810,N_27967);
nor U30466 (N_30466,N_29205,N_29969);
or U30467 (N_30467,N_28319,N_29434);
nand U30468 (N_30468,N_27732,N_28112);
and U30469 (N_30469,N_29745,N_29404);
xor U30470 (N_30470,N_28311,N_29613);
or U30471 (N_30471,N_28015,N_29784);
and U30472 (N_30472,N_29327,N_28977);
xnor U30473 (N_30473,N_28192,N_29946);
and U30474 (N_30474,N_27828,N_27857);
nand U30475 (N_30475,N_29164,N_28326);
xnor U30476 (N_30476,N_28392,N_29595);
xnor U30477 (N_30477,N_29245,N_28289);
nand U30478 (N_30478,N_29505,N_28149);
and U30479 (N_30479,N_28204,N_27806);
or U30480 (N_30480,N_28553,N_29133);
and U30481 (N_30481,N_28220,N_28767);
xnor U30482 (N_30482,N_29895,N_28916);
or U30483 (N_30483,N_27892,N_28408);
nand U30484 (N_30484,N_29375,N_27922);
nand U30485 (N_30485,N_29748,N_28180);
xor U30486 (N_30486,N_28264,N_27704);
nand U30487 (N_30487,N_29715,N_29518);
nor U30488 (N_30488,N_29599,N_29055);
or U30489 (N_30489,N_28649,N_27571);
nand U30490 (N_30490,N_28358,N_29687);
and U30491 (N_30491,N_27740,N_29659);
xnor U30492 (N_30492,N_28505,N_29445);
nand U30493 (N_30493,N_29112,N_28312);
nor U30494 (N_30494,N_29443,N_29209);
nor U30495 (N_30495,N_28380,N_28531);
nor U30496 (N_30496,N_27870,N_29058);
xor U30497 (N_30497,N_29958,N_29703);
and U30498 (N_30498,N_27502,N_29041);
nand U30499 (N_30499,N_29308,N_29902);
nand U30500 (N_30500,N_29883,N_29349);
nand U30501 (N_30501,N_27973,N_29195);
or U30502 (N_30502,N_28900,N_29502);
nor U30503 (N_30503,N_29768,N_29835);
and U30504 (N_30504,N_27852,N_28759);
xor U30505 (N_30505,N_29385,N_29355);
xor U30506 (N_30506,N_29213,N_29169);
xor U30507 (N_30507,N_29528,N_28747);
nand U30508 (N_30508,N_29160,N_27527);
or U30509 (N_30509,N_28208,N_28755);
nor U30510 (N_30510,N_27757,N_28812);
xor U30511 (N_30511,N_28483,N_28560);
nand U30512 (N_30512,N_29829,N_29087);
and U30513 (N_30513,N_29774,N_28571);
xnor U30514 (N_30514,N_29729,N_28337);
or U30515 (N_30515,N_29306,N_28890);
xor U30516 (N_30516,N_28328,N_29458);
xor U30517 (N_30517,N_27893,N_27559);
nand U30518 (N_30518,N_28581,N_28860);
xor U30519 (N_30519,N_28252,N_28217);
and U30520 (N_30520,N_28779,N_27801);
nand U30521 (N_30521,N_28258,N_27871);
and U30522 (N_30522,N_29521,N_27589);
and U30523 (N_30523,N_29473,N_29858);
nand U30524 (N_30524,N_27682,N_28057);
or U30525 (N_30525,N_28991,N_29672);
or U30526 (N_30526,N_29491,N_28623);
nor U30527 (N_30527,N_27896,N_29351);
nand U30528 (N_30528,N_27966,N_28011);
nand U30529 (N_30529,N_29723,N_29022);
nand U30530 (N_30530,N_29309,N_28907);
and U30531 (N_30531,N_28254,N_29573);
or U30532 (N_30532,N_27909,N_28728);
xnor U30533 (N_30533,N_28506,N_28714);
and U30534 (N_30534,N_28309,N_28766);
or U30535 (N_30535,N_28822,N_29553);
nor U30536 (N_30536,N_29487,N_28166);
nand U30537 (N_30537,N_29243,N_28818);
nand U30538 (N_30538,N_28159,N_29452);
nor U30539 (N_30539,N_28452,N_28840);
nand U30540 (N_30540,N_29853,N_27520);
and U30541 (N_30541,N_28065,N_29286);
xor U30542 (N_30542,N_29839,N_28455);
nor U30543 (N_30543,N_28294,N_28663);
or U30544 (N_30544,N_29727,N_27962);
or U30545 (N_30545,N_29137,N_27636);
and U30546 (N_30546,N_27851,N_27677);
or U30547 (N_30547,N_28503,N_27953);
or U30548 (N_30548,N_28385,N_29323);
xnor U30549 (N_30549,N_29864,N_28652);
nand U30550 (N_30550,N_28195,N_28903);
xor U30551 (N_30551,N_29945,N_27679);
and U30552 (N_30552,N_29111,N_28590);
nand U30553 (N_30553,N_27501,N_29891);
and U30554 (N_30554,N_28332,N_28734);
xor U30555 (N_30555,N_28666,N_27842);
xor U30556 (N_30556,N_27776,N_29132);
and U30557 (N_30557,N_29789,N_29407);
and U30558 (N_30558,N_28706,N_27816);
nor U30559 (N_30559,N_29807,N_28572);
xor U30560 (N_30560,N_29201,N_29670);
xor U30561 (N_30561,N_29105,N_28934);
xnor U30562 (N_30562,N_29654,N_28817);
nand U30563 (N_30563,N_28325,N_27702);
and U30564 (N_30564,N_28148,N_29485);
nand U30565 (N_30565,N_29671,N_29031);
xor U30566 (N_30566,N_28282,N_27557);
xor U30567 (N_30567,N_29755,N_27919);
and U30568 (N_30568,N_29312,N_27992);
nand U30569 (N_30569,N_28598,N_27654);
nand U30570 (N_30570,N_28446,N_28816);
nor U30571 (N_30571,N_29696,N_28067);
and U30572 (N_30572,N_27689,N_29393);
nand U30573 (N_30573,N_27946,N_27519);
nor U30574 (N_30574,N_28828,N_29212);
or U30575 (N_30575,N_29224,N_27998);
xnor U30576 (N_30576,N_28041,N_28495);
nand U30577 (N_30577,N_29417,N_28889);
xor U30578 (N_30578,N_27572,N_28295);
xnor U30579 (N_30579,N_28178,N_29268);
nand U30580 (N_30580,N_28073,N_27934);
nand U30581 (N_30581,N_29526,N_27849);
xor U30582 (N_30582,N_29529,N_27718);
and U30583 (N_30583,N_27749,N_29382);
nor U30584 (N_30584,N_29076,N_28076);
and U30585 (N_30585,N_29800,N_29808);
or U30586 (N_30586,N_29996,N_27758);
or U30587 (N_30587,N_28191,N_28491);
nor U30588 (N_30588,N_28570,N_29806);
and U30589 (N_30589,N_28461,N_29456);
xnor U30590 (N_30590,N_27800,N_28188);
and U30591 (N_30591,N_28330,N_27575);
xnor U30592 (N_30592,N_28654,N_29976);
or U30593 (N_30593,N_27547,N_27976);
xor U30594 (N_30594,N_29402,N_28284);
nand U30595 (N_30595,N_28764,N_28811);
or U30596 (N_30596,N_29889,N_29822);
and U30597 (N_30597,N_29812,N_28966);
nor U30598 (N_30598,N_29153,N_28970);
or U30599 (N_30599,N_29693,N_29691);
or U30600 (N_30600,N_28293,N_28858);
or U30601 (N_30601,N_28847,N_28034);
nand U30602 (N_30602,N_28756,N_28901);
nand U30603 (N_30603,N_27592,N_27558);
xor U30604 (N_30604,N_29906,N_29167);
xor U30605 (N_30605,N_28693,N_28917);
nor U30606 (N_30606,N_28740,N_27703);
xor U30607 (N_30607,N_29377,N_27783);
and U30608 (N_30608,N_29825,N_28049);
nor U30609 (N_30609,N_29903,N_29805);
or U30610 (N_30610,N_28565,N_28987);
nor U30611 (N_30611,N_29795,N_29690);
nor U30612 (N_30612,N_29280,N_28952);
and U30613 (N_30613,N_27591,N_29409);
and U30614 (N_30614,N_29904,N_29416);
nand U30615 (N_30615,N_29342,N_27787);
xnor U30616 (N_30616,N_29004,N_29427);
xor U30617 (N_30617,N_29556,N_28942);
xor U30618 (N_30618,N_29477,N_28138);
xnor U30619 (N_30619,N_28474,N_27815);
xnor U30620 (N_30620,N_29277,N_27712);
or U30621 (N_30621,N_28262,N_28874);
nand U30622 (N_30622,N_29956,N_29712);
nor U30623 (N_30623,N_28110,N_29550);
xnor U30624 (N_30624,N_28182,N_29490);
and U30625 (N_30625,N_28580,N_28119);
and U30626 (N_30626,N_28125,N_28723);
or U30627 (N_30627,N_28419,N_28009);
and U30628 (N_30628,N_28241,N_28494);
and U30629 (N_30629,N_28128,N_28790);
xnor U30630 (N_30630,N_28792,N_28402);
nand U30631 (N_30631,N_29934,N_28904);
xor U30632 (N_30632,N_29147,N_29992);
or U30633 (N_30633,N_27597,N_29179);
nand U30634 (N_30634,N_29860,N_28425);
xnor U30635 (N_30635,N_28416,N_29589);
xor U30636 (N_30636,N_29381,N_28808);
nor U30637 (N_30637,N_27517,N_28179);
or U30638 (N_30638,N_29587,N_27644);
xor U30639 (N_30639,N_27540,N_28202);
or U30640 (N_30640,N_29887,N_29517);
nand U30641 (N_30641,N_29128,N_28514);
xnor U30642 (N_30642,N_28861,N_28162);
and U30643 (N_30643,N_27657,N_28060);
or U30644 (N_30644,N_28484,N_29281);
nor U30645 (N_30645,N_27700,N_27550);
or U30646 (N_30646,N_29717,N_29472);
nand U30647 (N_30647,N_29065,N_29600);
and U30648 (N_30648,N_28184,N_28657);
nand U30649 (N_30649,N_29325,N_29846);
and U30650 (N_30650,N_28719,N_27683);
nor U30651 (N_30651,N_28859,N_27568);
nand U30652 (N_30652,N_28177,N_28717);
xnor U30653 (N_30653,N_29731,N_27691);
nor U30654 (N_30654,N_29937,N_27876);
or U30655 (N_30655,N_29917,N_29433);
nor U30656 (N_30656,N_27862,N_28399);
or U30657 (N_30657,N_28787,N_28019);
xor U30658 (N_30658,N_28945,N_27918);
nand U30659 (N_30659,N_28307,N_29009);
nand U30660 (N_30660,N_27629,N_28524);
and U30661 (N_30661,N_29582,N_28424);
nand U30662 (N_30662,N_29890,N_29796);
nor U30663 (N_30663,N_29307,N_28142);
nand U30664 (N_30664,N_27724,N_28718);
and U30665 (N_30665,N_28660,N_28201);
xnor U30666 (N_30666,N_29136,N_29174);
and U30667 (N_30667,N_28618,N_28345);
and U30668 (N_30668,N_27715,N_27555);
nor U30669 (N_30669,N_29983,N_27609);
and U30670 (N_30670,N_29188,N_29561);
nand U30671 (N_30671,N_29240,N_27685);
nor U30672 (N_30672,N_29116,N_28193);
nand U30673 (N_30673,N_28117,N_29360);
xor U30674 (N_30674,N_28568,N_27971);
nand U30675 (N_30675,N_28815,N_27945);
nor U30676 (N_30676,N_28614,N_27570);
xor U30677 (N_30677,N_29085,N_29624);
nor U30678 (N_30678,N_29643,N_28857);
or U30679 (N_30679,N_28784,N_27623);
and U30680 (N_30680,N_29214,N_27773);
or U30681 (N_30681,N_29664,N_28554);
nor U30682 (N_30682,N_27777,N_29797);
nor U30683 (N_30683,N_27747,N_29466);
xor U30684 (N_30684,N_27832,N_29196);
or U30685 (N_30685,N_27886,N_29370);
and U30686 (N_30686,N_27544,N_29366);
and U30687 (N_30687,N_27538,N_28669);
nor U30688 (N_30688,N_29994,N_28410);
and U30689 (N_30689,N_29075,N_28457);
nor U30690 (N_30690,N_28869,N_27549);
nand U30691 (N_30691,N_29056,N_27714);
or U30692 (N_30692,N_28914,N_27746);
nor U30693 (N_30693,N_28780,N_29339);
xor U30694 (N_30694,N_27761,N_27665);
or U30695 (N_30695,N_27821,N_27915);
or U30696 (N_30696,N_29291,N_29158);
xor U30697 (N_30697,N_28502,N_28927);
nand U30698 (N_30698,N_27716,N_28959);
nand U30699 (N_30699,N_29305,N_28689);
nand U30700 (N_30700,N_28423,N_28370);
xor U30701 (N_30701,N_29516,N_28163);
nor U30702 (N_30702,N_28679,N_28605);
nor U30703 (N_30703,N_29231,N_28189);
nand U30704 (N_30704,N_29176,N_29758);
or U30705 (N_30705,N_29123,N_28304);
and U30706 (N_30706,N_28229,N_29720);
or U30707 (N_30707,N_28694,N_29285);
or U30708 (N_30708,N_27739,N_29682);
xnor U30709 (N_30709,N_28567,N_28508);
or U30710 (N_30710,N_28951,N_27867);
nand U30711 (N_30711,N_28575,N_27611);
or U30712 (N_30712,N_28534,N_28681);
or U30713 (N_30713,N_29562,N_29798);
nor U30714 (N_30714,N_29936,N_29053);
or U30715 (N_30715,N_27838,N_27561);
nand U30716 (N_30716,N_27692,N_28692);
nand U30717 (N_30717,N_29483,N_29879);
xnor U30718 (N_30718,N_28075,N_29482);
nand U30719 (N_30719,N_27755,N_28938);
nor U30720 (N_30720,N_28648,N_27752);
nand U30721 (N_30721,N_28277,N_27941);
nor U30722 (N_30722,N_29352,N_28318);
nand U30723 (N_30723,N_29138,N_28939);
or U30724 (N_30724,N_28420,N_27764);
or U30725 (N_30725,N_29508,N_29386);
xnor U30726 (N_30726,N_27595,N_29982);
nand U30727 (N_30727,N_28527,N_28606);
nor U30728 (N_30728,N_27793,N_29203);
nor U30729 (N_30729,N_27676,N_28308);
nor U30730 (N_30730,N_29583,N_29751);
or U30731 (N_30731,N_28518,N_28079);
nand U30732 (N_30732,N_27723,N_29484);
nand U30733 (N_30733,N_28821,N_28673);
nor U30734 (N_30734,N_28324,N_27914);
xnor U30735 (N_30735,N_28650,N_28141);
xnor U30736 (N_30736,N_28776,N_27722);
and U30737 (N_30737,N_29965,N_29615);
and U30738 (N_30738,N_29859,N_29699);
or U30739 (N_30739,N_28107,N_28617);
xnor U30740 (N_30740,N_28549,N_29469);
or U30741 (N_30741,N_28757,N_27791);
or U30742 (N_30742,N_29294,N_27935);
nor U30743 (N_30743,N_29481,N_29199);
nand U30744 (N_30744,N_27653,N_29989);
nand U30745 (N_30745,N_28350,N_27996);
nand U30746 (N_30746,N_28678,N_28335);
and U30747 (N_30747,N_28146,N_28004);
or U30748 (N_30748,N_29446,N_29998);
or U30749 (N_30749,N_28968,N_27628);
xor U30750 (N_30750,N_29151,N_28088);
nor U30751 (N_30751,N_29942,N_28482);
xnor U30752 (N_30752,N_28120,N_29344);
nand U30753 (N_30753,N_29092,N_29008);
or U30754 (N_30754,N_29029,N_28243);
and U30755 (N_30755,N_29938,N_29088);
xor U30756 (N_30756,N_27813,N_29614);
nand U30757 (N_30757,N_29555,N_28653);
and U30758 (N_30758,N_29941,N_28932);
nor U30759 (N_30759,N_29656,N_28449);
xnor U30760 (N_30760,N_29826,N_28843);
nor U30761 (N_30761,N_28247,N_29892);
nand U30762 (N_30762,N_29079,N_28823);
xnor U30763 (N_30763,N_29981,N_27614);
nand U30764 (N_30764,N_28063,N_28724);
xor U30765 (N_30765,N_29554,N_27794);
xnor U30766 (N_30766,N_29995,N_29492);
nor U30767 (N_30767,N_29959,N_27798);
nand U30768 (N_30768,N_28152,N_28371);
xor U30769 (N_30769,N_28207,N_29548);
and U30770 (N_30770,N_28445,N_28033);
nor U30771 (N_30771,N_28758,N_27987);
xor U30772 (N_30772,N_28428,N_28748);
xor U30773 (N_30773,N_27839,N_29586);
nor U30774 (N_30774,N_29157,N_29646);
nor U30775 (N_30775,N_29525,N_29028);
or U30776 (N_30776,N_29384,N_29489);
nand U30777 (N_30777,N_29113,N_29125);
nor U30778 (N_30778,N_29782,N_29171);
or U30779 (N_30779,N_28633,N_28504);
and U30780 (N_30780,N_28539,N_29265);
xor U30781 (N_30781,N_29674,N_29604);
and U30782 (N_30782,N_29632,N_28727);
and U30783 (N_30783,N_27610,N_27663);
or U30784 (N_30784,N_28819,N_29638);
nor U30785 (N_30785,N_29606,N_28165);
nand U30786 (N_30786,N_28522,N_28682);
nand U30787 (N_30787,N_27780,N_28200);
xnor U30788 (N_30788,N_29637,N_28133);
or U30789 (N_30789,N_29259,N_28443);
xnor U30790 (N_30790,N_27535,N_28955);
nor U30791 (N_30791,N_28379,N_27984);
nand U30792 (N_30792,N_28242,N_28559);
nor U30793 (N_30793,N_27778,N_29818);
xor U30794 (N_30794,N_28134,N_28194);
nor U30795 (N_30795,N_29052,N_28171);
and U30796 (N_30796,N_27875,N_27903);
nor U30797 (N_30797,N_28487,N_29777);
nor U30798 (N_30798,N_27983,N_28233);
or U30799 (N_30799,N_29269,N_28376);
and U30800 (N_30800,N_28155,N_28087);
nor U30801 (N_30801,N_27515,N_27660);
nor U30802 (N_30802,N_28082,N_28384);
or U30803 (N_30803,N_28027,N_29520);
xnor U30804 (N_30804,N_28109,N_27961);
nand U30805 (N_30805,N_27933,N_29068);
or U30806 (N_30806,N_29893,N_27937);
or U30807 (N_30807,N_28377,N_29424);
and U30808 (N_30808,N_28038,N_28670);
or U30809 (N_30809,N_28881,N_27541);
nand U30810 (N_30810,N_28564,N_28266);
and U30811 (N_30811,N_28030,N_29635);
nand U30812 (N_30812,N_28078,N_29495);
nand U30813 (N_30813,N_28074,N_28281);
or U30814 (N_30814,N_27859,N_28974);
nor U30815 (N_30815,N_28829,N_28135);
xnor U30816 (N_30816,N_28997,N_27970);
and U30817 (N_30817,N_28892,N_28933);
nand U30818 (N_30818,N_28507,N_27762);
xor U30819 (N_30819,N_28555,N_27887);
or U30820 (N_30820,N_29331,N_28260);
xor U30821 (N_30821,N_29037,N_28750);
nand U30822 (N_30822,N_27939,N_28852);
xnor U30823 (N_30823,N_27883,N_27504);
nand U30824 (N_30824,N_28516,N_29252);
or U30825 (N_30825,N_27735,N_28400);
and U30826 (N_30826,N_29256,N_29432);
and U30827 (N_30827,N_28103,N_29757);
nor U30828 (N_30828,N_28796,N_29064);
nor U30829 (N_30829,N_29641,N_29216);
and U30830 (N_30830,N_29571,N_29261);
xnor U30831 (N_30831,N_28646,N_28794);
nor U30832 (N_30832,N_29662,N_28250);
or U30833 (N_30833,N_29038,N_28137);
xnor U30834 (N_30834,N_29510,N_28885);
nand U30835 (N_30835,N_29161,N_29684);
xnor U30836 (N_30836,N_28677,N_29110);
nor U30837 (N_30837,N_29882,N_27648);
xor U30838 (N_30838,N_27774,N_28285);
or U30839 (N_30839,N_29332,N_29610);
xor U30840 (N_30840,N_27845,N_29728);
xnor U30841 (N_30841,N_27756,N_28636);
and U30842 (N_30842,N_27880,N_29172);
xnor U30843 (N_30843,N_29317,N_28941);
nor U30844 (N_30844,N_29837,N_27514);
nor U30845 (N_30845,N_28418,N_29817);
nand U30846 (N_30846,N_28950,N_29149);
or U30847 (N_30847,N_28070,N_28867);
nor U30848 (N_30848,N_28702,N_29232);
or U30849 (N_30849,N_29591,N_29488);
xor U30850 (N_30850,N_28357,N_27638);
and U30851 (N_30851,N_28346,N_29211);
or U30852 (N_30852,N_29338,N_28593);
or U30853 (N_30853,N_28059,N_28464);
xor U30854 (N_30854,N_28629,N_29103);
xor U30855 (N_30855,N_28925,N_28733);
xnor U30856 (N_30856,N_28458,N_29390);
xnor U30857 (N_30857,N_27975,N_28226);
xnor U30858 (N_30858,N_27674,N_28267);
nor U30859 (N_30859,N_29326,N_29993);
or U30860 (N_30860,N_29726,N_28320);
and U30861 (N_30861,N_29913,N_29884);
or U30862 (N_30862,N_27706,N_28069);
xor U30863 (N_30863,N_27524,N_28072);
nor U30864 (N_30864,N_28039,N_28280);
nor U30865 (N_30865,N_27765,N_28140);
nor U30866 (N_30866,N_28104,N_28291);
xor U30867 (N_30867,N_28053,N_27512);
nor U30868 (N_30868,N_29910,N_29051);
nor U30869 (N_30869,N_29827,N_27770);
or U30870 (N_30870,N_29912,N_28046);
and U30871 (N_30871,N_28651,N_29815);
nor U30872 (N_30872,N_29300,N_28983);
or U30873 (N_30873,N_28800,N_27864);
and U30874 (N_30874,N_27807,N_29026);
and U30875 (N_30875,N_29459,N_28232);
and U30876 (N_30876,N_29310,N_28715);
xnor U30877 (N_30877,N_29732,N_29241);
nor U30878 (N_30878,N_27869,N_29032);
nor U30879 (N_30879,N_27769,N_28499);
nor U30880 (N_30880,N_27710,N_29457);
nor U30881 (N_30881,N_28417,N_29925);
nor U30882 (N_30882,N_28971,N_27618);
nor U30883 (N_30883,N_27565,N_29465);
nand U30884 (N_30884,N_28665,N_28042);
nand U30885 (N_30885,N_28830,N_28196);
xnor U30886 (N_30886,N_27797,N_28013);
nor U30887 (N_30887,N_28122,N_27693);
xor U30888 (N_30888,N_29888,N_28185);
or U30889 (N_30889,N_28389,N_28465);
nor U30890 (N_30890,N_29474,N_29328);
xnor U30891 (N_30891,N_29478,N_28037);
nor U30892 (N_30892,N_29044,N_28225);
xnor U30893 (N_30893,N_28958,N_29131);
or U30894 (N_30894,N_27528,N_29062);
nand U30895 (N_30895,N_27824,N_28632);
nor U30896 (N_30896,N_28701,N_29094);
nand U30897 (N_30897,N_28170,N_29928);
nor U30898 (N_30898,N_28640,N_29830);
and U30899 (N_30899,N_29392,N_29311);
or U30900 (N_30900,N_28360,N_27661);
or U30901 (N_30901,N_28500,N_28883);
nand U30902 (N_30902,N_29183,N_28485);
and U30903 (N_30903,N_29933,N_27854);
nand U30904 (N_30904,N_27562,N_27542);
or U30905 (N_30905,N_28050,N_29546);
xor U30906 (N_30906,N_29383,N_28647);
nor U30907 (N_30907,N_29660,N_28375);
xnor U30908 (N_30908,N_29811,N_27789);
nand U30909 (N_30909,N_27912,N_29924);
nand U30910 (N_30910,N_29793,N_29838);
xnor U30911 (N_30911,N_29547,N_28454);
xnor U30912 (N_30912,N_27968,N_29270);
and U30913 (N_30913,N_28855,N_27612);
nand U30914 (N_30914,N_28334,N_29535);
nor U30915 (N_30915,N_27799,N_27678);
and U30916 (N_30916,N_29845,N_29043);
and U30917 (N_30917,N_27860,N_27872);
or U30918 (N_30918,N_29095,N_29150);
nand U30919 (N_30919,N_29834,N_27921);
and U30920 (N_30920,N_28965,N_27868);
nor U30921 (N_30921,N_29364,N_29718);
nand U30922 (N_30922,N_28244,N_27948);
and U30923 (N_30923,N_28587,N_28535);
and U30924 (N_30924,N_28848,N_29229);
and U30925 (N_30925,N_28569,N_28496);
xnor U30926 (N_30926,N_29184,N_28394);
nand U30927 (N_30927,N_27811,N_29885);
or U30928 (N_30928,N_28390,N_29235);
nor U30929 (N_30929,N_28915,N_27694);
and U30930 (N_30930,N_28761,N_28556);
and U30931 (N_30931,N_28980,N_27743);
nor U30932 (N_30932,N_28845,N_29415);
nor U30933 (N_30933,N_29401,N_29070);
xnor U30934 (N_30934,N_27808,N_28884);
and U30935 (N_30935,N_29997,N_27655);
xnor U30936 (N_30936,N_27725,N_27759);
nand U30937 (N_30937,N_27878,N_28584);
nor U30938 (N_30938,N_29460,N_28749);
nand U30939 (N_30939,N_27632,N_29371);
or U30940 (N_30940,N_29697,N_27647);
and U30941 (N_30941,N_29810,N_28466);
nor U30942 (N_30942,N_27944,N_29142);
nor U30943 (N_30943,N_27879,N_27916);
or U30944 (N_30944,N_28993,N_28551);
nor U30945 (N_30945,N_28426,N_29651);
nor U30946 (N_30946,N_28415,N_27926);
xor U30947 (N_30947,N_28721,N_27858);
and U30948 (N_30948,N_29527,N_28437);
nor U30949 (N_30949,N_27507,N_29673);
nand U30950 (N_30950,N_29194,N_28842);
nand U30951 (N_30951,N_29962,N_29515);
xor U30952 (N_30952,N_28012,N_28943);
nand U30953 (N_30953,N_29266,N_28257);
or U30954 (N_30954,N_29724,N_28259);
nor U30955 (N_30955,N_28000,N_28773);
nand U30956 (N_30956,N_27989,N_29753);
nand U30957 (N_30957,N_29321,N_29922);
and U30958 (N_30958,N_27730,N_27882);
and U30959 (N_30959,N_28713,N_29977);
or U30960 (N_30960,N_29781,N_29953);
nand U30961 (N_30961,N_28611,N_28558);
nor U30962 (N_30962,N_29403,N_28984);
nor U30963 (N_30963,N_29023,N_28305);
nor U30964 (N_30964,N_27993,N_28752);
and U30965 (N_30965,N_28348,N_28479);
nand U30966 (N_30966,N_29260,N_27701);
and U30967 (N_30967,N_29683,N_29856);
or U30968 (N_30968,N_29944,N_29500);
and U30969 (N_30969,N_28533,N_27913);
nand U30970 (N_30970,N_28621,N_27532);
or U30971 (N_30971,N_29005,N_28206);
nor U30972 (N_30972,N_28409,N_28105);
nand U30973 (N_30973,N_29497,N_27578);
nand U30974 (N_30974,N_27656,N_29900);
nor U30975 (N_30975,N_29219,N_28221);
nor U30976 (N_30976,N_29980,N_29626);
and U30977 (N_30977,N_28999,N_27988);
nor U30978 (N_30978,N_27598,N_29760);
or U30979 (N_30979,N_28596,N_28960);
xor U30980 (N_30980,N_29322,N_28174);
and U30981 (N_30981,N_29387,N_28906);
nor U30982 (N_30982,N_27709,N_29074);
nand U30983 (N_30983,N_29948,N_28691);
nor U30984 (N_30984,N_28365,N_27583);
nor U30985 (N_30985,N_29388,N_28872);
or U30986 (N_30986,N_29929,N_28986);
nor U30987 (N_30987,N_29335,N_28374);
nor U30988 (N_30988,N_29741,N_28230);
xnor U30989 (N_30989,N_28709,N_27943);
or U30990 (N_30990,N_28725,N_27518);
and U30991 (N_30991,N_29739,N_28707);
and U30992 (N_30992,N_28139,N_28680);
nand U30993 (N_30993,N_27748,N_28902);
or U30994 (N_30994,N_28878,N_28936);
xor U30995 (N_30995,N_28856,N_28369);
xnor U30996 (N_30996,N_28807,N_27949);
or U30997 (N_30997,N_28227,N_29663);
nand U30998 (N_30998,N_29145,N_28003);
nand U30999 (N_30999,N_28908,N_29363);
xor U31000 (N_31000,N_27785,N_28331);
and U31001 (N_31001,N_29939,N_28827);
nand U31002 (N_31002,N_29356,N_29464);
and U31003 (N_31003,N_29791,N_28278);
xor U31004 (N_31004,N_28493,N_27573);
and U31005 (N_31005,N_29947,N_29776);
nor U31006 (N_31006,N_28785,N_27826);
or U31007 (N_31007,N_28940,N_28263);
xnor U31008 (N_31008,N_28912,N_28722);
or U31009 (N_31009,N_27631,N_27775);
or U31010 (N_31010,N_29783,N_28131);
or U31011 (N_31011,N_29089,N_27605);
nor U31012 (N_31012,N_28920,N_29950);
nand U31013 (N_31013,N_28688,N_28025);
or U31014 (N_31014,N_28467,N_28853);
nor U31015 (N_31015,N_28540,N_28820);
and U31016 (N_31016,N_27954,N_29450);
xnor U31017 (N_31017,N_29503,N_29479);
nand U31018 (N_31018,N_29389,N_29421);
nand U31019 (N_31019,N_29986,N_29653);
nor U31020 (N_31020,N_28302,N_28382);
or U31021 (N_31021,N_27554,N_27947);
or U31022 (N_31022,N_29501,N_28091);
nand U31023 (N_31023,N_29175,N_27525);
and U31024 (N_31024,N_27885,N_28154);
and U31025 (N_31025,N_29742,N_27645);
and U31026 (N_31026,N_29915,N_28525);
nor U31027 (N_31027,N_28754,N_27894);
or U31028 (N_31028,N_27979,N_29850);
or U31029 (N_31029,N_29006,N_28777);
nor U31030 (N_31030,N_29000,N_28741);
and U31031 (N_31031,N_27810,N_28745);
nand U31032 (N_31032,N_29391,N_29570);
nor U31033 (N_31033,N_28686,N_27666);
nand U31034 (N_31034,N_29451,N_27978);
and U31035 (N_31035,N_28297,N_29581);
nor U31036 (N_31036,N_28683,N_28478);
or U31037 (N_31037,N_29833,N_29288);
xnor U31038 (N_31038,N_29315,N_29930);
nor U31039 (N_31039,N_27955,N_27792);
nand U31040 (N_31040,N_29752,N_28450);
xnor U31041 (N_31041,N_28438,N_28697);
nand U31042 (N_31042,N_27819,N_28851);
xor U31043 (N_31043,N_29773,N_28671);
or U31044 (N_31044,N_28044,N_28497);
and U31045 (N_31045,N_29943,N_27596);
xnor U31046 (N_31046,N_29013,N_29551);
nor U31047 (N_31047,N_29847,N_28832);
nor U31048 (N_31048,N_28994,N_29120);
or U31049 (N_31049,N_29545,N_29405);
nor U31050 (N_31050,N_27803,N_29237);
xor U31051 (N_31051,N_28604,N_27888);
and U31052 (N_31052,N_28342,N_29073);
nand U31053 (N_31053,N_28047,N_29441);
nand U31054 (N_31054,N_29247,N_29565);
nand U31055 (N_31055,N_27642,N_29361);
nor U31056 (N_31056,N_29714,N_28704);
nand U31057 (N_31057,N_29139,N_28972);
nand U31058 (N_31058,N_27788,N_28573);
nand U31059 (N_31059,N_28106,N_27942);
and U31060 (N_31060,N_29657,N_28430);
nand U31061 (N_31061,N_29576,N_28603);
or U31062 (N_31062,N_29642,N_28566);
or U31063 (N_31063,N_28753,N_29447);
and U31064 (N_31064,N_27957,N_29857);
and U31065 (N_31065,N_29336,N_28218);
and U31066 (N_31066,N_27634,N_28427);
or U31067 (N_31067,N_29106,N_29353);
xnor U31068 (N_31068,N_29086,N_29621);
nor U31069 (N_31069,N_29010,N_28453);
xnor U31070 (N_31070,N_28469,N_28099);
and U31071 (N_31071,N_28730,N_29287);
nor U31072 (N_31072,N_27690,N_28622);
nand U31073 (N_31073,N_28298,N_29486);
nor U31074 (N_31074,N_29011,N_28737);
xor U31075 (N_31075,N_28804,N_29177);
xor U31076 (N_31076,N_29625,N_29081);
nand U31077 (N_31077,N_29192,N_29754);
nor U31078 (N_31078,N_29530,N_28098);
nor U31079 (N_31079,N_28199,N_27556);
nor U31080 (N_31080,N_29940,N_29494);
and U31081 (N_31081,N_27736,N_27779);
nand U31082 (N_31082,N_29298,N_28786);
or U31083 (N_31083,N_28608,N_29057);
xor U31084 (N_31084,N_27951,N_28809);
or U31085 (N_31085,N_29423,N_29302);
xor U31086 (N_31086,N_29590,N_28463);
nand U31087 (N_31087,N_28321,N_28949);
and U31088 (N_31088,N_29524,N_29350);
xor U31089 (N_31089,N_28798,N_27920);
nand U31090 (N_31090,N_28197,N_29608);
xnor U31091 (N_31091,N_28909,N_28471);
xnor U31092 (N_31092,N_28781,N_28597);
or U31093 (N_31093,N_29955,N_29873);
xor U31094 (N_31094,N_27545,N_28615);
xnor U31095 (N_31095,N_29914,N_28381);
and U31096 (N_31096,N_28288,N_29640);
nor U31097 (N_31097,N_27837,N_28351);
or U31098 (N_31098,N_28198,N_28020);
or U31099 (N_31099,N_29348,N_28547);
xnor U31100 (N_31100,N_27846,N_27917);
and U31101 (N_31101,N_29831,N_28726);
nand U31102 (N_31102,N_28979,N_27781);
and U31103 (N_31103,N_28187,N_29193);
or U31104 (N_31104,N_29379,N_29187);
xnor U31105 (N_31105,N_27652,N_29279);
and U31106 (N_31106,N_29639,N_29836);
nor U31107 (N_31107,N_29957,N_29597);
or U31108 (N_31108,N_28976,N_28296);
and U31109 (N_31109,N_28978,N_29066);
nor U31110 (N_31110,N_28782,N_29429);
nor U31111 (N_31111,N_29650,N_29228);
nand U31112 (N_31112,N_28711,N_27995);
and U31113 (N_31113,N_28771,N_28235);
nor U31114 (N_31114,N_28084,N_29054);
and U31115 (N_31115,N_27537,N_29162);
xnor U31116 (N_31116,N_29764,N_28489);
xor U31117 (N_31117,N_29685,N_29400);
nor U31118 (N_31118,N_28367,N_28961);
nand U31119 (N_31119,N_29511,N_27805);
xor U31120 (N_31120,N_28124,N_28928);
nor U31121 (N_31121,N_29373,N_29734);
and U31122 (N_31122,N_28698,N_28769);
nand U31123 (N_31123,N_28398,N_29426);
or U31124 (N_31124,N_27853,N_28386);
and U31125 (N_31125,N_27897,N_29722);
nor U31126 (N_31126,N_28395,N_29772);
nand U31127 (N_31127,N_29999,N_29292);
nor U31128 (N_31128,N_29647,N_28990);
and U31129 (N_31129,N_28739,N_27930);
nor U31130 (N_31130,N_28136,N_29814);
nor U31131 (N_31131,N_29289,N_27825);
and U31132 (N_31132,N_28440,N_29018);
xor U31133 (N_31133,N_28882,N_27529);
or U31134 (N_31134,N_29221,N_28448);
and U31135 (N_31135,N_28659,N_27766);
or U31136 (N_31136,N_27831,N_28589);
nand U31137 (N_31137,N_29329,N_28310);
xor U31138 (N_31138,N_29649,N_29334);
nor U31139 (N_31139,N_29061,N_28429);
nor U31140 (N_31140,N_28488,N_29019);
or U31141 (N_31141,N_27982,N_29878);
nand U31142 (N_31142,N_27809,N_28396);
and U31143 (N_31143,N_28238,N_29869);
xnor U31144 (N_31144,N_29078,N_29048);
and U31145 (N_31145,N_29821,N_27991);
xor U31146 (N_31146,N_27977,N_29463);
or U31147 (N_31147,N_28006,N_28720);
xor U31148 (N_31148,N_29788,N_28172);
nor U31149 (N_31149,N_29242,N_28316);
nor U31150 (N_31150,N_29991,N_28891);
nor U31151 (N_31151,N_29558,N_28303);
and U31152 (N_31152,N_29376,N_28272);
nor U31153 (N_31153,N_28052,N_28022);
nor U31154 (N_31154,N_27900,N_27567);
nor U31155 (N_31155,N_29357,N_28875);
xnor U31156 (N_31156,N_27898,N_29108);
nor U31157 (N_31157,N_28850,N_29420);
and U31158 (N_31158,N_27697,N_29909);
and U31159 (N_31159,N_29897,N_29689);
or U31160 (N_31160,N_28490,N_28926);
xor U31161 (N_31161,N_29234,N_27508);
and U31162 (N_31162,N_29437,N_29763);
nor U31163 (N_31163,N_28301,N_28523);
nand U31164 (N_31164,N_28077,N_28601);
and U31165 (N_31165,N_28173,N_29410);
and U31166 (N_31166,N_28101,N_29206);
nor U31167 (N_31167,N_29675,N_28864);
nand U31168 (N_31168,N_28441,N_28014);
xor U31169 (N_31169,N_27924,N_29218);
nor U31170 (N_31170,N_29552,N_28151);
nor U31171 (N_31171,N_28638,N_28846);
and U31172 (N_31172,N_29215,N_28276);
nand U31173 (N_31173,N_27974,N_29588);
xor U31174 (N_31174,N_29636,N_28433);
or U31175 (N_31175,N_29985,N_29134);
and U31176 (N_31176,N_29124,N_28393);
xnor U31177 (N_31177,N_28849,N_29096);
nor U31178 (N_31178,N_27782,N_27510);
or U31179 (N_31179,N_29406,N_29083);
xnor U31180 (N_31180,N_28528,N_28213);
or U31181 (N_31181,N_28879,N_29333);
and U31182 (N_31182,N_29823,N_29346);
nor U31183 (N_31183,N_29872,N_28368);
and U31184 (N_31184,N_29628,N_29042);
or U31185 (N_31185,N_28762,N_29761);
or U31186 (N_31186,N_28839,N_28083);
xor U31187 (N_31187,N_27877,N_28361);
and U31188 (N_31188,N_28738,N_28066);
and U31189 (N_31189,N_29907,N_28814);
or U31190 (N_31190,N_29541,N_27874);
nand U31191 (N_31191,N_28513,N_28992);
nand U31192 (N_31192,N_29816,N_27843);
and U31193 (N_31193,N_28032,N_29567);
or U31194 (N_31194,N_29117,N_28529);
xor U31195 (N_31195,N_28512,N_28862);
nor U31196 (N_31196,N_29785,N_28521);
nand U31197 (N_31197,N_27750,N_29238);
nand U31198 (N_31198,N_29733,N_29645);
nor U31199 (N_31199,N_28548,N_28317);
nand U31200 (N_31200,N_29620,N_28803);
and U31201 (N_31201,N_27986,N_29047);
or U31202 (N_31202,N_29012,N_27684);
and U31203 (N_31203,N_28602,N_28477);
or U31204 (N_31204,N_29744,N_27651);
nor U31205 (N_31205,N_29677,N_28871);
nand U31206 (N_31206,N_27574,N_28359);
xor U31207 (N_31207,N_29413,N_29563);
nand U31208 (N_31208,N_28043,N_29678);
xor U31209 (N_31209,N_29109,N_28456);
nor U31210 (N_31210,N_28588,N_29439);
and U31211 (N_31211,N_27539,N_27582);
nor U31212 (N_31212,N_29918,N_27908);
or U31213 (N_31213,N_28210,N_29121);
and U31214 (N_31214,N_28511,N_29533);
and U31215 (N_31215,N_29963,N_28080);
nand U31216 (N_31216,N_28205,N_28870);
and U31217 (N_31217,N_27910,N_28071);
xor U31218 (N_31218,N_27999,N_28834);
xnor U31219 (N_31219,N_28216,N_29609);
nor U31220 (N_31220,N_29658,N_28609);
xnor U31221 (N_31221,N_28114,N_27619);
xnor U31222 (N_31222,N_29173,N_28667);
nor U31223 (N_31223,N_28176,N_27509);
and U31224 (N_31224,N_28274,N_29809);
nand U31225 (N_31225,N_29874,N_27763);
xnor U31226 (N_31226,N_29743,N_29060);
and U31227 (N_31227,N_28460,N_27680);
or U31228 (N_31228,N_29498,N_28562);
xor U31229 (N_31229,N_29540,N_28509);
nand U31230 (N_31230,N_29003,N_27889);
or U31231 (N_31231,N_29273,N_28962);
nor U31232 (N_31232,N_28286,N_29299);
nand U31233 (N_31233,N_27772,N_28353);
nand U31234 (N_31234,N_29523,N_29971);
xor U31235 (N_31235,N_28347,N_28270);
and U31236 (N_31236,N_29779,N_27940);
nor U31237 (N_31237,N_28097,N_28035);
nand U31238 (N_31238,N_28292,N_29695);
nor U31239 (N_31239,N_27673,N_28186);
nor U31240 (N_31240,N_29154,N_29318);
xnor U31241 (N_31241,N_29455,N_27627);
and U31242 (N_31242,N_29186,N_28175);
or U31243 (N_31243,N_29852,N_29842);
and U31244 (N_31244,N_28366,N_28492);
nor U31245 (N_31245,N_29185,N_27626);
xor U31246 (N_31246,N_28563,N_27884);
nor U31247 (N_31247,N_28150,N_27861);
nand U31248 (N_31248,N_29440,N_27617);
nand U31249 (N_31249,N_28058,N_29612);
xnor U31250 (N_31250,N_29224,N_28466);
and U31251 (N_31251,N_28783,N_27501);
and U31252 (N_31252,N_29701,N_27686);
nor U31253 (N_31253,N_27889,N_29910);
or U31254 (N_31254,N_28388,N_29180);
nand U31255 (N_31255,N_29421,N_28455);
xor U31256 (N_31256,N_29575,N_28026);
nand U31257 (N_31257,N_28585,N_29606);
and U31258 (N_31258,N_27986,N_29901);
xnor U31259 (N_31259,N_29370,N_29746);
and U31260 (N_31260,N_28241,N_29297);
xor U31261 (N_31261,N_28311,N_28630);
and U31262 (N_31262,N_28888,N_29437);
xnor U31263 (N_31263,N_29912,N_28845);
nand U31264 (N_31264,N_29980,N_29446);
and U31265 (N_31265,N_28238,N_29505);
xnor U31266 (N_31266,N_29082,N_29711);
or U31267 (N_31267,N_29589,N_27833);
xnor U31268 (N_31268,N_29372,N_28138);
nand U31269 (N_31269,N_29033,N_27718);
xor U31270 (N_31270,N_29411,N_29198);
xnor U31271 (N_31271,N_28612,N_27692);
and U31272 (N_31272,N_27586,N_28823);
nand U31273 (N_31273,N_29179,N_28466);
nand U31274 (N_31274,N_28795,N_28955);
and U31275 (N_31275,N_29303,N_28972);
and U31276 (N_31276,N_29751,N_29230);
and U31277 (N_31277,N_27879,N_28234);
nor U31278 (N_31278,N_29890,N_27868);
nand U31279 (N_31279,N_27872,N_29192);
nor U31280 (N_31280,N_28190,N_29634);
nand U31281 (N_31281,N_29891,N_29863);
nand U31282 (N_31282,N_29621,N_29386);
xor U31283 (N_31283,N_28431,N_28726);
or U31284 (N_31284,N_27779,N_27994);
nand U31285 (N_31285,N_29375,N_29028);
nand U31286 (N_31286,N_28717,N_28311);
nand U31287 (N_31287,N_28855,N_29696);
xnor U31288 (N_31288,N_29386,N_28897);
and U31289 (N_31289,N_27669,N_27899);
nand U31290 (N_31290,N_28405,N_29314);
nor U31291 (N_31291,N_27713,N_27894);
nor U31292 (N_31292,N_27572,N_28570);
or U31293 (N_31293,N_29926,N_27892);
nand U31294 (N_31294,N_27936,N_27509);
nor U31295 (N_31295,N_28635,N_29986);
and U31296 (N_31296,N_28200,N_28973);
nand U31297 (N_31297,N_27784,N_29330);
nor U31298 (N_31298,N_28415,N_27624);
xnor U31299 (N_31299,N_27546,N_27802);
nand U31300 (N_31300,N_27975,N_27834);
or U31301 (N_31301,N_28212,N_27646);
xnor U31302 (N_31302,N_28160,N_28818);
xnor U31303 (N_31303,N_29754,N_28446);
nor U31304 (N_31304,N_28016,N_28641);
xor U31305 (N_31305,N_29125,N_29130);
nor U31306 (N_31306,N_29993,N_29689);
or U31307 (N_31307,N_28520,N_28155);
nor U31308 (N_31308,N_29659,N_29916);
and U31309 (N_31309,N_27528,N_27986);
and U31310 (N_31310,N_29959,N_27855);
xnor U31311 (N_31311,N_27970,N_29750);
nand U31312 (N_31312,N_28291,N_28625);
or U31313 (N_31313,N_28155,N_27561);
nand U31314 (N_31314,N_28124,N_29363);
and U31315 (N_31315,N_28286,N_29235);
xor U31316 (N_31316,N_29051,N_29583);
xnor U31317 (N_31317,N_29671,N_28158);
nor U31318 (N_31318,N_27797,N_28316);
and U31319 (N_31319,N_29839,N_27683);
nor U31320 (N_31320,N_28519,N_29107);
nor U31321 (N_31321,N_27766,N_27531);
xnor U31322 (N_31322,N_28609,N_29127);
xnor U31323 (N_31323,N_29094,N_28216);
nor U31324 (N_31324,N_29528,N_28254);
nor U31325 (N_31325,N_28725,N_28255);
and U31326 (N_31326,N_28151,N_29484);
nand U31327 (N_31327,N_28047,N_27830);
nand U31328 (N_31328,N_29192,N_28391);
nor U31329 (N_31329,N_28752,N_28288);
or U31330 (N_31330,N_29717,N_29946);
nor U31331 (N_31331,N_29065,N_29548);
or U31332 (N_31332,N_29236,N_27688);
and U31333 (N_31333,N_28226,N_28349);
nand U31334 (N_31334,N_28008,N_27508);
xor U31335 (N_31335,N_27823,N_28489);
or U31336 (N_31336,N_28680,N_28532);
nor U31337 (N_31337,N_29621,N_27649);
xnor U31338 (N_31338,N_28699,N_28380);
nor U31339 (N_31339,N_29617,N_28088);
nand U31340 (N_31340,N_28832,N_29884);
or U31341 (N_31341,N_28927,N_29986);
nor U31342 (N_31342,N_28682,N_28179);
and U31343 (N_31343,N_29448,N_28892);
xnor U31344 (N_31344,N_29755,N_29368);
xor U31345 (N_31345,N_27537,N_29570);
nor U31346 (N_31346,N_29080,N_29694);
xor U31347 (N_31347,N_27644,N_28352);
or U31348 (N_31348,N_28892,N_29777);
or U31349 (N_31349,N_28163,N_27721);
nor U31350 (N_31350,N_28599,N_28736);
xor U31351 (N_31351,N_29521,N_28727);
nand U31352 (N_31352,N_29916,N_28673);
and U31353 (N_31353,N_27816,N_28945);
and U31354 (N_31354,N_28841,N_27622);
nand U31355 (N_31355,N_28983,N_29614);
nand U31356 (N_31356,N_29145,N_27903);
nand U31357 (N_31357,N_28544,N_27790);
or U31358 (N_31358,N_27634,N_29649);
and U31359 (N_31359,N_28318,N_28793);
xnor U31360 (N_31360,N_27759,N_28169);
nor U31361 (N_31361,N_28122,N_28483);
or U31362 (N_31362,N_27873,N_29433);
or U31363 (N_31363,N_29148,N_29335);
or U31364 (N_31364,N_29326,N_27511);
and U31365 (N_31365,N_27568,N_29370);
and U31366 (N_31366,N_27899,N_28024);
nor U31367 (N_31367,N_29548,N_29729);
or U31368 (N_31368,N_29794,N_28783);
or U31369 (N_31369,N_28914,N_28915);
and U31370 (N_31370,N_28711,N_29337);
and U31371 (N_31371,N_29728,N_29084);
nor U31372 (N_31372,N_28252,N_29389);
nand U31373 (N_31373,N_28613,N_29602);
or U31374 (N_31374,N_28082,N_29210);
and U31375 (N_31375,N_27520,N_27929);
or U31376 (N_31376,N_28134,N_29835);
or U31377 (N_31377,N_29002,N_28456);
or U31378 (N_31378,N_27961,N_28714);
nor U31379 (N_31379,N_29334,N_28033);
nand U31380 (N_31380,N_28679,N_29591);
or U31381 (N_31381,N_28687,N_28174);
and U31382 (N_31382,N_28016,N_28546);
xor U31383 (N_31383,N_29610,N_29629);
xnor U31384 (N_31384,N_28480,N_29272);
nor U31385 (N_31385,N_27710,N_28839);
nand U31386 (N_31386,N_29065,N_29228);
nand U31387 (N_31387,N_27548,N_27756);
nand U31388 (N_31388,N_28146,N_27744);
or U31389 (N_31389,N_29793,N_29049);
nor U31390 (N_31390,N_27817,N_27643);
xnor U31391 (N_31391,N_28105,N_29533);
xnor U31392 (N_31392,N_28695,N_28626);
and U31393 (N_31393,N_29169,N_29098);
nand U31394 (N_31394,N_27697,N_28048);
xor U31395 (N_31395,N_29900,N_28781);
nor U31396 (N_31396,N_27963,N_28824);
or U31397 (N_31397,N_27921,N_29867);
and U31398 (N_31398,N_28320,N_28742);
xnor U31399 (N_31399,N_28342,N_28539);
nand U31400 (N_31400,N_28387,N_29595);
nor U31401 (N_31401,N_28688,N_29586);
and U31402 (N_31402,N_29342,N_27959);
xor U31403 (N_31403,N_29761,N_27584);
xnor U31404 (N_31404,N_29430,N_28283);
or U31405 (N_31405,N_28848,N_29728);
or U31406 (N_31406,N_28691,N_29290);
nor U31407 (N_31407,N_29667,N_28330);
and U31408 (N_31408,N_28076,N_29306);
nor U31409 (N_31409,N_29033,N_29263);
or U31410 (N_31410,N_29819,N_29015);
xor U31411 (N_31411,N_27688,N_27598);
and U31412 (N_31412,N_27597,N_28697);
nor U31413 (N_31413,N_28249,N_28646);
or U31414 (N_31414,N_29899,N_27580);
or U31415 (N_31415,N_27835,N_28952);
xnor U31416 (N_31416,N_28007,N_29529);
nand U31417 (N_31417,N_28722,N_27803);
or U31418 (N_31418,N_29131,N_28026);
nand U31419 (N_31419,N_29759,N_29935);
xnor U31420 (N_31420,N_28940,N_27676);
and U31421 (N_31421,N_28500,N_29579);
nor U31422 (N_31422,N_29550,N_27549);
nand U31423 (N_31423,N_29345,N_29677);
nor U31424 (N_31424,N_27844,N_28260);
nand U31425 (N_31425,N_27959,N_28352);
nand U31426 (N_31426,N_28167,N_29121);
and U31427 (N_31427,N_28370,N_27921);
nand U31428 (N_31428,N_27939,N_29165);
or U31429 (N_31429,N_27887,N_27581);
xnor U31430 (N_31430,N_29175,N_28167);
and U31431 (N_31431,N_29978,N_28959);
nor U31432 (N_31432,N_29067,N_28507);
nand U31433 (N_31433,N_29931,N_28987);
xnor U31434 (N_31434,N_28151,N_29309);
and U31435 (N_31435,N_27913,N_28558);
xor U31436 (N_31436,N_29375,N_29378);
nor U31437 (N_31437,N_28646,N_28869);
nand U31438 (N_31438,N_27813,N_28086);
nor U31439 (N_31439,N_29128,N_29517);
nand U31440 (N_31440,N_29878,N_29073);
and U31441 (N_31441,N_29193,N_27763);
nand U31442 (N_31442,N_27837,N_27861);
xnor U31443 (N_31443,N_28547,N_27532);
nor U31444 (N_31444,N_27835,N_28979);
and U31445 (N_31445,N_28493,N_29833);
nand U31446 (N_31446,N_29747,N_28590);
or U31447 (N_31447,N_29697,N_27696);
nor U31448 (N_31448,N_28465,N_29238);
nor U31449 (N_31449,N_28214,N_29883);
and U31450 (N_31450,N_29813,N_27548);
and U31451 (N_31451,N_29732,N_28202);
nor U31452 (N_31452,N_28763,N_28592);
nor U31453 (N_31453,N_29945,N_29553);
and U31454 (N_31454,N_28634,N_29867);
nor U31455 (N_31455,N_27926,N_28132);
nor U31456 (N_31456,N_29448,N_29509);
nand U31457 (N_31457,N_27673,N_28238);
nand U31458 (N_31458,N_28962,N_28852);
nand U31459 (N_31459,N_29915,N_28247);
nand U31460 (N_31460,N_27575,N_28336);
and U31461 (N_31461,N_29695,N_28789);
nor U31462 (N_31462,N_28775,N_29041);
xnor U31463 (N_31463,N_28613,N_29051);
and U31464 (N_31464,N_27669,N_28274);
nor U31465 (N_31465,N_29286,N_27979);
and U31466 (N_31466,N_29850,N_29333);
or U31467 (N_31467,N_28944,N_28872);
nor U31468 (N_31468,N_29487,N_29411);
nor U31469 (N_31469,N_29215,N_28578);
or U31470 (N_31470,N_28258,N_29629);
xor U31471 (N_31471,N_28621,N_29656);
or U31472 (N_31472,N_28781,N_29870);
nand U31473 (N_31473,N_27931,N_29266);
nand U31474 (N_31474,N_28482,N_28179);
or U31475 (N_31475,N_27874,N_29931);
or U31476 (N_31476,N_28134,N_27529);
xor U31477 (N_31477,N_28412,N_29209);
nand U31478 (N_31478,N_29078,N_29673);
nor U31479 (N_31479,N_27912,N_28732);
xor U31480 (N_31480,N_28421,N_29728);
nand U31481 (N_31481,N_28421,N_29257);
xnor U31482 (N_31482,N_28255,N_29589);
nor U31483 (N_31483,N_29520,N_27899);
or U31484 (N_31484,N_28687,N_29990);
or U31485 (N_31485,N_29491,N_28189);
nand U31486 (N_31486,N_29656,N_29979);
nand U31487 (N_31487,N_27938,N_27971);
nand U31488 (N_31488,N_29947,N_28403);
xnor U31489 (N_31489,N_28224,N_27810);
or U31490 (N_31490,N_28489,N_28822);
nor U31491 (N_31491,N_29973,N_29448);
xnor U31492 (N_31492,N_28260,N_28986);
or U31493 (N_31493,N_27851,N_27521);
nand U31494 (N_31494,N_27598,N_29586);
and U31495 (N_31495,N_29784,N_28585);
xor U31496 (N_31496,N_28581,N_29961);
xor U31497 (N_31497,N_28693,N_28904);
and U31498 (N_31498,N_29476,N_28285);
nor U31499 (N_31499,N_27776,N_29253);
nand U31500 (N_31500,N_27866,N_29063);
and U31501 (N_31501,N_28826,N_29203);
nor U31502 (N_31502,N_28991,N_27680);
xor U31503 (N_31503,N_29836,N_27759);
xor U31504 (N_31504,N_28446,N_28288);
xor U31505 (N_31505,N_29538,N_29188);
xor U31506 (N_31506,N_29232,N_27908);
and U31507 (N_31507,N_28230,N_29641);
and U31508 (N_31508,N_29642,N_28259);
nand U31509 (N_31509,N_29797,N_29560);
or U31510 (N_31510,N_28401,N_28801);
nand U31511 (N_31511,N_27702,N_27601);
or U31512 (N_31512,N_27791,N_28594);
xor U31513 (N_31513,N_27905,N_27875);
xnor U31514 (N_31514,N_28175,N_29316);
and U31515 (N_31515,N_28406,N_27501);
nor U31516 (N_31516,N_29421,N_27725);
or U31517 (N_31517,N_27900,N_29864);
nand U31518 (N_31518,N_27828,N_29701);
xor U31519 (N_31519,N_27512,N_27856);
nand U31520 (N_31520,N_29623,N_29691);
nand U31521 (N_31521,N_27767,N_28800);
nor U31522 (N_31522,N_29763,N_29621);
nor U31523 (N_31523,N_29847,N_29350);
nand U31524 (N_31524,N_28264,N_27676);
and U31525 (N_31525,N_29024,N_28672);
nand U31526 (N_31526,N_29344,N_29196);
nor U31527 (N_31527,N_29998,N_28346);
nor U31528 (N_31528,N_28543,N_27700);
or U31529 (N_31529,N_29236,N_28590);
nor U31530 (N_31530,N_29303,N_28528);
nand U31531 (N_31531,N_29541,N_29613);
xor U31532 (N_31532,N_28880,N_28502);
or U31533 (N_31533,N_28511,N_27872);
xnor U31534 (N_31534,N_29848,N_29862);
and U31535 (N_31535,N_28105,N_28936);
and U31536 (N_31536,N_28237,N_28076);
xor U31537 (N_31537,N_29656,N_29939);
or U31538 (N_31538,N_29284,N_28008);
nor U31539 (N_31539,N_29140,N_29583);
nand U31540 (N_31540,N_27530,N_29951);
xor U31541 (N_31541,N_28267,N_28418);
xor U31542 (N_31542,N_28622,N_29425);
nand U31543 (N_31543,N_28839,N_29916);
nor U31544 (N_31544,N_27869,N_28985);
xor U31545 (N_31545,N_28714,N_28093);
nor U31546 (N_31546,N_28673,N_28649);
nand U31547 (N_31547,N_28367,N_28900);
nor U31548 (N_31548,N_28248,N_28012);
xor U31549 (N_31549,N_27597,N_29835);
nor U31550 (N_31550,N_28319,N_27985);
nand U31551 (N_31551,N_28078,N_29992);
or U31552 (N_31552,N_29312,N_28269);
nand U31553 (N_31553,N_29652,N_29266);
xor U31554 (N_31554,N_27979,N_27515);
nand U31555 (N_31555,N_28748,N_29802);
nand U31556 (N_31556,N_29478,N_29822);
and U31557 (N_31557,N_29098,N_28015);
or U31558 (N_31558,N_28035,N_27989);
or U31559 (N_31559,N_28738,N_27766);
or U31560 (N_31560,N_28911,N_27789);
nor U31561 (N_31561,N_28544,N_28343);
xnor U31562 (N_31562,N_27740,N_29493);
and U31563 (N_31563,N_27883,N_28632);
nand U31564 (N_31564,N_27859,N_27604);
or U31565 (N_31565,N_28716,N_29188);
nand U31566 (N_31566,N_27882,N_27998);
nand U31567 (N_31567,N_28630,N_28274);
nor U31568 (N_31568,N_28037,N_29495);
and U31569 (N_31569,N_29810,N_28011);
nand U31570 (N_31570,N_28525,N_29877);
xor U31571 (N_31571,N_29668,N_28357);
nor U31572 (N_31572,N_28823,N_29324);
nand U31573 (N_31573,N_29608,N_28927);
nand U31574 (N_31574,N_29116,N_27583);
nor U31575 (N_31575,N_28531,N_29062);
xnor U31576 (N_31576,N_27685,N_29204);
nor U31577 (N_31577,N_27837,N_28970);
and U31578 (N_31578,N_28300,N_27695);
and U31579 (N_31579,N_28184,N_29268);
nand U31580 (N_31580,N_29073,N_27910);
xnor U31581 (N_31581,N_27694,N_27542);
nand U31582 (N_31582,N_29858,N_29965);
nand U31583 (N_31583,N_28560,N_28270);
and U31584 (N_31584,N_28679,N_27765);
nand U31585 (N_31585,N_28458,N_28931);
xor U31586 (N_31586,N_28390,N_29007);
nor U31587 (N_31587,N_28244,N_29370);
xnor U31588 (N_31588,N_27772,N_28757);
xor U31589 (N_31589,N_27644,N_29636);
xor U31590 (N_31590,N_29307,N_28879);
and U31591 (N_31591,N_28417,N_27564);
or U31592 (N_31592,N_28132,N_28884);
nor U31593 (N_31593,N_29336,N_28841);
xnor U31594 (N_31594,N_29952,N_29917);
nor U31595 (N_31595,N_28663,N_29857);
xnor U31596 (N_31596,N_28213,N_28652);
or U31597 (N_31597,N_28548,N_28169);
and U31598 (N_31598,N_28796,N_29229);
or U31599 (N_31599,N_29234,N_28712);
or U31600 (N_31600,N_28555,N_28711);
nand U31601 (N_31601,N_27952,N_27778);
nor U31602 (N_31602,N_28261,N_28355);
or U31603 (N_31603,N_28035,N_29115);
nor U31604 (N_31604,N_28137,N_28219);
or U31605 (N_31605,N_28713,N_29250);
and U31606 (N_31606,N_29377,N_29615);
nand U31607 (N_31607,N_29571,N_28624);
and U31608 (N_31608,N_28883,N_29911);
xor U31609 (N_31609,N_28770,N_28542);
or U31610 (N_31610,N_28711,N_29655);
and U31611 (N_31611,N_29827,N_29815);
or U31612 (N_31612,N_28620,N_27756);
and U31613 (N_31613,N_28756,N_28673);
xnor U31614 (N_31614,N_29019,N_29976);
nand U31615 (N_31615,N_29775,N_28447);
nand U31616 (N_31616,N_28761,N_28409);
and U31617 (N_31617,N_29303,N_27708);
nor U31618 (N_31618,N_29792,N_29143);
xnor U31619 (N_31619,N_28986,N_28102);
or U31620 (N_31620,N_28345,N_29492);
and U31621 (N_31621,N_29667,N_28611);
nor U31622 (N_31622,N_29503,N_27666);
nor U31623 (N_31623,N_28786,N_28129);
nand U31624 (N_31624,N_28174,N_29618);
xor U31625 (N_31625,N_27768,N_28306);
or U31626 (N_31626,N_28544,N_27903);
or U31627 (N_31627,N_27820,N_29271);
nor U31628 (N_31628,N_29101,N_29002);
or U31629 (N_31629,N_28687,N_29660);
nand U31630 (N_31630,N_27643,N_29597);
or U31631 (N_31631,N_28070,N_28019);
or U31632 (N_31632,N_27933,N_28789);
or U31633 (N_31633,N_29651,N_28181);
nor U31634 (N_31634,N_29255,N_29235);
xor U31635 (N_31635,N_28186,N_27581);
xor U31636 (N_31636,N_29567,N_28782);
or U31637 (N_31637,N_28823,N_28775);
xor U31638 (N_31638,N_28655,N_28665);
or U31639 (N_31639,N_29570,N_27569);
or U31640 (N_31640,N_28687,N_29290);
or U31641 (N_31641,N_29438,N_28532);
or U31642 (N_31642,N_28682,N_27758);
and U31643 (N_31643,N_29769,N_29245);
xor U31644 (N_31644,N_27702,N_29160);
or U31645 (N_31645,N_29680,N_28137);
xnor U31646 (N_31646,N_28300,N_29868);
nor U31647 (N_31647,N_28106,N_29384);
xnor U31648 (N_31648,N_29404,N_28475);
xor U31649 (N_31649,N_27715,N_29546);
nor U31650 (N_31650,N_28442,N_28029);
nor U31651 (N_31651,N_29402,N_27901);
nor U31652 (N_31652,N_28116,N_27537);
nand U31653 (N_31653,N_27563,N_29042);
or U31654 (N_31654,N_28130,N_28917);
xor U31655 (N_31655,N_29935,N_29969);
nand U31656 (N_31656,N_29615,N_27564);
nor U31657 (N_31657,N_28925,N_28222);
nor U31658 (N_31658,N_27740,N_29390);
xnor U31659 (N_31659,N_29934,N_29314);
or U31660 (N_31660,N_29284,N_29638);
nor U31661 (N_31661,N_28552,N_29390);
and U31662 (N_31662,N_29998,N_29105);
or U31663 (N_31663,N_29052,N_29515);
and U31664 (N_31664,N_27623,N_28996);
nand U31665 (N_31665,N_28408,N_28538);
and U31666 (N_31666,N_27563,N_27765);
nand U31667 (N_31667,N_29519,N_29797);
xnor U31668 (N_31668,N_29959,N_29354);
nor U31669 (N_31669,N_28794,N_28919);
xnor U31670 (N_31670,N_29296,N_29494);
nor U31671 (N_31671,N_29853,N_28623);
nand U31672 (N_31672,N_27877,N_29252);
nor U31673 (N_31673,N_29537,N_29568);
nor U31674 (N_31674,N_29912,N_28115);
or U31675 (N_31675,N_29101,N_29434);
and U31676 (N_31676,N_29576,N_27571);
nand U31677 (N_31677,N_29959,N_29569);
xnor U31678 (N_31678,N_29015,N_27818);
nand U31679 (N_31679,N_28228,N_27775);
nor U31680 (N_31680,N_29056,N_27923);
or U31681 (N_31681,N_27669,N_29715);
and U31682 (N_31682,N_28357,N_29458);
nor U31683 (N_31683,N_29417,N_29860);
nor U31684 (N_31684,N_29161,N_29861);
and U31685 (N_31685,N_28906,N_29989);
nor U31686 (N_31686,N_27922,N_28954);
nor U31687 (N_31687,N_28714,N_29516);
xnor U31688 (N_31688,N_28166,N_27681);
and U31689 (N_31689,N_28054,N_28818);
nor U31690 (N_31690,N_27639,N_28978);
and U31691 (N_31691,N_28869,N_27646);
nor U31692 (N_31692,N_29164,N_27981);
nand U31693 (N_31693,N_28942,N_29639);
and U31694 (N_31694,N_28362,N_27812);
nor U31695 (N_31695,N_28683,N_27988);
and U31696 (N_31696,N_29999,N_28917);
or U31697 (N_31697,N_28369,N_28555);
nor U31698 (N_31698,N_29497,N_27967);
xnor U31699 (N_31699,N_28656,N_28197);
nor U31700 (N_31700,N_29488,N_28065);
xor U31701 (N_31701,N_27804,N_29053);
xnor U31702 (N_31702,N_28440,N_28041);
and U31703 (N_31703,N_28887,N_27770);
and U31704 (N_31704,N_29669,N_29222);
and U31705 (N_31705,N_29414,N_28887);
nand U31706 (N_31706,N_27874,N_29350);
or U31707 (N_31707,N_27634,N_27589);
xnor U31708 (N_31708,N_29395,N_29165);
nor U31709 (N_31709,N_29927,N_27767);
xnor U31710 (N_31710,N_28341,N_29041);
nand U31711 (N_31711,N_28810,N_27996);
nand U31712 (N_31712,N_28763,N_28705);
nand U31713 (N_31713,N_29125,N_29044);
or U31714 (N_31714,N_27622,N_28767);
nor U31715 (N_31715,N_29760,N_28528);
or U31716 (N_31716,N_29106,N_29866);
nor U31717 (N_31717,N_27798,N_27715);
xor U31718 (N_31718,N_29135,N_28988);
xor U31719 (N_31719,N_27795,N_29395);
nor U31720 (N_31720,N_28831,N_27816);
and U31721 (N_31721,N_28215,N_28457);
or U31722 (N_31722,N_28476,N_28086);
nand U31723 (N_31723,N_28508,N_29655);
xnor U31724 (N_31724,N_28946,N_28305);
or U31725 (N_31725,N_28236,N_28207);
xor U31726 (N_31726,N_29196,N_28588);
and U31727 (N_31727,N_27503,N_28052);
xnor U31728 (N_31728,N_28444,N_29957);
nand U31729 (N_31729,N_28687,N_28464);
nand U31730 (N_31730,N_29791,N_29291);
xor U31731 (N_31731,N_28668,N_27696);
or U31732 (N_31732,N_28037,N_29353);
xnor U31733 (N_31733,N_28045,N_28081);
nand U31734 (N_31734,N_29274,N_28301);
or U31735 (N_31735,N_28031,N_29029);
nand U31736 (N_31736,N_28166,N_29707);
nor U31737 (N_31737,N_29373,N_28766);
nor U31738 (N_31738,N_27965,N_28882);
and U31739 (N_31739,N_27707,N_28889);
xor U31740 (N_31740,N_29417,N_27825);
nand U31741 (N_31741,N_27794,N_29866);
or U31742 (N_31742,N_29518,N_29914);
nand U31743 (N_31743,N_29738,N_28964);
nand U31744 (N_31744,N_29927,N_27722);
xor U31745 (N_31745,N_28128,N_29948);
or U31746 (N_31746,N_29969,N_28790);
xnor U31747 (N_31747,N_29447,N_29117);
and U31748 (N_31748,N_29010,N_28548);
and U31749 (N_31749,N_29876,N_29764);
or U31750 (N_31750,N_28063,N_29661);
xor U31751 (N_31751,N_28067,N_28617);
nand U31752 (N_31752,N_29973,N_29831);
and U31753 (N_31753,N_28994,N_29846);
and U31754 (N_31754,N_29782,N_29005);
xnor U31755 (N_31755,N_29883,N_29036);
and U31756 (N_31756,N_29304,N_29272);
nor U31757 (N_31757,N_29100,N_27545);
nor U31758 (N_31758,N_29939,N_28943);
xnor U31759 (N_31759,N_29630,N_28158);
nor U31760 (N_31760,N_29407,N_28756);
xnor U31761 (N_31761,N_28078,N_28262);
or U31762 (N_31762,N_28310,N_29404);
nand U31763 (N_31763,N_28443,N_29635);
nand U31764 (N_31764,N_28449,N_27698);
xnor U31765 (N_31765,N_28990,N_29701);
and U31766 (N_31766,N_28492,N_28819);
nor U31767 (N_31767,N_29426,N_29055);
or U31768 (N_31768,N_29379,N_29161);
or U31769 (N_31769,N_28047,N_28365);
and U31770 (N_31770,N_28195,N_27694);
and U31771 (N_31771,N_28012,N_29379);
xnor U31772 (N_31772,N_28846,N_28319);
or U31773 (N_31773,N_28479,N_28419);
nand U31774 (N_31774,N_28412,N_28388);
xnor U31775 (N_31775,N_28284,N_29248);
nand U31776 (N_31776,N_28394,N_29419);
nand U31777 (N_31777,N_27587,N_28893);
or U31778 (N_31778,N_28867,N_29464);
nor U31779 (N_31779,N_28146,N_29337);
and U31780 (N_31780,N_27733,N_28265);
and U31781 (N_31781,N_28868,N_27881);
or U31782 (N_31782,N_29160,N_29395);
nand U31783 (N_31783,N_27678,N_29709);
nand U31784 (N_31784,N_29099,N_28552);
nand U31785 (N_31785,N_28061,N_28014);
nand U31786 (N_31786,N_27533,N_29666);
xnor U31787 (N_31787,N_27567,N_29355);
xnor U31788 (N_31788,N_29085,N_28718);
nand U31789 (N_31789,N_29364,N_27719);
nor U31790 (N_31790,N_28108,N_27893);
xnor U31791 (N_31791,N_28995,N_29367);
and U31792 (N_31792,N_28377,N_28770);
xnor U31793 (N_31793,N_27567,N_29838);
xnor U31794 (N_31794,N_27833,N_28200);
and U31795 (N_31795,N_27755,N_28591);
or U31796 (N_31796,N_29176,N_29574);
nand U31797 (N_31797,N_28166,N_28712);
nor U31798 (N_31798,N_28843,N_28507);
or U31799 (N_31799,N_28468,N_28974);
nor U31800 (N_31800,N_29625,N_29443);
or U31801 (N_31801,N_29224,N_29689);
nand U31802 (N_31802,N_27743,N_29558);
xnor U31803 (N_31803,N_28774,N_29774);
or U31804 (N_31804,N_28530,N_28425);
nor U31805 (N_31805,N_28287,N_28245);
nand U31806 (N_31806,N_28256,N_29063);
or U31807 (N_31807,N_28058,N_28875);
or U31808 (N_31808,N_29809,N_29292);
nor U31809 (N_31809,N_29384,N_28150);
or U31810 (N_31810,N_29600,N_27659);
nand U31811 (N_31811,N_27911,N_28559);
and U31812 (N_31812,N_28010,N_29139);
xor U31813 (N_31813,N_29916,N_29167);
and U31814 (N_31814,N_27690,N_29470);
and U31815 (N_31815,N_29894,N_28143);
and U31816 (N_31816,N_28612,N_28114);
or U31817 (N_31817,N_28376,N_28929);
nor U31818 (N_31818,N_27985,N_29622);
nor U31819 (N_31819,N_28166,N_28121);
nor U31820 (N_31820,N_27560,N_29753);
nor U31821 (N_31821,N_28011,N_29255);
nor U31822 (N_31822,N_29625,N_29927);
nand U31823 (N_31823,N_28990,N_29287);
nor U31824 (N_31824,N_28211,N_28822);
nand U31825 (N_31825,N_27769,N_29387);
xor U31826 (N_31826,N_29391,N_28552);
nor U31827 (N_31827,N_28741,N_28262);
or U31828 (N_31828,N_28111,N_28400);
nor U31829 (N_31829,N_28411,N_29523);
or U31830 (N_31830,N_29333,N_27756);
nand U31831 (N_31831,N_29523,N_27530);
and U31832 (N_31832,N_28701,N_28950);
xor U31833 (N_31833,N_29015,N_29602);
xor U31834 (N_31834,N_28246,N_29173);
nand U31835 (N_31835,N_27613,N_28167);
xor U31836 (N_31836,N_29925,N_28926);
nand U31837 (N_31837,N_27761,N_28721);
and U31838 (N_31838,N_29677,N_29820);
nand U31839 (N_31839,N_27516,N_29152);
nor U31840 (N_31840,N_29150,N_29829);
or U31841 (N_31841,N_28040,N_28072);
nand U31842 (N_31842,N_27942,N_28170);
xor U31843 (N_31843,N_29273,N_28412);
or U31844 (N_31844,N_27722,N_28188);
and U31845 (N_31845,N_28321,N_28813);
and U31846 (N_31846,N_29180,N_28155);
and U31847 (N_31847,N_28325,N_29141);
nor U31848 (N_31848,N_28588,N_28333);
or U31849 (N_31849,N_29581,N_29176);
nand U31850 (N_31850,N_28648,N_28551);
or U31851 (N_31851,N_28628,N_28799);
or U31852 (N_31852,N_27972,N_29472);
xnor U31853 (N_31853,N_29187,N_28245);
or U31854 (N_31854,N_28572,N_28047);
or U31855 (N_31855,N_29046,N_27586);
and U31856 (N_31856,N_29167,N_27775);
xnor U31857 (N_31857,N_27889,N_28910);
and U31858 (N_31858,N_29372,N_29861);
nand U31859 (N_31859,N_29983,N_27708);
nor U31860 (N_31860,N_29893,N_29286);
nor U31861 (N_31861,N_29585,N_28272);
nand U31862 (N_31862,N_29499,N_29503);
and U31863 (N_31863,N_29552,N_29465);
nand U31864 (N_31864,N_28437,N_27539);
nor U31865 (N_31865,N_28065,N_28445);
or U31866 (N_31866,N_28819,N_28065);
or U31867 (N_31867,N_29529,N_27703);
and U31868 (N_31868,N_29214,N_29487);
xor U31869 (N_31869,N_29759,N_28000);
and U31870 (N_31870,N_28423,N_29678);
nand U31871 (N_31871,N_28297,N_27887);
xor U31872 (N_31872,N_28009,N_29558);
xnor U31873 (N_31873,N_29075,N_29053);
nand U31874 (N_31874,N_28090,N_28782);
nor U31875 (N_31875,N_29465,N_28347);
nor U31876 (N_31876,N_28805,N_29950);
xnor U31877 (N_31877,N_28147,N_28752);
nor U31878 (N_31878,N_29511,N_29993);
nand U31879 (N_31879,N_28900,N_29712);
nand U31880 (N_31880,N_28778,N_29507);
nand U31881 (N_31881,N_28648,N_28967);
nor U31882 (N_31882,N_28333,N_29654);
nor U31883 (N_31883,N_28544,N_29553);
xnor U31884 (N_31884,N_27649,N_29064);
nor U31885 (N_31885,N_29176,N_27944);
and U31886 (N_31886,N_28226,N_28094);
and U31887 (N_31887,N_29040,N_28076);
nor U31888 (N_31888,N_29066,N_28833);
xnor U31889 (N_31889,N_29495,N_28535);
or U31890 (N_31890,N_28262,N_29270);
xnor U31891 (N_31891,N_29069,N_28465);
or U31892 (N_31892,N_29920,N_28226);
or U31893 (N_31893,N_28548,N_27757);
and U31894 (N_31894,N_28868,N_28669);
nor U31895 (N_31895,N_27738,N_28286);
nor U31896 (N_31896,N_27903,N_28597);
and U31897 (N_31897,N_28351,N_28083);
xnor U31898 (N_31898,N_28727,N_28566);
nand U31899 (N_31899,N_29692,N_27696);
xnor U31900 (N_31900,N_27514,N_29847);
and U31901 (N_31901,N_28976,N_27501);
xor U31902 (N_31902,N_29897,N_29274);
and U31903 (N_31903,N_28164,N_28747);
nor U31904 (N_31904,N_29339,N_29832);
or U31905 (N_31905,N_29836,N_27757);
and U31906 (N_31906,N_29566,N_29252);
xnor U31907 (N_31907,N_29348,N_29977);
or U31908 (N_31908,N_29827,N_29324);
or U31909 (N_31909,N_27895,N_28227);
nand U31910 (N_31910,N_29652,N_28877);
or U31911 (N_31911,N_28671,N_29969);
and U31912 (N_31912,N_27503,N_29903);
nand U31913 (N_31913,N_27765,N_29065);
or U31914 (N_31914,N_29160,N_27983);
nor U31915 (N_31915,N_29308,N_28510);
nor U31916 (N_31916,N_27970,N_29532);
and U31917 (N_31917,N_27921,N_29033);
nor U31918 (N_31918,N_27537,N_28202);
nand U31919 (N_31919,N_27914,N_27606);
nor U31920 (N_31920,N_29093,N_28254);
or U31921 (N_31921,N_28949,N_28402);
nand U31922 (N_31922,N_29109,N_28648);
nor U31923 (N_31923,N_28719,N_28771);
xnor U31924 (N_31924,N_29783,N_28741);
nor U31925 (N_31925,N_28394,N_28583);
nand U31926 (N_31926,N_28967,N_28733);
nor U31927 (N_31927,N_28925,N_28237);
nor U31928 (N_31928,N_29148,N_28047);
xor U31929 (N_31929,N_28112,N_28084);
nor U31930 (N_31930,N_29649,N_28781);
nand U31931 (N_31931,N_27638,N_29707);
and U31932 (N_31932,N_29665,N_27820);
and U31933 (N_31933,N_29342,N_28111);
and U31934 (N_31934,N_28433,N_28695);
and U31935 (N_31935,N_28739,N_29168);
and U31936 (N_31936,N_28821,N_27996);
and U31937 (N_31937,N_28527,N_28085);
nor U31938 (N_31938,N_28170,N_28112);
and U31939 (N_31939,N_27821,N_29877);
xnor U31940 (N_31940,N_28561,N_28107);
xor U31941 (N_31941,N_28825,N_29745);
nand U31942 (N_31942,N_28517,N_29142);
xnor U31943 (N_31943,N_28405,N_28907);
nand U31944 (N_31944,N_29204,N_29564);
and U31945 (N_31945,N_27830,N_28870);
nand U31946 (N_31946,N_27621,N_29484);
and U31947 (N_31947,N_28489,N_27543);
xnor U31948 (N_31948,N_29840,N_28055);
xor U31949 (N_31949,N_29959,N_28922);
xnor U31950 (N_31950,N_27998,N_29015);
nand U31951 (N_31951,N_29927,N_29828);
and U31952 (N_31952,N_27704,N_29879);
nor U31953 (N_31953,N_28558,N_28315);
or U31954 (N_31954,N_29430,N_28926);
xor U31955 (N_31955,N_27944,N_29572);
nand U31956 (N_31956,N_29444,N_28757);
nor U31957 (N_31957,N_28239,N_29880);
and U31958 (N_31958,N_29673,N_28473);
xnor U31959 (N_31959,N_27957,N_28117);
nor U31960 (N_31960,N_27606,N_29973);
nand U31961 (N_31961,N_29209,N_28117);
nor U31962 (N_31962,N_29001,N_27627);
or U31963 (N_31963,N_27977,N_27593);
nor U31964 (N_31964,N_27783,N_29774);
and U31965 (N_31965,N_28873,N_27894);
or U31966 (N_31966,N_27825,N_29116);
nand U31967 (N_31967,N_28891,N_29329);
nand U31968 (N_31968,N_28047,N_28580);
and U31969 (N_31969,N_28441,N_28636);
nor U31970 (N_31970,N_27861,N_28101);
and U31971 (N_31971,N_28197,N_29539);
or U31972 (N_31972,N_29710,N_28620);
or U31973 (N_31973,N_28643,N_27800);
nor U31974 (N_31974,N_28693,N_27742);
nand U31975 (N_31975,N_28292,N_27990);
xnor U31976 (N_31976,N_28131,N_29414);
nand U31977 (N_31977,N_28840,N_29948);
and U31978 (N_31978,N_27864,N_29917);
nor U31979 (N_31979,N_29490,N_28567);
nand U31980 (N_31980,N_28735,N_28126);
or U31981 (N_31981,N_28713,N_28127);
and U31982 (N_31982,N_29108,N_28100);
and U31983 (N_31983,N_29487,N_29191);
or U31984 (N_31984,N_29345,N_27904);
nand U31985 (N_31985,N_28610,N_27624);
and U31986 (N_31986,N_27991,N_28138);
nor U31987 (N_31987,N_28676,N_29757);
or U31988 (N_31988,N_29685,N_29087);
nand U31989 (N_31989,N_29454,N_29619);
nor U31990 (N_31990,N_27689,N_28172);
or U31991 (N_31991,N_27743,N_28857);
nand U31992 (N_31992,N_29478,N_29960);
xor U31993 (N_31993,N_29360,N_28475);
nor U31994 (N_31994,N_29492,N_28160);
xnor U31995 (N_31995,N_27851,N_29326);
nand U31996 (N_31996,N_28806,N_29963);
xnor U31997 (N_31997,N_27836,N_28270);
or U31998 (N_31998,N_29052,N_28997);
xnor U31999 (N_31999,N_27747,N_28716);
nor U32000 (N_32000,N_28112,N_28283);
nor U32001 (N_32001,N_29683,N_29896);
or U32002 (N_32002,N_28465,N_28660);
and U32003 (N_32003,N_29542,N_29164);
nand U32004 (N_32004,N_28178,N_29835);
nor U32005 (N_32005,N_28703,N_28153);
or U32006 (N_32006,N_27771,N_28755);
nor U32007 (N_32007,N_29272,N_27626);
or U32008 (N_32008,N_27672,N_29488);
xor U32009 (N_32009,N_29412,N_27611);
nor U32010 (N_32010,N_28089,N_29748);
nor U32011 (N_32011,N_27501,N_28657);
nor U32012 (N_32012,N_28839,N_29120);
nand U32013 (N_32013,N_27857,N_28750);
nor U32014 (N_32014,N_27820,N_29378);
and U32015 (N_32015,N_29727,N_27882);
nor U32016 (N_32016,N_28077,N_27754);
nand U32017 (N_32017,N_27956,N_29007);
nor U32018 (N_32018,N_29810,N_27782);
or U32019 (N_32019,N_28168,N_29947);
or U32020 (N_32020,N_27821,N_29505);
nor U32021 (N_32021,N_28912,N_28574);
and U32022 (N_32022,N_27969,N_29112);
nor U32023 (N_32023,N_29914,N_29444);
xnor U32024 (N_32024,N_28784,N_28414);
and U32025 (N_32025,N_28407,N_28663);
and U32026 (N_32026,N_27841,N_27757);
or U32027 (N_32027,N_29414,N_29622);
nor U32028 (N_32028,N_28442,N_29289);
nand U32029 (N_32029,N_29097,N_27948);
nand U32030 (N_32030,N_27729,N_27824);
and U32031 (N_32031,N_28436,N_29441);
and U32032 (N_32032,N_28344,N_29860);
nor U32033 (N_32033,N_29322,N_29097);
xor U32034 (N_32034,N_29279,N_27846);
and U32035 (N_32035,N_28703,N_29829);
or U32036 (N_32036,N_28259,N_29005);
nand U32037 (N_32037,N_28696,N_29054);
nand U32038 (N_32038,N_28203,N_29370);
nand U32039 (N_32039,N_29578,N_28130);
nor U32040 (N_32040,N_28710,N_28966);
nand U32041 (N_32041,N_28715,N_27797);
xor U32042 (N_32042,N_27706,N_29197);
and U32043 (N_32043,N_29315,N_29778);
nor U32044 (N_32044,N_29042,N_27861);
and U32045 (N_32045,N_27726,N_29374);
nand U32046 (N_32046,N_28187,N_29497);
xnor U32047 (N_32047,N_29818,N_28088);
and U32048 (N_32048,N_29899,N_28523);
or U32049 (N_32049,N_29233,N_29489);
nor U32050 (N_32050,N_27961,N_29637);
nor U32051 (N_32051,N_27965,N_28890);
and U32052 (N_32052,N_28881,N_29849);
xnor U32053 (N_32053,N_28723,N_29795);
nor U32054 (N_32054,N_28110,N_28946);
and U32055 (N_32055,N_27550,N_28984);
nand U32056 (N_32056,N_28822,N_29357);
nor U32057 (N_32057,N_29257,N_27867);
nand U32058 (N_32058,N_28449,N_27824);
xnor U32059 (N_32059,N_29963,N_28898);
nor U32060 (N_32060,N_27563,N_29071);
nand U32061 (N_32061,N_27773,N_27869);
and U32062 (N_32062,N_29405,N_29788);
nand U32063 (N_32063,N_28750,N_28621);
or U32064 (N_32064,N_29469,N_28666);
xor U32065 (N_32065,N_28129,N_27636);
or U32066 (N_32066,N_28541,N_27501);
or U32067 (N_32067,N_28144,N_27958);
and U32068 (N_32068,N_27650,N_29166);
xor U32069 (N_32069,N_27759,N_28234);
xnor U32070 (N_32070,N_27888,N_28688);
or U32071 (N_32071,N_29199,N_29672);
and U32072 (N_32072,N_29538,N_28391);
nand U32073 (N_32073,N_28379,N_29431);
nor U32074 (N_32074,N_29102,N_28115);
xnor U32075 (N_32075,N_27809,N_28468);
xor U32076 (N_32076,N_27705,N_28857);
nor U32077 (N_32077,N_28280,N_28769);
xor U32078 (N_32078,N_28284,N_27863);
nor U32079 (N_32079,N_28860,N_28700);
or U32080 (N_32080,N_28055,N_29811);
and U32081 (N_32081,N_29512,N_28731);
xnor U32082 (N_32082,N_28191,N_29321);
nand U32083 (N_32083,N_28270,N_27788);
nand U32084 (N_32084,N_27606,N_29229);
xnor U32085 (N_32085,N_29983,N_28159);
nor U32086 (N_32086,N_27568,N_28840);
and U32087 (N_32087,N_29074,N_29785);
or U32088 (N_32088,N_29145,N_29373);
nand U32089 (N_32089,N_28314,N_28131);
nor U32090 (N_32090,N_28511,N_28084);
xnor U32091 (N_32091,N_29306,N_29087);
and U32092 (N_32092,N_28050,N_27677);
xor U32093 (N_32093,N_28830,N_29398);
nand U32094 (N_32094,N_27865,N_29286);
or U32095 (N_32095,N_28705,N_28401);
and U32096 (N_32096,N_29765,N_29753);
nand U32097 (N_32097,N_27851,N_27896);
nand U32098 (N_32098,N_29333,N_29813);
xor U32099 (N_32099,N_28632,N_29931);
nor U32100 (N_32100,N_28095,N_28716);
and U32101 (N_32101,N_28962,N_28276);
nand U32102 (N_32102,N_27545,N_29438);
xor U32103 (N_32103,N_28801,N_29857);
and U32104 (N_32104,N_28545,N_29037);
and U32105 (N_32105,N_28231,N_29761);
nor U32106 (N_32106,N_29818,N_28225);
or U32107 (N_32107,N_28777,N_29963);
nor U32108 (N_32108,N_29726,N_29809);
nand U32109 (N_32109,N_29882,N_29200);
and U32110 (N_32110,N_29481,N_29949);
and U32111 (N_32111,N_27591,N_28336);
nor U32112 (N_32112,N_28127,N_29369);
xor U32113 (N_32113,N_29700,N_28690);
nand U32114 (N_32114,N_27993,N_29290);
xor U32115 (N_32115,N_28075,N_27974);
and U32116 (N_32116,N_27907,N_29631);
or U32117 (N_32117,N_27794,N_28866);
and U32118 (N_32118,N_29198,N_27581);
nor U32119 (N_32119,N_29005,N_27711);
and U32120 (N_32120,N_29200,N_29926);
and U32121 (N_32121,N_29713,N_28661);
or U32122 (N_32122,N_27931,N_28333);
or U32123 (N_32123,N_27558,N_28946);
or U32124 (N_32124,N_29137,N_28807);
xnor U32125 (N_32125,N_28631,N_28552);
nand U32126 (N_32126,N_29713,N_29311);
xor U32127 (N_32127,N_29927,N_28180);
nand U32128 (N_32128,N_29171,N_29393);
nor U32129 (N_32129,N_28733,N_28116);
nand U32130 (N_32130,N_27629,N_29728);
xnor U32131 (N_32131,N_29836,N_27874);
xor U32132 (N_32132,N_28115,N_27510);
and U32133 (N_32133,N_27895,N_27614);
and U32134 (N_32134,N_27741,N_29368);
xnor U32135 (N_32135,N_28492,N_28137);
nand U32136 (N_32136,N_28456,N_29594);
xor U32137 (N_32137,N_29666,N_29381);
nor U32138 (N_32138,N_28901,N_29291);
nor U32139 (N_32139,N_28079,N_28054);
and U32140 (N_32140,N_28533,N_28287);
and U32141 (N_32141,N_27937,N_29234);
xor U32142 (N_32142,N_29117,N_28437);
or U32143 (N_32143,N_29393,N_28330);
and U32144 (N_32144,N_27519,N_29913);
and U32145 (N_32145,N_29511,N_28693);
or U32146 (N_32146,N_28692,N_28933);
and U32147 (N_32147,N_29608,N_29730);
or U32148 (N_32148,N_28980,N_29564);
xnor U32149 (N_32149,N_29799,N_29240);
and U32150 (N_32150,N_29557,N_28880);
and U32151 (N_32151,N_28052,N_28062);
or U32152 (N_32152,N_28753,N_29772);
and U32153 (N_32153,N_29550,N_29299);
or U32154 (N_32154,N_29248,N_28909);
or U32155 (N_32155,N_29063,N_27980);
or U32156 (N_32156,N_28498,N_29996);
or U32157 (N_32157,N_29948,N_28216);
and U32158 (N_32158,N_29921,N_27647);
nand U32159 (N_32159,N_28472,N_28073);
or U32160 (N_32160,N_28789,N_27752);
nand U32161 (N_32161,N_29660,N_29902);
or U32162 (N_32162,N_29883,N_27800);
nand U32163 (N_32163,N_27970,N_28899);
nor U32164 (N_32164,N_28953,N_29578);
and U32165 (N_32165,N_28133,N_28982);
nor U32166 (N_32166,N_27820,N_28542);
nand U32167 (N_32167,N_28443,N_29477);
xor U32168 (N_32168,N_29971,N_28706);
or U32169 (N_32169,N_28827,N_28857);
or U32170 (N_32170,N_27757,N_28806);
nand U32171 (N_32171,N_28578,N_27640);
xnor U32172 (N_32172,N_29749,N_28419);
and U32173 (N_32173,N_28973,N_29298);
xor U32174 (N_32174,N_28229,N_28462);
and U32175 (N_32175,N_28307,N_27500);
nor U32176 (N_32176,N_27624,N_28598);
or U32177 (N_32177,N_29097,N_28687);
and U32178 (N_32178,N_29139,N_27946);
nand U32179 (N_32179,N_28338,N_28778);
or U32180 (N_32180,N_28421,N_28565);
nor U32181 (N_32181,N_29327,N_29132);
and U32182 (N_32182,N_28865,N_28520);
nor U32183 (N_32183,N_29182,N_29229);
and U32184 (N_32184,N_28651,N_29467);
and U32185 (N_32185,N_29922,N_28765);
or U32186 (N_32186,N_29322,N_28277);
or U32187 (N_32187,N_27685,N_29129);
xor U32188 (N_32188,N_29534,N_27946);
or U32189 (N_32189,N_28796,N_29182);
xor U32190 (N_32190,N_27830,N_27938);
nor U32191 (N_32191,N_28015,N_28461);
or U32192 (N_32192,N_28355,N_29842);
nor U32193 (N_32193,N_29688,N_29813);
xnor U32194 (N_32194,N_29906,N_27964);
and U32195 (N_32195,N_28117,N_28662);
and U32196 (N_32196,N_28744,N_29795);
nand U32197 (N_32197,N_27990,N_27839);
nand U32198 (N_32198,N_28193,N_28545);
or U32199 (N_32199,N_28829,N_28871);
or U32200 (N_32200,N_27820,N_28972);
xnor U32201 (N_32201,N_27763,N_27596);
or U32202 (N_32202,N_29295,N_28661);
or U32203 (N_32203,N_29001,N_28644);
nand U32204 (N_32204,N_27775,N_29826);
or U32205 (N_32205,N_27603,N_29690);
nor U32206 (N_32206,N_28932,N_28828);
or U32207 (N_32207,N_29869,N_29066);
xor U32208 (N_32208,N_29332,N_27946);
xor U32209 (N_32209,N_27782,N_29211);
xnor U32210 (N_32210,N_29219,N_28725);
nor U32211 (N_32211,N_28926,N_29347);
or U32212 (N_32212,N_29606,N_29889);
or U32213 (N_32213,N_28263,N_28268);
and U32214 (N_32214,N_27993,N_27843);
nand U32215 (N_32215,N_29697,N_28375);
nor U32216 (N_32216,N_28412,N_28435);
and U32217 (N_32217,N_29513,N_28962);
nand U32218 (N_32218,N_29882,N_27688);
or U32219 (N_32219,N_29009,N_28012);
xnor U32220 (N_32220,N_28674,N_28873);
and U32221 (N_32221,N_29402,N_27717);
or U32222 (N_32222,N_29822,N_27787);
nor U32223 (N_32223,N_29009,N_28338);
nor U32224 (N_32224,N_27742,N_27806);
and U32225 (N_32225,N_28320,N_27841);
nand U32226 (N_32226,N_27765,N_27739);
nor U32227 (N_32227,N_27932,N_28446);
nand U32228 (N_32228,N_27516,N_28017);
and U32229 (N_32229,N_29441,N_28986);
nor U32230 (N_32230,N_28290,N_28679);
nand U32231 (N_32231,N_27553,N_29602);
nand U32232 (N_32232,N_27563,N_29329);
xnor U32233 (N_32233,N_27678,N_29731);
nand U32234 (N_32234,N_28571,N_29172);
or U32235 (N_32235,N_28582,N_29197);
xor U32236 (N_32236,N_28596,N_29142);
or U32237 (N_32237,N_29798,N_29968);
or U32238 (N_32238,N_27881,N_28018);
or U32239 (N_32239,N_28725,N_29358);
or U32240 (N_32240,N_27823,N_28924);
nor U32241 (N_32241,N_27916,N_29090);
or U32242 (N_32242,N_29023,N_29782);
xor U32243 (N_32243,N_28946,N_28557);
xnor U32244 (N_32244,N_29140,N_28196);
nand U32245 (N_32245,N_28249,N_28321);
and U32246 (N_32246,N_29045,N_29020);
or U32247 (N_32247,N_28485,N_28372);
xor U32248 (N_32248,N_29782,N_29914);
and U32249 (N_32249,N_27576,N_29189);
nand U32250 (N_32250,N_28000,N_28096);
xnor U32251 (N_32251,N_27898,N_28424);
or U32252 (N_32252,N_28463,N_28717);
xnor U32253 (N_32253,N_29580,N_28138);
xnor U32254 (N_32254,N_29919,N_29201);
nor U32255 (N_32255,N_28146,N_29232);
nand U32256 (N_32256,N_28055,N_28537);
nand U32257 (N_32257,N_28238,N_27983);
nand U32258 (N_32258,N_28792,N_29912);
nand U32259 (N_32259,N_27696,N_29637);
xor U32260 (N_32260,N_28010,N_27729);
nand U32261 (N_32261,N_29092,N_29894);
or U32262 (N_32262,N_29064,N_29306);
and U32263 (N_32263,N_28971,N_28973);
nand U32264 (N_32264,N_28019,N_28619);
xor U32265 (N_32265,N_28080,N_29203);
and U32266 (N_32266,N_27778,N_28086);
xnor U32267 (N_32267,N_28720,N_27546);
xnor U32268 (N_32268,N_27677,N_29310);
and U32269 (N_32269,N_29509,N_29419);
or U32270 (N_32270,N_27975,N_28023);
and U32271 (N_32271,N_29273,N_29709);
nor U32272 (N_32272,N_28090,N_29160);
and U32273 (N_32273,N_29248,N_29102);
or U32274 (N_32274,N_27949,N_28352);
or U32275 (N_32275,N_27719,N_29097);
nand U32276 (N_32276,N_27735,N_29444);
nand U32277 (N_32277,N_29834,N_28302);
and U32278 (N_32278,N_28357,N_29985);
or U32279 (N_32279,N_27959,N_28214);
nor U32280 (N_32280,N_28730,N_29016);
or U32281 (N_32281,N_27573,N_27999);
xor U32282 (N_32282,N_28738,N_28057);
xor U32283 (N_32283,N_29149,N_29847);
nand U32284 (N_32284,N_29110,N_28244);
nor U32285 (N_32285,N_29074,N_28554);
xnor U32286 (N_32286,N_29286,N_28497);
nor U32287 (N_32287,N_29323,N_29766);
nor U32288 (N_32288,N_28281,N_28814);
xnor U32289 (N_32289,N_28177,N_28108);
nand U32290 (N_32290,N_27874,N_29147);
nand U32291 (N_32291,N_29256,N_29931);
xor U32292 (N_32292,N_28582,N_29145);
nor U32293 (N_32293,N_28121,N_29868);
nand U32294 (N_32294,N_27501,N_28139);
and U32295 (N_32295,N_27952,N_29427);
or U32296 (N_32296,N_28139,N_28918);
xor U32297 (N_32297,N_28057,N_27909);
or U32298 (N_32298,N_28630,N_29463);
or U32299 (N_32299,N_29042,N_28618);
nor U32300 (N_32300,N_27664,N_29360);
or U32301 (N_32301,N_29065,N_28617);
and U32302 (N_32302,N_27721,N_29297);
or U32303 (N_32303,N_27852,N_28198);
nand U32304 (N_32304,N_29468,N_29898);
and U32305 (N_32305,N_29823,N_28582);
and U32306 (N_32306,N_29815,N_28675);
and U32307 (N_32307,N_28922,N_29045);
xor U32308 (N_32308,N_29075,N_28757);
or U32309 (N_32309,N_28797,N_29325);
nor U32310 (N_32310,N_28372,N_27511);
or U32311 (N_32311,N_28049,N_29529);
nor U32312 (N_32312,N_28029,N_29467);
nor U32313 (N_32313,N_28662,N_27723);
nand U32314 (N_32314,N_27826,N_28320);
xor U32315 (N_32315,N_28325,N_29608);
and U32316 (N_32316,N_29452,N_29034);
or U32317 (N_32317,N_27819,N_27690);
nand U32318 (N_32318,N_28810,N_29690);
nor U32319 (N_32319,N_28070,N_27979);
or U32320 (N_32320,N_28327,N_27687);
nand U32321 (N_32321,N_28491,N_28121);
nor U32322 (N_32322,N_29958,N_29355);
nand U32323 (N_32323,N_29454,N_28426);
and U32324 (N_32324,N_29278,N_28102);
or U32325 (N_32325,N_29962,N_28783);
nand U32326 (N_32326,N_29154,N_29557);
or U32327 (N_32327,N_29610,N_28433);
xor U32328 (N_32328,N_29124,N_29984);
nand U32329 (N_32329,N_27681,N_27784);
nand U32330 (N_32330,N_29478,N_28808);
or U32331 (N_32331,N_29845,N_29140);
nand U32332 (N_32332,N_28362,N_28375);
nand U32333 (N_32333,N_29364,N_29955);
and U32334 (N_32334,N_28108,N_28982);
nand U32335 (N_32335,N_29634,N_29961);
nand U32336 (N_32336,N_28169,N_29707);
or U32337 (N_32337,N_27982,N_28113);
nand U32338 (N_32338,N_29397,N_29916);
or U32339 (N_32339,N_28452,N_29747);
nor U32340 (N_32340,N_29590,N_27512);
and U32341 (N_32341,N_28229,N_27725);
nor U32342 (N_32342,N_28139,N_27876);
or U32343 (N_32343,N_28150,N_28996);
or U32344 (N_32344,N_28087,N_27676);
nand U32345 (N_32345,N_28353,N_28572);
nand U32346 (N_32346,N_28981,N_29992);
or U32347 (N_32347,N_28972,N_27515);
xnor U32348 (N_32348,N_29811,N_29351);
and U32349 (N_32349,N_29669,N_29573);
or U32350 (N_32350,N_28555,N_27806);
and U32351 (N_32351,N_29546,N_29047);
or U32352 (N_32352,N_27856,N_28155);
nand U32353 (N_32353,N_29828,N_29034);
and U32354 (N_32354,N_27742,N_28732);
nor U32355 (N_32355,N_28921,N_29845);
nor U32356 (N_32356,N_29572,N_27934);
and U32357 (N_32357,N_28448,N_27792);
and U32358 (N_32358,N_28271,N_29525);
nand U32359 (N_32359,N_29899,N_29903);
nor U32360 (N_32360,N_28427,N_29109);
or U32361 (N_32361,N_29731,N_28926);
xnor U32362 (N_32362,N_28513,N_28109);
xor U32363 (N_32363,N_29503,N_29012);
and U32364 (N_32364,N_28252,N_27718);
nand U32365 (N_32365,N_28385,N_27944);
or U32366 (N_32366,N_28357,N_28303);
and U32367 (N_32367,N_29717,N_27527);
xnor U32368 (N_32368,N_29150,N_29890);
nand U32369 (N_32369,N_28319,N_28537);
nand U32370 (N_32370,N_28178,N_28729);
nor U32371 (N_32371,N_29414,N_27808);
and U32372 (N_32372,N_29545,N_27676);
nand U32373 (N_32373,N_28335,N_29957);
and U32374 (N_32374,N_28684,N_27660);
xnor U32375 (N_32375,N_29867,N_29312);
and U32376 (N_32376,N_28902,N_29659);
xnor U32377 (N_32377,N_29850,N_28745);
xor U32378 (N_32378,N_29453,N_29976);
nand U32379 (N_32379,N_28110,N_28898);
xor U32380 (N_32380,N_29338,N_27727);
nor U32381 (N_32381,N_29570,N_29070);
and U32382 (N_32382,N_28786,N_28582);
nand U32383 (N_32383,N_28280,N_28174);
or U32384 (N_32384,N_28259,N_28713);
nor U32385 (N_32385,N_28189,N_29130);
or U32386 (N_32386,N_29359,N_28903);
nand U32387 (N_32387,N_28729,N_27767);
or U32388 (N_32388,N_29226,N_29363);
nand U32389 (N_32389,N_29745,N_27899);
nor U32390 (N_32390,N_28193,N_29709);
nand U32391 (N_32391,N_27605,N_29113);
nand U32392 (N_32392,N_27928,N_28010);
nand U32393 (N_32393,N_29762,N_28052);
and U32394 (N_32394,N_29661,N_29152);
and U32395 (N_32395,N_28782,N_28571);
xor U32396 (N_32396,N_28513,N_29895);
nor U32397 (N_32397,N_29508,N_28251);
xor U32398 (N_32398,N_29822,N_29626);
nand U32399 (N_32399,N_28382,N_29722);
nor U32400 (N_32400,N_29219,N_28898);
or U32401 (N_32401,N_29120,N_28542);
or U32402 (N_32402,N_28172,N_27704);
nor U32403 (N_32403,N_28847,N_29179);
and U32404 (N_32404,N_29926,N_29939);
nor U32405 (N_32405,N_28786,N_28134);
or U32406 (N_32406,N_27797,N_29087);
nand U32407 (N_32407,N_29158,N_27958);
or U32408 (N_32408,N_27532,N_28320);
and U32409 (N_32409,N_28833,N_28008);
nand U32410 (N_32410,N_28445,N_27584);
nand U32411 (N_32411,N_28860,N_28230);
xor U32412 (N_32412,N_28897,N_29377);
xor U32413 (N_32413,N_29117,N_28005);
or U32414 (N_32414,N_27815,N_29848);
and U32415 (N_32415,N_29959,N_28528);
and U32416 (N_32416,N_29666,N_29304);
nand U32417 (N_32417,N_27678,N_29932);
nor U32418 (N_32418,N_27817,N_27760);
xor U32419 (N_32419,N_29358,N_28722);
xnor U32420 (N_32420,N_29578,N_27742);
nand U32421 (N_32421,N_28271,N_28290);
nor U32422 (N_32422,N_29628,N_28955);
or U32423 (N_32423,N_27697,N_28483);
or U32424 (N_32424,N_29278,N_28253);
or U32425 (N_32425,N_29302,N_29568);
nand U32426 (N_32426,N_28167,N_29567);
nor U32427 (N_32427,N_28703,N_29580);
nand U32428 (N_32428,N_28961,N_29846);
and U32429 (N_32429,N_29886,N_29843);
nand U32430 (N_32430,N_28375,N_29117);
xor U32431 (N_32431,N_29052,N_29295);
or U32432 (N_32432,N_29564,N_27992);
nand U32433 (N_32433,N_27971,N_29365);
nor U32434 (N_32434,N_28501,N_29607);
xnor U32435 (N_32435,N_28779,N_29452);
nand U32436 (N_32436,N_29660,N_29808);
or U32437 (N_32437,N_27791,N_29952);
nor U32438 (N_32438,N_27894,N_27828);
nand U32439 (N_32439,N_27900,N_28604);
nand U32440 (N_32440,N_28093,N_27628);
nor U32441 (N_32441,N_29319,N_28018);
xnor U32442 (N_32442,N_29455,N_29860);
and U32443 (N_32443,N_29934,N_28678);
nand U32444 (N_32444,N_27741,N_29732);
or U32445 (N_32445,N_29610,N_28926);
xor U32446 (N_32446,N_28924,N_27773);
or U32447 (N_32447,N_27610,N_28384);
or U32448 (N_32448,N_29002,N_29899);
nand U32449 (N_32449,N_28412,N_27800);
xor U32450 (N_32450,N_28024,N_29475);
and U32451 (N_32451,N_28714,N_29972);
nor U32452 (N_32452,N_28913,N_27513);
and U32453 (N_32453,N_29249,N_29892);
xor U32454 (N_32454,N_28498,N_29398);
nand U32455 (N_32455,N_29840,N_27603);
or U32456 (N_32456,N_28139,N_29192);
or U32457 (N_32457,N_28997,N_28023);
and U32458 (N_32458,N_28888,N_27866);
nor U32459 (N_32459,N_28802,N_28900);
and U32460 (N_32460,N_28403,N_28010);
nand U32461 (N_32461,N_29217,N_29252);
nor U32462 (N_32462,N_28212,N_29018);
and U32463 (N_32463,N_29816,N_28880);
and U32464 (N_32464,N_28896,N_29356);
xor U32465 (N_32465,N_27576,N_28031);
nor U32466 (N_32466,N_29495,N_29020);
or U32467 (N_32467,N_29996,N_29659);
or U32468 (N_32468,N_28167,N_28926);
or U32469 (N_32469,N_28947,N_29417);
xnor U32470 (N_32470,N_29326,N_28013);
nand U32471 (N_32471,N_28175,N_28263);
nand U32472 (N_32472,N_29205,N_27778);
nand U32473 (N_32473,N_28760,N_27943);
and U32474 (N_32474,N_28500,N_28957);
and U32475 (N_32475,N_28427,N_29325);
or U32476 (N_32476,N_27958,N_29935);
and U32477 (N_32477,N_28668,N_28161);
and U32478 (N_32478,N_29840,N_29379);
or U32479 (N_32479,N_29511,N_29657);
or U32480 (N_32480,N_28296,N_29739);
nor U32481 (N_32481,N_29745,N_28231);
or U32482 (N_32482,N_27806,N_29986);
xnor U32483 (N_32483,N_29816,N_29901);
or U32484 (N_32484,N_29330,N_27520);
nand U32485 (N_32485,N_29338,N_29482);
xor U32486 (N_32486,N_27733,N_29289);
and U32487 (N_32487,N_28769,N_28868);
nor U32488 (N_32488,N_28462,N_27798);
xor U32489 (N_32489,N_29511,N_29682);
xor U32490 (N_32490,N_27878,N_29288);
nor U32491 (N_32491,N_28679,N_27977);
nor U32492 (N_32492,N_28306,N_29467);
and U32493 (N_32493,N_29663,N_28375);
or U32494 (N_32494,N_29735,N_27791);
xor U32495 (N_32495,N_28305,N_28021);
or U32496 (N_32496,N_28519,N_29142);
or U32497 (N_32497,N_29416,N_27969);
nor U32498 (N_32498,N_29110,N_29205);
and U32499 (N_32499,N_29995,N_28105);
xnor U32500 (N_32500,N_30830,N_31180);
xnor U32501 (N_32501,N_31011,N_31104);
nor U32502 (N_32502,N_30752,N_32397);
nand U32503 (N_32503,N_32053,N_31502);
nand U32504 (N_32504,N_31302,N_31666);
xor U32505 (N_32505,N_31267,N_31137);
nand U32506 (N_32506,N_31798,N_30472);
nor U32507 (N_32507,N_30702,N_32278);
and U32508 (N_32508,N_31009,N_30464);
nor U32509 (N_32509,N_32434,N_30844);
nand U32510 (N_32510,N_30477,N_31187);
or U32511 (N_32511,N_31990,N_30398);
nor U32512 (N_32512,N_31437,N_31958);
nand U32513 (N_32513,N_31877,N_31116);
xnor U32514 (N_32514,N_31290,N_32047);
and U32515 (N_32515,N_31475,N_31670);
nor U32516 (N_32516,N_32445,N_30971);
xor U32517 (N_32517,N_30358,N_30671);
nor U32518 (N_32518,N_31146,N_31166);
or U32519 (N_32519,N_32155,N_30575);
xor U32520 (N_32520,N_30680,N_31381);
xnor U32521 (N_32521,N_31681,N_32080);
nand U32522 (N_32522,N_32476,N_30037);
nand U32523 (N_32523,N_31047,N_31677);
nor U32524 (N_32524,N_31350,N_30587);
nand U32525 (N_32525,N_30317,N_30743);
or U32526 (N_32526,N_30879,N_31592);
or U32527 (N_32527,N_31625,N_30474);
xor U32528 (N_32528,N_31838,N_30019);
nand U32529 (N_32529,N_30406,N_31477);
and U32530 (N_32530,N_32052,N_30824);
nand U32531 (N_32531,N_32045,N_31496);
nand U32532 (N_32532,N_31804,N_32348);
and U32533 (N_32533,N_32470,N_30742);
or U32534 (N_32534,N_32163,N_31227);
nor U32535 (N_32535,N_30336,N_32316);
xor U32536 (N_32536,N_31490,N_30664);
nand U32537 (N_32537,N_31080,N_31360);
xor U32538 (N_32538,N_32036,N_32106);
or U32539 (N_32539,N_31195,N_31012);
and U32540 (N_32540,N_30940,N_30488);
nor U32541 (N_32541,N_30013,N_30583);
nor U32542 (N_32542,N_31777,N_31675);
nor U32543 (N_32543,N_32289,N_30321);
xnor U32544 (N_32544,N_30465,N_30224);
nand U32545 (N_32545,N_31521,N_31067);
and U32546 (N_32546,N_32023,N_31595);
or U32547 (N_32547,N_30952,N_31183);
xor U32548 (N_32548,N_32439,N_30517);
nand U32549 (N_32549,N_31782,N_30399);
xnor U32550 (N_32550,N_31509,N_30443);
or U32551 (N_32551,N_31332,N_30648);
or U32552 (N_32552,N_32478,N_30293);
or U32553 (N_32553,N_30288,N_30056);
xnor U32554 (N_32554,N_31366,N_30350);
or U32555 (N_32555,N_30341,N_31357);
or U32556 (N_32556,N_30910,N_32220);
and U32557 (N_32557,N_30335,N_30894);
and U32558 (N_32558,N_30163,N_31096);
xnor U32559 (N_32559,N_31701,N_30397);
nand U32560 (N_32560,N_30951,N_30802);
and U32561 (N_32561,N_32229,N_30751);
or U32562 (N_32562,N_31388,N_31072);
xor U32563 (N_32563,N_32062,N_30820);
nor U32564 (N_32564,N_30964,N_31452);
xor U32565 (N_32565,N_32097,N_30209);
xor U32566 (N_32566,N_30057,N_30716);
nand U32567 (N_32567,N_31462,N_30106);
nor U32568 (N_32568,N_32083,N_30093);
nand U32569 (N_32569,N_31400,N_32124);
nor U32570 (N_32570,N_30721,N_30495);
nor U32571 (N_32571,N_31486,N_30549);
and U32572 (N_32572,N_32302,N_32255);
xnor U32573 (N_32573,N_32184,N_30214);
or U32574 (N_32574,N_31880,N_30467);
xor U32575 (N_32575,N_32252,N_32328);
nor U32576 (N_32576,N_31539,N_30707);
and U32577 (N_32577,N_31805,N_31766);
xor U32578 (N_32578,N_30065,N_31780);
nor U32579 (N_32579,N_31121,N_31225);
or U32580 (N_32580,N_32017,N_31278);
xor U32581 (N_32581,N_30788,N_31045);
nor U32582 (N_32582,N_30231,N_31476);
xor U32583 (N_32583,N_30923,N_31075);
or U32584 (N_32584,N_30098,N_30731);
and U32585 (N_32585,N_30318,N_30957);
nand U32586 (N_32586,N_30502,N_31313);
or U32587 (N_32587,N_30208,N_30083);
or U32588 (N_32588,N_31402,N_31193);
nand U32589 (N_32589,N_30251,N_32313);
and U32590 (N_32590,N_31663,N_31175);
and U32591 (N_32591,N_31404,N_31752);
and U32592 (N_32592,N_30927,N_30486);
and U32593 (N_32593,N_31079,N_30260);
xnor U32594 (N_32594,N_30221,N_32341);
nor U32595 (N_32595,N_31272,N_31082);
nand U32596 (N_32596,N_30794,N_31478);
and U32597 (N_32597,N_30897,N_30361);
xor U32598 (N_32598,N_32419,N_30058);
nor U32599 (N_32599,N_31176,N_30503);
xor U32600 (N_32600,N_32007,N_32485);
nand U32601 (N_32601,N_30976,N_31337);
xnor U32602 (N_32602,N_30255,N_30049);
nand U32603 (N_32603,N_31600,N_32162);
and U32604 (N_32604,N_30855,N_30681);
nand U32605 (N_32605,N_30124,N_32072);
and U32606 (N_32606,N_31436,N_31140);
nand U32607 (N_32607,N_32076,N_31020);
or U32608 (N_32608,N_32411,N_31441);
or U32609 (N_32609,N_30813,N_30781);
nor U32610 (N_32610,N_31247,N_31453);
nor U32611 (N_32611,N_30603,N_30369);
and U32612 (N_32612,N_31824,N_32379);
or U32613 (N_32613,N_30890,N_30111);
nand U32614 (N_32614,N_31786,N_30330);
or U32615 (N_32615,N_30339,N_31529);
or U32616 (N_32616,N_30627,N_31370);
nor U32617 (N_32617,N_31390,N_30446);
nand U32618 (N_32618,N_32139,N_30798);
nor U32619 (N_32619,N_31073,N_32116);
nor U32620 (N_32620,N_30407,N_32333);
and U32621 (N_32621,N_31908,N_30157);
nor U32622 (N_32622,N_32081,N_31499);
or U32623 (N_32623,N_31724,N_31467);
and U32624 (N_32624,N_31434,N_30693);
nand U32625 (N_32625,N_30195,N_30316);
and U32626 (N_32626,N_31841,N_32268);
nor U32627 (N_32627,N_31565,N_30101);
or U32628 (N_32628,N_30484,N_32132);
nor U32629 (N_32629,N_30179,N_30092);
xnor U32630 (N_32630,N_31374,N_30705);
and U32631 (N_32631,N_30168,N_30104);
and U32632 (N_32632,N_31288,N_30212);
nand U32633 (N_32633,N_31488,N_30711);
and U32634 (N_32634,N_30972,N_31318);
or U32635 (N_32635,N_30701,N_31001);
xor U32636 (N_32636,N_30310,N_32234);
and U32637 (N_32637,N_30079,N_32195);
xnor U32638 (N_32638,N_30823,N_30021);
xnor U32639 (N_32639,N_32054,N_31362);
or U32640 (N_32640,N_30076,N_30827);
nand U32641 (N_32641,N_31937,N_30814);
xor U32642 (N_32642,N_32179,N_31553);
xnor U32643 (N_32643,N_31036,N_30918);
and U32644 (N_32644,N_31888,N_30980);
or U32645 (N_32645,N_32457,N_30557);
xor U32646 (N_32646,N_31796,N_30937);
nand U32647 (N_32647,N_30419,N_32211);
or U32648 (N_32648,N_32405,N_30966);
nor U32649 (N_32649,N_31693,N_31523);
xor U32650 (N_32650,N_30613,N_31783);
and U32651 (N_32651,N_31062,N_30478);
nand U32652 (N_32652,N_31519,N_30757);
xor U32653 (N_32653,N_30803,N_31525);
xnor U32654 (N_32654,N_31627,N_32094);
nor U32655 (N_32655,N_30385,N_31471);
nor U32656 (N_32656,N_31720,N_30508);
nor U32657 (N_32657,N_31760,N_31793);
or U32658 (N_32658,N_32322,N_30044);
nand U32659 (N_32659,N_32198,N_32145);
nand U32660 (N_32660,N_30097,N_30619);
xnor U32661 (N_32661,N_32304,N_30302);
or U32662 (N_32662,N_30417,N_32366);
xor U32663 (N_32663,N_30975,N_30566);
nand U32664 (N_32664,N_31095,N_30708);
nand U32665 (N_32665,N_31754,N_31207);
nand U32666 (N_32666,N_31644,N_30158);
nor U32667 (N_32667,N_30760,N_32260);
or U32668 (N_32668,N_30663,N_30012);
or U32669 (N_32669,N_32086,N_30642);
nand U32670 (N_32670,N_32060,N_30942);
xnor U32671 (N_32671,N_30235,N_31161);
or U32672 (N_32672,N_32059,N_31244);
xor U32673 (N_32673,N_31678,N_31006);
and U32674 (N_32674,N_30256,N_31491);
nand U32675 (N_32675,N_31427,N_32368);
nor U32676 (N_32676,N_31409,N_30732);
or U32677 (N_32677,N_30052,N_31930);
or U32678 (N_32678,N_31098,N_31713);
or U32679 (N_32679,N_30838,N_30299);
and U32680 (N_32680,N_30073,N_30120);
nor U32681 (N_32681,N_30935,N_31301);
nor U32682 (N_32682,N_30074,N_30659);
nand U32683 (N_32683,N_30329,N_32236);
nand U32684 (N_32684,N_31781,N_30762);
and U32685 (N_32685,N_31673,N_32185);
nand U32686 (N_32686,N_30748,N_31065);
xor U32687 (N_32687,N_31587,N_31588);
and U32688 (N_32688,N_31349,N_30261);
and U32689 (N_32689,N_30997,N_32219);
xnor U32690 (N_32690,N_30833,N_30623);
and U32691 (N_32691,N_30876,N_30002);
or U32692 (N_32692,N_30018,N_31929);
nor U32693 (N_32693,N_31931,N_32320);
xnor U32694 (N_32694,N_30230,N_30257);
xor U32695 (N_32695,N_30969,N_32259);
nand U32696 (N_32696,N_30694,N_30600);
and U32697 (N_32697,N_30840,N_32373);
nand U32698 (N_32698,N_31808,N_32100);
and U32699 (N_32699,N_31719,N_30775);
and U32700 (N_32700,N_30143,N_31384);
and U32701 (N_32701,N_32374,N_30034);
xnor U32702 (N_32702,N_31863,N_31992);
nor U32703 (N_32703,N_30679,N_32009);
nand U32704 (N_32704,N_30550,N_30423);
nand U32705 (N_32705,N_31778,N_31199);
nor U32706 (N_32706,N_31163,N_31858);
nand U32707 (N_32707,N_32074,N_31108);
nor U32708 (N_32708,N_31051,N_31895);
and U32709 (N_32709,N_31603,N_30872);
xnor U32710 (N_32710,N_30411,N_31642);
nor U32711 (N_32711,N_30384,N_30948);
and U32712 (N_32712,N_30943,N_30063);
xor U32713 (N_32713,N_31165,N_32228);
xor U32714 (N_32714,N_30574,N_31469);
and U32715 (N_32715,N_30602,N_30095);
xor U32716 (N_32716,N_31764,N_31076);
and U32717 (N_32717,N_30780,N_31691);
xor U32718 (N_32718,N_31910,N_30887);
xor U32719 (N_32719,N_30658,N_30882);
xor U32720 (N_32720,N_30354,N_31159);
and U32721 (N_32721,N_31413,N_31300);
or U32722 (N_32722,N_31394,N_30447);
xnor U32723 (N_32723,N_31218,N_30277);
xnor U32724 (N_32724,N_30886,N_31917);
and U32725 (N_32725,N_31470,N_30936);
xnor U32726 (N_32726,N_31152,N_31083);
and U32727 (N_32727,N_31255,N_30046);
nor U32728 (N_32728,N_30215,N_31368);
or U32729 (N_32729,N_30071,N_31634);
nand U32730 (N_32730,N_30722,N_30278);
or U32731 (N_32731,N_30624,N_30677);
xnor U32732 (N_32732,N_31927,N_30345);
and U32733 (N_32733,N_31396,N_31262);
nor U32734 (N_32734,N_30473,N_31739);
nand U32735 (N_32735,N_32004,N_30959);
nor U32736 (N_32736,N_31329,N_30586);
or U32737 (N_32737,N_31352,N_32262);
nor U32738 (N_32738,N_31348,N_30118);
and U32739 (N_32739,N_32150,N_32077);
or U32740 (N_32740,N_32484,N_31316);
nor U32741 (N_32741,N_31391,N_30510);
or U32742 (N_32742,N_31758,N_30629);
nor U32743 (N_32743,N_31881,N_31148);
and U32744 (N_32744,N_31221,N_31530);
or U32745 (N_32745,N_30558,N_31298);
and U32746 (N_32746,N_31795,N_32144);
nor U32747 (N_32747,N_32256,N_31056);
nor U32748 (N_32748,N_31331,N_32308);
nand U32749 (N_32749,N_31321,N_31621);
and U32750 (N_32750,N_30616,N_31043);
nor U32751 (N_32751,N_30675,N_31944);
xor U32752 (N_32752,N_30818,N_31535);
and U32753 (N_32753,N_30242,N_30933);
xor U32754 (N_32754,N_32026,N_32334);
xor U32755 (N_32755,N_31527,N_32258);
xor U32756 (N_32756,N_30553,N_30008);
and U32757 (N_32757,N_31052,N_30159);
and U32758 (N_32758,N_32424,N_31576);
nor U32759 (N_32759,N_32444,N_31585);
or U32760 (N_32760,N_30281,N_32188);
and U32761 (N_32761,N_31103,N_31905);
xor U32762 (N_32762,N_32156,N_30800);
or U32763 (N_32763,N_31772,N_30432);
xor U32764 (N_32764,N_30615,N_30804);
or U32765 (N_32765,N_31308,N_31878);
xor U32766 (N_32766,N_32046,N_30921);
xor U32767 (N_32767,N_32315,N_31834);
or U32768 (N_32768,N_30469,N_31609);
or U32769 (N_32769,N_30598,N_31936);
xor U32770 (N_32770,N_32107,N_31344);
and U32771 (N_32771,N_31860,N_32013);
nand U32772 (N_32772,N_31984,N_30344);
xor U32773 (N_32773,N_30402,N_31042);
and U32774 (N_32774,N_31179,N_31144);
or U32775 (N_32775,N_30753,N_31698);
and U32776 (N_32776,N_32340,N_31069);
or U32777 (N_32777,N_31981,N_32460);
nor U32778 (N_32778,N_31828,N_30950);
or U32779 (N_32779,N_32474,N_30403);
nor U32780 (N_32780,N_30107,N_30949);
or U32781 (N_32781,N_31971,N_32117);
xnor U32782 (N_32782,N_30254,N_31431);
xor U32783 (N_32783,N_31216,N_31306);
or U32784 (N_32784,N_32396,N_30893);
nand U32785 (N_32785,N_30301,N_30229);
or U32786 (N_32786,N_30489,N_32431);
and U32787 (N_32787,N_31816,N_30584);
nor U32788 (N_32788,N_30730,N_30851);
nand U32789 (N_32789,N_31951,N_31641);
xor U32790 (N_32790,N_30033,N_30173);
and U32791 (N_32791,N_31983,N_30703);
and U32792 (N_32792,N_32199,N_30082);
xor U32793 (N_32793,N_31122,N_30248);
nor U32794 (N_32794,N_31265,N_31729);
and U32795 (N_32795,N_30090,N_31970);
nor U32796 (N_32796,N_30607,N_31188);
nand U32797 (N_32797,N_30915,N_31091);
nor U32798 (N_32798,N_31451,N_31653);
and U32799 (N_32799,N_30456,N_30713);
and U32800 (N_32800,N_30968,N_30868);
nor U32801 (N_32801,N_31946,N_30956);
xor U32802 (N_32802,N_30320,N_31645);
nor U32803 (N_32803,N_31210,N_31147);
nand U32804 (N_32804,N_32449,N_31715);
nand U32805 (N_32805,N_31546,N_31989);
nor U32806 (N_32806,N_32443,N_32427);
and U32807 (N_32807,N_32183,N_31259);
nor U32808 (N_32808,N_32129,N_31597);
or U32809 (N_32809,N_30691,N_30723);
and U32810 (N_32810,N_32490,N_32465);
xnor U32811 (N_32811,N_32486,N_31767);
nand U32812 (N_32812,N_32468,N_31656);
and U32813 (N_32813,N_32064,N_30391);
nand U32814 (N_32814,N_31733,N_30871);
or U32815 (N_32815,N_31143,N_31215);
and U32816 (N_32816,N_31005,N_30852);
or U32817 (N_32817,N_31817,N_31775);
nand U32818 (N_32818,N_30688,N_30548);
and U32819 (N_32819,N_32051,N_30847);
nor U32820 (N_32820,N_31177,N_31369);
xnor U32821 (N_32821,N_31866,N_32420);
nand U32822 (N_32822,N_31571,N_30494);
nand U32823 (N_32823,N_32393,N_32137);
nor U32824 (N_32824,N_31234,N_31128);
and U32825 (N_32825,N_31567,N_30777);
nand U32826 (N_32826,N_31867,N_31030);
and U32827 (N_32827,N_32001,N_30131);
and U32828 (N_32828,N_31872,N_32038);
xnor U32829 (N_32829,N_32164,N_31743);
and U32830 (N_32830,N_31900,N_31061);
nor U32831 (N_32831,N_32141,N_32391);
xor U32832 (N_32832,N_30072,N_31174);
and U32833 (N_32833,N_31070,N_32428);
xnor U32834 (N_32834,N_31765,N_30304);
nor U32835 (N_32835,N_30706,N_31696);
or U32836 (N_32836,N_30005,N_32096);
xor U32837 (N_32837,N_30001,N_30116);
or U32838 (N_32838,N_30130,N_32121);
xnor U32839 (N_32839,N_31706,N_31150);
nor U32840 (N_32840,N_30853,N_32016);
xnor U32841 (N_32841,N_30645,N_31555);
and U32842 (N_32842,N_31317,N_30126);
nand U32843 (N_32843,N_30110,N_30576);
xor U32844 (N_32844,N_31432,N_30259);
or U32845 (N_32845,N_31735,N_30690);
and U32846 (N_32846,N_32135,N_32002);
nand U32847 (N_32847,N_31498,N_30306);
xor U32848 (N_32848,N_30979,N_32147);
nand U32849 (N_32849,N_30776,N_32346);
or U32850 (N_32850,N_31230,N_31168);
nor U32851 (N_32851,N_32497,N_31500);
nand U32852 (N_32852,N_31154,N_31996);
or U32853 (N_32853,N_30865,N_31551);
nor U32854 (N_32854,N_31818,N_32288);
and U32855 (N_32855,N_31566,N_31497);
or U32856 (N_32856,N_32380,N_31223);
xor U32857 (N_32857,N_31721,N_30528);
nor U32858 (N_32858,N_31934,N_31066);
nand U32859 (N_32859,N_30920,N_30866);
nor U32860 (N_32860,N_30389,N_31768);
nand U32861 (N_32861,N_30040,N_30274);
and U32862 (N_32862,N_32435,N_32222);
xnor U32863 (N_32863,N_31307,N_32386);
xor U32864 (N_32864,N_31287,N_31246);
nor U32865 (N_32865,N_31723,N_31945);
nand U32866 (N_32866,N_32394,N_30601);
nand U32867 (N_32867,N_31843,N_30286);
nor U32868 (N_32868,N_31607,N_31049);
nor U32869 (N_32869,N_31660,N_31756);
and U32870 (N_32870,N_32453,N_31113);
nor U32871 (N_32871,N_30699,N_30468);
nor U32872 (N_32872,N_32338,N_30010);
xnor U32873 (N_32873,N_31444,N_30009);
nor U32874 (N_32874,N_30460,N_30377);
xnor U32875 (N_32875,N_30636,N_31842);
nand U32876 (N_32876,N_31209,N_31563);
xor U32877 (N_32877,N_32296,N_31372);
xor U32878 (N_32878,N_31543,N_30889);
nor U32879 (N_32879,N_31871,N_30068);
xnor U32880 (N_32880,N_30653,N_31568);
and U32881 (N_32881,N_31868,N_31710);
xor U32882 (N_32882,N_32012,N_31658);
nor U32883 (N_32883,N_31652,N_32310);
xor U32884 (N_32884,N_31189,N_31319);
nor U32885 (N_32885,N_31186,N_30408);
or U32886 (N_32886,N_32114,N_30400);
and U32887 (N_32887,N_30480,N_30630);
and U32888 (N_32888,N_31697,N_31776);
nand U32889 (N_32889,N_31325,N_30487);
and U32890 (N_32890,N_31510,N_31809);
nor U32891 (N_32891,N_31340,N_32403);
or U32892 (N_32892,N_31248,N_31633);
nand U32893 (N_32893,N_32172,N_31687);
and U32894 (N_32894,N_30036,N_31728);
nand U32895 (N_32895,N_30799,N_30485);
or U32896 (N_32896,N_30139,N_31851);
or U32897 (N_32897,N_32003,N_31613);
and U32898 (N_32898,N_31039,N_30911);
and U32899 (N_32899,N_30471,N_31922);
xnor U32900 (N_32900,N_31662,N_30991);
nor U32901 (N_32901,N_30129,N_30367);
nor U32902 (N_32902,N_30618,N_31483);
nor U32903 (N_32903,N_31800,N_30178);
or U32904 (N_32904,N_30386,N_32058);
nor U32905 (N_32905,N_31229,N_30265);
and U32906 (N_32906,N_30631,N_32105);
nor U32907 (N_32907,N_31727,N_32407);
nor U32908 (N_32908,N_30570,N_32385);
nor U32909 (N_32909,N_30622,N_30401);
nor U32910 (N_32910,N_31802,N_30873);
nor U32911 (N_32911,N_31578,N_32082);
or U32912 (N_32912,N_32138,N_31770);
or U32913 (N_32913,N_31655,N_30342);
nor U32914 (N_32914,N_31356,N_31909);
nor U32915 (N_32915,N_30849,N_31425);
or U32916 (N_32916,N_30481,N_30839);
xnor U32917 (N_32917,N_31460,N_31387);
nor U32918 (N_32918,N_30053,N_31884);
or U32919 (N_32919,N_30081,N_30426);
nand U32920 (N_32920,N_31220,N_30592);
or U32921 (N_32921,N_30112,N_30704);
nand U32922 (N_32922,N_32178,N_31725);
or U32923 (N_32923,N_31968,N_31852);
nand U32924 (N_32924,N_30733,N_32475);
nor U32925 (N_32925,N_30533,N_31395);
and U32926 (N_32926,N_31286,N_31506);
xor U32927 (N_32927,N_31414,N_30507);
or U32928 (N_32928,N_31417,N_30294);
nand U32929 (N_32929,N_30099,N_31938);
xnor U32930 (N_32930,N_32267,N_30205);
xnor U32931 (N_32931,N_31988,N_30782);
nor U32932 (N_32932,N_32111,N_32378);
xor U32933 (N_32933,N_30767,N_31115);
nor U32934 (N_32934,N_31085,N_30669);
nor U32935 (N_32935,N_32237,N_31022);
nor U32936 (N_32936,N_31547,N_30222);
nor U32937 (N_32937,N_31790,N_30220);
and U32938 (N_32938,N_31669,N_31918);
nand U32939 (N_32939,N_30199,N_31980);
nand U32940 (N_32940,N_32277,N_31053);
nand U32941 (N_32941,N_31338,N_30543);
nand U32942 (N_32942,N_31648,N_31593);
nand U32943 (N_32943,N_31015,N_30638);
or U32944 (N_32944,N_31242,N_30709);
nor U32945 (N_32945,N_31038,N_30148);
xor U32946 (N_32946,N_31579,N_30685);
nand U32947 (N_32947,N_31791,N_30884);
xor U32948 (N_32948,N_31398,N_32048);
xnor U32949 (N_32949,N_31716,N_30461);
nor U32950 (N_32950,N_31416,N_31392);
or U32951 (N_32951,N_30944,N_30994);
nand U32952 (N_32952,N_32142,N_30526);
nand U32953 (N_32953,N_30060,N_30102);
xor U32954 (N_32954,N_31774,N_32112);
nand U32955 (N_32955,N_30774,N_30182);
and U32956 (N_32956,N_31826,N_30515);
nor U32957 (N_32957,N_30719,N_30821);
nand U32958 (N_32958,N_30992,N_30521);
nor U32959 (N_32959,N_32270,N_30346);
and U32960 (N_32960,N_30393,N_32173);
nand U32961 (N_32961,N_31750,N_30922);
nor U32962 (N_32962,N_30564,N_30357);
or U32963 (N_32963,N_32362,N_31882);
nor U32964 (N_32964,N_31173,N_31273);
xnor U32965 (N_32965,N_31222,N_32287);
nand U32966 (N_32966,N_31745,N_31311);
xnor U32967 (N_32967,N_31389,N_31487);
xor U32968 (N_32968,N_30878,N_30275);
and U32969 (N_32969,N_30308,N_31380);
and U32970 (N_32970,N_32271,N_32073);
and U32971 (N_32971,N_30903,N_32022);
nand U32972 (N_32972,N_31953,N_32305);
and U32973 (N_32973,N_31589,N_31463);
nand U32974 (N_32974,N_30877,N_31604);
or U32975 (N_32975,N_31952,N_30571);
nor U32976 (N_32976,N_31266,N_31494);
xnor U32977 (N_32977,N_31068,N_30166);
and U32978 (N_32978,N_31700,N_31894);
nand U32979 (N_32979,N_31505,N_31747);
or U32980 (N_32980,N_31197,N_31468);
nand U32981 (N_32981,N_31423,N_30739);
nand U32982 (N_32982,N_30902,N_32454);
xnor U32983 (N_32983,N_30764,N_32212);
and U32984 (N_32984,N_31446,N_30412);
nor U32985 (N_32985,N_31077,N_30689);
or U32986 (N_32986,N_30712,N_31397);
nor U32987 (N_32987,N_31455,N_30449);
and U32988 (N_32988,N_31461,N_31458);
xor U32989 (N_32989,N_31580,N_30476);
nor U32990 (N_32990,N_30007,N_32487);
and U32991 (N_32991,N_31245,N_32110);
nand U32992 (N_32992,N_32087,N_32451);
and U32993 (N_32993,N_31393,N_31586);
nor U32994 (N_32994,N_30267,N_31619);
nor U32995 (N_32995,N_30128,N_30458);
nor U32996 (N_32996,N_31692,N_31861);
xnor U32997 (N_32997,N_30756,N_32175);
nor U32998 (N_32998,N_30559,N_32126);
or U32999 (N_32999,N_32015,N_32230);
nor U33000 (N_33000,N_30309,N_32342);
and U33001 (N_33001,N_31919,N_30191);
nor U33002 (N_33002,N_32495,N_31459);
nand U33003 (N_33003,N_31562,N_31848);
nor U33004 (N_33004,N_31442,N_31797);
xor U33005 (N_33005,N_31276,N_30715);
nor U33006 (N_33006,N_30547,N_31825);
xor U33007 (N_33007,N_31702,N_31985);
and U33008 (N_33008,N_32167,N_30505);
nand U33009 (N_33009,N_30088,N_30810);
and U33010 (N_33010,N_30953,N_32415);
or U33011 (N_33011,N_32447,N_32351);
xor U33012 (N_33012,N_30300,N_31335);
and U33013 (N_33013,N_32430,N_31964);
xnor U33014 (N_33014,N_30684,N_31044);
or U33015 (N_33015,N_31732,N_30904);
nor U33016 (N_33016,N_32246,N_32067);
or U33017 (N_33017,N_30410,N_31829);
or U33018 (N_33018,N_31133,N_32160);
or U33019 (N_33019,N_31637,N_32063);
or U33020 (N_33020,N_31058,N_31041);
nand U33021 (N_33021,N_32225,N_30815);
or U33022 (N_33022,N_31703,N_31602);
nand U33023 (N_33023,N_32187,N_32194);
and U33024 (N_33024,N_30239,N_30499);
nand U33025 (N_33025,N_32233,N_32243);
xnor U33026 (N_33026,N_30899,N_30497);
and U33027 (N_33027,N_30193,N_30243);
or U33028 (N_33028,N_30250,N_31741);
and U33029 (N_33029,N_31837,N_30283);
or U33030 (N_33030,N_30811,N_30812);
and U33031 (N_33031,N_31890,N_30125);
and U33032 (N_33032,N_32196,N_32471);
and U33033 (N_33033,N_30226,N_32425);
and U33034 (N_33034,N_30817,N_30854);
and U33035 (N_33035,N_31684,N_32332);
nor U33036 (N_33036,N_31126,N_31614);
xnor U33037 (N_33037,N_32031,N_31081);
xor U33038 (N_33038,N_30024,N_32149);
and U33039 (N_33039,N_31239,N_31134);
or U33040 (N_33040,N_31528,N_30155);
nand U33041 (N_33041,N_32413,N_31029);
nand U33042 (N_33042,N_32350,N_31202);
and U33043 (N_33043,N_30087,N_30634);
or U33044 (N_33044,N_30789,N_31254);
xor U33045 (N_33045,N_31688,N_30962);
nor U33046 (N_33046,N_32400,N_31192);
nand U33047 (N_33047,N_31640,N_30234);
nor U33048 (N_33048,N_31591,N_30652);
or U33049 (N_33049,N_31856,N_31679);
nor U33050 (N_33050,N_30219,N_30042);
nand U33051 (N_33051,N_31516,N_31862);
nor U33052 (N_33052,N_30981,N_30343);
nand U33053 (N_33053,N_30883,N_30761);
nor U33054 (N_33054,N_30778,N_31690);
and U33055 (N_33055,N_30045,N_30758);
and U33056 (N_33056,N_30032,N_30181);
or U33057 (N_33057,N_32266,N_31667);
or U33058 (N_33058,N_30977,N_30651);
or U33059 (N_33059,N_31811,N_30896);
or U33060 (N_33060,N_30655,N_30773);
and U33061 (N_33061,N_31023,N_30555);
nor U33062 (N_33062,N_30122,N_30483);
nor U33063 (N_33063,N_30405,N_32075);
and U33064 (N_33064,N_30160,N_30916);
nand U33065 (N_33065,N_32301,N_31059);
nand U33066 (N_33066,N_31473,N_32377);
nor U33067 (N_33067,N_31367,N_32197);
nand U33068 (N_33068,N_30608,N_31124);
and U33069 (N_33069,N_31063,N_31084);
xnor U33070 (N_33070,N_30470,N_31003);
or U33071 (N_33071,N_30563,N_32130);
nand U33072 (N_33072,N_30387,N_32232);
and U33073 (N_33073,N_31346,N_31846);
and U33074 (N_33074,N_31608,N_30491);
or U33075 (N_33075,N_30784,N_30945);
nand U33076 (N_33076,N_30569,N_30579);
xor U33077 (N_33077,N_30596,N_31445);
xnor U33078 (N_33078,N_31885,N_30946);
or U33079 (N_33079,N_31206,N_31185);
nor U33080 (N_33080,N_31541,N_32410);
and U33081 (N_33081,N_31999,N_30463);
nand U33082 (N_33082,N_31088,N_30183);
and U33083 (N_33083,N_30963,N_31064);
or U33084 (N_33084,N_31501,N_30436);
nor U33085 (N_33085,N_30825,N_30271);
and U33086 (N_33086,N_31575,N_31522);
and U33087 (N_33087,N_32034,N_31190);
nor U33088 (N_33088,N_31365,N_31671);
nand U33089 (N_33089,N_32307,N_30552);
or U33090 (N_33090,N_30059,N_31016);
nand U33091 (N_33091,N_32244,N_32161);
xnor U33092 (N_33092,N_31991,N_30961);
xnor U33093 (N_33093,N_30835,N_30990);
nand U33094 (N_33094,N_30416,N_30674);
or U33095 (N_33095,N_30791,N_30796);
xor U33096 (N_33096,N_31194,N_31995);
nor U33097 (N_33097,N_31665,N_32104);
xnor U33098 (N_33098,N_32049,N_31712);
or U33099 (N_33099,N_32241,N_30174);
or U33100 (N_33100,N_32037,N_30809);
or U33101 (N_33101,N_31151,N_31426);
or U33102 (N_33102,N_31954,N_31034);
or U33103 (N_33103,N_30745,N_30355);
or U33104 (N_33104,N_30206,N_31736);
nand U33105 (N_33105,N_31260,N_30974);
and U33106 (N_33106,N_30885,N_32203);
and U33107 (N_33107,N_30289,N_31751);
and U33108 (N_33108,N_30617,N_31156);
nor U33109 (N_33109,N_31630,N_32349);
nand U33110 (N_33110,N_32452,N_30770);
nand U33111 (N_33111,N_31605,N_31833);
xor U33112 (N_33112,N_32043,N_32298);
and U33113 (N_33113,N_30171,N_31659);
nand U33114 (N_33114,N_31911,N_31017);
and U33115 (N_33115,N_30086,N_31507);
or U33116 (N_33116,N_30925,N_32193);
and U33117 (N_33117,N_31916,N_30801);
xnor U33118 (N_33118,N_30881,N_32458);
nor U33119 (N_33119,N_31013,N_30030);
and U33120 (N_33120,N_31236,N_31167);
or U33121 (N_33121,N_31717,N_30292);
nand U33122 (N_33122,N_32192,N_30246);
nand U33123 (N_33123,N_30718,N_30614);
nand U33124 (N_33124,N_31010,N_31261);
nor U33125 (N_33125,N_30768,N_31515);
or U33126 (N_33126,N_31611,N_32103);
and U33127 (N_33127,N_31896,N_31942);
nor U33128 (N_33128,N_30187,N_32216);
or U33129 (N_33129,N_30700,N_32108);
nor U33130 (N_33130,N_32249,N_30728);
or U33131 (N_33131,N_31212,N_32214);
xor U33132 (N_33132,N_32325,N_31564);
nor U33133 (N_33133,N_31106,N_31819);
xor U33134 (N_33134,N_30077,N_32098);
nor U33135 (N_33135,N_31726,N_32181);
nand U33136 (N_33136,N_30540,N_31859);
xor U33137 (N_33137,N_32020,N_30572);
nand U33138 (N_33138,N_32323,N_32493);
xnor U33139 (N_33139,N_30459,N_32274);
xnor U33140 (N_33140,N_32027,N_30268);
and U33141 (N_33141,N_31258,N_30932);
or U33142 (N_33142,N_30577,N_31975);
and U33143 (N_33143,N_30437,N_30931);
or U33144 (N_33144,N_30660,N_30434);
nand U33145 (N_33145,N_31415,N_30066);
nand U33146 (N_33146,N_30117,N_30984);
and U33147 (N_33147,N_31364,N_32078);
xor U33148 (N_33148,N_30797,N_32446);
nand U33149 (N_33149,N_30857,N_31599);
or U33150 (N_33150,N_31960,N_31289);
xnor U33151 (N_33151,N_30146,N_31326);
and U33152 (N_33152,N_32438,N_30720);
nand U33153 (N_33153,N_32005,N_30611);
xor U33154 (N_33154,N_30192,N_32019);
nor U33155 (N_33155,N_32303,N_30051);
and U33156 (N_33156,N_30698,N_31788);
nand U33157 (N_33157,N_31709,N_31296);
or U33158 (N_33158,N_31028,N_30518);
nand U33159 (N_33159,N_31762,N_30448);
or U33160 (N_33160,N_31035,N_32285);
or U33161 (N_33161,N_30319,N_30207);
nor U33162 (N_33162,N_31672,N_32044);
or U33163 (N_33163,N_31447,N_30466);
and U33164 (N_33164,N_31171,N_31864);
and U33165 (N_33165,N_30185,N_30114);
and U33166 (N_33166,N_31920,N_32295);
nand U33167 (N_33167,N_31887,N_30779);
or U33168 (N_33168,N_31792,N_31378);
nand U33169 (N_33169,N_32190,N_31966);
and U33170 (N_33170,N_31518,N_30198);
or U33171 (N_33171,N_31722,N_32109);
nand U33172 (N_33172,N_32032,N_30285);
nand U33173 (N_33173,N_31172,N_31214);
nor U33174 (N_33174,N_31440,N_30573);
and U33175 (N_33175,N_31050,N_30697);
nor U33176 (N_33176,N_30356,N_31406);
nor U33177 (N_33177,N_31508,N_30496);
nand U33178 (N_33178,N_32384,N_32498);
and U33179 (N_33179,N_31004,N_31830);
xnor U33180 (N_33180,N_30172,N_31731);
nand U33181 (N_33181,N_31142,N_32056);
xnor U33182 (N_33182,N_31574,N_31162);
and U33183 (N_33183,N_30783,N_30123);
nor U33184 (N_33184,N_32251,N_32140);
or U33185 (N_33185,N_31297,N_30223);
or U33186 (N_33186,N_30149,N_31689);
nand U33187 (N_33187,N_30625,N_32127);
nand U33188 (N_33188,N_31341,N_30368);
nor U33189 (N_33189,N_30338,N_31657);
nand U33190 (N_33190,N_31421,N_30091);
and U33191 (N_33191,N_31794,N_31320);
and U33192 (N_33192,N_30029,N_32223);
and U33193 (N_33193,N_31583,N_32448);
and U33194 (N_33194,N_31554,N_30280);
nor U33195 (N_33195,N_30973,N_31503);
nand U33196 (N_33196,N_31324,N_32010);
xnor U33197 (N_33197,N_31274,N_32422);
nand U33198 (N_33198,N_32180,N_31046);
nor U33199 (N_33199,N_30258,N_30427);
nor U33200 (N_33200,N_30808,N_31661);
nand U33201 (N_33201,N_31734,N_31027);
nor U33202 (N_33202,N_32433,N_31897);
nand U33203 (N_33203,N_31074,N_32025);
or U33204 (N_33204,N_30127,N_30360);
nand U33205 (N_33205,N_32264,N_31465);
and U33206 (N_33206,N_30919,N_32169);
and U33207 (N_33207,N_32240,N_31631);
nor U33208 (N_33208,N_31957,N_31008);
nor U33209 (N_33209,N_30989,N_31870);
nand U33210 (N_33210,N_31814,N_30067);
xnor U33211 (N_33211,N_31969,N_32360);
nand U33212 (N_33212,N_31285,N_32235);
or U33213 (N_33213,N_30177,N_32151);
or U33214 (N_33214,N_30983,N_31226);
or U33215 (N_33215,N_31213,N_32335);
xnor U33216 (N_33216,N_31994,N_32207);
nor U33217 (N_33217,N_31594,N_31883);
nor U33218 (N_33218,N_32029,N_30532);
nand U33219 (N_33219,N_31914,N_30504);
and U33220 (N_33220,N_32174,N_30011);
nor U33221 (N_33221,N_32416,N_30190);
nand U33222 (N_33222,N_31803,N_31196);
or U33223 (N_33223,N_31204,N_31363);
and U33224 (N_33224,N_30431,N_31385);
nor U33225 (N_33225,N_31454,N_30023);
nand U33226 (N_33226,N_32221,N_30754);
xor U33227 (N_33227,N_32464,N_30475);
nor U33228 (N_33228,N_31322,N_30831);
nand U33229 (N_33229,N_30837,N_32412);
or U33230 (N_33230,N_30985,N_30594);
nor U33231 (N_33231,N_31757,N_32356);
and U33232 (N_33232,N_30870,N_30295);
and U33233 (N_33233,N_30151,N_30683);
xnor U33234 (N_33234,N_31827,N_30740);
and U33235 (N_33235,N_31354,N_30589);
nor U33236 (N_33236,N_31823,N_31686);
and U33237 (N_33237,N_31928,N_32292);
xnor U33238 (N_33238,N_30597,N_30864);
and U33239 (N_33239,N_32463,N_30539);
or U33240 (N_33240,N_30218,N_30506);
and U33241 (N_33241,N_31865,N_30892);
or U33242 (N_33242,N_31558,N_32071);
and U33243 (N_33243,N_31129,N_31618);
and U33244 (N_33244,N_31117,N_31466);
and U33245 (N_33245,N_31328,N_30912);
and U33246 (N_33246,N_30006,N_32006);
xnor U33247 (N_33247,N_32189,N_30270);
nor U33248 (N_33248,N_30015,N_31749);
nand U33249 (N_33249,N_32324,N_32050);
nor U33250 (N_33250,N_30136,N_30834);
nor U33251 (N_33251,N_31674,N_32263);
and U33252 (N_33252,N_30856,N_30070);
nor U33253 (N_33253,N_30666,N_30395);
xor U33254 (N_33254,N_32361,N_31753);
nor U33255 (N_33255,N_32272,N_31131);
and U33256 (N_33256,N_30103,N_31787);
or U33257 (N_33257,N_32441,N_31303);
and U33258 (N_33258,N_32409,N_31130);
xor U33259 (N_33259,N_31224,N_31109);
nor U33260 (N_33260,N_30353,N_30202);
xor U33261 (N_33261,N_30245,N_31915);
xor U33262 (N_33262,N_31590,N_31596);
or U33263 (N_33263,N_31853,N_31420);
nor U33264 (N_33264,N_30816,N_31649);
or U33265 (N_33265,N_31511,N_30089);
nor U33266 (N_33266,N_30519,N_30201);
nand U33267 (N_33267,N_32300,N_31107);
and U33268 (N_33268,N_32265,N_32337);
xnor U33269 (N_33269,N_31606,N_31810);
nand U33270 (N_33270,N_31323,N_30939);
and U33271 (N_33271,N_31921,N_31294);
xnor U33272 (N_33272,N_30734,N_30726);
and U33273 (N_33273,N_30374,N_31208);
and U33274 (N_33274,N_30941,N_30806);
and U33275 (N_33275,N_32242,N_32000);
nor U33276 (N_33276,N_30490,N_31577);
or U33277 (N_33277,N_32417,N_30514);
nor U33278 (N_33278,N_31799,N_31164);
xnor U33279 (N_33279,N_32148,N_32085);
nand U33280 (N_33280,N_32294,N_31099);
nand U33281 (N_33281,N_30637,N_31000);
or U33282 (N_33282,N_30084,N_31026);
or U33283 (N_33283,N_32279,N_32101);
or U33284 (N_33284,N_31836,N_31901);
or U33285 (N_33285,N_30137,N_30909);
or U33286 (N_33286,N_31987,N_31869);
and U33287 (N_33287,N_31235,N_30264);
nor U33288 (N_33288,N_30492,N_31993);
xnor U33289 (N_33289,N_30988,N_30326);
nor U33290 (N_33290,N_31333,N_30900);
and U33291 (N_33291,N_32462,N_30438);
or U33292 (N_33292,N_32068,N_31998);
nor U33293 (N_33293,N_32134,N_32432);
nand U33294 (N_33294,N_31959,N_32011);
or U33295 (N_33295,N_30888,N_31548);
nand U33296 (N_33296,N_32345,N_32157);
nand U33297 (N_33297,N_30807,N_31635);
xnor U33298 (N_33298,N_31241,N_32191);
xor U33299 (N_33299,N_31110,N_32170);
nor U33300 (N_33300,N_31623,N_31545);
or U33301 (N_33301,N_30513,N_31977);
or U33302 (N_33302,N_31145,N_31184);
nor U33303 (N_33303,N_30444,N_31250);
nand U33304 (N_33304,N_31304,N_31912);
and U33305 (N_33305,N_30562,N_31399);
and U33306 (N_33306,N_31559,N_31435);
nand U33307 (N_33307,N_30861,N_31240);
nor U33308 (N_33308,N_30591,N_30891);
nor U33309 (N_33309,N_31705,N_30247);
and U33310 (N_33310,N_30523,N_31449);
or U33311 (N_33311,N_30392,N_30150);
xnor U33312 (N_33312,N_31092,N_31903);
or U33313 (N_33313,N_30455,N_31252);
nor U33314 (N_33314,N_32239,N_32482);
or U33315 (N_33315,N_32477,N_30017);
nor U33316 (N_33316,N_30200,N_30331);
or U33317 (N_33317,N_31685,N_30759);
and U33318 (N_33318,N_30305,N_31032);
and U33319 (N_33319,N_32408,N_32177);
xor U33320 (N_33320,N_32488,N_30863);
nor U33321 (N_33321,N_30189,N_30641);
and U33322 (N_33322,N_31448,N_30272);
xor U33323 (N_33323,N_30273,N_31283);
nand U33324 (N_33324,N_32143,N_32079);
nand U33325 (N_33325,N_31293,N_31141);
and U33326 (N_33326,N_30364,N_30428);
nand U33327 (N_33327,N_30588,N_31643);
and U33328 (N_33328,N_31118,N_31514);
and U33329 (N_33329,N_30237,N_31182);
xnor U33330 (N_33330,N_31178,N_30425);
nor U33331 (N_33331,N_30435,N_31200);
nand U33332 (N_33332,N_31493,N_30161);
nor U33333 (N_33333,N_30646,N_31263);
nand U33334 (N_33334,N_30832,N_32200);
nand U33335 (N_33335,N_32339,N_31581);
nand U33336 (N_33336,N_31761,N_31330);
nand U33337 (N_33337,N_31299,N_31615);
nand U33338 (N_33338,N_30901,N_31755);
xor U33339 (N_33339,N_31676,N_30819);
xnor U33340 (N_33340,N_32442,N_30236);
or U33341 (N_33341,N_31935,N_30934);
nor U33342 (N_33342,N_32273,N_32297);
nand U33343 (N_33343,N_32275,N_30987);
nand U33344 (N_33344,N_32227,N_30696);
or U33345 (N_33345,N_31682,N_32231);
or U33346 (N_33346,N_32355,N_30240);
or U33347 (N_33347,N_32014,N_31405);
or U33348 (N_33348,N_31622,N_32414);
or U33349 (N_33349,N_32461,N_30055);
xor U33350 (N_33350,N_30895,N_32091);
nor U33351 (N_33351,N_31845,N_30441);
xnor U33352 (N_33352,N_30498,N_30414);
nor U33353 (N_33353,N_32253,N_30108);
nand U33354 (N_33354,N_31480,N_32311);
or U33355 (N_33355,N_30372,N_30312);
xnor U33356 (N_33356,N_30147,N_30452);
xnor U33357 (N_33357,N_31886,N_30153);
nor U33358 (N_33358,N_30445,N_32306);
xor U33359 (N_33359,N_30105,N_31054);
and U33360 (N_33360,N_31310,N_32154);
and U33361 (N_33361,N_30140,N_32095);
nand U33362 (N_33362,N_30580,N_32248);
nand U33363 (N_33363,N_31123,N_31251);
xnor U33364 (N_33364,N_32450,N_32469);
nor U33365 (N_33365,N_30144,N_32473);
xnor U33366 (N_33366,N_31840,N_30786);
or U33367 (N_33367,N_32357,N_30662);
and U33368 (N_33368,N_31695,N_31158);
or U33369 (N_33369,N_30323,N_32426);
nand U33370 (N_33370,N_30371,N_32314);
xor U33371 (N_33371,N_30249,N_31439);
or U33372 (N_33372,N_31639,N_31489);
nand U33373 (N_33373,N_31629,N_32215);
nand U33374 (N_33374,N_30717,N_31746);
xor U33375 (N_33375,N_31801,N_31377);
nor U33376 (N_33376,N_31874,N_30197);
or U33377 (N_33377,N_31233,N_30829);
and U33378 (N_33378,N_31191,N_30028);
nor U33379 (N_33379,N_32371,N_31281);
xor U33380 (N_33380,N_30735,N_31481);
xor U33381 (N_33381,N_30027,N_32466);
xnor U33382 (N_33382,N_32057,N_31933);
and U33383 (N_33383,N_32389,N_30850);
nand U33384 (N_33384,N_31773,N_32171);
xnor U33385 (N_33385,N_31504,N_30035);
xor U33386 (N_33386,N_30048,N_30233);
or U33387 (N_33387,N_32282,N_30620);
nand U33388 (N_33388,N_32455,N_30695);
nand U33389 (N_33389,N_31334,N_31714);
and U33390 (N_33390,N_31014,N_31383);
nand U33391 (N_33391,N_31114,N_31718);
or U33392 (N_33392,N_31135,N_31443);
and U33393 (N_33393,N_30156,N_30593);
nand U33394 (N_33394,N_32312,N_31021);
xnor U33395 (N_33395,N_32336,N_30599);
nand U33396 (N_33396,N_30661,N_31636);
xor U33397 (N_33397,N_31950,N_30541);
or U33398 (N_33398,N_30993,N_32070);
nor U33399 (N_33399,N_30692,N_31275);
nand U33400 (N_33400,N_30375,N_31264);
or U33401 (N_33401,N_32209,N_30359);
and U33402 (N_33402,N_32329,N_30710);
xor U33403 (N_33403,N_30291,N_30133);
nand U33404 (N_33404,N_32042,N_31704);
and U33405 (N_33405,N_31358,N_31664);
nand U33406 (N_33406,N_30038,N_31632);
nand U33407 (N_33407,N_31359,N_32021);
and U33408 (N_33408,N_30094,N_30378);
nor U33409 (N_33409,N_31102,N_30322);
and U33410 (N_33410,N_30649,N_30628);
or U33411 (N_33411,N_30763,N_31955);
xor U33412 (N_33412,N_32299,N_31057);
or U33413 (N_33413,N_31071,N_30311);
xnor U33414 (N_33414,N_30194,N_31779);
nor U33415 (N_33415,N_30004,N_31336);
and U33416 (N_33416,N_30039,N_32120);
and U33417 (N_33417,N_30500,N_30535);
or U33418 (N_33418,N_30875,N_32061);
nor U33419 (N_33419,N_31291,N_32125);
and U33420 (N_33420,N_30290,N_30433);
or U33421 (N_33421,N_31097,N_31219);
xnor U33422 (N_33422,N_31127,N_31759);
and U33423 (N_33423,N_30388,N_30000);
xor U33424 (N_33424,N_31513,N_32418);
nor U33425 (N_33425,N_32028,N_32284);
nor U33426 (N_33426,N_30747,N_32089);
or U33427 (N_33427,N_30244,N_31292);
or U33428 (N_33428,N_31155,N_31517);
or U33429 (N_33429,N_31484,N_30328);
nand U33430 (N_33430,N_32066,N_30429);
xnor U33431 (N_33431,N_32290,N_30682);
or U33432 (N_33432,N_30665,N_32283);
nand U33433 (N_33433,N_30724,N_30366);
nand U33434 (N_33434,N_30805,N_30217);
nor U33435 (N_33435,N_32358,N_30793);
or U33436 (N_33436,N_31315,N_30737);
nand U33437 (N_33437,N_30567,N_32254);
nor U33438 (N_33438,N_31312,N_31923);
nor U33439 (N_33439,N_31228,N_31351);
or U33440 (N_33440,N_30269,N_30982);
or U33441 (N_33441,N_30204,N_32040);
nand U33442 (N_33442,N_31485,N_31926);
xor U33443 (N_33443,N_30188,N_30612);
or U33444 (N_33444,N_30016,N_32421);
nor U33445 (N_33445,N_31201,N_30228);
xor U33446 (N_33446,N_31738,N_30582);
nor U33447 (N_33447,N_31892,N_31282);
nor U33448 (N_33448,N_30738,N_30568);
nor U33449 (N_33449,N_31019,N_30373);
or U33450 (N_33450,N_31552,N_32365);
or U33451 (N_33451,N_30213,N_31295);
xnor U33452 (N_33452,N_30115,N_31412);
xnor U33453 (N_33453,N_31584,N_32217);
nor U33454 (N_33454,N_30729,N_32280);
nand U33455 (N_33455,N_32165,N_32202);
and U33456 (N_33456,N_32456,N_30746);
xnor U33457 (N_33457,N_30479,N_31533);
nand U33458 (N_33458,N_32372,N_32359);
nor U33459 (N_33459,N_32321,N_31974);
xor U33460 (N_33460,N_31835,N_32370);
nor U33461 (N_33461,N_31430,N_30609);
and U33462 (N_33462,N_31948,N_30003);
nand U33463 (N_33463,N_30282,N_31737);
or U33464 (N_33464,N_31422,N_31132);
and U33465 (N_33465,N_30454,N_31598);
and U33466 (N_33466,N_31450,N_30880);
nor U33467 (N_33467,N_30929,N_31807);
xor U33468 (N_33468,N_31526,N_31238);
nor U33469 (N_33469,N_30913,N_30686);
or U33470 (N_33470,N_31812,N_30164);
nor U33471 (N_33471,N_31474,N_32213);
xor U33472 (N_33472,N_31007,N_31680);
xor U33473 (N_33473,N_31962,N_31269);
and U33474 (N_33474,N_31031,N_30965);
or U33475 (N_33475,N_31268,N_31327);
nand U33476 (N_33476,N_32090,N_32317);
or U33477 (N_33477,N_31339,N_30657);
xnor U33478 (N_33478,N_30678,N_30530);
or U33479 (N_33479,N_31361,N_32492);
nand U33480 (N_33480,N_32102,N_30232);
or U33481 (N_33481,N_30069,N_31820);
nor U33482 (N_33482,N_30442,N_32039);
and U33483 (N_33483,N_32353,N_30512);
nor U33484 (N_33484,N_30749,N_32238);
and U33485 (N_33485,N_30180,N_32245);
and U33486 (N_33486,N_30522,N_31347);
nor U33487 (N_33487,N_30379,N_30238);
and U33488 (N_33488,N_30266,N_31025);
nand U33489 (N_33489,N_32099,N_30050);
or U33490 (N_33490,N_32206,N_30836);
and U33491 (N_33491,N_30654,N_31557);
xnor U33492 (N_33492,N_31973,N_30263);
or U33493 (N_33493,N_30216,N_30842);
and U33494 (N_33494,N_30031,N_31963);
nor U33495 (N_33495,N_30324,N_32479);
or U33496 (N_33496,N_31699,N_30142);
nand U33497 (N_33497,N_32483,N_31342);
and U33498 (N_33498,N_31040,N_31956);
and U33499 (N_33499,N_30307,N_31650);
and U33500 (N_33500,N_31616,N_31309);
or U33501 (N_33501,N_31534,N_31353);
and U33502 (N_33502,N_30370,N_30656);
nand U33503 (N_33503,N_32065,N_30225);
nor U33504 (N_33504,N_31769,N_31105);
nand U33505 (N_33505,N_30766,N_30415);
nor U33506 (N_33506,N_30141,N_32344);
nand U33507 (N_33507,N_30332,N_30365);
and U33508 (N_33508,N_31763,N_30352);
xnor U33509 (N_33509,N_30383,N_30930);
nor U33510 (N_33510,N_30955,N_30175);
and U33511 (N_33511,N_31857,N_32269);
nand U33512 (N_33512,N_30874,N_31708);
nand U33513 (N_33513,N_30348,N_31170);
and U33514 (N_33514,N_31924,N_30297);
nor U33515 (N_33515,N_31037,N_31873);
nor U33516 (N_33516,N_31256,N_32153);
xor U33517 (N_33517,N_30560,N_31237);
nand U33518 (N_33518,N_31433,N_30349);
nor U33519 (N_33519,N_30078,N_32276);
and U33520 (N_33520,N_30062,N_31544);
and U33521 (N_33521,N_31492,N_31119);
xor U33522 (N_33522,N_30362,N_32331);
and U33523 (N_33523,N_30822,N_31139);
xnor U33524 (N_33524,N_30581,N_32387);
nor U33525 (N_33525,N_32363,N_30313);
nand U33526 (N_33526,N_32204,N_31087);
or U33527 (N_33527,N_31855,N_31407);
nand U33528 (N_33528,N_30907,N_31879);
and U33529 (N_33529,N_32402,N_30826);
nand U33530 (N_33530,N_31160,N_31231);
nor U33531 (N_33531,N_31850,N_32088);
xor U33532 (N_33532,N_30453,N_30337);
and U33533 (N_33533,N_31899,N_31002);
xor U33534 (N_33534,N_30075,N_30859);
and U33535 (N_33535,N_31060,N_30621);
xor U33536 (N_33536,N_30999,N_30121);
nor U33537 (N_33537,N_31375,N_31411);
nand U33538 (N_33538,N_31771,N_30924);
or U33539 (N_33539,N_30315,N_31694);
nor U33540 (N_33540,N_31371,N_30914);
xnor U33541 (N_33541,N_30138,N_32024);
or U33542 (N_33542,N_31961,N_30556);
nand U33543 (N_33543,N_31540,N_30154);
nand U33544 (N_33544,N_30413,N_31169);
xor U33545 (N_33545,N_30351,N_30382);
and U33546 (N_33546,N_30995,N_30736);
xnor U33547 (N_33547,N_32146,N_31902);
and U33548 (N_33548,N_30162,N_31628);
nand U33549 (N_33549,N_32388,N_31556);
nor U33550 (N_33550,N_30546,N_31889);
and U33551 (N_33551,N_31401,N_32330);
nand U33552 (N_33552,N_32401,N_30841);
nand U33553 (N_33553,N_30867,N_31089);
or U33554 (N_33554,N_31744,N_31740);
and U33555 (N_33555,N_32496,N_30418);
or U33556 (N_33556,N_30529,N_30908);
or U33557 (N_33557,N_30727,N_31094);
and U33558 (N_33558,N_31986,N_31280);
or U33559 (N_33559,N_31822,N_31806);
and U33560 (N_33560,N_30635,N_30135);
nor U33561 (N_33561,N_32381,N_32030);
or U33562 (N_33562,N_31904,N_30347);
and U33563 (N_33563,N_31582,N_31711);
nand U33564 (N_33564,N_32437,N_30064);
and U33565 (N_33565,N_31048,N_31345);
nor U33566 (N_33566,N_30772,N_32293);
nand U33567 (N_33567,N_30451,N_30769);
nor U33568 (N_33568,N_32367,N_31789);
nand U33569 (N_33569,N_32472,N_31271);
nand U33570 (N_33570,N_31284,N_30626);
xor U33571 (N_33571,N_32158,N_30440);
nand U33572 (N_33572,N_31438,N_32480);
and U33573 (N_33573,N_31646,N_31542);
and U33574 (N_33574,N_32399,N_31549);
and U33575 (N_33575,N_32218,N_31601);
and U33576 (N_33576,N_32033,N_30169);
and U33577 (N_33577,N_31854,N_30422);
nand U33578 (N_33578,N_30869,N_30917);
nand U33579 (N_33579,N_31537,N_31785);
xnor U33580 (N_33580,N_32347,N_31386);
and U33581 (N_33581,N_31181,N_30673);
xnor U33582 (N_33582,N_31839,N_31524);
or U33583 (N_33583,N_31813,N_32382);
and U33584 (N_33584,N_30967,N_31205);
nand U33585 (N_33585,N_30152,N_31913);
and U33586 (N_33586,N_31875,N_30390);
xnor U33587 (N_33587,N_31898,N_30520);
and U33588 (N_33588,N_31495,N_32489);
and U33589 (N_33589,N_31120,N_30928);
nor U33590 (N_33590,N_30595,N_30296);
and U33591 (N_33591,N_30639,N_31101);
xor U33592 (N_33592,N_30545,N_30409);
xor U33593 (N_33593,N_30845,N_32131);
or U33594 (N_33594,N_31090,N_31078);
and U33595 (N_33595,N_31638,N_32440);
nor U33596 (N_33596,N_32247,N_30333);
xor U33597 (N_33597,N_32326,N_31626);
or U33598 (N_33598,N_31844,N_30327);
and U33599 (N_33599,N_30113,N_32008);
and U33600 (N_33600,N_30020,N_30376);
or U33601 (N_33601,N_30846,N_32168);
or U33602 (N_33602,N_30279,N_30672);
or U33603 (N_33603,N_30176,N_32201);
and U33604 (N_33604,N_30186,N_31279);
nor U33605 (N_33605,N_30536,N_30145);
nor U33606 (N_33606,N_30978,N_32398);
and U33607 (N_33607,N_31997,N_31086);
and U33608 (N_33608,N_31949,N_31876);
nor U33609 (N_33609,N_30047,N_32069);
and U33610 (N_33610,N_31932,N_31428);
or U33611 (N_33611,N_30043,N_32352);
nand U33612 (N_33612,N_30022,N_30843);
xor U33613 (N_33613,N_31112,N_30926);
xor U33614 (N_33614,N_30862,N_31482);
nand U33615 (N_33615,N_30668,N_31707);
xor U33616 (N_33616,N_32364,N_30755);
nand U33617 (N_33617,N_30795,N_30252);
nand U33618 (N_33618,N_30096,N_32119);
nor U33619 (N_33619,N_31849,N_30787);
nor U33620 (N_33620,N_30578,N_30714);
xnor U33621 (N_33621,N_32309,N_31249);
and U33622 (N_33622,N_31617,N_30632);
and U33623 (N_33623,N_30054,N_32250);
and U33624 (N_33624,N_30184,N_32406);
and U33625 (N_33625,N_30303,N_32208);
nand U33626 (N_33626,N_32084,N_31536);
or U33627 (N_33627,N_30109,N_31610);
nand U33628 (N_33628,N_32390,N_30421);
nor U33629 (N_33629,N_31217,N_31314);
nand U33630 (N_33630,N_32182,N_31138);
and U33631 (N_33631,N_31343,N_30516);
xor U33632 (N_33632,N_31972,N_30298);
nand U33633 (N_33633,N_31683,N_31538);
nor U33634 (N_33634,N_30848,N_32375);
or U33635 (N_33635,N_32093,N_30424);
nand U33636 (N_33636,N_30640,N_31982);
nor U33637 (N_33637,N_30858,N_30561);
nand U33638 (N_33638,N_30667,N_30606);
and U33639 (N_33639,N_32186,N_31612);
and U33640 (N_33640,N_31243,N_31967);
nand U33641 (N_33641,N_30986,N_30542);
or U33642 (N_33642,N_31742,N_31153);
or U33643 (N_33643,N_31832,N_32055);
nand U33644 (N_33644,N_31253,N_32286);
and U33645 (N_33645,N_32226,N_32159);
and U33646 (N_33646,N_31560,N_30860);
nor U33647 (N_33647,N_31379,N_32499);
xnor U33648 (N_33648,N_31561,N_32376);
xor U33649 (N_33649,N_31429,N_32092);
and U33650 (N_33650,N_31257,N_30544);
or U33651 (N_33651,N_31024,N_30551);
nor U33652 (N_33652,N_30165,N_32383);
nor U33653 (N_33653,N_31668,N_30041);
and U33654 (N_33654,N_31373,N_32115);
nor U33655 (N_33655,N_30590,N_32354);
xor U33656 (N_33656,N_31947,N_31620);
and U33657 (N_33657,N_30394,N_32392);
nor U33658 (N_33658,N_31149,N_31550);
nor U33659 (N_33659,N_30196,N_32018);
and U33660 (N_33660,N_30771,N_30643);
nand U33661 (N_33661,N_31410,N_30334);
and U33662 (N_33662,N_31940,N_32166);
and U33663 (N_33663,N_30167,N_31815);
and U33664 (N_33664,N_32210,N_32395);
nand U33665 (N_33665,N_32319,N_31941);
and U33666 (N_33666,N_31512,N_30905);
nand U33667 (N_33667,N_32152,N_30276);
or U33668 (N_33668,N_32122,N_32494);
xor U33669 (N_33669,N_30898,N_30262);
or U33670 (N_33670,N_31419,N_30605);
xor U33671 (N_33671,N_30524,N_30119);
and U33672 (N_33672,N_31355,N_31100);
and U33673 (N_33673,N_30538,N_31831);
or U33674 (N_33674,N_31570,N_31157);
xor U33675 (N_33675,N_31979,N_31647);
or U33676 (N_33676,N_32113,N_30380);
nor U33677 (N_33677,N_30482,N_30687);
or U33678 (N_33678,N_30958,N_31305);
nand U33679 (N_33679,N_31943,N_30785);
and U33680 (N_33680,N_32429,N_30960);
or U33681 (N_33681,N_31925,N_32491);
and U33682 (N_33682,N_30284,N_31821);
xnor U33683 (N_33683,N_31418,N_30996);
and U33684 (N_33684,N_30287,N_31464);
or U33685 (N_33685,N_32343,N_31624);
and U33686 (N_33686,N_32481,N_30644);
xor U33687 (N_33687,N_31939,N_32423);
nand U33688 (N_33688,N_31730,N_31893);
xor U33689 (N_33689,N_30314,N_31907);
or U33690 (N_33690,N_30610,N_30765);
or U33691 (N_33691,N_30210,N_30650);
xor U33692 (N_33692,N_30501,N_30404);
nand U33693 (N_33693,N_30938,N_30085);
or U33694 (N_33694,N_31532,N_31376);
and U33695 (N_33695,N_30947,N_30906);
and U33696 (N_33696,N_30450,N_31211);
xor U33697 (N_33697,N_30132,N_30462);
xor U33698 (N_33698,N_31965,N_30585);
or U33699 (N_33699,N_31125,N_30744);
or U33700 (N_33700,N_30170,N_32467);
or U33701 (N_33701,N_32224,N_31978);
nor U33702 (N_33702,N_32291,N_30670);
xor U33703 (N_33703,N_31847,N_30203);
xnor U33704 (N_33704,N_31573,N_30790);
or U33705 (N_33705,N_31891,N_31976);
nand U33706 (N_33706,N_30025,N_30565);
nand U33707 (N_33707,N_30750,N_32136);
nor U33708 (N_33708,N_31479,N_32436);
nand U33709 (N_33709,N_30604,N_31520);
nand U33710 (N_33710,N_30493,N_30420);
or U33711 (N_33711,N_32318,N_32261);
and U33712 (N_33712,N_30363,N_30100);
nor U33713 (N_33713,N_30080,N_30970);
xor U33714 (N_33714,N_31382,N_30430);
nand U33715 (N_33715,N_31457,N_31569);
nand U33716 (N_33716,N_30241,N_30537);
nor U33717 (N_33717,N_30014,N_30647);
nand U33718 (N_33718,N_30396,N_30227);
nor U33719 (N_33719,N_30525,N_30457);
nand U33720 (N_33720,N_32035,N_32205);
or U33721 (N_33721,N_32041,N_31424);
and U33722 (N_33722,N_30061,N_30828);
nor U33723 (N_33723,N_32123,N_32257);
or U33724 (N_33724,N_32404,N_30792);
or U33725 (N_33725,N_32118,N_31203);
xor U33726 (N_33726,N_30511,N_32133);
xor U33727 (N_33727,N_31198,N_31572);
or U33728 (N_33728,N_30725,N_31270);
nor U33729 (N_33729,N_31906,N_30509);
and U33730 (N_33730,N_30741,N_32281);
xor U33731 (N_33731,N_30954,N_31531);
nand U33732 (N_33732,N_32128,N_32459);
xor U33733 (N_33733,N_31232,N_31055);
and U33734 (N_33734,N_30998,N_30633);
and U33735 (N_33735,N_32176,N_30527);
nand U33736 (N_33736,N_31408,N_31654);
nor U33737 (N_33737,N_30026,N_30676);
or U33738 (N_33738,N_30325,N_31136);
xnor U33739 (N_33739,N_30253,N_31277);
and U33740 (N_33740,N_31456,N_31403);
nand U33741 (N_33741,N_30340,N_31784);
nor U33742 (N_33742,N_30381,N_31472);
or U33743 (N_33743,N_30531,N_30134);
or U33744 (N_33744,N_32327,N_31111);
and U33745 (N_33745,N_31018,N_31093);
nand U33746 (N_33746,N_30534,N_31033);
nor U33747 (N_33747,N_32369,N_31651);
nand U33748 (N_33748,N_31748,N_30554);
and U33749 (N_33749,N_30211,N_30439);
nand U33750 (N_33750,N_31713,N_32451);
nor U33751 (N_33751,N_31174,N_32447);
or U33752 (N_33752,N_31743,N_30116);
nor U33753 (N_33753,N_30705,N_30343);
xnor U33754 (N_33754,N_32095,N_32186);
and U33755 (N_33755,N_31941,N_30059);
and U33756 (N_33756,N_31896,N_32310);
xor U33757 (N_33757,N_30988,N_31270);
nor U33758 (N_33758,N_30545,N_31764);
or U33759 (N_33759,N_32142,N_31551);
nor U33760 (N_33760,N_31125,N_31548);
xor U33761 (N_33761,N_30686,N_30043);
or U33762 (N_33762,N_31667,N_32430);
nand U33763 (N_33763,N_30488,N_30221);
nand U33764 (N_33764,N_32007,N_30922);
xnor U33765 (N_33765,N_30680,N_31752);
nand U33766 (N_33766,N_30858,N_32285);
or U33767 (N_33767,N_31226,N_30469);
and U33768 (N_33768,N_32198,N_31036);
nor U33769 (N_33769,N_31507,N_31434);
nor U33770 (N_33770,N_30737,N_30405);
nor U33771 (N_33771,N_32034,N_31610);
and U33772 (N_33772,N_30242,N_32283);
xnor U33773 (N_33773,N_31659,N_30754);
nor U33774 (N_33774,N_31666,N_31527);
and U33775 (N_33775,N_31533,N_32033);
and U33776 (N_33776,N_31259,N_31902);
and U33777 (N_33777,N_30767,N_31900);
nand U33778 (N_33778,N_31210,N_31690);
nor U33779 (N_33779,N_31518,N_30340);
nand U33780 (N_33780,N_30554,N_31730);
and U33781 (N_33781,N_31135,N_31769);
nand U33782 (N_33782,N_30040,N_31760);
or U33783 (N_33783,N_30631,N_31505);
or U33784 (N_33784,N_32331,N_31625);
nor U33785 (N_33785,N_32458,N_31577);
nand U33786 (N_33786,N_32384,N_30658);
nor U33787 (N_33787,N_30161,N_30950);
or U33788 (N_33788,N_30734,N_30569);
xnor U33789 (N_33789,N_31632,N_32125);
nand U33790 (N_33790,N_31454,N_31721);
nor U33791 (N_33791,N_31300,N_30280);
nor U33792 (N_33792,N_30952,N_32420);
nor U33793 (N_33793,N_32445,N_30830);
nand U33794 (N_33794,N_31432,N_31348);
and U33795 (N_33795,N_30951,N_30534);
and U33796 (N_33796,N_31588,N_31060);
nand U33797 (N_33797,N_30066,N_30392);
or U33798 (N_33798,N_30561,N_31873);
nor U33799 (N_33799,N_30901,N_32146);
or U33800 (N_33800,N_31515,N_31689);
and U33801 (N_33801,N_30392,N_31192);
xnor U33802 (N_33802,N_30746,N_30681);
nand U33803 (N_33803,N_30579,N_32475);
nor U33804 (N_33804,N_31583,N_31338);
and U33805 (N_33805,N_32227,N_30141);
nor U33806 (N_33806,N_30038,N_30432);
xor U33807 (N_33807,N_30258,N_30881);
and U33808 (N_33808,N_32089,N_30832);
or U33809 (N_33809,N_32369,N_30350);
xnor U33810 (N_33810,N_30058,N_30700);
nor U33811 (N_33811,N_32219,N_31700);
nand U33812 (N_33812,N_32494,N_30061);
and U33813 (N_33813,N_31330,N_30408);
xnor U33814 (N_33814,N_30349,N_30258);
xnor U33815 (N_33815,N_31272,N_30844);
or U33816 (N_33816,N_31229,N_32356);
xor U33817 (N_33817,N_30324,N_32420);
and U33818 (N_33818,N_31911,N_31455);
nand U33819 (N_33819,N_32227,N_30801);
nor U33820 (N_33820,N_30537,N_31681);
xnor U33821 (N_33821,N_31733,N_31147);
nor U33822 (N_33822,N_31329,N_31953);
and U33823 (N_33823,N_32319,N_30994);
nand U33824 (N_33824,N_31225,N_32062);
nor U33825 (N_33825,N_31872,N_31574);
or U33826 (N_33826,N_32181,N_32486);
nor U33827 (N_33827,N_32424,N_30724);
nand U33828 (N_33828,N_31114,N_30815);
nor U33829 (N_33829,N_30024,N_31398);
or U33830 (N_33830,N_32145,N_30255);
nand U33831 (N_33831,N_30525,N_31769);
or U33832 (N_33832,N_32324,N_31119);
xnor U33833 (N_33833,N_30536,N_31189);
nor U33834 (N_33834,N_31122,N_30852);
xnor U33835 (N_33835,N_32168,N_30810);
nand U33836 (N_33836,N_32156,N_32389);
and U33837 (N_33837,N_31065,N_31408);
or U33838 (N_33838,N_32027,N_31819);
and U33839 (N_33839,N_30336,N_30527);
xnor U33840 (N_33840,N_31780,N_30834);
nor U33841 (N_33841,N_31693,N_31155);
nor U33842 (N_33842,N_31188,N_31074);
and U33843 (N_33843,N_30607,N_32050);
nor U33844 (N_33844,N_31989,N_30833);
nor U33845 (N_33845,N_31746,N_32453);
or U33846 (N_33846,N_30520,N_31830);
nand U33847 (N_33847,N_31985,N_32112);
xor U33848 (N_33848,N_32362,N_32401);
nor U33849 (N_33849,N_31912,N_32082);
and U33850 (N_33850,N_31103,N_32326);
nand U33851 (N_33851,N_32418,N_31662);
and U33852 (N_33852,N_30075,N_30966);
or U33853 (N_33853,N_31640,N_31061);
and U33854 (N_33854,N_30050,N_30792);
nor U33855 (N_33855,N_31150,N_31532);
nor U33856 (N_33856,N_30256,N_30083);
nand U33857 (N_33857,N_31337,N_32158);
xnor U33858 (N_33858,N_31790,N_31326);
xnor U33859 (N_33859,N_31282,N_30108);
and U33860 (N_33860,N_30710,N_30866);
or U33861 (N_33861,N_31964,N_31564);
nor U33862 (N_33862,N_31391,N_31507);
nor U33863 (N_33863,N_30307,N_32429);
or U33864 (N_33864,N_31118,N_31699);
and U33865 (N_33865,N_32154,N_30316);
nor U33866 (N_33866,N_31679,N_31106);
or U33867 (N_33867,N_30059,N_30757);
nor U33868 (N_33868,N_32484,N_31453);
nor U33869 (N_33869,N_32168,N_31457);
and U33870 (N_33870,N_30580,N_31188);
nand U33871 (N_33871,N_32020,N_31638);
nand U33872 (N_33872,N_30189,N_30852);
nand U33873 (N_33873,N_30953,N_30347);
xnor U33874 (N_33874,N_31297,N_31992);
nand U33875 (N_33875,N_30573,N_30434);
xnor U33876 (N_33876,N_31567,N_31130);
and U33877 (N_33877,N_30689,N_30060);
or U33878 (N_33878,N_31116,N_32451);
xnor U33879 (N_33879,N_30080,N_31930);
nand U33880 (N_33880,N_31887,N_30478);
or U33881 (N_33881,N_31918,N_30801);
nand U33882 (N_33882,N_31529,N_30125);
xnor U33883 (N_33883,N_30549,N_32154);
and U33884 (N_33884,N_30573,N_31369);
nor U33885 (N_33885,N_32341,N_30278);
or U33886 (N_33886,N_32363,N_31108);
nor U33887 (N_33887,N_30019,N_31638);
xor U33888 (N_33888,N_31811,N_31699);
nand U33889 (N_33889,N_30919,N_30602);
and U33890 (N_33890,N_32278,N_31786);
nor U33891 (N_33891,N_30074,N_30071);
or U33892 (N_33892,N_30033,N_32010);
nor U33893 (N_33893,N_30130,N_31000);
nand U33894 (N_33894,N_31606,N_31969);
nor U33895 (N_33895,N_31617,N_32339);
nand U33896 (N_33896,N_31252,N_31177);
nor U33897 (N_33897,N_31140,N_32263);
nand U33898 (N_33898,N_32166,N_31161);
nor U33899 (N_33899,N_30201,N_32422);
nand U33900 (N_33900,N_30500,N_31090);
and U33901 (N_33901,N_32256,N_31059);
and U33902 (N_33902,N_30076,N_31862);
xor U33903 (N_33903,N_30871,N_30997);
and U33904 (N_33904,N_30113,N_31895);
or U33905 (N_33905,N_31617,N_31235);
nor U33906 (N_33906,N_32377,N_30925);
nor U33907 (N_33907,N_31335,N_31155);
nand U33908 (N_33908,N_31907,N_31813);
xor U33909 (N_33909,N_31946,N_31575);
nand U33910 (N_33910,N_31819,N_31565);
or U33911 (N_33911,N_30795,N_30090);
or U33912 (N_33912,N_30139,N_30853);
nor U33913 (N_33913,N_32305,N_31808);
nor U33914 (N_33914,N_30986,N_31996);
nand U33915 (N_33915,N_31737,N_30738);
xor U33916 (N_33916,N_32050,N_30063);
nor U33917 (N_33917,N_31980,N_32231);
nand U33918 (N_33918,N_31782,N_31552);
nor U33919 (N_33919,N_32068,N_30863);
or U33920 (N_33920,N_30501,N_31459);
nand U33921 (N_33921,N_32040,N_31016);
or U33922 (N_33922,N_31564,N_31905);
and U33923 (N_33923,N_31350,N_32321);
nand U33924 (N_33924,N_31775,N_30023);
xnor U33925 (N_33925,N_31870,N_31878);
nand U33926 (N_33926,N_31991,N_30103);
nand U33927 (N_33927,N_30981,N_30772);
or U33928 (N_33928,N_30001,N_31077);
nand U33929 (N_33929,N_30496,N_30895);
and U33930 (N_33930,N_32101,N_32355);
nand U33931 (N_33931,N_31627,N_30696);
and U33932 (N_33932,N_30809,N_31016);
or U33933 (N_33933,N_31222,N_31120);
or U33934 (N_33934,N_30589,N_32034);
xnor U33935 (N_33935,N_31355,N_30782);
or U33936 (N_33936,N_30738,N_31608);
nor U33937 (N_33937,N_31768,N_32317);
and U33938 (N_33938,N_30402,N_31246);
or U33939 (N_33939,N_30994,N_32287);
nor U33940 (N_33940,N_30989,N_31440);
and U33941 (N_33941,N_30240,N_31492);
nand U33942 (N_33942,N_31184,N_31177);
nor U33943 (N_33943,N_31339,N_32111);
or U33944 (N_33944,N_30660,N_32181);
xor U33945 (N_33945,N_32115,N_32142);
nor U33946 (N_33946,N_31348,N_31010);
and U33947 (N_33947,N_30545,N_30174);
nor U33948 (N_33948,N_31845,N_31368);
and U33949 (N_33949,N_32357,N_32014);
xor U33950 (N_33950,N_32105,N_30527);
or U33951 (N_33951,N_31530,N_31687);
xnor U33952 (N_33952,N_31965,N_30392);
nand U33953 (N_33953,N_30007,N_31582);
nand U33954 (N_33954,N_30134,N_30859);
nand U33955 (N_33955,N_32383,N_30619);
or U33956 (N_33956,N_30385,N_30783);
nand U33957 (N_33957,N_31446,N_31973);
xnor U33958 (N_33958,N_31152,N_32077);
nand U33959 (N_33959,N_30976,N_32292);
xor U33960 (N_33960,N_30823,N_32391);
and U33961 (N_33961,N_31594,N_31804);
xor U33962 (N_33962,N_30533,N_30540);
xor U33963 (N_33963,N_31096,N_31750);
and U33964 (N_33964,N_30382,N_30891);
and U33965 (N_33965,N_31682,N_31373);
nand U33966 (N_33966,N_32124,N_32463);
and U33967 (N_33967,N_31471,N_30053);
nand U33968 (N_33968,N_30501,N_31481);
and U33969 (N_33969,N_30498,N_30222);
nor U33970 (N_33970,N_31562,N_30824);
nand U33971 (N_33971,N_30467,N_30180);
nand U33972 (N_33972,N_30925,N_31634);
nor U33973 (N_33973,N_30540,N_32419);
xnor U33974 (N_33974,N_31295,N_30849);
nand U33975 (N_33975,N_31232,N_30079);
or U33976 (N_33976,N_30890,N_31998);
nor U33977 (N_33977,N_30515,N_30658);
or U33978 (N_33978,N_31475,N_31807);
xor U33979 (N_33979,N_30645,N_30658);
or U33980 (N_33980,N_30186,N_31535);
nand U33981 (N_33981,N_31090,N_31834);
xnor U33982 (N_33982,N_31692,N_31583);
xnor U33983 (N_33983,N_31783,N_32237);
nor U33984 (N_33984,N_30319,N_30992);
nor U33985 (N_33985,N_31937,N_30188);
nand U33986 (N_33986,N_30714,N_32309);
nor U33987 (N_33987,N_31538,N_30032);
nand U33988 (N_33988,N_30767,N_31668);
or U33989 (N_33989,N_30795,N_31487);
xnor U33990 (N_33990,N_31723,N_31589);
or U33991 (N_33991,N_31678,N_31460);
nand U33992 (N_33992,N_30867,N_31871);
xor U33993 (N_33993,N_31591,N_30534);
xnor U33994 (N_33994,N_30867,N_31553);
xor U33995 (N_33995,N_32480,N_30805);
xor U33996 (N_33996,N_30035,N_32272);
nand U33997 (N_33997,N_30596,N_30843);
nor U33998 (N_33998,N_31107,N_31530);
and U33999 (N_33999,N_30721,N_31018);
nand U34000 (N_34000,N_32498,N_30994);
nand U34001 (N_34001,N_31514,N_31141);
and U34002 (N_34002,N_31750,N_30908);
xnor U34003 (N_34003,N_31605,N_31520);
xor U34004 (N_34004,N_32101,N_31108);
xor U34005 (N_34005,N_31012,N_31055);
xor U34006 (N_34006,N_31258,N_30868);
and U34007 (N_34007,N_30826,N_30462);
and U34008 (N_34008,N_32212,N_30776);
nor U34009 (N_34009,N_30397,N_32030);
xor U34010 (N_34010,N_30534,N_31823);
xnor U34011 (N_34011,N_31151,N_31543);
nand U34012 (N_34012,N_30268,N_30244);
nor U34013 (N_34013,N_31245,N_30545);
or U34014 (N_34014,N_30070,N_30864);
nand U34015 (N_34015,N_30837,N_31373);
nor U34016 (N_34016,N_31760,N_30804);
or U34017 (N_34017,N_30763,N_30095);
or U34018 (N_34018,N_30315,N_31321);
nand U34019 (N_34019,N_31516,N_31213);
or U34020 (N_34020,N_30983,N_32210);
nand U34021 (N_34021,N_31249,N_30416);
xor U34022 (N_34022,N_32100,N_31594);
or U34023 (N_34023,N_31430,N_32143);
nor U34024 (N_34024,N_31917,N_31102);
nor U34025 (N_34025,N_31856,N_32268);
nor U34026 (N_34026,N_30175,N_30915);
xnor U34027 (N_34027,N_30457,N_32170);
nand U34028 (N_34028,N_31859,N_32234);
nor U34029 (N_34029,N_31442,N_30314);
and U34030 (N_34030,N_30553,N_30911);
or U34031 (N_34031,N_30065,N_31964);
nor U34032 (N_34032,N_30460,N_30814);
nor U34033 (N_34033,N_31099,N_30742);
nand U34034 (N_34034,N_30000,N_30284);
nand U34035 (N_34035,N_31133,N_31717);
nand U34036 (N_34036,N_30562,N_31385);
or U34037 (N_34037,N_30683,N_32463);
nand U34038 (N_34038,N_32465,N_30446);
nand U34039 (N_34039,N_30389,N_31747);
xor U34040 (N_34040,N_31425,N_32195);
nand U34041 (N_34041,N_30925,N_31639);
and U34042 (N_34042,N_31065,N_31386);
nand U34043 (N_34043,N_30862,N_30534);
xor U34044 (N_34044,N_31963,N_30755);
nand U34045 (N_34045,N_32028,N_30824);
and U34046 (N_34046,N_30226,N_32348);
nor U34047 (N_34047,N_30903,N_31488);
and U34048 (N_34048,N_31786,N_31887);
and U34049 (N_34049,N_31530,N_31864);
nand U34050 (N_34050,N_31585,N_31721);
and U34051 (N_34051,N_30803,N_32000);
nand U34052 (N_34052,N_30543,N_31176);
nor U34053 (N_34053,N_30191,N_30188);
nor U34054 (N_34054,N_31572,N_31064);
xnor U34055 (N_34055,N_30044,N_30901);
or U34056 (N_34056,N_30867,N_30840);
xnor U34057 (N_34057,N_31514,N_31559);
xor U34058 (N_34058,N_31270,N_32406);
nor U34059 (N_34059,N_31830,N_30589);
and U34060 (N_34060,N_32058,N_30517);
and U34061 (N_34061,N_32114,N_31772);
nor U34062 (N_34062,N_32200,N_32232);
xnor U34063 (N_34063,N_32485,N_30351);
or U34064 (N_34064,N_30146,N_30365);
or U34065 (N_34065,N_31359,N_31426);
xnor U34066 (N_34066,N_31927,N_30706);
nand U34067 (N_34067,N_32065,N_31799);
xor U34068 (N_34068,N_31552,N_32493);
nand U34069 (N_34069,N_31732,N_32413);
xor U34070 (N_34070,N_30344,N_30466);
or U34071 (N_34071,N_30032,N_31320);
and U34072 (N_34072,N_30138,N_30617);
xor U34073 (N_34073,N_32385,N_31584);
nor U34074 (N_34074,N_30859,N_31044);
nor U34075 (N_34075,N_32294,N_30751);
and U34076 (N_34076,N_30683,N_30311);
and U34077 (N_34077,N_30104,N_30323);
nor U34078 (N_34078,N_30453,N_30949);
xor U34079 (N_34079,N_30509,N_31440);
xor U34080 (N_34080,N_31473,N_30728);
and U34081 (N_34081,N_31004,N_32433);
xor U34082 (N_34082,N_32194,N_31817);
nor U34083 (N_34083,N_30117,N_30752);
nor U34084 (N_34084,N_30567,N_30438);
nand U34085 (N_34085,N_31688,N_30376);
xor U34086 (N_34086,N_31836,N_31079);
xor U34087 (N_34087,N_30898,N_31895);
and U34088 (N_34088,N_30936,N_31998);
xnor U34089 (N_34089,N_30583,N_31999);
and U34090 (N_34090,N_31332,N_31268);
and U34091 (N_34091,N_32181,N_31831);
nor U34092 (N_34092,N_30060,N_32426);
or U34093 (N_34093,N_32434,N_30088);
nand U34094 (N_34094,N_32371,N_32357);
nand U34095 (N_34095,N_32393,N_31688);
and U34096 (N_34096,N_32369,N_30621);
or U34097 (N_34097,N_31388,N_32458);
nand U34098 (N_34098,N_31221,N_32171);
xnor U34099 (N_34099,N_30894,N_32045);
nor U34100 (N_34100,N_30201,N_30268);
or U34101 (N_34101,N_31402,N_31097);
nand U34102 (N_34102,N_30988,N_30635);
and U34103 (N_34103,N_32498,N_31435);
and U34104 (N_34104,N_30009,N_30538);
nand U34105 (N_34105,N_30184,N_31824);
xnor U34106 (N_34106,N_32159,N_30482);
nand U34107 (N_34107,N_30777,N_30823);
nor U34108 (N_34108,N_30727,N_30664);
and U34109 (N_34109,N_30798,N_30514);
and U34110 (N_34110,N_30652,N_32011);
xnor U34111 (N_34111,N_31220,N_31869);
nand U34112 (N_34112,N_32207,N_30892);
nand U34113 (N_34113,N_31296,N_32403);
xor U34114 (N_34114,N_31042,N_32341);
nand U34115 (N_34115,N_30088,N_30491);
or U34116 (N_34116,N_32498,N_31019);
or U34117 (N_34117,N_32129,N_32324);
and U34118 (N_34118,N_31214,N_30575);
and U34119 (N_34119,N_31524,N_30472);
nand U34120 (N_34120,N_30363,N_32408);
and U34121 (N_34121,N_31439,N_30317);
nand U34122 (N_34122,N_32435,N_30447);
nor U34123 (N_34123,N_31490,N_30469);
and U34124 (N_34124,N_30407,N_32474);
xor U34125 (N_34125,N_30280,N_30396);
nor U34126 (N_34126,N_32209,N_31376);
and U34127 (N_34127,N_30149,N_32266);
or U34128 (N_34128,N_30576,N_32134);
nor U34129 (N_34129,N_31571,N_31820);
nor U34130 (N_34130,N_30765,N_32389);
nor U34131 (N_34131,N_31687,N_30530);
and U34132 (N_34132,N_30699,N_30897);
or U34133 (N_34133,N_30656,N_31846);
or U34134 (N_34134,N_30759,N_32379);
nand U34135 (N_34135,N_31787,N_31257);
nor U34136 (N_34136,N_31483,N_31448);
or U34137 (N_34137,N_32250,N_31120);
and U34138 (N_34138,N_31569,N_30186);
nand U34139 (N_34139,N_30863,N_31232);
nor U34140 (N_34140,N_31219,N_32498);
xor U34141 (N_34141,N_31433,N_31017);
and U34142 (N_34142,N_31935,N_31524);
nor U34143 (N_34143,N_31446,N_30663);
or U34144 (N_34144,N_30002,N_31456);
and U34145 (N_34145,N_30844,N_32201);
or U34146 (N_34146,N_31459,N_31187);
xor U34147 (N_34147,N_30082,N_30965);
or U34148 (N_34148,N_32076,N_31130);
nor U34149 (N_34149,N_30079,N_30378);
nand U34150 (N_34150,N_31076,N_31276);
or U34151 (N_34151,N_32284,N_31998);
xor U34152 (N_34152,N_31022,N_30113);
or U34153 (N_34153,N_32005,N_32444);
nor U34154 (N_34154,N_30061,N_30264);
nor U34155 (N_34155,N_32067,N_31545);
xnor U34156 (N_34156,N_32404,N_30883);
nor U34157 (N_34157,N_32341,N_30881);
nor U34158 (N_34158,N_31894,N_30082);
nand U34159 (N_34159,N_31441,N_30092);
nor U34160 (N_34160,N_32031,N_30237);
xnor U34161 (N_34161,N_31888,N_30990);
or U34162 (N_34162,N_32065,N_30774);
nand U34163 (N_34163,N_32231,N_32352);
xor U34164 (N_34164,N_31957,N_31066);
nand U34165 (N_34165,N_31457,N_30488);
nand U34166 (N_34166,N_30899,N_30091);
xnor U34167 (N_34167,N_32387,N_30625);
nor U34168 (N_34168,N_31792,N_31506);
xor U34169 (N_34169,N_32277,N_31459);
and U34170 (N_34170,N_32293,N_31046);
or U34171 (N_34171,N_32098,N_30310);
nor U34172 (N_34172,N_32141,N_31374);
and U34173 (N_34173,N_30404,N_30650);
and U34174 (N_34174,N_31074,N_31464);
xor U34175 (N_34175,N_31880,N_31432);
nand U34176 (N_34176,N_30042,N_32215);
nor U34177 (N_34177,N_31508,N_30853);
nand U34178 (N_34178,N_30558,N_31993);
or U34179 (N_34179,N_31262,N_30720);
nand U34180 (N_34180,N_30914,N_31610);
nand U34181 (N_34181,N_32493,N_32211);
and U34182 (N_34182,N_31532,N_31643);
nand U34183 (N_34183,N_31701,N_31083);
nor U34184 (N_34184,N_30963,N_30600);
nand U34185 (N_34185,N_31491,N_31432);
nor U34186 (N_34186,N_30862,N_30154);
and U34187 (N_34187,N_31258,N_32278);
nand U34188 (N_34188,N_32242,N_30601);
xor U34189 (N_34189,N_30513,N_32220);
xnor U34190 (N_34190,N_30788,N_30001);
nand U34191 (N_34191,N_32478,N_32441);
nor U34192 (N_34192,N_32017,N_30959);
xnor U34193 (N_34193,N_31294,N_30547);
nor U34194 (N_34194,N_31152,N_30390);
or U34195 (N_34195,N_30850,N_32203);
xnor U34196 (N_34196,N_31024,N_31619);
nor U34197 (N_34197,N_30446,N_30234);
xnor U34198 (N_34198,N_30191,N_31683);
or U34199 (N_34199,N_31663,N_31237);
xnor U34200 (N_34200,N_32063,N_30581);
or U34201 (N_34201,N_32073,N_32423);
nand U34202 (N_34202,N_31019,N_31551);
or U34203 (N_34203,N_31181,N_31917);
nand U34204 (N_34204,N_30828,N_32172);
and U34205 (N_34205,N_30497,N_31887);
or U34206 (N_34206,N_31680,N_32088);
or U34207 (N_34207,N_31877,N_30558);
nand U34208 (N_34208,N_31917,N_30139);
nand U34209 (N_34209,N_30331,N_30929);
or U34210 (N_34210,N_32243,N_31116);
nand U34211 (N_34211,N_30602,N_30064);
nand U34212 (N_34212,N_31384,N_31288);
nand U34213 (N_34213,N_30824,N_31289);
nand U34214 (N_34214,N_32180,N_32016);
and U34215 (N_34215,N_31752,N_30871);
nor U34216 (N_34216,N_32272,N_31821);
or U34217 (N_34217,N_32454,N_32040);
or U34218 (N_34218,N_30959,N_32403);
nor U34219 (N_34219,N_30357,N_32061);
or U34220 (N_34220,N_30115,N_31006);
and U34221 (N_34221,N_31009,N_32340);
nand U34222 (N_34222,N_30764,N_31863);
xnor U34223 (N_34223,N_32036,N_31710);
nor U34224 (N_34224,N_32258,N_30137);
xnor U34225 (N_34225,N_32225,N_31529);
or U34226 (N_34226,N_31893,N_32391);
or U34227 (N_34227,N_31790,N_30238);
nor U34228 (N_34228,N_31914,N_30297);
nand U34229 (N_34229,N_30161,N_30021);
xor U34230 (N_34230,N_31406,N_31498);
nand U34231 (N_34231,N_30220,N_30779);
xnor U34232 (N_34232,N_31921,N_30287);
xor U34233 (N_34233,N_31024,N_32381);
nand U34234 (N_34234,N_32190,N_30736);
nor U34235 (N_34235,N_32192,N_30828);
and U34236 (N_34236,N_31943,N_32424);
and U34237 (N_34237,N_30150,N_30619);
xnor U34238 (N_34238,N_30354,N_31997);
and U34239 (N_34239,N_30124,N_30859);
or U34240 (N_34240,N_31236,N_31762);
or U34241 (N_34241,N_30735,N_30740);
xnor U34242 (N_34242,N_30221,N_30305);
or U34243 (N_34243,N_31737,N_31937);
nand U34244 (N_34244,N_31426,N_32009);
nor U34245 (N_34245,N_32187,N_30467);
nand U34246 (N_34246,N_30716,N_30301);
nand U34247 (N_34247,N_32028,N_32191);
and U34248 (N_34248,N_31678,N_32139);
nand U34249 (N_34249,N_30251,N_31888);
nand U34250 (N_34250,N_32240,N_31484);
nand U34251 (N_34251,N_31418,N_30563);
nor U34252 (N_34252,N_30531,N_31618);
nor U34253 (N_34253,N_30246,N_32266);
or U34254 (N_34254,N_32382,N_31995);
nor U34255 (N_34255,N_31540,N_30450);
and U34256 (N_34256,N_31049,N_30786);
or U34257 (N_34257,N_30167,N_31292);
xnor U34258 (N_34258,N_32355,N_31443);
or U34259 (N_34259,N_30632,N_31364);
or U34260 (N_34260,N_31274,N_30096);
and U34261 (N_34261,N_31174,N_30077);
and U34262 (N_34262,N_30246,N_31335);
or U34263 (N_34263,N_31131,N_30100);
nand U34264 (N_34264,N_31913,N_30328);
or U34265 (N_34265,N_31507,N_32060);
and U34266 (N_34266,N_31805,N_31681);
and U34267 (N_34267,N_31257,N_31392);
xor U34268 (N_34268,N_30034,N_30949);
nor U34269 (N_34269,N_30588,N_30107);
xor U34270 (N_34270,N_32196,N_32164);
nor U34271 (N_34271,N_30011,N_32267);
nand U34272 (N_34272,N_31880,N_32299);
and U34273 (N_34273,N_30802,N_31026);
and U34274 (N_34274,N_32461,N_32315);
and U34275 (N_34275,N_30915,N_30978);
nand U34276 (N_34276,N_31707,N_31976);
nand U34277 (N_34277,N_30602,N_31626);
or U34278 (N_34278,N_30697,N_31474);
xnor U34279 (N_34279,N_31648,N_32047);
nand U34280 (N_34280,N_32070,N_30375);
nor U34281 (N_34281,N_32205,N_32447);
nor U34282 (N_34282,N_32005,N_30144);
or U34283 (N_34283,N_30287,N_30800);
nand U34284 (N_34284,N_32465,N_32321);
nor U34285 (N_34285,N_30946,N_30461);
xor U34286 (N_34286,N_31595,N_30408);
nor U34287 (N_34287,N_32294,N_32482);
xor U34288 (N_34288,N_31484,N_31744);
nor U34289 (N_34289,N_31011,N_32360);
nand U34290 (N_34290,N_30508,N_32122);
xor U34291 (N_34291,N_32460,N_31429);
nand U34292 (N_34292,N_31478,N_30918);
nor U34293 (N_34293,N_30999,N_30250);
xnor U34294 (N_34294,N_30253,N_30655);
and U34295 (N_34295,N_31111,N_31387);
nor U34296 (N_34296,N_32352,N_31814);
xor U34297 (N_34297,N_30460,N_32288);
xor U34298 (N_34298,N_30211,N_32432);
or U34299 (N_34299,N_31769,N_31167);
nand U34300 (N_34300,N_30703,N_32147);
nand U34301 (N_34301,N_32416,N_30059);
nor U34302 (N_34302,N_30990,N_30108);
nand U34303 (N_34303,N_31168,N_31891);
xnor U34304 (N_34304,N_32298,N_31156);
xnor U34305 (N_34305,N_31523,N_31450);
nand U34306 (N_34306,N_32120,N_30217);
nor U34307 (N_34307,N_32193,N_30786);
nand U34308 (N_34308,N_30892,N_32144);
nor U34309 (N_34309,N_31804,N_31171);
or U34310 (N_34310,N_31530,N_32151);
and U34311 (N_34311,N_30373,N_32200);
and U34312 (N_34312,N_31954,N_30117);
and U34313 (N_34313,N_31631,N_32193);
or U34314 (N_34314,N_30838,N_31543);
and U34315 (N_34315,N_30461,N_30491);
xor U34316 (N_34316,N_32125,N_31081);
nand U34317 (N_34317,N_31650,N_31391);
nand U34318 (N_34318,N_31864,N_30086);
nand U34319 (N_34319,N_30099,N_30049);
xnor U34320 (N_34320,N_30452,N_31615);
xnor U34321 (N_34321,N_32489,N_31620);
nor U34322 (N_34322,N_31438,N_32095);
or U34323 (N_34323,N_31883,N_30555);
and U34324 (N_34324,N_30452,N_30704);
and U34325 (N_34325,N_32433,N_32466);
nand U34326 (N_34326,N_31302,N_30883);
nor U34327 (N_34327,N_32288,N_31618);
or U34328 (N_34328,N_31082,N_31930);
and U34329 (N_34329,N_31085,N_30092);
xnor U34330 (N_34330,N_30867,N_31762);
xor U34331 (N_34331,N_30838,N_31080);
xor U34332 (N_34332,N_32307,N_30862);
nand U34333 (N_34333,N_32357,N_31556);
xnor U34334 (N_34334,N_31561,N_32124);
or U34335 (N_34335,N_31962,N_31393);
or U34336 (N_34336,N_31350,N_30031);
and U34337 (N_34337,N_31342,N_31009);
xor U34338 (N_34338,N_32354,N_30317);
nand U34339 (N_34339,N_30824,N_30526);
or U34340 (N_34340,N_32062,N_30789);
nand U34341 (N_34341,N_31183,N_31336);
and U34342 (N_34342,N_30152,N_31737);
and U34343 (N_34343,N_31674,N_32067);
xnor U34344 (N_34344,N_32213,N_30525);
or U34345 (N_34345,N_32184,N_32414);
nand U34346 (N_34346,N_31842,N_30098);
nor U34347 (N_34347,N_30020,N_31146);
nor U34348 (N_34348,N_30302,N_31813);
nand U34349 (N_34349,N_30541,N_31755);
nand U34350 (N_34350,N_31781,N_30794);
xor U34351 (N_34351,N_30518,N_31719);
nand U34352 (N_34352,N_31661,N_30193);
xor U34353 (N_34353,N_30162,N_31978);
or U34354 (N_34354,N_31324,N_30790);
nor U34355 (N_34355,N_30653,N_31664);
or U34356 (N_34356,N_30881,N_30328);
nand U34357 (N_34357,N_30879,N_30331);
nor U34358 (N_34358,N_31250,N_32435);
xnor U34359 (N_34359,N_30754,N_30102);
and U34360 (N_34360,N_30142,N_31250);
xor U34361 (N_34361,N_32375,N_32097);
xnor U34362 (N_34362,N_31143,N_31520);
and U34363 (N_34363,N_30008,N_31269);
nand U34364 (N_34364,N_31743,N_31081);
and U34365 (N_34365,N_30370,N_30069);
and U34366 (N_34366,N_30024,N_30779);
nor U34367 (N_34367,N_30096,N_31968);
or U34368 (N_34368,N_30109,N_31264);
or U34369 (N_34369,N_32122,N_31237);
xor U34370 (N_34370,N_31262,N_30469);
nand U34371 (N_34371,N_30116,N_30976);
and U34372 (N_34372,N_30997,N_31966);
xnor U34373 (N_34373,N_30343,N_32035);
xor U34374 (N_34374,N_31525,N_30169);
or U34375 (N_34375,N_32102,N_31711);
and U34376 (N_34376,N_30061,N_31444);
or U34377 (N_34377,N_31265,N_31392);
xor U34378 (N_34378,N_31500,N_31478);
xor U34379 (N_34379,N_31825,N_32205);
or U34380 (N_34380,N_31741,N_31553);
and U34381 (N_34381,N_30968,N_30561);
or U34382 (N_34382,N_31908,N_30826);
nand U34383 (N_34383,N_30326,N_30194);
and U34384 (N_34384,N_32174,N_32288);
xor U34385 (N_34385,N_30701,N_30158);
xnor U34386 (N_34386,N_30263,N_30433);
and U34387 (N_34387,N_30549,N_32067);
and U34388 (N_34388,N_30232,N_30179);
nand U34389 (N_34389,N_32456,N_31774);
nand U34390 (N_34390,N_31220,N_30262);
xnor U34391 (N_34391,N_30372,N_32390);
nand U34392 (N_34392,N_30730,N_32164);
nand U34393 (N_34393,N_31366,N_31862);
and U34394 (N_34394,N_30356,N_30305);
nor U34395 (N_34395,N_30302,N_31641);
xnor U34396 (N_34396,N_31657,N_31501);
nand U34397 (N_34397,N_31940,N_31166);
nor U34398 (N_34398,N_31397,N_31196);
nand U34399 (N_34399,N_31585,N_30677);
nand U34400 (N_34400,N_32042,N_31355);
or U34401 (N_34401,N_32194,N_30686);
nor U34402 (N_34402,N_30862,N_32197);
xor U34403 (N_34403,N_30366,N_31426);
nand U34404 (N_34404,N_31693,N_30634);
nor U34405 (N_34405,N_30760,N_31155);
xor U34406 (N_34406,N_30727,N_31179);
or U34407 (N_34407,N_30738,N_32323);
xor U34408 (N_34408,N_31932,N_30080);
and U34409 (N_34409,N_31838,N_31771);
nand U34410 (N_34410,N_31005,N_30019);
nor U34411 (N_34411,N_31903,N_30793);
nor U34412 (N_34412,N_31060,N_32044);
nor U34413 (N_34413,N_30720,N_30492);
or U34414 (N_34414,N_30026,N_31067);
and U34415 (N_34415,N_31080,N_31182);
nand U34416 (N_34416,N_31056,N_30279);
nor U34417 (N_34417,N_31918,N_32481);
nand U34418 (N_34418,N_32017,N_30050);
nor U34419 (N_34419,N_32418,N_30778);
or U34420 (N_34420,N_31796,N_30335);
nand U34421 (N_34421,N_31621,N_31123);
xnor U34422 (N_34422,N_30760,N_31377);
xor U34423 (N_34423,N_30157,N_31740);
xor U34424 (N_34424,N_30916,N_31428);
and U34425 (N_34425,N_32264,N_32024);
xor U34426 (N_34426,N_30199,N_31062);
nor U34427 (N_34427,N_31511,N_30977);
nor U34428 (N_34428,N_32054,N_30012);
and U34429 (N_34429,N_31180,N_32193);
or U34430 (N_34430,N_30879,N_31748);
xnor U34431 (N_34431,N_31546,N_32382);
and U34432 (N_34432,N_30238,N_31246);
and U34433 (N_34433,N_32043,N_30902);
xor U34434 (N_34434,N_31536,N_30086);
and U34435 (N_34435,N_31555,N_32177);
nor U34436 (N_34436,N_30018,N_31424);
xor U34437 (N_34437,N_31611,N_32047);
nand U34438 (N_34438,N_31606,N_31950);
and U34439 (N_34439,N_30340,N_31469);
and U34440 (N_34440,N_31151,N_30288);
or U34441 (N_34441,N_30744,N_30096);
or U34442 (N_34442,N_31603,N_30307);
and U34443 (N_34443,N_30261,N_30152);
xnor U34444 (N_34444,N_31154,N_31618);
nand U34445 (N_34445,N_32291,N_31582);
nor U34446 (N_34446,N_32349,N_31165);
nand U34447 (N_34447,N_30931,N_32271);
nand U34448 (N_34448,N_31469,N_30857);
nand U34449 (N_34449,N_32307,N_32112);
nand U34450 (N_34450,N_31151,N_30871);
nand U34451 (N_34451,N_32412,N_32205);
and U34452 (N_34452,N_32413,N_32159);
nor U34453 (N_34453,N_30406,N_31942);
nor U34454 (N_34454,N_30930,N_31603);
xor U34455 (N_34455,N_30828,N_31152);
nor U34456 (N_34456,N_30178,N_31293);
or U34457 (N_34457,N_30392,N_31441);
or U34458 (N_34458,N_30018,N_30488);
nand U34459 (N_34459,N_31015,N_30363);
nor U34460 (N_34460,N_31811,N_31351);
and U34461 (N_34461,N_30303,N_32137);
xnor U34462 (N_34462,N_31439,N_32384);
nor U34463 (N_34463,N_32353,N_30375);
xnor U34464 (N_34464,N_32430,N_30701);
xnor U34465 (N_34465,N_31046,N_31009);
and U34466 (N_34466,N_30990,N_30127);
xor U34467 (N_34467,N_31255,N_32076);
nor U34468 (N_34468,N_30191,N_30542);
and U34469 (N_34469,N_30169,N_30355);
or U34470 (N_34470,N_32492,N_30707);
nand U34471 (N_34471,N_31925,N_30081);
and U34472 (N_34472,N_32323,N_30244);
nand U34473 (N_34473,N_31870,N_31348);
or U34474 (N_34474,N_31669,N_32024);
and U34475 (N_34475,N_32479,N_31955);
and U34476 (N_34476,N_31832,N_30555);
or U34477 (N_34477,N_31407,N_32398);
or U34478 (N_34478,N_32237,N_31430);
or U34479 (N_34479,N_31617,N_31074);
nand U34480 (N_34480,N_31214,N_31535);
nor U34481 (N_34481,N_31012,N_32215);
nand U34482 (N_34482,N_32117,N_31471);
or U34483 (N_34483,N_31619,N_30484);
or U34484 (N_34484,N_30187,N_32034);
xor U34485 (N_34485,N_32414,N_31192);
or U34486 (N_34486,N_32214,N_30486);
and U34487 (N_34487,N_30575,N_30435);
or U34488 (N_34488,N_31868,N_31225);
xnor U34489 (N_34489,N_31165,N_30774);
or U34490 (N_34490,N_32415,N_32490);
and U34491 (N_34491,N_31661,N_31632);
nor U34492 (N_34492,N_32177,N_31557);
nor U34493 (N_34493,N_30584,N_30099);
or U34494 (N_34494,N_31407,N_30508);
nor U34495 (N_34495,N_30896,N_30487);
and U34496 (N_34496,N_32186,N_31085);
nor U34497 (N_34497,N_30542,N_30930);
nand U34498 (N_34498,N_32307,N_31624);
or U34499 (N_34499,N_31588,N_31367);
xor U34500 (N_34500,N_30557,N_31660);
or U34501 (N_34501,N_30847,N_31072);
xor U34502 (N_34502,N_32089,N_32180);
nor U34503 (N_34503,N_30555,N_30035);
nand U34504 (N_34504,N_31499,N_30382);
nand U34505 (N_34505,N_32127,N_31827);
and U34506 (N_34506,N_31506,N_30775);
or U34507 (N_34507,N_30934,N_30905);
xor U34508 (N_34508,N_32459,N_30004);
nand U34509 (N_34509,N_30061,N_32408);
nor U34510 (N_34510,N_30284,N_32231);
and U34511 (N_34511,N_30917,N_30187);
nor U34512 (N_34512,N_31147,N_31051);
nor U34513 (N_34513,N_31172,N_31695);
xnor U34514 (N_34514,N_32191,N_32473);
and U34515 (N_34515,N_31419,N_32376);
nand U34516 (N_34516,N_31656,N_32025);
or U34517 (N_34517,N_32266,N_32436);
nand U34518 (N_34518,N_31913,N_32095);
and U34519 (N_34519,N_32375,N_31837);
and U34520 (N_34520,N_31105,N_32073);
xnor U34521 (N_34521,N_30019,N_31384);
and U34522 (N_34522,N_31694,N_30565);
xnor U34523 (N_34523,N_31225,N_31794);
and U34524 (N_34524,N_30578,N_30833);
or U34525 (N_34525,N_31789,N_30870);
and U34526 (N_34526,N_30077,N_30344);
nor U34527 (N_34527,N_32242,N_30421);
nand U34528 (N_34528,N_30339,N_32122);
nand U34529 (N_34529,N_32472,N_32351);
nand U34530 (N_34530,N_31152,N_31714);
or U34531 (N_34531,N_30356,N_31476);
or U34532 (N_34532,N_31924,N_31219);
or U34533 (N_34533,N_30174,N_32362);
nand U34534 (N_34534,N_32258,N_31528);
nand U34535 (N_34535,N_30277,N_30128);
or U34536 (N_34536,N_31426,N_31382);
or U34537 (N_34537,N_31097,N_30879);
nand U34538 (N_34538,N_31034,N_30195);
nand U34539 (N_34539,N_31910,N_32351);
xor U34540 (N_34540,N_30776,N_31625);
and U34541 (N_34541,N_31256,N_31603);
or U34542 (N_34542,N_32178,N_32356);
and U34543 (N_34543,N_32273,N_30885);
and U34544 (N_34544,N_30136,N_30950);
nand U34545 (N_34545,N_31264,N_30000);
xor U34546 (N_34546,N_31819,N_30063);
or U34547 (N_34547,N_31355,N_30917);
nor U34548 (N_34548,N_31987,N_31785);
and U34549 (N_34549,N_31918,N_31752);
nor U34550 (N_34550,N_30958,N_31860);
and U34551 (N_34551,N_30130,N_31447);
nand U34552 (N_34552,N_31254,N_31571);
and U34553 (N_34553,N_30470,N_30551);
and U34554 (N_34554,N_31614,N_31763);
and U34555 (N_34555,N_30173,N_30784);
and U34556 (N_34556,N_32134,N_31995);
nand U34557 (N_34557,N_30725,N_32326);
nand U34558 (N_34558,N_31125,N_30588);
nor U34559 (N_34559,N_30070,N_32406);
nor U34560 (N_34560,N_30571,N_32421);
nand U34561 (N_34561,N_31389,N_31828);
nand U34562 (N_34562,N_32122,N_31827);
nor U34563 (N_34563,N_30186,N_30157);
and U34564 (N_34564,N_30206,N_32012);
nand U34565 (N_34565,N_31851,N_31232);
nand U34566 (N_34566,N_31019,N_30506);
nand U34567 (N_34567,N_32476,N_30968);
or U34568 (N_34568,N_31068,N_32331);
or U34569 (N_34569,N_32454,N_31670);
and U34570 (N_34570,N_31574,N_30162);
nor U34571 (N_34571,N_30545,N_30042);
or U34572 (N_34572,N_31319,N_30842);
xnor U34573 (N_34573,N_30299,N_30820);
xnor U34574 (N_34574,N_30507,N_32333);
nand U34575 (N_34575,N_31323,N_30144);
nor U34576 (N_34576,N_31501,N_32071);
nor U34577 (N_34577,N_30134,N_30439);
and U34578 (N_34578,N_31701,N_30834);
nand U34579 (N_34579,N_32001,N_30597);
or U34580 (N_34580,N_32078,N_30204);
nor U34581 (N_34581,N_32177,N_32393);
nor U34582 (N_34582,N_31296,N_31644);
nor U34583 (N_34583,N_31151,N_32383);
and U34584 (N_34584,N_32120,N_30931);
nor U34585 (N_34585,N_31338,N_31368);
xnor U34586 (N_34586,N_31033,N_32173);
or U34587 (N_34587,N_32011,N_31128);
and U34588 (N_34588,N_30010,N_31311);
or U34589 (N_34589,N_32045,N_31029);
and U34590 (N_34590,N_30621,N_31396);
nor U34591 (N_34591,N_31036,N_30821);
and U34592 (N_34592,N_32211,N_30490);
nand U34593 (N_34593,N_31122,N_31306);
or U34594 (N_34594,N_30321,N_30700);
nand U34595 (N_34595,N_32145,N_31018);
nor U34596 (N_34596,N_30944,N_30135);
nor U34597 (N_34597,N_30620,N_31122);
or U34598 (N_34598,N_31742,N_30894);
nand U34599 (N_34599,N_31613,N_30813);
or U34600 (N_34600,N_32194,N_30122);
and U34601 (N_34601,N_31249,N_31271);
nand U34602 (N_34602,N_31329,N_32041);
nor U34603 (N_34603,N_30975,N_30322);
nor U34604 (N_34604,N_31254,N_31910);
or U34605 (N_34605,N_32475,N_32183);
nor U34606 (N_34606,N_31640,N_32495);
and U34607 (N_34607,N_32238,N_32278);
or U34608 (N_34608,N_30872,N_31127);
or U34609 (N_34609,N_31899,N_32392);
nand U34610 (N_34610,N_30850,N_31608);
xnor U34611 (N_34611,N_31351,N_30935);
and U34612 (N_34612,N_31853,N_30566);
nor U34613 (N_34613,N_32042,N_30889);
or U34614 (N_34614,N_32428,N_30707);
xor U34615 (N_34615,N_31203,N_30519);
or U34616 (N_34616,N_30795,N_30985);
xnor U34617 (N_34617,N_30985,N_31411);
and U34618 (N_34618,N_30553,N_30022);
and U34619 (N_34619,N_31039,N_31296);
nand U34620 (N_34620,N_31195,N_31482);
xnor U34621 (N_34621,N_31185,N_31970);
nor U34622 (N_34622,N_32277,N_31724);
nand U34623 (N_34623,N_30610,N_32437);
and U34624 (N_34624,N_31609,N_30891);
nand U34625 (N_34625,N_32483,N_32109);
and U34626 (N_34626,N_31365,N_32329);
nor U34627 (N_34627,N_30213,N_30092);
and U34628 (N_34628,N_31313,N_31703);
nor U34629 (N_34629,N_30845,N_32313);
and U34630 (N_34630,N_30413,N_30923);
nor U34631 (N_34631,N_30694,N_30835);
or U34632 (N_34632,N_30759,N_31772);
and U34633 (N_34633,N_31706,N_30338);
xor U34634 (N_34634,N_32081,N_32471);
and U34635 (N_34635,N_30908,N_32334);
xnor U34636 (N_34636,N_31392,N_31005);
or U34637 (N_34637,N_32197,N_31646);
and U34638 (N_34638,N_32409,N_31129);
and U34639 (N_34639,N_32156,N_31606);
or U34640 (N_34640,N_31713,N_31642);
and U34641 (N_34641,N_31375,N_30578);
nor U34642 (N_34642,N_31590,N_32280);
or U34643 (N_34643,N_31092,N_32417);
or U34644 (N_34644,N_30962,N_30396);
and U34645 (N_34645,N_31470,N_32305);
nand U34646 (N_34646,N_30574,N_32332);
nand U34647 (N_34647,N_32296,N_30030);
and U34648 (N_34648,N_32372,N_30292);
or U34649 (N_34649,N_30496,N_30758);
nand U34650 (N_34650,N_31990,N_30387);
nor U34651 (N_34651,N_31618,N_30176);
and U34652 (N_34652,N_31062,N_30703);
xor U34653 (N_34653,N_31729,N_30804);
nor U34654 (N_34654,N_31921,N_30679);
or U34655 (N_34655,N_31162,N_30727);
or U34656 (N_34656,N_30772,N_31467);
nor U34657 (N_34657,N_31605,N_30180);
and U34658 (N_34658,N_30021,N_30893);
nand U34659 (N_34659,N_31866,N_30114);
or U34660 (N_34660,N_31749,N_31884);
nand U34661 (N_34661,N_31249,N_32070);
and U34662 (N_34662,N_31540,N_31396);
and U34663 (N_34663,N_31624,N_32061);
xor U34664 (N_34664,N_30708,N_30176);
nor U34665 (N_34665,N_30515,N_31804);
nand U34666 (N_34666,N_30070,N_32085);
nand U34667 (N_34667,N_30695,N_32134);
and U34668 (N_34668,N_32397,N_30760);
nor U34669 (N_34669,N_30097,N_31439);
or U34670 (N_34670,N_31313,N_30187);
nor U34671 (N_34671,N_30609,N_30734);
xnor U34672 (N_34672,N_31128,N_32117);
or U34673 (N_34673,N_30753,N_32116);
and U34674 (N_34674,N_30557,N_30143);
nand U34675 (N_34675,N_30660,N_30990);
nand U34676 (N_34676,N_30724,N_31610);
or U34677 (N_34677,N_31288,N_30390);
and U34678 (N_34678,N_30768,N_31994);
or U34679 (N_34679,N_30341,N_30422);
or U34680 (N_34680,N_30534,N_30690);
or U34681 (N_34681,N_32349,N_31053);
nand U34682 (N_34682,N_31152,N_30933);
and U34683 (N_34683,N_31879,N_32123);
nand U34684 (N_34684,N_32013,N_31816);
nand U34685 (N_34685,N_30320,N_31902);
or U34686 (N_34686,N_31873,N_30540);
nor U34687 (N_34687,N_31529,N_31457);
xor U34688 (N_34688,N_30845,N_32345);
and U34689 (N_34689,N_31718,N_31994);
and U34690 (N_34690,N_31183,N_31995);
nor U34691 (N_34691,N_30576,N_31896);
nor U34692 (N_34692,N_30251,N_30921);
nor U34693 (N_34693,N_30507,N_30823);
xnor U34694 (N_34694,N_31613,N_32006);
nand U34695 (N_34695,N_31283,N_31731);
nand U34696 (N_34696,N_32350,N_32052);
and U34697 (N_34697,N_31798,N_30706);
or U34698 (N_34698,N_30874,N_32208);
nand U34699 (N_34699,N_31960,N_32284);
nor U34700 (N_34700,N_30436,N_30801);
nor U34701 (N_34701,N_30297,N_30841);
xnor U34702 (N_34702,N_31810,N_32063);
or U34703 (N_34703,N_31671,N_31229);
or U34704 (N_34704,N_32036,N_32293);
or U34705 (N_34705,N_31079,N_32476);
or U34706 (N_34706,N_31456,N_30867);
and U34707 (N_34707,N_30116,N_30423);
or U34708 (N_34708,N_31883,N_30394);
or U34709 (N_34709,N_30654,N_30300);
and U34710 (N_34710,N_30037,N_30656);
nor U34711 (N_34711,N_32159,N_31728);
nand U34712 (N_34712,N_30787,N_31375);
xnor U34713 (N_34713,N_31516,N_31452);
xnor U34714 (N_34714,N_31618,N_32015);
nor U34715 (N_34715,N_31627,N_32486);
xnor U34716 (N_34716,N_30558,N_32158);
or U34717 (N_34717,N_30161,N_32333);
and U34718 (N_34718,N_31814,N_31617);
xor U34719 (N_34719,N_32076,N_31808);
xor U34720 (N_34720,N_30175,N_32097);
nand U34721 (N_34721,N_30336,N_32392);
xnor U34722 (N_34722,N_30431,N_32284);
nand U34723 (N_34723,N_30389,N_32110);
nand U34724 (N_34724,N_31959,N_30406);
nand U34725 (N_34725,N_32155,N_32020);
xor U34726 (N_34726,N_31289,N_32169);
and U34727 (N_34727,N_32049,N_31191);
nand U34728 (N_34728,N_31236,N_30442);
xnor U34729 (N_34729,N_32307,N_30291);
and U34730 (N_34730,N_30889,N_31680);
and U34731 (N_34731,N_30719,N_30857);
and U34732 (N_34732,N_30718,N_32201);
or U34733 (N_34733,N_31632,N_30702);
or U34734 (N_34734,N_32048,N_32162);
or U34735 (N_34735,N_31644,N_30075);
nand U34736 (N_34736,N_30076,N_30342);
or U34737 (N_34737,N_30676,N_30181);
or U34738 (N_34738,N_30847,N_31580);
nand U34739 (N_34739,N_30976,N_30451);
or U34740 (N_34740,N_30248,N_31613);
and U34741 (N_34741,N_30098,N_30343);
nand U34742 (N_34742,N_31591,N_32358);
nor U34743 (N_34743,N_30841,N_30356);
xor U34744 (N_34744,N_31915,N_31628);
and U34745 (N_34745,N_31951,N_32045);
nor U34746 (N_34746,N_32032,N_31466);
nand U34747 (N_34747,N_30138,N_31659);
and U34748 (N_34748,N_32067,N_31919);
xnor U34749 (N_34749,N_31787,N_30158);
nand U34750 (N_34750,N_30569,N_30022);
and U34751 (N_34751,N_31859,N_30255);
or U34752 (N_34752,N_32091,N_31056);
nor U34753 (N_34753,N_30921,N_31700);
xnor U34754 (N_34754,N_31684,N_31048);
or U34755 (N_34755,N_31315,N_31035);
or U34756 (N_34756,N_30920,N_30060);
and U34757 (N_34757,N_31482,N_30340);
xor U34758 (N_34758,N_32301,N_30525);
or U34759 (N_34759,N_32450,N_31019);
nor U34760 (N_34760,N_31902,N_31403);
and U34761 (N_34761,N_31139,N_31839);
nor U34762 (N_34762,N_32475,N_32053);
xor U34763 (N_34763,N_31083,N_31122);
nor U34764 (N_34764,N_32302,N_31659);
or U34765 (N_34765,N_32484,N_31106);
and U34766 (N_34766,N_31665,N_31722);
nand U34767 (N_34767,N_32245,N_30848);
nand U34768 (N_34768,N_30303,N_31781);
nor U34769 (N_34769,N_31894,N_31385);
xor U34770 (N_34770,N_31444,N_32426);
nand U34771 (N_34771,N_31346,N_32342);
and U34772 (N_34772,N_31222,N_31105);
xnor U34773 (N_34773,N_30688,N_30753);
or U34774 (N_34774,N_31389,N_31211);
nor U34775 (N_34775,N_30004,N_30686);
or U34776 (N_34776,N_31086,N_31696);
or U34777 (N_34777,N_30960,N_30166);
nor U34778 (N_34778,N_30540,N_32444);
nand U34779 (N_34779,N_30150,N_31597);
xor U34780 (N_34780,N_31201,N_30140);
xor U34781 (N_34781,N_30781,N_31123);
and U34782 (N_34782,N_32141,N_30091);
nand U34783 (N_34783,N_30605,N_30980);
or U34784 (N_34784,N_31050,N_31380);
nand U34785 (N_34785,N_30802,N_32229);
or U34786 (N_34786,N_30700,N_31924);
or U34787 (N_34787,N_32421,N_30732);
or U34788 (N_34788,N_32296,N_31006);
nand U34789 (N_34789,N_31151,N_30182);
nor U34790 (N_34790,N_31550,N_30411);
nor U34791 (N_34791,N_32262,N_30227);
xnor U34792 (N_34792,N_31657,N_30797);
nor U34793 (N_34793,N_30113,N_31291);
and U34794 (N_34794,N_30271,N_32116);
xor U34795 (N_34795,N_31380,N_31089);
nand U34796 (N_34796,N_32370,N_32427);
or U34797 (N_34797,N_32110,N_30062);
xnor U34798 (N_34798,N_31040,N_32082);
nand U34799 (N_34799,N_31339,N_30603);
or U34800 (N_34800,N_31605,N_31156);
and U34801 (N_34801,N_31249,N_31463);
xor U34802 (N_34802,N_31712,N_32388);
xnor U34803 (N_34803,N_32411,N_32401);
and U34804 (N_34804,N_31008,N_31285);
or U34805 (N_34805,N_32433,N_32103);
nor U34806 (N_34806,N_32130,N_32079);
or U34807 (N_34807,N_30154,N_31089);
and U34808 (N_34808,N_31088,N_32460);
or U34809 (N_34809,N_32234,N_30115);
or U34810 (N_34810,N_30696,N_30779);
and U34811 (N_34811,N_30060,N_31868);
or U34812 (N_34812,N_30270,N_32152);
or U34813 (N_34813,N_30791,N_31904);
xnor U34814 (N_34814,N_31896,N_31104);
or U34815 (N_34815,N_30182,N_32131);
nand U34816 (N_34816,N_32452,N_31175);
or U34817 (N_34817,N_31837,N_31114);
nor U34818 (N_34818,N_32430,N_30034);
nor U34819 (N_34819,N_30718,N_30356);
nor U34820 (N_34820,N_30540,N_32400);
xnor U34821 (N_34821,N_30939,N_31899);
xnor U34822 (N_34822,N_31572,N_30418);
and U34823 (N_34823,N_30394,N_32163);
nand U34824 (N_34824,N_31969,N_32396);
xor U34825 (N_34825,N_30819,N_31740);
xnor U34826 (N_34826,N_30433,N_32140);
and U34827 (N_34827,N_30045,N_31969);
nand U34828 (N_34828,N_30075,N_30833);
and U34829 (N_34829,N_32102,N_30156);
nor U34830 (N_34830,N_31703,N_30109);
or U34831 (N_34831,N_31802,N_31796);
nor U34832 (N_34832,N_31566,N_32243);
and U34833 (N_34833,N_31970,N_30970);
xnor U34834 (N_34834,N_30016,N_30887);
or U34835 (N_34835,N_30294,N_31867);
nor U34836 (N_34836,N_32208,N_31061);
nand U34837 (N_34837,N_31313,N_31054);
or U34838 (N_34838,N_30924,N_32408);
nand U34839 (N_34839,N_30562,N_30822);
or U34840 (N_34840,N_30841,N_30846);
or U34841 (N_34841,N_30348,N_30449);
xnor U34842 (N_34842,N_30930,N_30718);
xor U34843 (N_34843,N_31746,N_31026);
and U34844 (N_34844,N_32161,N_31937);
and U34845 (N_34845,N_30607,N_32422);
and U34846 (N_34846,N_32316,N_32076);
and U34847 (N_34847,N_32007,N_30571);
nand U34848 (N_34848,N_31873,N_31340);
or U34849 (N_34849,N_30116,N_30143);
or U34850 (N_34850,N_31432,N_30154);
and U34851 (N_34851,N_32438,N_32497);
or U34852 (N_34852,N_32257,N_31844);
or U34853 (N_34853,N_30899,N_32087);
nor U34854 (N_34854,N_30407,N_32246);
nand U34855 (N_34855,N_30800,N_31631);
xor U34856 (N_34856,N_31233,N_32057);
xor U34857 (N_34857,N_31083,N_32432);
nor U34858 (N_34858,N_31086,N_30189);
or U34859 (N_34859,N_30957,N_30525);
nand U34860 (N_34860,N_31801,N_31665);
or U34861 (N_34861,N_31076,N_30050);
nor U34862 (N_34862,N_30204,N_30739);
or U34863 (N_34863,N_31694,N_30793);
or U34864 (N_34864,N_31545,N_31206);
nor U34865 (N_34865,N_32430,N_30973);
xnor U34866 (N_34866,N_31805,N_30467);
or U34867 (N_34867,N_31115,N_31699);
nor U34868 (N_34868,N_30971,N_31537);
nor U34869 (N_34869,N_31622,N_31252);
or U34870 (N_34870,N_31677,N_30917);
or U34871 (N_34871,N_30732,N_32347);
xnor U34872 (N_34872,N_30899,N_32281);
nor U34873 (N_34873,N_30510,N_32003);
and U34874 (N_34874,N_32055,N_30079);
and U34875 (N_34875,N_30596,N_32474);
and U34876 (N_34876,N_30262,N_32419);
nor U34877 (N_34877,N_31232,N_31445);
nand U34878 (N_34878,N_31362,N_30739);
and U34879 (N_34879,N_31876,N_30815);
nor U34880 (N_34880,N_31823,N_31015);
xor U34881 (N_34881,N_30969,N_31794);
nor U34882 (N_34882,N_30719,N_30196);
nand U34883 (N_34883,N_30890,N_30008);
and U34884 (N_34884,N_31206,N_31934);
and U34885 (N_34885,N_32348,N_30316);
and U34886 (N_34886,N_31532,N_31776);
nand U34887 (N_34887,N_31361,N_32005);
nor U34888 (N_34888,N_31252,N_30357);
and U34889 (N_34889,N_30994,N_30769);
and U34890 (N_34890,N_31401,N_31528);
nor U34891 (N_34891,N_30676,N_30079);
xor U34892 (N_34892,N_30311,N_32405);
xor U34893 (N_34893,N_30320,N_31755);
nand U34894 (N_34894,N_30614,N_32214);
nand U34895 (N_34895,N_31136,N_30804);
and U34896 (N_34896,N_30645,N_31856);
nand U34897 (N_34897,N_31104,N_30827);
xor U34898 (N_34898,N_30347,N_30975);
nand U34899 (N_34899,N_31266,N_31706);
or U34900 (N_34900,N_30484,N_30396);
nand U34901 (N_34901,N_32448,N_30928);
or U34902 (N_34902,N_31002,N_31129);
nand U34903 (N_34903,N_31182,N_31404);
nor U34904 (N_34904,N_31231,N_31244);
nor U34905 (N_34905,N_31812,N_31751);
nor U34906 (N_34906,N_32294,N_32087);
xnor U34907 (N_34907,N_31056,N_31545);
or U34908 (N_34908,N_31760,N_31640);
nor U34909 (N_34909,N_30504,N_31384);
and U34910 (N_34910,N_30856,N_31376);
xnor U34911 (N_34911,N_30925,N_32108);
xnor U34912 (N_34912,N_31699,N_30197);
nor U34913 (N_34913,N_30184,N_31703);
nor U34914 (N_34914,N_30525,N_32185);
nand U34915 (N_34915,N_30108,N_32426);
and U34916 (N_34916,N_31510,N_32082);
or U34917 (N_34917,N_31634,N_31856);
xor U34918 (N_34918,N_32047,N_30899);
or U34919 (N_34919,N_32112,N_30994);
nand U34920 (N_34920,N_30564,N_31919);
and U34921 (N_34921,N_30534,N_32438);
and U34922 (N_34922,N_31120,N_31721);
nor U34923 (N_34923,N_31903,N_30912);
xor U34924 (N_34924,N_30569,N_32133);
nand U34925 (N_34925,N_30790,N_32432);
and U34926 (N_34926,N_30500,N_31958);
and U34927 (N_34927,N_30677,N_30289);
or U34928 (N_34928,N_30720,N_30202);
or U34929 (N_34929,N_31574,N_31930);
or U34930 (N_34930,N_30974,N_30380);
xor U34931 (N_34931,N_31822,N_31669);
xor U34932 (N_34932,N_31607,N_30705);
or U34933 (N_34933,N_30201,N_30892);
or U34934 (N_34934,N_30076,N_30854);
or U34935 (N_34935,N_30887,N_30029);
or U34936 (N_34936,N_32092,N_30300);
nor U34937 (N_34937,N_31149,N_30840);
or U34938 (N_34938,N_32118,N_32341);
nand U34939 (N_34939,N_31246,N_31430);
nor U34940 (N_34940,N_31512,N_31828);
nand U34941 (N_34941,N_31707,N_31351);
and U34942 (N_34942,N_31255,N_31478);
nor U34943 (N_34943,N_31001,N_31445);
xnor U34944 (N_34944,N_30559,N_31873);
or U34945 (N_34945,N_30225,N_32295);
or U34946 (N_34946,N_31560,N_31711);
xnor U34947 (N_34947,N_31520,N_32490);
xnor U34948 (N_34948,N_31274,N_32063);
and U34949 (N_34949,N_32199,N_32318);
nand U34950 (N_34950,N_31830,N_31250);
nor U34951 (N_34951,N_30731,N_32181);
and U34952 (N_34952,N_30034,N_30954);
and U34953 (N_34953,N_30623,N_31729);
and U34954 (N_34954,N_30826,N_30128);
xnor U34955 (N_34955,N_31502,N_31345);
nand U34956 (N_34956,N_30357,N_30207);
and U34957 (N_34957,N_31659,N_31299);
nand U34958 (N_34958,N_30732,N_32334);
and U34959 (N_34959,N_30874,N_31506);
or U34960 (N_34960,N_30158,N_31941);
nor U34961 (N_34961,N_30756,N_30497);
nand U34962 (N_34962,N_31602,N_30717);
and U34963 (N_34963,N_30823,N_30116);
xnor U34964 (N_34964,N_32442,N_30054);
or U34965 (N_34965,N_32149,N_30973);
and U34966 (N_34966,N_30176,N_31553);
nand U34967 (N_34967,N_30774,N_31135);
nand U34968 (N_34968,N_31498,N_31560);
and U34969 (N_34969,N_31613,N_31268);
nor U34970 (N_34970,N_30895,N_30821);
nand U34971 (N_34971,N_32099,N_31729);
nor U34972 (N_34972,N_31323,N_32460);
nand U34973 (N_34973,N_31274,N_30962);
nor U34974 (N_34974,N_31647,N_31279);
nor U34975 (N_34975,N_30034,N_31385);
and U34976 (N_34976,N_30295,N_32015);
nor U34977 (N_34977,N_31892,N_32187);
nor U34978 (N_34978,N_31062,N_30958);
xnor U34979 (N_34979,N_30755,N_30877);
or U34980 (N_34980,N_32291,N_31878);
and U34981 (N_34981,N_32207,N_30286);
xor U34982 (N_34982,N_30002,N_30149);
and U34983 (N_34983,N_31630,N_30989);
xor U34984 (N_34984,N_30442,N_31025);
nand U34985 (N_34985,N_32217,N_31932);
nor U34986 (N_34986,N_32176,N_30858);
nor U34987 (N_34987,N_31833,N_32250);
nand U34988 (N_34988,N_31785,N_30899);
or U34989 (N_34989,N_32153,N_30391);
xnor U34990 (N_34990,N_31974,N_30289);
or U34991 (N_34991,N_31370,N_31436);
xor U34992 (N_34992,N_31649,N_31100);
or U34993 (N_34993,N_31009,N_31274);
and U34994 (N_34994,N_31940,N_30159);
nor U34995 (N_34995,N_30999,N_30800);
nand U34996 (N_34996,N_30215,N_30071);
nand U34997 (N_34997,N_31294,N_31625);
and U34998 (N_34998,N_30312,N_31145);
nand U34999 (N_34999,N_32483,N_30896);
nand U35000 (N_35000,N_34700,N_33107);
or U35001 (N_35001,N_33694,N_34157);
and U35002 (N_35002,N_32923,N_34757);
or U35003 (N_35003,N_33366,N_33248);
nand U35004 (N_35004,N_33231,N_33307);
nor U35005 (N_35005,N_33762,N_32889);
nor U35006 (N_35006,N_33162,N_34169);
nand U35007 (N_35007,N_33190,N_34775);
and U35008 (N_35008,N_34866,N_33939);
nand U35009 (N_35009,N_33625,N_32806);
xor U35010 (N_35010,N_34779,N_32868);
and U35011 (N_35011,N_33518,N_33673);
xnor U35012 (N_35012,N_34140,N_34831);
nor U35013 (N_35013,N_33166,N_32662);
and U35014 (N_35014,N_34354,N_33665);
nand U35015 (N_35015,N_33770,N_33956);
nor U35016 (N_35016,N_34351,N_34171);
xnor U35017 (N_35017,N_34980,N_33968);
nand U35018 (N_35018,N_34764,N_34395);
nand U35019 (N_35019,N_33328,N_33500);
xnor U35020 (N_35020,N_33083,N_33360);
nor U35021 (N_35021,N_34122,N_34071);
and U35022 (N_35022,N_32879,N_33646);
xor U35023 (N_35023,N_33460,N_33918);
nand U35024 (N_35024,N_32911,N_33268);
nor U35025 (N_35025,N_34698,N_33846);
nand U35026 (N_35026,N_32731,N_34227);
xor U35027 (N_35027,N_34151,N_34417);
nand U35028 (N_35028,N_34943,N_33041);
and U35029 (N_35029,N_32636,N_34902);
nand U35030 (N_35030,N_34492,N_33862);
or U35031 (N_35031,N_34975,N_32899);
or U35032 (N_35032,N_33908,N_33821);
xnor U35033 (N_35033,N_32577,N_33005);
xnor U35034 (N_35034,N_34162,N_32690);
nor U35035 (N_35035,N_33829,N_32574);
xnor U35036 (N_35036,N_33783,N_33937);
or U35037 (N_35037,N_34655,N_33733);
nor U35038 (N_35038,N_34020,N_33828);
or U35039 (N_35039,N_34285,N_34794);
nand U35040 (N_35040,N_34480,N_33418);
xor U35041 (N_35041,N_32721,N_32750);
nor U35042 (N_35042,N_33597,N_33156);
nand U35043 (N_35043,N_32648,N_34997);
nand U35044 (N_35044,N_32743,N_32878);
and U35045 (N_35045,N_32762,N_32964);
and U35046 (N_35046,N_34042,N_33557);
xor U35047 (N_35047,N_34188,N_34015);
nor U35048 (N_35048,N_33061,N_32931);
and U35049 (N_35049,N_32585,N_34881);
nor U35050 (N_35050,N_34561,N_34033);
or U35051 (N_35051,N_34334,N_34663);
nand U35052 (N_35052,N_32999,N_33046);
and U35053 (N_35053,N_34961,N_34130);
or U35054 (N_35054,N_34359,N_33697);
nor U35055 (N_35055,N_34010,N_33115);
nand U35056 (N_35056,N_34954,N_32759);
nand U35057 (N_35057,N_33075,N_34948);
xor U35058 (N_35058,N_33813,N_33320);
or U35059 (N_35059,N_33359,N_33613);
and U35060 (N_35060,N_33066,N_33547);
and U35061 (N_35061,N_33852,N_32726);
xor U35062 (N_35062,N_34703,N_32888);
or U35063 (N_35063,N_32920,N_34725);
and U35064 (N_35064,N_33870,N_34360);
xnor U35065 (N_35065,N_34545,N_33837);
nor U35066 (N_35066,N_34059,N_33825);
xor U35067 (N_35067,N_32967,N_34898);
and U35068 (N_35068,N_32781,N_33634);
xnor U35069 (N_35069,N_33093,N_34910);
nand U35070 (N_35070,N_33630,N_34892);
xnor U35071 (N_35071,N_34842,N_34267);
and U35072 (N_35072,N_33163,N_34614);
nand U35073 (N_35073,N_34812,N_33244);
xnor U35074 (N_35074,N_33324,N_34032);
or U35075 (N_35075,N_34949,N_34308);
nor U35076 (N_35076,N_34502,N_34557);
or U35077 (N_35077,N_32563,N_34973);
nand U35078 (N_35078,N_34235,N_34255);
nand U35079 (N_35079,N_33384,N_32504);
nand U35080 (N_35080,N_34826,N_33127);
xor U35081 (N_35081,N_33032,N_32582);
or U35082 (N_35082,N_34891,N_33759);
nand U35083 (N_35083,N_33310,N_33144);
or U35084 (N_35084,N_33885,N_34079);
or U35085 (N_35085,N_33406,N_34011);
or U35086 (N_35086,N_34905,N_34486);
xnor U35087 (N_35087,N_33443,N_33065);
xnor U35088 (N_35088,N_34497,N_33602);
xor U35089 (N_35089,N_34542,N_33021);
or U35090 (N_35090,N_32604,N_34560);
and U35091 (N_35091,N_34265,N_34202);
and U35092 (N_35092,N_34726,N_34860);
nor U35093 (N_35093,N_32699,N_33534);
nor U35094 (N_35094,N_34463,N_33844);
nor U35095 (N_35095,N_33346,N_34924);
nand U35096 (N_35096,N_32698,N_32768);
xor U35097 (N_35097,N_33209,N_32561);
nand U35098 (N_35098,N_33139,N_34719);
and U35099 (N_35099,N_32834,N_33708);
nand U35100 (N_35100,N_33342,N_34735);
xnor U35101 (N_35101,N_33578,N_34107);
xor U35102 (N_35102,N_34294,N_34582);
and U35103 (N_35103,N_34134,N_32681);
nand U35104 (N_35104,N_32847,N_32505);
nand U35105 (N_35105,N_33878,N_34078);
and U35106 (N_35106,N_33680,N_33619);
nand U35107 (N_35107,N_33028,N_33364);
and U35108 (N_35108,N_34843,N_34028);
nor U35109 (N_35109,N_34476,N_33283);
nor U35110 (N_35110,N_34013,N_32988);
or U35111 (N_35111,N_32831,N_34765);
nor U35112 (N_35112,N_33415,N_34581);
xor U35113 (N_35113,N_34318,N_33659);
xor U35114 (N_35114,N_33398,N_34710);
nor U35115 (N_35115,N_34408,N_33174);
xnor U35116 (N_35116,N_34845,N_33370);
or U35117 (N_35117,N_32620,N_33650);
and U35118 (N_35118,N_34858,N_34341);
nand U35119 (N_35119,N_34063,N_34236);
nor U35120 (N_35120,N_33161,N_33411);
nor U35121 (N_35121,N_34682,N_33027);
nand U35122 (N_35122,N_34196,N_34337);
xor U35123 (N_35123,N_34742,N_32863);
nand U35124 (N_35124,N_34529,N_34409);
nor U35125 (N_35125,N_32668,N_33631);
or U35126 (N_35126,N_34402,N_33591);
or U35127 (N_35127,N_34238,N_33254);
nand U35128 (N_35128,N_32793,N_33259);
or U35129 (N_35129,N_33577,N_32646);
nor U35130 (N_35130,N_33096,N_34664);
or U35131 (N_35131,N_33233,N_34615);
and U35132 (N_35132,N_33198,N_33172);
or U35133 (N_35133,N_33438,N_33258);
or U35134 (N_35134,N_32718,N_33405);
nor U35135 (N_35135,N_32894,N_33998);
and U35136 (N_35136,N_34180,N_33015);
xnor U35137 (N_35137,N_33285,N_33620);
xnor U35138 (N_35138,N_33347,N_33530);
nor U35139 (N_35139,N_34737,N_32785);
nor U35140 (N_35140,N_33805,N_34343);
xor U35141 (N_35141,N_32993,N_33593);
nor U35142 (N_35142,N_33736,N_34370);
nand U35143 (N_35143,N_33655,N_34142);
nand U35144 (N_35144,N_32776,N_34816);
nand U35145 (N_35145,N_32586,N_34548);
nand U35146 (N_35146,N_33705,N_34407);
or U35147 (N_35147,N_33752,N_33234);
or U35148 (N_35148,N_32873,N_33780);
or U35149 (N_35149,N_34984,N_32789);
xor U35150 (N_35150,N_34194,N_32805);
nand U35151 (N_35151,N_33463,N_32757);
nand U35152 (N_35152,N_34602,N_34822);
nor U35153 (N_35153,N_34808,N_33982);
nor U35154 (N_35154,N_34859,N_34484);
and U35155 (N_35155,N_34758,N_32573);
nor U35156 (N_35156,N_34031,N_33587);
nor U35157 (N_35157,N_34657,N_34190);
xnor U35158 (N_35158,N_33987,N_34218);
or U35159 (N_35159,N_34840,N_33187);
xor U35160 (N_35160,N_32675,N_34406);
nor U35161 (N_35161,N_34841,N_34524);
nand U35162 (N_35162,N_34959,N_32588);
nor U35163 (N_35163,N_34195,N_34623);
or U35164 (N_35164,N_34996,N_34897);
nor U35165 (N_35165,N_34233,N_33089);
xor U35166 (N_35166,N_33595,N_32772);
xnor U35167 (N_35167,N_34272,N_33175);
nor U35168 (N_35168,N_32915,N_32810);
or U35169 (N_35169,N_33961,N_33446);
and U35170 (N_35170,N_33922,N_33407);
or U35171 (N_35171,N_34451,N_33444);
xnor U35172 (N_35172,N_33815,N_34108);
nand U35173 (N_35173,N_33365,N_32853);
xnor U35174 (N_35174,N_33727,N_33910);
xor U35175 (N_35175,N_34818,N_34374);
nor U35176 (N_35176,N_33600,N_34823);
xor U35177 (N_35177,N_33873,N_33135);
xor U35178 (N_35178,N_34544,N_32867);
xnor U35179 (N_35179,N_33570,N_33473);
nor U35180 (N_35180,N_34471,N_33251);
xnor U35181 (N_35181,N_34029,N_33011);
and U35182 (N_35182,N_33349,N_34900);
nor U35183 (N_35183,N_32556,N_33303);
and U35184 (N_35184,N_33158,N_32942);
nand U35185 (N_35185,N_34634,N_33851);
or U35186 (N_35186,N_34639,N_33799);
or U35187 (N_35187,N_33062,N_34419);
nand U35188 (N_35188,N_33754,N_34391);
xor U35189 (N_35189,N_32935,N_34004);
and U35190 (N_35190,N_34378,N_34832);
or U35191 (N_35191,N_32859,N_34317);
nand U35192 (N_35192,N_32553,N_32602);
xor U35193 (N_35193,N_33865,N_33421);
xor U35194 (N_35194,N_33563,N_34938);
nand U35195 (N_35195,N_33753,N_33820);
nor U35196 (N_35196,N_33236,N_32749);
or U35197 (N_35197,N_33657,N_32579);
or U35198 (N_35198,N_34516,N_32877);
nand U35199 (N_35199,N_33008,N_33901);
or U35200 (N_35200,N_33986,N_34345);
nand U35201 (N_35201,N_33375,N_32539);
and U35202 (N_35202,N_33441,N_33566);
or U35203 (N_35203,N_34738,N_33401);
xor U35204 (N_35204,N_34751,N_33465);
xnor U35205 (N_35205,N_33149,N_33495);
nor U35206 (N_35206,N_32575,N_32804);
nand U35207 (N_35207,N_33179,N_32621);
nand U35208 (N_35208,N_34073,N_33911);
and U35209 (N_35209,N_34690,N_32732);
or U35210 (N_35210,N_32569,N_34076);
nor U35211 (N_35211,N_34104,N_32865);
or U35212 (N_35212,N_34643,N_34181);
nand U35213 (N_35213,N_33085,N_33105);
and U35214 (N_35214,N_34752,N_32947);
or U35215 (N_35215,N_33549,N_32609);
or U35216 (N_35216,N_33410,N_32565);
nor U35217 (N_35217,N_33608,N_33081);
nor U35218 (N_35218,N_32815,N_33648);
xnor U35219 (N_35219,N_32896,N_33408);
nand U35220 (N_35220,N_32850,N_34717);
nand U35221 (N_35221,N_32538,N_32811);
or U35222 (N_35222,N_34410,N_33433);
or U35223 (N_35223,N_34521,N_33833);
or U35224 (N_35224,N_33035,N_32783);
nor U35225 (N_35225,N_34509,N_33684);
or U35226 (N_35226,N_34712,N_33618);
and U35227 (N_35227,N_34929,N_32876);
nor U35228 (N_35228,N_33624,N_32858);
nor U35229 (N_35229,N_33314,N_33876);
or U35230 (N_35230,N_34242,N_34799);
nand U35231 (N_35231,N_34875,N_33031);
xnor U35232 (N_35232,N_34759,N_33138);
xor U35233 (N_35233,N_33100,N_33984);
nor U35234 (N_35234,N_33861,N_32827);
nand U35235 (N_35235,N_32832,N_34495);
or U35236 (N_35236,N_32587,N_32897);
and U35237 (N_35237,N_32734,N_32996);
nand U35238 (N_35238,N_34711,N_34763);
and U35239 (N_35239,N_33636,N_33670);
nor U35240 (N_35240,N_32821,N_32644);
and U35241 (N_35241,N_32851,N_33237);
and U35242 (N_35242,N_32818,N_33834);
nand U35243 (N_35243,N_34571,N_33751);
xor U35244 (N_35244,N_34393,N_34413);
xor U35245 (N_35245,N_32580,N_34443);
or U35246 (N_35246,N_33743,N_34479);
and U35247 (N_35247,N_34043,N_32870);
xor U35248 (N_35248,N_32583,N_32541);
and U35249 (N_35249,N_34784,N_33681);
and U35250 (N_35250,N_32963,N_33272);
xnor U35251 (N_35251,N_32977,N_32590);
nor U35252 (N_35252,N_33502,N_34780);
and U35253 (N_35253,N_32738,N_34999);
nand U35254 (N_35254,N_34325,N_32607);
or U35255 (N_35255,N_34120,N_34191);
nand U35256 (N_35256,N_33380,N_34065);
nor U35257 (N_35257,N_32930,N_33424);
xnor U35258 (N_35258,N_33275,N_32921);
nand U35259 (N_35259,N_33189,N_33420);
or U35260 (N_35260,N_34149,N_32519);
nor U35261 (N_35261,N_34610,N_33568);
and U35262 (N_35262,N_33044,N_34695);
or U35263 (N_35263,N_34767,N_34844);
nor U35264 (N_35264,N_33160,N_33353);
xnor U35265 (N_35265,N_34907,N_33909);
or U35266 (N_35266,N_34000,N_32518);
xnor U35267 (N_35267,N_33476,N_33839);
nor U35268 (N_35268,N_33094,N_34470);
nor U35269 (N_35269,N_33351,N_33579);
nor U35270 (N_35270,N_33131,N_32506);
nor U35271 (N_35271,N_33440,N_33246);
xor U35272 (N_35272,N_34716,N_34350);
nand U35273 (N_35273,N_32746,N_34981);
xnor U35274 (N_35274,N_33461,N_33567);
nand U35275 (N_35275,N_34885,N_34991);
nor U35276 (N_35276,N_33295,N_32702);
xor U35277 (N_35277,N_32927,N_32976);
nand U35278 (N_35278,N_33668,N_33777);
xor U35279 (N_35279,N_32562,N_34754);
and U35280 (N_35280,N_33504,N_33087);
and U35281 (N_35281,N_33039,N_34773);
xor U35282 (N_35282,N_33491,N_32720);
nand U35283 (N_35283,N_33776,N_34683);
and U35284 (N_35284,N_34290,N_32552);
nor U35285 (N_35285,N_32697,N_34675);
or U35286 (N_35286,N_32864,N_33835);
nand U35287 (N_35287,N_34075,N_33464);
xnor U35288 (N_35288,N_32844,N_33760);
and U35289 (N_35289,N_33626,N_33824);
or U35290 (N_35290,N_32535,N_34361);
nand U35291 (N_35291,N_32802,N_34913);
nor U35292 (N_35292,N_34173,N_33522);
xor U35293 (N_35293,N_34864,N_32660);
or U35294 (N_35294,N_33279,N_32592);
nand U35295 (N_35295,N_33981,N_34894);
and U35296 (N_35296,N_32980,N_34868);
nand U35297 (N_35297,N_32638,N_33999);
xor U35298 (N_35298,N_32756,N_33012);
and U35299 (N_35299,N_34048,N_34743);
nor U35300 (N_35300,N_33790,N_32900);
xor U35301 (N_35301,N_33706,N_32857);
or U35302 (N_35302,N_34925,N_32625);
xor U35303 (N_35303,N_32994,N_33963);
xnor U35304 (N_35304,N_34331,N_33419);
xnor U35305 (N_35305,N_32817,N_33068);
xnor U35306 (N_35306,N_33397,N_34183);
and U35307 (N_35307,N_34003,N_34454);
nor U35308 (N_35308,N_33853,N_33545);
nor U35309 (N_35309,N_34951,N_34204);
nand U35310 (N_35310,N_34126,N_33101);
nor U35311 (N_35311,N_34650,N_33583);
xor U35312 (N_35312,N_33073,N_34448);
xor U35313 (N_35313,N_34645,N_33651);
nor U35314 (N_35314,N_32689,N_33306);
and U35315 (N_35315,N_33084,N_34704);
xor U35316 (N_35316,N_34209,N_33764);
and U35317 (N_35317,N_33490,N_33818);
nand U35318 (N_35318,N_32528,N_34908);
nand U35319 (N_35319,N_34270,N_33304);
or U35320 (N_35320,N_34302,N_32544);
nor U35321 (N_35321,N_33123,N_33399);
nor U35322 (N_35322,N_34652,N_33535);
xor U35323 (N_35323,N_34187,N_34006);
or U35324 (N_35324,N_34261,N_34498);
xor U35325 (N_35325,N_34276,N_32595);
nand U35326 (N_35326,N_32924,N_34423);
or U35327 (N_35327,N_34117,N_34896);
or U35328 (N_35328,N_34568,N_32622);
nand U35329 (N_35329,N_33007,N_32839);
xnor U35330 (N_35330,N_32651,N_33803);
xnor U35331 (N_35331,N_33948,N_34632);
and U35332 (N_35332,N_32650,N_33675);
xnor U35333 (N_35333,N_34111,N_34802);
nor U35334 (N_35334,N_34340,N_33109);
and U35335 (N_35335,N_33677,N_33195);
xor U35336 (N_35336,N_33693,N_32707);
and U35337 (N_35337,N_33262,N_34356);
and U35338 (N_35338,N_33641,N_34586);
xnor U35339 (N_35339,N_34168,N_33121);
or U35340 (N_35340,N_34396,N_32502);
nand U35341 (N_35341,N_34186,N_34312);
nor U35342 (N_35342,N_33585,N_32775);
nor U35343 (N_35343,N_34329,N_33836);
xnor U35344 (N_35344,N_33886,N_32581);
nand U35345 (N_35345,N_33276,N_33991);
and U35346 (N_35346,N_32616,N_34430);
or U35347 (N_35347,N_33352,N_33294);
xnor U35348 (N_35348,N_33750,N_34167);
and U35349 (N_35349,N_33972,N_34333);
or U35350 (N_35350,N_32943,N_32658);
xor U35351 (N_35351,N_34640,N_34205);
nor U35352 (N_35352,N_34293,N_33746);
and U35353 (N_35353,N_34274,N_33962);
and U35354 (N_35354,N_33594,N_34332);
and U35355 (N_35355,N_33996,N_33792);
nand U35356 (N_35356,N_34551,N_34292);
nor U35357 (N_35357,N_34806,N_33967);
or U35358 (N_35358,N_34531,N_34523);
nand U35359 (N_35359,N_33219,N_32950);
nand U35360 (N_35360,N_33556,N_32531);
nor U35361 (N_35361,N_32686,N_34365);
nor U35362 (N_35362,N_32751,N_33945);
xnor U35363 (N_35363,N_33528,N_34254);
nor U35364 (N_35364,N_33270,N_34876);
xnor U35365 (N_35365,N_32797,N_34313);
or U35366 (N_35366,N_34347,N_32525);
and U35367 (N_35367,N_34110,N_34936);
nor U35368 (N_35368,N_34755,N_33337);
nand U35369 (N_35369,N_34785,N_33327);
nand U35370 (N_35370,N_34172,N_34095);
nand U35371 (N_35371,N_33652,N_34491);
and U35372 (N_35372,N_32706,N_33687);
and U35373 (N_35373,N_32796,N_34611);
nor U35374 (N_35374,N_33560,N_33954);
nand U35375 (N_35375,N_33212,N_33923);
xor U35376 (N_35376,N_34791,N_33800);
nand U35377 (N_35377,N_33590,N_33218);
xor U35378 (N_35378,N_32813,N_33763);
and U35379 (N_35379,N_34501,N_32514);
xnor U35380 (N_35380,N_34884,N_34930);
xnor U35381 (N_35381,N_32624,N_34661);
nor U35382 (N_35382,N_34715,N_34556);
xor U35383 (N_35383,N_33868,N_34621);
and U35384 (N_35384,N_33863,N_33915);
xor U35385 (N_35385,N_33305,N_34215);
or U35386 (N_35386,N_33511,N_34328);
or U35387 (N_35387,N_34965,N_33286);
and U35388 (N_35388,N_32856,N_32849);
xnor U35389 (N_35389,N_32882,N_34141);
nand U35390 (N_35390,N_34982,N_32803);
nor U35391 (N_35391,N_34554,N_33289);
nand U35392 (N_35392,N_34403,N_34239);
nor U35393 (N_35393,N_32778,N_33459);
nand U35394 (N_35394,N_34886,N_34024);
xnor U35395 (N_35395,N_32664,N_32767);
and U35396 (N_35396,N_34260,N_33113);
xnor U35397 (N_35397,N_33225,N_32559);
nor U35398 (N_35398,N_33313,N_32961);
or U35399 (N_35399,N_33730,N_34459);
and U35400 (N_35400,N_34899,N_33023);
nand U35401 (N_35401,N_34041,N_33335);
xor U35402 (N_35402,N_34072,N_33050);
or U35403 (N_35403,N_33729,N_33150);
nor U35404 (N_35404,N_33333,N_33637);
or U35405 (N_35405,N_32560,N_32808);
or U35406 (N_35406,N_33720,N_34462);
and U35407 (N_35407,N_32902,N_34916);
xor U35408 (N_35408,N_33284,N_34603);
nor U35409 (N_35409,N_32934,N_34833);
or U35410 (N_35410,N_33884,N_34390);
and U35411 (N_35411,N_32529,N_32536);
xor U35412 (N_35412,N_33060,N_32968);
xor U35413 (N_35413,N_33822,N_34879);
nor U35414 (N_35414,N_32672,N_33080);
and U35415 (N_35415,N_32833,N_33124);
or U35416 (N_35416,N_33321,N_32669);
or U35417 (N_35417,N_34164,N_33572);
nor U35418 (N_35418,N_32761,N_34852);
xnor U35419 (N_35419,N_34444,N_34414);
and U35420 (N_35420,N_33311,N_34871);
and U35421 (N_35421,N_33831,N_34372);
nand U35422 (N_35422,N_32945,N_33079);
and U35423 (N_35423,N_32615,N_34198);
nand U35424 (N_35424,N_32983,N_33809);
nor U35425 (N_35425,N_34804,N_33816);
and U35426 (N_35426,N_33819,N_33422);
and U35427 (N_35427,N_34051,N_33088);
xor U35428 (N_35428,N_33930,N_33718);
or U35429 (N_35429,N_33091,N_34979);
or U35430 (N_35430,N_34601,N_33728);
nor U35431 (N_35431,N_34320,N_33340);
nand U35432 (N_35432,N_34796,N_33747);
nor U35433 (N_35433,N_33806,N_33177);
or U35434 (N_35434,N_32752,N_33788);
or U35435 (N_35435,N_33723,N_34608);
nand U35436 (N_35436,N_34694,N_33848);
and U35437 (N_35437,N_33202,N_33781);
nor U35438 (N_35438,N_32954,N_34045);
xnor U35439 (N_35439,N_34283,N_33243);
nor U35440 (N_35440,N_34228,N_32612);
xnor U35441 (N_35441,N_33437,N_33067);
nand U35442 (N_35442,N_33377,N_33935);
and U35443 (N_35443,N_33389,N_34163);
nor U35444 (N_35444,N_34635,N_33741);
nor U35445 (N_35445,N_32830,N_33486);
xor U35446 (N_35446,N_32744,N_33562);
nor U35447 (N_35447,N_33374,N_34424);
or U35448 (N_35448,N_33971,N_34957);
xnor U35449 (N_35449,N_34809,N_33165);
or U35450 (N_35450,N_34555,N_34469);
nor U35451 (N_35451,N_33503,N_34125);
or U35452 (N_35452,N_33235,N_33390);
nor U35453 (N_35453,N_33843,N_33501);
or U35454 (N_35454,N_33735,N_33038);
nand U35455 (N_35455,N_34427,N_32820);
or U35456 (N_35456,N_32584,N_33558);
or U35457 (N_35457,N_32542,N_34705);
or U35458 (N_35458,N_34803,N_34506);
nand U35459 (N_35459,N_33581,N_34547);
and U35460 (N_35460,N_33249,N_33134);
and U35461 (N_35461,N_33238,N_34734);
and U35462 (N_35462,N_34097,N_34256);
and U35463 (N_35463,N_34622,N_34087);
and U35464 (N_35464,N_34849,N_33802);
nor U35465 (N_35465,N_32628,N_34418);
or U35466 (N_35466,N_33704,N_34231);
and U35467 (N_35467,N_34626,N_33462);
and U35468 (N_35468,N_34353,N_34472);
xor U35469 (N_35469,N_32769,N_34768);
nand U35470 (N_35470,N_34512,N_34566);
and U35471 (N_35471,N_34219,N_33951);
nor U35472 (N_35472,N_33940,N_33118);
or U35473 (N_35473,N_34727,N_34086);
and U35474 (N_35474,N_33457,N_34857);
or U35475 (N_35475,N_33055,N_33941);
nand U35476 (N_35476,N_32895,N_33669);
xor U35477 (N_35477,N_34932,N_33755);
xnor U35478 (N_35478,N_32957,N_33355);
and U35479 (N_35479,N_34373,N_34433);
or U35480 (N_35480,N_32667,N_32855);
xnor U35481 (N_35481,N_32666,N_34550);
and U35482 (N_35482,N_33223,N_34827);
nor U35483 (N_35483,N_32719,N_32837);
nor U35484 (N_35484,N_34128,N_34580);
nand U35485 (N_35485,N_34179,N_34289);
and U35486 (N_35486,N_34956,N_33309);
nor U35487 (N_35487,N_33858,N_33667);
and U35488 (N_35488,N_33542,N_34739);
nand U35489 (N_35489,N_32979,N_34678);
nand U35490 (N_35490,N_34624,N_34252);
and U35491 (N_35491,N_33879,N_33758);
and U35492 (N_35492,N_34945,N_34552);
nand U35493 (N_35493,N_34821,N_33932);
or U35494 (N_35494,N_34503,N_33512);
or U35495 (N_35495,N_34203,N_34952);
and U35496 (N_35496,N_34438,N_34940);
or U35497 (N_35497,N_33188,N_34025);
xnor U35498 (N_35498,N_32995,N_34528);
and U35499 (N_35499,N_33111,N_32825);
nand U35500 (N_35500,N_33707,N_33506);
xnor U35501 (N_35501,N_33642,N_34460);
nand U35502 (N_35502,N_33204,N_32645);
xor U35503 (N_35503,N_34339,N_33317);
xnor U35504 (N_35504,N_32774,N_34660);
nand U35505 (N_35505,N_34835,N_34654);
or U35506 (N_35506,N_33378,N_32986);
nor U35507 (N_35507,N_33871,N_34950);
and U35508 (N_35508,N_33510,N_32521);
or U35509 (N_35509,N_34686,N_33297);
nand U35510 (N_35510,N_34797,N_34279);
nor U35511 (N_35511,N_32543,N_33148);
and U35512 (N_35512,N_33617,N_34428);
nand U35513 (N_35513,N_34208,N_32677);
and U35514 (N_35514,N_34193,N_33756);
nand U35515 (N_35515,N_34630,N_34850);
nand U35516 (N_35516,N_33786,N_32619);
nor U35517 (N_35517,N_34371,N_32845);
nand U35518 (N_35518,N_32617,N_33523);
xnor U35519 (N_35519,N_34175,N_33592);
or U35520 (N_35520,N_33970,N_32601);
nor U35521 (N_35521,N_33344,N_34116);
or U35522 (N_35522,N_32652,N_33607);
xor U35523 (N_35523,N_34525,N_34605);
nand U35524 (N_35524,N_33287,N_34211);
nand U35525 (N_35525,N_34429,N_33348);
xnor U35526 (N_35526,N_33498,N_33966);
nor U35527 (N_35527,N_34490,N_34221);
and U35528 (N_35528,N_34310,N_34220);
nor U35529 (N_35529,N_33447,N_33383);
nand U35530 (N_35530,N_32630,N_33480);
and U35531 (N_35531,N_34667,N_34520);
nor U35532 (N_35532,N_33417,N_34536);
and U35533 (N_35533,N_34398,N_34250);
and U35534 (N_35534,N_34475,N_32823);
and U35535 (N_35535,N_32891,N_33382);
or U35536 (N_35536,N_33766,N_33678);
nand U35537 (N_35537,N_32912,N_33529);
or U35538 (N_35538,N_34919,N_32764);
xor U35539 (N_35539,N_34064,N_33125);
nand U35540 (N_35540,N_34201,N_34616);
nor U35541 (N_35541,N_34400,N_34848);
and U35542 (N_35542,N_34606,N_33725);
and U35543 (N_35543,N_34781,N_33610);
and U35544 (N_35544,N_32723,N_34062);
or U35545 (N_35545,N_32883,N_33404);
and U35546 (N_35546,N_34101,N_34699);
xor U35547 (N_35547,N_33102,N_34617);
nor U35548 (N_35548,N_34307,N_34507);
nor U35549 (N_35549,N_33748,N_33004);
and U35550 (N_35550,N_32936,N_32674);
or U35551 (N_35551,N_34129,N_33467);
xor U35552 (N_35552,N_34578,N_34264);
nand U35553 (N_35553,N_34185,N_34707);
nand U35554 (N_35554,N_32557,N_32753);
and U35555 (N_35555,N_32807,N_34105);
nand U35556 (N_35556,N_34970,N_32654);
xnor U35557 (N_35557,N_32773,N_34273);
nand U35558 (N_35558,N_32819,N_33092);
or U35559 (N_35559,N_33745,N_33672);
and U35560 (N_35560,N_33508,N_34156);
xnor U35561 (N_35561,N_34939,N_34769);
xor U35562 (N_35562,N_33639,N_34795);
and U35563 (N_35563,N_33881,N_33958);
xor U35564 (N_35564,N_34019,N_33025);
or U35565 (N_35565,N_32836,N_33864);
and U35566 (N_35566,N_33431,N_33278);
and U35567 (N_35567,N_34904,N_34364);
nand U35568 (N_35568,N_33450,N_34597);
xor U35569 (N_35569,N_34839,N_33663);
or U35570 (N_35570,N_32948,N_34213);
and U35571 (N_35571,N_34918,N_32969);
and U35572 (N_35572,N_33120,N_33964);
nor U35573 (N_35573,N_33676,N_33738);
and U35574 (N_35574,N_33331,N_34096);
nor U35575 (N_35575,N_34511,N_33173);
or U35576 (N_35576,N_32510,N_34680);
or U35577 (N_35577,N_32568,N_33761);
or U35578 (N_35578,N_34862,N_34044);
xor U35579 (N_35579,N_34587,N_33924);
xor U35580 (N_35580,N_33037,N_33367);
nand U35581 (N_35581,N_34311,N_34629);
nor U35582 (N_35582,N_34993,N_32974);
or U35583 (N_35583,N_33892,N_34455);
xnor U35584 (N_35584,N_34647,N_32729);
nor U35585 (N_35585,N_32787,N_32655);
nor U35586 (N_35586,N_32939,N_34701);
xor U35587 (N_35587,N_33622,N_32633);
xnor U35588 (N_35588,N_34434,N_33255);
or U35589 (N_35589,N_34483,N_34888);
nand U35590 (N_35590,N_34914,N_33721);
nor U35591 (N_35591,N_33596,N_33070);
nor U35592 (N_35592,N_34729,N_34057);
nor U35593 (N_35593,N_33214,N_34106);
or U35594 (N_35594,N_32500,N_34061);
and U35595 (N_35595,N_34607,N_33856);
xor U35596 (N_35596,N_34431,N_33427);
nor U35597 (N_35597,N_32545,N_33538);
xnor U35598 (N_35598,N_34281,N_33022);
nor U35599 (N_35599,N_32591,N_34596);
or U35600 (N_35600,N_34612,N_33726);
and U35601 (N_35601,N_33213,N_33638);
xnor U35602 (N_35602,N_34756,N_34671);
or U35603 (N_35603,N_34026,N_34405);
and U35604 (N_35604,N_33606,N_33053);
or U35605 (N_35605,N_32940,N_33614);
nand U35606 (N_35606,N_33564,N_32755);
nand U35607 (N_35607,N_33994,N_34466);
nor U35608 (N_35608,N_34633,N_34732);
xnor U35609 (N_35609,N_34314,N_33488);
xnor U35610 (N_35610,N_33507,N_34309);
xnor U35611 (N_35611,N_34184,N_34066);
nor U35612 (N_35612,N_32880,N_32599);
nand U35613 (N_35613,N_34745,N_33713);
xor U35614 (N_35614,N_34085,N_33778);
and U35615 (N_35615,N_34054,N_34324);
or U35616 (N_35616,N_33387,N_33656);
or U35617 (N_35617,N_34001,N_32712);
or U35618 (N_35618,N_32843,N_33904);
nor U35619 (N_35619,N_33559,N_33171);
nand U35620 (N_35620,N_34872,N_34553);
or U35621 (N_35621,N_34214,N_32840);
nor U35622 (N_35622,N_33773,N_34146);
nor U35623 (N_35623,N_33413,N_33629);
and U35624 (N_35624,N_33301,N_34911);
nor U35625 (N_35625,N_33808,N_33095);
nor U35626 (N_35626,N_34182,N_33553);
nand U35627 (N_35627,N_34200,N_33071);
or U35628 (N_35628,N_33797,N_33042);
xor U35629 (N_35629,N_34549,N_32709);
and U35630 (N_35630,N_34666,N_34793);
nor U35631 (N_35631,N_34144,N_33731);
nand U35632 (N_35632,N_34800,N_32786);
and U35633 (N_35633,N_34599,N_33040);
and U35634 (N_35634,N_32593,N_33811);
or U35635 (N_35635,N_34246,N_34411);
xnor U35636 (N_35636,N_32713,N_34224);
or U35637 (N_35637,N_34636,N_34225);
xnor U35638 (N_35638,N_33143,N_33318);
nand U35639 (N_35639,N_34247,N_32741);
or U35640 (N_35640,N_32779,N_33580);
and U35641 (N_35641,N_33152,N_33700);
or U35642 (N_35642,N_33526,N_33900);
or U35643 (N_35643,N_34790,N_34969);
xnor U35644 (N_35644,N_32716,N_34517);
xor U35645 (N_35645,N_33855,N_34977);
or U35646 (N_35646,N_33423,N_32605);
or U35647 (N_35647,N_32784,N_33322);
nand U35648 (N_35648,N_33154,N_34148);
xnor U35649 (N_35649,N_32606,N_34232);
nor U35650 (N_35650,N_32949,N_34047);
or U35651 (N_35651,N_33182,N_34197);
nand U35652 (N_35652,N_33122,N_33810);
and U35653 (N_35653,N_34216,N_34113);
or U35654 (N_35654,N_34592,N_32670);
or U35655 (N_35655,N_33169,N_33226);
xnor U35656 (N_35656,N_33787,N_34305);
xnor U35657 (N_35657,N_34967,N_34514);
xor U35658 (N_35658,N_33944,N_34522);
nor U35659 (N_35659,N_32696,N_34641);
nand U35660 (N_35660,N_34008,N_34383);
nand U35661 (N_35661,N_34697,N_32507);
and U35662 (N_35662,N_33034,N_34138);
nor U35663 (N_35663,N_34733,N_34222);
nor U35664 (N_35664,N_33859,N_34420);
nand U35665 (N_35665,N_34882,N_34335);
xor U35666 (N_35666,N_34159,N_32814);
xor U35667 (N_35667,N_34384,N_33099);
xnor U35668 (N_35668,N_32710,N_34619);
xnor U35669 (N_35669,N_34212,N_34338);
and U35670 (N_35670,N_34326,N_32649);
nor U35671 (N_35671,N_33782,N_34367);
nor U35672 (N_35672,N_33576,N_32910);
nand U35673 (N_35673,N_34090,N_34016);
or U35674 (N_35674,N_33645,N_33357);
xor U35675 (N_35675,N_34099,N_33319);
nor U35676 (N_35676,N_34718,N_32922);
xnor U35677 (N_35677,N_34357,N_33582);
nand U35678 (N_35678,N_32608,N_33605);
or U35679 (N_35679,N_34493,N_33076);
nor U35680 (N_35680,N_34810,N_33376);
or U35681 (N_35681,N_33477,N_34576);
xor U35682 (N_35682,N_33795,N_33975);
and U35683 (N_35683,N_32705,N_34838);
nand U35684 (N_35684,N_32941,N_32929);
nor U35685 (N_35685,N_34853,N_33448);
and U35686 (N_35686,N_34268,N_34994);
or U35687 (N_35687,N_33906,N_33045);
and U35688 (N_35688,N_33789,N_33882);
or U35689 (N_35689,N_34206,N_34668);
nor U35690 (N_35690,N_34154,N_32687);
and U35691 (N_35691,N_33009,N_33356);
and U35692 (N_35692,N_34692,N_33548);
and U35693 (N_35693,N_34934,N_32801);
nand U35694 (N_35694,N_34263,N_34135);
nand U35695 (N_35695,N_34753,N_34487);
nand U35696 (N_35696,N_34777,N_34449);
nand U35697 (N_35697,N_33300,N_33264);
xor U35698 (N_35698,N_34296,N_34591);
xnor U35699 (N_35699,N_34673,N_34983);
and U35700 (N_35700,N_32511,N_33184);
nor U35701 (N_35701,N_34713,N_33628);
nand U35702 (N_35702,N_33658,N_33888);
nor U35703 (N_35703,N_34771,N_34145);
nor U35704 (N_35704,N_33779,N_32892);
or U35705 (N_35705,N_33221,N_33838);
or U35706 (N_35706,N_33997,N_34659);
xor U35707 (N_35707,N_33867,N_34518);
xnor U35708 (N_35708,N_33992,N_33897);
or U35709 (N_35709,N_34249,N_33361);
xor U35710 (N_35710,N_34458,N_34942);
nor U35711 (N_35711,N_33960,N_34342);
xor U35712 (N_35712,N_33203,N_33555);
nor U35713 (N_35713,N_32862,N_33449);
and U35714 (N_35714,N_34778,N_32736);
nand U35715 (N_35715,N_32551,N_33929);
and U35716 (N_35716,N_32975,N_33719);
or U35717 (N_35717,N_33242,N_33716);
or U35718 (N_35718,N_34869,N_33271);
nor U35719 (N_35719,N_33117,N_34160);
xnor U35720 (N_35720,N_33442,N_34579);
or U35721 (N_35721,N_34161,N_33372);
and U35722 (N_35722,N_34322,N_34241);
or U35723 (N_35723,N_32635,N_34052);
or U35724 (N_35724,N_33739,N_33493);
or U35725 (N_35725,N_33126,N_34344);
or U35726 (N_35726,N_33018,N_34123);
nor U35727 (N_35727,N_34895,N_33640);
nor U35728 (N_35728,N_34112,N_33426);
xor U35729 (N_35729,N_33691,N_33540);
nand U35730 (N_35730,N_34432,N_32860);
nor U35731 (N_35731,N_33296,N_34955);
and U35732 (N_35732,N_34789,N_33765);
nor U35733 (N_35733,N_34102,N_33842);
nor U35734 (N_35734,N_32523,N_33823);
nand U35735 (N_35735,N_34585,N_33920);
or U35736 (N_35736,N_33230,N_32788);
xnor U35737 (N_35737,N_32984,N_34829);
or U35738 (N_35738,N_33492,N_32770);
nor U35739 (N_35739,N_34741,N_33280);
or U35740 (N_35740,N_33841,N_33191);
xnor U35741 (N_35741,N_33598,N_32626);
nand U35742 (N_35742,N_33985,N_33452);
nand U35743 (N_35743,N_34702,N_34262);
nor U35744 (N_35744,N_34288,N_33489);
nor U35745 (N_35745,N_33260,N_34681);
nand U35746 (N_35746,N_33524,N_34127);
and U35747 (N_35747,N_33388,N_34750);
or U35748 (N_35748,N_34620,N_32515);
and U35749 (N_35749,N_33051,N_33153);
nand U35750 (N_35750,N_34847,N_34192);
and U35751 (N_35751,N_33277,N_33394);
nor U35752 (N_35752,N_33588,N_32991);
nand U35753 (N_35753,N_33481,N_34189);
xor U35754 (N_35754,N_33653,N_34590);
and U35755 (N_35755,N_33519,N_33575);
xnor U35756 (N_35756,N_32846,N_34389);
xor U35757 (N_35757,N_33181,N_33108);
and U35758 (N_35758,N_32763,N_33024);
xor U35759 (N_35759,N_33057,N_33474);
and U35760 (N_35760,N_34909,N_33895);
nand U35761 (N_35761,N_33902,N_34820);
nor U35762 (N_35762,N_32627,N_33141);
and U35763 (N_35763,N_33217,N_32597);
nor U35764 (N_35764,N_33543,N_32678);
nor U35765 (N_35765,N_34230,N_34685);
or U35766 (N_35766,N_32632,N_32639);
xnor U35767 (N_35767,N_33774,N_34399);
or U35768 (N_35768,N_34447,N_32998);
and U35769 (N_35769,N_34446,N_34022);
nand U35770 (N_35770,N_34837,N_34094);
xnor U35771 (N_35771,N_32997,N_32509);
and U35772 (N_35772,N_34226,N_34987);
xor U35773 (N_35773,N_34243,N_33054);
nand U35774 (N_35774,N_32904,N_32503);
or U35775 (N_35775,N_34985,N_34473);
xnor U35776 (N_35776,N_32671,N_32566);
nand U35777 (N_35777,N_34093,N_32916);
xnor U35778 (N_35778,N_32693,N_32682);
or U35779 (N_35779,N_34388,N_32780);
nor U35780 (N_35780,N_33724,N_33257);
nor U35781 (N_35781,N_33468,N_33332);
and U35782 (N_35782,N_33827,N_33647);
and U35783 (N_35783,N_32659,N_34824);
nand U35784 (N_35784,N_33159,N_34060);
nor U35785 (N_35785,N_34917,N_34880);
xor U35786 (N_35786,N_34382,N_33064);
xor U35787 (N_35787,N_33281,N_33969);
nor U35788 (N_35788,N_33471,N_33403);
xor U35789 (N_35789,N_33216,N_32647);
and U35790 (N_35790,N_34662,N_33400);
nand U35791 (N_35791,N_33458,N_33905);
xnor U35792 (N_35792,N_33269,N_33402);
xor U35793 (N_35793,N_33058,N_32946);
nor U35794 (N_35794,N_34723,N_32717);
xnor U35795 (N_35795,N_34257,N_34836);
or U35796 (N_35796,N_32782,N_34762);
and U35797 (N_35797,N_34761,N_34494);
nand U35798 (N_35798,N_34363,N_32962);
xor U35799 (N_35799,N_34152,N_32951);
nor U35800 (N_35800,N_32533,N_34595);
xnor U35801 (N_35801,N_33010,N_32903);
nand U35802 (N_35802,N_32727,N_34990);
and U35803 (N_35803,N_34121,N_32596);
or U35804 (N_35804,N_34366,N_32637);
and U35805 (N_35805,N_32676,N_33206);
and U35806 (N_35806,N_33469,N_34968);
xor U35807 (N_35807,N_33699,N_33049);
or U35808 (N_35808,N_34574,N_34223);
and U35809 (N_35809,N_33455,N_33052);
or U35810 (N_35810,N_34251,N_34485);
or U35811 (N_35811,N_34628,N_32982);
nor U35812 (N_35812,N_32854,N_34385);
xnor U35813 (N_35813,N_33913,N_33949);
or U35814 (N_35814,N_32826,N_33514);
and U35815 (N_35815,N_33315,N_34721);
and U35816 (N_35816,N_34131,N_34035);
nor U35817 (N_35817,N_33494,N_33302);
xor U35818 (N_35818,N_33925,N_33282);
nor U35819 (N_35819,N_33196,N_33688);
and U35820 (N_35820,N_32684,N_33439);
and U35821 (N_35821,N_33537,N_34327);
or U35822 (N_35822,N_33048,N_34625);
nand U35823 (N_35823,N_34137,N_33683);
or U35824 (N_35824,N_33267,N_32866);
nor U35825 (N_35825,N_33893,N_33561);
and U35826 (N_35826,N_33703,N_33266);
xnor U35827 (N_35827,N_33715,N_34558);
nor U35828 (N_35828,N_34627,N_33934);
xnor U35829 (N_35829,N_33544,N_34319);
or U35830 (N_35830,N_33955,N_33654);
xnor U35831 (N_35831,N_34760,N_33136);
nor U35832 (N_35832,N_33354,N_33976);
nor U35833 (N_35833,N_34946,N_33176);
nand U35834 (N_35834,N_32703,N_32598);
xnor U35835 (N_35835,N_32932,N_33466);
nor U35836 (N_35836,N_32800,N_34068);
xor U35837 (N_35837,N_34564,N_34677);
or U35838 (N_35838,N_33074,N_32908);
nand U35839 (N_35839,N_32971,N_33695);
nor U35840 (N_35840,N_34863,N_34380);
and U35841 (N_35841,N_32848,N_33199);
nor U35842 (N_35842,N_34807,N_34266);
and U35843 (N_35843,N_34854,N_34166);
nand U35844 (N_35844,N_33412,N_33527);
nand U35845 (N_35845,N_34783,N_33785);
or U35846 (N_35846,N_33090,N_34304);
nor U35847 (N_35847,N_34280,N_33261);
and U35848 (N_35848,N_34567,N_32642);
and U35849 (N_35849,N_32835,N_34375);
nand U35850 (N_35850,N_33145,N_34637);
or U35851 (N_35851,N_34259,N_32547);
or U35852 (N_35852,N_34002,N_32663);
and U35853 (N_35853,N_33409,N_34642);
or U35854 (N_35854,N_34034,N_34284);
nor U35855 (N_35855,N_33686,N_33767);
xor U35856 (N_35856,N_34609,N_33586);
xor U35857 (N_35857,N_34992,N_33180);
xor U35858 (N_35858,N_33146,N_33019);
nor U35859 (N_35859,N_32919,N_33211);
nand U35860 (N_35860,N_33814,N_34234);
and U35861 (N_35861,N_33849,N_32516);
or U35862 (N_35862,N_32838,N_33293);
and U35863 (N_35863,N_33616,N_33621);
nor U35864 (N_35864,N_33157,N_32754);
and U35865 (N_35865,N_32680,N_33599);
and U35866 (N_35866,N_33325,N_33186);
nor U35867 (N_35867,N_33740,N_34986);
and U35868 (N_35868,N_34543,N_34788);
or U35869 (N_35869,N_33644,N_33880);
nand U35870 (N_35870,N_34786,N_34776);
and U35871 (N_35871,N_33336,N_32603);
nand U35872 (N_35872,N_32555,N_33696);
and U35873 (N_35873,N_34050,N_34133);
or U35874 (N_35874,N_33036,N_33957);
nor U35875 (N_35875,N_33479,N_34749);
or U35876 (N_35876,N_34923,N_34040);
nand U35877 (N_35877,N_34541,N_32685);
nor U35878 (N_35878,N_32989,N_33170);
nand U35879 (N_35879,N_33980,N_34153);
and U35880 (N_35880,N_33482,N_34488);
nand U35881 (N_35881,N_33717,N_32885);
nand U35882 (N_35882,N_34787,N_33082);
and U35883 (N_35883,N_34962,N_32990);
xor U35884 (N_35884,N_34770,N_33928);
xnor U35885 (N_35885,N_33456,N_34593);
nor U35886 (N_35886,N_34736,N_33771);
nor U35887 (N_35887,N_32909,N_33988);
nand U35888 (N_35888,N_32972,N_33429);
nand U35889 (N_35889,N_34282,N_34510);
nand U35890 (N_35890,N_34974,N_34883);
and U35891 (N_35891,N_34588,N_34387);
or U35892 (N_35892,N_34158,N_33505);
and U35893 (N_35893,N_34728,N_33569);
and U35894 (N_35894,N_32907,N_33006);
xor U35895 (N_35895,N_34248,N_33395);
or U35896 (N_35896,N_34297,N_33002);
nand U35897 (N_35897,N_32799,N_34277);
or U35898 (N_35898,N_34782,N_34067);
nor U35899 (N_35899,N_33993,N_32589);
nor U35900 (N_35900,N_33445,N_32643);
xnor U35901 (N_35901,N_34489,N_34477);
xnor U35902 (N_35902,N_33205,N_33483);
nor U35903 (N_35903,N_33907,N_34442);
nor U35904 (N_35904,N_32890,N_33943);
nand U35905 (N_35905,N_33478,N_33874);
or U35906 (N_35906,N_34150,N_33298);
and U35907 (N_35907,N_34348,N_33983);
nand U35908 (N_35908,N_34530,N_34709);
or U35909 (N_35909,N_34538,N_34316);
nor U35910 (N_35910,N_33872,N_33509);
or U35911 (N_35911,N_34439,N_32558);
and U35912 (N_35912,N_33017,N_34963);
nand U35913 (N_35913,N_34689,N_33151);
and U35914 (N_35914,N_34873,N_34537);
or U35915 (N_35915,N_34798,N_33072);
nand U35916 (N_35916,N_34539,N_33817);
xnor U35917 (N_35917,N_33714,N_34583);
nand U35918 (N_35918,N_33147,N_32917);
and U35919 (N_35919,N_33611,N_33129);
or U35920 (N_35920,N_34825,N_33916);
xor U35921 (N_35921,N_33485,N_34014);
nand U35922 (N_35922,N_34656,N_32640);
and U35923 (N_35923,N_34766,N_33428);
nor U35924 (N_35924,N_34527,N_32540);
or U35925 (N_35925,N_34174,N_33210);
and U35926 (N_35926,N_33973,N_33536);
or U35927 (N_35927,N_33043,N_34500);
xnor U35928 (N_35928,N_34613,N_34935);
and U35929 (N_35929,N_32520,N_34964);
and U35930 (N_35930,N_34594,N_34830);
nand U35931 (N_35931,N_33860,N_34253);
or U35932 (N_35932,N_32711,N_33030);
nor U35933 (N_35933,N_33950,N_33722);
xor U35934 (N_35934,N_34513,N_33430);
or U35935 (N_35935,N_34714,N_32944);
or U35936 (N_35936,N_34083,N_32841);
nand U35937 (N_35937,N_33551,N_32937);
and U35938 (N_35938,N_34377,N_34115);
nand U35939 (N_35939,N_34017,N_33168);
nand U35940 (N_35940,N_32634,N_32673);
and U35941 (N_35941,N_34275,N_34465);
or U35942 (N_35942,N_33350,N_33845);
xor U35943 (N_35943,N_34426,N_32955);
or U35944 (N_35944,N_33573,N_32735);
nand U35945 (N_35945,N_32795,N_32965);
nand U35946 (N_35946,N_33784,N_34998);
nor U35947 (N_35947,N_33252,N_33227);
nand U35948 (N_35948,N_32576,N_32522);
xnor U35949 (N_35949,N_34648,N_32960);
or U35950 (N_35950,N_33541,N_33097);
nand U35951 (N_35951,N_33671,N_33875);
nand U35952 (N_35952,N_33178,N_32884);
xnor U35953 (N_35953,N_34653,N_32874);
xnor U35954 (N_35954,N_34958,N_32905);
or U35955 (N_35955,N_33308,N_32881);
nor U35956 (N_35956,N_33215,N_33604);
xor U35957 (N_35957,N_32715,N_32708);
and U35958 (N_35958,N_32724,N_33959);
nand U35959 (N_35959,N_34920,N_32747);
or U35960 (N_35960,N_34394,N_33323);
xnor U35961 (N_35961,N_33942,N_34893);
nor U35962 (N_35962,N_33253,N_34688);
and U35963 (N_35963,N_34496,N_34291);
and U35964 (N_35964,N_33830,N_34358);
nand U35965 (N_35965,N_32614,N_34889);
or U35966 (N_35966,N_34132,N_33208);
or U35967 (N_35967,N_34672,N_33220);
and U35968 (N_35968,N_34481,N_32926);
nand U35969 (N_35969,N_32953,N_34912);
xnor U35970 (N_35970,N_33130,N_33358);
nand U35971 (N_35971,N_33453,N_33183);
or U35972 (N_35972,N_34676,N_34828);
or U35973 (N_35973,N_33167,N_32661);
xnor U35974 (N_35974,N_33768,N_32737);
nand U35975 (N_35975,N_34092,N_33240);
nand U35976 (N_35976,N_32739,N_34240);
xnor U35977 (N_35977,N_34009,N_32992);
nor U35978 (N_35978,N_34834,N_33917);
nand U35979 (N_35979,N_34244,N_33386);
and U35980 (N_35980,N_33393,N_34415);
and U35981 (N_35981,N_33373,N_34646);
nand U35982 (N_35982,N_33086,N_32554);
or U35983 (N_35983,N_32887,N_32567);
or U35984 (N_35984,N_32623,N_32546);
and U35985 (N_35985,N_33069,N_34404);
xnor U35986 (N_35986,N_33571,N_32760);
nor U35987 (N_35987,N_34928,N_33200);
and U35988 (N_35988,N_33931,N_34177);
nand U35989 (N_35989,N_33539,N_33470);
xnor U35990 (N_35990,N_33106,N_32594);
nor U35991 (N_35991,N_33273,N_34084);
xor U35992 (N_35992,N_34478,N_34056);
and U35993 (N_35993,N_33194,N_34526);
xor U35994 (N_35994,N_32537,N_32901);
and U35995 (N_35995,N_34878,N_33112);
xnor U35996 (N_35996,N_34575,N_32549);
nand U35997 (N_35997,N_33119,N_32842);
xor U35998 (N_35998,N_34301,N_34468);
nor U35999 (N_35999,N_34425,N_33516);
and U36000 (N_36000,N_34303,N_32524);
and U36001 (N_36001,N_32824,N_32914);
nor U36002 (N_36002,N_32527,N_34631);
nand U36003 (N_36003,N_32798,N_33487);
nor U36004 (N_36004,N_33000,N_33475);
nor U36005 (N_36005,N_33565,N_34401);
and U36006 (N_36006,N_33692,N_34801);
nand U36007 (N_36007,N_33685,N_33104);
or U36008 (N_36008,N_33978,N_33245);
or U36009 (N_36009,N_33635,N_34504);
xor U36010 (N_36010,N_32771,N_32701);
xor U36011 (N_36011,N_34598,N_33103);
and U36012 (N_36012,N_33222,N_34012);
nor U36013 (N_36013,N_33114,N_34947);
and U36014 (N_36014,N_34330,N_32700);
nand U36015 (N_36015,N_34467,N_32572);
or U36016 (N_36016,N_33927,N_34482);
or U36017 (N_36017,N_32790,N_34901);
or U36018 (N_36018,N_32657,N_34437);
xnor U36019 (N_36019,N_34944,N_33734);
and U36020 (N_36020,N_33265,N_33520);
or U36021 (N_36021,N_33749,N_33291);
xor U36022 (N_36022,N_33737,N_34210);
nand U36023 (N_36023,N_33496,N_34708);
and U36024 (N_36024,N_32611,N_34805);
or U36025 (N_36025,N_34971,N_34369);
or U36026 (N_36026,N_34819,N_32913);
nand U36027 (N_36027,N_32526,N_32683);
xor U36028 (N_36028,N_34589,N_33334);
and U36029 (N_36029,N_33250,N_32722);
and U36030 (N_36030,N_33921,N_34368);
and U36031 (N_36031,N_33912,N_33142);
and U36032 (N_36032,N_34865,N_34315);
or U36033 (N_36033,N_33769,N_32688);
nor U36034 (N_36034,N_33026,N_33381);
nor U36035 (N_36035,N_33371,N_33603);
and U36036 (N_36036,N_33385,N_34147);
or U36037 (N_36037,N_34346,N_33247);
or U36038 (N_36038,N_33533,N_33702);
or U36039 (N_36039,N_34731,N_33001);
xor U36040 (N_36040,N_34665,N_34573);
nor U36041 (N_36041,N_32981,N_33938);
nor U36042 (N_36042,N_33363,N_34114);
nand U36043 (N_36043,N_34546,N_34505);
xnor U36044 (N_36044,N_34036,N_33232);
xor U36045 (N_36045,N_32641,N_33059);
nor U36046 (N_36046,N_33627,N_33263);
xor U36047 (N_36047,N_32872,N_34058);
nand U36048 (N_36048,N_34021,N_34813);
xor U36049 (N_36049,N_34397,N_33379);
nand U36050 (N_36050,N_34381,N_34815);
nand U36051 (N_36051,N_34461,N_33894);
and U36052 (N_36052,N_32875,N_33193);
and U36053 (N_36053,N_32618,N_34669);
xor U36054 (N_36054,N_34746,N_33840);
xnor U36055 (N_36055,N_34299,N_33343);
or U36056 (N_36056,N_33137,N_33229);
or U36057 (N_36057,N_34499,N_32777);
xor U36058 (N_36058,N_32629,N_34569);
xnor U36059 (N_36059,N_34091,N_34867);
and U36060 (N_36060,N_32973,N_34534);
and U36061 (N_36061,N_34855,N_32548);
or U36062 (N_36062,N_34978,N_33682);
or U36063 (N_36063,N_33432,N_34453);
xnor U36064 (N_36064,N_32829,N_34903);
nor U36065 (N_36065,N_33292,N_33228);
or U36066 (N_36066,N_33898,N_33133);
or U36067 (N_36067,N_34421,N_33609);
and U36068 (N_36068,N_34861,N_32694);
or U36069 (N_36069,N_34456,N_34604);
and U36070 (N_36070,N_33003,N_34074);
nor U36071 (N_36071,N_34355,N_33077);
and U36072 (N_36072,N_32966,N_34870);
nor U36073 (N_36073,N_34298,N_33965);
and U36074 (N_36074,N_33451,N_34508);
nand U36075 (N_36075,N_34445,N_33857);
xor U36076 (N_36076,N_34748,N_33742);
xnor U36077 (N_36077,N_34972,N_34089);
nand U36078 (N_36078,N_34814,N_34519);
nand U36079 (N_36079,N_34271,N_34321);
nand U36080 (N_36080,N_33063,N_33974);
nand U36081 (N_36081,N_32714,N_33589);
nor U36082 (N_36082,N_34287,N_34098);
or U36083 (N_36083,N_33643,N_32631);
xor U36084 (N_36084,N_33056,N_34450);
or U36085 (N_36085,N_33391,N_33601);
xor U36086 (N_36086,N_33869,N_34295);
and U36087 (N_36087,N_34772,N_33701);
nand U36088 (N_36088,N_34258,N_33029);
xor U36089 (N_36089,N_32508,N_32653);
or U36090 (N_36090,N_32578,N_33812);
nand U36091 (N_36091,N_34687,N_33339);
nor U36092 (N_36092,N_34744,N_33484);
nor U36093 (N_36093,N_34720,N_33995);
and U36094 (N_36094,N_33047,N_33926);
nor U36095 (N_36095,N_33517,N_32534);
xnor U36096 (N_36096,N_34540,N_33632);
and U36097 (N_36097,N_33497,N_34535);
nor U36098 (N_36098,N_33532,N_33574);
nand U36099 (N_36099,N_34436,N_34651);
xor U36100 (N_36100,N_33513,N_33989);
nand U36101 (N_36101,N_32958,N_33661);
and U36102 (N_36102,N_32656,N_34452);
nand U36103 (N_36103,N_34435,N_33796);
nor U36104 (N_36104,N_34600,N_33854);
nand U36105 (N_36105,N_32550,N_33312);
and U36106 (N_36106,N_33531,N_32987);
nand U36107 (N_36107,N_34976,N_33241);
or U36108 (N_36108,N_32970,N_33435);
xnor U36109 (N_36109,N_33896,N_34740);
or U36110 (N_36110,N_34926,N_34136);
or U36111 (N_36111,N_33164,N_34100);
and U36112 (N_36112,N_34269,N_32513);
nand U36113 (N_36113,N_34670,N_32725);
or U36114 (N_36114,N_34199,N_33016);
and U36115 (N_36115,N_33369,N_33710);
and U36116 (N_36116,N_33525,N_34724);
or U36117 (N_36117,N_34927,N_34995);
xor U36118 (N_36118,N_33414,N_32501);
nor U36119 (N_36119,N_32740,N_33274);
or U36120 (N_36120,N_34207,N_33078);
and U36121 (N_36121,N_34440,N_34792);
or U36122 (N_36122,N_32906,N_33979);
and U36123 (N_36123,N_32695,N_32938);
and U36124 (N_36124,N_33368,N_33887);
or U36125 (N_36125,N_32517,N_33192);
nand U36126 (N_36126,N_33711,N_34464);
or U36127 (N_36127,N_34046,N_32816);
nor U36128 (N_36128,N_33877,N_33847);
or U36129 (N_36129,N_33936,N_33890);
nor U36130 (N_36130,N_32613,N_33801);
nand U36131 (N_36131,N_33649,N_34693);
and U36132 (N_36132,N_33014,N_34937);
xnor U36133 (N_36133,N_34379,N_33914);
and U36134 (N_36134,N_33804,N_34856);
nand U36135 (N_36135,N_32925,N_34577);
nand U36136 (N_36136,N_34877,N_33207);
xor U36137 (N_36137,N_33850,N_32861);
and U36138 (N_36138,N_34412,N_34921);
xnor U36139 (N_36139,N_32570,N_34649);
or U36140 (N_36140,N_33546,N_34037);
nand U36141 (N_36141,N_34070,N_34018);
xnor U36142 (N_36142,N_32959,N_33615);
or U36143 (N_36143,N_32852,N_34570);
nor U36144 (N_36144,N_33794,N_32765);
nor U36145 (N_36145,N_32728,N_34245);
nand U36146 (N_36146,N_32794,N_33709);
xor U36147 (N_36147,N_32745,N_34532);
nand U36148 (N_36148,N_34915,N_33140);
or U36149 (N_36149,N_34416,N_34696);
nand U36150 (N_36150,N_32691,N_34077);
nor U36151 (N_36151,N_34080,N_33757);
xor U36152 (N_36152,N_34306,N_33826);
xnor U36153 (N_36153,N_33919,N_34563);
and U36154 (N_36154,N_33454,N_33889);
or U36155 (N_36155,N_33633,N_34081);
xnor U36156 (N_36156,N_34644,N_34109);
nand U36157 (N_36157,N_34178,N_33330);
xnor U36158 (N_36158,N_33155,N_33550);
or U36159 (N_36159,N_33832,N_34286);
nor U36160 (N_36160,N_33947,N_32610);
nand U36161 (N_36161,N_33185,N_33866);
nor U36162 (N_36162,N_34039,N_34027);
or U36163 (N_36163,N_33807,N_34584);
and U36164 (N_36164,N_34055,N_33698);
nor U36165 (N_36165,N_33392,N_34722);
xor U36166 (N_36166,N_32933,N_32733);
nor U36167 (N_36167,N_32512,N_34941);
nor U36168 (N_36168,N_34165,N_33662);
or U36169 (N_36169,N_33033,N_33883);
nand U36170 (N_36170,N_34730,N_34572);
nand U36171 (N_36171,N_33116,N_34846);
nand U36172 (N_36172,N_32665,N_32978);
xor U36173 (N_36173,N_34217,N_34515);
or U36174 (N_36174,N_34392,N_33256);
nand U36175 (N_36175,N_34005,N_34082);
xor U36176 (N_36176,N_33201,N_34103);
and U36177 (N_36177,N_34376,N_32952);
xor U36178 (N_36178,N_33933,N_34562);
nor U36179 (N_36179,N_34906,N_34155);
and U36180 (N_36180,N_33013,N_33288);
nand U36181 (N_36181,N_32898,N_33674);
nor U36182 (N_36182,N_33791,N_34674);
or U36183 (N_36183,N_33666,N_34747);
nand U36184 (N_36184,N_32766,N_33396);
xor U36185 (N_36185,N_32812,N_34170);
xor U36186 (N_36186,N_34874,N_34922);
or U36187 (N_36187,N_32886,N_32758);
xor U36188 (N_36188,N_34887,N_34422);
nor U36189 (N_36189,N_32692,N_34229);
or U36190 (N_36190,N_34139,N_32564);
xor U36191 (N_36191,N_33554,N_32809);
xnor U36192 (N_36192,N_34007,N_34474);
or U36193 (N_36193,N_33132,N_33425);
nor U36194 (N_36194,N_34684,N_32985);
xnor U36195 (N_36195,N_32893,N_34336);
nand U36196 (N_36196,N_32792,N_34679);
xnor U36197 (N_36197,N_34023,N_33299);
nor U36198 (N_36198,N_33345,N_34989);
nand U36199 (N_36199,N_32791,N_32600);
nand U36200 (N_36200,N_32822,N_33798);
nand U36201 (N_36201,N_33472,N_34691);
or U36202 (N_36202,N_33362,N_33793);
xor U36203 (N_36203,N_33434,N_34300);
nand U36204 (N_36204,N_33552,N_33712);
nor U36205 (N_36205,N_34658,N_34811);
nor U36206 (N_36206,N_32571,N_33952);
nand U36207 (N_36207,N_33128,N_34176);
and U36208 (N_36208,N_34069,N_33903);
nand U36209 (N_36209,N_34124,N_33584);
xnor U36210 (N_36210,N_33690,N_34386);
xor U36211 (N_36211,N_32532,N_33953);
xnor U36212 (N_36212,N_34237,N_34851);
xnor U36213 (N_36213,N_33326,N_33197);
nor U36214 (N_36214,N_33416,N_34118);
nand U36215 (N_36215,N_34441,N_32748);
nand U36216 (N_36216,N_34457,N_34774);
nand U36217 (N_36217,N_33899,N_33977);
and U36218 (N_36218,N_34565,N_33664);
xor U36219 (N_36219,N_33290,N_34966);
nand U36220 (N_36220,N_33224,N_33338);
or U36221 (N_36221,N_32742,N_34323);
nand U36222 (N_36222,N_32918,N_34349);
and U36223 (N_36223,N_32871,N_34559);
or U36224 (N_36224,N_33020,N_34890);
nand U36225 (N_36225,N_34038,N_33744);
nand U36226 (N_36226,N_33891,N_33772);
xnor U36227 (N_36227,N_33499,N_34988);
xor U36228 (N_36228,N_33623,N_33689);
or U36229 (N_36229,N_34533,N_33521);
xor U36230 (N_36230,N_32704,N_34049);
or U36231 (N_36231,N_32869,N_34278);
xor U36232 (N_36232,N_34143,N_34088);
nor U36233 (N_36233,N_33679,N_33239);
xor U36234 (N_36234,N_33775,N_34618);
xnor U36235 (N_36235,N_33732,N_34030);
nand U36236 (N_36236,N_32828,N_32956);
or U36237 (N_36237,N_34960,N_33990);
and U36238 (N_36238,N_33329,N_34931);
xnor U36239 (N_36239,N_32730,N_34953);
or U36240 (N_36240,N_33316,N_34053);
and U36241 (N_36241,N_34706,N_33612);
nand U36242 (N_36242,N_34817,N_33098);
nand U36243 (N_36243,N_33110,N_34362);
nor U36244 (N_36244,N_34119,N_32530);
nor U36245 (N_36245,N_34638,N_33436);
and U36246 (N_36246,N_33660,N_32679);
or U36247 (N_36247,N_32928,N_33946);
nand U36248 (N_36248,N_33515,N_34933);
xnor U36249 (N_36249,N_33341,N_34352);
and U36250 (N_36250,N_33014,N_34086);
nand U36251 (N_36251,N_33836,N_34859);
or U36252 (N_36252,N_33823,N_34074);
nand U36253 (N_36253,N_34138,N_34149);
nand U36254 (N_36254,N_34275,N_32852);
xnor U36255 (N_36255,N_32911,N_34979);
and U36256 (N_36256,N_34203,N_32634);
xor U36257 (N_36257,N_34441,N_34763);
nand U36258 (N_36258,N_33424,N_33229);
and U36259 (N_36259,N_34852,N_32505);
nor U36260 (N_36260,N_33365,N_34369);
or U36261 (N_36261,N_33557,N_33760);
xnor U36262 (N_36262,N_32986,N_32746);
or U36263 (N_36263,N_32719,N_32681);
or U36264 (N_36264,N_34543,N_32547);
nor U36265 (N_36265,N_32971,N_34476);
xor U36266 (N_36266,N_33346,N_34165);
nor U36267 (N_36267,N_33225,N_34811);
xnor U36268 (N_36268,N_34377,N_34203);
nor U36269 (N_36269,N_33927,N_33038);
xor U36270 (N_36270,N_33781,N_34805);
xnor U36271 (N_36271,N_33341,N_32713);
and U36272 (N_36272,N_32585,N_33770);
nand U36273 (N_36273,N_33097,N_34189);
nand U36274 (N_36274,N_34861,N_33300);
nand U36275 (N_36275,N_34783,N_33452);
nor U36276 (N_36276,N_34837,N_33492);
xor U36277 (N_36277,N_34283,N_34974);
or U36278 (N_36278,N_33375,N_33250);
nor U36279 (N_36279,N_33791,N_33969);
and U36280 (N_36280,N_33339,N_34710);
or U36281 (N_36281,N_33926,N_32992);
nand U36282 (N_36282,N_34221,N_34606);
nor U36283 (N_36283,N_32916,N_33336);
or U36284 (N_36284,N_33499,N_34139);
and U36285 (N_36285,N_32993,N_32699);
nand U36286 (N_36286,N_34183,N_34570);
xnor U36287 (N_36287,N_34714,N_33603);
xnor U36288 (N_36288,N_33973,N_32804);
xor U36289 (N_36289,N_34599,N_33360);
xnor U36290 (N_36290,N_32894,N_33786);
nand U36291 (N_36291,N_33536,N_33724);
xor U36292 (N_36292,N_33940,N_33506);
xnor U36293 (N_36293,N_34351,N_33727);
and U36294 (N_36294,N_34363,N_34494);
nor U36295 (N_36295,N_34302,N_33462);
or U36296 (N_36296,N_33919,N_34463);
xor U36297 (N_36297,N_32950,N_33466);
nand U36298 (N_36298,N_32716,N_33221);
nor U36299 (N_36299,N_33172,N_32785);
nand U36300 (N_36300,N_33567,N_32988);
or U36301 (N_36301,N_32928,N_33975);
xnor U36302 (N_36302,N_34494,N_33409);
nor U36303 (N_36303,N_34884,N_33227);
xor U36304 (N_36304,N_34783,N_33659);
and U36305 (N_36305,N_33435,N_32859);
or U36306 (N_36306,N_34570,N_34992);
xor U36307 (N_36307,N_34682,N_33819);
xor U36308 (N_36308,N_32932,N_34656);
nand U36309 (N_36309,N_34511,N_33872);
nand U36310 (N_36310,N_33985,N_34131);
nor U36311 (N_36311,N_33365,N_34573);
nor U36312 (N_36312,N_33041,N_33086);
and U36313 (N_36313,N_34315,N_32547);
nor U36314 (N_36314,N_33194,N_33388);
nor U36315 (N_36315,N_33233,N_33343);
and U36316 (N_36316,N_33305,N_33619);
nor U36317 (N_36317,N_33323,N_32951);
xor U36318 (N_36318,N_33128,N_34121);
and U36319 (N_36319,N_33941,N_33392);
or U36320 (N_36320,N_34619,N_33298);
and U36321 (N_36321,N_32556,N_34342);
nor U36322 (N_36322,N_33292,N_34960);
or U36323 (N_36323,N_34357,N_34477);
or U36324 (N_36324,N_34097,N_34412);
nand U36325 (N_36325,N_34000,N_34421);
and U36326 (N_36326,N_34037,N_34609);
and U36327 (N_36327,N_34739,N_34378);
nand U36328 (N_36328,N_34606,N_32666);
xor U36329 (N_36329,N_33723,N_32925);
nand U36330 (N_36330,N_34690,N_34572);
xnor U36331 (N_36331,N_34797,N_32830);
xor U36332 (N_36332,N_34562,N_33416);
and U36333 (N_36333,N_32646,N_33120);
or U36334 (N_36334,N_34130,N_32567);
nor U36335 (N_36335,N_32609,N_33504);
xor U36336 (N_36336,N_32921,N_34347);
and U36337 (N_36337,N_34965,N_32733);
xnor U36338 (N_36338,N_33158,N_34015);
nor U36339 (N_36339,N_33722,N_32570);
nand U36340 (N_36340,N_33055,N_32756);
nor U36341 (N_36341,N_32578,N_34153);
or U36342 (N_36342,N_33299,N_32827);
nor U36343 (N_36343,N_34163,N_33622);
and U36344 (N_36344,N_34937,N_33573);
or U36345 (N_36345,N_34438,N_33951);
nand U36346 (N_36346,N_34477,N_32550);
nor U36347 (N_36347,N_32688,N_34663);
and U36348 (N_36348,N_34369,N_33863);
nor U36349 (N_36349,N_32824,N_33954);
and U36350 (N_36350,N_32679,N_32524);
xor U36351 (N_36351,N_34983,N_33086);
or U36352 (N_36352,N_34386,N_32847);
or U36353 (N_36353,N_32862,N_33257);
and U36354 (N_36354,N_33788,N_32791);
nor U36355 (N_36355,N_33386,N_32886);
or U36356 (N_36356,N_33795,N_33534);
nand U36357 (N_36357,N_33609,N_34902);
or U36358 (N_36358,N_34702,N_34437);
nor U36359 (N_36359,N_34378,N_34746);
nor U36360 (N_36360,N_34397,N_33075);
or U36361 (N_36361,N_34005,N_33127);
nand U36362 (N_36362,N_33373,N_33935);
or U36363 (N_36363,N_33987,N_33470);
or U36364 (N_36364,N_34952,N_33588);
nor U36365 (N_36365,N_33467,N_32873);
nand U36366 (N_36366,N_33526,N_34492);
or U36367 (N_36367,N_33486,N_33027);
or U36368 (N_36368,N_33019,N_32843);
nor U36369 (N_36369,N_32708,N_32739);
nand U36370 (N_36370,N_33650,N_34687);
nor U36371 (N_36371,N_34104,N_33606);
xor U36372 (N_36372,N_32519,N_34095);
xnor U36373 (N_36373,N_32704,N_32764);
or U36374 (N_36374,N_34518,N_34704);
nor U36375 (N_36375,N_34407,N_34883);
and U36376 (N_36376,N_34639,N_33130);
and U36377 (N_36377,N_33298,N_34008);
or U36378 (N_36378,N_33678,N_33442);
or U36379 (N_36379,N_34336,N_33786);
xor U36380 (N_36380,N_34959,N_33498);
or U36381 (N_36381,N_33107,N_34220);
xnor U36382 (N_36382,N_32664,N_32700);
or U36383 (N_36383,N_34974,N_32619);
nor U36384 (N_36384,N_33971,N_33261);
nand U36385 (N_36385,N_34751,N_33415);
and U36386 (N_36386,N_34467,N_34116);
xor U36387 (N_36387,N_34407,N_33621);
and U36388 (N_36388,N_34381,N_34658);
nor U36389 (N_36389,N_34964,N_34785);
nor U36390 (N_36390,N_34575,N_32593);
or U36391 (N_36391,N_34521,N_33619);
xor U36392 (N_36392,N_33943,N_33165);
xnor U36393 (N_36393,N_32820,N_34135);
nor U36394 (N_36394,N_33121,N_34722);
or U36395 (N_36395,N_32667,N_34239);
or U36396 (N_36396,N_34885,N_33845);
or U36397 (N_36397,N_33689,N_33177);
xnor U36398 (N_36398,N_34066,N_32830);
or U36399 (N_36399,N_33525,N_33985);
or U36400 (N_36400,N_34033,N_33953);
xnor U36401 (N_36401,N_33463,N_32524);
or U36402 (N_36402,N_32951,N_34054);
or U36403 (N_36403,N_32550,N_34168);
nand U36404 (N_36404,N_33387,N_33392);
and U36405 (N_36405,N_34862,N_34259);
and U36406 (N_36406,N_33311,N_34572);
xnor U36407 (N_36407,N_32852,N_33752);
and U36408 (N_36408,N_32773,N_32958);
nor U36409 (N_36409,N_33597,N_34758);
xnor U36410 (N_36410,N_32722,N_34539);
nand U36411 (N_36411,N_34817,N_33012);
nand U36412 (N_36412,N_34629,N_33879);
nand U36413 (N_36413,N_32782,N_33476);
nor U36414 (N_36414,N_33477,N_34809);
or U36415 (N_36415,N_34320,N_33573);
xnor U36416 (N_36416,N_33546,N_34045);
and U36417 (N_36417,N_33542,N_33147);
and U36418 (N_36418,N_33761,N_33203);
or U36419 (N_36419,N_33022,N_34332);
xor U36420 (N_36420,N_33958,N_32795);
and U36421 (N_36421,N_34396,N_33666);
nor U36422 (N_36422,N_33045,N_33951);
or U36423 (N_36423,N_33187,N_33306);
nor U36424 (N_36424,N_33116,N_34902);
and U36425 (N_36425,N_33766,N_33316);
and U36426 (N_36426,N_33640,N_32917);
nand U36427 (N_36427,N_34434,N_33141);
nor U36428 (N_36428,N_32884,N_32974);
nand U36429 (N_36429,N_34460,N_34023);
and U36430 (N_36430,N_34871,N_32808);
nor U36431 (N_36431,N_34581,N_34533);
and U36432 (N_36432,N_32891,N_33482);
and U36433 (N_36433,N_33238,N_32745);
and U36434 (N_36434,N_32985,N_34702);
or U36435 (N_36435,N_34355,N_33216);
nand U36436 (N_36436,N_34168,N_34394);
nand U36437 (N_36437,N_32728,N_34580);
nand U36438 (N_36438,N_33111,N_32701);
xnor U36439 (N_36439,N_34414,N_33786);
xor U36440 (N_36440,N_34841,N_33120);
or U36441 (N_36441,N_34391,N_33894);
xor U36442 (N_36442,N_33879,N_33622);
nand U36443 (N_36443,N_34719,N_34388);
nand U36444 (N_36444,N_34758,N_33775);
nor U36445 (N_36445,N_33863,N_33150);
and U36446 (N_36446,N_33551,N_34409);
nand U36447 (N_36447,N_33029,N_34211);
and U36448 (N_36448,N_34714,N_34769);
or U36449 (N_36449,N_33616,N_33818);
and U36450 (N_36450,N_33751,N_33794);
xor U36451 (N_36451,N_33443,N_33775);
nand U36452 (N_36452,N_33017,N_33866);
and U36453 (N_36453,N_34997,N_33112);
nor U36454 (N_36454,N_33332,N_33339);
and U36455 (N_36455,N_34309,N_33921);
nor U36456 (N_36456,N_32887,N_34025);
nor U36457 (N_36457,N_33022,N_34010);
nor U36458 (N_36458,N_34774,N_34082);
xor U36459 (N_36459,N_34719,N_33977);
xor U36460 (N_36460,N_33885,N_33543);
nand U36461 (N_36461,N_34211,N_34837);
xor U36462 (N_36462,N_33721,N_34849);
nand U36463 (N_36463,N_33653,N_34731);
nand U36464 (N_36464,N_33473,N_33464);
and U36465 (N_36465,N_32674,N_33416);
and U36466 (N_36466,N_34051,N_34383);
nand U36467 (N_36467,N_34900,N_34610);
nor U36468 (N_36468,N_34506,N_33677);
nand U36469 (N_36469,N_34338,N_34682);
nand U36470 (N_36470,N_33667,N_33337);
nor U36471 (N_36471,N_33860,N_33056);
nand U36472 (N_36472,N_33649,N_32941);
or U36473 (N_36473,N_33222,N_33821);
and U36474 (N_36474,N_34050,N_34932);
xnor U36475 (N_36475,N_34522,N_32944);
nor U36476 (N_36476,N_34749,N_33821);
nand U36477 (N_36477,N_32819,N_34371);
nor U36478 (N_36478,N_32897,N_32692);
or U36479 (N_36479,N_33385,N_32753);
xnor U36480 (N_36480,N_34558,N_34894);
and U36481 (N_36481,N_33307,N_34923);
nor U36482 (N_36482,N_33756,N_34300);
and U36483 (N_36483,N_34658,N_33336);
and U36484 (N_36484,N_34749,N_32714);
nand U36485 (N_36485,N_33116,N_33216);
xnor U36486 (N_36486,N_34956,N_33915);
xor U36487 (N_36487,N_32928,N_33305);
nor U36488 (N_36488,N_32501,N_34810);
and U36489 (N_36489,N_33019,N_33250);
nor U36490 (N_36490,N_32982,N_34820);
nor U36491 (N_36491,N_33520,N_32736);
and U36492 (N_36492,N_33688,N_34422);
nor U36493 (N_36493,N_32927,N_34000);
xor U36494 (N_36494,N_33552,N_34440);
and U36495 (N_36495,N_33601,N_34453);
and U36496 (N_36496,N_33571,N_33325);
nor U36497 (N_36497,N_33610,N_32863);
nand U36498 (N_36498,N_34542,N_34223);
xor U36499 (N_36499,N_34256,N_32764);
nor U36500 (N_36500,N_34348,N_32552);
nand U36501 (N_36501,N_32507,N_34378);
xor U36502 (N_36502,N_33854,N_33791);
nand U36503 (N_36503,N_34355,N_33718);
xor U36504 (N_36504,N_33163,N_33001);
xor U36505 (N_36505,N_33871,N_32794);
or U36506 (N_36506,N_33112,N_33995);
nand U36507 (N_36507,N_33967,N_32923);
nand U36508 (N_36508,N_32560,N_32708);
nor U36509 (N_36509,N_33145,N_32667);
nor U36510 (N_36510,N_34232,N_32639);
nor U36511 (N_36511,N_32855,N_34311);
nor U36512 (N_36512,N_34090,N_34624);
nand U36513 (N_36513,N_34812,N_33446);
xnor U36514 (N_36514,N_34513,N_32642);
or U36515 (N_36515,N_34543,N_34614);
xnor U36516 (N_36516,N_33620,N_34678);
nand U36517 (N_36517,N_34708,N_34212);
nor U36518 (N_36518,N_34839,N_34870);
and U36519 (N_36519,N_34115,N_33593);
nand U36520 (N_36520,N_32549,N_32756);
nand U36521 (N_36521,N_34958,N_33761);
or U36522 (N_36522,N_33112,N_34103);
nand U36523 (N_36523,N_33532,N_34994);
and U36524 (N_36524,N_33558,N_32822);
or U36525 (N_36525,N_32623,N_33170);
nand U36526 (N_36526,N_33581,N_33474);
nand U36527 (N_36527,N_34417,N_33841);
and U36528 (N_36528,N_32739,N_34066);
nand U36529 (N_36529,N_32663,N_34744);
and U36530 (N_36530,N_34026,N_34397);
nor U36531 (N_36531,N_34121,N_32750);
nand U36532 (N_36532,N_33889,N_34953);
and U36533 (N_36533,N_34420,N_34693);
or U36534 (N_36534,N_33653,N_32885);
xor U36535 (N_36535,N_34382,N_33370);
nand U36536 (N_36536,N_34595,N_34308);
or U36537 (N_36537,N_33224,N_34691);
xor U36538 (N_36538,N_34645,N_33102);
xnor U36539 (N_36539,N_34445,N_34102);
nor U36540 (N_36540,N_34945,N_34232);
nand U36541 (N_36541,N_33929,N_33742);
nor U36542 (N_36542,N_34124,N_34770);
nand U36543 (N_36543,N_34332,N_34627);
nand U36544 (N_36544,N_34817,N_32632);
xnor U36545 (N_36545,N_34063,N_34320);
nor U36546 (N_36546,N_34419,N_34661);
xor U36547 (N_36547,N_33669,N_34575);
xor U36548 (N_36548,N_34151,N_33704);
xor U36549 (N_36549,N_33600,N_33196);
nor U36550 (N_36550,N_32549,N_32527);
nor U36551 (N_36551,N_33672,N_34400);
or U36552 (N_36552,N_33491,N_33786);
nor U36553 (N_36553,N_33589,N_33335);
or U36554 (N_36554,N_34384,N_33428);
xnor U36555 (N_36555,N_32587,N_34072);
nor U36556 (N_36556,N_34841,N_32887);
and U36557 (N_36557,N_34468,N_33604);
nand U36558 (N_36558,N_34281,N_33869);
xor U36559 (N_36559,N_33490,N_32637);
nor U36560 (N_36560,N_33404,N_33588);
or U36561 (N_36561,N_32906,N_33475);
nor U36562 (N_36562,N_34397,N_34987);
and U36563 (N_36563,N_34550,N_32874);
or U36564 (N_36564,N_33888,N_32616);
and U36565 (N_36565,N_34288,N_34545);
nand U36566 (N_36566,N_32587,N_33409);
xnor U36567 (N_36567,N_33364,N_33700);
nor U36568 (N_36568,N_33983,N_34744);
or U36569 (N_36569,N_34003,N_33729);
xor U36570 (N_36570,N_34712,N_33766);
xor U36571 (N_36571,N_32516,N_32668);
and U36572 (N_36572,N_34984,N_32527);
nand U36573 (N_36573,N_34554,N_34935);
and U36574 (N_36574,N_33941,N_33445);
xor U36575 (N_36575,N_34973,N_32569);
nor U36576 (N_36576,N_32538,N_33255);
nor U36577 (N_36577,N_34452,N_34467);
or U36578 (N_36578,N_33282,N_33042);
and U36579 (N_36579,N_33186,N_34438);
or U36580 (N_36580,N_32962,N_34390);
nand U36581 (N_36581,N_33299,N_33270);
xnor U36582 (N_36582,N_33030,N_33124);
xor U36583 (N_36583,N_32511,N_34787);
nand U36584 (N_36584,N_33394,N_33583);
nor U36585 (N_36585,N_33789,N_34627);
or U36586 (N_36586,N_34531,N_33305);
and U36587 (N_36587,N_34193,N_33239);
and U36588 (N_36588,N_34823,N_33885);
and U36589 (N_36589,N_34994,N_34718);
nand U36590 (N_36590,N_33182,N_33789);
xnor U36591 (N_36591,N_34677,N_32777);
xor U36592 (N_36592,N_33321,N_34133);
xnor U36593 (N_36593,N_33655,N_34195);
nor U36594 (N_36594,N_32876,N_33116);
nor U36595 (N_36595,N_33134,N_33979);
or U36596 (N_36596,N_33808,N_32899);
and U36597 (N_36597,N_34599,N_32568);
and U36598 (N_36598,N_33899,N_34748);
and U36599 (N_36599,N_33154,N_32657);
nand U36600 (N_36600,N_32982,N_34715);
xnor U36601 (N_36601,N_33789,N_32751);
and U36602 (N_36602,N_33394,N_34486);
xor U36603 (N_36603,N_34845,N_32682);
nor U36604 (N_36604,N_34166,N_32718);
nand U36605 (N_36605,N_32723,N_32533);
and U36606 (N_36606,N_32845,N_32855);
nand U36607 (N_36607,N_33415,N_32980);
nand U36608 (N_36608,N_33046,N_34577);
and U36609 (N_36609,N_34000,N_34747);
nor U36610 (N_36610,N_34514,N_34748);
nand U36611 (N_36611,N_33065,N_33710);
xnor U36612 (N_36612,N_33529,N_34872);
xor U36613 (N_36613,N_34972,N_33515);
or U36614 (N_36614,N_34002,N_33932);
nor U36615 (N_36615,N_34967,N_34734);
or U36616 (N_36616,N_34297,N_32916);
nand U36617 (N_36617,N_34911,N_33428);
nor U36618 (N_36618,N_34651,N_34737);
or U36619 (N_36619,N_33557,N_34156);
xor U36620 (N_36620,N_32621,N_33091);
and U36621 (N_36621,N_33574,N_34300);
or U36622 (N_36622,N_32858,N_33757);
xor U36623 (N_36623,N_34225,N_34435);
and U36624 (N_36624,N_34650,N_33529);
and U36625 (N_36625,N_32898,N_33466);
xnor U36626 (N_36626,N_33338,N_34795);
xor U36627 (N_36627,N_32900,N_34430);
and U36628 (N_36628,N_34277,N_33399);
nand U36629 (N_36629,N_33409,N_32804);
or U36630 (N_36630,N_33870,N_32902);
and U36631 (N_36631,N_32970,N_32878);
or U36632 (N_36632,N_33432,N_32772);
and U36633 (N_36633,N_33077,N_32678);
nand U36634 (N_36634,N_34263,N_32733);
xnor U36635 (N_36635,N_33887,N_32578);
nor U36636 (N_36636,N_33355,N_34000);
nand U36637 (N_36637,N_33415,N_33855);
xnor U36638 (N_36638,N_34121,N_33906);
nor U36639 (N_36639,N_33114,N_34581);
or U36640 (N_36640,N_33548,N_32970);
or U36641 (N_36641,N_32645,N_34803);
or U36642 (N_36642,N_32960,N_33812);
xnor U36643 (N_36643,N_34958,N_34518);
or U36644 (N_36644,N_33380,N_34543);
nor U36645 (N_36645,N_34446,N_34389);
nand U36646 (N_36646,N_33275,N_33730);
or U36647 (N_36647,N_34249,N_33668);
or U36648 (N_36648,N_33010,N_34323);
nand U36649 (N_36649,N_33122,N_33529);
xnor U36650 (N_36650,N_34381,N_33068);
and U36651 (N_36651,N_32735,N_34852);
or U36652 (N_36652,N_34406,N_33449);
nor U36653 (N_36653,N_32778,N_34488);
nor U36654 (N_36654,N_34075,N_32812);
nor U36655 (N_36655,N_34866,N_33791);
xor U36656 (N_36656,N_33526,N_34469);
nor U36657 (N_36657,N_33831,N_32842);
nand U36658 (N_36658,N_34402,N_33937);
nand U36659 (N_36659,N_33134,N_32559);
nor U36660 (N_36660,N_33791,N_34893);
or U36661 (N_36661,N_34091,N_34456);
xnor U36662 (N_36662,N_34489,N_32996);
and U36663 (N_36663,N_33709,N_34667);
and U36664 (N_36664,N_34712,N_34272);
nor U36665 (N_36665,N_33122,N_32702);
and U36666 (N_36666,N_33739,N_34537);
nor U36667 (N_36667,N_32880,N_33155);
or U36668 (N_36668,N_33657,N_32793);
nand U36669 (N_36669,N_32609,N_34678);
xor U36670 (N_36670,N_32963,N_32856);
nand U36671 (N_36671,N_33166,N_33183);
or U36672 (N_36672,N_34881,N_34478);
xor U36673 (N_36673,N_33812,N_34522);
or U36674 (N_36674,N_32812,N_34247);
and U36675 (N_36675,N_33018,N_34058);
and U36676 (N_36676,N_33059,N_34110);
xnor U36677 (N_36677,N_34313,N_34217);
and U36678 (N_36678,N_34968,N_32929);
nor U36679 (N_36679,N_34312,N_34159);
nor U36680 (N_36680,N_34051,N_32633);
xor U36681 (N_36681,N_33761,N_33499);
nor U36682 (N_36682,N_33472,N_32584);
or U36683 (N_36683,N_34432,N_32569);
nand U36684 (N_36684,N_32666,N_34219);
xnor U36685 (N_36685,N_32990,N_33074);
nor U36686 (N_36686,N_33741,N_34303);
or U36687 (N_36687,N_34535,N_33633);
xor U36688 (N_36688,N_34485,N_34672);
and U36689 (N_36689,N_33247,N_34521);
or U36690 (N_36690,N_33486,N_33651);
or U36691 (N_36691,N_32870,N_34071);
and U36692 (N_36692,N_33784,N_34703);
nor U36693 (N_36693,N_32721,N_34560);
nor U36694 (N_36694,N_32664,N_33692);
nand U36695 (N_36695,N_32726,N_33612);
and U36696 (N_36696,N_33618,N_32838);
and U36697 (N_36697,N_34692,N_34040);
xnor U36698 (N_36698,N_34352,N_33822);
or U36699 (N_36699,N_34562,N_32565);
and U36700 (N_36700,N_34161,N_34089);
nor U36701 (N_36701,N_33805,N_34563);
xor U36702 (N_36702,N_32531,N_32683);
and U36703 (N_36703,N_34564,N_33981);
nand U36704 (N_36704,N_32512,N_32577);
and U36705 (N_36705,N_33704,N_33332);
nand U36706 (N_36706,N_34995,N_34931);
nor U36707 (N_36707,N_32930,N_34088);
xnor U36708 (N_36708,N_32776,N_34075);
nand U36709 (N_36709,N_32713,N_33066);
and U36710 (N_36710,N_32986,N_33836);
and U36711 (N_36711,N_32618,N_33623);
or U36712 (N_36712,N_34966,N_33185);
and U36713 (N_36713,N_33666,N_34081);
xnor U36714 (N_36714,N_34971,N_33982);
nand U36715 (N_36715,N_33864,N_34468);
xor U36716 (N_36716,N_34915,N_33020);
or U36717 (N_36717,N_33894,N_33767);
xor U36718 (N_36718,N_32848,N_32892);
or U36719 (N_36719,N_34470,N_34933);
xnor U36720 (N_36720,N_33575,N_34402);
or U36721 (N_36721,N_33346,N_34573);
nor U36722 (N_36722,N_33837,N_32629);
and U36723 (N_36723,N_34691,N_33544);
or U36724 (N_36724,N_34039,N_34092);
xnor U36725 (N_36725,N_33454,N_34415);
and U36726 (N_36726,N_33616,N_33742);
xor U36727 (N_36727,N_32914,N_34961);
nand U36728 (N_36728,N_34689,N_34204);
nor U36729 (N_36729,N_34417,N_33981);
xnor U36730 (N_36730,N_32564,N_32751);
xnor U36731 (N_36731,N_33623,N_33636);
or U36732 (N_36732,N_32570,N_33163);
and U36733 (N_36733,N_34778,N_33027);
xnor U36734 (N_36734,N_32817,N_34654);
nor U36735 (N_36735,N_34047,N_32718);
or U36736 (N_36736,N_33940,N_32549);
or U36737 (N_36737,N_33478,N_34203);
or U36738 (N_36738,N_33191,N_34315);
xor U36739 (N_36739,N_34759,N_32586);
or U36740 (N_36740,N_34365,N_32774);
nand U36741 (N_36741,N_33406,N_33283);
or U36742 (N_36742,N_34106,N_33013);
xor U36743 (N_36743,N_33715,N_34121);
and U36744 (N_36744,N_33062,N_32664);
xor U36745 (N_36745,N_34137,N_34343);
or U36746 (N_36746,N_34667,N_33865);
xor U36747 (N_36747,N_32694,N_34238);
nor U36748 (N_36748,N_33571,N_33423);
or U36749 (N_36749,N_34298,N_33656);
and U36750 (N_36750,N_34705,N_33258);
nor U36751 (N_36751,N_33242,N_33957);
and U36752 (N_36752,N_34312,N_33099);
xnor U36753 (N_36753,N_33041,N_34622);
xnor U36754 (N_36754,N_33357,N_32818);
nor U36755 (N_36755,N_33014,N_33433);
xor U36756 (N_36756,N_33086,N_33815);
nand U36757 (N_36757,N_33507,N_34162);
or U36758 (N_36758,N_33056,N_34723);
nand U36759 (N_36759,N_34736,N_34087);
nand U36760 (N_36760,N_33875,N_34364);
or U36761 (N_36761,N_33360,N_33912);
nor U36762 (N_36762,N_34803,N_34852);
or U36763 (N_36763,N_33805,N_32816);
and U36764 (N_36764,N_33451,N_34733);
nand U36765 (N_36765,N_33780,N_32802);
or U36766 (N_36766,N_33687,N_33393);
or U36767 (N_36767,N_33025,N_34782);
nor U36768 (N_36768,N_32524,N_34732);
nor U36769 (N_36769,N_34728,N_33617);
nor U36770 (N_36770,N_34708,N_32801);
nor U36771 (N_36771,N_34525,N_33217);
and U36772 (N_36772,N_34058,N_34071);
nor U36773 (N_36773,N_34824,N_34784);
nand U36774 (N_36774,N_32877,N_33375);
xnor U36775 (N_36775,N_33891,N_32650);
xnor U36776 (N_36776,N_34778,N_33897);
nor U36777 (N_36777,N_33691,N_32760);
or U36778 (N_36778,N_34833,N_33842);
nand U36779 (N_36779,N_33248,N_34905);
nor U36780 (N_36780,N_32870,N_32653);
nand U36781 (N_36781,N_33919,N_34865);
nand U36782 (N_36782,N_33850,N_33256);
xor U36783 (N_36783,N_34454,N_32556);
and U36784 (N_36784,N_32639,N_34499);
nor U36785 (N_36785,N_32936,N_33303);
and U36786 (N_36786,N_33394,N_34623);
and U36787 (N_36787,N_33540,N_32811);
and U36788 (N_36788,N_34648,N_33879);
and U36789 (N_36789,N_34254,N_34720);
xnor U36790 (N_36790,N_32696,N_33494);
or U36791 (N_36791,N_34486,N_33018);
nor U36792 (N_36792,N_32672,N_34100);
and U36793 (N_36793,N_34252,N_34006);
or U36794 (N_36794,N_34696,N_33924);
and U36795 (N_36795,N_34020,N_33327);
and U36796 (N_36796,N_32961,N_34674);
nand U36797 (N_36797,N_33455,N_32639);
nor U36798 (N_36798,N_34834,N_33049);
or U36799 (N_36799,N_32724,N_33585);
and U36800 (N_36800,N_33014,N_32894);
nand U36801 (N_36801,N_33539,N_33593);
xnor U36802 (N_36802,N_34693,N_34924);
and U36803 (N_36803,N_34272,N_33375);
or U36804 (N_36804,N_34566,N_33574);
and U36805 (N_36805,N_34968,N_33923);
and U36806 (N_36806,N_34045,N_34923);
and U36807 (N_36807,N_33023,N_33031);
or U36808 (N_36808,N_33086,N_33703);
and U36809 (N_36809,N_32502,N_34533);
or U36810 (N_36810,N_33497,N_32774);
and U36811 (N_36811,N_34965,N_33782);
nor U36812 (N_36812,N_34078,N_32755);
nand U36813 (N_36813,N_34152,N_32595);
and U36814 (N_36814,N_34574,N_33548);
nor U36815 (N_36815,N_33599,N_33283);
xnor U36816 (N_36816,N_34318,N_34064);
xor U36817 (N_36817,N_34950,N_33446);
and U36818 (N_36818,N_33618,N_33462);
nand U36819 (N_36819,N_33160,N_34130);
or U36820 (N_36820,N_33298,N_34343);
nand U36821 (N_36821,N_33816,N_34344);
nor U36822 (N_36822,N_34864,N_33282);
nor U36823 (N_36823,N_34203,N_32932);
nand U36824 (N_36824,N_33811,N_32548);
nand U36825 (N_36825,N_33249,N_33798);
or U36826 (N_36826,N_34748,N_34361);
nor U36827 (N_36827,N_34533,N_34945);
nor U36828 (N_36828,N_34925,N_32514);
nand U36829 (N_36829,N_34541,N_33041);
xnor U36830 (N_36830,N_34973,N_34161);
xor U36831 (N_36831,N_33394,N_32703);
nand U36832 (N_36832,N_33420,N_33367);
nor U36833 (N_36833,N_34778,N_33682);
xor U36834 (N_36834,N_34237,N_34936);
nor U36835 (N_36835,N_33203,N_34107);
nor U36836 (N_36836,N_32741,N_34856);
nor U36837 (N_36837,N_34745,N_33503);
nor U36838 (N_36838,N_34501,N_34525);
xor U36839 (N_36839,N_34811,N_33909);
nand U36840 (N_36840,N_33070,N_34475);
nor U36841 (N_36841,N_33255,N_34796);
and U36842 (N_36842,N_32824,N_32799);
xor U36843 (N_36843,N_33876,N_33683);
or U36844 (N_36844,N_33257,N_34711);
nor U36845 (N_36845,N_32583,N_33036);
nand U36846 (N_36846,N_33663,N_32966);
or U36847 (N_36847,N_33857,N_34323);
nor U36848 (N_36848,N_33672,N_34482);
nor U36849 (N_36849,N_33459,N_34672);
and U36850 (N_36850,N_33244,N_33842);
nand U36851 (N_36851,N_32982,N_34893);
nor U36852 (N_36852,N_34304,N_34266);
nand U36853 (N_36853,N_33686,N_34105);
nor U36854 (N_36854,N_33910,N_33650);
or U36855 (N_36855,N_33229,N_32983);
xor U36856 (N_36856,N_32971,N_32850);
or U36857 (N_36857,N_34948,N_34974);
xor U36858 (N_36858,N_32938,N_33135);
and U36859 (N_36859,N_33451,N_33642);
and U36860 (N_36860,N_34380,N_33259);
and U36861 (N_36861,N_34405,N_33293);
or U36862 (N_36862,N_34939,N_32660);
xor U36863 (N_36863,N_33110,N_34413);
and U36864 (N_36864,N_34027,N_34934);
nor U36865 (N_36865,N_32768,N_32569);
xnor U36866 (N_36866,N_34806,N_33134);
xnor U36867 (N_36867,N_32784,N_34098);
or U36868 (N_36868,N_34935,N_34042);
or U36869 (N_36869,N_34078,N_33192);
and U36870 (N_36870,N_34009,N_34395);
nor U36871 (N_36871,N_32959,N_32642);
xnor U36872 (N_36872,N_32736,N_34759);
or U36873 (N_36873,N_33198,N_32502);
or U36874 (N_36874,N_32554,N_34661);
nor U36875 (N_36875,N_32528,N_32730);
nand U36876 (N_36876,N_33863,N_32540);
nand U36877 (N_36877,N_34334,N_33586);
xnor U36878 (N_36878,N_33470,N_34246);
and U36879 (N_36879,N_33222,N_34721);
nand U36880 (N_36880,N_34224,N_33449);
nor U36881 (N_36881,N_34942,N_32981);
xor U36882 (N_36882,N_32766,N_34959);
nor U36883 (N_36883,N_33235,N_33403);
xnor U36884 (N_36884,N_33266,N_34008);
and U36885 (N_36885,N_34480,N_32831);
and U36886 (N_36886,N_33866,N_34630);
nor U36887 (N_36887,N_33136,N_34270);
nand U36888 (N_36888,N_33344,N_33754);
and U36889 (N_36889,N_33565,N_34302);
xnor U36890 (N_36890,N_34072,N_33298);
or U36891 (N_36891,N_33510,N_33650);
nand U36892 (N_36892,N_34339,N_34905);
xnor U36893 (N_36893,N_33306,N_34521);
nand U36894 (N_36894,N_33261,N_34665);
nand U36895 (N_36895,N_34532,N_34233);
xnor U36896 (N_36896,N_34344,N_32635);
xnor U36897 (N_36897,N_34119,N_33315);
or U36898 (N_36898,N_34494,N_33674);
and U36899 (N_36899,N_34175,N_34108);
nand U36900 (N_36900,N_33148,N_33011);
nand U36901 (N_36901,N_32579,N_34902);
and U36902 (N_36902,N_32621,N_33244);
or U36903 (N_36903,N_33189,N_33916);
and U36904 (N_36904,N_32620,N_32966);
xnor U36905 (N_36905,N_32913,N_34948);
xnor U36906 (N_36906,N_33137,N_33407);
nand U36907 (N_36907,N_34668,N_32824);
or U36908 (N_36908,N_33522,N_34868);
xor U36909 (N_36909,N_33442,N_32757);
and U36910 (N_36910,N_34717,N_34356);
xor U36911 (N_36911,N_34174,N_34938);
nand U36912 (N_36912,N_32644,N_34756);
xor U36913 (N_36913,N_33012,N_33062);
xnor U36914 (N_36914,N_34775,N_33578);
xnor U36915 (N_36915,N_34090,N_34720);
nand U36916 (N_36916,N_32769,N_34559);
xnor U36917 (N_36917,N_32888,N_34022);
xor U36918 (N_36918,N_34594,N_34524);
or U36919 (N_36919,N_33474,N_34652);
and U36920 (N_36920,N_34567,N_34494);
and U36921 (N_36921,N_34045,N_33338);
nand U36922 (N_36922,N_33921,N_33679);
xnor U36923 (N_36923,N_33716,N_33931);
nor U36924 (N_36924,N_34031,N_34791);
nor U36925 (N_36925,N_32519,N_33278);
or U36926 (N_36926,N_34107,N_33744);
nand U36927 (N_36927,N_33000,N_33210);
nor U36928 (N_36928,N_34106,N_34054);
nor U36929 (N_36929,N_34609,N_33008);
nand U36930 (N_36930,N_33579,N_33325);
and U36931 (N_36931,N_34457,N_33468);
or U36932 (N_36932,N_34696,N_33174);
xnor U36933 (N_36933,N_33690,N_32998);
and U36934 (N_36934,N_32557,N_33965);
or U36935 (N_36935,N_34817,N_32798);
and U36936 (N_36936,N_34181,N_34186);
and U36937 (N_36937,N_32942,N_34510);
nand U36938 (N_36938,N_33420,N_33086);
nand U36939 (N_36939,N_34216,N_33573);
xor U36940 (N_36940,N_33738,N_34821);
and U36941 (N_36941,N_33806,N_34342);
nand U36942 (N_36942,N_33304,N_34553);
xor U36943 (N_36943,N_33397,N_34521);
nor U36944 (N_36944,N_32695,N_34790);
xnor U36945 (N_36945,N_33036,N_33245);
or U36946 (N_36946,N_34484,N_33016);
or U36947 (N_36947,N_32597,N_33062);
and U36948 (N_36948,N_32574,N_34756);
and U36949 (N_36949,N_34890,N_34584);
xnor U36950 (N_36950,N_34998,N_32814);
or U36951 (N_36951,N_34967,N_34324);
and U36952 (N_36952,N_33477,N_34478);
or U36953 (N_36953,N_33365,N_34125);
nor U36954 (N_36954,N_34335,N_34137);
nand U36955 (N_36955,N_34291,N_33740);
and U36956 (N_36956,N_32894,N_33231);
nor U36957 (N_36957,N_34897,N_32948);
and U36958 (N_36958,N_32788,N_34977);
and U36959 (N_36959,N_34696,N_34029);
or U36960 (N_36960,N_34327,N_34825);
and U36961 (N_36961,N_32990,N_34875);
or U36962 (N_36962,N_32699,N_34642);
and U36963 (N_36963,N_34624,N_32661);
xor U36964 (N_36964,N_32951,N_34629);
or U36965 (N_36965,N_32809,N_34568);
and U36966 (N_36966,N_34006,N_34105);
nand U36967 (N_36967,N_33967,N_34805);
xor U36968 (N_36968,N_32622,N_34562);
xnor U36969 (N_36969,N_34987,N_32537);
and U36970 (N_36970,N_33838,N_33683);
or U36971 (N_36971,N_34268,N_33188);
xor U36972 (N_36972,N_34614,N_34991);
nor U36973 (N_36973,N_34146,N_33293);
nor U36974 (N_36974,N_32558,N_33557);
or U36975 (N_36975,N_33434,N_33202);
nand U36976 (N_36976,N_34440,N_33977);
and U36977 (N_36977,N_34630,N_33533);
nand U36978 (N_36978,N_33849,N_33991);
nor U36979 (N_36979,N_33767,N_33180);
nor U36980 (N_36980,N_34745,N_32976);
and U36981 (N_36981,N_34971,N_33844);
nand U36982 (N_36982,N_33448,N_33158);
and U36983 (N_36983,N_34362,N_33077);
nor U36984 (N_36984,N_33573,N_32784);
xor U36985 (N_36985,N_34766,N_34178);
xnor U36986 (N_36986,N_34424,N_33766);
and U36987 (N_36987,N_33241,N_33283);
or U36988 (N_36988,N_34587,N_33059);
xor U36989 (N_36989,N_33451,N_33317);
xnor U36990 (N_36990,N_33389,N_34514);
and U36991 (N_36991,N_34362,N_32916);
nand U36992 (N_36992,N_33147,N_33151);
and U36993 (N_36993,N_32699,N_34786);
or U36994 (N_36994,N_33676,N_32976);
xnor U36995 (N_36995,N_34328,N_33657);
and U36996 (N_36996,N_34433,N_34311);
xor U36997 (N_36997,N_33495,N_34213);
nand U36998 (N_36998,N_33423,N_34391);
xnor U36999 (N_36999,N_33517,N_32688);
and U37000 (N_37000,N_34382,N_34034);
nor U37001 (N_37001,N_33345,N_34888);
and U37002 (N_37002,N_34386,N_33715);
and U37003 (N_37003,N_32998,N_34321);
nand U37004 (N_37004,N_33233,N_33602);
and U37005 (N_37005,N_34746,N_34449);
or U37006 (N_37006,N_33139,N_33448);
nand U37007 (N_37007,N_33370,N_32781);
or U37008 (N_37008,N_33760,N_32985);
nor U37009 (N_37009,N_32772,N_32731);
nor U37010 (N_37010,N_32964,N_34162);
and U37011 (N_37011,N_34714,N_33820);
and U37012 (N_37012,N_34012,N_32530);
and U37013 (N_37013,N_33497,N_34563);
xor U37014 (N_37014,N_34870,N_33104);
or U37015 (N_37015,N_33651,N_33529);
nor U37016 (N_37016,N_32653,N_34427);
nor U37017 (N_37017,N_34768,N_34594);
xor U37018 (N_37018,N_33677,N_34573);
and U37019 (N_37019,N_33867,N_33527);
or U37020 (N_37020,N_32758,N_34150);
nand U37021 (N_37021,N_34406,N_32602);
nor U37022 (N_37022,N_33273,N_32937);
nor U37023 (N_37023,N_33662,N_34878);
nor U37024 (N_37024,N_34855,N_33147);
xnor U37025 (N_37025,N_34673,N_32712);
xor U37026 (N_37026,N_33856,N_33737);
nand U37027 (N_37027,N_34982,N_34361);
xor U37028 (N_37028,N_32676,N_34245);
nor U37029 (N_37029,N_32789,N_33940);
nand U37030 (N_37030,N_32526,N_33476);
xnor U37031 (N_37031,N_34771,N_33589);
or U37032 (N_37032,N_33765,N_32834);
nor U37033 (N_37033,N_34084,N_33189);
nand U37034 (N_37034,N_34731,N_33093);
nor U37035 (N_37035,N_33354,N_34808);
or U37036 (N_37036,N_34259,N_32635);
or U37037 (N_37037,N_34141,N_33188);
or U37038 (N_37038,N_33201,N_33229);
and U37039 (N_37039,N_34022,N_33966);
nor U37040 (N_37040,N_32953,N_33449);
nor U37041 (N_37041,N_33080,N_34104);
and U37042 (N_37042,N_33772,N_32899);
nand U37043 (N_37043,N_34726,N_34856);
or U37044 (N_37044,N_34978,N_32854);
nor U37045 (N_37045,N_34783,N_33865);
or U37046 (N_37046,N_33913,N_33746);
nor U37047 (N_37047,N_33474,N_34972);
and U37048 (N_37048,N_33466,N_34910);
and U37049 (N_37049,N_34634,N_34651);
and U37050 (N_37050,N_33458,N_33818);
or U37051 (N_37051,N_33236,N_34399);
or U37052 (N_37052,N_34626,N_34725);
nand U37053 (N_37053,N_33448,N_34226);
nor U37054 (N_37054,N_32862,N_32516);
nand U37055 (N_37055,N_34683,N_33314);
or U37056 (N_37056,N_34651,N_33940);
nor U37057 (N_37057,N_34687,N_34848);
nor U37058 (N_37058,N_33225,N_32905);
xnor U37059 (N_37059,N_33121,N_34444);
or U37060 (N_37060,N_33722,N_34789);
nor U37061 (N_37061,N_33173,N_33480);
and U37062 (N_37062,N_33920,N_34228);
and U37063 (N_37063,N_34784,N_33001);
xor U37064 (N_37064,N_33830,N_32931);
and U37065 (N_37065,N_34944,N_32540);
nand U37066 (N_37066,N_34692,N_33962);
xnor U37067 (N_37067,N_34214,N_34786);
xor U37068 (N_37068,N_33790,N_33136);
nand U37069 (N_37069,N_34266,N_32681);
nor U37070 (N_37070,N_34915,N_33893);
xor U37071 (N_37071,N_34794,N_34106);
xor U37072 (N_37072,N_34599,N_34087);
nor U37073 (N_37073,N_33876,N_32879);
xnor U37074 (N_37074,N_34062,N_34838);
nor U37075 (N_37075,N_32789,N_32768);
or U37076 (N_37076,N_32645,N_32911);
nor U37077 (N_37077,N_34610,N_34865);
and U37078 (N_37078,N_34735,N_33211);
and U37079 (N_37079,N_33786,N_33132);
and U37080 (N_37080,N_33620,N_33972);
xnor U37081 (N_37081,N_33442,N_32775);
nand U37082 (N_37082,N_33353,N_34836);
nor U37083 (N_37083,N_34666,N_32706);
nor U37084 (N_37084,N_32539,N_34966);
xnor U37085 (N_37085,N_32607,N_34291);
nand U37086 (N_37086,N_33414,N_34137);
nand U37087 (N_37087,N_34951,N_33766);
nand U37088 (N_37088,N_34538,N_34194);
nor U37089 (N_37089,N_33119,N_33351);
xor U37090 (N_37090,N_34198,N_32697);
nor U37091 (N_37091,N_34821,N_33156);
nor U37092 (N_37092,N_33205,N_33241);
and U37093 (N_37093,N_33532,N_34374);
nand U37094 (N_37094,N_33806,N_34703);
xor U37095 (N_37095,N_34203,N_32945);
nor U37096 (N_37096,N_33202,N_33717);
nor U37097 (N_37097,N_34985,N_34415);
nor U37098 (N_37098,N_33070,N_33815);
nor U37099 (N_37099,N_34334,N_33260);
or U37100 (N_37100,N_32645,N_34137);
xor U37101 (N_37101,N_33536,N_34160);
and U37102 (N_37102,N_32739,N_33402);
and U37103 (N_37103,N_34240,N_34349);
nor U37104 (N_37104,N_34148,N_33985);
nor U37105 (N_37105,N_33443,N_34848);
and U37106 (N_37106,N_34733,N_34113);
and U37107 (N_37107,N_33602,N_34506);
or U37108 (N_37108,N_34286,N_34216);
nor U37109 (N_37109,N_33871,N_32999);
or U37110 (N_37110,N_32755,N_34115);
and U37111 (N_37111,N_33087,N_32778);
nor U37112 (N_37112,N_34519,N_33440);
and U37113 (N_37113,N_34448,N_34818);
or U37114 (N_37114,N_32708,N_32582);
or U37115 (N_37115,N_33809,N_32712);
nand U37116 (N_37116,N_32841,N_33894);
nand U37117 (N_37117,N_33425,N_34048);
nand U37118 (N_37118,N_33180,N_32711);
and U37119 (N_37119,N_34402,N_32760);
xor U37120 (N_37120,N_34277,N_34240);
or U37121 (N_37121,N_32533,N_33982);
and U37122 (N_37122,N_34059,N_32821);
nor U37123 (N_37123,N_33287,N_32642);
and U37124 (N_37124,N_33248,N_34900);
xnor U37125 (N_37125,N_34019,N_34682);
nand U37126 (N_37126,N_34232,N_34250);
and U37127 (N_37127,N_34139,N_33870);
xor U37128 (N_37128,N_33745,N_33093);
nand U37129 (N_37129,N_33675,N_33354);
nor U37130 (N_37130,N_32836,N_32612);
and U37131 (N_37131,N_33306,N_32618);
nor U37132 (N_37132,N_32597,N_32565);
xor U37133 (N_37133,N_34698,N_33433);
nor U37134 (N_37134,N_32955,N_33949);
or U37135 (N_37135,N_34459,N_34468);
or U37136 (N_37136,N_32994,N_34345);
nand U37137 (N_37137,N_33613,N_33304);
xnor U37138 (N_37138,N_33016,N_34310);
and U37139 (N_37139,N_32911,N_33585);
and U37140 (N_37140,N_33543,N_34108);
xnor U37141 (N_37141,N_33252,N_34416);
nand U37142 (N_37142,N_34318,N_34398);
and U37143 (N_37143,N_33826,N_33498);
nor U37144 (N_37144,N_33884,N_33419);
or U37145 (N_37145,N_34112,N_32641);
and U37146 (N_37146,N_32860,N_34255);
or U37147 (N_37147,N_33223,N_32543);
nand U37148 (N_37148,N_32933,N_33679);
nand U37149 (N_37149,N_33100,N_34118);
and U37150 (N_37150,N_33225,N_33082);
or U37151 (N_37151,N_34101,N_33354);
and U37152 (N_37152,N_32673,N_34174);
nor U37153 (N_37153,N_34642,N_34854);
xnor U37154 (N_37154,N_33390,N_33631);
nor U37155 (N_37155,N_34946,N_34226);
or U37156 (N_37156,N_32595,N_33945);
nand U37157 (N_37157,N_33783,N_32723);
or U37158 (N_37158,N_33289,N_33421);
or U37159 (N_37159,N_32609,N_34033);
nor U37160 (N_37160,N_34458,N_32612);
or U37161 (N_37161,N_33429,N_32512);
nand U37162 (N_37162,N_34890,N_32730);
and U37163 (N_37163,N_34390,N_32579);
xor U37164 (N_37164,N_33598,N_33305);
xnor U37165 (N_37165,N_32537,N_33787);
nor U37166 (N_37166,N_32952,N_33012);
and U37167 (N_37167,N_33579,N_33438);
nor U37168 (N_37168,N_32885,N_33162);
or U37169 (N_37169,N_34571,N_33498);
nand U37170 (N_37170,N_33906,N_34957);
nor U37171 (N_37171,N_33989,N_32883);
nand U37172 (N_37172,N_33839,N_33333);
and U37173 (N_37173,N_34279,N_34024);
nand U37174 (N_37174,N_33419,N_33964);
and U37175 (N_37175,N_34701,N_33921);
or U37176 (N_37176,N_32649,N_33239);
xor U37177 (N_37177,N_32902,N_33593);
nor U37178 (N_37178,N_32555,N_32780);
or U37179 (N_37179,N_33255,N_34990);
nor U37180 (N_37180,N_33013,N_34773);
or U37181 (N_37181,N_34618,N_34973);
or U37182 (N_37182,N_34348,N_33442);
nor U37183 (N_37183,N_33678,N_33465);
nand U37184 (N_37184,N_33821,N_34476);
and U37185 (N_37185,N_33144,N_33316);
xnor U37186 (N_37186,N_33908,N_33297);
and U37187 (N_37187,N_33385,N_32968);
or U37188 (N_37188,N_32935,N_32642);
nand U37189 (N_37189,N_34402,N_34588);
nor U37190 (N_37190,N_33360,N_33325);
nor U37191 (N_37191,N_33768,N_32766);
nor U37192 (N_37192,N_34573,N_34519);
or U37193 (N_37193,N_33698,N_34529);
xor U37194 (N_37194,N_33997,N_33915);
nand U37195 (N_37195,N_33363,N_33344);
or U37196 (N_37196,N_33373,N_34584);
xor U37197 (N_37197,N_34213,N_32722);
nor U37198 (N_37198,N_34369,N_34541);
xor U37199 (N_37199,N_34956,N_33139);
nor U37200 (N_37200,N_34038,N_33370);
xor U37201 (N_37201,N_34368,N_33720);
and U37202 (N_37202,N_32691,N_33883);
nor U37203 (N_37203,N_32780,N_32797);
and U37204 (N_37204,N_34939,N_33218);
xnor U37205 (N_37205,N_33781,N_32533);
and U37206 (N_37206,N_34332,N_32538);
or U37207 (N_37207,N_34536,N_33767);
and U37208 (N_37208,N_34249,N_34024);
xor U37209 (N_37209,N_34673,N_34094);
nand U37210 (N_37210,N_32522,N_34497);
nand U37211 (N_37211,N_33738,N_32607);
nor U37212 (N_37212,N_34592,N_33195);
xor U37213 (N_37213,N_33906,N_34365);
and U37214 (N_37214,N_34359,N_34558);
and U37215 (N_37215,N_33282,N_34218);
and U37216 (N_37216,N_32519,N_34026);
nand U37217 (N_37217,N_33078,N_33736);
xnor U37218 (N_37218,N_34837,N_33552);
and U37219 (N_37219,N_34143,N_34287);
nor U37220 (N_37220,N_34602,N_34682);
or U37221 (N_37221,N_34660,N_32818);
or U37222 (N_37222,N_34639,N_32673);
nand U37223 (N_37223,N_34967,N_34848);
nor U37224 (N_37224,N_32633,N_34179);
nor U37225 (N_37225,N_33969,N_32930);
nor U37226 (N_37226,N_34253,N_32780);
nand U37227 (N_37227,N_33561,N_33348);
xnor U37228 (N_37228,N_34910,N_34655);
xor U37229 (N_37229,N_33777,N_34481);
xor U37230 (N_37230,N_32665,N_33043);
nand U37231 (N_37231,N_32556,N_34386);
nor U37232 (N_37232,N_33765,N_34487);
nand U37233 (N_37233,N_34321,N_32531);
and U37234 (N_37234,N_33712,N_34960);
and U37235 (N_37235,N_33293,N_33437);
xor U37236 (N_37236,N_32720,N_32661);
or U37237 (N_37237,N_34706,N_33602);
nand U37238 (N_37238,N_32538,N_34209);
nor U37239 (N_37239,N_33564,N_33563);
nor U37240 (N_37240,N_33333,N_34066);
or U37241 (N_37241,N_34225,N_32660);
xnor U37242 (N_37242,N_34917,N_34685);
xor U37243 (N_37243,N_32564,N_34501);
xor U37244 (N_37244,N_32929,N_33577);
and U37245 (N_37245,N_34177,N_32538);
or U37246 (N_37246,N_34001,N_32623);
and U37247 (N_37247,N_34545,N_34936);
or U37248 (N_37248,N_34293,N_34231);
nor U37249 (N_37249,N_33938,N_34901);
nor U37250 (N_37250,N_33559,N_32718);
xnor U37251 (N_37251,N_33339,N_33539);
xnor U37252 (N_37252,N_34287,N_33256);
xnor U37253 (N_37253,N_34547,N_33978);
or U37254 (N_37254,N_34378,N_32615);
nor U37255 (N_37255,N_34413,N_33951);
xnor U37256 (N_37256,N_32792,N_32925);
or U37257 (N_37257,N_34370,N_34064);
nor U37258 (N_37258,N_33599,N_34468);
nor U37259 (N_37259,N_34836,N_33674);
nor U37260 (N_37260,N_32607,N_32588);
or U37261 (N_37261,N_33344,N_32792);
and U37262 (N_37262,N_34078,N_34502);
or U37263 (N_37263,N_34868,N_33730);
and U37264 (N_37264,N_32528,N_34457);
nand U37265 (N_37265,N_34572,N_34593);
and U37266 (N_37266,N_33382,N_33103);
nand U37267 (N_37267,N_34646,N_33020);
nand U37268 (N_37268,N_34618,N_34577);
nand U37269 (N_37269,N_32797,N_33918);
nor U37270 (N_37270,N_34010,N_32772);
xor U37271 (N_37271,N_32976,N_32996);
nor U37272 (N_37272,N_33562,N_34590);
xor U37273 (N_37273,N_33918,N_32868);
and U37274 (N_37274,N_34792,N_32709);
or U37275 (N_37275,N_32893,N_34010);
and U37276 (N_37276,N_34865,N_34463);
or U37277 (N_37277,N_34332,N_33353);
nor U37278 (N_37278,N_33212,N_33665);
nand U37279 (N_37279,N_33490,N_33634);
or U37280 (N_37280,N_32766,N_33293);
nor U37281 (N_37281,N_34892,N_34587);
nor U37282 (N_37282,N_32551,N_34892);
and U37283 (N_37283,N_33272,N_34493);
nor U37284 (N_37284,N_34687,N_33736);
nand U37285 (N_37285,N_34254,N_34825);
nor U37286 (N_37286,N_33709,N_34445);
nor U37287 (N_37287,N_32524,N_32727);
nand U37288 (N_37288,N_34306,N_33855);
or U37289 (N_37289,N_34993,N_34019);
or U37290 (N_37290,N_34482,N_33295);
nor U37291 (N_37291,N_34957,N_34272);
and U37292 (N_37292,N_32778,N_33472);
and U37293 (N_37293,N_33231,N_33281);
nor U37294 (N_37294,N_33791,N_33338);
nand U37295 (N_37295,N_33987,N_34691);
xor U37296 (N_37296,N_33325,N_34462);
nor U37297 (N_37297,N_33756,N_33769);
nand U37298 (N_37298,N_32540,N_32641);
nand U37299 (N_37299,N_34887,N_33221);
nor U37300 (N_37300,N_33754,N_32753);
nand U37301 (N_37301,N_32945,N_32642);
xor U37302 (N_37302,N_34504,N_33416);
nand U37303 (N_37303,N_34522,N_34148);
and U37304 (N_37304,N_33448,N_33022);
or U37305 (N_37305,N_33822,N_32816);
and U37306 (N_37306,N_34755,N_33547);
and U37307 (N_37307,N_32545,N_34314);
xnor U37308 (N_37308,N_34478,N_34361);
nor U37309 (N_37309,N_33429,N_33555);
nand U37310 (N_37310,N_34064,N_33793);
nand U37311 (N_37311,N_33436,N_34412);
xor U37312 (N_37312,N_33614,N_34935);
and U37313 (N_37313,N_34802,N_32690);
xor U37314 (N_37314,N_33376,N_34613);
xor U37315 (N_37315,N_33350,N_33583);
xnor U37316 (N_37316,N_34561,N_33396);
nand U37317 (N_37317,N_33872,N_33340);
and U37318 (N_37318,N_34323,N_33826);
and U37319 (N_37319,N_32634,N_33653);
or U37320 (N_37320,N_33801,N_33205);
nor U37321 (N_37321,N_34875,N_32714);
xor U37322 (N_37322,N_33926,N_33282);
xnor U37323 (N_37323,N_34361,N_33570);
xnor U37324 (N_37324,N_34028,N_33674);
nand U37325 (N_37325,N_33465,N_34994);
nand U37326 (N_37326,N_32903,N_33252);
and U37327 (N_37327,N_34126,N_33196);
nand U37328 (N_37328,N_32745,N_33543);
nand U37329 (N_37329,N_34081,N_34419);
nand U37330 (N_37330,N_33458,N_34809);
xnor U37331 (N_37331,N_34476,N_33931);
or U37332 (N_37332,N_34163,N_33327);
or U37333 (N_37333,N_34941,N_33027);
xor U37334 (N_37334,N_33384,N_34799);
nand U37335 (N_37335,N_32677,N_32597);
nor U37336 (N_37336,N_32792,N_33859);
nor U37337 (N_37337,N_34683,N_33533);
xnor U37338 (N_37338,N_32674,N_34811);
and U37339 (N_37339,N_34272,N_34315);
nand U37340 (N_37340,N_32931,N_34467);
and U37341 (N_37341,N_32648,N_33488);
xnor U37342 (N_37342,N_32843,N_32702);
nor U37343 (N_37343,N_33252,N_33960);
or U37344 (N_37344,N_33964,N_33804);
and U37345 (N_37345,N_34604,N_33730);
xor U37346 (N_37346,N_33823,N_33737);
nand U37347 (N_37347,N_32734,N_33487);
nor U37348 (N_37348,N_34331,N_34299);
nor U37349 (N_37349,N_34660,N_34331);
nand U37350 (N_37350,N_32869,N_32752);
nor U37351 (N_37351,N_32816,N_34508);
xnor U37352 (N_37352,N_34729,N_34645);
xor U37353 (N_37353,N_34455,N_32730);
nand U37354 (N_37354,N_34336,N_34299);
or U37355 (N_37355,N_33503,N_33444);
and U37356 (N_37356,N_34864,N_32907);
and U37357 (N_37357,N_33005,N_33213);
nor U37358 (N_37358,N_33170,N_34850);
and U37359 (N_37359,N_33208,N_34142);
or U37360 (N_37360,N_32571,N_34789);
or U37361 (N_37361,N_33607,N_33394);
nand U37362 (N_37362,N_32642,N_33978);
nand U37363 (N_37363,N_34785,N_33239);
nor U37364 (N_37364,N_34266,N_33400);
nand U37365 (N_37365,N_32577,N_33521);
nor U37366 (N_37366,N_34840,N_33236);
and U37367 (N_37367,N_33751,N_32633);
nand U37368 (N_37368,N_33538,N_34065);
nand U37369 (N_37369,N_33481,N_32577);
and U37370 (N_37370,N_34856,N_34195);
xnor U37371 (N_37371,N_34624,N_33555);
and U37372 (N_37372,N_32588,N_32684);
nor U37373 (N_37373,N_34646,N_34184);
nor U37374 (N_37374,N_33800,N_33927);
nand U37375 (N_37375,N_33011,N_34035);
or U37376 (N_37376,N_33008,N_34849);
and U37377 (N_37377,N_33792,N_34299);
xor U37378 (N_37378,N_32844,N_33426);
nor U37379 (N_37379,N_33042,N_32688);
nand U37380 (N_37380,N_33207,N_33928);
or U37381 (N_37381,N_34471,N_34443);
nor U37382 (N_37382,N_34234,N_34468);
xnor U37383 (N_37383,N_34476,N_33675);
nor U37384 (N_37384,N_33401,N_33297);
nor U37385 (N_37385,N_33670,N_32788);
or U37386 (N_37386,N_33156,N_34206);
nor U37387 (N_37387,N_33122,N_33612);
and U37388 (N_37388,N_34603,N_33108);
nand U37389 (N_37389,N_33103,N_32827);
nor U37390 (N_37390,N_33958,N_34618);
and U37391 (N_37391,N_34311,N_33726);
and U37392 (N_37392,N_33206,N_32641);
and U37393 (N_37393,N_33754,N_33581);
and U37394 (N_37394,N_34836,N_33112);
nand U37395 (N_37395,N_34844,N_32661);
nor U37396 (N_37396,N_34481,N_33459);
nor U37397 (N_37397,N_34441,N_34954);
or U37398 (N_37398,N_33435,N_34545);
or U37399 (N_37399,N_32667,N_33045);
nand U37400 (N_37400,N_32732,N_33981);
nand U37401 (N_37401,N_34007,N_34345);
nor U37402 (N_37402,N_33370,N_34708);
and U37403 (N_37403,N_32980,N_33814);
nor U37404 (N_37404,N_34482,N_33240);
nor U37405 (N_37405,N_33212,N_33659);
and U37406 (N_37406,N_33298,N_34427);
xnor U37407 (N_37407,N_34752,N_33887);
nor U37408 (N_37408,N_34973,N_33669);
nand U37409 (N_37409,N_34058,N_34427);
and U37410 (N_37410,N_33589,N_33286);
nor U37411 (N_37411,N_34883,N_33746);
and U37412 (N_37412,N_34079,N_34567);
nor U37413 (N_37413,N_34657,N_34353);
or U37414 (N_37414,N_33788,N_33523);
xor U37415 (N_37415,N_34360,N_34472);
nand U37416 (N_37416,N_33762,N_32782);
nor U37417 (N_37417,N_34529,N_33719);
and U37418 (N_37418,N_34176,N_33383);
nand U37419 (N_37419,N_34255,N_33929);
or U37420 (N_37420,N_33771,N_34169);
xor U37421 (N_37421,N_34180,N_32923);
and U37422 (N_37422,N_34253,N_34665);
or U37423 (N_37423,N_34379,N_34124);
nor U37424 (N_37424,N_34063,N_34350);
or U37425 (N_37425,N_33886,N_32866);
nor U37426 (N_37426,N_33567,N_33379);
and U37427 (N_37427,N_33161,N_34345);
and U37428 (N_37428,N_33114,N_34416);
nand U37429 (N_37429,N_33466,N_33695);
xor U37430 (N_37430,N_34882,N_34144);
and U37431 (N_37431,N_34041,N_33577);
or U37432 (N_37432,N_32666,N_33419);
nor U37433 (N_37433,N_34208,N_33929);
or U37434 (N_37434,N_34241,N_32559);
and U37435 (N_37435,N_33938,N_33108);
nand U37436 (N_37436,N_34444,N_33124);
nand U37437 (N_37437,N_34721,N_34880);
nand U37438 (N_37438,N_33894,N_32877);
nand U37439 (N_37439,N_33658,N_32649);
or U37440 (N_37440,N_34136,N_34050);
or U37441 (N_37441,N_32543,N_32989);
and U37442 (N_37442,N_32528,N_34368);
nor U37443 (N_37443,N_33715,N_34671);
or U37444 (N_37444,N_34857,N_32757);
nor U37445 (N_37445,N_33285,N_33466);
nor U37446 (N_37446,N_34085,N_34421);
and U37447 (N_37447,N_33052,N_33284);
xor U37448 (N_37448,N_32757,N_33294);
nor U37449 (N_37449,N_32739,N_33431);
and U37450 (N_37450,N_34174,N_34790);
nor U37451 (N_37451,N_32825,N_34063);
nor U37452 (N_37452,N_32812,N_33032);
nor U37453 (N_37453,N_34187,N_33187);
xnor U37454 (N_37454,N_32695,N_33095);
or U37455 (N_37455,N_34170,N_33896);
xor U37456 (N_37456,N_32850,N_34763);
nor U37457 (N_37457,N_34023,N_34574);
or U37458 (N_37458,N_33073,N_34468);
nor U37459 (N_37459,N_32964,N_33317);
and U37460 (N_37460,N_34286,N_34174);
nor U37461 (N_37461,N_34179,N_33068);
and U37462 (N_37462,N_34130,N_33928);
and U37463 (N_37463,N_34770,N_33264);
nand U37464 (N_37464,N_34225,N_33563);
or U37465 (N_37465,N_33036,N_34802);
nand U37466 (N_37466,N_33369,N_33489);
or U37467 (N_37467,N_34168,N_33428);
and U37468 (N_37468,N_34280,N_32765);
or U37469 (N_37469,N_33732,N_33723);
nor U37470 (N_37470,N_33936,N_33911);
nand U37471 (N_37471,N_34211,N_32789);
nor U37472 (N_37472,N_32923,N_33190);
nor U37473 (N_37473,N_33753,N_32659);
nand U37474 (N_37474,N_33276,N_32775);
or U37475 (N_37475,N_34828,N_33364);
nor U37476 (N_37476,N_33543,N_34076);
nand U37477 (N_37477,N_34524,N_32667);
xor U37478 (N_37478,N_34873,N_34939);
xnor U37479 (N_37479,N_32854,N_34020);
nand U37480 (N_37480,N_34222,N_34316);
nor U37481 (N_37481,N_34163,N_33282);
and U37482 (N_37482,N_33413,N_34900);
and U37483 (N_37483,N_32989,N_34600);
nand U37484 (N_37484,N_34008,N_34182);
and U37485 (N_37485,N_33237,N_34499);
or U37486 (N_37486,N_33480,N_33055);
nand U37487 (N_37487,N_33255,N_34105);
nand U37488 (N_37488,N_34575,N_33924);
nor U37489 (N_37489,N_33258,N_32587);
and U37490 (N_37490,N_34094,N_32644);
and U37491 (N_37491,N_32654,N_34896);
and U37492 (N_37492,N_34661,N_33485);
and U37493 (N_37493,N_33623,N_34031);
nand U37494 (N_37494,N_33551,N_34900);
nand U37495 (N_37495,N_33562,N_34483);
nand U37496 (N_37496,N_32950,N_33914);
nor U37497 (N_37497,N_33067,N_34886);
xnor U37498 (N_37498,N_34108,N_33455);
xnor U37499 (N_37499,N_34756,N_34644);
xnor U37500 (N_37500,N_37059,N_36696);
or U37501 (N_37501,N_35632,N_36801);
nand U37502 (N_37502,N_36665,N_36055);
nor U37503 (N_37503,N_35428,N_37462);
or U37504 (N_37504,N_35437,N_37172);
nor U37505 (N_37505,N_37427,N_36941);
or U37506 (N_37506,N_35596,N_35448);
nor U37507 (N_37507,N_35942,N_36682);
nor U37508 (N_37508,N_36384,N_36205);
nor U37509 (N_37509,N_36853,N_36934);
xnor U37510 (N_37510,N_35918,N_35493);
and U37511 (N_37511,N_35525,N_35466);
and U37512 (N_37512,N_36813,N_35575);
xor U37513 (N_37513,N_36578,N_37282);
or U37514 (N_37514,N_36058,N_35584);
xnor U37515 (N_37515,N_36117,N_36534);
nand U37516 (N_37516,N_35974,N_36294);
nand U37517 (N_37517,N_36845,N_35194);
xor U37518 (N_37518,N_35391,N_36353);
and U37519 (N_37519,N_35890,N_36479);
nor U37520 (N_37520,N_35435,N_36252);
nand U37521 (N_37521,N_35908,N_35321);
or U37522 (N_37522,N_36102,N_37486);
or U37523 (N_37523,N_36131,N_37146);
nand U37524 (N_37524,N_36257,N_35062);
nand U37525 (N_37525,N_36328,N_35993);
nand U37526 (N_37526,N_37339,N_36745);
xor U37527 (N_37527,N_35181,N_37474);
nor U37528 (N_37528,N_36130,N_36907);
nor U37529 (N_37529,N_35604,N_35560);
or U37530 (N_37530,N_37034,N_35196);
nand U37531 (N_37531,N_36575,N_36768);
and U37532 (N_37532,N_36604,N_37260);
nor U37533 (N_37533,N_36608,N_35098);
nor U37534 (N_37534,N_35000,N_35893);
nor U37535 (N_37535,N_36126,N_37307);
nor U37536 (N_37536,N_37110,N_35231);
nor U37537 (N_37537,N_35654,N_36743);
and U37538 (N_37538,N_36654,N_36963);
or U37539 (N_37539,N_36798,N_35283);
or U37540 (N_37540,N_36793,N_36748);
nand U37541 (N_37541,N_36705,N_36574);
nor U37542 (N_37542,N_35426,N_36098);
and U37543 (N_37543,N_36546,N_35923);
or U37544 (N_37544,N_35191,N_37297);
and U37545 (N_37545,N_37069,N_36060);
xor U37546 (N_37546,N_36762,N_35701);
and U37547 (N_37547,N_35216,N_36515);
xor U37548 (N_37548,N_35707,N_36557);
xnor U37549 (N_37549,N_36185,N_36389);
xnor U37550 (N_37550,N_37460,N_36022);
and U37551 (N_37551,N_35367,N_36410);
or U37552 (N_37552,N_35325,N_35861);
nor U37553 (N_37553,N_35483,N_36071);
or U37554 (N_37554,N_37021,N_36900);
nand U37555 (N_37555,N_35690,N_35931);
xor U37556 (N_37556,N_36331,N_37176);
or U37557 (N_37557,N_35622,N_37085);
nor U37558 (N_37558,N_35883,N_35223);
and U37559 (N_37559,N_36645,N_37210);
or U37560 (N_37560,N_36489,N_35425);
nor U37561 (N_37561,N_37457,N_37479);
and U37562 (N_37562,N_35753,N_37302);
nor U37563 (N_37563,N_35839,N_36712);
or U37564 (N_37564,N_37405,N_37407);
nor U37565 (N_37565,N_36524,N_36050);
or U37566 (N_37566,N_35869,N_36224);
and U37567 (N_37567,N_35922,N_35468);
or U37568 (N_37568,N_35474,N_35809);
xnor U37569 (N_37569,N_35482,N_35950);
xor U37570 (N_37570,N_35440,N_35305);
and U37571 (N_37571,N_37323,N_37214);
or U37572 (N_37572,N_36258,N_35757);
nand U37573 (N_37573,N_35116,N_37161);
nor U37574 (N_37574,N_35771,N_37006);
and U37575 (N_37575,N_35135,N_37331);
nor U37576 (N_37576,N_36279,N_37100);
or U37577 (N_37577,N_35540,N_35731);
xnor U37578 (N_37578,N_35368,N_36721);
xnor U37579 (N_37579,N_35379,N_37349);
xnor U37580 (N_37580,N_35949,N_36116);
xor U37581 (N_37581,N_35610,N_36263);
or U37582 (N_37582,N_35782,N_35767);
and U37583 (N_37583,N_35306,N_37274);
and U37584 (N_37584,N_36584,N_37238);
xor U37585 (N_37585,N_37099,N_35377);
or U37586 (N_37586,N_36095,N_36713);
nor U37587 (N_37587,N_36357,N_36327);
xor U37588 (N_37588,N_35301,N_36554);
nand U37589 (N_37589,N_36309,N_36520);
nand U37590 (N_37590,N_35565,N_36417);
xor U37591 (N_37591,N_36540,N_36254);
nor U37592 (N_37592,N_35447,N_36732);
and U37593 (N_37593,N_35322,N_35381);
xnor U37594 (N_37594,N_35928,N_35968);
xnor U37595 (N_37595,N_35759,N_35794);
and U37596 (N_37596,N_35095,N_35746);
nand U37597 (N_37597,N_36396,N_36607);
or U37598 (N_37598,N_35834,N_35264);
nand U37599 (N_37599,N_36716,N_37004);
or U37600 (N_37600,N_37228,N_35108);
nand U37601 (N_37601,N_35775,N_36538);
xor U37602 (N_37602,N_35516,N_36037);
nand U37603 (N_37603,N_35197,N_36306);
xor U37604 (N_37604,N_37366,N_36483);
and U37605 (N_37605,N_36218,N_35154);
or U37606 (N_37606,N_35595,N_36985);
nand U37607 (N_37607,N_36502,N_36176);
or U37608 (N_37608,N_37338,N_35518);
and U37609 (N_37609,N_36231,N_36191);
xor U37610 (N_37610,N_35532,N_35768);
or U37611 (N_37611,N_35157,N_36916);
or U37612 (N_37612,N_36339,N_36455);
nand U37613 (N_37613,N_36457,N_37488);
nand U37614 (N_37614,N_35339,N_35290);
nor U37615 (N_37615,N_36882,N_35805);
or U37616 (N_37616,N_37009,N_37163);
nand U37617 (N_37617,N_35599,N_35681);
and U37618 (N_37618,N_36655,N_37361);
or U37619 (N_37619,N_37375,N_36175);
and U37620 (N_37620,N_37255,N_35851);
and U37621 (N_37621,N_36507,N_36173);
or U37622 (N_37622,N_35469,N_35708);
xor U37623 (N_37623,N_35970,N_35549);
xor U37624 (N_37624,N_36246,N_35651);
nand U37625 (N_37625,N_36307,N_36083);
xnor U37626 (N_37626,N_36987,N_36349);
and U37627 (N_37627,N_36045,N_36372);
xnor U37628 (N_37628,N_37154,N_36454);
nand U37629 (N_37629,N_35750,N_37045);
nor U37630 (N_37630,N_36319,N_36487);
and U37631 (N_37631,N_36204,N_36089);
nand U37632 (N_37632,N_35462,N_35854);
nand U37633 (N_37633,N_37064,N_35311);
nor U37634 (N_37634,N_35100,N_35323);
nand U37635 (N_37635,N_37352,N_35357);
and U37636 (N_37636,N_35300,N_36125);
nand U37637 (N_37637,N_35998,N_35760);
and U37638 (N_37638,N_35395,N_36458);
xnor U37639 (N_37639,N_36613,N_36780);
or U37640 (N_37640,N_37434,N_36829);
nor U37641 (N_37641,N_36562,N_35074);
and U37642 (N_37642,N_37308,N_36409);
nand U37643 (N_37643,N_35199,N_37256);
xnor U37644 (N_37644,N_35667,N_36572);
nor U37645 (N_37645,N_36838,N_36744);
xnor U37646 (N_37646,N_36332,N_35378);
and U37647 (N_37647,N_37396,N_36035);
nor U37648 (N_37648,N_37335,N_35067);
xor U37649 (N_37649,N_37314,N_37092);
nand U37650 (N_37650,N_35173,N_37478);
and U37651 (N_37651,N_36844,N_35491);
and U37652 (N_37652,N_37429,N_36430);
nor U37653 (N_37653,N_37079,N_35414);
nor U37654 (N_37654,N_37195,N_37327);
or U37655 (N_37655,N_35939,N_36761);
nor U37656 (N_37656,N_35871,N_36817);
and U37657 (N_37657,N_35886,N_36677);
xor U37658 (N_37658,N_35788,N_37179);
xor U37659 (N_37659,N_35719,N_35246);
nor U37660 (N_37660,N_36955,N_36898);
nor U37661 (N_37661,N_36397,N_35606);
xnor U37662 (N_37662,N_36542,N_35398);
nand U37663 (N_37663,N_37048,N_36108);
nor U37664 (N_37664,N_36788,N_36657);
or U37665 (N_37665,N_35802,N_36912);
or U37666 (N_37666,N_37395,N_37261);
nor U37667 (N_37667,N_36196,N_35025);
nand U37668 (N_37668,N_35592,N_35644);
or U37669 (N_37669,N_35119,N_35044);
or U37670 (N_37670,N_36565,N_36596);
or U37671 (N_37671,N_36106,N_36541);
nor U37672 (N_37672,N_35253,N_37053);
or U37673 (N_37673,N_36476,N_36425);
nor U37674 (N_37674,N_37270,N_35914);
xor U37675 (N_37675,N_36449,N_36025);
nor U37676 (N_37676,N_37466,N_36787);
and U37677 (N_37677,N_35542,N_36105);
nand U37678 (N_37678,N_36200,N_36090);
and U37679 (N_37679,N_36895,N_36351);
nand U37680 (N_37680,N_37286,N_36730);
xor U37681 (N_37681,N_36627,N_36300);
or U37682 (N_37682,N_35046,N_36513);
and U37683 (N_37683,N_36234,N_35724);
xor U37684 (N_37684,N_37216,N_36874);
nor U37685 (N_37685,N_35977,N_36031);
nand U37686 (N_37686,N_36765,N_35415);
nor U37687 (N_37687,N_36301,N_35439);
nand U37688 (N_37688,N_35084,N_35385);
or U37689 (N_37689,N_36796,N_35783);
or U37690 (N_37690,N_36411,N_35093);
nand U37691 (N_37691,N_35781,N_36889);
xnor U37692 (N_37692,N_36774,N_35504);
xor U37693 (N_37693,N_36690,N_35139);
xnor U37694 (N_37694,N_35294,N_37249);
or U37695 (N_37695,N_37277,N_35513);
or U37696 (N_37696,N_37469,N_35992);
xnor U37697 (N_37697,N_35186,N_35444);
or U37698 (N_37698,N_36533,N_35740);
or U37699 (N_37699,N_35699,N_37357);
or U37700 (N_37700,N_37083,N_35501);
nand U37701 (N_37701,N_36352,N_35778);
xnor U37702 (N_37702,N_36436,N_35296);
nor U37703 (N_37703,N_36333,N_35387);
and U37704 (N_37704,N_36904,N_35240);
and U37705 (N_37705,N_36381,N_37119);
nor U37706 (N_37706,N_35383,N_36752);
nand U37707 (N_37707,N_35929,N_36511);
nand U37708 (N_37708,N_37380,N_36982);
or U37709 (N_37709,N_37328,N_35784);
nand U37710 (N_37710,N_37279,N_36265);
xor U37711 (N_37711,N_36441,N_36662);
xor U37712 (N_37712,N_37337,N_35293);
nor U37713 (N_37713,N_37171,N_36416);
nand U37714 (N_37714,N_37485,N_36085);
and U37715 (N_37715,N_36617,N_36529);
or U37716 (N_37716,N_37444,N_35487);
xor U37717 (N_37717,N_36018,N_35571);
and U37718 (N_37718,N_35944,N_36851);
and U37719 (N_37719,N_35113,N_35582);
and U37720 (N_37720,N_36532,N_37467);
or U37721 (N_37721,N_35262,N_36104);
and U37722 (N_37722,N_35676,N_35517);
nor U37723 (N_37723,N_35099,N_36836);
nor U37724 (N_37724,N_36053,N_35712);
or U37725 (N_37725,N_35049,N_36870);
nor U37726 (N_37726,N_35075,N_35018);
nor U37727 (N_37727,N_37437,N_35665);
xor U37728 (N_37728,N_37203,N_36118);
xnor U37729 (N_37729,N_35351,N_35408);
xnor U37730 (N_37730,N_35506,N_35967);
and U37731 (N_37731,N_36274,N_35524);
xor U37732 (N_37732,N_36506,N_35069);
and U37733 (N_37733,N_35105,N_35058);
or U37734 (N_37734,N_35616,N_35983);
nor U37735 (N_37735,N_36114,N_36247);
nor U37736 (N_37736,N_35765,N_36299);
nand U37737 (N_37737,N_36858,N_36868);
and U37738 (N_37738,N_37186,N_35295);
and U37739 (N_37739,N_35123,N_36147);
xnor U37740 (N_37740,N_35239,N_37109);
xor U37741 (N_37741,N_35176,N_35243);
or U37742 (N_37742,N_35146,N_37042);
xor U37743 (N_37743,N_35118,N_36791);
and U37744 (N_37744,N_36717,N_36886);
nand U37745 (N_37745,N_36504,N_35530);
nor U37746 (N_37746,N_35898,N_35894);
nand U37747 (N_37747,N_37231,N_37017);
nor U37748 (N_37748,N_37329,N_35177);
nand U37749 (N_37749,N_35636,N_35973);
xnor U37750 (N_37750,N_37152,N_36275);
xor U37751 (N_37751,N_35372,N_36350);
nand U37752 (N_37752,N_35637,N_36129);
or U37753 (N_37753,N_36293,N_35688);
nor U37754 (N_37754,N_36818,N_37254);
xor U37755 (N_37755,N_36312,N_36977);
and U37756 (N_37756,N_36920,N_36624);
and U37757 (N_37757,N_36519,N_36924);
nand U37758 (N_37758,N_36028,N_35892);
or U37759 (N_37759,N_35235,N_37304);
and U37760 (N_37760,N_36827,N_35954);
or U37761 (N_37761,N_35732,N_37298);
or U37762 (N_37762,N_36637,N_36576);
and U37763 (N_37763,N_36004,N_36582);
or U37764 (N_37764,N_36623,N_36733);
or U37765 (N_37765,N_37465,N_35334);
nand U37766 (N_37766,N_35124,N_35526);
or U37767 (N_37767,N_36133,N_36424);
xor U37768 (N_37768,N_35583,N_35836);
and U37769 (N_37769,N_36428,N_36297);
and U37770 (N_37770,N_36531,N_35319);
xnor U37771 (N_37771,N_35111,N_37322);
xor U37772 (N_37772,N_35745,N_36505);
or U37773 (N_37773,N_35029,N_36356);
xnor U37774 (N_37774,N_37359,N_36390);
or U37775 (N_37775,N_36481,N_37477);
nor U37776 (N_37776,N_36544,N_36651);
nor U37777 (N_37777,N_36824,N_37105);
nand U37778 (N_37778,N_37062,N_35133);
and U37779 (N_37779,N_37019,N_35060);
nand U37780 (N_37780,N_35373,N_35608);
nor U37781 (N_37781,N_36440,N_37334);
nor U37782 (N_37782,N_36587,N_35503);
or U37783 (N_37783,N_35885,N_37011);
and U37784 (N_37784,N_36634,N_36686);
and U37785 (N_37785,N_35866,N_35442);
nor U37786 (N_37786,N_36268,N_37002);
xnor U37787 (N_37787,N_36940,N_36992);
xnor U37788 (N_37788,N_37187,N_36650);
nand U37789 (N_37789,N_36986,N_35849);
xor U37790 (N_37790,N_35392,N_36049);
xnor U37791 (N_37791,N_36860,N_36629);
nand U37792 (N_37792,N_35590,N_37393);
nand U37793 (N_37793,N_37151,N_36567);
nand U37794 (N_37794,N_35159,N_37050);
nand U37795 (N_37795,N_35835,N_36610);
xor U37796 (N_37796,N_37257,N_36719);
or U37797 (N_37797,N_35508,N_35292);
nor U37798 (N_37798,N_35104,N_36722);
or U37799 (N_37799,N_36280,N_37184);
or U37800 (N_37800,N_37449,N_35635);
xor U37801 (N_37801,N_35572,N_36073);
or U37802 (N_37802,N_36221,N_35451);
and U37803 (N_37803,N_36207,N_35152);
or U37804 (N_37804,N_36571,N_35634);
nor U37805 (N_37805,N_35975,N_36526);
or U37806 (N_37806,N_35936,N_37311);
and U37807 (N_37807,N_36959,N_35902);
and U37808 (N_37808,N_36242,N_36566);
nand U37809 (N_37809,N_36849,N_36426);
or U37810 (N_37810,N_36805,N_36387);
xor U37811 (N_37811,N_36290,N_37497);
nand U37812 (N_37812,N_35536,N_35207);
xor U37813 (N_37813,N_35271,N_36121);
and U37814 (N_37814,N_36543,N_35945);
or U37815 (N_37815,N_36020,N_35711);
nor U37816 (N_37816,N_37007,N_36096);
or U37817 (N_37817,N_37026,N_36194);
and U37818 (N_37818,N_35999,N_35338);
nand U37819 (N_37819,N_37234,N_36420);
nor U37820 (N_37820,N_37267,N_36676);
nor U37821 (N_37821,N_35495,N_35416);
and U37822 (N_37822,N_35820,N_36151);
nand U37823 (N_37823,N_37262,N_35318);
xor U37824 (N_37824,N_37354,N_35882);
or U37825 (N_37825,N_36742,N_35958);
nor U37826 (N_37826,N_35865,N_35255);
xor U37827 (N_37827,N_35934,N_36876);
nor U37828 (N_37828,N_35369,N_35042);
nand U37829 (N_37829,N_36172,N_37067);
xnor U37830 (N_37830,N_35718,N_36418);
or U37831 (N_37831,N_36896,N_36235);
xnor U37832 (N_37832,N_35136,N_37072);
nor U37833 (N_37833,N_35407,N_35717);
and U37834 (N_37834,N_37039,N_36379);
or U37835 (N_37835,N_35714,N_36517);
xnor U37836 (N_37836,N_36848,N_35988);
and U37837 (N_37837,N_35204,N_36021);
xnor U37838 (N_37838,N_37223,N_37197);
and U37839 (N_37839,N_35022,N_35940);
or U37840 (N_37840,N_36163,N_37020);
nand U37841 (N_37841,N_36412,N_35182);
and U37842 (N_37842,N_35057,N_35709);
xnor U37843 (N_37843,N_36974,N_35241);
nor U37844 (N_37844,N_35404,N_35484);
xor U37845 (N_37845,N_35863,N_37406);
or U37846 (N_37846,N_37480,N_35336);
nor U37847 (N_37847,N_37446,N_36972);
xnor U37848 (N_37848,N_36497,N_35997);
xor U37849 (N_37849,N_37420,N_36820);
xor U37850 (N_37850,N_35303,N_35964);
xnor U37851 (N_37851,N_36148,N_35629);
xor U37852 (N_37852,N_37247,N_35638);
nor U37853 (N_37853,N_35756,N_35680);
xnor U37854 (N_37854,N_36447,N_35662);
xor U37855 (N_37855,N_36112,N_35003);
nand U37856 (N_37856,N_37229,N_36983);
nor U37857 (N_37857,N_36318,N_36086);
and U37858 (N_37858,N_35742,N_35803);
xnor U37859 (N_37859,N_36622,N_37350);
or U37860 (N_37860,N_35653,N_35147);
and U37861 (N_37861,N_35800,N_35647);
nand U37862 (N_37862,N_37213,N_35926);
nor U37863 (N_37863,N_35424,N_36530);
xor U37864 (N_37864,N_36468,N_36181);
nor U37865 (N_37865,N_36282,N_35729);
or U37866 (N_37866,N_36228,N_35762);
nor U37867 (N_37867,N_35669,N_35256);
nor U37868 (N_37868,N_36249,N_35683);
and U37869 (N_37869,N_35457,N_35804);
nor U37870 (N_37870,N_36781,N_35728);
and U37871 (N_37871,N_35278,N_36678);
nand U37872 (N_37872,N_37374,N_36570);
nor U37873 (N_37873,N_37284,N_36388);
and U37874 (N_37874,N_37381,N_37095);
or U37875 (N_37875,N_36492,N_37028);
xnor U37876 (N_37876,N_35780,N_35382);
nand U37877 (N_37877,N_35153,N_35808);
or U37878 (N_37878,N_37456,N_35073);
xnor U37879 (N_37879,N_35848,N_36832);
and U37880 (N_37880,N_35826,N_35024);
nor U37881 (N_37881,N_37343,N_36407);
or U37882 (N_37882,N_37201,N_37453);
nor U37883 (N_37883,N_35043,N_36270);
xnor U37884 (N_37884,N_35365,N_36585);
or U37885 (N_37885,N_35642,N_36731);
and U37886 (N_37886,N_35556,N_35006);
nor U37887 (N_37887,N_36683,N_36673);
nor U37888 (N_37888,N_35257,N_35823);
nor U37889 (N_37889,N_35916,N_36495);
nor U37890 (N_37890,N_35071,N_36843);
xor U37891 (N_37891,N_35456,N_36638);
and U37892 (N_37892,N_37190,N_35393);
xnor U37893 (N_37893,N_36128,N_36099);
nand U37894 (N_37894,N_35219,N_35737);
or U37895 (N_37895,N_36559,N_35646);
and U37896 (N_37896,N_37130,N_36999);
nor U37897 (N_37897,N_37475,N_36536);
nand U37898 (N_37898,N_35769,N_37271);
xnor U37899 (N_37899,N_35314,N_35758);
nand U37900 (N_37900,N_36210,N_35661);
or U37901 (N_37901,N_35289,N_36736);
and U37902 (N_37902,N_36925,N_36630);
xnor U37903 (N_37903,N_36808,N_35577);
and U37904 (N_37904,N_35664,N_35362);
nor U37905 (N_37905,N_35692,N_36041);
and U37906 (N_37906,N_36758,N_36757);
or U37907 (N_37907,N_35344,N_37060);
or U37908 (N_37908,N_35254,N_36819);
and U37909 (N_37909,N_37240,N_35534);
nor U37910 (N_37910,N_37442,N_35879);
nand U37911 (N_37911,N_35266,N_35041);
and U37912 (N_37912,N_36568,N_35412);
or U37913 (N_37913,N_37204,N_37040);
xnor U37914 (N_37914,N_37402,N_36222);
or U37915 (N_37915,N_35141,N_36563);
and U37916 (N_37916,N_35609,N_36369);
and U37917 (N_37917,N_37330,N_35706);
nand U37918 (N_37918,N_37386,N_35335);
or U37919 (N_37919,N_35340,N_36726);
and U37920 (N_37920,N_37394,N_35087);
nand U37921 (N_37921,N_35269,N_35380);
and U37922 (N_37922,N_36421,N_37022);
nand U37923 (N_37923,N_36165,N_36399);
xor U37924 (N_37924,N_37447,N_36550);
and U37925 (N_37925,N_37455,N_35063);
nor U37926 (N_37926,N_36913,N_36494);
nor U37927 (N_37927,N_37476,N_36291);
and U37928 (N_37928,N_36932,N_37180);
and U37929 (N_37929,N_36644,N_36398);
xor U37930 (N_37930,N_35109,N_35546);
and U37931 (N_37931,N_36363,N_36434);
or U37932 (N_37932,N_37142,N_36993);
nand U37933 (N_37933,N_37178,N_36149);
and U37934 (N_37934,N_36684,N_36144);
nor U37935 (N_37935,N_37451,N_36664);
and U37936 (N_37936,N_35443,N_36700);
or U37937 (N_37937,N_35224,N_35431);
nand U37938 (N_37938,N_35567,N_36179);
and U37939 (N_37939,N_37133,N_37324);
or U37940 (N_37940,N_36636,N_37463);
xnor U37941 (N_37941,N_37252,N_37183);
or U37942 (N_37942,N_36834,N_36602);
nand U37943 (N_37943,N_37244,N_36667);
and U37944 (N_37944,N_35110,N_37287);
nand U37945 (N_37945,N_37345,N_37208);
or U37946 (N_37946,N_35862,N_37086);
nor U37947 (N_37947,N_35117,N_35966);
nand U37948 (N_37948,N_36749,N_37077);
nor U37949 (N_37949,N_35170,N_36658);
xor U37950 (N_37950,N_37097,N_36463);
or U37951 (N_37951,N_37278,N_36770);
nor U37952 (N_37952,N_35817,N_35238);
xor U37953 (N_37953,N_35739,N_35617);
nor U37954 (N_37954,N_36219,N_35285);
or U37955 (N_37955,N_35354,N_35352);
or U37956 (N_37956,N_36152,N_36438);
nand U37957 (N_37957,N_36815,N_35502);
and U37958 (N_37958,N_37364,N_37242);
nor U37959 (N_37959,N_35402,N_36915);
xor U37960 (N_37960,N_37473,N_35920);
and U37961 (N_37961,N_37403,N_37108);
xnor U37962 (N_37962,N_36360,N_37090);
or U37963 (N_37963,N_35716,N_36718);
nor U37964 (N_37964,N_37448,N_36042);
xor U37965 (N_37965,N_37241,N_35735);
xnor U37966 (N_37966,N_36512,N_36954);
xnor U37967 (N_37967,N_36668,N_35030);
nand U37968 (N_37968,N_36267,N_35001);
nand U37969 (N_37969,N_35734,N_35976);
nand U37970 (N_37970,N_36694,N_35326);
nand U37971 (N_37971,N_36230,N_35593);
or U37972 (N_37972,N_35397,N_37325);
nor U37973 (N_37973,N_35023,N_35260);
nand U37974 (N_37974,N_37464,N_36475);
xnor U37975 (N_37975,N_35658,N_37112);
and U37976 (N_37976,N_36653,N_37399);
xnor U37977 (N_37977,N_36140,N_37008);
and U37978 (N_37978,N_35276,N_37232);
or U37979 (N_37979,N_35010,N_35088);
and U37980 (N_37980,N_36797,N_35671);
and U37981 (N_37981,N_36107,N_35052);
or U37982 (N_37982,N_36659,N_35247);
xnor U37983 (N_37983,N_35772,N_35843);
or U37984 (N_37984,N_36439,N_36317);
and U37985 (N_37985,N_36551,N_37319);
or U37986 (N_37986,N_36581,N_35366);
and U37987 (N_37987,N_36879,N_37088);
xor U37988 (N_37988,N_36897,N_37377);
nor U37989 (N_37989,N_36324,N_35488);
or U37990 (N_37990,N_36910,N_35656);
nor U37991 (N_37991,N_36437,N_37114);
nor U37992 (N_37992,N_35915,N_36253);
or U37993 (N_37993,N_37205,N_36064);
nand U37994 (N_37994,N_35150,N_36632);
nor U37995 (N_37995,N_35206,N_35055);
xnor U37996 (N_37996,N_37342,N_35037);
nor U37997 (N_37997,N_36887,N_37264);
xnor U37998 (N_37998,N_36579,N_37397);
xnor U37999 (N_37999,N_36609,N_37372);
or U38000 (N_38000,N_35703,N_35519);
and U38001 (N_38001,N_35065,N_36036);
nor U38002 (N_38002,N_37421,N_35568);
or U38003 (N_38003,N_37436,N_37189);
nor U38004 (N_38004,N_35685,N_36776);
nand U38005 (N_38005,N_37078,N_36588);
xnor U38006 (N_38006,N_35574,N_35905);
nand U38007 (N_38007,N_35014,N_37235);
nand U38008 (N_38008,N_37226,N_35467);
and U38009 (N_38009,N_35102,N_35528);
nand U38010 (N_38010,N_35704,N_35091);
xnor U38011 (N_38011,N_37376,N_36217);
or U38012 (N_38012,N_35573,N_36043);
xnor U38013 (N_38013,N_36600,N_37268);
and U38014 (N_38014,N_36334,N_36012);
nand U38015 (N_38015,N_36672,N_35092);
and U38016 (N_38016,N_35356,N_37344);
and U38017 (N_38017,N_37458,N_37428);
or U38018 (N_38018,N_36192,N_36141);
xnor U38019 (N_38019,N_35185,N_35831);
or U38020 (N_38020,N_35650,N_37459);
nor U38021 (N_38021,N_36288,N_37346);
nor U38022 (N_38022,N_35956,N_35396);
and U38023 (N_38023,N_37369,N_35315);
nor U38024 (N_38024,N_37104,N_36976);
and U38025 (N_38025,N_35012,N_37347);
nand U38026 (N_38026,N_36008,N_36866);
nor U38027 (N_38027,N_35148,N_36755);
nor U38028 (N_38028,N_36703,N_35844);
xor U38029 (N_38029,N_35189,N_35522);
nor U38030 (N_38030,N_36374,N_37248);
xnor U38031 (N_38031,N_35143,N_37415);
or U38032 (N_38032,N_36804,N_35492);
nor U38033 (N_38033,N_36990,N_37076);
or U38034 (N_38034,N_37117,N_35138);
nor U38035 (N_38035,N_35816,N_37082);
nor U38036 (N_38036,N_35050,N_36698);
xnor U38037 (N_38037,N_36273,N_36134);
nand U38038 (N_38038,N_36995,N_35543);
xnor U38039 (N_38039,N_37299,N_35245);
and U38040 (N_38040,N_35078,N_36038);
xnor U38041 (N_38041,N_35870,N_36044);
xnor U38042 (N_38042,N_36997,N_35188);
and U38043 (N_38043,N_37182,N_37222);
and U38044 (N_38044,N_35691,N_36209);
and U38045 (N_38045,N_35792,N_36782);
and U38046 (N_38046,N_37055,N_36652);
xnor U38047 (N_38047,N_36996,N_35770);
nor U38048 (N_38048,N_36891,N_37321);
nand U38049 (N_38049,N_35215,N_35162);
nand U38050 (N_38050,N_36097,N_37207);
xor U38051 (N_38051,N_37058,N_35218);
nor U38052 (N_38052,N_36244,N_35625);
and U38053 (N_38053,N_36320,N_35878);
and U38054 (N_38054,N_36178,N_37124);
nor U38055 (N_38055,N_36516,N_35490);
xnor U38056 (N_38056,N_37200,N_35569);
nand U38057 (N_38057,N_36281,N_36326);
nor U38058 (N_38058,N_36928,N_36861);
and U38059 (N_38059,N_35830,N_36078);
nand U38060 (N_38060,N_36942,N_36156);
nand U38061 (N_38061,N_35220,N_35566);
or U38062 (N_38062,N_37269,N_37418);
or U38063 (N_38063,N_35476,N_36456);
or U38064 (N_38064,N_36142,N_35059);
nand U38065 (N_38065,N_36867,N_36110);
nor U38066 (N_38066,N_35361,N_36186);
and U38067 (N_38067,N_36549,N_36278);
or U38068 (N_38068,N_36556,N_35747);
nand U38069 (N_38069,N_35722,N_36598);
nor U38070 (N_38070,N_35279,N_36182);
and U38071 (N_38071,N_35054,N_35013);
or U38072 (N_38072,N_37320,N_36965);
nand U38073 (N_38073,N_35535,N_35298);
nand U38074 (N_38074,N_36949,N_35537);
nor U38075 (N_38075,N_36558,N_35715);
nand U38076 (N_38076,N_36366,N_35790);
and U38077 (N_38077,N_37046,N_35700);
nor U38078 (N_38078,N_36792,N_36577);
nand U38079 (N_38079,N_35263,N_36966);
nor U38080 (N_38080,N_36295,N_36383);
and U38081 (N_38081,N_36767,N_36548);
nand U38082 (N_38082,N_36346,N_36052);
and U38083 (N_38083,N_36400,N_37236);
xor U38084 (N_38084,N_35873,N_35827);
and U38085 (N_38085,N_35570,N_35277);
or U38086 (N_38086,N_36701,N_35620);
and U38087 (N_38087,N_35164,N_36777);
nand U38088 (N_38088,N_35880,N_35748);
and U38089 (N_38089,N_35910,N_36612);
nor U38090 (N_38090,N_35364,N_36011);
nand U38091 (N_38091,N_37175,N_37051);
nor U38092 (N_38092,N_36302,N_35841);
xnor U38093 (N_38093,N_36337,N_36828);
and U38094 (N_38094,N_35019,N_36303);
or U38095 (N_38095,N_36378,N_35004);
nor U38096 (N_38096,N_37385,N_36408);
nand U38097 (N_38097,N_36880,N_35813);
nor U38098 (N_38098,N_36127,N_37181);
nand U38099 (N_38099,N_36074,N_37035);
and U38100 (N_38100,N_36922,N_37496);
or U38101 (N_38101,N_37360,N_36573);
xnor U38102 (N_38102,N_36030,N_36616);
and U38103 (N_38103,N_35581,N_35472);
and U38104 (N_38104,N_35209,N_36092);
xnor U38105 (N_38105,N_37378,N_35589);
or U38106 (N_38106,N_36856,N_36539);
nor U38107 (N_38107,N_35554,N_37266);
or U38108 (N_38108,N_36753,N_35579);
or U38109 (N_38109,N_35979,N_35829);
xnor U38110 (N_38110,N_35913,N_35270);
nor U38111 (N_38111,N_35932,N_35497);
nor U38112 (N_38112,N_37024,N_35273);
nand U38113 (N_38113,N_35461,N_36693);
xor U38114 (N_38114,N_35411,N_35796);
or U38115 (N_38115,N_36039,N_37016);
nand U38116 (N_38116,N_35896,N_35376);
or U38117 (N_38117,N_37111,N_36710);
nand U38118 (N_38118,N_35520,N_37071);
and U38119 (N_38119,N_36310,N_36935);
and U38120 (N_38120,N_35499,N_35114);
or U38121 (N_38121,N_36341,N_36795);
nor U38122 (N_38122,N_37013,N_35072);
or U38123 (N_38123,N_37296,N_37401);
or U38124 (N_38124,N_36518,N_37227);
xor U38125 (N_38125,N_37273,N_36462);
nor U38126 (N_38126,N_36474,N_36484);
xor U38127 (N_38127,N_35251,N_37313);
nand U38128 (N_38128,N_36523,N_35389);
xnor U38129 (N_38129,N_35384,N_36689);
nand U38130 (N_38130,N_35957,N_35132);
nand U38131 (N_38131,N_35666,N_37263);
nor U38132 (N_38132,N_36062,N_35248);
nand U38133 (N_38133,N_35810,N_36169);
nand U38134 (N_38134,N_37239,N_35496);
nand U38135 (N_38135,N_35807,N_37057);
or U38136 (N_38136,N_36066,N_36150);
or U38137 (N_38137,N_36075,N_35555);
nand U38138 (N_38138,N_36720,N_36227);
and U38139 (N_38139,N_37145,N_37103);
xor U38140 (N_38140,N_35452,N_35106);
nand U38141 (N_38141,N_35192,N_36211);
nand U38142 (N_38142,N_37276,N_35175);
nand U38143 (N_38143,N_36735,N_36451);
nand U38144 (N_38144,N_36248,N_35034);
nand U38145 (N_38145,N_35056,N_35470);
xor U38146 (N_38146,N_36422,N_35838);
nand U38147 (N_38147,N_36783,N_36271);
or U38148 (N_38148,N_36081,N_36803);
nand U38149 (N_38149,N_35847,N_35859);
xnor U38150 (N_38150,N_37162,N_35213);
nor U38151 (N_38151,N_36670,N_36296);
nor U38152 (N_38152,N_36766,N_36498);
xor U38153 (N_38153,N_36994,N_36100);
xnor U38154 (N_38154,N_35125,N_36206);
nand U38155 (N_38155,N_36260,N_37305);
or U38156 (N_38156,N_36404,N_36419);
xnor U38157 (N_38157,N_35374,N_35015);
and U38158 (N_38158,N_36485,N_36878);
nor U38159 (N_38159,N_35674,N_35252);
and U38160 (N_38160,N_36527,N_37440);
or U38161 (N_38161,N_35232,N_37233);
and U38162 (N_38162,N_35002,N_35811);
and U38163 (N_38163,N_37295,N_37259);
or U38164 (N_38164,N_36681,N_36431);
nor U38165 (N_38165,N_36823,N_35203);
nor U38166 (N_38166,N_36737,N_35302);
nor U38167 (N_38167,N_35070,N_36111);
nand U38168 (N_38168,N_35127,N_36939);
nor U38169 (N_38169,N_36979,N_36153);
nor U38170 (N_38170,N_36875,N_37202);
xnor U38171 (N_38171,N_36706,N_35801);
and U38172 (N_38172,N_36162,N_36646);
nor U38173 (N_38173,N_37414,N_36811);
nand U38174 (N_38174,N_36168,N_35234);
and U38175 (N_38175,N_36139,N_35359);
xnor U38176 (N_38176,N_36771,N_35621);
nor U38177 (N_38177,N_35268,N_35749);
nor U38178 (N_38178,N_37424,N_35134);
and U38179 (N_38179,N_36514,N_36382);
xor U38180 (N_38180,N_36229,N_36313);
or U38181 (N_38181,N_37192,N_35833);
nor U38182 (N_38182,N_35670,N_35587);
nand U38183 (N_38183,N_35464,N_37383);
or U38184 (N_38184,N_35272,N_37056);
nand U38185 (N_38185,N_36593,N_35422);
and U38186 (N_38186,N_35168,N_36830);
and U38187 (N_38187,N_36552,N_35562);
nand U38188 (N_38188,N_36998,N_37221);
xnor U38189 (N_38189,N_35190,N_36189);
and U38190 (N_38190,N_35872,N_36482);
xor U38191 (N_38191,N_35580,N_36591);
nor U38192 (N_38192,N_35948,N_35096);
or U38193 (N_38193,N_37315,N_35481);
nor U38194 (N_38194,N_35853,N_37294);
xnor U38195 (N_38195,N_36255,N_36814);
nand U38196 (N_38196,N_36873,N_36298);
xnor U38197 (N_38197,N_35333,N_35721);
nand U38198 (N_38198,N_35463,N_35846);
nor U38199 (N_38199,N_36927,N_35375);
and U38200 (N_38200,N_35040,N_35751);
xnor U38201 (N_38201,N_35094,N_36145);
or U38202 (N_38202,N_35971,N_36070);
xor U38203 (N_38203,N_37218,N_36699);
or U38204 (N_38204,N_35982,N_37126);
xor U38205 (N_38205,N_35287,N_35969);
or U38206 (N_38206,N_36902,N_36286);
xor U38207 (N_38207,N_35630,N_35479);
nand U38208 (N_38208,N_36340,N_36821);
xnor U38209 (N_38209,N_36013,N_35909);
and U38210 (N_38210,N_36981,N_37141);
and U38211 (N_38211,N_35837,N_36950);
xnor U38212 (N_38212,N_36358,N_35126);
or U38213 (N_38213,N_36119,N_36348);
nand U38214 (N_38214,N_35512,N_35510);
and U38215 (N_38215,N_35744,N_36330);
nand U38216 (N_38216,N_35618,N_36167);
nand U38217 (N_38217,N_37373,N_36946);
nand U38218 (N_38218,N_37164,N_37115);
nand U38219 (N_38219,N_35927,N_36812);
nand U38220 (N_38220,N_37290,N_36061);
nor U38221 (N_38221,N_35498,N_35349);
xnor U38222 (N_38222,N_35980,N_36921);
nor U38223 (N_38223,N_35614,N_36423);
nand U38224 (N_38224,N_35868,N_36738);
xor U38225 (N_38225,N_36007,N_36087);
nand U38226 (N_38226,N_35538,N_36459);
xor U38227 (N_38227,N_37454,N_35995);
xnor U38228 (N_38228,N_37159,N_37326);
nand U38229 (N_38229,N_35304,N_35005);
nand U38230 (N_38230,N_36314,N_35237);
nand U38231 (N_38231,N_36894,N_37143);
or U38232 (N_38232,N_36480,N_36989);
or U38233 (N_38233,N_36709,N_35605);
or U38234 (N_38234,N_36452,N_37155);
nand U38235 (N_38235,N_36138,N_37355);
nand U38236 (N_38236,N_35112,N_36839);
nor U38237 (N_38237,N_35332,N_36970);
or U38238 (N_38238,N_35947,N_35035);
nor U38239 (N_38239,N_36304,N_36594);
xnor U38240 (N_38240,N_35178,N_35128);
nor U38241 (N_38241,N_36315,N_36862);
and U38242 (N_38242,N_36695,N_35527);
and U38243 (N_38243,N_37470,N_36329);
xnor U38244 (N_38244,N_37435,N_36465);
or U38245 (N_38245,N_37220,N_36059);
nor U38246 (N_38246,N_35941,N_37445);
xnor U38247 (N_38247,N_35079,N_35663);
nor U38248 (N_38248,N_36660,N_36477);
xnor U38249 (N_38249,N_35904,N_35166);
nor U38250 (N_38250,N_35145,N_37047);
nand U38251 (N_38251,N_36671,N_35341);
xor U38252 (N_38252,N_35494,N_35624);
nand U38253 (N_38253,N_37493,N_36123);
and U38254 (N_38254,N_36197,N_35672);
or U38255 (N_38255,N_37398,N_35645);
xnor U38256 (N_38256,N_35856,N_36003);
xnor U38257 (N_38257,N_35163,N_35020);
xnor U38258 (N_38258,N_37362,N_36869);
and U38259 (N_38259,N_36470,N_36284);
and U38260 (N_38260,N_37209,N_36166);
nor U38261 (N_38261,N_37439,N_35195);
nor U38262 (N_38262,N_36250,N_36597);
or U38263 (N_38263,N_36347,N_37139);
nand U38264 (N_38264,N_37065,N_35140);
nor U38265 (N_38265,N_35930,N_36033);
or U38266 (N_38266,N_35563,N_36723);
nand U38267 (N_38267,N_37391,N_36764);
nand U38268 (N_38268,N_35924,N_35840);
xor U38269 (N_38269,N_35812,N_36091);
or U38270 (N_38270,N_36023,N_35281);
or U38271 (N_38271,N_37122,N_35938);
or U38272 (N_38272,N_36232,N_36964);
xor U38273 (N_38273,N_35386,N_35454);
or U38274 (N_38274,N_36124,N_35282);
or U38275 (N_38275,N_35684,N_36136);
and U38276 (N_38276,N_37165,N_35337);
and U38277 (N_38277,N_35500,N_35458);
nand U38278 (N_38278,N_36321,N_35743);
and U38279 (N_38279,N_36377,N_37215);
and U38280 (N_38280,N_37169,N_36857);
and U38281 (N_38281,N_35545,N_35951);
nand U38282 (N_38282,N_37471,N_35433);
nor U38283 (N_38283,N_35887,N_36002);
xnor U38284 (N_38284,N_35156,N_37245);
or U38285 (N_38285,N_37206,N_36239);
and U38286 (N_38286,N_35842,N_37156);
xnor U38287 (N_38287,N_36243,N_37049);
and U38288 (N_38288,N_35925,N_37487);
xnor U38289 (N_38289,N_36202,N_36583);
nor U38290 (N_38290,N_36491,N_35313);
xor U38291 (N_38291,N_37408,N_35427);
or U38292 (N_38292,N_37492,N_37089);
xor U38293 (N_38293,N_35445,N_36661);
nand U38294 (N_38294,N_36395,N_35891);
nor U38295 (N_38295,N_35881,N_35763);
nand U38296 (N_38296,N_37148,N_36406);
and U38297 (N_38297,N_36639,N_36171);
and U38298 (N_38298,N_35649,N_37000);
nand U38299 (N_38299,N_36855,N_37096);
or U38300 (N_38300,N_37219,N_37388);
or U38301 (N_38301,N_35511,N_37265);
nor U38302 (N_38302,N_35193,N_36756);
nand U38303 (N_38303,N_36806,N_36283);
nor U38304 (N_38304,N_35068,N_36135);
nor U38305 (N_38305,N_35212,N_35777);
and U38306 (N_38306,N_36892,N_36251);
and U38307 (N_38307,N_35987,N_35291);
nand U38308 (N_38308,N_35473,N_36739);
or U38309 (N_38309,N_36364,N_35202);
nor U38310 (N_38310,N_36241,N_35521);
and U38311 (N_38311,N_36865,N_35324);
nor U38312 (N_38312,N_37224,N_36589);
nor U38313 (N_38313,N_37167,N_35250);
or U38314 (N_38314,N_36432,N_35312);
or U38315 (N_38315,N_35888,N_37106);
nor U38316 (N_38316,N_36017,N_36094);
nor U38317 (N_38317,N_35955,N_35430);
and U38318 (N_38318,N_36760,N_35619);
xnor U38319 (N_38319,N_35480,N_36034);
and U38320 (N_38320,N_36599,N_37348);
and U38321 (N_38321,N_36375,N_35419);
nor U38322 (N_38322,N_35586,N_37170);
nor U38323 (N_38323,N_35284,N_35710);
or U38324 (N_38324,N_35564,N_36063);
nand U38325 (N_38325,N_35086,N_37389);
nand U38326 (N_38326,N_36187,N_35996);
and U38327 (N_38327,N_37491,N_35358);
nand U38328 (N_38328,N_36361,N_37125);
xnor U38329 (N_38329,N_35131,N_35171);
or U38330 (N_38330,N_36641,N_36488);
and U38331 (N_38331,N_35857,N_36201);
xnor U38332 (N_38332,N_35486,N_36054);
and U38333 (N_38333,N_35242,N_36272);
xnor U38334 (N_38334,N_35733,N_37194);
nor U38335 (N_38335,N_35066,N_37280);
or U38336 (N_38336,N_36918,N_36006);
or U38337 (N_38337,N_35961,N_37052);
xnor U38338 (N_38338,N_36947,N_35776);
nor U38339 (N_38339,N_35201,N_36864);
nor U38340 (N_38340,N_37230,N_37160);
xor U38341 (N_38341,N_36433,N_36984);
xnor U38342 (N_38342,N_36846,N_36893);
and U38343 (N_38343,N_35360,N_35981);
nor U38344 (N_38344,N_35819,N_36027);
xnor U38345 (N_38345,N_35130,N_36195);
xnor U38346 (N_38346,N_35149,N_35986);
or U38347 (N_38347,N_36615,N_35515);
or U38348 (N_38348,N_35031,N_35689);
nand U38349 (N_38349,N_36473,N_37370);
or U38350 (N_38350,N_36914,N_37353);
nor U38351 (N_38351,N_35754,N_35053);
or U38352 (N_38352,N_35652,N_36909);
and U38353 (N_38353,N_35541,N_37173);
or U38354 (N_38354,N_35552,N_35350);
or U38355 (N_38355,N_36807,N_36122);
or U38356 (N_38356,N_35226,N_36729);
nor U38357 (N_38357,N_37367,N_37001);
nor U38358 (N_38358,N_36960,N_35406);
nor U38359 (N_38359,N_35198,N_36213);
nor U38360 (N_38360,N_35935,N_36154);
xnor U38361 (N_38361,N_36852,N_35806);
and U38362 (N_38362,N_37118,N_36835);
xnor U38363 (N_38363,N_37291,N_35761);
xnor U38364 (N_38364,N_36026,N_36435);
xnor U38365 (N_38365,N_36014,N_37281);
or U38366 (N_38366,N_35401,N_35259);
nor U38367 (N_38367,N_37246,N_35167);
nor U38368 (N_38368,N_36642,N_36561);
and U38369 (N_38369,N_35697,N_37309);
xnor U38370 (N_38370,N_37494,N_37310);
nand U38371 (N_38371,N_35899,N_36944);
xnor U38372 (N_38372,N_36386,N_35288);
and U38373 (N_38373,N_37025,N_35786);
nor U38374 (N_38374,N_35455,N_36775);
and U38375 (N_38375,N_36442,N_36029);
nand U38376 (N_38376,N_35187,N_35818);
xor U38377 (N_38377,N_36472,N_35394);
nor U38378 (N_38378,N_36429,N_35420);
nand U38379 (N_38379,N_36747,N_37250);
and U38380 (N_38380,N_35702,N_35994);
nand U38381 (N_38381,N_36415,N_35330);
xnor U38382 (N_38382,N_37031,N_36779);
nand U38383 (N_38383,N_37490,N_35346);
nor U38384 (N_38384,N_35505,N_36628);
nor U38385 (N_38385,N_37023,N_36751);
nor U38386 (N_38386,N_35475,N_36233);
or U38387 (N_38387,N_35713,N_37258);
nor U38388 (N_38388,N_36076,N_36448);
or U38389 (N_38389,N_36592,N_35331);
nand U38390 (N_38390,N_36000,N_36528);
or U38391 (N_38391,N_35310,N_36170);
nand U38392 (N_38392,N_36537,N_37138);
xor U38393 (N_38393,N_35405,N_35172);
and U38394 (N_38394,N_36754,N_36414);
nor U38395 (N_38395,N_36380,N_35449);
nand U38396 (N_38396,N_35509,N_35657);
xnor U38397 (N_38397,N_35115,N_36343);
or U38398 (N_38398,N_35390,N_35698);
nor U38399 (N_38399,N_36460,N_37316);
nor U38400 (N_38400,N_35348,N_36789);
nor U38401 (N_38401,N_36115,N_36899);
nor U38402 (N_38402,N_37144,N_37093);
and U38403 (N_38403,N_36702,N_35907);
nand U38404 (N_38404,N_35911,N_35429);
and U38405 (N_38405,N_36287,N_36450);
xnor U38406 (N_38406,N_37312,N_36750);
and U38407 (N_38407,N_35978,N_36619);
or U38408 (N_38408,N_35355,N_36373);
xor U38409 (N_38409,N_36826,N_37081);
or U38410 (N_38410,N_35122,N_35200);
nand U38411 (N_38411,N_35083,N_37168);
or U38412 (N_38412,N_37012,N_35822);
nand U38413 (N_38413,N_35229,N_35421);
xor U38414 (N_38414,N_36508,N_35081);
or U38415 (N_38415,N_35900,N_35578);
and U38416 (N_38416,N_36938,N_37127);
or U38417 (N_38417,N_37498,N_35225);
and U38418 (N_38418,N_36991,N_35529);
nor U38419 (N_38419,N_36082,N_36822);
xnor U38420 (N_38420,N_35048,N_37289);
or U38421 (N_38421,N_35946,N_37301);
and U38422 (N_38422,N_37166,N_36680);
nor U38423 (N_38423,N_36881,N_35694);
and U38424 (N_38424,N_37135,N_35845);
nand U38425 (N_38425,N_36184,N_36603);
nand U38426 (N_38426,N_36688,N_35678);
and U38427 (N_38427,N_37044,N_36264);
nor U38428 (N_38428,N_36937,N_36164);
nand U38429 (N_38429,N_36708,N_36120);
or U38430 (N_38430,N_36019,N_36569);
and U38431 (N_38431,N_35655,N_37283);
or U38432 (N_38432,N_35453,N_35779);
xnor U38433 (N_38433,N_36226,N_36240);
xnor U38434 (N_38434,N_37120,N_35797);
or U38435 (N_38435,N_37332,N_36971);
nor U38436 (N_38436,N_36088,N_36466);
nor U38437 (N_38437,N_37251,N_35261);
or U38438 (N_38438,N_36649,N_37041);
or U38439 (N_38439,N_36262,N_35960);
or U38440 (N_38440,N_36725,N_35860);
or U38441 (N_38441,N_36056,N_35227);
nand U38442 (N_38442,N_36077,N_35008);
nand U38443 (N_38443,N_36355,N_36890);
or U38444 (N_38444,N_36746,N_35286);
nor U38445 (N_38445,N_35317,N_35623);
or U38446 (N_38446,N_35612,N_36633);
or U38447 (N_38447,N_37157,N_35471);
and U38448 (N_38448,N_35640,N_35989);
and U38449 (N_38449,N_35726,N_37128);
nor U38450 (N_38450,N_35047,N_37423);
xnor U38451 (N_38451,N_35400,N_35221);
or U38452 (N_38452,N_36486,N_35626);
xor U38453 (N_38453,N_36216,N_36322);
nand U38454 (N_38454,N_37356,N_35161);
nor U38455 (N_38455,N_35465,N_36917);
xor U38456 (N_38456,N_35007,N_36953);
and U38457 (N_38457,N_35696,N_35628);
xnor U38458 (N_38458,N_37285,N_36392);
xor U38459 (N_38459,N_35943,N_35990);
nand U38460 (N_38460,N_36394,N_36799);
nor U38461 (N_38461,N_37094,N_35917);
and U38462 (N_38462,N_35434,N_35815);
nand U38463 (N_38463,N_36715,N_37225);
and U38464 (N_38464,N_36285,N_36945);
and U38465 (N_38465,N_36198,N_36978);
and U38466 (N_38466,N_36635,N_36068);
or U38467 (N_38467,N_35165,N_37368);
nor U38468 (N_38468,N_36391,N_35875);
xor U38469 (N_38469,N_36605,N_35601);
and U38470 (N_38470,N_35342,N_37131);
or U38471 (N_38471,N_36103,N_36711);
nand U38472 (N_38472,N_36905,N_35603);
or U38473 (N_38473,N_37410,N_37005);
or U38474 (N_38474,N_36109,N_36009);
xnor U38475 (N_38475,N_35850,N_35675);
xor U38476 (N_38476,N_37382,N_35459);
xnor U38477 (N_38477,N_35972,N_36190);
xor U38478 (N_38478,N_36158,N_35345);
xor U38479 (N_38479,N_35307,N_36362);
or U38480 (N_38480,N_36951,N_37107);
xnor U38481 (N_38481,N_35602,N_36872);
or U38482 (N_38482,N_37481,N_36692);
or U38483 (N_38483,N_36010,N_36214);
nor U38484 (N_38484,N_37063,N_35155);
nand U38485 (N_38485,N_35799,N_37185);
nand U38486 (N_38486,N_35864,N_36962);
or U38487 (N_38487,N_35727,N_36269);
or U38488 (N_38488,N_35460,N_35309);
xnor U38489 (N_38489,N_36446,N_36047);
nand U38490 (N_38490,N_36183,N_37149);
xor U38491 (N_38491,N_36040,N_36906);
and U38492 (N_38492,N_36724,N_36393);
nor U38493 (N_38493,N_36365,N_35789);
or U38494 (N_38494,N_37188,N_36560);
nor U38495 (N_38495,N_36503,N_35142);
nor U38496 (N_38496,N_37288,N_36405);
xnor U38497 (N_38497,N_35021,N_37433);
xnor U38498 (N_38498,N_36810,N_35933);
or U38499 (N_38499,N_36471,N_36759);
xor U38500 (N_38500,N_35299,N_35544);
nor U38501 (N_38501,N_35764,N_36933);
and U38502 (N_38502,N_35011,N_37010);
or U38503 (N_38503,N_37495,N_36499);
nand U38504 (N_38504,N_35660,N_35895);
and U38505 (N_38505,N_36193,N_35275);
and U38506 (N_38506,N_36225,N_35308);
nor U38507 (N_38507,N_36825,N_36525);
xnor U38508 (N_38508,N_35208,N_36338);
nand U38509 (N_38509,N_35158,N_37113);
nor U38510 (N_38510,N_36215,N_36601);
or U38511 (N_38511,N_36132,N_37333);
or U38512 (N_38512,N_36080,N_35720);
and U38513 (N_38513,N_35591,N_35774);
and U38514 (N_38514,N_35963,N_37037);
nor U38515 (N_38515,N_37390,N_35752);
xor U38516 (N_38516,N_37029,N_35032);
nand U38517 (N_38517,N_35825,N_35594);
or U38518 (N_38518,N_37018,N_37198);
nand U38519 (N_38519,N_37275,N_35889);
or U38520 (N_38520,N_36510,N_36311);
or U38521 (N_38521,N_35160,N_36177);
and U38522 (N_38522,N_36675,N_35297);
nand U38523 (N_38523,N_36687,N_37137);
and U38524 (N_38524,N_35643,N_35210);
and U38525 (N_38525,N_35249,N_36496);
xnor U38526 (N_38526,N_37450,N_36884);
and U38527 (N_38527,N_35559,N_36188);
or U38528 (N_38528,N_35539,N_35409);
or U38529 (N_38529,N_36580,N_35787);
nor U38530 (N_38530,N_35921,N_36427);
nand U38531 (N_38531,N_36237,N_36001);
nand U38532 (N_38532,N_36445,N_35061);
or U38533 (N_38533,N_35611,N_37043);
nor U38534 (N_38534,N_35228,N_35090);
and U38535 (N_38535,N_36837,N_36763);
xor U38536 (N_38536,N_35673,N_35347);
xor U38537 (N_38537,N_37300,N_35169);
xor U38538 (N_38538,N_35410,N_35478);
nand U38539 (N_38539,N_35985,N_35755);
xor U38540 (N_38540,N_37091,N_36256);
nor U38541 (N_38541,N_37150,N_35919);
nor U38542 (N_38542,N_36305,N_36590);
xor U38543 (N_38543,N_37199,N_36956);
xnor U38544 (N_38544,N_36342,N_37123);
and U38545 (N_38545,N_36957,N_36919);
or U38546 (N_38546,N_35343,N_35077);
nand U38547 (N_38547,N_36500,N_37404);
xor U38548 (N_38548,N_35137,N_35423);
nand U38549 (N_38549,N_36266,N_35089);
nand U38550 (N_38550,N_37419,N_35026);
nor U38551 (N_38551,N_37416,N_37272);
and U38552 (N_38552,N_37432,N_36663);
and U38553 (N_38553,N_37438,N_35877);
nand U38554 (N_38554,N_36786,N_37038);
xor U38555 (N_38555,N_36336,N_35558);
or U38556 (N_38556,N_36911,N_37032);
or U38557 (N_38557,N_35884,N_36614);
or U38558 (N_38558,N_36146,N_36901);
or U38559 (N_38559,N_35677,N_35773);
and U38560 (N_38560,N_35320,N_35485);
nor U38561 (N_38561,N_36160,N_35561);
nand U38562 (N_38562,N_35450,N_36931);
or U38563 (N_38563,N_36236,N_35615);
nand U38564 (N_38564,N_35039,N_35129);
xor U38565 (N_38565,N_36521,N_35741);
or U38566 (N_38566,N_36785,N_37412);
xnor U38567 (N_38567,N_35821,N_36691);
or U38568 (N_38568,N_37003,N_36625);
xor U38569 (N_38569,N_37336,N_35533);
xor U38570 (N_38570,N_36016,N_36727);
xor U38571 (N_38571,N_36079,N_35798);
and U38572 (N_38572,N_37191,N_36469);
or U38573 (N_38573,N_37371,N_36611);
nor U38574 (N_38574,N_36403,N_36908);
nor U38575 (N_38575,N_36199,N_37358);
or U38576 (N_38576,N_36143,N_35316);
or U38577 (N_38577,N_37417,N_36174);
nor U38578 (N_38578,N_37363,N_37483);
or U38579 (N_38579,N_35267,N_35280);
nand U38580 (N_38580,N_37073,N_37243);
nor U38581 (N_38581,N_35222,N_36345);
nand U38582 (N_38582,N_36620,N_36926);
xnor U38583 (N_38583,N_35438,N_36930);
and U38584 (N_38584,N_35327,N_35852);
and U38585 (N_38585,N_36975,N_35828);
and U38586 (N_38586,N_36113,N_35144);
xnor U38587 (N_38587,N_37365,N_35151);
xor U38588 (N_38588,N_36769,N_35107);
and U38589 (N_38589,N_36401,N_35236);
and U38590 (N_38590,N_36952,N_35897);
xnor U38591 (N_38591,N_36370,N_36885);
and U38592 (N_38592,N_35265,N_36958);
xor U38593 (N_38593,N_36180,N_35388);
xnor U38594 (N_38594,N_35328,N_35585);
nand U38595 (N_38595,N_36784,N_35557);
or U38596 (N_38596,N_36648,N_35211);
nor U38597 (N_38597,N_36402,N_36155);
or U38598 (N_38598,N_35576,N_37061);
nand U38599 (N_38599,N_37129,N_37317);
or U38600 (N_38600,N_35824,N_35793);
nor U38601 (N_38601,N_36859,N_36842);
nor U38602 (N_38602,N_35659,N_37341);
nor U38603 (N_38603,N_37014,N_37193);
or U38604 (N_38604,N_37422,N_36220);
and U38605 (N_38605,N_35258,N_37468);
and U38606 (N_38606,N_35076,N_37066);
and U38607 (N_38607,N_37158,N_36453);
nand U38608 (N_38608,N_36621,N_35036);
or U38609 (N_38609,N_36968,N_37080);
nor U38610 (N_38610,N_36943,N_37030);
xnor U38611 (N_38611,N_36969,N_36586);
or U38612 (N_38612,N_36292,N_36359);
xnor U38613 (N_38613,N_36316,N_37306);
or U38614 (N_38614,N_35446,N_36883);
or U38615 (N_38615,N_35858,N_36547);
xnor U38616 (N_38616,N_35991,N_37054);
xnor U38617 (N_38617,N_35017,N_36203);
nand U38618 (N_38618,N_35738,N_36923);
nor U38619 (N_38619,N_35523,N_36545);
and U38620 (N_38620,N_36888,N_35477);
and U38621 (N_38621,N_37101,N_35553);
or U38622 (N_38622,N_36046,N_36704);
or U38623 (N_38623,N_36478,N_36065);
xor U38624 (N_38624,N_36137,N_36344);
nand U38625 (N_38625,N_35901,N_35370);
xnor U38626 (N_38626,N_36816,N_37431);
nor U38627 (N_38627,N_36461,N_35353);
nand U38628 (N_38628,N_35876,N_36101);
nor U38629 (N_38629,N_37452,N_35795);
nor U38630 (N_38630,N_36809,N_36032);
xor U38631 (N_38631,N_35103,N_36988);
and U38632 (N_38632,N_36595,N_35016);
nor U38633 (N_38633,N_37425,N_37074);
and U38634 (N_38634,N_37384,N_37430);
nand U38635 (N_38635,N_35906,N_36553);
and U38636 (N_38636,N_35045,N_36245);
xnor U38637 (N_38637,N_36877,N_36967);
nand U38638 (N_38638,N_36564,N_36259);
or U38639 (N_38639,N_35027,N_36005);
and U38640 (N_38640,N_35441,N_35489);
and U38641 (N_38641,N_37482,N_37292);
or U38642 (N_38642,N_36325,N_36072);
and U38643 (N_38643,N_37400,N_35855);
nor U38644 (N_38644,N_35736,N_37379);
nor U38645 (N_38645,N_35097,N_37136);
or U38646 (N_38646,N_35038,N_35120);
or U38647 (N_38647,N_35937,N_35631);
nand U38648 (N_38648,N_36772,N_36464);
or U38649 (N_38649,N_36794,N_35832);
nand U38650 (N_38650,N_36368,N_36961);
nand U38651 (N_38651,N_36948,N_36413);
or U38652 (N_38652,N_35598,N_37303);
and U38653 (N_38653,N_37033,N_36606);
and U38654 (N_38654,N_36841,N_36831);
and U38655 (N_38655,N_36024,N_37196);
xor U38656 (N_38656,N_37084,N_37499);
or U38657 (N_38657,N_36707,N_36850);
and U38658 (N_38658,N_36790,N_37489);
nor U38659 (N_38659,N_35399,N_36051);
or U38660 (N_38660,N_35600,N_35785);
xnor U38661 (N_38661,N_37293,N_37212);
and U38662 (N_38662,N_35867,N_36501);
nor U38663 (N_38663,N_37070,N_35233);
or U38664 (N_38664,N_36212,N_37134);
and U38665 (N_38665,N_37392,N_36385);
and U38666 (N_38666,N_36980,N_35639);
or U38667 (N_38667,N_35184,N_37472);
nor U38668 (N_38668,N_36509,N_36238);
nor U38669 (N_38669,N_37121,N_37409);
nor U38670 (N_38670,N_36354,N_35550);
nand U38671 (N_38671,N_35597,N_35679);
or U38672 (N_38672,N_35725,N_37140);
or U38673 (N_38673,N_36840,N_36863);
nor U38674 (N_38674,N_36679,N_36833);
and U38675 (N_38675,N_35965,N_36084);
nand U38676 (N_38676,N_35633,N_35531);
and U38677 (N_38677,N_35874,N_36936);
nand U38678 (N_38678,N_35418,N_37237);
nor U38679 (N_38679,N_36161,N_36289);
or U38680 (N_38680,N_36490,N_37461);
nor U38681 (N_38681,N_36367,N_36674);
xnor U38682 (N_38682,N_35766,N_36157);
xnor U38683 (N_38683,N_35682,N_35179);
and U38684 (N_38684,N_35962,N_36261);
and U38685 (N_38685,N_35959,N_37426);
or U38686 (N_38686,N_35082,N_35668);
or U38687 (N_38687,N_35033,N_35274);
or U38688 (N_38688,N_35051,N_37211);
and U38689 (N_38689,N_35028,N_36376);
nand U38690 (N_38690,N_35180,N_37147);
xnor U38691 (N_38691,N_37177,N_37174);
nor U38692 (N_38692,N_36929,N_36669);
nand U38693 (N_38693,N_36308,N_36973);
or U38694 (N_38694,N_35627,N_35641);
nor U38695 (N_38695,N_36685,N_35687);
xnor U38696 (N_38696,N_35607,N_35064);
or U38697 (N_38697,N_37132,N_36555);
nor U38698 (N_38698,N_37411,N_36666);
nor U38699 (N_38699,N_35121,N_36223);
or U38700 (N_38700,N_36854,N_35205);
nor U38701 (N_38701,N_35686,N_37036);
and U38702 (N_38702,N_36069,N_35230);
xor U38703 (N_38703,N_35080,N_36371);
xor U38704 (N_38704,N_35551,N_35507);
nor U38705 (N_38705,N_35693,N_35952);
and U38706 (N_38706,N_35648,N_36741);
and U38707 (N_38707,N_35436,N_36697);
nand U38708 (N_38708,N_37413,N_35548);
nand U38709 (N_38709,N_35514,N_37318);
or U38710 (N_38710,N_35723,N_36093);
and U38711 (N_38711,N_36159,N_36522);
or U38712 (N_38712,N_36640,N_35417);
nand U38713 (N_38713,N_35174,N_36728);
nand U38714 (N_38714,N_36015,N_36048);
xor U38715 (N_38715,N_37253,N_37087);
xor U38716 (N_38716,N_36802,N_35329);
xor U38717 (N_38717,N_36467,N_37153);
nand U38718 (N_38718,N_37027,N_37351);
and U38719 (N_38719,N_36444,N_36740);
nand U38720 (N_38720,N_37075,N_35547);
nand U38721 (N_38721,N_37068,N_36714);
nand U38722 (N_38722,N_37116,N_36643);
xnor U38723 (N_38723,N_37387,N_36734);
nand U38724 (N_38724,N_35217,N_35183);
xor U38725 (N_38725,N_36535,N_36493);
or U38726 (N_38726,N_37015,N_35695);
nand U38727 (N_38727,N_35613,N_36871);
and U38728 (N_38728,N_37102,N_35371);
xnor U38729 (N_38729,N_35009,N_36067);
and U38730 (N_38730,N_36631,N_35912);
nand U38731 (N_38731,N_35588,N_36618);
or U38732 (N_38732,N_36057,N_35705);
or U38733 (N_38733,N_35814,N_37098);
xnor U38734 (N_38734,N_36276,N_37484);
nand U38735 (N_38735,N_36903,N_35730);
nand U38736 (N_38736,N_36656,N_35214);
xnor U38737 (N_38737,N_35363,N_36778);
nor U38738 (N_38738,N_36847,N_37443);
nand U38739 (N_38739,N_36773,N_35413);
nand U38740 (N_38740,N_35791,N_36626);
nand U38741 (N_38741,N_35953,N_35432);
or U38742 (N_38742,N_36443,N_35403);
and U38743 (N_38743,N_35085,N_36277);
xor U38744 (N_38744,N_36647,N_35984);
and U38745 (N_38745,N_35244,N_36208);
xnor U38746 (N_38746,N_36335,N_35101);
and U38747 (N_38747,N_36323,N_37340);
nand U38748 (N_38748,N_35903,N_37217);
nand U38749 (N_38749,N_36800,N_37441);
nor U38750 (N_38750,N_36290,N_35211);
or U38751 (N_38751,N_36011,N_36614);
or U38752 (N_38752,N_36628,N_36880);
or U38753 (N_38753,N_35410,N_36611);
or U38754 (N_38754,N_36301,N_36145);
nor U38755 (N_38755,N_37367,N_35002);
nor U38756 (N_38756,N_37497,N_37287);
or U38757 (N_38757,N_35011,N_35119);
xor U38758 (N_38758,N_35504,N_36989);
and U38759 (N_38759,N_36043,N_37441);
nand U38760 (N_38760,N_35418,N_36387);
xor U38761 (N_38761,N_35598,N_35591);
nand U38762 (N_38762,N_35449,N_35901);
nor U38763 (N_38763,N_37098,N_35826);
or U38764 (N_38764,N_35522,N_36398);
xor U38765 (N_38765,N_37249,N_36891);
and U38766 (N_38766,N_35143,N_36521);
nand U38767 (N_38767,N_37189,N_35610);
and U38768 (N_38768,N_37071,N_36491);
and U38769 (N_38769,N_36038,N_36480);
xnor U38770 (N_38770,N_36995,N_36652);
nand U38771 (N_38771,N_36632,N_36687);
and U38772 (N_38772,N_36918,N_35364);
nor U38773 (N_38773,N_37173,N_36814);
nand U38774 (N_38774,N_37295,N_36427);
nor U38775 (N_38775,N_36727,N_36988);
xnor U38776 (N_38776,N_35642,N_35717);
or U38777 (N_38777,N_36916,N_37045);
nor U38778 (N_38778,N_36922,N_35077);
or U38779 (N_38779,N_36717,N_36916);
nor U38780 (N_38780,N_36330,N_35661);
nor U38781 (N_38781,N_35257,N_35794);
nand U38782 (N_38782,N_37127,N_36205);
xnor U38783 (N_38783,N_37448,N_36904);
xnor U38784 (N_38784,N_35786,N_35868);
xnor U38785 (N_38785,N_36306,N_35559);
nand U38786 (N_38786,N_36812,N_37161);
and U38787 (N_38787,N_35437,N_37364);
and U38788 (N_38788,N_36828,N_36941);
or U38789 (N_38789,N_36258,N_35322);
nor U38790 (N_38790,N_36710,N_36672);
xor U38791 (N_38791,N_35809,N_35131);
xor U38792 (N_38792,N_35276,N_35675);
xnor U38793 (N_38793,N_36852,N_35421);
xor U38794 (N_38794,N_35639,N_36510);
nor U38795 (N_38795,N_36107,N_36655);
nor U38796 (N_38796,N_37240,N_37216);
nor U38797 (N_38797,N_35108,N_36882);
nor U38798 (N_38798,N_37039,N_36131);
nor U38799 (N_38799,N_35020,N_35915);
nor U38800 (N_38800,N_37287,N_37223);
xor U38801 (N_38801,N_37077,N_36934);
nor U38802 (N_38802,N_37194,N_37453);
nor U38803 (N_38803,N_36973,N_35850);
and U38804 (N_38804,N_37343,N_36086);
nand U38805 (N_38805,N_37028,N_36826);
nor U38806 (N_38806,N_35241,N_35977);
xnor U38807 (N_38807,N_36955,N_37070);
and U38808 (N_38808,N_36350,N_35110);
and U38809 (N_38809,N_37475,N_36613);
nor U38810 (N_38810,N_35843,N_36237);
and U38811 (N_38811,N_36432,N_36107);
or U38812 (N_38812,N_36727,N_35273);
xnor U38813 (N_38813,N_35320,N_35835);
or U38814 (N_38814,N_36756,N_37348);
or U38815 (N_38815,N_37497,N_35984);
or U38816 (N_38816,N_36429,N_36979);
and U38817 (N_38817,N_36617,N_35600);
or U38818 (N_38818,N_36633,N_36537);
and U38819 (N_38819,N_35912,N_36896);
nand U38820 (N_38820,N_36935,N_35770);
nor U38821 (N_38821,N_36715,N_37467);
nor U38822 (N_38822,N_37486,N_35932);
or U38823 (N_38823,N_36206,N_35433);
nand U38824 (N_38824,N_36418,N_37131);
nand U38825 (N_38825,N_37324,N_36495);
and U38826 (N_38826,N_37291,N_37134);
and U38827 (N_38827,N_37449,N_35998);
nand U38828 (N_38828,N_35868,N_35564);
xnor U38829 (N_38829,N_36331,N_35997);
nand U38830 (N_38830,N_37426,N_36601);
nor U38831 (N_38831,N_36903,N_37088);
or U38832 (N_38832,N_35427,N_37167);
nor U38833 (N_38833,N_37052,N_35984);
or U38834 (N_38834,N_36114,N_37222);
xnor U38835 (N_38835,N_35683,N_36615);
nand U38836 (N_38836,N_36716,N_36361);
nand U38837 (N_38837,N_36417,N_35939);
nand U38838 (N_38838,N_35675,N_35888);
nand U38839 (N_38839,N_35096,N_35024);
xnor U38840 (N_38840,N_35523,N_36968);
and U38841 (N_38841,N_36968,N_37010);
nand U38842 (N_38842,N_35636,N_35980);
nor U38843 (N_38843,N_35341,N_35325);
xor U38844 (N_38844,N_37247,N_36021);
xnor U38845 (N_38845,N_36336,N_35035);
and U38846 (N_38846,N_37346,N_37106);
or U38847 (N_38847,N_37009,N_36623);
nor U38848 (N_38848,N_35553,N_35205);
nor U38849 (N_38849,N_35671,N_35757);
nand U38850 (N_38850,N_36274,N_35647);
xnor U38851 (N_38851,N_36666,N_36733);
and U38852 (N_38852,N_35228,N_36306);
xor U38853 (N_38853,N_36158,N_36033);
nor U38854 (N_38854,N_36080,N_36367);
xor U38855 (N_38855,N_37432,N_35254);
and U38856 (N_38856,N_36686,N_37177);
nand U38857 (N_38857,N_36200,N_35112);
xor U38858 (N_38858,N_37328,N_35915);
nor U38859 (N_38859,N_37140,N_35388);
nor U38860 (N_38860,N_35760,N_35336);
nand U38861 (N_38861,N_35399,N_35371);
or U38862 (N_38862,N_36867,N_37149);
and U38863 (N_38863,N_36326,N_35381);
and U38864 (N_38864,N_37242,N_37220);
or U38865 (N_38865,N_35728,N_35364);
nor U38866 (N_38866,N_36131,N_36455);
nand U38867 (N_38867,N_35709,N_36171);
xor U38868 (N_38868,N_35720,N_36609);
nand U38869 (N_38869,N_35902,N_35844);
nand U38870 (N_38870,N_36480,N_35518);
and U38871 (N_38871,N_37114,N_35855);
nor U38872 (N_38872,N_36346,N_36881);
and U38873 (N_38873,N_35256,N_36283);
nor U38874 (N_38874,N_35552,N_35499);
and U38875 (N_38875,N_36621,N_35863);
or U38876 (N_38876,N_35930,N_36582);
and U38877 (N_38877,N_36056,N_36799);
and U38878 (N_38878,N_35325,N_37418);
or U38879 (N_38879,N_35252,N_35451);
or U38880 (N_38880,N_35326,N_35414);
or U38881 (N_38881,N_37412,N_36019);
nand U38882 (N_38882,N_37234,N_36220);
or U38883 (N_38883,N_35827,N_36347);
nor U38884 (N_38884,N_36983,N_35415);
and U38885 (N_38885,N_35975,N_36989);
and U38886 (N_38886,N_37465,N_35697);
nand U38887 (N_38887,N_35087,N_36915);
nand U38888 (N_38888,N_35773,N_36411);
nand U38889 (N_38889,N_36607,N_35045);
xnor U38890 (N_38890,N_35862,N_36464);
and U38891 (N_38891,N_36933,N_37396);
nand U38892 (N_38892,N_36275,N_35227);
nor U38893 (N_38893,N_37379,N_36834);
or U38894 (N_38894,N_35863,N_37063);
and U38895 (N_38895,N_35323,N_35819);
or U38896 (N_38896,N_36854,N_36024);
nand U38897 (N_38897,N_35294,N_35776);
nand U38898 (N_38898,N_35584,N_36329);
xnor U38899 (N_38899,N_36176,N_37027);
nand U38900 (N_38900,N_37285,N_35443);
nand U38901 (N_38901,N_36682,N_35212);
nor U38902 (N_38902,N_35598,N_35458);
xor U38903 (N_38903,N_35253,N_35271);
xnor U38904 (N_38904,N_35173,N_36273);
or U38905 (N_38905,N_36249,N_36157);
nor U38906 (N_38906,N_35076,N_36188);
nand U38907 (N_38907,N_36046,N_37103);
nor U38908 (N_38908,N_35847,N_36463);
and U38909 (N_38909,N_36449,N_35650);
nand U38910 (N_38910,N_36779,N_37283);
nor U38911 (N_38911,N_35380,N_36835);
xor U38912 (N_38912,N_35058,N_35679);
nor U38913 (N_38913,N_35396,N_36766);
xnor U38914 (N_38914,N_35562,N_36339);
nand U38915 (N_38915,N_35972,N_37063);
nor U38916 (N_38916,N_36756,N_35631);
or U38917 (N_38917,N_36246,N_37250);
nor U38918 (N_38918,N_35067,N_35116);
or U38919 (N_38919,N_35613,N_36647);
and U38920 (N_38920,N_37090,N_36482);
nand U38921 (N_38921,N_35647,N_36915);
xor U38922 (N_38922,N_35599,N_35822);
nor U38923 (N_38923,N_37036,N_36734);
nand U38924 (N_38924,N_37137,N_35460);
nor U38925 (N_38925,N_35872,N_36040);
or U38926 (N_38926,N_36831,N_35722);
and U38927 (N_38927,N_35011,N_36803);
and U38928 (N_38928,N_35463,N_37430);
and U38929 (N_38929,N_36786,N_36393);
or U38930 (N_38930,N_36887,N_37068);
xnor U38931 (N_38931,N_35573,N_35475);
and U38932 (N_38932,N_36609,N_36992);
nor U38933 (N_38933,N_36641,N_36635);
or U38934 (N_38934,N_36747,N_36149);
nor U38935 (N_38935,N_35877,N_35586);
nor U38936 (N_38936,N_36554,N_35439);
nor U38937 (N_38937,N_35845,N_36212);
or U38938 (N_38938,N_36959,N_35113);
xor U38939 (N_38939,N_36274,N_36629);
nand U38940 (N_38940,N_36233,N_35818);
or U38941 (N_38941,N_36805,N_36939);
xor U38942 (N_38942,N_37200,N_35482);
nor U38943 (N_38943,N_36024,N_36611);
xor U38944 (N_38944,N_37342,N_35448);
nor U38945 (N_38945,N_37204,N_36583);
nor U38946 (N_38946,N_37052,N_36575);
nor U38947 (N_38947,N_35487,N_35511);
xnor U38948 (N_38948,N_35007,N_36853);
nand U38949 (N_38949,N_36623,N_37170);
xnor U38950 (N_38950,N_36210,N_36919);
or U38951 (N_38951,N_36298,N_36999);
nand U38952 (N_38952,N_36563,N_37483);
or U38953 (N_38953,N_36864,N_36573);
xnor U38954 (N_38954,N_35287,N_36076);
and U38955 (N_38955,N_36048,N_35026);
xnor U38956 (N_38956,N_36336,N_37008);
and U38957 (N_38957,N_36243,N_36556);
xnor U38958 (N_38958,N_35032,N_37491);
nor U38959 (N_38959,N_35792,N_35140);
and U38960 (N_38960,N_35619,N_37398);
nand U38961 (N_38961,N_35222,N_36301);
and U38962 (N_38962,N_36951,N_35356);
nand U38963 (N_38963,N_35228,N_36527);
or U38964 (N_38964,N_36373,N_35940);
or U38965 (N_38965,N_36158,N_35030);
xor U38966 (N_38966,N_37160,N_37213);
and U38967 (N_38967,N_35597,N_35428);
and U38968 (N_38968,N_35983,N_35620);
nor U38969 (N_38969,N_36211,N_37098);
nor U38970 (N_38970,N_37091,N_36572);
nand U38971 (N_38971,N_37490,N_36264);
or U38972 (N_38972,N_37282,N_36681);
xnor U38973 (N_38973,N_37349,N_37384);
nand U38974 (N_38974,N_36319,N_36831);
nor U38975 (N_38975,N_35755,N_37110);
xor U38976 (N_38976,N_36088,N_36123);
xor U38977 (N_38977,N_36232,N_36389);
nand U38978 (N_38978,N_35073,N_36008);
and U38979 (N_38979,N_37370,N_35565);
xnor U38980 (N_38980,N_36022,N_35001);
or U38981 (N_38981,N_35852,N_35262);
and U38982 (N_38982,N_35845,N_35677);
or U38983 (N_38983,N_35222,N_36821);
nor U38984 (N_38984,N_36620,N_35148);
nand U38985 (N_38985,N_37126,N_36183);
and U38986 (N_38986,N_36827,N_36628);
nand U38987 (N_38987,N_36809,N_35392);
nand U38988 (N_38988,N_35852,N_36415);
and U38989 (N_38989,N_35099,N_35974);
nor U38990 (N_38990,N_36081,N_37207);
and U38991 (N_38991,N_35235,N_37054);
nor U38992 (N_38992,N_35199,N_35821);
or U38993 (N_38993,N_36205,N_35940);
xnor U38994 (N_38994,N_35488,N_35111);
nand U38995 (N_38995,N_37246,N_35380);
xor U38996 (N_38996,N_37295,N_37215);
nor U38997 (N_38997,N_36596,N_35380);
or U38998 (N_38998,N_35397,N_37289);
nand U38999 (N_38999,N_35747,N_35085);
nor U39000 (N_39000,N_35422,N_37245);
or U39001 (N_39001,N_36366,N_35098);
and U39002 (N_39002,N_35390,N_36259);
or U39003 (N_39003,N_35175,N_37082);
nor U39004 (N_39004,N_35477,N_36587);
xor U39005 (N_39005,N_36740,N_35039);
nand U39006 (N_39006,N_35302,N_36830);
nand U39007 (N_39007,N_35511,N_36680);
xnor U39008 (N_39008,N_36035,N_36133);
or U39009 (N_39009,N_35534,N_37487);
xor U39010 (N_39010,N_36060,N_36798);
nand U39011 (N_39011,N_37209,N_35441);
and U39012 (N_39012,N_36371,N_35464);
nand U39013 (N_39013,N_37391,N_35224);
nand U39014 (N_39014,N_35323,N_35598);
or U39015 (N_39015,N_35605,N_36380);
nand U39016 (N_39016,N_35543,N_36426);
nor U39017 (N_39017,N_36028,N_36436);
nand U39018 (N_39018,N_36474,N_36991);
nor U39019 (N_39019,N_35713,N_35942);
and U39020 (N_39020,N_37355,N_35308);
nand U39021 (N_39021,N_36334,N_36565);
nand U39022 (N_39022,N_35049,N_37340);
nand U39023 (N_39023,N_35546,N_35069);
nand U39024 (N_39024,N_37470,N_35186);
xor U39025 (N_39025,N_37001,N_36165);
xor U39026 (N_39026,N_36664,N_36259);
xnor U39027 (N_39027,N_36719,N_36069);
xnor U39028 (N_39028,N_36979,N_35471);
and U39029 (N_39029,N_36443,N_36837);
and U39030 (N_39030,N_36199,N_35730);
and U39031 (N_39031,N_35331,N_35314);
and U39032 (N_39032,N_36565,N_35667);
xnor U39033 (N_39033,N_35169,N_36029);
nand U39034 (N_39034,N_36553,N_37083);
xor U39035 (N_39035,N_36678,N_36684);
and U39036 (N_39036,N_35727,N_35147);
nor U39037 (N_39037,N_35289,N_36580);
xor U39038 (N_39038,N_37289,N_37179);
nand U39039 (N_39039,N_35356,N_35874);
or U39040 (N_39040,N_37276,N_35453);
xor U39041 (N_39041,N_35426,N_35254);
nor U39042 (N_39042,N_36985,N_36480);
and U39043 (N_39043,N_35422,N_35753);
and U39044 (N_39044,N_35904,N_36015);
nand U39045 (N_39045,N_36887,N_35272);
xor U39046 (N_39046,N_36327,N_35663);
nor U39047 (N_39047,N_35147,N_35456);
or U39048 (N_39048,N_35895,N_36538);
nor U39049 (N_39049,N_35917,N_35995);
xor U39050 (N_39050,N_35609,N_37456);
nor U39051 (N_39051,N_36489,N_37056);
and U39052 (N_39052,N_36881,N_35851);
and U39053 (N_39053,N_36980,N_37116);
nor U39054 (N_39054,N_36091,N_35249);
xor U39055 (N_39055,N_36320,N_37158);
nor U39056 (N_39056,N_35097,N_35434);
or U39057 (N_39057,N_37034,N_37245);
nand U39058 (N_39058,N_36478,N_36727);
or U39059 (N_39059,N_36261,N_36430);
and U39060 (N_39060,N_36755,N_36731);
xnor U39061 (N_39061,N_36960,N_35349);
and U39062 (N_39062,N_37378,N_36195);
xnor U39063 (N_39063,N_35033,N_36038);
and U39064 (N_39064,N_35541,N_35515);
nand U39065 (N_39065,N_36365,N_35608);
or U39066 (N_39066,N_35408,N_36098);
and U39067 (N_39067,N_36668,N_35594);
and U39068 (N_39068,N_36992,N_35720);
nor U39069 (N_39069,N_35492,N_36138);
xor U39070 (N_39070,N_36884,N_35505);
or U39071 (N_39071,N_36562,N_35612);
xor U39072 (N_39072,N_35850,N_37094);
nor U39073 (N_39073,N_35169,N_36221);
nand U39074 (N_39074,N_37018,N_36830);
or U39075 (N_39075,N_36700,N_35568);
and U39076 (N_39076,N_37337,N_36663);
nand U39077 (N_39077,N_37154,N_35157);
or U39078 (N_39078,N_36160,N_35058);
nor U39079 (N_39079,N_36992,N_36048);
nand U39080 (N_39080,N_36229,N_36413);
and U39081 (N_39081,N_36992,N_36679);
or U39082 (N_39082,N_35092,N_36259);
or U39083 (N_39083,N_35801,N_35876);
or U39084 (N_39084,N_36382,N_35293);
and U39085 (N_39085,N_35881,N_36406);
and U39086 (N_39086,N_35603,N_37377);
nor U39087 (N_39087,N_36240,N_35920);
and U39088 (N_39088,N_35547,N_36051);
xnor U39089 (N_39089,N_36496,N_36703);
or U39090 (N_39090,N_36188,N_35484);
or U39091 (N_39091,N_36858,N_35073);
and U39092 (N_39092,N_35514,N_36080);
or U39093 (N_39093,N_35207,N_36022);
nand U39094 (N_39094,N_36601,N_35229);
and U39095 (N_39095,N_36676,N_35129);
nor U39096 (N_39096,N_36521,N_36861);
nand U39097 (N_39097,N_35765,N_35392);
xor U39098 (N_39098,N_36505,N_35095);
xor U39099 (N_39099,N_35863,N_35246);
xor U39100 (N_39100,N_36634,N_35312);
nor U39101 (N_39101,N_35476,N_37480);
nor U39102 (N_39102,N_36765,N_37175);
or U39103 (N_39103,N_35422,N_35991);
or U39104 (N_39104,N_35438,N_37112);
xor U39105 (N_39105,N_35895,N_35430);
or U39106 (N_39106,N_37391,N_35610);
nor U39107 (N_39107,N_37403,N_36080);
nand U39108 (N_39108,N_36774,N_36422);
or U39109 (N_39109,N_35890,N_36728);
and U39110 (N_39110,N_35296,N_36692);
nand U39111 (N_39111,N_36128,N_36256);
xor U39112 (N_39112,N_35897,N_37159);
xnor U39113 (N_39113,N_37008,N_35758);
and U39114 (N_39114,N_36374,N_36571);
nand U39115 (N_39115,N_35193,N_35130);
nand U39116 (N_39116,N_35919,N_35429);
nor U39117 (N_39117,N_35973,N_37218);
nor U39118 (N_39118,N_36707,N_36384);
and U39119 (N_39119,N_35685,N_35245);
xnor U39120 (N_39120,N_35011,N_36572);
or U39121 (N_39121,N_35039,N_35186);
xnor U39122 (N_39122,N_37492,N_35000);
nor U39123 (N_39123,N_35930,N_36601);
nand U39124 (N_39124,N_35903,N_36431);
and U39125 (N_39125,N_36982,N_35809);
nand U39126 (N_39126,N_37162,N_36566);
and U39127 (N_39127,N_35953,N_36521);
nand U39128 (N_39128,N_36855,N_37286);
nor U39129 (N_39129,N_37445,N_36695);
and U39130 (N_39130,N_35044,N_36406);
nand U39131 (N_39131,N_36396,N_35906);
nor U39132 (N_39132,N_36639,N_35855);
nand U39133 (N_39133,N_36119,N_35272);
or U39134 (N_39134,N_35432,N_35829);
nand U39135 (N_39135,N_36528,N_36269);
or U39136 (N_39136,N_36859,N_36307);
nand U39137 (N_39137,N_37485,N_35488);
and U39138 (N_39138,N_37464,N_35440);
nand U39139 (N_39139,N_35794,N_36858);
or U39140 (N_39140,N_35304,N_35960);
nand U39141 (N_39141,N_35038,N_35722);
and U39142 (N_39142,N_37123,N_35992);
nor U39143 (N_39143,N_36426,N_35433);
and U39144 (N_39144,N_37373,N_36722);
xor U39145 (N_39145,N_35382,N_35907);
nor U39146 (N_39146,N_35711,N_36320);
or U39147 (N_39147,N_36288,N_36732);
or U39148 (N_39148,N_37492,N_36087);
and U39149 (N_39149,N_36190,N_37041);
nor U39150 (N_39150,N_36670,N_35678);
nor U39151 (N_39151,N_37267,N_36704);
nand U39152 (N_39152,N_35041,N_36733);
xnor U39153 (N_39153,N_37399,N_37266);
or U39154 (N_39154,N_35283,N_35775);
nor U39155 (N_39155,N_35942,N_35594);
nor U39156 (N_39156,N_35076,N_36627);
and U39157 (N_39157,N_35159,N_36590);
nor U39158 (N_39158,N_36918,N_35306);
nand U39159 (N_39159,N_35924,N_37245);
nand U39160 (N_39160,N_35304,N_37217);
nand U39161 (N_39161,N_37337,N_35605);
and U39162 (N_39162,N_36274,N_35950);
nor U39163 (N_39163,N_35454,N_35911);
and U39164 (N_39164,N_37332,N_36592);
nand U39165 (N_39165,N_36353,N_36119);
and U39166 (N_39166,N_36477,N_36694);
or U39167 (N_39167,N_35168,N_35709);
or U39168 (N_39168,N_35700,N_37255);
xnor U39169 (N_39169,N_37004,N_36558);
nor U39170 (N_39170,N_37119,N_36424);
nand U39171 (N_39171,N_35280,N_35880);
xor U39172 (N_39172,N_35050,N_36901);
and U39173 (N_39173,N_36049,N_37027);
nand U39174 (N_39174,N_35777,N_35127);
nor U39175 (N_39175,N_37290,N_37245);
nor U39176 (N_39176,N_35079,N_36286);
nor U39177 (N_39177,N_36151,N_36599);
nand U39178 (N_39178,N_36349,N_35335);
xor U39179 (N_39179,N_37437,N_35955);
nor U39180 (N_39180,N_37497,N_37420);
xor U39181 (N_39181,N_36471,N_35580);
or U39182 (N_39182,N_36983,N_35492);
xnor U39183 (N_39183,N_35155,N_35683);
nand U39184 (N_39184,N_35015,N_36926);
nand U39185 (N_39185,N_35163,N_35786);
and U39186 (N_39186,N_36945,N_35313);
nand U39187 (N_39187,N_37012,N_36919);
or U39188 (N_39188,N_35602,N_36758);
nor U39189 (N_39189,N_37215,N_36028);
nand U39190 (N_39190,N_37316,N_37368);
xnor U39191 (N_39191,N_35577,N_35515);
and U39192 (N_39192,N_35625,N_36251);
nor U39193 (N_39193,N_35870,N_37315);
and U39194 (N_39194,N_37421,N_37259);
nand U39195 (N_39195,N_37043,N_36034);
nand U39196 (N_39196,N_35920,N_37350);
nand U39197 (N_39197,N_35463,N_36016);
and U39198 (N_39198,N_35131,N_36339);
nor U39199 (N_39199,N_35154,N_36655);
and U39200 (N_39200,N_35257,N_35299);
and U39201 (N_39201,N_36426,N_35087);
nand U39202 (N_39202,N_35163,N_36676);
and U39203 (N_39203,N_37372,N_37447);
nand U39204 (N_39204,N_36966,N_35296);
nor U39205 (N_39205,N_37142,N_36548);
and U39206 (N_39206,N_36684,N_36498);
nor U39207 (N_39207,N_36080,N_36296);
and U39208 (N_39208,N_35475,N_36828);
xor U39209 (N_39209,N_36732,N_35826);
and U39210 (N_39210,N_35120,N_35752);
nor U39211 (N_39211,N_35995,N_37035);
or U39212 (N_39212,N_37119,N_36350);
xor U39213 (N_39213,N_35358,N_37129);
nor U39214 (N_39214,N_35342,N_36226);
xnor U39215 (N_39215,N_36209,N_36272);
and U39216 (N_39216,N_35405,N_37462);
xor U39217 (N_39217,N_35513,N_37395);
nand U39218 (N_39218,N_35059,N_35269);
nor U39219 (N_39219,N_36176,N_35477);
nand U39220 (N_39220,N_37347,N_36336);
nor U39221 (N_39221,N_35042,N_36627);
or U39222 (N_39222,N_36707,N_35531);
nor U39223 (N_39223,N_36074,N_36642);
xnor U39224 (N_39224,N_35706,N_35640);
and U39225 (N_39225,N_36296,N_35456);
or U39226 (N_39226,N_35523,N_35601);
xor U39227 (N_39227,N_35167,N_35516);
xnor U39228 (N_39228,N_36724,N_36912);
or U39229 (N_39229,N_35283,N_35878);
xor U39230 (N_39230,N_36998,N_36065);
or U39231 (N_39231,N_36325,N_36308);
nand U39232 (N_39232,N_36874,N_35572);
xor U39233 (N_39233,N_35280,N_35707);
nor U39234 (N_39234,N_36616,N_36183);
nor U39235 (N_39235,N_35406,N_37204);
nand U39236 (N_39236,N_35343,N_35342);
nor U39237 (N_39237,N_36837,N_35554);
xor U39238 (N_39238,N_37307,N_37260);
nor U39239 (N_39239,N_35640,N_36477);
xor U39240 (N_39240,N_35047,N_36146);
or U39241 (N_39241,N_35796,N_36031);
nand U39242 (N_39242,N_37258,N_35481);
or U39243 (N_39243,N_36770,N_35576);
and U39244 (N_39244,N_35492,N_36617);
xnor U39245 (N_39245,N_35967,N_36346);
xor U39246 (N_39246,N_35322,N_36829);
and U39247 (N_39247,N_35431,N_35673);
nand U39248 (N_39248,N_37481,N_36032);
and U39249 (N_39249,N_36977,N_35859);
and U39250 (N_39250,N_36276,N_36776);
or U39251 (N_39251,N_36092,N_35795);
and U39252 (N_39252,N_35229,N_35430);
and U39253 (N_39253,N_35026,N_35206);
or U39254 (N_39254,N_35426,N_35084);
and U39255 (N_39255,N_37002,N_36274);
and U39256 (N_39256,N_35596,N_36343);
nor U39257 (N_39257,N_35402,N_35999);
or U39258 (N_39258,N_37311,N_35255);
nand U39259 (N_39259,N_35612,N_35431);
xnor U39260 (N_39260,N_36354,N_35518);
nand U39261 (N_39261,N_35465,N_35676);
xnor U39262 (N_39262,N_36133,N_35604);
nor U39263 (N_39263,N_37102,N_37187);
or U39264 (N_39264,N_37225,N_37369);
nor U39265 (N_39265,N_37129,N_36760);
nand U39266 (N_39266,N_37331,N_36552);
or U39267 (N_39267,N_35027,N_35611);
xnor U39268 (N_39268,N_35664,N_35242);
xor U39269 (N_39269,N_36314,N_36807);
xor U39270 (N_39270,N_36795,N_36911);
nor U39271 (N_39271,N_36139,N_35630);
or U39272 (N_39272,N_35636,N_35443);
and U39273 (N_39273,N_35481,N_37322);
nor U39274 (N_39274,N_37179,N_35875);
xnor U39275 (N_39275,N_36821,N_37084);
xor U39276 (N_39276,N_35995,N_36865);
nand U39277 (N_39277,N_36960,N_36174);
or U39278 (N_39278,N_36602,N_36062);
or U39279 (N_39279,N_35340,N_35442);
or U39280 (N_39280,N_35615,N_36988);
nor U39281 (N_39281,N_36844,N_36065);
xor U39282 (N_39282,N_35566,N_35980);
and U39283 (N_39283,N_35874,N_37344);
or U39284 (N_39284,N_36257,N_35915);
and U39285 (N_39285,N_36791,N_35451);
nor U39286 (N_39286,N_35458,N_36091);
nand U39287 (N_39287,N_35977,N_36332);
and U39288 (N_39288,N_36402,N_35415);
and U39289 (N_39289,N_35292,N_37260);
and U39290 (N_39290,N_37241,N_35520);
nor U39291 (N_39291,N_35287,N_36272);
or U39292 (N_39292,N_36231,N_36827);
or U39293 (N_39293,N_35930,N_35368);
nor U39294 (N_39294,N_36023,N_35827);
nor U39295 (N_39295,N_35449,N_36242);
and U39296 (N_39296,N_35303,N_36331);
xnor U39297 (N_39297,N_37110,N_37390);
or U39298 (N_39298,N_37009,N_36113);
and U39299 (N_39299,N_35151,N_36743);
xnor U39300 (N_39300,N_35758,N_37065);
nand U39301 (N_39301,N_35356,N_36227);
xnor U39302 (N_39302,N_37092,N_36244);
nor U39303 (N_39303,N_36656,N_36225);
nand U39304 (N_39304,N_36659,N_36316);
nand U39305 (N_39305,N_36824,N_36014);
nor U39306 (N_39306,N_35844,N_36067);
xor U39307 (N_39307,N_35265,N_35488);
nor U39308 (N_39308,N_36032,N_36293);
and U39309 (N_39309,N_36595,N_35734);
xnor U39310 (N_39310,N_36300,N_35235);
nor U39311 (N_39311,N_35348,N_35637);
xnor U39312 (N_39312,N_35894,N_35707);
xnor U39313 (N_39313,N_35284,N_37434);
nor U39314 (N_39314,N_35183,N_36634);
or U39315 (N_39315,N_35848,N_36041);
nor U39316 (N_39316,N_37139,N_36341);
nor U39317 (N_39317,N_35622,N_35575);
or U39318 (N_39318,N_35174,N_35884);
nand U39319 (N_39319,N_37194,N_35932);
nor U39320 (N_39320,N_35283,N_36898);
xnor U39321 (N_39321,N_36774,N_35820);
or U39322 (N_39322,N_36510,N_36655);
nand U39323 (N_39323,N_36537,N_36295);
or U39324 (N_39324,N_36840,N_36151);
nor U39325 (N_39325,N_36546,N_37059);
xor U39326 (N_39326,N_37250,N_37339);
and U39327 (N_39327,N_36290,N_35878);
nand U39328 (N_39328,N_36913,N_36723);
and U39329 (N_39329,N_36535,N_37313);
or U39330 (N_39330,N_35770,N_36988);
nand U39331 (N_39331,N_35718,N_36186);
xnor U39332 (N_39332,N_36610,N_36037);
or U39333 (N_39333,N_35551,N_35555);
and U39334 (N_39334,N_35689,N_36904);
and U39335 (N_39335,N_36951,N_35400);
nand U39336 (N_39336,N_36503,N_35299);
nor U39337 (N_39337,N_36146,N_37229);
nand U39338 (N_39338,N_36814,N_35077);
nand U39339 (N_39339,N_36677,N_35069);
and U39340 (N_39340,N_36714,N_36440);
nand U39341 (N_39341,N_37363,N_35878);
and U39342 (N_39342,N_36688,N_35578);
or U39343 (N_39343,N_37345,N_36102);
or U39344 (N_39344,N_35011,N_35751);
and U39345 (N_39345,N_37442,N_36488);
xnor U39346 (N_39346,N_35070,N_36089);
xnor U39347 (N_39347,N_37368,N_35268);
nand U39348 (N_39348,N_37138,N_37454);
xor U39349 (N_39349,N_37274,N_35907);
xnor U39350 (N_39350,N_36256,N_35134);
nor U39351 (N_39351,N_35080,N_37048);
and U39352 (N_39352,N_36619,N_37003);
nor U39353 (N_39353,N_36301,N_36312);
or U39354 (N_39354,N_36170,N_35938);
nor U39355 (N_39355,N_35167,N_37357);
and U39356 (N_39356,N_36998,N_36338);
nand U39357 (N_39357,N_35120,N_35093);
or U39358 (N_39358,N_36715,N_36207);
nor U39359 (N_39359,N_35376,N_36860);
nand U39360 (N_39360,N_36428,N_35954);
nor U39361 (N_39361,N_35811,N_36124);
xnor U39362 (N_39362,N_35206,N_37140);
nand U39363 (N_39363,N_35196,N_37312);
xnor U39364 (N_39364,N_37188,N_36486);
nand U39365 (N_39365,N_37306,N_37149);
and U39366 (N_39366,N_36224,N_36096);
nor U39367 (N_39367,N_35006,N_36876);
nor U39368 (N_39368,N_36524,N_36303);
xnor U39369 (N_39369,N_37140,N_36738);
and U39370 (N_39370,N_36094,N_36662);
nor U39371 (N_39371,N_36203,N_36310);
or U39372 (N_39372,N_35623,N_36043);
nand U39373 (N_39373,N_37294,N_37458);
and U39374 (N_39374,N_36948,N_37194);
nand U39375 (N_39375,N_36679,N_36036);
xor U39376 (N_39376,N_36286,N_35928);
nand U39377 (N_39377,N_36733,N_35039);
or U39378 (N_39378,N_35583,N_35439);
or U39379 (N_39379,N_37127,N_36658);
or U39380 (N_39380,N_35540,N_36655);
nor U39381 (N_39381,N_36840,N_35488);
nor U39382 (N_39382,N_37326,N_35779);
xor U39383 (N_39383,N_37005,N_37112);
or U39384 (N_39384,N_35724,N_37236);
nand U39385 (N_39385,N_35185,N_35899);
and U39386 (N_39386,N_36090,N_37152);
or U39387 (N_39387,N_36178,N_35997);
or U39388 (N_39388,N_35238,N_36660);
xnor U39389 (N_39389,N_37396,N_35706);
xor U39390 (N_39390,N_36169,N_35384);
and U39391 (N_39391,N_37063,N_36109);
nor U39392 (N_39392,N_36151,N_36770);
xnor U39393 (N_39393,N_36339,N_36556);
xor U39394 (N_39394,N_36149,N_36012);
xnor U39395 (N_39395,N_35186,N_37022);
or U39396 (N_39396,N_35192,N_37266);
nand U39397 (N_39397,N_35020,N_35860);
xnor U39398 (N_39398,N_36952,N_36010);
and U39399 (N_39399,N_37217,N_36663);
or U39400 (N_39400,N_37016,N_37010);
nor U39401 (N_39401,N_35179,N_37493);
nand U39402 (N_39402,N_35401,N_35187);
and U39403 (N_39403,N_36898,N_35897);
nand U39404 (N_39404,N_35758,N_36585);
nor U39405 (N_39405,N_36361,N_36730);
nor U39406 (N_39406,N_35256,N_36770);
or U39407 (N_39407,N_36331,N_35278);
or U39408 (N_39408,N_37299,N_35135);
xor U39409 (N_39409,N_35900,N_36839);
or U39410 (N_39410,N_35713,N_36339);
nand U39411 (N_39411,N_36350,N_36256);
or U39412 (N_39412,N_37090,N_37484);
nor U39413 (N_39413,N_35855,N_35247);
or U39414 (N_39414,N_36496,N_36513);
nand U39415 (N_39415,N_35117,N_35531);
and U39416 (N_39416,N_35235,N_35795);
nor U39417 (N_39417,N_36372,N_36353);
nand U39418 (N_39418,N_35786,N_36393);
xnor U39419 (N_39419,N_36493,N_35111);
nand U39420 (N_39420,N_35477,N_35312);
nor U39421 (N_39421,N_36805,N_35840);
nand U39422 (N_39422,N_35143,N_37091);
nor U39423 (N_39423,N_36306,N_37104);
xnor U39424 (N_39424,N_37179,N_37186);
xnor U39425 (N_39425,N_35750,N_36619);
and U39426 (N_39426,N_36581,N_37372);
and U39427 (N_39427,N_35334,N_35354);
xor U39428 (N_39428,N_35228,N_36541);
and U39429 (N_39429,N_35611,N_35311);
xnor U39430 (N_39430,N_36677,N_37345);
and U39431 (N_39431,N_35897,N_36322);
xor U39432 (N_39432,N_35742,N_36322);
and U39433 (N_39433,N_37252,N_35670);
nand U39434 (N_39434,N_35152,N_36503);
nor U39435 (N_39435,N_35568,N_36907);
or U39436 (N_39436,N_36512,N_36716);
or U39437 (N_39437,N_36737,N_36065);
nand U39438 (N_39438,N_36986,N_35050);
nand U39439 (N_39439,N_36367,N_36081);
nand U39440 (N_39440,N_36078,N_36979);
xor U39441 (N_39441,N_35157,N_36158);
xnor U39442 (N_39442,N_36797,N_35852);
nand U39443 (N_39443,N_36821,N_36031);
or U39444 (N_39444,N_35116,N_36496);
and U39445 (N_39445,N_36140,N_37175);
and U39446 (N_39446,N_36135,N_36053);
xnor U39447 (N_39447,N_36978,N_36664);
nor U39448 (N_39448,N_37437,N_36060);
nand U39449 (N_39449,N_35825,N_35979);
and U39450 (N_39450,N_35916,N_36266);
or U39451 (N_39451,N_35959,N_35143);
nand U39452 (N_39452,N_35322,N_35432);
nor U39453 (N_39453,N_36751,N_36507);
nand U39454 (N_39454,N_36642,N_35833);
or U39455 (N_39455,N_36650,N_37240);
xor U39456 (N_39456,N_35362,N_35759);
or U39457 (N_39457,N_35832,N_37488);
nand U39458 (N_39458,N_35493,N_36783);
xnor U39459 (N_39459,N_36169,N_35508);
nor U39460 (N_39460,N_35822,N_37379);
or U39461 (N_39461,N_36154,N_35996);
and U39462 (N_39462,N_37304,N_36827);
nor U39463 (N_39463,N_36787,N_36223);
and U39464 (N_39464,N_35571,N_36601);
xnor U39465 (N_39465,N_36911,N_36604);
nand U39466 (N_39466,N_35976,N_36587);
nor U39467 (N_39467,N_37131,N_36608);
and U39468 (N_39468,N_35578,N_36795);
or U39469 (N_39469,N_36510,N_35111);
and U39470 (N_39470,N_35974,N_35767);
and U39471 (N_39471,N_37382,N_35451);
nor U39472 (N_39472,N_36528,N_36861);
or U39473 (N_39473,N_36700,N_35662);
nand U39474 (N_39474,N_36403,N_36599);
or U39475 (N_39475,N_36306,N_36667);
nor U39476 (N_39476,N_35964,N_35141);
or U39477 (N_39477,N_36680,N_35971);
nand U39478 (N_39478,N_36047,N_36109);
nor U39479 (N_39479,N_36295,N_37382);
nand U39480 (N_39480,N_36837,N_36890);
nor U39481 (N_39481,N_37122,N_37315);
nor U39482 (N_39482,N_35744,N_35961);
nand U39483 (N_39483,N_36426,N_35647);
xor U39484 (N_39484,N_36725,N_37316);
or U39485 (N_39485,N_35251,N_35699);
xnor U39486 (N_39486,N_37088,N_36929);
or U39487 (N_39487,N_36196,N_36542);
nand U39488 (N_39488,N_36769,N_35379);
nor U39489 (N_39489,N_36411,N_37090);
nor U39490 (N_39490,N_37100,N_37202);
or U39491 (N_39491,N_35509,N_35228);
nand U39492 (N_39492,N_36905,N_36503);
nand U39493 (N_39493,N_35081,N_37079);
or U39494 (N_39494,N_36289,N_36091);
and U39495 (N_39495,N_37344,N_35391);
or U39496 (N_39496,N_35266,N_36270);
or U39497 (N_39497,N_35034,N_37013);
and U39498 (N_39498,N_37390,N_35046);
xnor U39499 (N_39499,N_36050,N_36307);
or U39500 (N_39500,N_35184,N_35007);
or U39501 (N_39501,N_35147,N_37377);
xnor U39502 (N_39502,N_36854,N_37161);
nand U39503 (N_39503,N_36379,N_37196);
or U39504 (N_39504,N_37404,N_36703);
and U39505 (N_39505,N_36138,N_35487);
or U39506 (N_39506,N_35488,N_36562);
xor U39507 (N_39507,N_35519,N_36251);
or U39508 (N_39508,N_36605,N_35723);
or U39509 (N_39509,N_37120,N_36856);
nor U39510 (N_39510,N_36430,N_35923);
nand U39511 (N_39511,N_36680,N_36042);
xor U39512 (N_39512,N_35683,N_36980);
xor U39513 (N_39513,N_36593,N_35133);
xnor U39514 (N_39514,N_37443,N_35945);
nand U39515 (N_39515,N_35055,N_36374);
nand U39516 (N_39516,N_35030,N_35488);
nor U39517 (N_39517,N_36773,N_35267);
nand U39518 (N_39518,N_36279,N_37474);
or U39519 (N_39519,N_36403,N_35557);
and U39520 (N_39520,N_36651,N_35038);
nand U39521 (N_39521,N_35288,N_36377);
nor U39522 (N_39522,N_35622,N_36883);
or U39523 (N_39523,N_37016,N_36035);
nor U39524 (N_39524,N_36753,N_36305);
nor U39525 (N_39525,N_35515,N_37024);
nor U39526 (N_39526,N_37261,N_35870);
xnor U39527 (N_39527,N_35322,N_36275);
and U39528 (N_39528,N_36240,N_36381);
nor U39529 (N_39529,N_36427,N_35734);
xor U39530 (N_39530,N_35116,N_36298);
nor U39531 (N_39531,N_36837,N_35168);
or U39532 (N_39532,N_37366,N_36756);
and U39533 (N_39533,N_36296,N_35193);
and U39534 (N_39534,N_35506,N_37242);
nand U39535 (N_39535,N_35957,N_37143);
nand U39536 (N_39536,N_36077,N_35540);
nand U39537 (N_39537,N_35717,N_35284);
nor U39538 (N_39538,N_36861,N_35388);
or U39539 (N_39539,N_37336,N_36369);
xnor U39540 (N_39540,N_35758,N_35773);
and U39541 (N_39541,N_36526,N_37028);
xnor U39542 (N_39542,N_35707,N_36572);
or U39543 (N_39543,N_35496,N_37391);
nand U39544 (N_39544,N_35038,N_37273);
nor U39545 (N_39545,N_35976,N_35526);
xor U39546 (N_39546,N_37257,N_36519);
nor U39547 (N_39547,N_36725,N_35572);
or U39548 (N_39548,N_37446,N_35002);
nand U39549 (N_39549,N_36006,N_36967);
or U39550 (N_39550,N_36372,N_36322);
or U39551 (N_39551,N_36943,N_35892);
xor U39552 (N_39552,N_36013,N_35021);
or U39553 (N_39553,N_35885,N_37205);
nand U39554 (N_39554,N_36283,N_36452);
or U39555 (N_39555,N_37127,N_35704);
xnor U39556 (N_39556,N_37232,N_36141);
and U39557 (N_39557,N_37419,N_36900);
and U39558 (N_39558,N_36608,N_35426);
or U39559 (N_39559,N_35554,N_35524);
and U39560 (N_39560,N_35387,N_36793);
nor U39561 (N_39561,N_35848,N_37335);
and U39562 (N_39562,N_37131,N_35875);
and U39563 (N_39563,N_36869,N_35085);
nor U39564 (N_39564,N_37397,N_35795);
nand U39565 (N_39565,N_35514,N_36618);
nand U39566 (N_39566,N_35742,N_35416);
xnor U39567 (N_39567,N_36697,N_36087);
or U39568 (N_39568,N_35839,N_35471);
and U39569 (N_39569,N_36987,N_37071);
nor U39570 (N_39570,N_35563,N_36961);
nand U39571 (N_39571,N_35486,N_36188);
nand U39572 (N_39572,N_35447,N_36693);
nor U39573 (N_39573,N_36688,N_36101);
nand U39574 (N_39574,N_36521,N_35266);
nand U39575 (N_39575,N_36100,N_35334);
nand U39576 (N_39576,N_35860,N_35096);
and U39577 (N_39577,N_37383,N_36158);
nand U39578 (N_39578,N_36640,N_35284);
xor U39579 (N_39579,N_37402,N_36299);
nor U39580 (N_39580,N_35495,N_36221);
and U39581 (N_39581,N_35405,N_36865);
and U39582 (N_39582,N_36733,N_37384);
or U39583 (N_39583,N_37439,N_36261);
nand U39584 (N_39584,N_35639,N_37174);
or U39585 (N_39585,N_35805,N_37131);
nor U39586 (N_39586,N_37441,N_36956);
xor U39587 (N_39587,N_36505,N_35256);
or U39588 (N_39588,N_35432,N_36398);
and U39589 (N_39589,N_36473,N_35723);
and U39590 (N_39590,N_36172,N_35834);
nand U39591 (N_39591,N_35373,N_36891);
or U39592 (N_39592,N_35803,N_36225);
nand U39593 (N_39593,N_35436,N_36902);
or U39594 (N_39594,N_36724,N_36567);
xor U39595 (N_39595,N_37112,N_35578);
xor U39596 (N_39596,N_35696,N_36421);
and U39597 (N_39597,N_36511,N_36622);
xnor U39598 (N_39598,N_35521,N_36278);
or U39599 (N_39599,N_36297,N_36941);
and U39600 (N_39600,N_36400,N_36106);
xnor U39601 (N_39601,N_36886,N_35090);
and U39602 (N_39602,N_36098,N_35974);
and U39603 (N_39603,N_37304,N_37141);
nor U39604 (N_39604,N_35845,N_36931);
xor U39605 (N_39605,N_37019,N_35318);
nand U39606 (N_39606,N_36610,N_37328);
and U39607 (N_39607,N_37023,N_35153);
nor U39608 (N_39608,N_37137,N_37275);
xnor U39609 (N_39609,N_35186,N_35814);
nor U39610 (N_39610,N_35592,N_35634);
and U39611 (N_39611,N_35550,N_37414);
or U39612 (N_39612,N_36295,N_35875);
nand U39613 (N_39613,N_36911,N_36509);
or U39614 (N_39614,N_36366,N_35874);
and U39615 (N_39615,N_36764,N_36030);
or U39616 (N_39616,N_37133,N_36509);
and U39617 (N_39617,N_36140,N_35675);
nor U39618 (N_39618,N_35462,N_36543);
xor U39619 (N_39619,N_35310,N_37305);
or U39620 (N_39620,N_36158,N_36866);
or U39621 (N_39621,N_36570,N_37338);
nand U39622 (N_39622,N_36822,N_35495);
nand U39623 (N_39623,N_37265,N_36744);
xnor U39624 (N_39624,N_36473,N_35416);
nand U39625 (N_39625,N_35655,N_37133);
nor U39626 (N_39626,N_36910,N_35720);
nand U39627 (N_39627,N_36855,N_37195);
xor U39628 (N_39628,N_36849,N_36725);
nand U39629 (N_39629,N_36755,N_36364);
and U39630 (N_39630,N_36649,N_37463);
and U39631 (N_39631,N_35570,N_37032);
nand U39632 (N_39632,N_37359,N_36935);
nand U39633 (N_39633,N_35875,N_35912);
nand U39634 (N_39634,N_36414,N_36887);
nand U39635 (N_39635,N_36591,N_36476);
xnor U39636 (N_39636,N_35594,N_36179);
or U39637 (N_39637,N_37239,N_36607);
and U39638 (N_39638,N_35804,N_36204);
and U39639 (N_39639,N_35149,N_36472);
nand U39640 (N_39640,N_37314,N_37361);
and U39641 (N_39641,N_36044,N_36016);
nor U39642 (N_39642,N_35730,N_35877);
and U39643 (N_39643,N_37417,N_37100);
and U39644 (N_39644,N_37462,N_36954);
or U39645 (N_39645,N_35454,N_36512);
xnor U39646 (N_39646,N_35412,N_35103);
xor U39647 (N_39647,N_36448,N_37406);
and U39648 (N_39648,N_35451,N_37051);
or U39649 (N_39649,N_37442,N_35881);
nand U39650 (N_39650,N_37066,N_35218);
and U39651 (N_39651,N_37412,N_36637);
nor U39652 (N_39652,N_35979,N_35938);
or U39653 (N_39653,N_36650,N_35854);
or U39654 (N_39654,N_36445,N_35199);
nand U39655 (N_39655,N_36408,N_37234);
or U39656 (N_39656,N_35310,N_37187);
nand U39657 (N_39657,N_36520,N_35763);
and U39658 (N_39658,N_35928,N_36559);
xor U39659 (N_39659,N_35585,N_35017);
or U39660 (N_39660,N_36188,N_35086);
and U39661 (N_39661,N_36369,N_37217);
nand U39662 (N_39662,N_37385,N_36353);
nand U39663 (N_39663,N_35331,N_35614);
and U39664 (N_39664,N_36944,N_37475);
nand U39665 (N_39665,N_35014,N_37140);
and U39666 (N_39666,N_36663,N_35493);
xnor U39667 (N_39667,N_35898,N_36672);
or U39668 (N_39668,N_36254,N_35122);
nand U39669 (N_39669,N_35229,N_36775);
and U39670 (N_39670,N_35588,N_36836);
nand U39671 (N_39671,N_36598,N_35731);
and U39672 (N_39672,N_35325,N_35646);
and U39673 (N_39673,N_36070,N_36832);
nand U39674 (N_39674,N_35474,N_36888);
or U39675 (N_39675,N_35443,N_37443);
and U39676 (N_39676,N_36620,N_35902);
xor U39677 (N_39677,N_35720,N_36307);
nor U39678 (N_39678,N_36249,N_37395);
and U39679 (N_39679,N_36085,N_35044);
or U39680 (N_39680,N_35866,N_36291);
or U39681 (N_39681,N_36389,N_36297);
and U39682 (N_39682,N_35703,N_36566);
or U39683 (N_39683,N_36113,N_37143);
nand U39684 (N_39684,N_36970,N_37458);
nor U39685 (N_39685,N_35145,N_35985);
nand U39686 (N_39686,N_35431,N_37386);
nand U39687 (N_39687,N_36671,N_36981);
and U39688 (N_39688,N_37217,N_35863);
nand U39689 (N_39689,N_36731,N_36415);
nor U39690 (N_39690,N_36019,N_35836);
nand U39691 (N_39691,N_35675,N_37064);
nor U39692 (N_39692,N_36470,N_37459);
or U39693 (N_39693,N_36763,N_36114);
nor U39694 (N_39694,N_36515,N_37192);
nand U39695 (N_39695,N_37493,N_35251);
xor U39696 (N_39696,N_35993,N_36977);
and U39697 (N_39697,N_35864,N_36435);
xor U39698 (N_39698,N_36776,N_37448);
or U39699 (N_39699,N_35832,N_36432);
and U39700 (N_39700,N_36353,N_36528);
or U39701 (N_39701,N_36443,N_36611);
nand U39702 (N_39702,N_35139,N_36937);
or U39703 (N_39703,N_36269,N_36199);
xnor U39704 (N_39704,N_36263,N_35353);
xor U39705 (N_39705,N_36055,N_36969);
or U39706 (N_39706,N_35528,N_35073);
nand U39707 (N_39707,N_36105,N_36025);
or U39708 (N_39708,N_36126,N_35149);
nor U39709 (N_39709,N_36066,N_35603);
or U39710 (N_39710,N_35639,N_37436);
and U39711 (N_39711,N_36580,N_35794);
nor U39712 (N_39712,N_36503,N_36320);
or U39713 (N_39713,N_35144,N_36810);
nor U39714 (N_39714,N_35055,N_37047);
nand U39715 (N_39715,N_35694,N_35863);
xor U39716 (N_39716,N_35158,N_36690);
or U39717 (N_39717,N_36586,N_36530);
nand U39718 (N_39718,N_37142,N_37497);
nand U39719 (N_39719,N_35542,N_35753);
nand U39720 (N_39720,N_36547,N_36004);
nor U39721 (N_39721,N_36129,N_37007);
xor U39722 (N_39722,N_35445,N_35157);
and U39723 (N_39723,N_35549,N_37399);
xor U39724 (N_39724,N_36258,N_35665);
nor U39725 (N_39725,N_35260,N_35139);
nand U39726 (N_39726,N_35167,N_36350);
xnor U39727 (N_39727,N_35056,N_35980);
nand U39728 (N_39728,N_37018,N_37184);
or U39729 (N_39729,N_36515,N_37087);
and U39730 (N_39730,N_35352,N_35999);
xnor U39731 (N_39731,N_35396,N_36790);
nor U39732 (N_39732,N_36740,N_36080);
or U39733 (N_39733,N_35871,N_35556);
xor U39734 (N_39734,N_36293,N_37171);
nand U39735 (N_39735,N_36915,N_36168);
nand U39736 (N_39736,N_35444,N_36609);
and U39737 (N_39737,N_36262,N_36193);
xor U39738 (N_39738,N_35350,N_37043);
nor U39739 (N_39739,N_35442,N_36616);
xnor U39740 (N_39740,N_35535,N_36181);
xor U39741 (N_39741,N_35795,N_36713);
or U39742 (N_39742,N_36567,N_35648);
and U39743 (N_39743,N_36703,N_36805);
xor U39744 (N_39744,N_37299,N_35210);
and U39745 (N_39745,N_36223,N_35227);
nor U39746 (N_39746,N_37209,N_35965);
xnor U39747 (N_39747,N_36305,N_37232);
or U39748 (N_39748,N_36184,N_36310);
and U39749 (N_39749,N_36018,N_36186);
nand U39750 (N_39750,N_35475,N_36761);
or U39751 (N_39751,N_36974,N_35795);
and U39752 (N_39752,N_37000,N_36265);
xor U39753 (N_39753,N_37353,N_36581);
and U39754 (N_39754,N_35623,N_36166);
xor U39755 (N_39755,N_36329,N_35952);
nand U39756 (N_39756,N_36760,N_37264);
xor U39757 (N_39757,N_35018,N_37397);
nor U39758 (N_39758,N_36297,N_36212);
nor U39759 (N_39759,N_37277,N_36750);
xnor U39760 (N_39760,N_36592,N_35427);
nor U39761 (N_39761,N_37492,N_35022);
or U39762 (N_39762,N_35586,N_37167);
nand U39763 (N_39763,N_35219,N_37055);
and U39764 (N_39764,N_36017,N_37066);
or U39765 (N_39765,N_36408,N_36591);
or U39766 (N_39766,N_37178,N_35026);
or U39767 (N_39767,N_36734,N_37136);
nor U39768 (N_39768,N_36388,N_35241);
nor U39769 (N_39769,N_37088,N_37375);
xnor U39770 (N_39770,N_35662,N_36325);
and U39771 (N_39771,N_36772,N_35187);
nand U39772 (N_39772,N_36626,N_36438);
nor U39773 (N_39773,N_36657,N_35562);
and U39774 (N_39774,N_36017,N_36334);
nand U39775 (N_39775,N_36400,N_35727);
or U39776 (N_39776,N_36273,N_35854);
or U39777 (N_39777,N_35633,N_35392);
and U39778 (N_39778,N_35124,N_37447);
or U39779 (N_39779,N_35500,N_37448);
xnor U39780 (N_39780,N_36436,N_37164);
nor U39781 (N_39781,N_37494,N_37095);
and U39782 (N_39782,N_36429,N_35683);
nor U39783 (N_39783,N_35959,N_36496);
and U39784 (N_39784,N_36652,N_35901);
and U39785 (N_39785,N_36142,N_37379);
and U39786 (N_39786,N_35074,N_35068);
nor U39787 (N_39787,N_37248,N_37356);
or U39788 (N_39788,N_35192,N_35987);
nor U39789 (N_39789,N_36681,N_35368);
nand U39790 (N_39790,N_36604,N_35274);
nor U39791 (N_39791,N_35290,N_35989);
nor U39792 (N_39792,N_36305,N_36698);
and U39793 (N_39793,N_35535,N_35239);
and U39794 (N_39794,N_35323,N_37434);
nor U39795 (N_39795,N_37444,N_35278);
and U39796 (N_39796,N_37426,N_35855);
or U39797 (N_39797,N_35812,N_35746);
or U39798 (N_39798,N_36725,N_35566);
nand U39799 (N_39799,N_36919,N_36142);
or U39800 (N_39800,N_35701,N_35559);
nand U39801 (N_39801,N_35432,N_35775);
nor U39802 (N_39802,N_37304,N_36946);
xnor U39803 (N_39803,N_36420,N_36969);
or U39804 (N_39804,N_36781,N_35871);
xor U39805 (N_39805,N_36320,N_37194);
xor U39806 (N_39806,N_36231,N_35717);
or U39807 (N_39807,N_35306,N_37350);
or U39808 (N_39808,N_36269,N_36416);
xor U39809 (N_39809,N_36764,N_37017);
xnor U39810 (N_39810,N_37045,N_36084);
xnor U39811 (N_39811,N_35905,N_37193);
nand U39812 (N_39812,N_35027,N_35024);
nor U39813 (N_39813,N_37079,N_35257);
nor U39814 (N_39814,N_36142,N_35683);
and U39815 (N_39815,N_37426,N_35055);
xnor U39816 (N_39816,N_37376,N_37481);
or U39817 (N_39817,N_37438,N_36620);
or U39818 (N_39818,N_36191,N_36081);
or U39819 (N_39819,N_36333,N_36805);
or U39820 (N_39820,N_36928,N_36457);
nand U39821 (N_39821,N_36153,N_36528);
xnor U39822 (N_39822,N_35381,N_35374);
or U39823 (N_39823,N_35438,N_36054);
nor U39824 (N_39824,N_36365,N_35553);
nand U39825 (N_39825,N_35941,N_35585);
and U39826 (N_39826,N_35907,N_37439);
nor U39827 (N_39827,N_36349,N_35937);
or U39828 (N_39828,N_35814,N_35651);
xnor U39829 (N_39829,N_36547,N_35644);
and U39830 (N_39830,N_37048,N_35226);
xnor U39831 (N_39831,N_35848,N_35354);
and U39832 (N_39832,N_36219,N_37238);
or U39833 (N_39833,N_37139,N_36213);
and U39834 (N_39834,N_35865,N_36458);
nor U39835 (N_39835,N_36234,N_37363);
and U39836 (N_39836,N_36458,N_35718);
or U39837 (N_39837,N_36116,N_35012);
nor U39838 (N_39838,N_37288,N_36186);
nor U39839 (N_39839,N_36864,N_35599);
and U39840 (N_39840,N_35148,N_36053);
xnor U39841 (N_39841,N_36240,N_36557);
or U39842 (N_39842,N_36476,N_35918);
and U39843 (N_39843,N_35708,N_37120);
nor U39844 (N_39844,N_36811,N_36184);
or U39845 (N_39845,N_36926,N_35598);
nor U39846 (N_39846,N_35365,N_35257);
and U39847 (N_39847,N_37111,N_36843);
nand U39848 (N_39848,N_37259,N_36083);
or U39849 (N_39849,N_35946,N_36422);
and U39850 (N_39850,N_36620,N_36301);
and U39851 (N_39851,N_37383,N_36445);
and U39852 (N_39852,N_37285,N_35245);
nand U39853 (N_39853,N_37407,N_35327);
xor U39854 (N_39854,N_37096,N_36214);
or U39855 (N_39855,N_35094,N_36207);
and U39856 (N_39856,N_35203,N_37490);
and U39857 (N_39857,N_36339,N_35345);
nand U39858 (N_39858,N_36242,N_35290);
nor U39859 (N_39859,N_36621,N_35506);
or U39860 (N_39860,N_36573,N_37146);
or U39861 (N_39861,N_37144,N_37088);
and U39862 (N_39862,N_35329,N_35945);
and U39863 (N_39863,N_36189,N_35833);
and U39864 (N_39864,N_37149,N_37169);
and U39865 (N_39865,N_35426,N_36920);
xnor U39866 (N_39866,N_35782,N_36866);
nand U39867 (N_39867,N_35962,N_36853);
nand U39868 (N_39868,N_37321,N_35844);
or U39869 (N_39869,N_36439,N_35793);
nand U39870 (N_39870,N_35587,N_35117);
or U39871 (N_39871,N_37193,N_35471);
xnor U39872 (N_39872,N_37190,N_36369);
and U39873 (N_39873,N_36161,N_37372);
and U39874 (N_39874,N_35513,N_35618);
nor U39875 (N_39875,N_36565,N_35454);
nand U39876 (N_39876,N_37197,N_37075);
nand U39877 (N_39877,N_37431,N_35319);
xnor U39878 (N_39878,N_36867,N_35237);
xnor U39879 (N_39879,N_36768,N_35721);
or U39880 (N_39880,N_36101,N_36815);
nor U39881 (N_39881,N_37188,N_35073);
or U39882 (N_39882,N_35435,N_35916);
and U39883 (N_39883,N_37036,N_36045);
nor U39884 (N_39884,N_36000,N_36809);
xor U39885 (N_39885,N_37172,N_36020);
or U39886 (N_39886,N_36363,N_35565);
or U39887 (N_39887,N_35968,N_36105);
or U39888 (N_39888,N_36763,N_35841);
xnor U39889 (N_39889,N_35918,N_36010);
xor U39890 (N_39890,N_35200,N_36908);
xor U39891 (N_39891,N_37143,N_35953);
and U39892 (N_39892,N_35001,N_35349);
xor U39893 (N_39893,N_36499,N_36517);
and U39894 (N_39894,N_36987,N_36623);
nor U39895 (N_39895,N_37192,N_35147);
nand U39896 (N_39896,N_36400,N_36050);
nor U39897 (N_39897,N_37215,N_35877);
or U39898 (N_39898,N_36495,N_35571);
nand U39899 (N_39899,N_36008,N_35013);
or U39900 (N_39900,N_35227,N_35386);
nand U39901 (N_39901,N_37261,N_37250);
xnor U39902 (N_39902,N_36697,N_35376);
and U39903 (N_39903,N_36347,N_35701);
or U39904 (N_39904,N_36337,N_36678);
nor U39905 (N_39905,N_35177,N_35107);
and U39906 (N_39906,N_36312,N_35842);
and U39907 (N_39907,N_35465,N_35122);
nor U39908 (N_39908,N_36071,N_37192);
nand U39909 (N_39909,N_37435,N_35509);
and U39910 (N_39910,N_37108,N_35080);
or U39911 (N_39911,N_36264,N_36169);
nor U39912 (N_39912,N_35740,N_36567);
or U39913 (N_39913,N_36365,N_35410);
xnor U39914 (N_39914,N_36243,N_35317);
or U39915 (N_39915,N_35094,N_35992);
or U39916 (N_39916,N_36095,N_36576);
or U39917 (N_39917,N_35741,N_37130);
nand U39918 (N_39918,N_36526,N_35041);
or U39919 (N_39919,N_36312,N_36648);
nand U39920 (N_39920,N_37137,N_35399);
nor U39921 (N_39921,N_37207,N_36382);
xnor U39922 (N_39922,N_36140,N_35724);
nand U39923 (N_39923,N_36037,N_35320);
nor U39924 (N_39924,N_35533,N_37490);
nor U39925 (N_39925,N_35823,N_36166);
nor U39926 (N_39926,N_35129,N_35212);
or U39927 (N_39927,N_36008,N_36155);
nand U39928 (N_39928,N_35249,N_36159);
or U39929 (N_39929,N_37363,N_35299);
nor U39930 (N_39930,N_35492,N_36160);
xnor U39931 (N_39931,N_35165,N_35127);
nor U39932 (N_39932,N_37132,N_36156);
xnor U39933 (N_39933,N_36647,N_36061);
and U39934 (N_39934,N_35140,N_35526);
xnor U39935 (N_39935,N_36205,N_35655);
nand U39936 (N_39936,N_36730,N_36875);
or U39937 (N_39937,N_35541,N_35868);
nor U39938 (N_39938,N_36569,N_36610);
nand U39939 (N_39939,N_35702,N_37199);
or U39940 (N_39940,N_35839,N_36769);
xnor U39941 (N_39941,N_36657,N_35401);
and U39942 (N_39942,N_36689,N_36062);
nand U39943 (N_39943,N_36154,N_36679);
or U39944 (N_39944,N_37349,N_35569);
xor U39945 (N_39945,N_35110,N_36335);
nor U39946 (N_39946,N_37005,N_35508);
nand U39947 (N_39947,N_37470,N_36192);
xor U39948 (N_39948,N_36080,N_36523);
and U39949 (N_39949,N_35667,N_35607);
nand U39950 (N_39950,N_36293,N_35470);
nand U39951 (N_39951,N_35290,N_35145);
xnor U39952 (N_39952,N_36693,N_37187);
or U39953 (N_39953,N_35542,N_36822);
xor U39954 (N_39954,N_35614,N_35210);
and U39955 (N_39955,N_36352,N_36381);
nor U39956 (N_39956,N_36941,N_35533);
or U39957 (N_39957,N_35750,N_35405);
nand U39958 (N_39958,N_35178,N_36030);
nand U39959 (N_39959,N_35045,N_35529);
or U39960 (N_39960,N_35033,N_36388);
or U39961 (N_39961,N_35805,N_35867);
xor U39962 (N_39962,N_37075,N_36479);
nand U39963 (N_39963,N_36654,N_36505);
nand U39964 (N_39964,N_37079,N_36808);
xnor U39965 (N_39965,N_37338,N_36240);
nor U39966 (N_39966,N_37170,N_36572);
or U39967 (N_39967,N_37466,N_35725);
or U39968 (N_39968,N_37442,N_37345);
xnor U39969 (N_39969,N_36554,N_37455);
xor U39970 (N_39970,N_35311,N_36042);
xor U39971 (N_39971,N_36723,N_36260);
xor U39972 (N_39972,N_36060,N_35809);
and U39973 (N_39973,N_35129,N_37385);
or U39974 (N_39974,N_35151,N_35586);
xnor U39975 (N_39975,N_35894,N_36053);
or U39976 (N_39976,N_37250,N_35625);
or U39977 (N_39977,N_36897,N_35484);
and U39978 (N_39978,N_35408,N_35564);
xor U39979 (N_39979,N_35621,N_35636);
or U39980 (N_39980,N_35372,N_35581);
nand U39981 (N_39981,N_35356,N_35255);
and U39982 (N_39982,N_37361,N_36014);
xnor U39983 (N_39983,N_36233,N_35950);
xnor U39984 (N_39984,N_36091,N_36728);
nand U39985 (N_39985,N_36834,N_36699);
or U39986 (N_39986,N_35392,N_35868);
xor U39987 (N_39987,N_36347,N_36357);
nor U39988 (N_39988,N_36481,N_36751);
nor U39989 (N_39989,N_35613,N_36023);
or U39990 (N_39990,N_36098,N_35175);
nor U39991 (N_39991,N_35691,N_37286);
nor U39992 (N_39992,N_36905,N_35349);
xnor U39993 (N_39993,N_37025,N_37419);
nand U39994 (N_39994,N_37397,N_36005);
xnor U39995 (N_39995,N_37212,N_36235);
or U39996 (N_39996,N_35213,N_36952);
nand U39997 (N_39997,N_37278,N_35029);
nand U39998 (N_39998,N_35987,N_37228);
nor U39999 (N_39999,N_36772,N_37060);
and U40000 (N_40000,N_38286,N_39548);
nor U40001 (N_40001,N_37689,N_39152);
nand U40002 (N_40002,N_38902,N_38601);
or U40003 (N_40003,N_37926,N_39444);
or U40004 (N_40004,N_38125,N_37573);
or U40005 (N_40005,N_39991,N_39573);
or U40006 (N_40006,N_39655,N_38031);
and U40007 (N_40007,N_39463,N_39569);
xnor U40008 (N_40008,N_37835,N_38237);
xor U40009 (N_40009,N_37788,N_39098);
or U40010 (N_40010,N_39172,N_39176);
and U40011 (N_40011,N_39097,N_38927);
and U40012 (N_40012,N_38058,N_39439);
xnor U40013 (N_40013,N_39344,N_39681);
nand U40014 (N_40014,N_39337,N_39686);
and U40015 (N_40015,N_37622,N_37724);
nand U40016 (N_40016,N_39206,N_38807);
nand U40017 (N_40017,N_38828,N_37790);
and U40018 (N_40018,N_37894,N_39046);
xnor U40019 (N_40019,N_38270,N_37557);
or U40020 (N_40020,N_38189,N_37729);
nor U40021 (N_40021,N_39066,N_38208);
nand U40022 (N_40022,N_38103,N_37702);
nor U40023 (N_40023,N_38203,N_38509);
nor U40024 (N_40024,N_39519,N_39168);
and U40025 (N_40025,N_39404,N_39630);
or U40026 (N_40026,N_38401,N_39671);
nand U40027 (N_40027,N_39282,N_38488);
or U40028 (N_40028,N_38354,N_39131);
nand U40029 (N_40029,N_38374,N_38154);
xor U40030 (N_40030,N_38141,N_38428);
nand U40031 (N_40031,N_37753,N_38541);
and U40032 (N_40032,N_38216,N_39242);
and U40033 (N_40033,N_39722,N_39451);
xor U40034 (N_40034,N_38266,N_38117);
and U40035 (N_40035,N_39564,N_38258);
and U40036 (N_40036,N_38062,N_39657);
nor U40037 (N_40037,N_38242,N_38655);
and U40038 (N_40038,N_38340,N_39408);
xor U40039 (N_40039,N_39579,N_39759);
nor U40040 (N_40040,N_38914,N_39906);
nand U40041 (N_40041,N_37635,N_37990);
and U40042 (N_40042,N_38254,N_39852);
nand U40043 (N_40043,N_37881,N_37576);
and U40044 (N_40044,N_38558,N_37909);
or U40045 (N_40045,N_38214,N_38536);
xnor U40046 (N_40046,N_37644,N_38371);
or U40047 (N_40047,N_38943,N_37930);
and U40048 (N_40048,N_38947,N_39224);
xnor U40049 (N_40049,N_39266,N_39188);
or U40050 (N_40050,N_39043,N_39780);
nand U40051 (N_40051,N_38637,N_38710);
xor U40052 (N_40052,N_38368,N_37738);
xor U40053 (N_40053,N_38730,N_39236);
nor U40054 (N_40054,N_39788,N_39592);
xnor U40055 (N_40055,N_39520,N_38308);
or U40056 (N_40056,N_38511,N_38200);
or U40057 (N_40057,N_38457,N_38543);
or U40058 (N_40058,N_37558,N_38232);
xor U40059 (N_40059,N_39305,N_38301);
and U40060 (N_40060,N_38048,N_37817);
xnor U40061 (N_40061,N_37665,N_37799);
xnor U40062 (N_40062,N_38491,N_38339);
nand U40063 (N_40063,N_39644,N_38900);
or U40064 (N_40064,N_39695,N_37652);
nor U40065 (N_40065,N_37785,N_38496);
nand U40066 (N_40066,N_39434,N_38960);
and U40067 (N_40067,N_39534,N_38582);
xnor U40068 (N_40068,N_38768,N_38241);
and U40069 (N_40069,N_37810,N_39251);
or U40070 (N_40070,N_38223,N_39248);
nand U40071 (N_40071,N_37636,N_37821);
xnor U40072 (N_40072,N_39608,N_38656);
nor U40073 (N_40073,N_39900,N_39698);
nor U40074 (N_40074,N_37730,N_39894);
and U40075 (N_40075,N_39376,N_37651);
and U40076 (N_40076,N_39688,N_38672);
nand U40077 (N_40077,N_38813,N_39233);
and U40078 (N_40078,N_37687,N_39616);
xnor U40079 (N_40079,N_39058,N_37594);
nand U40080 (N_40080,N_39099,N_38338);
nor U40081 (N_40081,N_39627,N_39810);
nor U40082 (N_40082,N_37684,N_38573);
or U40083 (N_40083,N_38936,N_38461);
and U40084 (N_40084,N_39379,N_38941);
nor U40085 (N_40085,N_37543,N_37596);
xor U40086 (N_40086,N_37677,N_38318);
nor U40087 (N_40087,N_39632,N_38205);
nor U40088 (N_40088,N_38050,N_39317);
xor U40089 (N_40089,N_38613,N_38282);
nand U40090 (N_40090,N_38268,N_38877);
nor U40091 (N_40091,N_39737,N_38378);
xor U40092 (N_40092,N_37941,N_38029);
or U40093 (N_40093,N_39901,N_37893);
and U40094 (N_40094,N_39908,N_38448);
nand U40095 (N_40095,N_39403,N_38330);
xnor U40096 (N_40096,N_37640,N_37661);
nor U40097 (N_40097,N_39117,N_38278);
nor U40098 (N_40098,N_39565,N_37998);
xor U40099 (N_40099,N_39280,N_38086);
or U40100 (N_40100,N_39588,N_37546);
and U40101 (N_40101,N_38411,N_39457);
xnor U40102 (N_40102,N_37623,N_39801);
xor U40103 (N_40103,N_39499,N_37595);
nand U40104 (N_40104,N_38171,N_39890);
and U40105 (N_40105,N_37597,N_39405);
nor U40106 (N_40106,N_38105,N_39691);
xor U40107 (N_40107,N_38412,N_37505);
xor U40108 (N_40108,N_38122,N_38638);
and U40109 (N_40109,N_39760,N_38824);
nor U40110 (N_40110,N_39470,N_38003);
nor U40111 (N_40111,N_39709,N_37883);
nor U40112 (N_40112,N_39910,N_39307);
or U40113 (N_40113,N_39940,N_39541);
nor U40114 (N_40114,N_38722,N_38153);
xor U40115 (N_40115,N_39703,N_39443);
and U40116 (N_40116,N_39203,N_38968);
nand U40117 (N_40117,N_37890,N_39963);
nor U40118 (N_40118,N_38781,N_38024);
or U40119 (N_40119,N_38734,N_39334);
and U40120 (N_40120,N_39765,N_37732);
or U40121 (N_40121,N_38964,N_37554);
xnor U40122 (N_40122,N_38084,N_38745);
nand U40123 (N_40123,N_38539,N_39918);
xnor U40124 (N_40124,N_38429,N_39078);
nand U40125 (N_40125,N_39198,N_39298);
nand U40126 (N_40126,N_38665,N_39515);
nor U40127 (N_40127,N_38966,N_39621);
xnor U40128 (N_40128,N_37964,N_38791);
nand U40129 (N_40129,N_37737,N_37791);
xor U40130 (N_40130,N_39934,N_37559);
xnor U40131 (N_40131,N_38094,N_38102);
or U40132 (N_40132,N_37924,N_39063);
nand U40133 (N_40133,N_37736,N_38996);
nor U40134 (N_40134,N_39868,N_37939);
nor U40135 (N_40135,N_38377,N_38077);
and U40136 (N_40136,N_37787,N_37742);
and U40137 (N_40137,N_38139,N_38871);
xnor U40138 (N_40138,N_38147,N_38986);
or U40139 (N_40139,N_39779,N_39407);
nor U40140 (N_40140,N_39436,N_38167);
xnor U40141 (N_40141,N_39892,N_37647);
nor U40142 (N_40142,N_39882,N_38454);
nor U40143 (N_40143,N_38503,N_39297);
or U40144 (N_40144,N_38812,N_38227);
nand U40145 (N_40145,N_38880,N_37952);
xor U40146 (N_40146,N_37758,N_38856);
nand U40147 (N_40147,N_39818,N_39861);
nand U40148 (N_40148,N_39100,N_37776);
xnor U40149 (N_40149,N_39757,N_39150);
and U40150 (N_40150,N_38177,N_39835);
xnor U40151 (N_40151,N_39060,N_39729);
nor U40152 (N_40152,N_39239,N_38743);
xnor U40153 (N_40153,N_39002,N_38417);
nor U40154 (N_40154,N_39567,N_39799);
nand U40155 (N_40155,N_39108,N_38973);
nor U40156 (N_40156,N_39093,N_38149);
or U40157 (N_40157,N_39116,N_38303);
nand U40158 (N_40158,N_38551,N_39666);
or U40159 (N_40159,N_39185,N_37832);
and U40160 (N_40160,N_37733,N_38133);
and U40161 (N_40161,N_37720,N_39898);
or U40162 (N_40162,N_39178,N_39595);
xnor U40163 (N_40163,N_39241,N_39422);
and U40164 (N_40164,N_38479,N_39391);
nor U40165 (N_40165,N_39068,N_38486);
or U40166 (N_40166,N_39095,N_38328);
nand U40167 (N_40167,N_37931,N_37759);
and U40168 (N_40168,N_39535,N_39276);
nor U40169 (N_40169,N_38366,N_39025);
nor U40170 (N_40170,N_39701,N_38886);
xnor U40171 (N_40171,N_39028,N_39518);
nand U40172 (N_40172,N_39006,N_37726);
and U40173 (N_40173,N_37813,N_38349);
and U40174 (N_40174,N_39855,N_38035);
and U40175 (N_40175,N_39106,N_38938);
or U40176 (N_40176,N_38184,N_38562);
or U40177 (N_40177,N_38593,N_38172);
xor U40178 (N_40178,N_38175,N_39731);
or U40179 (N_40179,N_39381,N_38712);
and U40180 (N_40180,N_38118,N_38542);
and U40181 (N_40181,N_38921,N_38005);
or U40182 (N_40182,N_37691,N_37937);
xor U40183 (N_40183,N_39926,N_38383);
xnor U40184 (N_40184,N_38676,N_39157);
and U40185 (N_40185,N_37854,N_39950);
nand U40186 (N_40186,N_37534,N_39358);
nor U40187 (N_40187,N_39195,N_37980);
nor U40188 (N_40188,N_38212,N_38481);
or U40189 (N_40189,N_39888,N_39387);
xor U40190 (N_40190,N_37648,N_38207);
nor U40191 (N_40191,N_38793,N_38680);
nand U40192 (N_40192,N_39916,N_38641);
nor U40193 (N_40193,N_38083,N_38019);
or U40194 (N_40194,N_37946,N_38046);
nor U40195 (N_40195,N_39009,N_38956);
nor U40196 (N_40196,N_38778,N_38809);
and U40197 (N_40197,N_39400,N_38057);
and U40198 (N_40198,N_38399,N_39617);
nand U40199 (N_40199,N_37641,N_39245);
or U40200 (N_40200,N_38579,N_38723);
and U40201 (N_40201,N_37711,N_39393);
xnor U40202 (N_40202,N_37763,N_39817);
xnor U40203 (N_40203,N_38838,N_38524);
xor U40204 (N_40204,N_39672,N_38478);
and U40205 (N_40205,N_37805,N_39600);
nor U40206 (N_40206,N_39896,N_39807);
nor U40207 (N_40207,N_37802,N_39335);
and U40208 (N_40208,N_38231,N_37632);
nand U40209 (N_40209,N_39190,N_39969);
or U40210 (N_40210,N_38826,N_39478);
xnor U40211 (N_40211,N_37947,N_38449);
xor U40212 (N_40212,N_39736,N_38040);
or U40213 (N_40213,N_39111,N_38742);
and U40214 (N_40214,N_39746,N_37847);
nor U40215 (N_40215,N_38044,N_39215);
nand U40216 (N_40216,N_39732,N_38619);
and U40217 (N_40217,N_39545,N_38114);
nand U40218 (N_40218,N_37697,N_39530);
xor U40219 (N_40219,N_38480,N_37556);
nand U40220 (N_40220,N_37816,N_39210);
and U40221 (N_40221,N_37713,N_38953);
and U40222 (N_40222,N_39667,N_39255);
xnor U40223 (N_40223,N_38213,N_38160);
xor U40224 (N_40224,N_38857,N_39314);
xor U40225 (N_40225,N_39476,N_39883);
xor U40226 (N_40226,N_39915,N_37765);
and U40227 (N_40227,N_39464,N_38135);
and U40228 (N_40228,N_37960,N_39488);
and U40229 (N_40229,N_38991,N_38521);
nor U40230 (N_40230,N_39792,N_39547);
nand U40231 (N_40231,N_38894,N_39468);
or U40232 (N_40232,N_39889,N_39183);
or U40233 (N_40233,N_38054,N_37927);
nor U40234 (N_40234,N_38097,N_39073);
nor U40235 (N_40235,N_38132,N_38915);
nand U40236 (N_40236,N_39563,N_37916);
xor U40237 (N_40237,N_39762,N_38247);
nor U40238 (N_40238,N_38595,N_38563);
nor U40239 (N_40239,N_37510,N_38369);
nor U40240 (N_40240,N_38787,N_39312);
nand U40241 (N_40241,N_39555,N_38611);
nor U40242 (N_40242,N_38599,N_38930);
or U40243 (N_40243,N_38190,N_38990);
xor U40244 (N_40244,N_38711,N_37950);
and U40245 (N_40245,N_37585,N_38219);
nor U40246 (N_40246,N_39585,N_39811);
and U40247 (N_40247,N_39920,N_37656);
xor U40248 (N_40248,N_37629,N_38821);
xnor U40249 (N_40249,N_37542,N_39273);
nor U40250 (N_40250,N_39459,N_37806);
nor U40251 (N_40251,N_39808,N_38835);
nand U40252 (N_40252,N_39700,N_38884);
nand U40253 (N_40253,N_37545,N_39214);
and U40254 (N_40254,N_37852,N_38398);
nand U40255 (N_40255,N_39989,N_39955);
nor U40256 (N_40256,N_38113,N_37646);
xnor U40257 (N_40257,N_38289,N_39069);
and U40258 (N_40258,N_38037,N_38435);
nand U40259 (N_40259,N_39286,N_38673);
and U40260 (N_40260,N_37945,N_38143);
and U40261 (N_40261,N_39634,N_37925);
nand U40262 (N_40262,N_38156,N_38505);
or U40263 (N_40263,N_38586,N_37658);
xnor U40264 (N_40264,N_39951,N_38179);
and U40265 (N_40265,N_39885,N_39558);
and U40266 (N_40266,N_39664,N_38774);
xnor U40267 (N_40267,N_39952,N_39181);
nor U40268 (N_40268,N_39749,N_37589);
xnor U40269 (N_40269,N_39458,N_38780);
nor U40270 (N_40270,N_38287,N_39891);
xor U40271 (N_40271,N_37611,N_39511);
or U40272 (N_40272,N_39734,N_37675);
nand U40273 (N_40273,N_39872,N_39018);
xnor U40274 (N_40274,N_39831,N_39716);
nand U40275 (N_40275,N_38587,N_38136);
nand U40276 (N_40276,N_39213,N_39201);
xnor U40277 (N_40277,N_39847,N_39038);
and U40278 (N_40278,N_39495,N_37654);
nor U40279 (N_40279,N_38967,N_38014);
and U40280 (N_40280,N_37723,N_38713);
xnor U40281 (N_40281,N_39570,N_37511);
xor U40282 (N_40282,N_38001,N_38531);
xnor U40283 (N_40283,N_37562,N_37957);
xor U40284 (N_40284,N_38972,N_37696);
and U40285 (N_40285,N_39256,N_39284);
and U40286 (N_40286,N_37803,N_39294);
nor U40287 (N_40287,N_38333,N_37989);
xnor U40288 (N_40288,N_39359,N_38570);
nor U40289 (N_40289,N_39869,N_38121);
and U40290 (N_40290,N_38396,N_39089);
nand U40291 (N_40291,N_39650,N_37685);
nand U40292 (N_40292,N_38999,N_39202);
and U40293 (N_40293,N_38802,N_39557);
nand U40294 (N_40294,N_38830,N_38052);
nor U40295 (N_40295,N_37686,N_39954);
nor U40296 (N_40296,N_37746,N_39733);
and U40297 (N_40297,N_38684,N_38529);
or U40298 (N_40298,N_38937,N_39021);
nor U40299 (N_40299,N_38923,N_37915);
or U40300 (N_40300,N_39921,N_39037);
nor U40301 (N_40301,N_38294,N_39022);
or U40302 (N_40302,N_38332,N_38440);
nor U40303 (N_40303,N_39866,N_38111);
nand U40304 (N_40304,N_37988,N_37507);
and U40305 (N_40305,N_37750,N_38272);
nand U40306 (N_40306,N_37918,N_37764);
xnor U40307 (N_40307,N_39821,N_38544);
nor U40308 (N_40308,N_38720,N_38430);
nor U40309 (N_40309,N_39139,N_39005);
and U40310 (N_40310,N_39961,N_38145);
nor U40311 (N_40311,N_38410,N_38770);
nor U40312 (N_40312,N_39594,N_37517);
nand U40313 (N_40313,N_39979,N_38935);
nand U40314 (N_40314,N_39930,N_38861);
or U40315 (N_40315,N_38422,N_38316);
nor U40316 (N_40316,N_37602,N_39756);
and U40317 (N_40317,N_39079,N_38186);
and U40318 (N_40318,N_38931,N_37999);
nand U40319 (N_40319,N_38725,N_39309);
xnor U40320 (N_40320,N_38546,N_37780);
and U40321 (N_40321,N_37541,N_39141);
and U40322 (N_40322,N_38790,N_39936);
xnor U40323 (N_40323,N_38977,N_38854);
nand U40324 (N_40324,N_38648,N_38554);
and U40325 (N_40325,N_39755,N_38079);
and U40326 (N_40326,N_37800,N_39658);
and U40327 (N_40327,N_38439,N_38896);
xnor U40328 (N_40328,N_38547,N_37530);
and U40329 (N_40329,N_38092,N_39625);
nor U40330 (N_40330,N_38169,N_38307);
or U40331 (N_40331,N_39212,N_38578);
nand U40332 (N_40332,N_38253,N_37568);
xnor U40333 (N_40333,N_37638,N_38068);
nand U40334 (N_40334,N_39272,N_38737);
nand U40335 (N_40335,N_39626,N_37954);
xnor U40336 (N_40336,N_39708,N_38438);
xor U40337 (N_40337,N_39778,N_37895);
xor U40338 (N_40338,N_38998,N_38696);
nor U40339 (N_40339,N_37979,N_38682);
nor U40340 (N_40340,N_38564,N_39014);
and U40341 (N_40341,N_38834,N_38384);
xnor U40342 (N_40342,N_38668,N_39997);
nand U40343 (N_40343,N_38708,N_38388);
and U40344 (N_40344,N_39717,N_39836);
nor U40345 (N_40345,N_39635,N_38997);
nor U40346 (N_40346,N_38291,N_38016);
or U40347 (N_40347,N_39467,N_39207);
nor U40348 (N_40348,N_39240,N_37527);
nor U40349 (N_40349,N_38724,N_38251);
nand U40350 (N_40350,N_38581,N_38875);
nand U40351 (N_40351,N_38091,N_38633);
or U40352 (N_40352,N_39639,N_37688);
or U40353 (N_40353,N_38845,N_38859);
and U40354 (N_40354,N_37607,N_39502);
and U40355 (N_40355,N_38508,N_39745);
nor U40356 (N_40356,N_37565,N_39678);
nand U40357 (N_40357,N_37571,N_37995);
and U40358 (N_40358,N_37627,N_37624);
nor U40359 (N_40359,N_38277,N_39120);
and U40360 (N_40360,N_39124,N_39296);
xor U40361 (N_40361,N_39875,N_38043);
and U40362 (N_40362,N_38475,N_37560);
or U40363 (N_40363,N_39123,N_37819);
nor U40364 (N_40364,N_37712,N_39591);
nor U40365 (N_40365,N_39791,N_38335);
xnor U40366 (N_40366,N_38907,N_39707);
or U40367 (N_40367,N_39340,N_39016);
nand U40368 (N_40368,N_39365,N_38034);
or U40369 (N_40369,N_37886,N_38472);
nand U40370 (N_40370,N_37555,N_38313);
nand U40371 (N_40371,N_38522,N_39175);
nor U40372 (N_40372,N_38703,N_39143);
xnor U40373 (N_40373,N_39263,N_39132);
and U40374 (N_40374,N_39489,N_38550);
nand U40375 (N_40375,N_38965,N_39927);
and U40376 (N_40376,N_37929,N_39102);
and U40377 (N_40377,N_39076,N_38878);
nand U40378 (N_40378,N_38858,N_39786);
or U40379 (N_40379,N_38402,N_39170);
nor U40380 (N_40380,N_37717,N_39739);
xnor U40381 (N_40381,N_37523,N_39829);
or U40382 (N_40382,N_38514,N_38606);
xnor U40383 (N_40383,N_38948,N_37912);
and U40384 (N_40384,N_37981,N_39122);
nand U40385 (N_40385,N_39349,N_39113);
and U40386 (N_40386,N_38218,N_38453);
nand U40387 (N_40387,N_39867,N_38124);
or U40388 (N_40388,N_38685,N_39094);
or U40389 (N_40389,N_39506,N_37725);
nor U40390 (N_40390,N_39946,N_39411);
and U40391 (N_40391,N_39775,N_37754);
or U40392 (N_40392,N_39324,N_37872);
or U40393 (N_40393,N_39226,N_39730);
nor U40394 (N_40394,N_38882,N_38356);
nand U40395 (N_40395,N_38992,N_37705);
and U40396 (N_40396,N_37621,N_39290);
and U40397 (N_40397,N_38506,N_39781);
xnor U40398 (N_40398,N_37671,N_39956);
nor U40399 (N_40399,N_38913,N_39486);
or U40400 (N_40400,N_37827,N_39983);
and U40401 (N_40401,N_38650,N_39711);
nand U40402 (N_40402,N_39024,N_38653);
or U40403 (N_40403,N_39516,N_37578);
nand U40404 (N_40404,N_39192,N_39039);
xor U40405 (N_40405,N_38530,N_39372);
nand U40406 (N_40406,N_37707,N_39415);
nand U40407 (N_40407,N_39809,N_38958);
or U40408 (N_40408,N_37716,N_38721);
nor U40409 (N_40409,N_38089,N_39352);
xor U40410 (N_40410,N_39845,N_39250);
nand U40411 (N_40411,N_39554,N_39416);
or U40412 (N_40412,N_39684,N_38502);
nor U40413 (N_40413,N_39421,N_38825);
or U40414 (N_40414,N_37550,N_38863);
or U40415 (N_40415,N_38596,N_39738);
xnor U40416 (N_40416,N_37767,N_37868);
or U40417 (N_40417,N_39694,N_37959);
nand U40418 (N_40418,N_38959,N_39619);
nor U40419 (N_40419,N_39562,N_38718);
or U40420 (N_40420,N_38876,N_38074);
nand U40421 (N_40421,N_37681,N_37955);
nand U40422 (N_40422,N_38906,N_38686);
xor U40423 (N_40423,N_37653,N_38030);
nand U40424 (N_40424,N_37863,N_39720);
nand U40425 (N_40425,N_38018,N_37986);
xnor U40426 (N_40426,N_37903,N_37569);
nor U40427 (N_40427,N_39507,N_38702);
or U40428 (N_40428,N_39741,N_38138);
and U40429 (N_40429,N_37951,N_38687);
nand U40430 (N_40430,N_39289,N_39902);
xor U40431 (N_40431,N_39982,N_38252);
nor U40432 (N_40432,N_37612,N_37613);
nand U40433 (N_40433,N_39070,N_37631);
or U40434 (N_40434,N_38772,N_38362);
nand U40435 (N_40435,N_38591,N_38561);
or U40436 (N_40436,N_37516,N_39813);
nor U40437 (N_40437,N_38583,N_39453);
nor U40438 (N_40438,N_39494,N_37940);
and U40439 (N_40439,N_38612,N_38466);
xnor U40440 (N_40440,N_38783,N_39587);
nand U40441 (N_40441,N_37880,N_37783);
or U40442 (N_40442,N_39360,N_37958);
xnor U40443 (N_40443,N_39268,N_39366);
nand U40444 (N_40444,N_38257,N_38885);
nand U40445 (N_40445,N_38944,N_38452);
xnor U40446 (N_40446,N_37591,N_39010);
xor U40447 (N_40447,N_38654,N_38163);
nor U40448 (N_40448,N_39086,N_38413);
and U40449 (N_40449,N_38442,N_39269);
or U40450 (N_40450,N_39714,N_39689);
nand U40451 (N_40451,N_39523,N_39820);
xor U40452 (N_40452,N_39696,N_38173);
or U40453 (N_40453,N_37804,N_37798);
or U40454 (N_40454,N_39347,N_39649);
or U40455 (N_40455,N_39061,N_39114);
or U40456 (N_40456,N_39622,N_39794);
and U40457 (N_40457,N_37820,N_39493);
xor U40458 (N_40458,N_37823,N_38817);
nand U40459 (N_40459,N_37855,N_38071);
nand U40460 (N_40460,N_39677,N_39128);
and U40461 (N_40461,N_39399,N_38615);
or U40462 (N_40462,N_39465,N_39692);
or U40463 (N_40463,N_38928,N_39721);
nand U40464 (N_40464,N_38553,N_38098);
nand U40465 (N_40465,N_38495,N_38540);
or U40466 (N_40466,N_39367,N_39396);
nor U40467 (N_40467,N_38211,N_39370);
nor U40468 (N_40468,N_38385,N_38236);
or U40469 (N_40469,N_37683,N_39522);
or U40470 (N_40470,N_38848,N_37766);
xnor U40471 (N_40471,N_37769,N_38598);
and U40472 (N_40472,N_39321,N_37876);
or U40473 (N_40473,N_37949,N_38534);
or U40474 (N_40474,N_37610,N_39832);
nand U40475 (N_40475,N_39253,N_38533);
nand U40476 (N_40476,N_39110,N_38326);
nor U40477 (N_40477,N_38974,N_38933);
and U40478 (N_40478,N_39578,N_39645);
nor U40479 (N_40479,N_38315,N_37818);
and U40480 (N_40480,N_38299,N_38201);
xnor U40481 (N_40481,N_37659,N_39914);
nand U40482 (N_40482,N_38759,N_37825);
or U40483 (N_40483,N_39221,N_37660);
or U40484 (N_40484,N_38849,N_39851);
xor U40485 (N_40485,N_39085,N_38300);
nor U40486 (N_40486,N_38159,N_38441);
nand U40487 (N_40487,N_37966,N_39196);
or U40488 (N_40488,N_39235,N_39462);
or U40489 (N_40489,N_38357,N_38652);
or U40490 (N_40490,N_38647,N_37532);
nand U40491 (N_40491,N_39219,N_37864);
nand U40492 (N_40492,N_38467,N_38271);
and U40493 (N_40493,N_39001,N_38127);
and U40494 (N_40494,N_37572,N_39977);
xor U40495 (N_40495,N_39299,N_39750);
or U40496 (N_40496,N_37830,N_39763);
nand U40497 (N_40497,N_38951,N_38822);
xor U40498 (N_40498,N_39042,N_39537);
nor U40499 (N_40499,N_39310,N_39990);
nor U40500 (N_40500,N_38865,N_39204);
xor U40501 (N_40501,N_38419,N_39127);
or U40502 (N_40502,N_38447,N_39624);
or U40503 (N_40503,N_37809,N_39521);
nor U40504 (N_40504,N_39023,N_38889);
or U40505 (N_40505,N_38975,N_39052);
or U40506 (N_40506,N_38445,N_39074);
nor U40507 (N_40507,N_37972,N_37814);
nor U40508 (N_40508,N_38940,N_38850);
and U40509 (N_40509,N_38594,N_37928);
nand U40510 (N_40510,N_39169,N_39133);
nor U40511 (N_40511,N_38761,N_39968);
or U40512 (N_40512,N_38920,N_38843);
nand U40513 (N_40513,N_37526,N_37843);
and U40514 (N_40514,N_39897,N_38994);
nand U40515 (N_40515,N_39633,N_39841);
or U40516 (N_40516,N_37536,N_39662);
nor U40517 (N_40517,N_39880,N_37519);
nand U40518 (N_40518,N_38754,N_39602);
or U40519 (N_40519,N_37902,N_37842);
and U40520 (N_40520,N_38022,N_38238);
xnor U40521 (N_40521,N_37882,N_39998);
and U40522 (N_40522,N_37889,N_39432);
and U40523 (N_40523,N_39978,N_39611);
nor U40524 (N_40524,N_37792,N_39225);
xnor U40525 (N_40525,N_38883,N_38952);
nor U40526 (N_40526,N_38690,N_39425);
nor U40527 (N_40527,N_38181,N_37898);
nor U40528 (N_40528,N_39077,N_39917);
or U40529 (N_40529,N_39160,N_39173);
and U40530 (N_40530,N_37502,N_38283);
nor U40531 (N_40531,N_39540,N_39744);
nor U40532 (N_40532,N_39568,N_38304);
and U40533 (N_40533,N_38075,N_39995);
nor U40534 (N_40534,N_39665,N_39967);
and U40535 (N_40535,N_39531,N_38110);
and U40536 (N_40536,N_38851,N_37975);
nand U40537 (N_40537,N_38698,N_38777);
and U40538 (N_40538,N_38651,N_37588);
nand U40539 (N_40539,N_38617,N_37727);
nand U40540 (N_40540,N_39603,N_37503);
or U40541 (N_40541,N_38789,N_38414);
nand U40542 (N_40542,N_39062,N_38864);
or U40543 (N_40543,N_39830,N_38577);
or U40544 (N_40544,N_38771,N_39345);
and U40545 (N_40545,N_38285,N_37779);
and U40546 (N_40546,N_39966,N_38738);
nor U40547 (N_40547,N_37710,N_39121);
nand U40548 (N_40548,N_37528,N_39401);
nor U40549 (N_40549,N_37978,N_39208);
nor U40550 (N_40550,N_38246,N_37564);
or U40551 (N_40551,N_39267,N_38082);
and U40552 (N_40552,N_39812,N_38694);
nor U40553 (N_40553,N_38348,N_39939);
nor U40554 (N_40554,N_38455,N_39311);
or U40555 (N_40555,N_39142,N_39674);
and U40556 (N_40556,N_37693,N_39782);
xnor U40557 (N_40557,N_38166,N_37561);
and U40558 (N_40558,N_37748,N_38995);
xnor U40559 (N_40559,N_39389,N_39532);
and U40560 (N_40560,N_39613,N_39727);
and U40561 (N_40561,N_37781,N_38220);
xor U40562 (N_40562,N_38989,N_38629);
xnor U40563 (N_40563,N_39975,N_37761);
or U40564 (N_40564,N_38255,N_39096);
or U40565 (N_40565,N_38164,N_37603);
and U40566 (N_40566,N_38642,N_38939);
or U40567 (N_40567,N_39394,N_39673);
nand U40568 (N_40568,N_39774,N_37551);
xor U40569 (N_40569,N_39580,N_37633);
and U40570 (N_40570,N_37795,N_38187);
and U40571 (N_40571,N_38380,N_39261);
or U40572 (N_40572,N_38460,N_37695);
xnor U40573 (N_40573,N_38752,N_39285);
and U40574 (N_40574,N_38833,N_38027);
or U40575 (N_40575,N_39996,N_38233);
and U40576 (N_40576,N_37600,N_39217);
or U40577 (N_40577,N_39125,N_38726);
nor U40578 (N_40578,N_38222,N_39824);
nand U40579 (N_40579,N_38130,N_39319);
or U40580 (N_40580,N_38729,N_39980);
nor U40581 (N_40581,N_39450,N_39984);
nor U40582 (N_40582,N_39252,N_39838);
xnor U40583 (N_40583,N_38060,N_38779);
xnor U40584 (N_40584,N_37662,N_39825);
nor U40585 (N_40585,N_38662,N_37812);
nor U40586 (N_40586,N_38235,N_39923);
and U40587 (N_40587,N_38059,N_37811);
nor U40588 (N_40588,N_39767,N_39469);
and U40589 (N_40589,N_38134,N_39533);
or U40590 (N_40590,N_39262,N_39406);
nor U40591 (N_40591,N_39232,N_39572);
xnor U40592 (N_40592,N_37581,N_38017);
or U40593 (N_40593,N_39332,N_39377);
nor U40594 (N_40594,N_38717,N_37772);
xor U40595 (N_40595,N_39275,N_37645);
xor U40596 (N_40596,N_39246,N_39743);
nand U40597 (N_40597,N_38887,N_39712);
nor U40598 (N_40598,N_39785,N_38855);
xnor U40599 (N_40599,N_38226,N_37857);
and U40600 (N_40600,N_38010,N_38576);
xor U40601 (N_40601,N_38548,N_39287);
and U40602 (N_40602,N_38667,N_37922);
and U40603 (N_40603,N_39690,N_38263);
nor U40604 (N_40604,N_39937,N_39596);
or U40605 (N_40605,N_37948,N_39859);
and U40606 (N_40606,N_38757,N_39773);
xor U40607 (N_40607,N_38185,N_38312);
or U40608 (N_40608,N_37752,N_37749);
nor U40609 (N_40609,N_39107,N_38012);
and U40610 (N_40610,N_39471,N_38618);
nand U40611 (N_40611,N_39472,N_38093);
and U40612 (N_40612,N_39856,N_39822);
nand U40613 (N_40613,N_39485,N_38191);
and U40614 (N_40614,N_38784,N_37982);
or U40615 (N_40615,N_37642,N_39816);
nor U40616 (N_40616,N_39374,N_39414);
nor U40617 (N_40617,N_38917,N_38969);
nor U40618 (N_40618,N_39036,N_39147);
or U40619 (N_40619,N_39402,N_37877);
or U40620 (N_40620,N_39566,N_38101);
xnor U40621 (N_40621,N_37782,N_38565);
or U40622 (N_40622,N_38510,N_39041);
nand U40623 (N_40623,N_38776,N_37614);
nor U40624 (N_40624,N_39970,N_39620);
or U40625 (N_40625,N_39259,N_39227);
or U40626 (N_40626,N_38107,N_37694);
and U40627 (N_40627,N_39191,N_37896);
and U40628 (N_40628,N_38217,N_39965);
nand U40629 (N_40629,N_38336,N_39959);
xor U40630 (N_40630,N_37878,N_38142);
xor U40631 (N_40631,N_39390,N_39539);
nor U40632 (N_40632,N_37910,N_38644);
and U40633 (N_40633,N_37971,N_37728);
nor U40634 (N_40634,N_37608,N_39230);
or U40635 (N_40635,N_38080,N_38585);
and U40636 (N_40636,N_39597,N_39103);
or U40637 (N_40637,N_38128,N_39800);
nand U40638 (N_40638,N_38425,N_38785);
xor U40639 (N_40639,N_38204,N_38640);
nor U40640 (N_40640,N_39336,N_38750);
and U40641 (N_40641,N_38926,N_37598);
or U40642 (N_40642,N_38026,N_38262);
and U40643 (N_40643,N_37848,N_37770);
nand U40644 (N_40644,N_38344,N_39544);
and U40645 (N_40645,N_38535,N_39895);
xor U40646 (N_40646,N_38358,N_38700);
and U40647 (N_40647,N_38056,N_39949);
nand U40648 (N_40648,N_37859,N_39487);
nor U40649 (N_40649,N_39960,N_39753);
and U40650 (N_40650,N_39091,N_39618);
xor U40651 (N_40651,N_39064,N_38727);
nor U40652 (N_40652,N_37703,N_39683);
and U40653 (N_40653,N_38451,N_38567);
nand U40654 (N_40654,N_38746,N_39322);
or U40655 (N_40655,N_38516,N_39543);
or U40656 (N_40656,N_39477,N_39162);
xor U40657 (N_40657,N_37906,N_39482);
nor U40658 (N_40658,N_38273,N_38760);
nand U40659 (N_40659,N_37721,N_38007);
nor U40660 (N_40660,N_39084,N_38608);
nor U40661 (N_40661,N_37773,N_38494);
xor U40662 (N_40662,N_38621,N_37888);
nor U40663 (N_40663,N_38047,N_39805);
and U40664 (N_40664,N_38275,N_37649);
and U40665 (N_40665,N_38195,N_38331);
nor U40666 (N_40666,N_38028,N_39642);
xor U40667 (N_40667,N_39333,N_37865);
or U40668 (N_40668,N_38626,N_37682);
and U40669 (N_40669,N_39161,N_39277);
nor U40670 (N_40670,N_38804,N_38070);
nor U40671 (N_40671,N_39601,N_38327);
or U40672 (N_40672,N_38363,N_38244);
nor U40673 (N_40673,N_38515,N_37994);
nand U40674 (N_40674,N_38376,N_38692);
nand U40675 (N_40675,N_38061,N_38984);
xor U40676 (N_40676,N_39197,N_38256);
and U40677 (N_40677,N_37709,N_39873);
or U40678 (N_40678,N_37796,N_37789);
nand U40679 (N_40679,N_38170,N_38697);
nor U40680 (N_40680,N_38786,N_38297);
nand U40681 (N_40681,N_39303,N_38847);
xor U40682 (N_40682,N_38837,N_38078);
xor U40683 (N_40683,N_37501,N_39031);
or U40684 (N_40684,N_39101,N_38881);
nor U40685 (N_40685,N_39826,N_37911);
xnor U40686 (N_40686,N_39607,N_38085);
nand U40687 (N_40687,N_39180,N_39104);
and U40688 (N_40688,N_39274,N_38660);
nand U40689 (N_40689,N_39135,N_38627);
and U40690 (N_40690,N_38182,N_38867);
xnor U40691 (N_40691,N_39527,N_39879);
and U40692 (N_40692,N_37664,N_38706);
and U40693 (N_40693,N_38683,N_37839);
xnor U40694 (N_40694,N_39151,N_38735);
xor U40695 (N_40695,N_38259,N_39860);
or U40696 (N_40696,N_38814,N_39905);
nand U40697 (N_40697,N_38773,N_39584);
xnor U40698 (N_40698,N_39247,N_37768);
xor U40699 (N_40699,N_38674,N_37917);
nor U40700 (N_40700,N_38088,N_37897);
and U40701 (N_40701,N_39935,N_39420);
or U40702 (N_40702,N_38903,N_38351);
nor U40703 (N_40703,N_38526,N_37815);
nand U40704 (N_40704,N_37735,N_39526);
or U40705 (N_40705,N_38193,N_38707);
xor U40706 (N_40706,N_39348,N_39735);
nor U40707 (N_40707,N_37666,N_38609);
xor U40708 (N_40708,N_39976,N_37574);
nand U40709 (N_40709,N_39065,N_39501);
or U40710 (N_40710,N_38749,N_37875);
or U40711 (N_40711,N_37985,N_37838);
nand U40712 (N_40712,N_39265,N_39492);
and U40713 (N_40713,N_39363,N_39382);
and U40714 (N_40714,N_39943,N_39281);
or U40715 (N_40715,N_37657,N_39300);
nor U40716 (N_40716,N_38387,N_38279);
and U40717 (N_40717,N_37549,N_37833);
or U40718 (N_40718,N_37871,N_39140);
xor U40719 (N_40719,N_37740,N_38350);
or U40720 (N_40720,N_39449,N_39030);
nor U40721 (N_40721,N_38635,N_38055);
xnor U40722 (N_40722,N_39839,N_37606);
nor U40723 (N_40723,N_38347,N_39035);
nand U40724 (N_40724,N_39136,N_38805);
nor U40725 (N_40725,N_38893,N_37892);
nand U40726 (N_40726,N_39497,N_38473);
or U40727 (N_40727,N_39675,N_37921);
nand U40728 (N_40728,N_37967,N_39638);
nand U40729 (N_40729,N_38891,N_39491);
or U40730 (N_40730,N_39166,N_38073);
nand U40731 (N_40731,N_38919,N_39876);
or U40732 (N_40732,N_38605,N_38065);
nand U40733 (N_40733,N_38924,N_37637);
xor U40734 (N_40734,N_38239,N_38215);
nand U40735 (N_40735,N_38245,N_39392);
nand U40736 (N_40736,N_39454,N_39747);
or U40737 (N_40737,N_39159,N_39342);
nor U40738 (N_40738,N_38643,N_39699);
and U40739 (N_40739,N_37885,N_38614);
or U40740 (N_40740,N_37913,N_39517);
xnor U40741 (N_40741,N_39609,N_39292);
xor U40742 (N_40742,N_38980,N_38688);
xnor U40743 (N_40743,N_39629,N_38311);
nor U40744 (N_40744,N_37953,N_37734);
xnor U40745 (N_40745,N_38504,N_39015);
and U40746 (N_40746,N_39631,N_38015);
and U40747 (N_40747,N_39440,N_38574);
nand U40748 (N_40748,N_38391,N_39445);
xnor U40749 (N_40749,N_39985,N_37757);
xor U40750 (N_40750,N_38150,N_38569);
xor U40751 (N_40751,N_39051,N_39270);
xor U40752 (N_40752,N_39524,N_37668);
nand U40753 (N_40753,N_39291,N_38459);
or U40754 (N_40754,N_37617,N_38701);
or U40755 (N_40755,N_39668,N_37616);
or U40756 (N_40756,N_38465,N_38152);
xnor U40757 (N_40757,N_38261,N_37655);
nor U40758 (N_40758,N_39479,N_38892);
and U40759 (N_40759,N_39509,N_37643);
nand U40760 (N_40760,N_38744,N_37879);
nand U40761 (N_40761,N_38584,N_39325);
nand U40762 (N_40762,N_38600,N_39182);
or U40763 (N_40763,N_38538,N_39827);
nor U40764 (N_40764,N_38288,N_37563);
or U40765 (N_40765,N_38832,N_39412);
or U40766 (N_40766,N_39048,N_39538);
nand U40767 (N_40767,N_38359,N_38677);
xnor U40768 (N_40768,N_38963,N_37582);
nand U40769 (N_40769,N_38069,N_38909);
or U40770 (N_40770,N_37943,N_37731);
xor U40771 (N_40771,N_39109,N_39082);
nand U40772 (N_40772,N_38860,N_37680);
or U40773 (N_40773,N_38306,N_38545);
nor U40774 (N_40774,N_38305,N_37824);
or U40775 (N_40775,N_37836,N_38981);
or U40776 (N_40776,N_39798,N_37933);
nor U40777 (N_40777,N_39442,N_39080);
xnor U40778 (N_40778,N_39490,N_38168);
or U40779 (N_40779,N_38115,N_37521);
nand U40780 (N_40780,N_37539,N_39770);
nor U40781 (N_40781,N_39766,N_38829);
xor U40782 (N_40782,N_38831,N_39874);
or U40783 (N_40783,N_39636,N_39870);
nand U40784 (N_40784,N_39819,N_37866);
or U40785 (N_40785,N_39907,N_38487);
and U40786 (N_40786,N_38794,N_39862);
or U40787 (N_40787,N_39599,N_39713);
nand U40788 (N_40788,N_39549,N_39346);
xor U40789 (N_40789,N_38590,N_38020);
and U40790 (N_40790,N_39508,N_39228);
nand U40791 (N_40791,N_38950,N_39158);
nor U40792 (N_40792,N_38341,N_39008);
nor U40793 (N_40793,N_38632,N_39725);
nor U40794 (N_40794,N_38260,N_38610);
and U40795 (N_40795,N_37714,N_38280);
xnor U40796 (N_40796,N_37525,N_39571);
xnor U40797 (N_40797,N_38816,N_39368);
nand U40798 (N_40798,N_37584,N_37663);
and U40799 (N_40799,N_37961,N_38971);
and U40800 (N_40800,N_38431,N_38345);
nand U40801 (N_40801,N_37634,N_38693);
nor U40802 (N_40802,N_38418,N_38527);
and U40803 (N_40803,N_39848,N_38290);
nor U40804 (N_40804,N_39126,N_37700);
and U40805 (N_40805,N_38916,N_38728);
nand U40806 (N_40806,N_37579,N_39339);
and U40807 (N_40807,N_38955,N_39288);
nor U40808 (N_40808,N_39019,N_38798);
and U40809 (N_40809,N_39007,N_37938);
xor U40810 (N_40810,N_37669,N_38276);
or U40811 (N_40811,N_39962,N_39858);
xnor U40812 (N_40812,N_39724,N_39646);
nor U40813 (N_40813,N_38604,N_39987);
or U40814 (N_40814,N_39323,N_38630);
or U40815 (N_40815,N_38389,N_38842);
and U40816 (N_40816,N_37756,N_39112);
and U40817 (N_40817,N_39186,N_37900);
nor U40818 (N_40818,N_39410,N_39764);
nand U40819 (N_40819,N_38556,N_38450);
xor U40820 (N_40820,N_39119,N_37618);
or U40821 (N_40821,N_39912,N_37760);
and U40822 (N_40822,N_38839,N_39238);
nor U40823 (N_40823,N_37566,N_37508);
or U40824 (N_40824,N_37524,N_38620);
xor U40825 (N_40825,N_39849,N_39218);
xnor U40826 (N_40826,N_37874,N_39473);
nor U40827 (N_40827,N_39771,N_37977);
nand U40828 (N_40828,N_38753,N_38957);
and U40829 (N_40829,N_38571,N_37509);
nand U40830 (N_40830,N_38174,N_37580);
or U40831 (N_40831,N_39652,N_37755);
nand U40832 (N_40832,N_38379,N_37807);
nand U40833 (N_40833,N_38224,N_38866);
nor U40834 (N_40834,N_37547,N_39237);
nand U40835 (N_40835,N_38360,N_39947);
nor U40836 (N_40836,N_38493,N_38407);
xor U40837 (N_40837,N_38658,N_38346);
nor U40838 (N_40838,N_37849,N_39209);
nand U40839 (N_40839,N_38370,N_39331);
nor U40840 (N_40840,N_38819,N_38264);
nor U40841 (N_40841,N_38528,N_39304);
xnor U40842 (N_40842,N_39748,N_38393);
nor U40843 (N_40843,N_37590,N_38888);
xnor U40844 (N_40844,N_39220,N_39529);
xnor U40845 (N_40845,N_39075,N_38555);
nor U40846 (N_40846,N_39452,N_39092);
xor U40847 (N_40847,N_38497,N_39398);
nor U40848 (N_40848,N_39145,N_39004);
nor U40849 (N_40849,N_38364,N_38284);
or U40850 (N_40850,N_39815,N_38560);
nor U40851 (N_40851,N_38426,N_39040);
xnor U40852 (N_40852,N_38416,N_39842);
or U40853 (N_40853,N_39863,N_39167);
nand U40854 (N_40854,N_38373,N_38978);
xor U40855 (N_40855,N_38664,N_38188);
nand U40856 (N_40856,N_39351,N_39071);
xnor U40857 (N_40857,N_38468,N_38747);
or U40858 (N_40858,N_39758,N_39257);
nand U40859 (N_40859,N_38011,N_39615);
nand U40860 (N_40860,N_39981,N_38400);
or U40861 (N_40861,N_37784,N_37552);
and U40862 (N_40862,N_38557,N_38922);
and U40863 (N_40863,N_38045,N_37771);
nor U40864 (N_40864,N_38292,N_39355);
and U40865 (N_40865,N_38962,N_38053);
or U40866 (N_40866,N_38912,N_39542);
xor U40867 (N_40867,N_37974,N_37932);
or U40868 (N_40868,N_38532,N_38616);
nand U40869 (N_40869,N_39877,N_39661);
nor U40870 (N_40870,N_38549,N_38309);
and U40871 (N_40871,N_37905,N_38970);
nor U40872 (N_40872,N_39525,N_39751);
and U40873 (N_40873,N_39053,N_38987);
xor U40874 (N_40874,N_39423,N_39418);
or U40875 (N_40875,N_38979,N_38325);
xnor U40876 (N_40876,N_39293,N_38456);
nand U40877 (N_40877,N_38049,N_39814);
and U40878 (N_40878,N_38403,N_39715);
xnor U40879 (N_40879,N_39419,N_39789);
or U40880 (N_40880,N_38803,N_38229);
or U40881 (N_40881,N_39448,N_37869);
or U40882 (N_40882,N_39011,N_38386);
and U40883 (N_40883,N_37701,N_37997);
and U40884 (N_40884,N_37520,N_38230);
nand U40885 (N_40885,N_37920,N_37793);
xor U40886 (N_40886,N_39330,N_39857);
xor U40887 (N_40887,N_38799,N_37858);
or U40888 (N_40888,N_39553,N_39948);
nand U40889 (N_40889,N_39993,N_39430);
xnor U40890 (N_40890,N_39067,N_37544);
nor U40891 (N_40891,N_38552,N_38715);
nor U40892 (N_40892,N_39386,N_37786);
xor U40893 (N_40893,N_38976,N_39590);
nor U40894 (N_40894,N_37719,N_38006);
or U40895 (N_40895,N_37984,N_39222);
xor U40896 (N_40896,N_37867,N_39045);
or U40897 (N_40897,N_37944,N_39154);
or U40898 (N_40898,N_38736,N_38872);
and U40899 (N_40899,N_39806,N_39498);
nand U40900 (N_40900,N_38323,N_39582);
and U40901 (N_40901,N_39528,N_39971);
or U40902 (N_40902,N_38151,N_39424);
nor U40903 (N_40903,N_39886,N_39648);
nand U40904 (N_40904,N_38810,N_39027);
and U40905 (N_40905,N_38993,N_39144);
nand U40906 (N_40906,N_39364,N_37907);
xor U40907 (N_40907,N_37599,N_37775);
xnor U40908 (N_40908,N_38801,N_39205);
nand U40909 (N_40909,N_38039,N_39865);
or U40910 (N_40910,N_39433,N_38394);
nor U40911 (N_40911,N_39258,N_38372);
nor U40912 (N_40912,N_39397,N_38895);
xor U40913 (N_40913,N_37533,N_39474);
nand U40914 (N_40914,N_39787,N_39059);
or U40915 (N_40915,N_37515,N_39480);
nand U40916 (N_40916,N_38437,N_39054);
or U40917 (N_40917,N_37884,N_39719);
nor U40918 (N_40918,N_37739,N_37639);
or U40919 (N_40919,N_37699,N_37667);
xor U40920 (N_40920,N_39081,N_38404);
xnor U40921 (N_40921,N_37970,N_37856);
nand U40922 (N_40922,N_38146,N_38095);
nor U40923 (N_40923,N_38898,N_37822);
or U40924 (N_40924,N_38901,N_37605);
nor U40925 (N_40925,N_39932,N_39941);
nor U40926 (N_40926,N_37969,N_38293);
nor U40927 (N_40927,N_38659,N_39586);
or U40928 (N_40928,N_38423,N_38766);
xnor U40929 (N_40929,N_39843,N_39659);
and U40930 (N_40930,N_39654,N_37965);
nor U40931 (N_40931,N_38482,N_38076);
nand U40932 (N_40932,N_38890,N_39413);
or U40933 (N_40933,N_37592,N_39223);
and U40934 (N_40934,N_39384,N_37923);
or U40935 (N_40935,N_39313,N_37744);
nor U40936 (N_40936,N_38041,N_38741);
xnor U40937 (N_40937,N_38470,N_38732);
nor U40938 (N_40938,N_37993,N_39797);
nand U40939 (N_40939,N_39427,N_38714);
and U40940 (N_40940,N_38352,N_38806);
and U40941 (N_40941,N_39003,N_38397);
nor U40942 (N_40942,N_38126,N_39637);
and U40943 (N_40943,N_38324,N_38210);
nand U40944 (N_40944,N_38666,N_38225);
or U40945 (N_40945,N_38434,N_38334);
or U40946 (N_40946,N_39574,N_37673);
and U40947 (N_40947,N_39034,N_38298);
nor U40948 (N_40948,N_39680,N_39823);
nand U40949 (N_40949,N_37956,N_39740);
nand U40950 (N_40950,N_38274,N_39710);
nand U40951 (N_40951,N_39354,N_39466);
or U40952 (N_40952,N_38689,N_39957);
nand U40953 (N_40953,N_38733,N_37887);
and U40954 (N_40954,N_38490,N_39651);
nand U40955 (N_40955,N_38657,N_37936);
nand U40956 (N_40956,N_38296,N_38202);
and U40957 (N_40957,N_37531,N_39174);
nor U40958 (N_40958,N_38769,N_38704);
or U40959 (N_40959,N_39090,N_38982);
nor U40960 (N_40960,N_38961,N_38489);
or U40961 (N_40961,N_39020,N_38206);
nor U40962 (N_40962,N_38036,N_39254);
nor U40963 (N_40963,N_38954,N_39643);
nor U40964 (N_40964,N_37987,N_39243);
or U40965 (N_40965,N_38782,N_39575);
or U40966 (N_40966,N_38106,N_39598);
xor U40967 (N_40967,N_39833,N_38483);
nor U40968 (N_40968,N_37996,N_38432);
or U40969 (N_40969,N_38155,N_39922);
and U40970 (N_40970,N_38929,N_38628);
nor U40971 (N_40971,N_39784,N_38140);
or U40972 (N_40972,N_39706,N_38361);
and U40973 (N_40973,N_38178,N_38458);
xor U40974 (N_40974,N_39589,N_39925);
nor U40975 (N_40975,N_39362,N_39350);
and U40976 (N_40976,N_39864,N_38099);
nand U40977 (N_40977,N_37908,N_39149);
xor U40978 (N_40978,N_38507,N_39013);
nor U40979 (N_40979,N_39343,N_38795);
xor U40980 (N_40980,N_39795,N_39137);
or U40981 (N_40981,N_37840,N_39899);
or U40982 (N_40982,N_38661,N_39320);
nand U40983 (N_40983,N_38846,N_38870);
and U40984 (N_40984,N_38517,N_39083);
and U40985 (N_40985,N_37630,N_38474);
or U40986 (N_40986,N_39840,N_38165);
and U40987 (N_40987,N_39768,N_39904);
nor U40988 (N_40988,N_39193,N_39164);
nand U40989 (N_40989,N_38090,N_39105);
nand U40990 (N_40990,N_39606,N_37973);
nand U40991 (N_40991,N_37674,N_38671);
or U40992 (N_40992,N_39171,N_39295);
nand U40993 (N_40993,N_39187,N_39850);
or U40994 (N_40994,N_39118,N_39972);
or U40995 (N_40995,N_38249,N_38592);
xor U40996 (N_40996,N_37860,N_38910);
or U40997 (N_40997,N_37777,N_39044);
nor U40998 (N_40998,N_39560,N_38853);
xnor U40999 (N_40999,N_39844,N_39329);
and U41000 (N_41000,N_38319,N_38196);
nand U41001 (N_41001,N_38067,N_38751);
nand U41002 (N_41002,N_37718,N_39942);
nand U41003 (N_41003,N_37615,N_39887);
and U41004 (N_41004,N_39944,N_38183);
nor U41005 (N_41005,N_38691,N_39279);
or U41006 (N_41006,N_39153,N_37715);
nor U41007 (N_41007,N_38679,N_38112);
and U41008 (N_41008,N_39033,N_37548);
and U41009 (N_41009,N_39029,N_39994);
and U41010 (N_41010,N_39278,N_39878);
and U41011 (N_41011,N_38157,N_38607);
nand U41012 (N_41012,N_38123,N_37670);
nor U41013 (N_41013,N_38109,N_38267);
xnor U41014 (N_41014,N_39318,N_39338);
nand U41015 (N_41015,N_38575,N_39958);
nor U41016 (N_41016,N_38879,N_38949);
or U41017 (N_41017,N_37862,N_37829);
xor U41018 (N_41018,N_38815,N_39301);
nor U41019 (N_41019,N_39854,N_38827);
nand U41020 (N_41020,N_39610,N_37676);
xnor U41021 (N_41021,N_38932,N_37834);
or U41022 (N_41022,N_39371,N_37620);
and U41023 (N_41023,N_37976,N_38197);
or U41024 (N_41024,N_39426,N_37968);
nand U41025 (N_41025,N_38646,N_39115);
and U41026 (N_41026,N_39148,N_37540);
nand U41027 (N_41027,N_39853,N_38675);
xor U41028 (N_41028,N_38862,N_39000);
and U41029 (N_41029,N_38004,N_38897);
and U41030 (N_41030,N_37934,N_39697);
or U41031 (N_41031,N_38988,N_38874);
nand U41032 (N_41032,N_37801,N_39546);
nand U41033 (N_41033,N_38000,N_38634);
and U41034 (N_41034,N_38985,N_39628);
xor U41035 (N_41035,N_38580,N_38192);
nand U41036 (N_41036,N_37828,N_37570);
or U41037 (N_41037,N_38645,N_38705);
nand U41038 (N_41038,N_38678,N_38699);
and U41039 (N_41039,N_39496,N_39357);
nand U41040 (N_41040,N_38622,N_38463);
nand U41041 (N_41041,N_39380,N_39593);
or U41042 (N_41042,N_39561,N_39361);
or U41043 (N_41043,N_38281,N_38243);
and U41044 (N_41044,N_37518,N_39903);
and U41045 (N_41045,N_38365,N_38568);
nor U41046 (N_41046,N_37538,N_38382);
and U41047 (N_41047,N_38763,N_37762);
and U41048 (N_41048,N_39973,N_38087);
and U41049 (N_41049,N_38624,N_39660);
and U41050 (N_41050,N_37831,N_38537);
and U41051 (N_41051,N_38623,N_38137);
and U41052 (N_41052,N_37514,N_37963);
xor U41053 (N_41053,N_38844,N_38911);
or U41054 (N_41054,N_38096,N_38120);
or U41055 (N_41055,N_39802,N_39846);
or U41056 (N_41056,N_39327,N_39184);
xor U41057 (N_41057,N_37672,N_37851);
xor U41058 (N_41058,N_39679,N_38485);
nor U41059 (N_41059,N_38063,N_38484);
nand U41060 (N_41060,N_38589,N_39437);
nor U41061 (N_41061,N_37506,N_38424);
xor U41062 (N_41062,N_38797,N_39964);
or U41063 (N_41063,N_37891,N_38559);
xnor U41064 (N_41064,N_39356,N_38198);
nor U41065 (N_41065,N_38669,N_38443);
xor U41066 (N_41066,N_37794,N_38250);
xor U41067 (N_41067,N_38100,N_39234);
and U41068 (N_41068,N_39837,N_37942);
and U41069 (N_41069,N_37962,N_38023);
nand U41070 (N_41070,N_38572,N_39156);
nand U41071 (N_41071,N_38755,N_38462);
and U41072 (N_41072,N_38176,N_39481);
xor U41073 (N_41073,N_39138,N_38800);
xnor U41074 (N_41074,N_39718,N_39328);
and U41075 (N_41075,N_39988,N_38199);
nand U41076 (N_41076,N_38408,N_39244);
and U41077 (N_41077,N_38603,N_38209);
xnor U41078 (N_41078,N_38317,N_39913);
and U41079 (N_41079,N_39050,N_39032);
xnor U41080 (N_41080,N_38934,N_37797);
or U41081 (N_41081,N_38469,N_37722);
and U41082 (N_41082,N_39461,N_39460);
nor U41083 (N_41083,N_37826,N_37873);
or U41084 (N_41084,N_39828,N_38476);
xor U41085 (N_41085,N_38116,N_38228);
nor U41086 (N_41086,N_39056,N_37690);
or U41087 (N_41087,N_39012,N_39928);
and U41088 (N_41088,N_39163,N_38775);
xnor U41089 (N_41089,N_38946,N_38695);
nand U41090 (N_41090,N_37992,N_39428);
nor U41091 (N_41091,N_38840,N_39260);
nor U41092 (N_41092,N_38518,N_38329);
or U41093 (N_41093,N_39155,N_39656);
nand U41094 (N_41094,N_38739,N_38796);
xor U41095 (N_41095,N_38719,N_37850);
xor U41096 (N_41096,N_38421,N_39924);
or U41097 (N_41097,N_39306,N_38248);
or U41098 (N_41098,N_38108,N_39693);
xnor U41099 (N_41099,N_37692,N_38492);
nand U41100 (N_41100,N_38748,N_38756);
nand U41101 (N_41101,N_38355,N_38636);
xor U41102 (N_41102,N_37845,N_37747);
nor U41103 (N_41103,N_37628,N_39931);
and U41104 (N_41104,N_38716,N_39614);
xor U41105 (N_41105,N_38420,N_39026);
nor U41106 (N_41106,N_39088,N_39315);
and U41107 (N_41107,N_38983,N_39441);
and U41108 (N_41108,N_39369,N_39742);
nor U41109 (N_41109,N_38477,N_39938);
xor U41110 (N_41110,N_38367,N_39055);
xor U41111 (N_41111,N_39395,N_37935);
nor U41112 (N_41112,N_39429,N_38740);
and U41113 (N_41113,N_38836,N_39919);
xnor U41114 (N_41114,N_38194,N_39640);
nand U41115 (N_41115,N_38390,N_38823);
xnor U41116 (N_41116,N_39723,N_37751);
xor U41117 (N_41117,N_38663,N_39484);
nand U41118 (N_41118,N_37625,N_38523);
xor U41119 (N_41119,N_39353,N_39647);
or U41120 (N_41120,N_39500,N_38731);
or U41121 (N_41121,N_39456,N_37500);
nor U41122 (N_41122,N_37504,N_38588);
xnor U41123 (N_41123,N_37914,N_39375);
xor U41124 (N_41124,N_39676,N_37708);
nor U41125 (N_41125,N_39945,N_39881);
nand U41126 (N_41126,N_37586,N_38119);
nand U41127 (N_41127,N_38498,N_37583);
nand U41128 (N_41128,N_38148,N_38002);
or U41129 (N_41129,N_38234,N_39933);
xor U41130 (N_41130,N_38631,N_37853);
nand U41131 (N_41131,N_37861,N_37704);
and U41132 (N_41132,N_39049,N_38945);
nor U41133 (N_41133,N_39385,N_38161);
xor U41134 (N_41134,N_38295,N_37626);
xor U41135 (N_41135,N_39893,N_38602);
or U41136 (N_41136,N_38681,N_38269);
and U41137 (N_41137,N_39728,N_38158);
or U41138 (N_41138,N_39447,N_37678);
nand U41139 (N_41139,N_39388,N_39341);
nand U41140 (N_41140,N_38639,N_38265);
nand U41141 (N_41141,N_37741,N_39483);
xor U41142 (N_41142,N_38788,N_37513);
and U41143 (N_41143,N_37601,N_38409);
and U41144 (N_41144,N_39211,N_38765);
nor U41145 (N_41145,N_38767,N_38392);
or U41146 (N_41146,N_38021,N_38009);
and U41147 (N_41147,N_37650,N_38104);
and U41148 (N_41148,N_37983,N_38512);
nor U41149 (N_41149,N_37841,N_38008);
nor U41150 (N_41150,N_39177,N_38353);
nand U41151 (N_41151,N_38464,N_39704);
nand U41152 (N_41152,N_39834,N_39087);
or U41153 (N_41153,N_39682,N_37778);
and U41154 (N_41154,N_39551,N_39475);
or U41155 (N_41155,N_39641,N_38321);
xnor U41156 (N_41156,N_39200,N_39302);
or U41157 (N_41157,N_38918,N_37706);
or U41158 (N_41158,N_38525,N_38566);
nor U41159 (N_41159,N_39271,N_39783);
xor U41160 (N_41160,N_39803,N_39409);
and U41161 (N_41161,N_39772,N_37991);
xnor U41162 (N_41162,N_39612,N_39229);
nor U41163 (N_41163,N_38129,N_37844);
nor U41164 (N_41164,N_38899,N_38433);
nor U41165 (N_41165,N_38499,N_39326);
nor U41166 (N_41166,N_39754,N_39685);
xor U41167 (N_41167,N_39373,N_39911);
nand U41168 (N_41168,N_38427,N_37575);
xor U41169 (N_41169,N_38625,N_39455);
nor U41170 (N_41170,N_39999,N_38905);
or U41171 (N_41171,N_38500,N_39308);
nand U41172 (N_41172,N_39581,N_39796);
nand U41173 (N_41173,N_39130,N_38808);
or U41174 (N_41174,N_38405,N_39790);
nand U41175 (N_41175,N_37901,N_37535);
nand U41176 (N_41176,N_39583,N_39776);
or U41177 (N_41177,N_37837,N_38649);
nand U41178 (N_41178,N_39179,N_39417);
nand U41179 (N_41179,N_39804,N_37522);
nand U41180 (N_41180,N_38072,N_39446);
nor U41181 (N_41181,N_39536,N_37870);
nor U41182 (N_41182,N_38762,N_39669);
xor U41183 (N_41183,N_37743,N_39194);
and U41184 (N_41184,N_38501,N_39929);
nor U41185 (N_41185,N_37904,N_39653);
and U41186 (N_41186,N_39438,N_38709);
nand U41187 (N_41187,N_38314,N_38032);
and U41188 (N_41188,N_38162,N_38942);
or U41189 (N_41189,N_39992,N_39871);
or U41190 (N_41190,N_39761,N_38337);
xnor U41191 (N_41191,N_37698,N_39017);
and U41192 (N_41192,N_37619,N_39316);
or U41193 (N_41193,N_38852,N_37587);
or U41194 (N_41194,N_39769,N_38131);
or U41195 (N_41195,N_39504,N_39057);
xnor U41196 (N_41196,N_39556,N_38240);
xor U41197 (N_41197,N_38811,N_38033);
nor U41198 (N_41198,N_38869,N_39189);
xor U41199 (N_41199,N_38415,N_39072);
or U41200 (N_41200,N_39146,N_39510);
xnor U41201 (N_41201,N_37593,N_39777);
nor U41202 (N_41202,N_38081,N_37553);
nand U41203 (N_41203,N_38322,N_39047);
xnor U41204 (N_41204,N_39974,N_39687);
xor U41205 (N_41205,N_38051,N_38444);
xor U41206 (N_41206,N_39503,N_38520);
or U41207 (N_41207,N_38792,N_37609);
and U41208 (N_41208,N_39264,N_37846);
and U41209 (N_41209,N_38343,N_37567);
nor U41210 (N_41210,N_37899,N_38873);
nand U41211 (N_41211,N_39726,N_39702);
nand U41212 (N_41212,N_39909,N_39283);
nand U41213 (N_41213,N_38042,N_38320);
and U41214 (N_41214,N_39663,N_39513);
nand U41215 (N_41215,N_38670,N_38038);
xor U41216 (N_41216,N_39953,N_37529);
xor U41217 (N_41217,N_38310,N_39199);
and U41218 (N_41218,N_39559,N_39505);
nand U41219 (N_41219,N_39216,N_37679);
and U41220 (N_41220,N_37604,N_38868);
nor U41221 (N_41221,N_37537,N_38597);
or U41222 (N_41222,N_38925,N_38820);
or U41223 (N_41223,N_37919,N_38064);
xnor U41224 (N_41224,N_38904,N_39670);
and U41225 (N_41225,N_39552,N_38841);
and U41226 (N_41226,N_39435,N_38519);
nand U41227 (N_41227,N_38381,N_39623);
or U41228 (N_41228,N_38342,N_39605);
nand U41229 (N_41229,N_37774,N_37577);
nor U41230 (N_41230,N_38302,N_38375);
or U41231 (N_41231,N_39550,N_39705);
nand U41232 (N_41232,N_38013,N_39512);
nand U41233 (N_41233,N_39576,N_38471);
xnor U41234 (N_41234,N_39577,N_38025);
nor U41235 (N_41235,N_38406,N_39793);
nand U41236 (N_41236,N_39165,N_38395);
or U41237 (N_41237,N_39431,N_38818);
and U41238 (N_41238,N_38180,N_39383);
nand U41239 (N_41239,N_38446,N_37808);
or U41240 (N_41240,N_38513,N_37745);
nand U41241 (N_41241,N_39884,N_38758);
and U41242 (N_41242,N_39378,N_38908);
nand U41243 (N_41243,N_38066,N_39129);
nor U41244 (N_41244,N_39514,N_39231);
or U41245 (N_41245,N_38221,N_39249);
nor U41246 (N_41246,N_38764,N_39134);
nand U41247 (N_41247,N_37512,N_38144);
xnor U41248 (N_41248,N_39986,N_39604);
and U41249 (N_41249,N_39752,N_38436);
xnor U41250 (N_41250,N_38330,N_38941);
nor U41251 (N_41251,N_38094,N_39985);
xnor U41252 (N_41252,N_38272,N_38783);
xor U41253 (N_41253,N_38355,N_38747);
nand U41254 (N_41254,N_38522,N_37875);
xnor U41255 (N_41255,N_39384,N_38002);
or U41256 (N_41256,N_38046,N_38335);
nor U41257 (N_41257,N_38915,N_38457);
xnor U41258 (N_41258,N_38481,N_37524);
and U41259 (N_41259,N_39314,N_38185);
and U41260 (N_41260,N_38454,N_39920);
or U41261 (N_41261,N_38504,N_39945);
nand U41262 (N_41262,N_38422,N_39143);
and U41263 (N_41263,N_39632,N_38436);
and U41264 (N_41264,N_38498,N_39283);
and U41265 (N_41265,N_39751,N_39548);
or U41266 (N_41266,N_39878,N_39647);
xor U41267 (N_41267,N_37527,N_39324);
and U41268 (N_41268,N_39959,N_38833);
nand U41269 (N_41269,N_38309,N_38930);
or U41270 (N_41270,N_39432,N_39983);
and U41271 (N_41271,N_39165,N_38457);
and U41272 (N_41272,N_39245,N_37950);
or U41273 (N_41273,N_39279,N_38148);
or U41274 (N_41274,N_38721,N_39929);
nor U41275 (N_41275,N_38925,N_37585);
nand U41276 (N_41276,N_38260,N_39039);
xor U41277 (N_41277,N_38512,N_39373);
nand U41278 (N_41278,N_38420,N_37689);
or U41279 (N_41279,N_37627,N_38643);
and U41280 (N_41280,N_38977,N_39796);
and U41281 (N_41281,N_39392,N_38835);
and U41282 (N_41282,N_39550,N_38004);
nand U41283 (N_41283,N_39795,N_37574);
and U41284 (N_41284,N_39887,N_39442);
and U41285 (N_41285,N_37577,N_38734);
xnor U41286 (N_41286,N_38304,N_38265);
xor U41287 (N_41287,N_39209,N_38090);
nor U41288 (N_41288,N_39842,N_38152);
xnor U41289 (N_41289,N_38498,N_38879);
and U41290 (N_41290,N_37529,N_39180);
xor U41291 (N_41291,N_38628,N_39050);
xnor U41292 (N_41292,N_39520,N_39219);
and U41293 (N_41293,N_38006,N_37817);
xnor U41294 (N_41294,N_39256,N_38532);
nor U41295 (N_41295,N_39322,N_39291);
nand U41296 (N_41296,N_39876,N_37632);
or U41297 (N_41297,N_38982,N_39086);
xnor U41298 (N_41298,N_38689,N_37520);
xor U41299 (N_41299,N_39138,N_39123);
or U41300 (N_41300,N_37815,N_38694);
nor U41301 (N_41301,N_38906,N_38750);
and U41302 (N_41302,N_39591,N_38869);
or U41303 (N_41303,N_39494,N_38512);
and U41304 (N_41304,N_38090,N_37529);
nor U41305 (N_41305,N_39458,N_38509);
xor U41306 (N_41306,N_39743,N_39167);
nor U41307 (N_41307,N_39905,N_38031);
xor U41308 (N_41308,N_37627,N_39526);
nand U41309 (N_41309,N_39463,N_38442);
nand U41310 (N_41310,N_38101,N_39122);
nor U41311 (N_41311,N_38424,N_38202);
or U41312 (N_41312,N_38025,N_39030);
nor U41313 (N_41313,N_37533,N_38638);
and U41314 (N_41314,N_39039,N_37981);
xnor U41315 (N_41315,N_37962,N_39810);
nor U41316 (N_41316,N_39245,N_38036);
xnor U41317 (N_41317,N_39601,N_39895);
or U41318 (N_41318,N_38539,N_37649);
nand U41319 (N_41319,N_37747,N_39868);
nand U41320 (N_41320,N_38350,N_39194);
and U41321 (N_41321,N_39564,N_39800);
nand U41322 (N_41322,N_39233,N_38097);
nand U41323 (N_41323,N_39566,N_39211);
or U41324 (N_41324,N_37585,N_38591);
or U41325 (N_41325,N_38316,N_38729);
and U41326 (N_41326,N_39823,N_37809);
nor U41327 (N_41327,N_39844,N_39112);
and U41328 (N_41328,N_38438,N_37795);
xor U41329 (N_41329,N_38231,N_39345);
and U41330 (N_41330,N_37984,N_38439);
and U41331 (N_41331,N_39466,N_38928);
xor U41332 (N_41332,N_39863,N_37696);
nand U41333 (N_41333,N_39238,N_38341);
nand U41334 (N_41334,N_39019,N_38832);
nand U41335 (N_41335,N_39839,N_39579);
xor U41336 (N_41336,N_39468,N_38426);
nand U41337 (N_41337,N_38737,N_39558);
nor U41338 (N_41338,N_39027,N_37883);
and U41339 (N_41339,N_39073,N_39199);
nor U41340 (N_41340,N_38005,N_39579);
nor U41341 (N_41341,N_37683,N_38180);
xnor U41342 (N_41342,N_39609,N_39643);
or U41343 (N_41343,N_37933,N_37839);
nand U41344 (N_41344,N_37656,N_38846);
or U41345 (N_41345,N_38669,N_39791);
or U41346 (N_41346,N_37694,N_37753);
or U41347 (N_41347,N_38093,N_39737);
xor U41348 (N_41348,N_39269,N_38215);
and U41349 (N_41349,N_39384,N_38831);
nand U41350 (N_41350,N_39368,N_39246);
nor U41351 (N_41351,N_39832,N_38889);
nand U41352 (N_41352,N_37996,N_38362);
xor U41353 (N_41353,N_39311,N_39281);
or U41354 (N_41354,N_38819,N_39104);
nor U41355 (N_41355,N_39118,N_37723);
xor U41356 (N_41356,N_37679,N_39615);
nor U41357 (N_41357,N_37827,N_37741);
xnor U41358 (N_41358,N_38935,N_39625);
xnor U41359 (N_41359,N_39792,N_37521);
nand U41360 (N_41360,N_38375,N_39982);
xor U41361 (N_41361,N_38318,N_38017);
nand U41362 (N_41362,N_38505,N_37617);
xnor U41363 (N_41363,N_39620,N_39148);
xnor U41364 (N_41364,N_37781,N_39033);
nor U41365 (N_41365,N_39329,N_38953);
nor U41366 (N_41366,N_38746,N_39632);
and U41367 (N_41367,N_39909,N_39359);
xnor U41368 (N_41368,N_39675,N_37825);
xnor U41369 (N_41369,N_38131,N_38828);
nor U41370 (N_41370,N_39216,N_37730);
nand U41371 (N_41371,N_37925,N_39732);
xnor U41372 (N_41372,N_39856,N_37944);
xnor U41373 (N_41373,N_38110,N_39371);
nand U41374 (N_41374,N_39483,N_39724);
or U41375 (N_41375,N_39315,N_38805);
and U41376 (N_41376,N_37871,N_39859);
xor U41377 (N_41377,N_37718,N_39346);
and U41378 (N_41378,N_37600,N_38821);
and U41379 (N_41379,N_38472,N_38387);
and U41380 (N_41380,N_38432,N_39860);
or U41381 (N_41381,N_38743,N_39112);
nand U41382 (N_41382,N_39862,N_38315);
nand U41383 (N_41383,N_37956,N_39819);
xor U41384 (N_41384,N_39920,N_38182);
nor U41385 (N_41385,N_39107,N_39659);
nand U41386 (N_41386,N_38147,N_38769);
and U41387 (N_41387,N_37715,N_38798);
nand U41388 (N_41388,N_39264,N_39093);
xnor U41389 (N_41389,N_39310,N_37549);
nor U41390 (N_41390,N_39788,N_37806);
xor U41391 (N_41391,N_38555,N_37826);
nand U41392 (N_41392,N_37959,N_38305);
nand U41393 (N_41393,N_37551,N_38221);
nor U41394 (N_41394,N_37653,N_38622);
nand U41395 (N_41395,N_38010,N_39858);
xnor U41396 (N_41396,N_37868,N_37663);
nor U41397 (N_41397,N_39788,N_38671);
nand U41398 (N_41398,N_37735,N_38003);
or U41399 (N_41399,N_38819,N_38170);
nand U41400 (N_41400,N_39119,N_38535);
xor U41401 (N_41401,N_38229,N_39313);
nand U41402 (N_41402,N_37595,N_37509);
or U41403 (N_41403,N_39810,N_38945);
xnor U41404 (N_41404,N_38162,N_37902);
or U41405 (N_41405,N_39244,N_38700);
xor U41406 (N_41406,N_39346,N_38411);
and U41407 (N_41407,N_38198,N_38409);
nor U41408 (N_41408,N_39903,N_39241);
xnor U41409 (N_41409,N_37598,N_39293);
xnor U41410 (N_41410,N_37508,N_39368);
or U41411 (N_41411,N_39932,N_37556);
xnor U41412 (N_41412,N_39338,N_37544);
and U41413 (N_41413,N_39080,N_38338);
nand U41414 (N_41414,N_37604,N_37896);
or U41415 (N_41415,N_38393,N_39614);
and U41416 (N_41416,N_39739,N_37667);
nor U41417 (N_41417,N_37829,N_37962);
xor U41418 (N_41418,N_39490,N_37549);
and U41419 (N_41419,N_38614,N_39441);
or U41420 (N_41420,N_39597,N_37807);
or U41421 (N_41421,N_38617,N_38174);
nand U41422 (N_41422,N_39866,N_39943);
xnor U41423 (N_41423,N_38247,N_39717);
and U41424 (N_41424,N_39695,N_38099);
and U41425 (N_41425,N_39588,N_37793);
nor U41426 (N_41426,N_38588,N_38698);
and U41427 (N_41427,N_39691,N_39531);
and U41428 (N_41428,N_38449,N_39829);
nand U41429 (N_41429,N_38638,N_37930);
and U41430 (N_41430,N_38192,N_38909);
xor U41431 (N_41431,N_37780,N_39678);
xnor U41432 (N_41432,N_38752,N_37697);
or U41433 (N_41433,N_39089,N_39662);
nor U41434 (N_41434,N_38632,N_39349);
nand U41435 (N_41435,N_38543,N_38273);
or U41436 (N_41436,N_37790,N_39139);
or U41437 (N_41437,N_39786,N_39993);
nor U41438 (N_41438,N_38725,N_37795);
xor U41439 (N_41439,N_38821,N_39147);
nor U41440 (N_41440,N_39659,N_39411);
nand U41441 (N_41441,N_39439,N_38625);
or U41442 (N_41442,N_38036,N_39186);
nor U41443 (N_41443,N_37880,N_38632);
or U41444 (N_41444,N_38041,N_38980);
xnor U41445 (N_41445,N_39635,N_37777);
nor U41446 (N_41446,N_38467,N_38922);
nand U41447 (N_41447,N_37962,N_38757);
and U41448 (N_41448,N_37755,N_37641);
and U41449 (N_41449,N_38518,N_39648);
nor U41450 (N_41450,N_39664,N_37932);
nor U41451 (N_41451,N_37939,N_38868);
xor U41452 (N_41452,N_38710,N_37652);
nor U41453 (N_41453,N_39155,N_39294);
xor U41454 (N_41454,N_39479,N_37591);
xnor U41455 (N_41455,N_37576,N_39143);
nand U41456 (N_41456,N_38390,N_39611);
nor U41457 (N_41457,N_39885,N_38526);
or U41458 (N_41458,N_38234,N_39314);
xnor U41459 (N_41459,N_39853,N_38349);
nor U41460 (N_41460,N_39068,N_39570);
nand U41461 (N_41461,N_39359,N_39066);
nor U41462 (N_41462,N_39915,N_39040);
xnor U41463 (N_41463,N_38758,N_37729);
or U41464 (N_41464,N_38891,N_37661);
xnor U41465 (N_41465,N_38664,N_39669);
nor U41466 (N_41466,N_37630,N_38707);
nor U41467 (N_41467,N_37827,N_39568);
nor U41468 (N_41468,N_37739,N_38452);
xor U41469 (N_41469,N_38137,N_39180);
and U41470 (N_41470,N_39308,N_37581);
nor U41471 (N_41471,N_39385,N_37621);
and U41472 (N_41472,N_37788,N_38530);
nand U41473 (N_41473,N_38211,N_38389);
nor U41474 (N_41474,N_38942,N_39370);
nand U41475 (N_41475,N_38540,N_39222);
or U41476 (N_41476,N_38044,N_37992);
xnor U41477 (N_41477,N_38434,N_37841);
and U41478 (N_41478,N_38926,N_38927);
nor U41479 (N_41479,N_38733,N_38009);
xor U41480 (N_41480,N_39771,N_39747);
xnor U41481 (N_41481,N_37750,N_38164);
and U41482 (N_41482,N_39320,N_38676);
nand U41483 (N_41483,N_39679,N_39822);
nand U41484 (N_41484,N_38203,N_38661);
or U41485 (N_41485,N_37542,N_38398);
xnor U41486 (N_41486,N_38975,N_38831);
or U41487 (N_41487,N_38031,N_38671);
or U41488 (N_41488,N_39233,N_37623);
nor U41489 (N_41489,N_39774,N_38302);
or U41490 (N_41490,N_38016,N_39538);
nor U41491 (N_41491,N_38360,N_38555);
and U41492 (N_41492,N_39224,N_39179);
and U41493 (N_41493,N_38508,N_39924);
and U41494 (N_41494,N_38268,N_39689);
and U41495 (N_41495,N_38437,N_37614);
nand U41496 (N_41496,N_39543,N_37975);
and U41497 (N_41497,N_37559,N_37535);
and U41498 (N_41498,N_39945,N_39025);
xor U41499 (N_41499,N_38790,N_38858);
nand U41500 (N_41500,N_38513,N_39867);
xnor U41501 (N_41501,N_38116,N_39973);
nand U41502 (N_41502,N_39602,N_39176);
nor U41503 (N_41503,N_38828,N_37675);
xnor U41504 (N_41504,N_37925,N_38100);
and U41505 (N_41505,N_37526,N_37758);
nor U41506 (N_41506,N_39984,N_39547);
or U41507 (N_41507,N_38379,N_39728);
or U41508 (N_41508,N_38345,N_38670);
or U41509 (N_41509,N_37617,N_38982);
xor U41510 (N_41510,N_39836,N_39901);
nor U41511 (N_41511,N_39121,N_39805);
nor U41512 (N_41512,N_39413,N_39370);
or U41513 (N_41513,N_37802,N_38224);
xnor U41514 (N_41514,N_38549,N_38987);
or U41515 (N_41515,N_37563,N_37953);
nand U41516 (N_41516,N_39882,N_39547);
xnor U41517 (N_41517,N_38651,N_38869);
nor U41518 (N_41518,N_39258,N_39396);
nor U41519 (N_41519,N_39920,N_38550);
xnor U41520 (N_41520,N_39591,N_38988);
xor U41521 (N_41521,N_39324,N_37776);
xnor U41522 (N_41522,N_39645,N_38401);
or U41523 (N_41523,N_38796,N_38403);
and U41524 (N_41524,N_37841,N_38957);
and U41525 (N_41525,N_39250,N_39929);
nor U41526 (N_41526,N_39920,N_38522);
or U41527 (N_41527,N_37652,N_39946);
and U41528 (N_41528,N_39536,N_39339);
or U41529 (N_41529,N_39534,N_39460);
nand U41530 (N_41530,N_39648,N_38097);
and U41531 (N_41531,N_39301,N_38323);
xnor U41532 (N_41532,N_37839,N_38204);
or U41533 (N_41533,N_38591,N_39030);
or U41534 (N_41534,N_38497,N_39204);
or U41535 (N_41535,N_38998,N_37935);
or U41536 (N_41536,N_38373,N_38747);
and U41537 (N_41537,N_38577,N_39085);
nor U41538 (N_41538,N_38446,N_37526);
xor U41539 (N_41539,N_39903,N_38644);
and U41540 (N_41540,N_37877,N_39825);
or U41541 (N_41541,N_37844,N_39440);
and U41542 (N_41542,N_37875,N_37825);
nor U41543 (N_41543,N_39915,N_38234);
and U41544 (N_41544,N_37622,N_38722);
nor U41545 (N_41545,N_37543,N_39269);
nand U41546 (N_41546,N_39223,N_39429);
xor U41547 (N_41547,N_38613,N_37553);
and U41548 (N_41548,N_38044,N_37603);
nand U41549 (N_41549,N_38925,N_39824);
and U41550 (N_41550,N_38099,N_39796);
and U41551 (N_41551,N_37751,N_38435);
nor U41552 (N_41552,N_39211,N_38024);
xor U41553 (N_41553,N_37885,N_39377);
nor U41554 (N_41554,N_37586,N_38546);
and U41555 (N_41555,N_38431,N_38715);
nor U41556 (N_41556,N_39079,N_37784);
nor U41557 (N_41557,N_39896,N_37771);
and U41558 (N_41558,N_38919,N_39523);
and U41559 (N_41559,N_37671,N_39679);
nor U41560 (N_41560,N_39498,N_39305);
or U41561 (N_41561,N_37705,N_39920);
xor U41562 (N_41562,N_37734,N_38095);
nor U41563 (N_41563,N_38357,N_39282);
or U41564 (N_41564,N_37528,N_39880);
nand U41565 (N_41565,N_39257,N_39826);
and U41566 (N_41566,N_39034,N_37800);
nand U41567 (N_41567,N_38849,N_38985);
nand U41568 (N_41568,N_37547,N_38635);
nand U41569 (N_41569,N_38321,N_39783);
or U41570 (N_41570,N_37883,N_38350);
nand U41571 (N_41571,N_38409,N_38822);
xor U41572 (N_41572,N_38185,N_38155);
xnor U41573 (N_41573,N_38853,N_37627);
xor U41574 (N_41574,N_39966,N_38578);
or U41575 (N_41575,N_37801,N_39765);
and U41576 (N_41576,N_37858,N_38763);
and U41577 (N_41577,N_39651,N_38604);
nor U41578 (N_41578,N_38520,N_38459);
or U41579 (N_41579,N_39886,N_38468);
xnor U41580 (N_41580,N_39791,N_37606);
nor U41581 (N_41581,N_37710,N_37573);
xnor U41582 (N_41582,N_38135,N_39454);
nand U41583 (N_41583,N_39264,N_37607);
and U41584 (N_41584,N_38773,N_38215);
or U41585 (N_41585,N_39564,N_38377);
and U41586 (N_41586,N_38547,N_37554);
xor U41587 (N_41587,N_37973,N_37617);
nor U41588 (N_41588,N_37823,N_37896);
nand U41589 (N_41589,N_39298,N_38436);
nor U41590 (N_41590,N_39231,N_38132);
xor U41591 (N_41591,N_37759,N_39833);
nor U41592 (N_41592,N_39437,N_38930);
nand U41593 (N_41593,N_39925,N_37848);
nor U41594 (N_41594,N_38157,N_39675);
nor U41595 (N_41595,N_37896,N_39407);
xor U41596 (N_41596,N_37746,N_38486);
nor U41597 (N_41597,N_38917,N_37951);
xor U41598 (N_41598,N_39480,N_38197);
nand U41599 (N_41599,N_39397,N_38210);
or U41600 (N_41600,N_39967,N_39673);
and U41601 (N_41601,N_38300,N_37918);
nand U41602 (N_41602,N_38764,N_38534);
and U41603 (N_41603,N_39069,N_39774);
and U41604 (N_41604,N_39841,N_39381);
xnor U41605 (N_41605,N_38342,N_39558);
nor U41606 (N_41606,N_39210,N_39232);
nor U41607 (N_41607,N_37924,N_38780);
or U41608 (N_41608,N_39213,N_39078);
xnor U41609 (N_41609,N_38775,N_38917);
nor U41610 (N_41610,N_37584,N_39003);
nor U41611 (N_41611,N_37646,N_37504);
nand U41612 (N_41612,N_39663,N_38531);
nand U41613 (N_41613,N_37936,N_39377);
nor U41614 (N_41614,N_38008,N_37810);
or U41615 (N_41615,N_38656,N_38864);
or U41616 (N_41616,N_39437,N_39992);
nor U41617 (N_41617,N_39613,N_39164);
and U41618 (N_41618,N_39027,N_38733);
nor U41619 (N_41619,N_38898,N_39437);
and U41620 (N_41620,N_37511,N_37917);
xnor U41621 (N_41621,N_38427,N_38641);
or U41622 (N_41622,N_38218,N_37861);
nand U41623 (N_41623,N_38760,N_39576);
xor U41624 (N_41624,N_38831,N_39512);
and U41625 (N_41625,N_38088,N_38152);
nor U41626 (N_41626,N_37845,N_38327);
nand U41627 (N_41627,N_39125,N_39433);
or U41628 (N_41628,N_38857,N_38495);
nand U41629 (N_41629,N_39737,N_38155);
and U41630 (N_41630,N_37629,N_38746);
xor U41631 (N_41631,N_38649,N_38242);
and U41632 (N_41632,N_38270,N_38057);
nor U41633 (N_41633,N_37573,N_39618);
or U41634 (N_41634,N_37535,N_39504);
or U41635 (N_41635,N_38445,N_39302);
or U41636 (N_41636,N_38588,N_38269);
and U41637 (N_41637,N_38655,N_38013);
xnor U41638 (N_41638,N_39855,N_38823);
nor U41639 (N_41639,N_39647,N_39722);
nand U41640 (N_41640,N_38171,N_39158);
and U41641 (N_41641,N_38689,N_38418);
nor U41642 (N_41642,N_37945,N_38252);
and U41643 (N_41643,N_38935,N_39087);
and U41644 (N_41644,N_39976,N_37850);
or U41645 (N_41645,N_37750,N_37657);
xnor U41646 (N_41646,N_38704,N_38096);
nor U41647 (N_41647,N_38169,N_39647);
and U41648 (N_41648,N_38835,N_39961);
nor U41649 (N_41649,N_39785,N_37516);
nor U41650 (N_41650,N_38739,N_39319);
nor U41651 (N_41651,N_39859,N_38254);
or U41652 (N_41652,N_37661,N_38654);
or U41653 (N_41653,N_37829,N_37710);
xnor U41654 (N_41654,N_38388,N_39690);
or U41655 (N_41655,N_39110,N_38195);
nor U41656 (N_41656,N_39243,N_39175);
xor U41657 (N_41657,N_39616,N_37578);
nor U41658 (N_41658,N_39315,N_38150);
nand U41659 (N_41659,N_38394,N_38759);
xnor U41660 (N_41660,N_38043,N_39925);
nand U41661 (N_41661,N_39170,N_38489);
nor U41662 (N_41662,N_38051,N_39659);
nor U41663 (N_41663,N_39945,N_39808);
or U41664 (N_41664,N_39508,N_37606);
nor U41665 (N_41665,N_39539,N_39008);
and U41666 (N_41666,N_39986,N_38248);
nand U41667 (N_41667,N_38439,N_38745);
or U41668 (N_41668,N_38191,N_39963);
nor U41669 (N_41669,N_37545,N_38317);
nand U41670 (N_41670,N_39498,N_37957);
or U41671 (N_41671,N_37598,N_39993);
or U41672 (N_41672,N_37709,N_39409);
nor U41673 (N_41673,N_37946,N_38161);
nand U41674 (N_41674,N_38112,N_37533);
and U41675 (N_41675,N_39077,N_39905);
xnor U41676 (N_41676,N_38205,N_39987);
nor U41677 (N_41677,N_39239,N_39222);
nor U41678 (N_41678,N_38285,N_38512);
xor U41679 (N_41679,N_39927,N_38647);
nand U41680 (N_41680,N_38538,N_39626);
and U41681 (N_41681,N_39537,N_38766);
or U41682 (N_41682,N_39431,N_39309);
nor U41683 (N_41683,N_38923,N_38609);
nand U41684 (N_41684,N_39478,N_38297);
and U41685 (N_41685,N_37597,N_38780);
xor U41686 (N_41686,N_38766,N_38556);
and U41687 (N_41687,N_37522,N_39065);
and U41688 (N_41688,N_39513,N_39127);
and U41689 (N_41689,N_39897,N_37840);
and U41690 (N_41690,N_37907,N_38942);
nor U41691 (N_41691,N_38592,N_39882);
nor U41692 (N_41692,N_38949,N_37967);
xnor U41693 (N_41693,N_38233,N_38689);
or U41694 (N_41694,N_38709,N_37792);
nand U41695 (N_41695,N_39095,N_37520);
and U41696 (N_41696,N_38698,N_39334);
or U41697 (N_41697,N_39255,N_37579);
nor U41698 (N_41698,N_39051,N_38839);
and U41699 (N_41699,N_38180,N_38283);
xnor U41700 (N_41700,N_38140,N_38729);
xor U41701 (N_41701,N_37923,N_37642);
xnor U41702 (N_41702,N_38765,N_37882);
nand U41703 (N_41703,N_37503,N_39026);
nand U41704 (N_41704,N_39330,N_39266);
nor U41705 (N_41705,N_37831,N_37852);
nand U41706 (N_41706,N_38553,N_38549);
or U41707 (N_41707,N_38843,N_38161);
and U41708 (N_41708,N_37624,N_37590);
and U41709 (N_41709,N_39983,N_38636);
nand U41710 (N_41710,N_38669,N_39740);
nand U41711 (N_41711,N_39490,N_37865);
xnor U41712 (N_41712,N_37967,N_37683);
nand U41713 (N_41713,N_39192,N_37507);
xnor U41714 (N_41714,N_37913,N_38263);
nor U41715 (N_41715,N_38965,N_37681);
or U41716 (N_41716,N_38069,N_38279);
nand U41717 (N_41717,N_37748,N_39838);
or U41718 (N_41718,N_39972,N_37500);
xor U41719 (N_41719,N_37822,N_39770);
xnor U41720 (N_41720,N_39503,N_37543);
or U41721 (N_41721,N_39658,N_38626);
or U41722 (N_41722,N_39195,N_37680);
or U41723 (N_41723,N_38164,N_39493);
nand U41724 (N_41724,N_38909,N_39514);
or U41725 (N_41725,N_39659,N_39758);
xnor U41726 (N_41726,N_38812,N_38399);
xor U41727 (N_41727,N_38289,N_38328);
xor U41728 (N_41728,N_39344,N_38352);
and U41729 (N_41729,N_38952,N_38603);
or U41730 (N_41730,N_39734,N_37532);
or U41731 (N_41731,N_38627,N_38750);
and U41732 (N_41732,N_38699,N_38365);
or U41733 (N_41733,N_39349,N_39312);
or U41734 (N_41734,N_37577,N_39000);
xnor U41735 (N_41735,N_39481,N_39294);
and U41736 (N_41736,N_39423,N_37872);
xor U41737 (N_41737,N_39635,N_39882);
xnor U41738 (N_41738,N_39065,N_39594);
or U41739 (N_41739,N_37926,N_37972);
or U41740 (N_41740,N_39666,N_38398);
or U41741 (N_41741,N_39650,N_39165);
nand U41742 (N_41742,N_37529,N_39959);
nor U41743 (N_41743,N_39970,N_38950);
or U41744 (N_41744,N_38886,N_38991);
nor U41745 (N_41745,N_39894,N_37745);
xor U41746 (N_41746,N_38271,N_38981);
xor U41747 (N_41747,N_39275,N_39717);
or U41748 (N_41748,N_39137,N_38355);
nand U41749 (N_41749,N_38877,N_39214);
nor U41750 (N_41750,N_39588,N_39994);
nand U41751 (N_41751,N_38053,N_38676);
and U41752 (N_41752,N_39944,N_38501);
nor U41753 (N_41753,N_38554,N_39315);
nand U41754 (N_41754,N_39153,N_38551);
xnor U41755 (N_41755,N_39797,N_38202);
and U41756 (N_41756,N_39047,N_37868);
and U41757 (N_41757,N_38242,N_39376);
and U41758 (N_41758,N_39688,N_38247);
nor U41759 (N_41759,N_39295,N_38941);
or U41760 (N_41760,N_38254,N_39822);
or U41761 (N_41761,N_39547,N_38122);
nand U41762 (N_41762,N_39143,N_39299);
xor U41763 (N_41763,N_39043,N_37603);
and U41764 (N_41764,N_37542,N_39321);
and U41765 (N_41765,N_37514,N_38831);
nor U41766 (N_41766,N_38394,N_39067);
nand U41767 (N_41767,N_39138,N_37952);
or U41768 (N_41768,N_39605,N_38879);
xor U41769 (N_41769,N_39170,N_37855);
or U41770 (N_41770,N_39481,N_39760);
or U41771 (N_41771,N_38221,N_39825);
and U41772 (N_41772,N_39129,N_39695);
and U41773 (N_41773,N_39007,N_38308);
and U41774 (N_41774,N_39202,N_37675);
and U41775 (N_41775,N_39829,N_39819);
xnor U41776 (N_41776,N_37716,N_39876);
and U41777 (N_41777,N_38655,N_39421);
xor U41778 (N_41778,N_38664,N_38403);
and U41779 (N_41779,N_39736,N_39181);
xnor U41780 (N_41780,N_39718,N_39675);
nand U41781 (N_41781,N_38890,N_38671);
nand U41782 (N_41782,N_38442,N_39488);
and U41783 (N_41783,N_38378,N_39623);
nor U41784 (N_41784,N_39849,N_39168);
nand U41785 (N_41785,N_39522,N_39147);
xor U41786 (N_41786,N_38577,N_38546);
xnor U41787 (N_41787,N_38490,N_39780);
and U41788 (N_41788,N_38111,N_37807);
or U41789 (N_41789,N_39698,N_39571);
or U41790 (N_41790,N_39345,N_38446);
or U41791 (N_41791,N_38549,N_39928);
or U41792 (N_41792,N_39281,N_39362);
nand U41793 (N_41793,N_38793,N_39655);
nand U41794 (N_41794,N_38458,N_39812);
nand U41795 (N_41795,N_38745,N_38858);
xnor U41796 (N_41796,N_39460,N_37530);
nor U41797 (N_41797,N_38236,N_39977);
nand U41798 (N_41798,N_39377,N_38074);
nand U41799 (N_41799,N_37645,N_38576);
or U41800 (N_41800,N_37999,N_38388);
xor U41801 (N_41801,N_39406,N_39028);
and U41802 (N_41802,N_38666,N_37648);
nand U41803 (N_41803,N_37657,N_38860);
or U41804 (N_41804,N_38268,N_38652);
nor U41805 (N_41805,N_37977,N_37608);
nor U41806 (N_41806,N_39669,N_39465);
nor U41807 (N_41807,N_38262,N_39296);
or U41808 (N_41808,N_38089,N_37534);
xnor U41809 (N_41809,N_38626,N_38230);
or U41810 (N_41810,N_37676,N_38211);
or U41811 (N_41811,N_39462,N_38918);
nor U41812 (N_41812,N_39101,N_37782);
nand U41813 (N_41813,N_37581,N_37797);
nor U41814 (N_41814,N_38050,N_39797);
nand U41815 (N_41815,N_39575,N_39416);
nor U41816 (N_41816,N_39201,N_38529);
and U41817 (N_41817,N_39957,N_37973);
or U41818 (N_41818,N_38358,N_37705);
or U41819 (N_41819,N_38773,N_38430);
nand U41820 (N_41820,N_39382,N_38746);
nand U41821 (N_41821,N_39960,N_37952);
nand U41822 (N_41822,N_38256,N_38806);
xnor U41823 (N_41823,N_37546,N_39162);
nor U41824 (N_41824,N_39900,N_37897);
nor U41825 (N_41825,N_38983,N_37987);
nand U41826 (N_41826,N_38156,N_39941);
and U41827 (N_41827,N_39365,N_38476);
xnor U41828 (N_41828,N_38876,N_39391);
nor U41829 (N_41829,N_38726,N_37817);
nand U41830 (N_41830,N_39775,N_38840);
nand U41831 (N_41831,N_37813,N_38846);
nand U41832 (N_41832,N_38073,N_38230);
xor U41833 (N_41833,N_38152,N_38154);
nand U41834 (N_41834,N_37980,N_38273);
xor U41835 (N_41835,N_38426,N_39597);
nor U41836 (N_41836,N_38732,N_39129);
nand U41837 (N_41837,N_38569,N_39340);
xnor U41838 (N_41838,N_37558,N_39983);
or U41839 (N_41839,N_38401,N_39791);
and U41840 (N_41840,N_38533,N_39943);
nor U41841 (N_41841,N_39927,N_38288);
or U41842 (N_41842,N_39618,N_39734);
or U41843 (N_41843,N_37815,N_38679);
nor U41844 (N_41844,N_37950,N_39038);
and U41845 (N_41845,N_39843,N_38390);
nor U41846 (N_41846,N_38671,N_38475);
and U41847 (N_41847,N_38207,N_38001);
or U41848 (N_41848,N_38280,N_38007);
and U41849 (N_41849,N_37726,N_38560);
and U41850 (N_41850,N_38820,N_38865);
xor U41851 (N_41851,N_39885,N_39175);
or U41852 (N_41852,N_37591,N_38257);
or U41853 (N_41853,N_39612,N_38370);
or U41854 (N_41854,N_38360,N_37857);
xor U41855 (N_41855,N_39748,N_37860);
and U41856 (N_41856,N_39383,N_39565);
nor U41857 (N_41857,N_39354,N_38149);
or U41858 (N_41858,N_38584,N_37714);
and U41859 (N_41859,N_37774,N_38921);
nor U41860 (N_41860,N_39433,N_39047);
xnor U41861 (N_41861,N_37777,N_39759);
or U41862 (N_41862,N_39626,N_38195);
nor U41863 (N_41863,N_39045,N_37826);
nand U41864 (N_41864,N_38412,N_38891);
nor U41865 (N_41865,N_38803,N_37640);
or U41866 (N_41866,N_38680,N_37994);
xnor U41867 (N_41867,N_38273,N_38001);
and U41868 (N_41868,N_39828,N_39700);
or U41869 (N_41869,N_38715,N_38445);
or U41870 (N_41870,N_39091,N_38340);
nand U41871 (N_41871,N_38478,N_39175);
xor U41872 (N_41872,N_38970,N_38791);
xor U41873 (N_41873,N_37694,N_38437);
nor U41874 (N_41874,N_38604,N_39188);
and U41875 (N_41875,N_38253,N_38742);
and U41876 (N_41876,N_39411,N_38156);
xor U41877 (N_41877,N_38408,N_38295);
nand U41878 (N_41878,N_39962,N_37635);
nor U41879 (N_41879,N_38027,N_39484);
nor U41880 (N_41880,N_39753,N_39104);
nor U41881 (N_41881,N_37940,N_38223);
xnor U41882 (N_41882,N_38923,N_37580);
xor U41883 (N_41883,N_39730,N_37583);
nand U41884 (N_41884,N_38228,N_39515);
xnor U41885 (N_41885,N_38953,N_38653);
nand U41886 (N_41886,N_38445,N_39029);
nand U41887 (N_41887,N_38107,N_39576);
nand U41888 (N_41888,N_38008,N_38006);
nor U41889 (N_41889,N_39138,N_39260);
nor U41890 (N_41890,N_38418,N_37501);
and U41891 (N_41891,N_39370,N_39479);
and U41892 (N_41892,N_39634,N_38837);
nor U41893 (N_41893,N_38937,N_39087);
nand U41894 (N_41894,N_39652,N_37826);
and U41895 (N_41895,N_37892,N_38926);
nand U41896 (N_41896,N_37702,N_38672);
and U41897 (N_41897,N_39766,N_38550);
nand U41898 (N_41898,N_39923,N_38996);
nor U41899 (N_41899,N_39752,N_37829);
or U41900 (N_41900,N_39067,N_38798);
and U41901 (N_41901,N_39401,N_39175);
or U41902 (N_41902,N_39122,N_39302);
xor U41903 (N_41903,N_39909,N_37869);
or U41904 (N_41904,N_38144,N_39465);
nor U41905 (N_41905,N_39418,N_38630);
and U41906 (N_41906,N_39390,N_37649);
nand U41907 (N_41907,N_38364,N_38812);
nor U41908 (N_41908,N_39693,N_38079);
xnor U41909 (N_41909,N_38276,N_38483);
xor U41910 (N_41910,N_39460,N_39636);
nand U41911 (N_41911,N_39931,N_39118);
nand U41912 (N_41912,N_38908,N_37684);
or U41913 (N_41913,N_38725,N_38994);
or U41914 (N_41914,N_39745,N_38877);
and U41915 (N_41915,N_37538,N_38830);
or U41916 (N_41916,N_37635,N_38591);
and U41917 (N_41917,N_38238,N_37800);
xor U41918 (N_41918,N_37604,N_39236);
nand U41919 (N_41919,N_37956,N_38898);
and U41920 (N_41920,N_39650,N_38269);
nand U41921 (N_41921,N_38383,N_38289);
nand U41922 (N_41922,N_37597,N_39309);
nor U41923 (N_41923,N_38154,N_38255);
xor U41924 (N_41924,N_38119,N_38913);
nand U41925 (N_41925,N_39726,N_39907);
nand U41926 (N_41926,N_38661,N_39218);
and U41927 (N_41927,N_39909,N_39513);
or U41928 (N_41928,N_38122,N_39214);
nor U41929 (N_41929,N_39414,N_38519);
nand U41930 (N_41930,N_39269,N_38787);
xnor U41931 (N_41931,N_37872,N_39196);
or U41932 (N_41932,N_37762,N_39219);
xor U41933 (N_41933,N_39685,N_39677);
nand U41934 (N_41934,N_39939,N_37521);
and U41935 (N_41935,N_37615,N_38474);
nand U41936 (N_41936,N_38492,N_38942);
or U41937 (N_41937,N_38042,N_39165);
xor U41938 (N_41938,N_37994,N_39509);
or U41939 (N_41939,N_39104,N_39665);
xor U41940 (N_41940,N_39085,N_39245);
or U41941 (N_41941,N_37652,N_39303);
xnor U41942 (N_41942,N_37769,N_38309);
nor U41943 (N_41943,N_37819,N_38517);
nor U41944 (N_41944,N_38836,N_39591);
and U41945 (N_41945,N_38527,N_39329);
xnor U41946 (N_41946,N_38942,N_39341);
and U41947 (N_41947,N_39177,N_37897);
nand U41948 (N_41948,N_38393,N_39464);
nor U41949 (N_41949,N_37634,N_39389);
or U41950 (N_41950,N_39316,N_39912);
or U41951 (N_41951,N_38411,N_39975);
nor U41952 (N_41952,N_38013,N_37780);
nor U41953 (N_41953,N_39673,N_37984);
or U41954 (N_41954,N_39863,N_39626);
or U41955 (N_41955,N_37572,N_37671);
xnor U41956 (N_41956,N_38241,N_39263);
and U41957 (N_41957,N_39250,N_37859);
and U41958 (N_41958,N_39347,N_38642);
xnor U41959 (N_41959,N_39634,N_39348);
nor U41960 (N_41960,N_39306,N_39577);
nor U41961 (N_41961,N_38480,N_38292);
nand U41962 (N_41962,N_38950,N_39940);
or U41963 (N_41963,N_38630,N_37829);
and U41964 (N_41964,N_38828,N_37928);
nor U41965 (N_41965,N_38827,N_39361);
nand U41966 (N_41966,N_38491,N_38288);
or U41967 (N_41967,N_37595,N_39338);
nand U41968 (N_41968,N_38967,N_37856);
nor U41969 (N_41969,N_38313,N_37534);
and U41970 (N_41970,N_39547,N_39648);
and U41971 (N_41971,N_38299,N_37636);
nor U41972 (N_41972,N_38403,N_39413);
nor U41973 (N_41973,N_38701,N_39444);
and U41974 (N_41974,N_38352,N_39499);
xor U41975 (N_41975,N_37859,N_39446);
or U41976 (N_41976,N_39428,N_39407);
and U41977 (N_41977,N_38140,N_37836);
nor U41978 (N_41978,N_39859,N_37591);
nand U41979 (N_41979,N_38881,N_39741);
nor U41980 (N_41980,N_39013,N_39324);
and U41981 (N_41981,N_38670,N_39278);
nand U41982 (N_41982,N_39784,N_38644);
nand U41983 (N_41983,N_39080,N_38281);
nor U41984 (N_41984,N_38216,N_39140);
xor U41985 (N_41985,N_38393,N_37723);
xnor U41986 (N_41986,N_38081,N_38723);
or U41987 (N_41987,N_38161,N_39225);
nand U41988 (N_41988,N_39007,N_38968);
or U41989 (N_41989,N_39624,N_38860);
nand U41990 (N_41990,N_39743,N_38681);
or U41991 (N_41991,N_38144,N_38746);
and U41992 (N_41992,N_37698,N_37931);
nor U41993 (N_41993,N_37933,N_37968);
and U41994 (N_41994,N_37793,N_37824);
xnor U41995 (N_41995,N_39330,N_38597);
and U41996 (N_41996,N_37997,N_39317);
xor U41997 (N_41997,N_38699,N_37786);
or U41998 (N_41998,N_39132,N_39338);
and U41999 (N_41999,N_38700,N_39204);
nor U42000 (N_42000,N_38688,N_39442);
xnor U42001 (N_42001,N_39600,N_38316);
nor U42002 (N_42002,N_38518,N_38867);
and U42003 (N_42003,N_37840,N_38103);
nor U42004 (N_42004,N_38729,N_37854);
nand U42005 (N_42005,N_39705,N_39348);
nand U42006 (N_42006,N_39959,N_38507);
nor U42007 (N_42007,N_39443,N_37846);
and U42008 (N_42008,N_39775,N_39717);
xnor U42009 (N_42009,N_39621,N_38459);
nor U42010 (N_42010,N_38168,N_39989);
and U42011 (N_42011,N_37556,N_39742);
and U42012 (N_42012,N_38688,N_38659);
xnor U42013 (N_42013,N_39940,N_39281);
nand U42014 (N_42014,N_38159,N_38955);
nand U42015 (N_42015,N_39180,N_39665);
and U42016 (N_42016,N_37814,N_38061);
nor U42017 (N_42017,N_39982,N_39275);
nand U42018 (N_42018,N_39314,N_39781);
and U42019 (N_42019,N_39918,N_39764);
and U42020 (N_42020,N_37664,N_38269);
nor U42021 (N_42021,N_38740,N_39455);
xnor U42022 (N_42022,N_38571,N_38401);
or U42023 (N_42023,N_38240,N_38218);
and U42024 (N_42024,N_39729,N_39710);
or U42025 (N_42025,N_38986,N_39891);
and U42026 (N_42026,N_39908,N_39773);
nand U42027 (N_42027,N_39076,N_38065);
or U42028 (N_42028,N_39145,N_37642);
nor U42029 (N_42029,N_39364,N_38330);
xor U42030 (N_42030,N_38175,N_38351);
and U42031 (N_42031,N_38437,N_38271);
nand U42032 (N_42032,N_39190,N_38715);
or U42033 (N_42033,N_39356,N_37706);
and U42034 (N_42034,N_37572,N_39958);
xnor U42035 (N_42035,N_39718,N_38062);
and U42036 (N_42036,N_39204,N_38710);
nand U42037 (N_42037,N_38915,N_38246);
or U42038 (N_42038,N_38343,N_38915);
or U42039 (N_42039,N_38587,N_39427);
nor U42040 (N_42040,N_38806,N_38141);
or U42041 (N_42041,N_37798,N_38691);
and U42042 (N_42042,N_37995,N_39789);
nor U42043 (N_42043,N_37973,N_39532);
xnor U42044 (N_42044,N_39226,N_38734);
and U42045 (N_42045,N_38588,N_38857);
nor U42046 (N_42046,N_39629,N_39685);
nor U42047 (N_42047,N_37840,N_38014);
nand U42048 (N_42048,N_38363,N_39194);
or U42049 (N_42049,N_39201,N_38416);
or U42050 (N_42050,N_39580,N_38146);
and U42051 (N_42051,N_39524,N_37947);
or U42052 (N_42052,N_37983,N_39283);
xnor U42053 (N_42053,N_38851,N_38309);
xnor U42054 (N_42054,N_38086,N_38726);
xnor U42055 (N_42055,N_39354,N_39445);
nand U42056 (N_42056,N_38625,N_38571);
nand U42057 (N_42057,N_39452,N_37801);
nor U42058 (N_42058,N_37823,N_39304);
and U42059 (N_42059,N_38331,N_39822);
xor U42060 (N_42060,N_39551,N_39875);
and U42061 (N_42061,N_37729,N_38840);
nor U42062 (N_42062,N_39156,N_38471);
xnor U42063 (N_42063,N_39812,N_37563);
xnor U42064 (N_42064,N_38340,N_39003);
nand U42065 (N_42065,N_38327,N_39809);
nor U42066 (N_42066,N_38087,N_38895);
nor U42067 (N_42067,N_37620,N_38879);
and U42068 (N_42068,N_39072,N_37566);
and U42069 (N_42069,N_37940,N_39809);
xnor U42070 (N_42070,N_39428,N_38751);
or U42071 (N_42071,N_38973,N_37896);
or U42072 (N_42072,N_39332,N_39717);
nand U42073 (N_42073,N_39740,N_39470);
and U42074 (N_42074,N_37653,N_38297);
and U42075 (N_42075,N_38159,N_38376);
nand U42076 (N_42076,N_38697,N_39463);
nand U42077 (N_42077,N_38718,N_38433);
nor U42078 (N_42078,N_39965,N_38410);
or U42079 (N_42079,N_37836,N_38742);
or U42080 (N_42080,N_37789,N_37957);
or U42081 (N_42081,N_38767,N_38232);
xor U42082 (N_42082,N_39217,N_39317);
nor U42083 (N_42083,N_37999,N_38115);
or U42084 (N_42084,N_38161,N_38428);
nand U42085 (N_42085,N_38989,N_39798);
nand U42086 (N_42086,N_39004,N_38272);
and U42087 (N_42087,N_38744,N_38962);
nor U42088 (N_42088,N_39519,N_38451);
and U42089 (N_42089,N_37822,N_39384);
xnor U42090 (N_42090,N_38645,N_38723);
nor U42091 (N_42091,N_39700,N_38924);
xor U42092 (N_42092,N_39317,N_38090);
and U42093 (N_42093,N_38869,N_38804);
or U42094 (N_42094,N_39626,N_39044);
or U42095 (N_42095,N_38477,N_39726);
xor U42096 (N_42096,N_38605,N_37934);
and U42097 (N_42097,N_38031,N_39174);
nor U42098 (N_42098,N_37664,N_38797);
nand U42099 (N_42099,N_39949,N_38637);
or U42100 (N_42100,N_37673,N_37524);
or U42101 (N_42101,N_37620,N_39839);
nor U42102 (N_42102,N_38090,N_39325);
nand U42103 (N_42103,N_39397,N_38295);
xnor U42104 (N_42104,N_37564,N_39408);
xnor U42105 (N_42105,N_37638,N_38305);
nor U42106 (N_42106,N_37585,N_38400);
xnor U42107 (N_42107,N_39873,N_38031);
nand U42108 (N_42108,N_38246,N_38641);
xnor U42109 (N_42109,N_37515,N_39179);
xnor U42110 (N_42110,N_38116,N_39039);
xor U42111 (N_42111,N_37781,N_39111);
nor U42112 (N_42112,N_38727,N_39412);
or U42113 (N_42113,N_38697,N_39356);
nor U42114 (N_42114,N_39248,N_38172);
nand U42115 (N_42115,N_38770,N_38563);
xnor U42116 (N_42116,N_38653,N_37835);
or U42117 (N_42117,N_38754,N_39683);
and U42118 (N_42118,N_39261,N_37740);
nor U42119 (N_42119,N_38785,N_38997);
nor U42120 (N_42120,N_38374,N_37696);
and U42121 (N_42121,N_37577,N_37633);
nor U42122 (N_42122,N_37537,N_39333);
xor U42123 (N_42123,N_37601,N_38697);
nand U42124 (N_42124,N_39430,N_37690);
xor U42125 (N_42125,N_37963,N_37624);
nand U42126 (N_42126,N_39930,N_39864);
and U42127 (N_42127,N_37835,N_39835);
xor U42128 (N_42128,N_37754,N_38189);
or U42129 (N_42129,N_39469,N_37771);
nor U42130 (N_42130,N_38027,N_37704);
nor U42131 (N_42131,N_39200,N_39684);
or U42132 (N_42132,N_38965,N_38975);
or U42133 (N_42133,N_39182,N_37830);
and U42134 (N_42134,N_39495,N_38054);
or U42135 (N_42135,N_39601,N_39292);
nand U42136 (N_42136,N_38084,N_37628);
or U42137 (N_42137,N_38574,N_37783);
xnor U42138 (N_42138,N_37573,N_39127);
nand U42139 (N_42139,N_38096,N_38855);
and U42140 (N_42140,N_38417,N_38907);
and U42141 (N_42141,N_38423,N_39248);
nand U42142 (N_42142,N_39428,N_39038);
or U42143 (N_42143,N_37553,N_37506);
nor U42144 (N_42144,N_38633,N_37962);
or U42145 (N_42145,N_38277,N_38427);
and U42146 (N_42146,N_38718,N_39123);
and U42147 (N_42147,N_38399,N_38282);
xor U42148 (N_42148,N_39629,N_38158);
nor U42149 (N_42149,N_37971,N_37949);
xnor U42150 (N_42150,N_38563,N_39705);
or U42151 (N_42151,N_38758,N_39535);
nand U42152 (N_42152,N_38754,N_39564);
xor U42153 (N_42153,N_38682,N_39513);
and U42154 (N_42154,N_39958,N_37762);
nand U42155 (N_42155,N_37508,N_38734);
xor U42156 (N_42156,N_39871,N_39850);
and U42157 (N_42157,N_38815,N_39097);
xor U42158 (N_42158,N_38982,N_39412);
nor U42159 (N_42159,N_39873,N_39970);
and U42160 (N_42160,N_38880,N_37932);
and U42161 (N_42161,N_38111,N_39936);
or U42162 (N_42162,N_38253,N_38119);
or U42163 (N_42163,N_38396,N_37865);
nor U42164 (N_42164,N_37808,N_37884);
or U42165 (N_42165,N_37894,N_38821);
and U42166 (N_42166,N_38876,N_39188);
or U42167 (N_42167,N_39609,N_39454);
nor U42168 (N_42168,N_38764,N_37675);
xor U42169 (N_42169,N_37819,N_39880);
and U42170 (N_42170,N_38306,N_39009);
nor U42171 (N_42171,N_37575,N_38972);
nand U42172 (N_42172,N_39704,N_37936);
or U42173 (N_42173,N_38226,N_39280);
and U42174 (N_42174,N_38487,N_37840);
or U42175 (N_42175,N_38009,N_39355);
nor U42176 (N_42176,N_39904,N_37737);
xor U42177 (N_42177,N_39788,N_37931);
and U42178 (N_42178,N_39602,N_39554);
nor U42179 (N_42179,N_38460,N_37578);
or U42180 (N_42180,N_38923,N_38452);
xnor U42181 (N_42181,N_38551,N_38652);
or U42182 (N_42182,N_39472,N_39095);
nor U42183 (N_42183,N_38353,N_38691);
and U42184 (N_42184,N_38135,N_38068);
and U42185 (N_42185,N_38015,N_39939);
nand U42186 (N_42186,N_39179,N_38440);
and U42187 (N_42187,N_39095,N_39671);
nand U42188 (N_42188,N_37507,N_38405);
xor U42189 (N_42189,N_39799,N_38080);
xnor U42190 (N_42190,N_39535,N_38406);
or U42191 (N_42191,N_37644,N_37763);
nor U42192 (N_42192,N_39455,N_38057);
xnor U42193 (N_42193,N_39735,N_39948);
nor U42194 (N_42194,N_39409,N_37657);
nand U42195 (N_42195,N_39421,N_37716);
or U42196 (N_42196,N_38512,N_39817);
xnor U42197 (N_42197,N_38666,N_37880);
and U42198 (N_42198,N_37688,N_37675);
nor U42199 (N_42199,N_39583,N_38473);
nand U42200 (N_42200,N_37617,N_37763);
and U42201 (N_42201,N_39391,N_38888);
or U42202 (N_42202,N_38049,N_38967);
nand U42203 (N_42203,N_37807,N_39556);
nand U42204 (N_42204,N_38785,N_39764);
or U42205 (N_42205,N_37802,N_38403);
and U42206 (N_42206,N_39781,N_39684);
and U42207 (N_42207,N_37647,N_38605);
nor U42208 (N_42208,N_37573,N_39682);
and U42209 (N_42209,N_39688,N_39552);
and U42210 (N_42210,N_37685,N_38862);
xor U42211 (N_42211,N_38828,N_39297);
and U42212 (N_42212,N_38720,N_38928);
xor U42213 (N_42213,N_39457,N_38338);
or U42214 (N_42214,N_37727,N_39097);
nand U42215 (N_42215,N_37677,N_39361);
nand U42216 (N_42216,N_38664,N_38839);
or U42217 (N_42217,N_38456,N_39417);
and U42218 (N_42218,N_39159,N_38248);
xor U42219 (N_42219,N_38201,N_38501);
xor U42220 (N_42220,N_39993,N_39645);
nor U42221 (N_42221,N_39147,N_37654);
xor U42222 (N_42222,N_39831,N_38673);
and U42223 (N_42223,N_38719,N_38360);
nor U42224 (N_42224,N_38485,N_37938);
or U42225 (N_42225,N_37940,N_38686);
or U42226 (N_42226,N_39306,N_39359);
nor U42227 (N_42227,N_39293,N_37923);
and U42228 (N_42228,N_38745,N_38391);
nor U42229 (N_42229,N_38828,N_38670);
nor U42230 (N_42230,N_39128,N_38500);
xnor U42231 (N_42231,N_39638,N_38395);
xor U42232 (N_42232,N_39183,N_38990);
nand U42233 (N_42233,N_39653,N_37605);
or U42234 (N_42234,N_37507,N_37570);
or U42235 (N_42235,N_39846,N_38815);
nor U42236 (N_42236,N_38210,N_38610);
nor U42237 (N_42237,N_38896,N_38232);
or U42238 (N_42238,N_39164,N_39662);
xnor U42239 (N_42239,N_37613,N_38658);
and U42240 (N_42240,N_37546,N_39470);
and U42241 (N_42241,N_38406,N_39108);
or U42242 (N_42242,N_39594,N_38552);
xnor U42243 (N_42243,N_38843,N_38111);
or U42244 (N_42244,N_38697,N_38613);
and U42245 (N_42245,N_37770,N_38495);
nor U42246 (N_42246,N_39255,N_39423);
nor U42247 (N_42247,N_38346,N_39209);
or U42248 (N_42248,N_38315,N_39673);
nand U42249 (N_42249,N_37937,N_37618);
nand U42250 (N_42250,N_39430,N_39792);
nand U42251 (N_42251,N_37825,N_38839);
nor U42252 (N_42252,N_39037,N_37675);
or U42253 (N_42253,N_39289,N_37606);
or U42254 (N_42254,N_38061,N_38656);
and U42255 (N_42255,N_39505,N_37631);
or U42256 (N_42256,N_39208,N_38010);
nand U42257 (N_42257,N_39883,N_38022);
nor U42258 (N_42258,N_38518,N_39819);
nor U42259 (N_42259,N_38677,N_37818);
nor U42260 (N_42260,N_39635,N_38996);
nor U42261 (N_42261,N_38863,N_38458);
xor U42262 (N_42262,N_38879,N_39599);
xor U42263 (N_42263,N_38085,N_39508);
or U42264 (N_42264,N_37682,N_38968);
and U42265 (N_42265,N_38867,N_39532);
and U42266 (N_42266,N_39296,N_38931);
nand U42267 (N_42267,N_37544,N_38796);
nand U42268 (N_42268,N_38511,N_38921);
nor U42269 (N_42269,N_37672,N_37845);
or U42270 (N_42270,N_39359,N_39789);
xnor U42271 (N_42271,N_38119,N_38967);
nand U42272 (N_42272,N_37830,N_38372);
nor U42273 (N_42273,N_39199,N_39692);
or U42274 (N_42274,N_39744,N_39039);
xor U42275 (N_42275,N_38446,N_39030);
or U42276 (N_42276,N_37580,N_39248);
nor U42277 (N_42277,N_37584,N_37841);
nand U42278 (N_42278,N_38975,N_38664);
and U42279 (N_42279,N_37668,N_38861);
nor U42280 (N_42280,N_37728,N_39445);
or U42281 (N_42281,N_37995,N_38459);
and U42282 (N_42282,N_39316,N_39575);
nand U42283 (N_42283,N_38060,N_39916);
nor U42284 (N_42284,N_38081,N_38942);
and U42285 (N_42285,N_39707,N_39142);
xnor U42286 (N_42286,N_38543,N_37876);
nor U42287 (N_42287,N_37961,N_38844);
and U42288 (N_42288,N_39773,N_39878);
or U42289 (N_42289,N_39492,N_39656);
nand U42290 (N_42290,N_38423,N_37704);
nand U42291 (N_42291,N_39551,N_39632);
xor U42292 (N_42292,N_38544,N_39319);
or U42293 (N_42293,N_38178,N_39806);
nand U42294 (N_42294,N_38258,N_37774);
and U42295 (N_42295,N_38141,N_38812);
or U42296 (N_42296,N_39430,N_37510);
nor U42297 (N_42297,N_37824,N_37529);
and U42298 (N_42298,N_37789,N_39335);
xnor U42299 (N_42299,N_39210,N_38253);
nand U42300 (N_42300,N_39616,N_38946);
xnor U42301 (N_42301,N_38635,N_38126);
or U42302 (N_42302,N_38328,N_39364);
or U42303 (N_42303,N_38442,N_38091);
nor U42304 (N_42304,N_39183,N_39762);
or U42305 (N_42305,N_39933,N_37653);
and U42306 (N_42306,N_38198,N_38051);
nor U42307 (N_42307,N_37933,N_39251);
xnor U42308 (N_42308,N_38406,N_37945);
xor U42309 (N_42309,N_39348,N_39000);
and U42310 (N_42310,N_38129,N_39335);
nand U42311 (N_42311,N_37537,N_39606);
xnor U42312 (N_42312,N_37892,N_38364);
xor U42313 (N_42313,N_39054,N_38038);
nand U42314 (N_42314,N_37758,N_38962);
xnor U42315 (N_42315,N_37938,N_38859);
or U42316 (N_42316,N_38648,N_38704);
or U42317 (N_42317,N_38954,N_39134);
or U42318 (N_42318,N_38502,N_39404);
or U42319 (N_42319,N_39446,N_38665);
nor U42320 (N_42320,N_39362,N_38246);
nor U42321 (N_42321,N_38708,N_39088);
or U42322 (N_42322,N_39765,N_38549);
nor U42323 (N_42323,N_38243,N_39260);
and U42324 (N_42324,N_39268,N_37998);
or U42325 (N_42325,N_38555,N_38553);
nand U42326 (N_42326,N_39144,N_38326);
or U42327 (N_42327,N_39216,N_38872);
and U42328 (N_42328,N_39186,N_39119);
or U42329 (N_42329,N_38914,N_39162);
nand U42330 (N_42330,N_37612,N_39458);
xnor U42331 (N_42331,N_38552,N_38314);
and U42332 (N_42332,N_38144,N_38817);
nand U42333 (N_42333,N_39960,N_38790);
nor U42334 (N_42334,N_38441,N_39121);
or U42335 (N_42335,N_38208,N_39864);
nor U42336 (N_42336,N_38328,N_39918);
xnor U42337 (N_42337,N_38523,N_38367);
nand U42338 (N_42338,N_39255,N_39767);
xor U42339 (N_42339,N_39624,N_38158);
xor U42340 (N_42340,N_38278,N_38858);
xor U42341 (N_42341,N_38645,N_38887);
nor U42342 (N_42342,N_37632,N_37541);
or U42343 (N_42343,N_38716,N_39584);
xnor U42344 (N_42344,N_39637,N_39142);
xor U42345 (N_42345,N_39707,N_39373);
xnor U42346 (N_42346,N_39152,N_38527);
nor U42347 (N_42347,N_37970,N_39444);
xnor U42348 (N_42348,N_37511,N_38633);
or U42349 (N_42349,N_39379,N_37541);
or U42350 (N_42350,N_39690,N_39085);
nor U42351 (N_42351,N_39498,N_39532);
nor U42352 (N_42352,N_39595,N_38408);
xnor U42353 (N_42353,N_38804,N_38019);
xor U42354 (N_42354,N_39803,N_38897);
nand U42355 (N_42355,N_39770,N_38838);
nor U42356 (N_42356,N_39727,N_38959);
or U42357 (N_42357,N_38380,N_38114);
nor U42358 (N_42358,N_39084,N_37823);
or U42359 (N_42359,N_39520,N_39515);
and U42360 (N_42360,N_39764,N_38167);
and U42361 (N_42361,N_38368,N_39754);
nor U42362 (N_42362,N_37809,N_37960);
nor U42363 (N_42363,N_39894,N_39514);
xor U42364 (N_42364,N_37886,N_37879);
and U42365 (N_42365,N_38603,N_39672);
and U42366 (N_42366,N_38965,N_37504);
or U42367 (N_42367,N_37722,N_39705);
and U42368 (N_42368,N_38237,N_38270);
nor U42369 (N_42369,N_38046,N_39781);
and U42370 (N_42370,N_39239,N_38647);
xnor U42371 (N_42371,N_37614,N_39378);
xnor U42372 (N_42372,N_39327,N_38449);
nor U42373 (N_42373,N_38394,N_38040);
xnor U42374 (N_42374,N_39825,N_39272);
nand U42375 (N_42375,N_39328,N_39769);
nor U42376 (N_42376,N_39242,N_39787);
or U42377 (N_42377,N_39549,N_38957);
xor U42378 (N_42378,N_39107,N_37988);
nor U42379 (N_42379,N_39939,N_38605);
xnor U42380 (N_42380,N_37664,N_37840);
and U42381 (N_42381,N_38939,N_38626);
or U42382 (N_42382,N_39750,N_38375);
and U42383 (N_42383,N_39497,N_37951);
and U42384 (N_42384,N_38277,N_38776);
nand U42385 (N_42385,N_38771,N_39710);
nand U42386 (N_42386,N_37666,N_38742);
and U42387 (N_42387,N_39963,N_37786);
nand U42388 (N_42388,N_37620,N_39909);
xor U42389 (N_42389,N_38437,N_38111);
and U42390 (N_42390,N_37861,N_38026);
and U42391 (N_42391,N_37984,N_39256);
xor U42392 (N_42392,N_38696,N_38219);
or U42393 (N_42393,N_39881,N_37909);
or U42394 (N_42394,N_39093,N_38823);
or U42395 (N_42395,N_38466,N_37887);
xnor U42396 (N_42396,N_39745,N_39810);
or U42397 (N_42397,N_39385,N_39774);
or U42398 (N_42398,N_38215,N_39165);
nand U42399 (N_42399,N_39480,N_39806);
nor U42400 (N_42400,N_39448,N_39638);
or U42401 (N_42401,N_38041,N_37796);
nand U42402 (N_42402,N_37735,N_38520);
or U42403 (N_42403,N_38195,N_38790);
xor U42404 (N_42404,N_39143,N_39869);
xor U42405 (N_42405,N_37792,N_38574);
or U42406 (N_42406,N_37673,N_37543);
nor U42407 (N_42407,N_38813,N_39897);
nand U42408 (N_42408,N_39417,N_39309);
xor U42409 (N_42409,N_38426,N_37541);
xnor U42410 (N_42410,N_37806,N_37831);
xnor U42411 (N_42411,N_39897,N_38325);
nand U42412 (N_42412,N_37833,N_39849);
and U42413 (N_42413,N_38454,N_39372);
xor U42414 (N_42414,N_39723,N_39449);
or U42415 (N_42415,N_37638,N_38321);
or U42416 (N_42416,N_37735,N_39315);
nand U42417 (N_42417,N_37926,N_39637);
and U42418 (N_42418,N_39775,N_37916);
nand U42419 (N_42419,N_39756,N_37633);
nand U42420 (N_42420,N_37924,N_39998);
and U42421 (N_42421,N_38598,N_38696);
or U42422 (N_42422,N_38182,N_38016);
or U42423 (N_42423,N_38629,N_38163);
and U42424 (N_42424,N_39656,N_39828);
nor U42425 (N_42425,N_37847,N_38095);
xor U42426 (N_42426,N_38010,N_38833);
or U42427 (N_42427,N_38558,N_39724);
nor U42428 (N_42428,N_39379,N_39078);
or U42429 (N_42429,N_38990,N_38128);
nor U42430 (N_42430,N_37700,N_39794);
and U42431 (N_42431,N_37938,N_38468);
nor U42432 (N_42432,N_37818,N_38399);
nor U42433 (N_42433,N_39163,N_38715);
nor U42434 (N_42434,N_38463,N_39820);
or U42435 (N_42435,N_38604,N_39193);
nor U42436 (N_42436,N_38759,N_38271);
nor U42437 (N_42437,N_39867,N_39674);
and U42438 (N_42438,N_39902,N_39618);
or U42439 (N_42439,N_39512,N_39765);
nand U42440 (N_42440,N_38735,N_38327);
or U42441 (N_42441,N_38628,N_39130);
nor U42442 (N_42442,N_39473,N_37831);
xnor U42443 (N_42443,N_38510,N_39979);
or U42444 (N_42444,N_37626,N_38654);
nand U42445 (N_42445,N_38747,N_39381);
or U42446 (N_42446,N_39668,N_39545);
xnor U42447 (N_42447,N_37514,N_39998);
and U42448 (N_42448,N_39839,N_38460);
nand U42449 (N_42449,N_38629,N_39733);
or U42450 (N_42450,N_38359,N_39190);
xor U42451 (N_42451,N_38720,N_38187);
nor U42452 (N_42452,N_38040,N_38321);
nand U42453 (N_42453,N_37742,N_38630);
or U42454 (N_42454,N_38949,N_39165);
nand U42455 (N_42455,N_37574,N_37772);
nand U42456 (N_42456,N_39053,N_39108);
nand U42457 (N_42457,N_39059,N_38645);
or U42458 (N_42458,N_39378,N_39628);
or U42459 (N_42459,N_37754,N_38092);
and U42460 (N_42460,N_37804,N_37668);
or U42461 (N_42461,N_38669,N_38794);
or U42462 (N_42462,N_37989,N_37910);
or U42463 (N_42463,N_39545,N_38505);
and U42464 (N_42464,N_39549,N_39128);
xnor U42465 (N_42465,N_38094,N_38701);
nor U42466 (N_42466,N_39974,N_37582);
xnor U42467 (N_42467,N_39003,N_39389);
xnor U42468 (N_42468,N_39379,N_37589);
xor U42469 (N_42469,N_39311,N_39173);
and U42470 (N_42470,N_37830,N_39023);
nor U42471 (N_42471,N_38124,N_37851);
and U42472 (N_42472,N_39879,N_37711);
or U42473 (N_42473,N_39615,N_39528);
and U42474 (N_42474,N_39528,N_37561);
xor U42475 (N_42475,N_39833,N_39823);
nor U42476 (N_42476,N_38667,N_39018);
and U42477 (N_42477,N_39086,N_39503);
nor U42478 (N_42478,N_38132,N_38040);
or U42479 (N_42479,N_38856,N_38335);
nand U42480 (N_42480,N_39602,N_38288);
xor U42481 (N_42481,N_39495,N_37826);
nand U42482 (N_42482,N_39072,N_38144);
and U42483 (N_42483,N_39059,N_39735);
nor U42484 (N_42484,N_39525,N_38495);
and U42485 (N_42485,N_39218,N_37775);
and U42486 (N_42486,N_38824,N_39002);
nand U42487 (N_42487,N_39508,N_37659);
and U42488 (N_42488,N_37794,N_38444);
nand U42489 (N_42489,N_38200,N_38986);
nor U42490 (N_42490,N_38381,N_38992);
or U42491 (N_42491,N_39545,N_39711);
and U42492 (N_42492,N_39455,N_39717);
and U42493 (N_42493,N_38385,N_38735);
nand U42494 (N_42494,N_39087,N_39685);
nand U42495 (N_42495,N_37986,N_38474);
xor U42496 (N_42496,N_39465,N_39776);
or U42497 (N_42497,N_39662,N_38502);
and U42498 (N_42498,N_39160,N_39020);
nor U42499 (N_42499,N_39131,N_38970);
nor U42500 (N_42500,N_40354,N_41279);
nand U42501 (N_42501,N_41821,N_40782);
and U42502 (N_42502,N_42161,N_42244);
and U42503 (N_42503,N_41131,N_40463);
xnor U42504 (N_42504,N_41252,N_41349);
or U42505 (N_42505,N_42223,N_41341);
xor U42506 (N_42506,N_42346,N_40734);
xor U42507 (N_42507,N_40449,N_41222);
or U42508 (N_42508,N_40604,N_40661);
xnor U42509 (N_42509,N_42114,N_41264);
nor U42510 (N_42510,N_41840,N_40718);
or U42511 (N_42511,N_41515,N_41853);
xnor U42512 (N_42512,N_41561,N_41670);
xnor U42513 (N_42513,N_41908,N_42145);
and U42514 (N_42514,N_40248,N_41461);
nor U42515 (N_42515,N_40885,N_40528);
nor U42516 (N_42516,N_42224,N_41790);
or U42517 (N_42517,N_41391,N_41717);
xnor U42518 (N_42518,N_40769,N_40890);
or U42519 (N_42519,N_42280,N_42379);
and U42520 (N_42520,N_41620,N_40429);
or U42521 (N_42521,N_40222,N_41224);
xnor U42522 (N_42522,N_41204,N_42478);
xnor U42523 (N_42523,N_40450,N_40113);
nor U42524 (N_42524,N_41291,N_40492);
or U42525 (N_42525,N_40610,N_40818);
nor U42526 (N_42526,N_41812,N_42019);
xnor U42527 (N_42527,N_40922,N_41275);
nor U42528 (N_42528,N_40807,N_40733);
nand U42529 (N_42529,N_41991,N_42493);
or U42530 (N_42530,N_40617,N_42476);
nand U42531 (N_42531,N_40259,N_40746);
or U42532 (N_42532,N_41307,N_40561);
nor U42533 (N_42533,N_40434,N_40020);
nor U42534 (N_42534,N_40220,N_41859);
or U42535 (N_42535,N_42182,N_42207);
nand U42536 (N_42536,N_40192,N_40419);
or U42537 (N_42537,N_41591,N_40983);
and U42538 (N_42538,N_41419,N_40501);
xor U42539 (N_42539,N_42459,N_40652);
or U42540 (N_42540,N_40148,N_40452);
nand U42541 (N_42541,N_40611,N_40189);
and U42542 (N_42542,N_41069,N_41094);
nor U42543 (N_42543,N_41874,N_41711);
xnor U42544 (N_42544,N_40815,N_41796);
or U42545 (N_42545,N_40755,N_42196);
nor U42546 (N_42546,N_42366,N_41541);
and U42547 (N_42547,N_42219,N_40977);
nor U42548 (N_42548,N_41406,N_42110);
xor U42549 (N_42549,N_41677,N_40163);
or U42550 (N_42550,N_42386,N_40962);
xor U42551 (N_42551,N_41707,N_42230);
xor U42552 (N_42552,N_42056,N_41046);
or U42553 (N_42553,N_40062,N_42358);
or U42554 (N_42554,N_41987,N_41443);
or U42555 (N_42555,N_40286,N_42337);
and U42556 (N_42556,N_41892,N_40888);
or U42557 (N_42557,N_41301,N_40064);
xor U42558 (N_42558,N_41640,N_41522);
or U42559 (N_42559,N_42263,N_41937);
or U42560 (N_42560,N_41453,N_40093);
nand U42561 (N_42561,N_42170,N_41034);
or U42562 (N_42562,N_41811,N_40010);
nor U42563 (N_42563,N_40297,N_41241);
nand U42564 (N_42564,N_42037,N_41184);
nand U42565 (N_42565,N_40421,N_40787);
or U42566 (N_42566,N_41495,N_41862);
xnor U42567 (N_42567,N_41190,N_41535);
nor U42568 (N_42568,N_42333,N_41834);
and U42569 (N_42569,N_40088,N_40477);
nand U42570 (N_42570,N_42365,N_41078);
xor U42571 (N_42571,N_40892,N_40041);
or U42572 (N_42572,N_41837,N_41858);
xnor U42573 (N_42573,N_41102,N_42240);
or U42574 (N_42574,N_40210,N_40442);
and U42575 (N_42575,N_40871,N_41693);
nor U42576 (N_42576,N_40155,N_40811);
xnor U42577 (N_42577,N_42347,N_41753);
and U42578 (N_42578,N_41676,N_40848);
and U42579 (N_42579,N_42010,N_41829);
xnor U42580 (N_42580,N_41295,N_40038);
nor U42581 (N_42581,N_41182,N_41942);
nor U42582 (N_42582,N_40496,N_41254);
and U42583 (N_42583,N_42312,N_40271);
or U42584 (N_42584,N_41333,N_42177);
or U42585 (N_42585,N_40771,N_41319);
and U42586 (N_42586,N_42495,N_41985);
or U42587 (N_42587,N_40785,N_40412);
nor U42588 (N_42588,N_40567,N_40318);
xor U42589 (N_42589,N_41146,N_40999);
nand U42590 (N_42590,N_40373,N_40986);
or U42591 (N_42591,N_40876,N_40312);
and U42592 (N_42592,N_41695,N_40550);
nor U42593 (N_42593,N_41183,N_40670);
or U42594 (N_42594,N_40711,N_40676);
nand U42595 (N_42595,N_40569,N_41962);
and U42596 (N_42596,N_41323,N_42143);
nor U42597 (N_42597,N_40397,N_42176);
nand U42598 (N_42598,N_40277,N_40873);
or U42599 (N_42599,N_41526,N_41806);
or U42600 (N_42600,N_40000,N_41557);
nor U42601 (N_42601,N_41532,N_42301);
and U42602 (N_42602,N_42189,N_40531);
nand U42603 (N_42603,N_42107,N_40680);
and U42604 (N_42604,N_41718,N_40039);
or U42605 (N_42605,N_41313,N_40383);
or U42606 (N_42606,N_41053,N_40984);
xor U42607 (N_42607,N_41366,N_41473);
nor U42608 (N_42608,N_40651,N_41000);
nand U42609 (N_42609,N_42348,N_41126);
nand U42610 (N_42610,N_41478,N_41995);
xnor U42611 (N_42611,N_40003,N_41001);
and U42612 (N_42612,N_42443,N_40294);
nor U42613 (N_42613,N_40539,N_40518);
xnor U42614 (N_42614,N_40936,N_40262);
and U42615 (N_42615,N_41090,N_40058);
and U42616 (N_42616,N_40773,N_40594);
xnor U42617 (N_42617,N_41467,N_42133);
and U42618 (N_42618,N_40001,N_40705);
xnor U42619 (N_42619,N_41855,N_40592);
nor U42620 (N_42620,N_42242,N_41506);
and U42621 (N_42621,N_41548,N_40346);
nor U42622 (N_42622,N_41353,N_41994);
or U42623 (N_42623,N_41003,N_40527);
nand U42624 (N_42624,N_42142,N_42105);
xor U42625 (N_42625,N_40370,N_40844);
xnor U42626 (N_42626,N_40647,N_41423);
xnor U42627 (N_42627,N_41340,N_41559);
or U42628 (N_42628,N_41822,N_40883);
and U42629 (N_42629,N_42368,N_41037);
nand U42630 (N_42630,N_40216,N_40517);
nor U42631 (N_42631,N_42456,N_40387);
or U42632 (N_42632,N_41881,N_40959);
nand U42633 (N_42633,N_41563,N_40468);
nor U42634 (N_42634,N_41481,N_42445);
and U42635 (N_42635,N_40034,N_40909);
nor U42636 (N_42636,N_40250,N_40066);
and U42637 (N_42637,N_41352,N_40196);
xor U42638 (N_42638,N_40448,N_40972);
xnor U42639 (N_42639,N_41121,N_42123);
and U42640 (N_42640,N_40514,N_41688);
xor U42641 (N_42641,N_41975,N_40016);
nand U42642 (N_42642,N_41984,N_41097);
and U42643 (N_42643,N_41487,N_40748);
or U42644 (N_42644,N_41629,N_41668);
xor U42645 (N_42645,N_40221,N_40076);
and U42646 (N_42646,N_41757,N_40245);
and U42647 (N_42647,N_41760,N_40745);
or U42648 (N_42648,N_40882,N_42474);
nand U42649 (N_42649,N_41059,N_40825);
nand U42650 (N_42650,N_40503,N_41068);
xnor U42651 (N_42651,N_41882,N_41215);
nand U42652 (N_42652,N_41095,N_42109);
xnor U42653 (N_42653,N_40126,N_40166);
or U42654 (N_42654,N_41597,N_42414);
nor U42655 (N_42655,N_40478,N_42178);
nand U42656 (N_42656,N_41347,N_40147);
xnor U42657 (N_42657,N_40994,N_42210);
nor U42658 (N_42658,N_41084,N_40684);
xor U42659 (N_42659,N_40123,N_40515);
nand U42660 (N_42660,N_40151,N_40841);
nor U42661 (N_42661,N_42141,N_40823);
or U42662 (N_42662,N_40935,N_40176);
nand U42663 (N_42663,N_42048,N_40507);
nand U42664 (N_42664,N_42441,N_42147);
nor U42665 (N_42665,N_42018,N_41221);
or U42666 (N_42666,N_41415,N_42423);
and U42667 (N_42667,N_40403,N_41007);
xor U42668 (N_42668,N_40961,N_41550);
or U42669 (N_42669,N_40854,N_42124);
or U42670 (N_42670,N_40654,N_41468);
nand U42671 (N_42671,N_40369,N_41031);
and U42672 (N_42672,N_40239,N_41165);
xor U42673 (N_42673,N_42231,N_41459);
xor U42674 (N_42674,N_41311,N_40764);
xor U42675 (N_42675,N_40568,N_40025);
or U42676 (N_42676,N_42465,N_40473);
nand U42677 (N_42677,N_41838,N_41267);
xor U42678 (N_42678,N_41449,N_42483);
or U42679 (N_42679,N_41079,N_41883);
nand U42680 (N_42680,N_41618,N_41742);
nand U42681 (N_42681,N_40122,N_40253);
xnor U42682 (N_42682,N_41334,N_40788);
nor U42683 (N_42683,N_42289,N_41286);
nor U42684 (N_42684,N_41450,N_40943);
nor U42685 (N_42685,N_40279,N_41705);
xnor U42686 (N_42686,N_41509,N_40632);
xor U42687 (N_42687,N_41242,N_41260);
or U42688 (N_42688,N_40278,N_40887);
xnor U42689 (N_42689,N_41163,N_42259);
and U42690 (N_42690,N_41475,N_41484);
and U42691 (N_42691,N_41910,N_41738);
and U42692 (N_42692,N_40668,N_40090);
xor U42693 (N_42693,N_41852,N_40141);
nand U42694 (N_42694,N_40585,N_40616);
or U42695 (N_42695,N_41781,N_40565);
or U42696 (N_42696,N_41581,N_40461);
nand U42697 (N_42697,N_41219,N_42357);
and U42698 (N_42698,N_42429,N_41022);
nor U42699 (N_42699,N_41844,N_40819);
nand U42700 (N_42700,N_40916,N_42430);
nand U42701 (N_42701,N_41486,N_41582);
nor U42702 (N_42702,N_40710,N_40698);
or U42703 (N_42703,N_40015,N_41565);
nand U42704 (N_42704,N_40886,N_41685);
or U42705 (N_42705,N_42269,N_41359);
nor U42706 (N_42706,N_41702,N_40260);
nor U42707 (N_42707,N_41015,N_40645);
and U42708 (N_42708,N_41240,N_40071);
or U42709 (N_42709,N_40197,N_42282);
xnor U42710 (N_42710,N_40095,N_41152);
xnor U42711 (N_42711,N_40047,N_40227);
or U42712 (N_42712,N_41873,N_41642);
nor U42713 (N_42713,N_42261,N_41657);
and U42714 (N_42714,N_40541,N_41813);
nor U42715 (N_42715,N_40355,N_40300);
and U42716 (N_42716,N_42045,N_42011);
and U42717 (N_42717,N_42071,N_42250);
nand U42718 (N_42718,N_40418,N_40415);
nor U42719 (N_42719,N_40454,N_42129);
or U42720 (N_42720,N_40979,N_40551);
and U42721 (N_42721,N_41592,N_40140);
nor U42722 (N_42722,N_40942,N_40441);
nor U42723 (N_42723,N_41516,N_40945);
xor U42724 (N_42724,N_41961,N_40362);
nand U42725 (N_42725,N_42460,N_40709);
or U42726 (N_42726,N_41201,N_41300);
nor U42727 (N_42727,N_42079,N_40004);
nor U42728 (N_42728,N_41040,N_42006);
nand U42729 (N_42729,N_40627,N_41886);
nor U42730 (N_42730,N_41730,N_40809);
xnor U42731 (N_42731,N_41610,N_40414);
nor U42732 (N_42732,N_42043,N_40570);
nor U42733 (N_42733,N_42398,N_40435);
or U42734 (N_42734,N_41703,N_41628);
nand U42735 (N_42735,N_40763,N_42464);
nand U42736 (N_42736,N_41198,N_40919);
nand U42737 (N_42737,N_41277,N_41715);
nand U42738 (N_42738,N_40267,N_41137);
xnor U42739 (N_42739,N_40455,N_41117);
xor U42740 (N_42740,N_41181,N_41505);
or U42741 (N_42741,N_40630,N_42197);
or U42742 (N_42742,N_41303,N_42050);
or U42743 (N_42743,N_40615,N_40814);
nand U42744 (N_42744,N_40862,N_40870);
nor U42745 (N_42745,N_40420,N_40662);
or U42746 (N_42746,N_40152,N_40111);
nand U42747 (N_42747,N_40756,N_41361);
nor U42748 (N_42748,N_41614,N_41250);
nand U42749 (N_42749,N_41116,N_40506);
nor U42750 (N_42750,N_42425,N_41316);
xor U42751 (N_42751,N_41868,N_42064);
and U42752 (N_42752,N_40603,N_42377);
nor U42753 (N_42753,N_40821,N_40067);
nor U42754 (N_42754,N_42059,N_40717);
or U42755 (N_42755,N_41997,N_42229);
nand U42756 (N_42756,N_40786,N_40775);
xnor U42757 (N_42757,N_42438,N_40036);
and U42758 (N_42758,N_42281,N_42283);
or U42759 (N_42759,N_40522,N_41590);
nor U42760 (N_42760,N_41722,N_41931);
and U42761 (N_42761,N_41047,N_40485);
or U42762 (N_42762,N_40860,N_41584);
and U42763 (N_42763,N_40700,N_41470);
or U42764 (N_42764,N_42299,N_41210);
and U42765 (N_42765,N_40874,N_42345);
and U42766 (N_42766,N_42111,N_40044);
nand U42767 (N_42767,N_41424,N_41740);
or U42768 (N_42768,N_42391,N_41355);
xnor U42769 (N_42769,N_40537,N_42354);
xor U42770 (N_42770,N_41570,N_41809);
or U42771 (N_42771,N_41220,N_41429);
nand U42772 (N_42772,N_41399,N_40149);
or U42773 (N_42773,N_41887,N_40526);
nand U42774 (N_42774,N_40164,N_40377);
nand U42775 (N_42775,N_41772,N_41365);
and U42776 (N_42776,N_41802,N_41294);
or U42777 (N_42777,N_42463,N_40317);
nand U42778 (N_42778,N_40857,N_41919);
or U42779 (N_42779,N_41482,N_42163);
or U42780 (N_42780,N_41589,N_41168);
nor U42781 (N_42781,N_40589,N_41662);
nand U42782 (N_42782,N_42093,N_40523);
nor U42783 (N_42783,N_40835,N_40658);
nand U42784 (N_42784,N_40491,N_40704);
or U42785 (N_42785,N_41872,N_42288);
nand U42786 (N_42786,N_41914,N_41587);
and U42787 (N_42787,N_40063,N_40946);
nor U42788 (N_42788,N_40779,N_41746);
nor U42789 (N_42789,N_40446,N_41777);
nor U42790 (N_42790,N_41368,N_41783);
nand U42791 (N_42791,N_41151,N_41343);
nor U42792 (N_42792,N_40366,N_40750);
nor U42793 (N_42793,N_42239,N_42336);
and U42794 (N_42794,N_40112,N_42328);
xor U42795 (N_42795,N_41636,N_41907);
and U42796 (N_42796,N_40017,N_40214);
nor U42797 (N_42797,N_40653,N_40213);
or U42798 (N_42798,N_41944,N_42304);
xnor U42799 (N_42799,N_40749,N_42297);
and U42800 (N_42800,N_42199,N_41965);
nand U42801 (N_42801,N_40107,N_40822);
nand U42802 (N_42802,N_42015,N_41042);
or U42803 (N_42803,N_41077,N_42317);
xnor U42804 (N_42804,N_40901,N_41776);
and U42805 (N_42805,N_42054,N_40060);
or U42806 (N_42806,N_41903,N_40263);
and U42807 (N_42807,N_42405,N_40465);
or U42808 (N_42808,N_40826,N_40538);
nor U42809 (N_42809,N_41594,N_41651);
or U42810 (N_42810,N_40856,N_42021);
or U42811 (N_42811,N_40070,N_41237);
nor U42812 (N_42812,N_42380,N_42130);
or U42813 (N_42813,N_41161,N_40343);
xnor U42814 (N_42814,N_40389,N_41915);
or U42815 (N_42815,N_41744,N_40520);
nand U42816 (N_42816,N_40323,N_41070);
nand U42817 (N_42817,N_41752,N_40046);
nand U42818 (N_42818,N_41876,N_41422);
and U42819 (N_42819,N_42321,N_41315);
xor U42820 (N_42820,N_41010,N_40382);
or U42821 (N_42821,N_40964,N_41169);
nand U42822 (N_42822,N_40327,N_41823);
nand U42823 (N_42823,N_42075,N_41114);
nand U42824 (N_42824,N_41476,N_40618);
nor U42825 (N_42825,N_42181,N_42081);
nand U42826 (N_42826,N_40667,N_40007);
and U42827 (N_42827,N_41463,N_41292);
nand U42828 (N_42828,N_40595,N_42324);
nand U42829 (N_42829,N_40659,N_41282);
xnor U42830 (N_42830,N_40881,N_40612);
nor U42831 (N_42831,N_40798,N_41649);
or U42832 (N_42832,N_41364,N_40283);
nand U42833 (N_42833,N_42432,N_41922);
xor U42834 (N_42834,N_41766,N_41839);
or U42835 (N_42835,N_40053,N_41411);
and U42836 (N_42836,N_41682,N_40768);
nand U42837 (N_42837,N_42490,N_42187);
and U42838 (N_42838,N_41342,N_40558);
nor U42839 (N_42839,N_40158,N_40981);
and U42840 (N_42840,N_41496,N_41596);
xor U42841 (N_42841,N_40921,N_40350);
nor U42842 (N_42842,N_41562,N_41005);
nor U42843 (N_42843,N_40693,N_41673);
and U42844 (N_42844,N_41118,N_41923);
xor U42845 (N_42845,N_40796,N_41524);
or U42846 (N_42846,N_40409,N_41020);
and U42847 (N_42847,N_41595,N_40619);
xor U42848 (N_42848,N_41281,N_40341);
nor U42849 (N_42849,N_40657,N_40085);
nor U42850 (N_42850,N_42096,N_41491);
or U42851 (N_42851,N_41879,N_41988);
xor U42852 (N_42852,N_41081,N_41832);
nand U42853 (N_42853,N_40708,N_40118);
xor U42854 (N_42854,N_42421,N_42251);
or U42855 (N_42855,N_41030,N_41326);
or U42856 (N_42856,N_40915,N_40715);
and U42857 (N_42857,N_41154,N_42060);
and U42858 (N_42858,N_41239,N_41363);
and U42859 (N_42859,N_41441,N_42258);
xor U42860 (N_42860,N_40406,N_42334);
and U42861 (N_42861,N_40035,N_42286);
or U42862 (N_42862,N_41141,N_42397);
or U42863 (N_42863,N_41064,N_42291);
xnor U42864 (N_42864,N_41608,N_40243);
xnor U42865 (N_42865,N_41058,N_42013);
nand U42866 (N_42866,N_41115,N_41556);
or U42867 (N_42867,N_42062,N_40019);
or U42868 (N_42868,N_41864,N_41356);
and U42869 (N_42869,N_41842,N_42226);
and U42870 (N_42870,N_41566,N_41085);
xor U42871 (N_42871,N_40891,N_40232);
and U42872 (N_42872,N_41004,N_42278);
xor U42873 (N_42873,N_42467,N_42007);
and U42874 (N_42874,N_41504,N_40702);
or U42875 (N_42875,N_41107,N_41389);
xor U42876 (N_42876,N_41045,N_42442);
nor U42877 (N_42877,N_42494,N_40257);
or U42878 (N_42878,N_42164,N_42100);
nor U42879 (N_42879,N_40689,N_41899);
nand U42880 (N_42880,N_40837,N_40102);
and U42881 (N_42881,N_40952,N_40519);
or U42882 (N_42882,N_40082,N_41701);
nor U42883 (N_42883,N_41272,N_41980);
xnor U42884 (N_42884,N_41061,N_40685);
or U42885 (N_42885,N_41472,N_41497);
and U42886 (N_42886,N_41113,N_40542);
and U42887 (N_42887,N_40666,N_40272);
xnor U42888 (N_42888,N_41884,N_40673);
or U42889 (N_42889,N_42042,N_41172);
xor U42890 (N_42890,N_42329,N_40172);
nand U42891 (N_42891,N_41626,N_41456);
nand U42892 (N_42892,N_41032,N_40813);
and U42893 (N_42893,N_41029,N_40622);
or U42894 (N_42894,N_40580,N_40349);
and U42895 (N_42895,N_41696,N_40606);
xor U42896 (N_42896,N_40476,N_41066);
and U42897 (N_42897,N_42491,N_40002);
nand U42898 (N_42898,N_40104,N_40106);
xor U42899 (N_42899,N_40131,N_42136);
nor U42900 (N_42900,N_41803,N_41328);
or U42901 (N_42901,N_41257,N_40344);
xnor U42902 (N_42902,N_41403,N_40803);
nor U42903 (N_42903,N_41293,N_42126);
nand U42904 (N_42904,N_40237,N_41191);
nor U42905 (N_42905,N_42447,N_42076);
xor U42906 (N_42906,N_40291,N_40225);
xnor U42907 (N_42907,N_40054,N_40411);
nor U42908 (N_42908,N_40398,N_41972);
xnor U42909 (N_42909,N_40400,N_42008);
and U42910 (N_42910,N_42194,N_41577);
xnor U42911 (N_42911,N_42449,N_40055);
nand U42912 (N_42912,N_42327,N_41351);
xnor U42913 (N_42913,N_41904,N_40948);
nor U42914 (N_42914,N_40600,N_42287);
or U42915 (N_42915,N_40895,N_40408);
or U42916 (N_42916,N_41951,N_42412);
nand U42917 (N_42917,N_41943,N_42482);
nand U42918 (N_42918,N_40867,N_41807);
nand U42919 (N_42919,N_41617,N_41451);
nand U42920 (N_42920,N_40974,N_41945);
or U42921 (N_42921,N_40439,N_40577);
or U42922 (N_42922,N_42470,N_40751);
xor U42923 (N_42923,N_40701,N_41253);
and U42924 (N_42924,N_40008,N_40256);
nor U42925 (N_42925,N_40049,N_40358);
and U42926 (N_42926,N_40674,N_41036);
nand U42927 (N_42927,N_42063,N_40505);
xnor U42928 (N_42928,N_42264,N_40425);
xnor U42929 (N_42929,N_41655,N_41551);
or U42930 (N_42930,N_40484,N_42069);
xnor U42931 (N_42931,N_40596,N_42012);
nand U42932 (N_42932,N_40557,N_41633);
and U42933 (N_42933,N_42370,N_42303);
and U42934 (N_42934,N_40820,N_40133);
and U42935 (N_42935,N_41157,N_40928);
or U42936 (N_42936,N_41329,N_41466);
or U42937 (N_42937,N_41309,N_40521);
nor U42938 (N_42938,N_41920,N_40879);
xnor U42939 (N_42939,N_42294,N_40296);
and U42940 (N_42940,N_42290,N_42022);
xor U42941 (N_42941,N_41687,N_41775);
nand U42942 (N_42942,N_40307,N_41231);
nand U42943 (N_42943,N_41479,N_40669);
xnor U42944 (N_42944,N_42462,N_40553);
nand U42945 (N_42945,N_41439,N_42375);
nand U42946 (N_42946,N_40242,N_40767);
nand U42947 (N_42947,N_40027,N_41700);
or U42948 (N_42948,N_41727,N_42162);
and U42949 (N_42949,N_42325,N_41162);
nand U42950 (N_42950,N_40009,N_41850);
xor U42951 (N_42951,N_42137,N_41269);
nand U42952 (N_42952,N_40437,N_42209);
and U42953 (N_42953,N_40937,N_41751);
xor U42954 (N_42954,N_42201,N_40261);
or U42955 (N_42955,N_41643,N_40543);
nor U42956 (N_42956,N_42131,N_41431);
and U42957 (N_42957,N_41549,N_40238);
xnor U42958 (N_42958,N_40934,N_42252);
nand U42959 (N_42959,N_41977,N_40097);
nor U42960 (N_42960,N_40828,N_40985);
xor U42961 (N_42961,N_42435,N_41893);
xor U42962 (N_42962,N_41789,N_40005);
nor U42963 (N_42963,N_40978,N_41421);
nor U42964 (N_42964,N_40638,N_40488);
and U42965 (N_42965,N_42422,N_42185);
nor U42966 (N_42966,N_42204,N_40467);
or U42967 (N_42967,N_41312,N_41845);
nor U42968 (N_42968,N_40736,N_41109);
and U42969 (N_42969,N_40091,N_41009);
or U42970 (N_42970,N_40479,N_40115);
nor U42971 (N_42971,N_40380,N_41974);
and U42972 (N_42972,N_40208,N_41499);
nand U42973 (N_42973,N_40579,N_42273);
and U42974 (N_42974,N_41507,N_40012);
nand U42975 (N_42975,N_40965,N_40805);
and U42976 (N_42976,N_41396,N_41178);
nor U42977 (N_42977,N_40849,N_41801);
or U42978 (N_42978,N_41989,N_42307);
nand U42979 (N_42979,N_42052,N_42341);
or U42980 (N_42980,N_40363,N_41318);
nor U42981 (N_42981,N_40422,N_40954);
xnor U42982 (N_42982,N_42426,N_41171);
nor U42983 (N_42983,N_40597,N_41830);
nor U42984 (N_42984,N_42039,N_41982);
and U42985 (N_42985,N_42340,N_40554);
and U42986 (N_42986,N_41375,N_40695);
nor U42987 (N_42987,N_42032,N_40546);
nor U42988 (N_42988,N_40493,N_42099);
nor U42989 (N_42989,N_42302,N_40340);
nand U42990 (N_42990,N_41205,N_41233);
nand U42991 (N_42991,N_40424,N_40599);
nand U42992 (N_42992,N_42104,N_40023);
nand U42993 (N_42993,N_40194,N_40995);
or U42994 (N_42994,N_41317,N_40404);
and U42995 (N_42995,N_40980,N_42198);
and U42996 (N_42996,N_40329,N_42077);
and U42997 (N_42997,N_40432,N_40218);
xor U42998 (N_42998,N_42309,N_40077);
nand U42999 (N_42999,N_40083,N_41276);
and U43000 (N_43000,N_41056,N_41196);
nor U43001 (N_43001,N_40065,N_41736);
xor U43002 (N_43002,N_40740,N_40646);
and U43003 (N_43003,N_41136,N_42024);
or U43004 (N_43004,N_40642,N_41949);
nand U43005 (N_43005,N_41946,N_42332);
nand U43006 (N_43006,N_41216,N_40832);
or U43007 (N_43007,N_40940,N_41265);
xor U43008 (N_43008,N_42256,N_41143);
or U43009 (N_43009,N_41393,N_42152);
and U43010 (N_43010,N_42125,N_41345);
nand U43011 (N_43011,N_42419,N_41111);
xnor U43012 (N_43012,N_40146,N_40753);
nand U43013 (N_43013,N_41814,N_40336);
nand U43014 (N_43014,N_41075,N_40401);
xnor U43015 (N_43015,N_40316,N_42311);
nor U43016 (N_43016,N_41409,N_40231);
and U43017 (N_43017,N_41716,N_42103);
or U43018 (N_43018,N_41638,N_40905);
nor U43019 (N_43019,N_42049,N_42167);
nor U43020 (N_43020,N_42343,N_40770);
nor U43021 (N_43021,N_40714,N_42179);
nor U43022 (N_43022,N_41519,N_41185);
nor U43023 (N_43023,N_41271,N_40258);
nand U43024 (N_43024,N_41878,N_40524);
nand U43025 (N_43025,N_41571,N_40722);
nor U43026 (N_43026,N_40688,N_41758);
nand U43027 (N_43027,N_41827,N_42392);
xnor U43028 (N_43028,N_42195,N_41268);
nand U43029 (N_43029,N_41660,N_42322);
nand U43030 (N_43030,N_40752,N_42439);
nor U43031 (N_43031,N_41854,N_41362);
and U43032 (N_43032,N_41728,N_41734);
nand U43033 (N_43033,N_40914,N_40188);
nand U43034 (N_43034,N_40804,N_41936);
nor U43035 (N_43035,N_42437,N_42051);
or U43036 (N_43036,N_42274,N_40620);
or U43037 (N_43037,N_40311,N_40760);
xnor U43038 (N_43038,N_40073,N_42030);
nand U43039 (N_43039,N_41960,N_40364);
and U43040 (N_43040,N_41970,N_41199);
or U43041 (N_43041,N_41433,N_42154);
nand U43042 (N_43042,N_40861,N_42314);
or U43043 (N_43043,N_40545,N_40802);
or U43044 (N_43044,N_42479,N_40966);
or U43045 (N_43045,N_40502,N_41442);
nor U43046 (N_43046,N_41933,N_41251);
and U43047 (N_43047,N_42276,N_42331);
nand U43048 (N_43048,N_42206,N_40361);
xnor U43049 (N_43049,N_40348,N_42268);
nand U43050 (N_43050,N_40834,N_40021);
xnor U43051 (N_43051,N_41699,N_40938);
and U43052 (N_43052,N_40792,N_41177);
xor U43053 (N_43053,N_41929,N_40119);
or U43054 (N_43054,N_42300,N_41767);
nand U43055 (N_43055,N_41469,N_41511);
nand U43056 (N_43056,N_40679,N_41860);
nand U43057 (N_43057,N_41140,N_41160);
nand U43058 (N_43058,N_41825,N_41055);
xor U43059 (N_43059,N_40894,N_40187);
nor U43060 (N_43060,N_41645,N_41420);
or U43061 (N_43061,N_42135,N_40687);
xor U43062 (N_43062,N_41739,N_41971);
or U43063 (N_43063,N_40840,N_42180);
nand U43064 (N_43064,N_42066,N_41395);
nor U43065 (N_43065,N_40947,N_40850);
and U43066 (N_43066,N_42356,N_42106);
and U43067 (N_43067,N_42101,N_42446);
nand U43068 (N_43068,N_40556,N_41555);
and U43069 (N_43069,N_41014,N_41381);
nor U43070 (N_43070,N_42497,N_41713);
or U43071 (N_43071,N_42450,N_41572);
xnor U43072 (N_43072,N_42436,N_41394);
nand U43073 (N_43073,N_42067,N_41932);
xnor U43074 (N_43074,N_40059,N_40174);
or U43075 (N_43075,N_40729,N_40100);
nor U43076 (N_43076,N_41071,N_42149);
or U43077 (N_43077,N_41390,N_41203);
nand U43078 (N_43078,N_41226,N_41073);
xor U43079 (N_43079,N_40293,N_40993);
xnor U43080 (N_43080,N_41086,N_41280);
xnor U43081 (N_43081,N_41132,N_41635);
nor U43082 (N_43082,N_40339,N_41028);
xnor U43083 (N_43083,N_40678,N_40285);
and U43084 (N_43084,N_40374,N_42184);
or U43085 (N_43085,N_41026,N_40384);
and U43086 (N_43086,N_41546,N_42480);
and U43087 (N_43087,N_41848,N_40395);
nand U43088 (N_43088,N_40292,N_41021);
or U43089 (N_43089,N_41290,N_41208);
xnor U43090 (N_43090,N_41622,N_40639);
and U43091 (N_43091,N_42144,N_40338);
xor U43092 (N_43092,N_41793,N_40741);
nor U43093 (N_43093,N_41335,N_41684);
nor U43094 (N_43094,N_40371,N_40089);
nor U43095 (N_43095,N_40649,N_41386);
xor U43096 (N_43096,N_40281,N_41875);
nor U43097 (N_43097,N_41101,N_42233);
nor U43098 (N_43098,N_41354,N_42339);
nor U43099 (N_43099,N_40359,N_41954);
and U43100 (N_43100,N_42487,N_41672);
nor U43101 (N_43101,N_41378,N_41173);
and U43102 (N_43102,N_40202,N_41935);
nand U43103 (N_43103,N_42190,N_40212);
nand U43104 (N_43104,N_41052,N_40853);
xor U43105 (N_43105,N_41819,N_41625);
nor U43106 (N_43106,N_41127,N_41158);
or U43107 (N_43107,N_40656,N_42222);
xor U43108 (N_43108,N_40951,N_41650);
xnor U43109 (N_43109,N_40162,N_40132);
and U43110 (N_43110,N_41678,N_40180);
and U43111 (N_43111,N_41631,N_41611);
and U43112 (N_43112,N_42014,N_41230);
or U43113 (N_43113,N_40912,N_40691);
and U43114 (N_43114,N_40953,N_40987);
nand U43115 (N_43115,N_40529,N_42061);
or U43116 (N_43116,N_40784,N_40254);
and U43117 (N_43117,N_42481,N_41457);
or U43118 (N_43118,N_41692,N_41474);
or U43119 (N_43119,N_41768,N_41338);
nand U43120 (N_43120,N_41054,N_40223);
and U43121 (N_43121,N_41437,N_41530);
or U43122 (N_43122,N_41831,N_40075);
and U43123 (N_43123,N_42087,N_40390);
nor U43124 (N_43124,N_42092,N_41992);
nor U43125 (N_43125,N_40516,N_40028);
xnor U43126 (N_43126,N_40394,N_40078);
and U43127 (N_43127,N_42241,N_41348);
or U43128 (N_43128,N_42372,N_40284);
and U43129 (N_43129,N_42085,N_40241);
nor U43130 (N_43130,N_41145,N_41480);
or U43131 (N_43131,N_42424,N_40137);
xnor U43132 (N_43132,N_40913,N_40407);
xor U43133 (N_43133,N_41953,N_42471);
nor U43134 (N_43134,N_41896,N_40845);
nand U43135 (N_43135,N_40200,N_40130);
nand U43136 (N_43136,N_42237,N_41986);
nor U43137 (N_43137,N_41489,N_41719);
and U43138 (N_43138,N_40416,N_41218);
nand U43139 (N_43139,N_41192,N_40320);
nor U43140 (N_43140,N_40094,N_41383);
and U43141 (N_43141,N_41287,N_41483);
xor U43142 (N_43142,N_42378,N_41427);
nand U43143 (N_43143,N_40607,N_40255);
nand U43144 (N_43144,N_41913,N_41501);
and U43145 (N_43145,N_41762,N_41720);
xor U43146 (N_43146,N_42120,N_41011);
nor U43147 (N_43147,N_42065,N_41520);
nor U43148 (N_43148,N_40635,N_41144);
nand U43149 (N_43149,N_40960,N_42047);
nand U43150 (N_43150,N_42305,N_41575);
xor U43151 (N_43151,N_41586,N_40530);
nor U43152 (N_43152,N_41304,N_40275);
or U43153 (N_43153,N_40108,N_42098);
nor U43154 (N_43154,N_41732,N_41634);
nor U43155 (N_43155,N_40217,N_41658);
xnor U43156 (N_43156,N_41704,N_41604);
xnor U43157 (N_43157,N_42046,N_42253);
xnor U43158 (N_43158,N_40806,N_40322);
xnor U43159 (N_43159,N_40963,N_40696);
nor U43160 (N_43160,N_40229,N_40812);
xor U43161 (N_43161,N_41755,N_41024);
and U43162 (N_43162,N_41018,N_41310);
or U43163 (N_43163,N_42157,N_42308);
nor U43164 (N_43164,N_40201,N_42228);
and U43165 (N_43165,N_41138,N_40236);
and U43166 (N_43166,N_41041,N_40923);
or U43167 (N_43167,N_42186,N_41710);
or U43168 (N_43168,N_40598,N_40280);
nand U43169 (N_43169,N_42385,N_41891);
and U43170 (N_43170,N_40637,N_40173);
nor U43171 (N_43171,N_40471,N_42035);
xnor U43172 (N_43172,N_41999,N_41297);
and U43173 (N_43173,N_41358,N_42472);
or U43174 (N_43174,N_41125,N_42454);
nand U43175 (N_43175,N_41843,N_40641);
or U43176 (N_43176,N_42083,N_40875);
nor U43177 (N_43177,N_40228,N_41462);
xor U43178 (N_43178,N_42338,N_42108);
xor U43179 (N_43179,N_41607,N_42394);
and U43180 (N_43180,N_42169,N_42213);
nand U43181 (N_43181,N_42434,N_41336);
nand U43182 (N_43182,N_40182,N_42451);
nand U43183 (N_43183,N_42475,N_40650);
nand U43184 (N_43184,N_41869,N_40510);
nor U43185 (N_43185,N_40308,N_40744);
nor U43186 (N_43186,N_40540,N_41538);
nor U43187 (N_43187,N_41159,N_41683);
and U43188 (N_43188,N_41099,N_40436);
or U43189 (N_43189,N_41067,N_41370);
nand U43190 (N_43190,N_40459,N_40671);
nor U43191 (N_43191,N_41308,N_40190);
or U43192 (N_43192,N_42026,N_40388);
nand U43193 (N_43193,N_40393,N_40712);
nand U43194 (N_43194,N_41373,N_41835);
nor U43195 (N_43195,N_40209,N_40234);
nand U43196 (N_43196,N_42216,N_40314);
nor U43197 (N_43197,N_41578,N_40778);
or U43198 (N_43198,N_41357,N_41273);
xor U43199 (N_43199,N_40464,N_41096);
xnor U43200 (N_43200,N_40544,N_40907);
xor U43201 (N_43201,N_41498,N_41653);
and U43202 (N_43202,N_42292,N_42265);
xor U43203 (N_43203,N_41554,N_41870);
nor U43204 (N_43204,N_40026,N_41939);
and U43205 (N_43205,N_40472,N_41969);
xnor U43206 (N_43206,N_41780,N_40833);
or U43207 (N_43207,N_42371,N_40103);
or U43208 (N_43208,N_41616,N_41890);
nor U43209 (N_43209,N_41564,N_41106);
nand U43210 (N_43210,N_40305,N_42140);
nand U43211 (N_43211,N_40481,N_40831);
and U43212 (N_43212,N_41110,N_40636);
and U43213 (N_43213,N_40014,N_42382);
and U43214 (N_43214,N_41130,N_41065);
nor U43215 (N_43215,N_42318,N_42349);
nand U43216 (N_43216,N_42433,N_41804);
nand U43217 (N_43217,N_42202,N_42005);
and U43218 (N_43218,N_41863,N_42127);
and U43219 (N_43219,N_41412,N_41180);
nand U43220 (N_43220,N_41376,N_41374);
or U43221 (N_43221,N_42102,N_42088);
nor U43222 (N_43222,N_42384,N_42469);
and U43223 (N_43223,N_40165,N_42212);
xor U43224 (N_43224,N_41038,N_41436);
nand U43225 (N_43225,N_41769,N_40817);
xnor U43226 (N_43226,N_41063,N_41761);
and U43227 (N_43227,N_40655,N_40313);
xor U43228 (N_43228,N_40274,N_40956);
xnor U43229 (N_43229,N_40303,N_41748);
or U43230 (N_43230,N_40037,N_41756);
xor U43231 (N_43231,N_41232,N_40992);
nor U43232 (N_43232,N_41553,N_41510);
nand U43233 (N_43233,N_41248,N_40765);
nor U43234 (N_43234,N_40941,N_41262);
nor U43235 (N_43235,N_42027,N_41770);
nand U43236 (N_43236,N_42496,N_41306);
nor U43237 (N_43237,N_40929,N_40511);
or U43238 (N_43238,N_42150,N_40625);
xnor U43239 (N_43239,N_42417,N_40092);
xor U43240 (N_43240,N_40660,N_40483);
nand U43241 (N_43241,N_41952,N_41380);
nor U43242 (N_43242,N_42492,N_40555);
or U43243 (N_43243,N_40489,N_40161);
or U43244 (N_43244,N_40170,N_41905);
or U43245 (N_43245,N_40051,N_40719);
and U43246 (N_43246,N_42477,N_42072);
and U43247 (N_43247,N_40533,N_40273);
nand U43248 (N_43248,N_42029,N_41917);
nand U43249 (N_43249,N_41093,N_40042);
xnor U43250 (N_43250,N_40663,N_40150);
and U43251 (N_43251,N_41747,N_40758);
or U43252 (N_43252,N_42306,N_40552);
and U43253 (N_43253,N_41754,N_40109);
or U43254 (N_43254,N_41128,N_42165);
nand U43255 (N_43255,N_40576,N_41918);
xor U43256 (N_43256,N_41664,N_42122);
nor U43257 (N_43257,N_40925,N_41214);
xnor U43258 (N_43258,N_42484,N_41135);
xnor U43259 (N_43259,N_41708,N_40289);
or U43260 (N_43260,N_41076,N_42159);
nor U43261 (N_43261,N_40375,N_40664);
nor U43262 (N_43262,N_41417,N_42452);
nand U43263 (N_43263,N_40105,N_41500);
nor U43264 (N_43264,N_40022,N_41189);
and U43265 (N_43265,N_40571,N_40298);
and U43266 (N_43266,N_41049,N_40240);
xnor U43267 (N_43267,N_41648,N_41087);
nand U43268 (N_43268,N_41593,N_40470);
nor U43269 (N_43269,N_42090,N_40048);
or U43270 (N_43270,N_40276,N_42431);
nor U43271 (N_43271,N_40969,N_40302);
or U43272 (N_43272,N_40018,N_41270);
nand U43273 (N_43273,N_40301,N_42214);
and U43274 (N_43274,N_40868,N_42246);
and U43275 (N_43275,N_41147,N_42016);
nand U43276 (N_43276,N_41889,N_41996);
and U43277 (N_43277,N_40582,N_42390);
nor U43278 (N_43278,N_40628,N_40950);
or U43279 (N_43279,N_41314,N_40626);
or U43280 (N_43280,N_40367,N_40135);
nor U43281 (N_43281,N_40774,N_41680);
nor U43282 (N_43282,N_42403,N_40904);
nand U43283 (N_43283,N_41369,N_40829);
nor U43284 (N_43284,N_41764,N_42270);
and U43285 (N_43285,N_40591,N_41344);
xnor U43286 (N_43286,N_42174,N_41967);
or U43287 (N_43287,N_41098,N_42070);
nor U43288 (N_43288,N_41371,N_40043);
or U43289 (N_43289,N_41866,N_42082);
and U43290 (N_43290,N_40509,N_42191);
xnor U43291 (N_43291,N_40462,N_41247);
nor U43292 (N_43292,N_41785,N_41797);
and U43293 (N_43293,N_40759,N_40052);
nor U43294 (N_43294,N_42295,N_41430);
nor U43295 (N_43295,N_41166,N_40675);
nand U43296 (N_43296,N_41824,N_40264);
xor U43297 (N_43297,N_40445,N_42298);
and U43298 (N_43298,N_42266,N_40244);
and U43299 (N_43299,N_41925,N_41170);
nor U43300 (N_43300,N_40443,N_40949);
xnor U43301 (N_43301,N_40379,N_41195);
nand U43302 (N_43302,N_41895,N_40139);
and U43303 (N_43303,N_40790,N_41129);
or U43304 (N_43304,N_40512,N_41346);
xnor U43305 (N_43305,N_41360,N_40057);
or U43306 (N_43306,N_41187,N_41298);
or U43307 (N_43307,N_41791,N_42400);
nand U43308 (N_43308,N_41569,N_41963);
or U43309 (N_43309,N_42146,N_40321);
or U43310 (N_43310,N_42468,N_42427);
or U43311 (N_43311,N_42310,N_41686);
nand U43312 (N_43312,N_41488,N_42498);
and U43313 (N_43313,N_40124,N_40793);
nand U43314 (N_43314,N_40842,N_41816);
or U43315 (N_43315,N_40178,N_40794);
or U43316 (N_43316,N_42260,N_40843);
and U43317 (N_43317,N_42396,N_42175);
nand U43318 (N_43318,N_42192,N_42402);
or U43319 (N_43319,N_41382,N_42009);
nand U43320 (N_43320,N_40996,N_42383);
nand U43321 (N_43321,N_40290,N_40998);
and U43322 (N_43322,N_40608,N_41148);
xnor U43323 (N_43323,N_42254,N_42353);
or U43324 (N_43324,N_41534,N_42203);
or U43325 (N_43325,N_42326,N_40906);
xor U43326 (N_43326,N_41950,N_41017);
xnor U43327 (N_43327,N_40824,N_41023);
nor U43328 (N_43328,N_41544,N_41175);
and U43329 (N_43329,N_40498,N_40640);
nand U43330 (N_43330,N_40345,N_41150);
or U43331 (N_43331,N_40006,N_40968);
and U43332 (N_43332,N_42461,N_40431);
xor U43333 (N_43333,N_40976,N_42172);
and U43334 (N_43334,N_42364,N_40683);
nor U43335 (N_43335,N_40504,N_40183);
nor U43336 (N_43336,N_40233,N_40944);
nand U43337 (N_43337,N_41630,N_41709);
xor U43338 (N_43338,N_40265,N_40475);
or U43339 (N_43339,N_40247,N_40356);
and U43340 (N_43340,N_40171,N_41492);
nand U43341 (N_43341,N_41209,N_41176);
and U43342 (N_43342,N_41885,N_41112);
or U43343 (N_43343,N_41641,N_42352);
and U43344 (N_43344,N_41533,N_42188);
or U43345 (N_43345,N_40392,N_40154);
xor U43346 (N_43346,N_40045,N_42389);
nor U43347 (N_43347,N_41414,N_40175);
and U43348 (N_43348,N_41243,N_41302);
or U43349 (N_43349,N_41606,N_40206);
xor U43350 (N_43350,N_40376,N_41523);
and U43351 (N_43351,N_40900,N_40351);
and U43352 (N_43352,N_40534,N_41778);
or U43353 (N_43353,N_40360,N_41959);
and U43354 (N_43354,N_40629,N_42418);
and U43355 (N_43355,N_41627,N_41588);
or U43356 (N_43356,N_42232,N_40215);
nor U43357 (N_43357,N_40706,N_40957);
and U43358 (N_43358,N_41938,N_41817);
nor U43359 (N_43359,N_42367,N_41725);
xnor U43360 (N_43360,N_41671,N_41773);
xor U43361 (N_43361,N_41846,N_41407);
xnor U43362 (N_43362,N_40830,N_40386);
nand U43363 (N_43363,N_41735,N_40086);
or U43364 (N_43364,N_41258,N_41082);
xor U43365 (N_43365,N_41539,N_40601);
xnor U43366 (N_43366,N_41255,N_40846);
and U43367 (N_43367,N_41729,N_40024);
nand U43368 (N_43368,N_40791,N_41615);
and U43369 (N_43369,N_41339,N_40144);
nor U43370 (N_43370,N_41083,N_42017);
nor U43371 (N_43371,N_40624,N_40880);
and U43372 (N_43372,N_40621,N_41123);
xor U43373 (N_43373,N_41465,N_41940);
nor U43374 (N_43374,N_41540,N_42227);
or U43375 (N_43375,N_41320,N_40486);
nor U43376 (N_43376,N_42078,N_40143);
nand U43377 (N_43377,N_41568,N_40199);
nand U43378 (N_43378,N_41976,N_42284);
nor U43379 (N_43379,N_40783,N_42004);
nor U43380 (N_43380,N_41613,N_42112);
xor U43381 (N_43381,N_41792,N_42097);
nor U43382 (N_43382,N_41337,N_40808);
nor U43383 (N_43383,N_41485,N_42410);
xor U43384 (N_43384,N_40138,N_42489);
nor U43385 (N_43385,N_41235,N_41921);
or U43386 (N_43386,N_41202,N_41558);
nor U43387 (N_43387,N_41493,N_40309);
nand U43388 (N_43388,N_41543,N_40762);
xor U43389 (N_43389,N_42361,N_42235);
and U43390 (N_43390,N_41669,N_41197);
xnor U43391 (N_43391,N_40851,N_42215);
or U43392 (N_43392,N_41261,N_41517);
or U43393 (N_43393,N_41392,N_41325);
xnor U43394 (N_43394,N_40453,N_41327);
xor U43395 (N_43395,N_42262,N_42381);
or U43396 (N_43396,N_40219,N_40855);
and U43397 (N_43397,N_41372,N_41800);
or U43398 (N_43398,N_40074,N_40378);
nand U43399 (N_43399,N_41513,N_40157);
xnor U43400 (N_43400,N_41828,N_41930);
xor U43401 (N_43401,N_42089,N_41508);
and U43402 (N_43402,N_40716,N_42399);
nand U43403 (N_43403,N_41019,N_40991);
nand U43404 (N_43404,N_40365,N_41901);
nand U43405 (N_43405,N_40186,N_42132);
and U43406 (N_43406,N_40069,N_40869);
nor U43407 (N_43407,N_41245,N_42234);
nor U43408 (N_43408,N_41602,N_42094);
or U43409 (N_43409,N_40593,N_40508);
and U43410 (N_43410,N_40737,N_42095);
xnor U43411 (N_43411,N_40988,N_40153);
nand U43412 (N_43412,N_42415,N_42025);
xnor U43413 (N_43413,N_42376,N_40156);
or U43414 (N_43414,N_40203,N_40742);
xnor U43415 (N_43415,N_42139,N_42115);
nand U43416 (N_43416,N_41012,N_41847);
nor U43417 (N_43417,N_41153,N_41644);
nor U43418 (N_43418,N_40893,N_40728);
or U43419 (N_43419,N_41926,N_41599);
xor U43420 (N_43420,N_41528,N_42401);
xor U43421 (N_43421,N_40780,N_40177);
xor U43422 (N_43422,N_41043,N_40686);
or U43423 (N_43423,N_40549,N_42020);
nor U43424 (N_43424,N_40342,N_40967);
nor U43425 (N_43425,N_41164,N_40410);
or U43426 (N_43426,N_41256,N_40971);
nor U43427 (N_43427,N_40050,N_41167);
xor U43428 (N_43428,N_40801,N_40863);
xnor U43429 (N_43429,N_41927,N_40899);
nor U43430 (N_43430,N_40816,N_41227);
nand U43431 (N_43431,N_42156,N_40495);
nand U43432 (N_43432,N_42166,N_41993);
or U43433 (N_43433,N_42073,N_41537);
or U43434 (N_43434,N_41880,N_41573);
nor U43435 (N_43435,N_42036,N_42023);
nor U43436 (N_43436,N_41877,N_41088);
nand U43437 (N_43437,N_41188,N_40079);
nor U43438 (N_43438,N_41238,N_41134);
nand U43439 (N_43439,N_40918,N_41894);
or U43440 (N_43440,N_41750,N_42293);
nor U43441 (N_43441,N_40800,N_40207);
or U43442 (N_43442,N_42001,N_40438);
or U43443 (N_43443,N_40587,N_41639);
nor U43444 (N_43444,N_40224,N_40474);
and U43445 (N_43445,N_40535,N_40525);
or U43446 (N_43446,N_41567,N_40332);
nand U43447 (N_43447,N_41016,N_40337);
nand U43448 (N_43448,N_41542,N_41091);
or U43449 (N_43449,N_42028,N_41771);
and U43450 (N_43450,N_40128,N_42053);
xor U43451 (N_43451,N_42040,N_40096);
or U43452 (N_43452,N_41039,N_41979);
nand U43453 (N_43453,N_41663,N_40644);
and U43454 (N_43454,N_41122,N_40084);
xnor U43455 (N_43455,N_41948,N_41737);
and U43456 (N_43456,N_40413,N_41916);
nand U43457 (N_43457,N_41048,N_40731);
and U43458 (N_43458,N_42211,N_41964);
or U43459 (N_43459,N_42041,N_41574);
nor U43460 (N_43460,N_40330,N_40482);
nor U43461 (N_43461,N_40757,N_40029);
and U43462 (N_43462,N_40724,N_41861);
xor U43463 (N_43463,N_40747,N_40878);
or U43464 (N_43464,N_40970,N_42044);
nor U43465 (N_43465,N_40665,N_42285);
or U43466 (N_43466,N_41956,N_42138);
or U43467 (N_43467,N_40975,N_40602);
or U43468 (N_43468,N_40494,N_42320);
nor U43469 (N_43469,N_41350,N_42330);
nand U43470 (N_43470,N_41051,N_41156);
and U43471 (N_43471,N_42247,N_41514);
nand U43472 (N_43472,N_40563,N_40500);
nor U43473 (N_43473,N_40572,N_41092);
or U43474 (N_43474,N_41690,N_42151);
and U43475 (N_43475,N_40852,N_41619);
nand U43476 (N_43476,N_42296,N_40578);
nand U43477 (N_43477,N_40469,N_42057);
nand U43478 (N_43478,N_41080,N_40692);
xnor U43479 (N_43479,N_41966,N_40428);
or U43480 (N_43480,N_41749,N_41155);
or U43481 (N_43481,N_40699,N_41397);
and U43482 (N_43482,N_42158,N_41621);
or U43483 (N_43483,N_40584,N_42279);
or U43484 (N_43484,N_40402,N_40575);
xor U43485 (N_43485,N_41799,N_41174);
or U43486 (N_43486,N_42121,N_42031);
and U43487 (N_43487,N_41206,N_41322);
nand U43488 (N_43488,N_40903,N_40497);
or U43489 (N_43489,N_41377,N_41654);
and U43490 (N_43490,N_40081,N_40697);
nand U43491 (N_43491,N_42245,N_40121);
xnor U43492 (N_43492,N_41408,N_41906);
and U43493 (N_43493,N_42168,N_40310);
xnor U43494 (N_43494,N_42116,N_42119);
or U43495 (N_43495,N_40926,N_40877);
xnor U43496 (N_43496,N_40211,N_40230);
xnor U43497 (N_43497,N_41527,N_40168);
and U43498 (N_43498,N_40743,N_41689);
nor U43499 (N_43499,N_41471,N_41385);
xnor U43500 (N_43500,N_42068,N_40013);
or U43501 (N_43501,N_42344,N_40583);
nor U43502 (N_43502,N_42267,N_42428);
xnor U43503 (N_43503,N_40795,N_41502);
nor U43504 (N_43504,N_41212,N_40836);
xnor U43505 (N_43505,N_41547,N_41089);
xnor U43506 (N_43506,N_40797,N_40099);
or U43507 (N_43507,N_42485,N_41841);
or U43508 (N_43508,N_41973,N_41401);
nand U43509 (N_43509,N_40490,N_42360);
or U43510 (N_43510,N_41600,N_40694);
or U43511 (N_43511,N_41211,N_42058);
nor U43512 (N_43512,N_40605,N_40333);
and U43513 (N_43513,N_41044,N_40559);
nand U43514 (N_43514,N_42002,N_40908);
xor U43515 (N_43515,N_40973,N_40352);
nor U43516 (N_43516,N_41460,N_42080);
nor U43517 (N_43517,N_40672,N_40614);
xnor U43518 (N_43518,N_40933,N_41612);
nand U43519 (N_43519,N_40827,N_40235);
and U43520 (N_43520,N_41691,N_41531);
or U43521 (N_43521,N_42160,N_41694);
nand U43522 (N_43522,N_40574,N_41416);
nand U43523 (N_43523,N_40456,N_41795);
nand U43524 (N_43524,N_40866,N_40847);
xor U43525 (N_43525,N_40080,N_41072);
xor U43526 (N_43526,N_41871,N_40732);
and U43527 (N_43527,N_40433,N_41656);
xnor U43528 (N_43528,N_41698,N_42218);
nor U43529 (N_43529,N_42488,N_41490);
nand U43530 (N_43530,N_42416,N_40911);
xor U43531 (N_43531,N_41246,N_42117);
nand U43532 (N_43532,N_41536,N_41448);
and U43533 (N_43533,N_41815,N_40739);
or U43534 (N_43534,N_41784,N_40864);
xnor U43535 (N_43535,N_41503,N_42407);
nand U43536 (N_43536,N_42362,N_41284);
xnor U43537 (N_43537,N_40142,N_41445);
xor U43538 (N_43538,N_41379,N_41025);
nand U43539 (N_43539,N_41330,N_40056);
xnor U43540 (N_43540,N_40101,N_40643);
xor U43541 (N_43541,N_42351,N_41912);
or U43542 (N_43542,N_40347,N_41100);
nand U43543 (N_43543,N_41900,N_41585);
nor U43544 (N_43544,N_41924,N_41119);
nand U43545 (N_43545,N_42033,N_41990);
or U43546 (N_43546,N_42255,N_42323);
nor U43547 (N_43547,N_40353,N_40295);
or U43548 (N_43548,N_40917,N_42155);
or U43549 (N_43549,N_41432,N_41139);
xnor U43550 (N_43550,N_42448,N_41332);
or U43551 (N_43551,N_41200,N_40723);
and U43552 (N_43552,N_42086,N_41402);
or U43553 (N_43553,N_40116,N_40129);
nor U43554 (N_43554,N_42458,N_42000);
xor U43555 (N_43555,N_41798,N_42091);
and U43556 (N_43556,N_41299,N_41249);
and U43557 (N_43557,N_42393,N_40609);
and U43558 (N_43558,N_40426,N_40588);
nor U43559 (N_43559,N_42388,N_42193);
or U43560 (N_43560,N_42404,N_41552);
nand U43561 (N_43561,N_41652,N_41186);
nand U43562 (N_43562,N_42387,N_40068);
or U43563 (N_43563,N_42406,N_41104);
or U43564 (N_43564,N_40910,N_40633);
xnor U43565 (N_43565,N_40924,N_41035);
and U43566 (N_43566,N_41731,N_41818);
nor U43567 (N_43567,N_42249,N_41661);
and U43568 (N_43568,N_40725,N_42183);
nand U43569 (N_43569,N_41228,N_40185);
nor U43570 (N_43570,N_42034,N_41438);
and U43571 (N_43571,N_40884,N_41851);
or U43572 (N_43572,N_40072,N_40677);
or U43573 (N_43573,N_41849,N_41968);
or U43574 (N_43574,N_40865,N_42319);
or U43575 (N_43575,N_41458,N_41400);
and U43576 (N_43576,N_41384,N_40430);
xnor U43577 (N_43577,N_41743,N_40838);
nand U43578 (N_43578,N_40989,N_40282);
or U43579 (N_43579,N_41659,N_40573);
and U43580 (N_43580,N_41646,N_41057);
or U43581 (N_43581,N_40799,N_41712);
or U43582 (N_43582,N_41244,N_41512);
and U43583 (N_43583,N_41647,N_41706);
nand U43584 (N_43584,N_42238,N_41957);
xor U43585 (N_43585,N_42272,N_41601);
xor U43586 (N_43586,N_40754,N_40703);
nor U43587 (N_43587,N_41637,N_41133);
nand U43588 (N_43588,N_40372,N_41826);
and U43589 (N_43589,N_41667,N_40990);
or U43590 (N_43590,N_41120,N_40939);
and U43591 (N_43591,N_40385,N_40761);
nand U43592 (N_43592,N_40098,N_40548);
and U43593 (N_43593,N_40160,N_41928);
xnor U43594 (N_43594,N_42473,N_41983);
xor U43595 (N_43595,N_41583,N_41217);
and U43596 (N_43596,N_40087,N_40136);
nand U43597 (N_43597,N_40781,N_41679);
nor U43598 (N_43598,N_40896,N_41632);
or U43599 (N_43599,N_40613,N_41278);
xor U43600 (N_43600,N_40889,N_41609);
and U43601 (N_43601,N_40246,N_40720);
xnor U43602 (N_43602,N_41529,N_40726);
nor U43603 (N_43603,N_41033,N_41697);
nor U43604 (N_43604,N_42355,N_41289);
or U43605 (N_43605,N_40226,N_40536);
nor U43606 (N_43606,N_41105,N_42038);
or U43607 (N_43607,N_41605,N_42440);
xnor U43608 (N_43608,N_41331,N_40982);
nor U43609 (N_43609,N_40634,N_41624);
or U43610 (N_43610,N_41074,N_42350);
or U43611 (N_43611,N_42499,N_42369);
and U43612 (N_43612,N_41263,N_41283);
xnor U43613 (N_43613,N_41225,N_40562);
xnor U43614 (N_43614,N_40266,N_41897);
nand U43615 (N_43615,N_41008,N_41426);
nand U43616 (N_43616,N_42420,N_40335);
and U43617 (N_43617,N_40682,N_41296);
nand U43618 (N_43618,N_40030,N_40648);
nor U43619 (N_43619,N_41288,N_41674);
and U43620 (N_43620,N_40032,N_40487);
and U43621 (N_43621,N_41274,N_40287);
and U43622 (N_43622,N_42173,N_42257);
nand U43623 (N_43623,N_40288,N_42486);
nor U43624 (N_43624,N_41418,N_40181);
and U43625 (N_43625,N_41193,N_40444);
nor U43626 (N_43626,N_40590,N_40931);
nand U43627 (N_43627,N_40331,N_42205);
xor U43628 (N_43628,N_40269,N_40191);
and U43629 (N_43629,N_41234,N_41941);
nor U43630 (N_43630,N_41998,N_41981);
xnor U43631 (N_43631,N_40958,N_40902);
nand U43632 (N_43632,N_40738,N_40932);
xnor U43633 (N_43633,N_40735,N_41413);
or U43634 (N_43634,N_42395,N_41108);
xor U43635 (N_43635,N_40810,N_41763);
and U43636 (N_43636,N_40547,N_41779);
nand U43637 (N_43637,N_40897,N_41213);
xnor U43638 (N_43638,N_40564,N_40730);
and U43639 (N_43639,N_42363,N_41958);
and U43640 (N_43640,N_40581,N_42457);
xor U43641 (N_43641,N_41788,N_42243);
xnor U43642 (N_43642,N_41947,N_41447);
xor U43643 (N_43643,N_41865,N_42208);
nor U43644 (N_43644,N_40249,N_41444);
and U43645 (N_43645,N_40396,N_40480);
xor U43646 (N_43646,N_42453,N_41733);
and U43647 (N_43647,N_41794,N_42315);
nand U43648 (N_43648,N_40368,N_41666);
nand U43649 (N_43649,N_42455,N_42359);
xnor U43650 (N_43650,N_41836,N_42153);
or U43651 (N_43651,N_40167,N_40195);
nand U43652 (N_43652,N_40859,N_41902);
xnor U43653 (N_43653,N_41410,N_41305);
xor U43654 (N_43654,N_41623,N_41103);
or U43655 (N_43655,N_41820,N_42225);
nor U43656 (N_43656,N_41805,N_40179);
and U43657 (N_43657,N_41867,N_41741);
nand U43658 (N_43658,N_40304,N_40328);
xor U43659 (N_43659,N_41525,N_40427);
or U43660 (N_43660,N_41013,N_42413);
xnor U43661 (N_43661,N_40930,N_40198);
nand U43662 (N_43662,N_41002,N_40898);
xor U43663 (N_43663,N_41236,N_40920);
or U43664 (N_43664,N_40315,N_41911);
and U43665 (N_43665,N_42236,N_42171);
and U43666 (N_43666,N_40566,N_40458);
nor U43667 (N_43667,N_41229,N_41062);
and U43668 (N_43668,N_41714,N_41545);
or U43669 (N_43669,N_40145,N_41518);
or U43670 (N_43670,N_40134,N_41909);
xor U43671 (N_43671,N_40560,N_40872);
nor U43672 (N_43672,N_41726,N_41857);
or U43673 (N_43673,N_42409,N_41560);
nor U43674 (N_43674,N_42084,N_41404);
and U43675 (N_43675,N_41434,N_42074);
nand U43676 (N_43676,N_40326,N_42444);
and U43677 (N_43677,N_42335,N_40721);
nor U43678 (N_43678,N_40586,N_41494);
xor U43679 (N_43679,N_40011,N_40839);
and U43680 (N_43680,N_40391,N_41723);
and U43681 (N_43681,N_42373,N_40325);
nor U43682 (N_43682,N_40466,N_42275);
nor U43683 (N_43683,N_40766,N_40789);
and U43684 (N_43684,N_41142,N_40440);
or U43685 (N_43685,N_41179,N_41898);
and U43686 (N_43686,N_40381,N_40777);
and U43687 (N_43687,N_42248,N_41266);
or U43688 (N_43688,N_40268,N_40184);
and U43689 (N_43689,N_40125,N_40399);
nand U43690 (N_43690,N_41787,N_42148);
and U43691 (N_43691,N_41978,N_41934);
xnor U43692 (N_43692,N_41428,N_41477);
or U43693 (N_43693,N_40319,N_42221);
and U43694 (N_43694,N_41223,N_41774);
xnor U43695 (N_43695,N_41440,N_42217);
xnor U43696 (N_43696,N_42466,N_41782);
nand U43697 (N_43697,N_42411,N_40927);
or U43698 (N_43698,N_40460,N_41454);
nand U43699 (N_43699,N_41665,N_41387);
nand U43700 (N_43700,N_42200,N_40499);
xor U43701 (N_43701,N_41810,N_41579);
xor U43702 (N_43702,N_40117,N_41888);
xnor U43703 (N_43703,N_40955,N_40252);
nand U43704 (N_43704,N_41435,N_41285);
or U43705 (N_43705,N_41194,N_41050);
nand U43706 (N_43706,N_41955,N_41681);
and U43707 (N_43707,N_40357,N_42134);
nand U43708 (N_43708,N_41745,N_40061);
nor U43709 (N_43709,N_40405,N_40251);
nand U43710 (N_43710,N_41259,N_41856);
or U43711 (N_43711,N_40270,N_40707);
nand U43712 (N_43712,N_40120,N_40451);
nand U43713 (N_43713,N_42055,N_41759);
or U43714 (N_43714,N_41446,N_40159);
and U43715 (N_43715,N_40169,N_41367);
xnor U43716 (N_43716,N_41124,N_40306);
nor U43717 (N_43717,N_41027,N_40631);
nor U43718 (N_43718,N_42277,N_40423);
or U43719 (N_43719,N_41452,N_40713);
xnor U43720 (N_43720,N_41675,N_40532);
nor U43721 (N_43721,N_42271,N_40776);
and U43722 (N_43722,N_42118,N_40040);
and U43723 (N_43723,N_41598,N_40457);
nor U43724 (N_43724,N_40727,N_41324);
and U43725 (N_43725,N_42003,N_41321);
or U43726 (N_43726,N_42342,N_41521);
and U43727 (N_43727,N_41576,N_41398);
or U43728 (N_43728,N_42113,N_41721);
xnor U43729 (N_43729,N_40681,N_40772);
nand U43730 (N_43730,N_41464,N_41006);
nor U43731 (N_43731,N_41808,N_41060);
nand U43732 (N_43732,N_40204,N_41149);
xnor U43733 (N_43733,N_40127,N_41425);
or U43734 (N_43734,N_41833,N_40447);
nor U43735 (N_43735,N_41455,N_40299);
and U43736 (N_43736,N_40690,N_40033);
or U43737 (N_43737,N_40110,N_42128);
and U43738 (N_43738,N_40513,N_40334);
and U43739 (N_43739,N_42374,N_40858);
or U43740 (N_43740,N_40114,N_42408);
xnor U43741 (N_43741,N_41724,N_42220);
nand U43742 (N_43742,N_40031,N_41207);
and U43743 (N_43743,N_42316,N_40205);
xnor U43744 (N_43744,N_41388,N_40324);
nor U43745 (N_43745,N_42313,N_41603);
xnor U43746 (N_43746,N_40997,N_40193);
or U43747 (N_43747,N_41580,N_41765);
xor U43748 (N_43748,N_41786,N_40623);
nand U43749 (N_43749,N_40417,N_41405);
nor U43750 (N_43750,N_40303,N_40851);
and U43751 (N_43751,N_40118,N_40494);
or U43752 (N_43752,N_41566,N_40373);
and U43753 (N_43753,N_42381,N_40077);
xor U43754 (N_43754,N_41075,N_42282);
nor U43755 (N_43755,N_41790,N_40445);
nor U43756 (N_43756,N_40819,N_42350);
and U43757 (N_43757,N_42144,N_42384);
xor U43758 (N_43758,N_41391,N_41022);
nand U43759 (N_43759,N_42390,N_40268);
xnor U43760 (N_43760,N_40788,N_40154);
or U43761 (N_43761,N_41191,N_40812);
and U43762 (N_43762,N_42079,N_41441);
and U43763 (N_43763,N_42066,N_42434);
and U43764 (N_43764,N_42175,N_40595);
and U43765 (N_43765,N_42120,N_40349);
nor U43766 (N_43766,N_41807,N_42039);
or U43767 (N_43767,N_42445,N_40981);
and U43768 (N_43768,N_42026,N_41986);
xor U43769 (N_43769,N_42100,N_40171);
and U43770 (N_43770,N_41147,N_41493);
nand U43771 (N_43771,N_40900,N_40305);
nand U43772 (N_43772,N_40290,N_42149);
xnor U43773 (N_43773,N_40130,N_42311);
and U43774 (N_43774,N_42002,N_40794);
nor U43775 (N_43775,N_41787,N_40000);
and U43776 (N_43776,N_41292,N_41017);
and U43777 (N_43777,N_42357,N_40857);
xor U43778 (N_43778,N_41057,N_40010);
and U43779 (N_43779,N_40398,N_42300);
nand U43780 (N_43780,N_40974,N_41481);
nand U43781 (N_43781,N_40165,N_42234);
nor U43782 (N_43782,N_40936,N_40552);
nand U43783 (N_43783,N_41917,N_40171);
nor U43784 (N_43784,N_40310,N_42222);
nor U43785 (N_43785,N_40926,N_41920);
nand U43786 (N_43786,N_40883,N_41605);
nand U43787 (N_43787,N_40057,N_40853);
nor U43788 (N_43788,N_42481,N_40196);
nand U43789 (N_43789,N_41173,N_40655);
and U43790 (N_43790,N_42342,N_40609);
xor U43791 (N_43791,N_41279,N_41717);
or U43792 (N_43792,N_41312,N_40668);
or U43793 (N_43793,N_40039,N_42237);
nor U43794 (N_43794,N_40798,N_40444);
xor U43795 (N_43795,N_41578,N_41992);
nand U43796 (N_43796,N_41150,N_40490);
nor U43797 (N_43797,N_42226,N_42340);
nand U43798 (N_43798,N_41595,N_41687);
nor U43799 (N_43799,N_40671,N_41822);
nor U43800 (N_43800,N_41337,N_40747);
nand U43801 (N_43801,N_41184,N_40679);
and U43802 (N_43802,N_40639,N_42278);
xor U43803 (N_43803,N_41207,N_41800);
or U43804 (N_43804,N_41583,N_40289);
nand U43805 (N_43805,N_42486,N_40225);
xnor U43806 (N_43806,N_41924,N_41348);
and U43807 (N_43807,N_41504,N_41026);
or U43808 (N_43808,N_40610,N_40968);
xor U43809 (N_43809,N_41537,N_40279);
or U43810 (N_43810,N_40238,N_40258);
or U43811 (N_43811,N_41769,N_41012);
nor U43812 (N_43812,N_41286,N_41122);
xor U43813 (N_43813,N_40611,N_41038);
nor U43814 (N_43814,N_41727,N_40590);
nor U43815 (N_43815,N_40800,N_42388);
and U43816 (N_43816,N_40344,N_40340);
nor U43817 (N_43817,N_41723,N_42101);
nor U43818 (N_43818,N_40045,N_40116);
and U43819 (N_43819,N_41608,N_40420);
nand U43820 (N_43820,N_41325,N_40856);
nor U43821 (N_43821,N_40734,N_42107);
or U43822 (N_43822,N_40676,N_40431);
and U43823 (N_43823,N_41209,N_40161);
and U43824 (N_43824,N_42004,N_41606);
or U43825 (N_43825,N_40111,N_41511);
nor U43826 (N_43826,N_41856,N_40520);
nor U43827 (N_43827,N_40556,N_41589);
and U43828 (N_43828,N_40488,N_41272);
nand U43829 (N_43829,N_41611,N_40323);
and U43830 (N_43830,N_40223,N_41593);
and U43831 (N_43831,N_40380,N_40026);
xor U43832 (N_43832,N_41288,N_41453);
nand U43833 (N_43833,N_40554,N_42494);
and U43834 (N_43834,N_42069,N_42206);
nor U43835 (N_43835,N_41688,N_41644);
nor U43836 (N_43836,N_41779,N_40066);
nand U43837 (N_43837,N_41699,N_41666);
xnor U43838 (N_43838,N_40563,N_41428);
and U43839 (N_43839,N_40823,N_41797);
nand U43840 (N_43840,N_40690,N_42093);
nor U43841 (N_43841,N_40241,N_41880);
xnor U43842 (N_43842,N_41253,N_41251);
or U43843 (N_43843,N_40595,N_40724);
nor U43844 (N_43844,N_41986,N_42448);
xnor U43845 (N_43845,N_40055,N_42143);
nand U43846 (N_43846,N_42316,N_40660);
xor U43847 (N_43847,N_42084,N_41367);
and U43848 (N_43848,N_41620,N_40082);
nand U43849 (N_43849,N_40300,N_41342);
or U43850 (N_43850,N_40576,N_41496);
xor U43851 (N_43851,N_40695,N_41898);
and U43852 (N_43852,N_42116,N_42020);
or U43853 (N_43853,N_40434,N_41571);
nor U43854 (N_43854,N_40210,N_40609);
nand U43855 (N_43855,N_40993,N_41560);
or U43856 (N_43856,N_40282,N_40421);
xor U43857 (N_43857,N_40673,N_41812);
and U43858 (N_43858,N_42166,N_41606);
and U43859 (N_43859,N_41929,N_40475);
or U43860 (N_43860,N_41394,N_41461);
and U43861 (N_43861,N_40032,N_40602);
nand U43862 (N_43862,N_40228,N_40182);
nor U43863 (N_43863,N_42039,N_42069);
or U43864 (N_43864,N_41068,N_41486);
nand U43865 (N_43865,N_40630,N_41253);
or U43866 (N_43866,N_40862,N_40772);
nand U43867 (N_43867,N_41376,N_40020);
xor U43868 (N_43868,N_42057,N_41359);
or U43869 (N_43869,N_40550,N_40103);
and U43870 (N_43870,N_41577,N_41323);
nand U43871 (N_43871,N_42227,N_40783);
nor U43872 (N_43872,N_41142,N_42196);
or U43873 (N_43873,N_40661,N_41948);
and U43874 (N_43874,N_41636,N_42253);
and U43875 (N_43875,N_41519,N_41285);
nand U43876 (N_43876,N_41373,N_40758);
or U43877 (N_43877,N_40073,N_40462);
xnor U43878 (N_43878,N_41924,N_41260);
xor U43879 (N_43879,N_40606,N_40459);
and U43880 (N_43880,N_41352,N_41236);
and U43881 (N_43881,N_41732,N_40229);
or U43882 (N_43882,N_40630,N_40113);
and U43883 (N_43883,N_41597,N_41231);
and U43884 (N_43884,N_40590,N_42490);
and U43885 (N_43885,N_40634,N_42452);
or U43886 (N_43886,N_41459,N_41763);
or U43887 (N_43887,N_42040,N_42067);
or U43888 (N_43888,N_41400,N_41896);
and U43889 (N_43889,N_40076,N_41843);
and U43890 (N_43890,N_40524,N_40938);
nor U43891 (N_43891,N_41316,N_40476);
or U43892 (N_43892,N_40320,N_41667);
nand U43893 (N_43893,N_40174,N_42277);
or U43894 (N_43894,N_40161,N_40397);
or U43895 (N_43895,N_40538,N_40488);
xnor U43896 (N_43896,N_40396,N_42075);
nor U43897 (N_43897,N_40985,N_41343);
nor U43898 (N_43898,N_42343,N_41543);
or U43899 (N_43899,N_41768,N_41032);
or U43900 (N_43900,N_42321,N_42242);
nor U43901 (N_43901,N_40355,N_42074);
or U43902 (N_43902,N_41230,N_41951);
xnor U43903 (N_43903,N_40713,N_41609);
and U43904 (N_43904,N_41014,N_40651);
xnor U43905 (N_43905,N_41341,N_40610);
and U43906 (N_43906,N_42464,N_41793);
and U43907 (N_43907,N_41205,N_41648);
nand U43908 (N_43908,N_41617,N_41024);
nor U43909 (N_43909,N_40568,N_42055);
and U43910 (N_43910,N_41296,N_40191);
or U43911 (N_43911,N_42399,N_40703);
and U43912 (N_43912,N_40373,N_41408);
and U43913 (N_43913,N_42429,N_41341);
xor U43914 (N_43914,N_41306,N_41392);
or U43915 (N_43915,N_42084,N_41197);
and U43916 (N_43916,N_40918,N_40390);
xor U43917 (N_43917,N_41084,N_42049);
or U43918 (N_43918,N_42289,N_41651);
xnor U43919 (N_43919,N_41527,N_41112);
and U43920 (N_43920,N_42018,N_40528);
nor U43921 (N_43921,N_42272,N_41827);
nor U43922 (N_43922,N_41488,N_42189);
or U43923 (N_43923,N_40302,N_40482);
nand U43924 (N_43924,N_40558,N_40001);
and U43925 (N_43925,N_42031,N_40353);
and U43926 (N_43926,N_40993,N_40180);
nor U43927 (N_43927,N_42150,N_40752);
nand U43928 (N_43928,N_41877,N_40131);
nand U43929 (N_43929,N_40915,N_42127);
nand U43930 (N_43930,N_40911,N_41314);
xor U43931 (N_43931,N_41407,N_41870);
xnor U43932 (N_43932,N_41273,N_41440);
nand U43933 (N_43933,N_41899,N_42290);
nor U43934 (N_43934,N_40699,N_42391);
nor U43935 (N_43935,N_41603,N_41463);
nand U43936 (N_43936,N_41463,N_40779);
nor U43937 (N_43937,N_42430,N_41260);
and U43938 (N_43938,N_40241,N_41886);
nand U43939 (N_43939,N_41073,N_40143);
nand U43940 (N_43940,N_40745,N_42017);
nor U43941 (N_43941,N_42093,N_41682);
nor U43942 (N_43942,N_40147,N_42309);
xnor U43943 (N_43943,N_42153,N_42494);
and U43944 (N_43944,N_40718,N_41655);
nand U43945 (N_43945,N_41908,N_42230);
and U43946 (N_43946,N_40073,N_40875);
xnor U43947 (N_43947,N_40202,N_40555);
and U43948 (N_43948,N_41179,N_41902);
nor U43949 (N_43949,N_41083,N_41898);
nand U43950 (N_43950,N_42224,N_41665);
xnor U43951 (N_43951,N_40702,N_40941);
nand U43952 (N_43952,N_41013,N_42197);
nor U43953 (N_43953,N_40159,N_41596);
and U43954 (N_43954,N_41639,N_41314);
or U43955 (N_43955,N_40286,N_41400);
and U43956 (N_43956,N_40710,N_40622);
or U43957 (N_43957,N_41455,N_42230);
or U43958 (N_43958,N_41243,N_40268);
nor U43959 (N_43959,N_40029,N_40675);
nor U43960 (N_43960,N_40396,N_41972);
xor U43961 (N_43961,N_42474,N_40514);
xnor U43962 (N_43962,N_40849,N_41982);
or U43963 (N_43963,N_40744,N_40419);
nor U43964 (N_43964,N_40781,N_40534);
nand U43965 (N_43965,N_42407,N_41467);
nand U43966 (N_43966,N_41733,N_41926);
xnor U43967 (N_43967,N_42205,N_41977);
nor U43968 (N_43968,N_41344,N_42349);
xor U43969 (N_43969,N_41545,N_42480);
and U43970 (N_43970,N_42165,N_40219);
nand U43971 (N_43971,N_41086,N_41138);
nor U43972 (N_43972,N_41973,N_42469);
and U43973 (N_43973,N_40971,N_40808);
xor U43974 (N_43974,N_41817,N_42496);
xnor U43975 (N_43975,N_40629,N_42015);
and U43976 (N_43976,N_41099,N_41613);
and U43977 (N_43977,N_40635,N_42032);
nor U43978 (N_43978,N_40113,N_42249);
or U43979 (N_43979,N_41527,N_40828);
or U43980 (N_43980,N_40345,N_40866);
nor U43981 (N_43981,N_42139,N_41432);
xnor U43982 (N_43982,N_42366,N_42489);
or U43983 (N_43983,N_41377,N_41090);
xor U43984 (N_43984,N_41711,N_40412);
and U43985 (N_43985,N_40777,N_40206);
and U43986 (N_43986,N_40039,N_41497);
or U43987 (N_43987,N_40425,N_41403);
and U43988 (N_43988,N_41938,N_42323);
xnor U43989 (N_43989,N_41024,N_42301);
nand U43990 (N_43990,N_40028,N_42336);
nand U43991 (N_43991,N_40455,N_42432);
nand U43992 (N_43992,N_40158,N_41997);
nor U43993 (N_43993,N_41414,N_42167);
or U43994 (N_43994,N_41144,N_41329);
and U43995 (N_43995,N_41798,N_42491);
or U43996 (N_43996,N_41131,N_42301);
nand U43997 (N_43997,N_41564,N_40722);
or U43998 (N_43998,N_40779,N_40490);
nand U43999 (N_43999,N_41201,N_41613);
xor U44000 (N_44000,N_40565,N_41558);
and U44001 (N_44001,N_40218,N_40930);
xnor U44002 (N_44002,N_41220,N_41573);
xnor U44003 (N_44003,N_40104,N_42025);
or U44004 (N_44004,N_40114,N_42136);
and U44005 (N_44005,N_41008,N_41039);
xor U44006 (N_44006,N_40988,N_40307);
xnor U44007 (N_44007,N_41567,N_41559);
nor U44008 (N_44008,N_40937,N_41983);
xnor U44009 (N_44009,N_42207,N_41405);
nand U44010 (N_44010,N_40354,N_41324);
nand U44011 (N_44011,N_42488,N_40428);
nand U44012 (N_44012,N_41087,N_40362);
or U44013 (N_44013,N_41521,N_41270);
nor U44014 (N_44014,N_42146,N_40908);
nand U44015 (N_44015,N_40778,N_41224);
or U44016 (N_44016,N_41718,N_40980);
and U44017 (N_44017,N_41486,N_42045);
xnor U44018 (N_44018,N_41340,N_40632);
or U44019 (N_44019,N_40296,N_40544);
or U44020 (N_44020,N_40775,N_40409);
and U44021 (N_44021,N_40470,N_40572);
or U44022 (N_44022,N_41184,N_40499);
or U44023 (N_44023,N_40061,N_41304);
or U44024 (N_44024,N_40415,N_41844);
nand U44025 (N_44025,N_40428,N_40510);
or U44026 (N_44026,N_41788,N_41503);
xnor U44027 (N_44027,N_40273,N_42409);
and U44028 (N_44028,N_41535,N_42429);
or U44029 (N_44029,N_42045,N_40456);
nor U44030 (N_44030,N_42122,N_41036);
xor U44031 (N_44031,N_40440,N_42250);
nor U44032 (N_44032,N_41388,N_40310);
nor U44033 (N_44033,N_40995,N_41327);
xnor U44034 (N_44034,N_41354,N_40352);
nand U44035 (N_44035,N_41969,N_41049);
or U44036 (N_44036,N_42310,N_41694);
and U44037 (N_44037,N_41195,N_42237);
xor U44038 (N_44038,N_41574,N_41356);
or U44039 (N_44039,N_40037,N_40940);
and U44040 (N_44040,N_40230,N_41895);
and U44041 (N_44041,N_41496,N_41115);
xnor U44042 (N_44042,N_40830,N_40638);
xnor U44043 (N_44043,N_41011,N_40170);
xnor U44044 (N_44044,N_42474,N_40195);
or U44045 (N_44045,N_41194,N_40517);
nor U44046 (N_44046,N_41086,N_42407);
nand U44047 (N_44047,N_40571,N_41780);
nor U44048 (N_44048,N_41096,N_42310);
nand U44049 (N_44049,N_42460,N_41506);
xnor U44050 (N_44050,N_41159,N_41139);
nor U44051 (N_44051,N_40891,N_42294);
nor U44052 (N_44052,N_41104,N_41851);
or U44053 (N_44053,N_42185,N_42122);
nand U44054 (N_44054,N_42306,N_42069);
and U44055 (N_44055,N_41449,N_41847);
and U44056 (N_44056,N_40172,N_41226);
xnor U44057 (N_44057,N_41330,N_40769);
nand U44058 (N_44058,N_41151,N_40929);
nor U44059 (N_44059,N_40483,N_41539);
xnor U44060 (N_44060,N_40673,N_40040);
nand U44061 (N_44061,N_40598,N_41249);
nor U44062 (N_44062,N_40229,N_41006);
xor U44063 (N_44063,N_40019,N_42232);
nand U44064 (N_44064,N_41189,N_41866);
nor U44065 (N_44065,N_40385,N_40842);
and U44066 (N_44066,N_40312,N_42003);
and U44067 (N_44067,N_40858,N_41417);
nand U44068 (N_44068,N_42244,N_40277);
or U44069 (N_44069,N_40035,N_41511);
and U44070 (N_44070,N_40868,N_41151);
nand U44071 (N_44071,N_40538,N_40959);
and U44072 (N_44072,N_40769,N_41351);
xnor U44073 (N_44073,N_40255,N_40825);
or U44074 (N_44074,N_41122,N_41959);
nor U44075 (N_44075,N_40224,N_42036);
nand U44076 (N_44076,N_42266,N_40475);
and U44077 (N_44077,N_40845,N_40701);
and U44078 (N_44078,N_40929,N_41381);
and U44079 (N_44079,N_40899,N_41231);
nand U44080 (N_44080,N_40472,N_40088);
nor U44081 (N_44081,N_42192,N_40686);
nor U44082 (N_44082,N_42055,N_40351);
nor U44083 (N_44083,N_42223,N_42486);
nand U44084 (N_44084,N_40691,N_42499);
nor U44085 (N_44085,N_40366,N_41229);
or U44086 (N_44086,N_42161,N_41593);
nor U44087 (N_44087,N_42490,N_40470);
nand U44088 (N_44088,N_41747,N_40985);
xor U44089 (N_44089,N_42310,N_40332);
nand U44090 (N_44090,N_40190,N_42154);
nor U44091 (N_44091,N_41896,N_40434);
or U44092 (N_44092,N_41295,N_42246);
and U44093 (N_44093,N_40727,N_40805);
nor U44094 (N_44094,N_40574,N_41701);
or U44095 (N_44095,N_42413,N_41851);
or U44096 (N_44096,N_40905,N_40184);
or U44097 (N_44097,N_41283,N_41511);
xor U44098 (N_44098,N_41559,N_42411);
nand U44099 (N_44099,N_41097,N_42122);
or U44100 (N_44100,N_41405,N_42465);
or U44101 (N_44101,N_41358,N_40228);
and U44102 (N_44102,N_42245,N_41740);
or U44103 (N_44103,N_40426,N_41109);
nor U44104 (N_44104,N_40372,N_40843);
nor U44105 (N_44105,N_41402,N_41815);
xor U44106 (N_44106,N_41176,N_41325);
nor U44107 (N_44107,N_41370,N_42263);
nand U44108 (N_44108,N_40094,N_41170);
nor U44109 (N_44109,N_41732,N_41800);
nand U44110 (N_44110,N_40756,N_40677);
and U44111 (N_44111,N_41193,N_42252);
or U44112 (N_44112,N_40957,N_41224);
nor U44113 (N_44113,N_40951,N_41220);
nand U44114 (N_44114,N_40650,N_42067);
nor U44115 (N_44115,N_40078,N_41661);
nor U44116 (N_44116,N_41340,N_42029);
xor U44117 (N_44117,N_41780,N_40825);
or U44118 (N_44118,N_42426,N_40327);
nand U44119 (N_44119,N_40953,N_40213);
and U44120 (N_44120,N_41999,N_41866);
xor U44121 (N_44121,N_40817,N_40842);
nand U44122 (N_44122,N_41449,N_40805);
xnor U44123 (N_44123,N_40963,N_41235);
xor U44124 (N_44124,N_40634,N_41115);
nand U44125 (N_44125,N_41221,N_40550);
and U44126 (N_44126,N_41172,N_40146);
xnor U44127 (N_44127,N_41147,N_41132);
nor U44128 (N_44128,N_42137,N_42272);
nor U44129 (N_44129,N_41092,N_41554);
xor U44130 (N_44130,N_40097,N_41595);
or U44131 (N_44131,N_41518,N_40028);
nand U44132 (N_44132,N_40815,N_40011);
nor U44133 (N_44133,N_40014,N_41412);
or U44134 (N_44134,N_41933,N_42098);
nor U44135 (N_44135,N_42275,N_40991);
or U44136 (N_44136,N_40187,N_40680);
nand U44137 (N_44137,N_40468,N_41414);
nand U44138 (N_44138,N_42079,N_40309);
nand U44139 (N_44139,N_40725,N_40754);
nand U44140 (N_44140,N_40911,N_40754);
or U44141 (N_44141,N_41555,N_40857);
or U44142 (N_44142,N_40504,N_41529);
nor U44143 (N_44143,N_42048,N_41115);
nor U44144 (N_44144,N_42358,N_41282);
xor U44145 (N_44145,N_41395,N_40215);
nand U44146 (N_44146,N_40697,N_40680);
xnor U44147 (N_44147,N_40227,N_40153);
or U44148 (N_44148,N_41098,N_41119);
xor U44149 (N_44149,N_41618,N_41365);
and U44150 (N_44150,N_41000,N_40498);
and U44151 (N_44151,N_40787,N_41135);
xor U44152 (N_44152,N_41069,N_40591);
or U44153 (N_44153,N_41903,N_41063);
nand U44154 (N_44154,N_40446,N_41474);
or U44155 (N_44155,N_40850,N_40050);
or U44156 (N_44156,N_41968,N_42135);
nor U44157 (N_44157,N_42393,N_41981);
xnor U44158 (N_44158,N_40325,N_41299);
or U44159 (N_44159,N_41705,N_40013);
and U44160 (N_44160,N_40280,N_41197);
and U44161 (N_44161,N_40458,N_40872);
nand U44162 (N_44162,N_40096,N_40972);
nand U44163 (N_44163,N_40363,N_40973);
xor U44164 (N_44164,N_42385,N_42243);
nor U44165 (N_44165,N_42013,N_40960);
nand U44166 (N_44166,N_40675,N_42169);
xnor U44167 (N_44167,N_42443,N_42324);
or U44168 (N_44168,N_42489,N_40037);
nor U44169 (N_44169,N_41889,N_42318);
xor U44170 (N_44170,N_41180,N_41702);
nor U44171 (N_44171,N_42219,N_41651);
and U44172 (N_44172,N_40472,N_42341);
or U44173 (N_44173,N_40407,N_42461);
or U44174 (N_44174,N_42318,N_41128);
and U44175 (N_44175,N_41518,N_41226);
nor U44176 (N_44176,N_40691,N_40166);
and U44177 (N_44177,N_41574,N_40598);
or U44178 (N_44178,N_40598,N_40692);
nand U44179 (N_44179,N_40853,N_41989);
nand U44180 (N_44180,N_40237,N_42127);
or U44181 (N_44181,N_40492,N_41947);
nand U44182 (N_44182,N_40386,N_40450);
nor U44183 (N_44183,N_41153,N_41473);
or U44184 (N_44184,N_41112,N_42437);
nor U44185 (N_44185,N_40529,N_41726);
xor U44186 (N_44186,N_41053,N_41519);
and U44187 (N_44187,N_40802,N_41395);
xnor U44188 (N_44188,N_41734,N_40060);
nand U44189 (N_44189,N_41840,N_40558);
and U44190 (N_44190,N_40942,N_42330);
or U44191 (N_44191,N_41527,N_42213);
and U44192 (N_44192,N_41019,N_41908);
nand U44193 (N_44193,N_42102,N_41490);
xnor U44194 (N_44194,N_41243,N_40935);
or U44195 (N_44195,N_41564,N_40961);
xnor U44196 (N_44196,N_40797,N_41641);
or U44197 (N_44197,N_42480,N_41208);
or U44198 (N_44198,N_41670,N_42278);
nand U44199 (N_44199,N_40191,N_40711);
nor U44200 (N_44200,N_42496,N_40967);
xnor U44201 (N_44201,N_40400,N_40714);
xnor U44202 (N_44202,N_41741,N_41930);
xnor U44203 (N_44203,N_40331,N_41830);
xnor U44204 (N_44204,N_41625,N_41235);
nand U44205 (N_44205,N_40301,N_40235);
nand U44206 (N_44206,N_41461,N_40842);
nor U44207 (N_44207,N_40185,N_40120);
xnor U44208 (N_44208,N_41228,N_41143);
or U44209 (N_44209,N_41496,N_41329);
and U44210 (N_44210,N_41327,N_40456);
xor U44211 (N_44211,N_41802,N_40337);
or U44212 (N_44212,N_40084,N_40994);
or U44213 (N_44213,N_41447,N_40178);
xnor U44214 (N_44214,N_40589,N_40621);
nor U44215 (N_44215,N_42426,N_40860);
nand U44216 (N_44216,N_40556,N_40899);
xor U44217 (N_44217,N_42299,N_40797);
xor U44218 (N_44218,N_41056,N_41821);
nand U44219 (N_44219,N_42410,N_42185);
nand U44220 (N_44220,N_41258,N_41459);
xnor U44221 (N_44221,N_41441,N_41111);
nand U44222 (N_44222,N_42152,N_41510);
and U44223 (N_44223,N_42136,N_42494);
and U44224 (N_44224,N_42077,N_40887);
nor U44225 (N_44225,N_42350,N_40608);
nand U44226 (N_44226,N_41965,N_41696);
nor U44227 (N_44227,N_41789,N_42279);
or U44228 (N_44228,N_41928,N_40277);
nor U44229 (N_44229,N_40114,N_42220);
xnor U44230 (N_44230,N_41299,N_42125);
nand U44231 (N_44231,N_41696,N_41635);
xor U44232 (N_44232,N_40625,N_41473);
xor U44233 (N_44233,N_41021,N_40922);
and U44234 (N_44234,N_41155,N_42365);
nand U44235 (N_44235,N_41412,N_40929);
xnor U44236 (N_44236,N_40960,N_42292);
nor U44237 (N_44237,N_41579,N_40185);
nand U44238 (N_44238,N_42046,N_42300);
nor U44239 (N_44239,N_40920,N_41626);
and U44240 (N_44240,N_40727,N_41815);
xor U44241 (N_44241,N_40774,N_40801);
nand U44242 (N_44242,N_42371,N_41737);
nor U44243 (N_44243,N_42366,N_40448);
and U44244 (N_44244,N_40335,N_41989);
nor U44245 (N_44245,N_42111,N_41507);
nor U44246 (N_44246,N_41327,N_41457);
nor U44247 (N_44247,N_41097,N_40578);
nand U44248 (N_44248,N_41135,N_40231);
or U44249 (N_44249,N_41819,N_40957);
or U44250 (N_44250,N_40386,N_42386);
xor U44251 (N_44251,N_41292,N_41457);
nor U44252 (N_44252,N_41644,N_40294);
and U44253 (N_44253,N_41185,N_40129);
nand U44254 (N_44254,N_41148,N_40950);
or U44255 (N_44255,N_41251,N_42226);
and U44256 (N_44256,N_40381,N_42274);
nor U44257 (N_44257,N_40513,N_41812);
nor U44258 (N_44258,N_40415,N_40535);
nor U44259 (N_44259,N_41754,N_40368);
nor U44260 (N_44260,N_41447,N_41881);
nor U44261 (N_44261,N_40456,N_40606);
nand U44262 (N_44262,N_41331,N_40812);
or U44263 (N_44263,N_40735,N_42261);
or U44264 (N_44264,N_40120,N_41566);
nand U44265 (N_44265,N_41996,N_40529);
nor U44266 (N_44266,N_42230,N_41143);
and U44267 (N_44267,N_42039,N_41549);
nor U44268 (N_44268,N_40458,N_40923);
xor U44269 (N_44269,N_41031,N_41370);
or U44270 (N_44270,N_41624,N_41636);
nor U44271 (N_44271,N_41527,N_41870);
nor U44272 (N_44272,N_42224,N_40351);
and U44273 (N_44273,N_40428,N_41948);
xor U44274 (N_44274,N_41750,N_40291);
or U44275 (N_44275,N_40682,N_40739);
nand U44276 (N_44276,N_41602,N_41239);
nand U44277 (N_44277,N_41281,N_42255);
xnor U44278 (N_44278,N_41487,N_40420);
and U44279 (N_44279,N_42483,N_41029);
nand U44280 (N_44280,N_40211,N_41813);
and U44281 (N_44281,N_42210,N_40163);
nand U44282 (N_44282,N_40901,N_40921);
and U44283 (N_44283,N_40162,N_41719);
or U44284 (N_44284,N_41160,N_41895);
nor U44285 (N_44285,N_41565,N_42135);
nor U44286 (N_44286,N_40998,N_42081);
nor U44287 (N_44287,N_40119,N_41198);
and U44288 (N_44288,N_41547,N_40275);
xor U44289 (N_44289,N_41558,N_41471);
and U44290 (N_44290,N_41870,N_42428);
nor U44291 (N_44291,N_41357,N_40749);
or U44292 (N_44292,N_42052,N_42380);
xor U44293 (N_44293,N_41923,N_41975);
or U44294 (N_44294,N_41122,N_41577);
and U44295 (N_44295,N_40020,N_40478);
nand U44296 (N_44296,N_42268,N_41612);
nand U44297 (N_44297,N_41478,N_41614);
xnor U44298 (N_44298,N_42100,N_40882);
nand U44299 (N_44299,N_40928,N_41826);
xor U44300 (N_44300,N_41772,N_41432);
xor U44301 (N_44301,N_42125,N_40108);
nor U44302 (N_44302,N_41495,N_40335);
nand U44303 (N_44303,N_41609,N_40175);
xor U44304 (N_44304,N_42322,N_40251);
nor U44305 (N_44305,N_41761,N_41766);
xor U44306 (N_44306,N_40174,N_41716);
nor U44307 (N_44307,N_40146,N_42006);
nor U44308 (N_44308,N_40349,N_40850);
and U44309 (N_44309,N_40279,N_41653);
xor U44310 (N_44310,N_40106,N_41272);
and U44311 (N_44311,N_41583,N_42065);
xnor U44312 (N_44312,N_42096,N_42467);
xnor U44313 (N_44313,N_42369,N_42273);
nand U44314 (N_44314,N_42102,N_41497);
and U44315 (N_44315,N_41978,N_40490);
xor U44316 (N_44316,N_40171,N_41793);
nand U44317 (N_44317,N_41246,N_40495);
and U44318 (N_44318,N_40230,N_40555);
or U44319 (N_44319,N_40501,N_42409);
or U44320 (N_44320,N_41409,N_41153);
or U44321 (N_44321,N_40091,N_41349);
nor U44322 (N_44322,N_41893,N_40190);
or U44323 (N_44323,N_42086,N_41607);
nand U44324 (N_44324,N_41353,N_40103);
and U44325 (N_44325,N_42120,N_41876);
xor U44326 (N_44326,N_41543,N_41409);
or U44327 (N_44327,N_41623,N_41523);
and U44328 (N_44328,N_40469,N_40286);
and U44329 (N_44329,N_41978,N_40815);
xnor U44330 (N_44330,N_41581,N_40486);
nor U44331 (N_44331,N_41453,N_40281);
and U44332 (N_44332,N_41800,N_41199);
and U44333 (N_44333,N_42080,N_40585);
nand U44334 (N_44334,N_40683,N_41155);
or U44335 (N_44335,N_41268,N_41197);
nand U44336 (N_44336,N_40510,N_40721);
nor U44337 (N_44337,N_42139,N_40167);
nand U44338 (N_44338,N_40532,N_42485);
and U44339 (N_44339,N_40291,N_40587);
or U44340 (N_44340,N_42166,N_41954);
nand U44341 (N_44341,N_41844,N_42320);
nor U44342 (N_44342,N_41232,N_41043);
and U44343 (N_44343,N_41016,N_42297);
xor U44344 (N_44344,N_42152,N_40352);
nand U44345 (N_44345,N_41669,N_42035);
and U44346 (N_44346,N_41302,N_41020);
nand U44347 (N_44347,N_41038,N_41290);
nor U44348 (N_44348,N_41152,N_42110);
xnor U44349 (N_44349,N_40295,N_41297);
nor U44350 (N_44350,N_42396,N_40941);
nor U44351 (N_44351,N_41915,N_41395);
nand U44352 (N_44352,N_41962,N_42422);
nor U44353 (N_44353,N_40879,N_40429);
nor U44354 (N_44354,N_41335,N_40384);
or U44355 (N_44355,N_41610,N_42101);
nor U44356 (N_44356,N_40060,N_40848);
nand U44357 (N_44357,N_42134,N_42318);
nor U44358 (N_44358,N_42257,N_40962);
xor U44359 (N_44359,N_41798,N_40440);
nand U44360 (N_44360,N_40903,N_40531);
or U44361 (N_44361,N_41399,N_40684);
or U44362 (N_44362,N_40548,N_41275);
nor U44363 (N_44363,N_40767,N_41302);
and U44364 (N_44364,N_41958,N_40251);
nor U44365 (N_44365,N_40077,N_40776);
xor U44366 (N_44366,N_41166,N_40284);
xor U44367 (N_44367,N_41984,N_41772);
xnor U44368 (N_44368,N_41394,N_40688);
nor U44369 (N_44369,N_42140,N_41479);
or U44370 (N_44370,N_40785,N_40637);
and U44371 (N_44371,N_40770,N_41386);
and U44372 (N_44372,N_40627,N_40904);
or U44373 (N_44373,N_42153,N_40277);
or U44374 (N_44374,N_41931,N_40108);
nand U44375 (N_44375,N_40714,N_40841);
or U44376 (N_44376,N_42448,N_42353);
or U44377 (N_44377,N_40798,N_40078);
xnor U44378 (N_44378,N_41566,N_40501);
nand U44379 (N_44379,N_41255,N_40428);
nand U44380 (N_44380,N_41276,N_40521);
and U44381 (N_44381,N_40500,N_40318);
and U44382 (N_44382,N_41088,N_41268);
and U44383 (N_44383,N_40694,N_40431);
or U44384 (N_44384,N_40284,N_41620);
nand U44385 (N_44385,N_41501,N_40972);
or U44386 (N_44386,N_40845,N_40252);
nor U44387 (N_44387,N_42040,N_41990);
or U44388 (N_44388,N_42255,N_42413);
nor U44389 (N_44389,N_41494,N_40316);
or U44390 (N_44390,N_40583,N_40995);
or U44391 (N_44391,N_41828,N_40652);
xnor U44392 (N_44392,N_41034,N_41409);
nor U44393 (N_44393,N_41494,N_40671);
and U44394 (N_44394,N_41253,N_42464);
nand U44395 (N_44395,N_40653,N_40478);
and U44396 (N_44396,N_41934,N_41952);
xnor U44397 (N_44397,N_41445,N_41013);
nor U44398 (N_44398,N_41930,N_42195);
and U44399 (N_44399,N_41652,N_41866);
nor U44400 (N_44400,N_41081,N_40233);
nand U44401 (N_44401,N_40401,N_41907);
or U44402 (N_44402,N_40306,N_41372);
xor U44403 (N_44403,N_40321,N_40632);
nand U44404 (N_44404,N_42089,N_41892);
nor U44405 (N_44405,N_40086,N_40223);
and U44406 (N_44406,N_42021,N_42224);
nor U44407 (N_44407,N_41083,N_42299);
nand U44408 (N_44408,N_40339,N_40109);
or U44409 (N_44409,N_41456,N_42180);
nand U44410 (N_44410,N_40854,N_41810);
nor U44411 (N_44411,N_42113,N_42062);
and U44412 (N_44412,N_40382,N_40748);
nor U44413 (N_44413,N_41012,N_41823);
nand U44414 (N_44414,N_40028,N_40571);
or U44415 (N_44415,N_42011,N_41329);
xor U44416 (N_44416,N_41239,N_41377);
or U44417 (N_44417,N_41377,N_41747);
xor U44418 (N_44418,N_40528,N_40508);
and U44419 (N_44419,N_41416,N_41829);
nand U44420 (N_44420,N_40540,N_40325);
nor U44421 (N_44421,N_40744,N_40176);
and U44422 (N_44422,N_41011,N_41437);
and U44423 (N_44423,N_41883,N_42111);
xor U44424 (N_44424,N_40701,N_42033);
and U44425 (N_44425,N_41980,N_41530);
and U44426 (N_44426,N_41444,N_40376);
xor U44427 (N_44427,N_40565,N_41197);
or U44428 (N_44428,N_41313,N_42119);
nor U44429 (N_44429,N_42075,N_42480);
and U44430 (N_44430,N_40382,N_40017);
xnor U44431 (N_44431,N_40825,N_42092);
or U44432 (N_44432,N_42303,N_40917);
or U44433 (N_44433,N_40346,N_40967);
nor U44434 (N_44434,N_40086,N_41027);
nor U44435 (N_44435,N_41540,N_40112);
or U44436 (N_44436,N_40996,N_40107);
and U44437 (N_44437,N_40626,N_40235);
nand U44438 (N_44438,N_42425,N_41423);
and U44439 (N_44439,N_41543,N_40141);
xor U44440 (N_44440,N_41488,N_40092);
nand U44441 (N_44441,N_42086,N_40540);
or U44442 (N_44442,N_40379,N_41626);
xnor U44443 (N_44443,N_42111,N_40345);
or U44444 (N_44444,N_41842,N_41474);
or U44445 (N_44445,N_42061,N_40672);
and U44446 (N_44446,N_41750,N_40668);
xor U44447 (N_44447,N_41642,N_40287);
or U44448 (N_44448,N_41004,N_40969);
or U44449 (N_44449,N_40635,N_40533);
and U44450 (N_44450,N_40488,N_42003);
xor U44451 (N_44451,N_40732,N_42096);
and U44452 (N_44452,N_41231,N_41648);
and U44453 (N_44453,N_40877,N_41417);
nor U44454 (N_44454,N_40190,N_42397);
and U44455 (N_44455,N_40415,N_40283);
xnor U44456 (N_44456,N_40504,N_40693);
and U44457 (N_44457,N_42150,N_41570);
or U44458 (N_44458,N_41412,N_42003);
nor U44459 (N_44459,N_41723,N_41093);
nand U44460 (N_44460,N_40455,N_41713);
nand U44461 (N_44461,N_42298,N_40359);
nor U44462 (N_44462,N_40168,N_40486);
nor U44463 (N_44463,N_41138,N_41832);
xor U44464 (N_44464,N_41357,N_40702);
or U44465 (N_44465,N_41172,N_40281);
or U44466 (N_44466,N_42109,N_40036);
nor U44467 (N_44467,N_42018,N_41552);
and U44468 (N_44468,N_40043,N_40774);
nand U44469 (N_44469,N_41049,N_41960);
xor U44470 (N_44470,N_40944,N_40207);
or U44471 (N_44471,N_41639,N_42027);
or U44472 (N_44472,N_41695,N_42272);
and U44473 (N_44473,N_40284,N_40532);
and U44474 (N_44474,N_40492,N_41372);
nand U44475 (N_44475,N_40267,N_40428);
xnor U44476 (N_44476,N_41271,N_40043);
and U44477 (N_44477,N_41265,N_40796);
and U44478 (N_44478,N_40356,N_41631);
nand U44479 (N_44479,N_40546,N_40374);
and U44480 (N_44480,N_42069,N_41184);
nand U44481 (N_44481,N_40951,N_40939);
or U44482 (N_44482,N_42450,N_40258);
or U44483 (N_44483,N_42394,N_40612);
nor U44484 (N_44484,N_40817,N_40839);
nand U44485 (N_44485,N_41957,N_40776);
and U44486 (N_44486,N_41936,N_40024);
xor U44487 (N_44487,N_41090,N_41030);
nand U44488 (N_44488,N_42257,N_40505);
nand U44489 (N_44489,N_40820,N_41309);
and U44490 (N_44490,N_42473,N_40510);
and U44491 (N_44491,N_41314,N_40001);
or U44492 (N_44492,N_40899,N_41058);
xnor U44493 (N_44493,N_42484,N_41978);
nand U44494 (N_44494,N_41301,N_42205);
and U44495 (N_44495,N_41418,N_40817);
and U44496 (N_44496,N_41384,N_40938);
nand U44497 (N_44497,N_40847,N_40890);
nor U44498 (N_44498,N_40928,N_40171);
or U44499 (N_44499,N_41904,N_42086);
or U44500 (N_44500,N_41477,N_42453);
nand U44501 (N_44501,N_41891,N_41126);
or U44502 (N_44502,N_40338,N_41048);
and U44503 (N_44503,N_40213,N_40478);
and U44504 (N_44504,N_41585,N_41571);
nor U44505 (N_44505,N_41366,N_41806);
nor U44506 (N_44506,N_41517,N_40021);
xor U44507 (N_44507,N_41413,N_41000);
xnor U44508 (N_44508,N_40320,N_41039);
nand U44509 (N_44509,N_40909,N_40100);
and U44510 (N_44510,N_40996,N_40126);
or U44511 (N_44511,N_41781,N_41333);
or U44512 (N_44512,N_41347,N_40992);
nor U44513 (N_44513,N_41556,N_40420);
nor U44514 (N_44514,N_40763,N_41911);
or U44515 (N_44515,N_42396,N_41299);
xor U44516 (N_44516,N_41993,N_42461);
or U44517 (N_44517,N_42481,N_40456);
nand U44518 (N_44518,N_41309,N_41257);
nor U44519 (N_44519,N_41529,N_42253);
or U44520 (N_44520,N_41971,N_40666);
and U44521 (N_44521,N_42212,N_42293);
nor U44522 (N_44522,N_40609,N_40228);
or U44523 (N_44523,N_42470,N_41088);
xnor U44524 (N_44524,N_40951,N_41512);
xor U44525 (N_44525,N_40597,N_42371);
and U44526 (N_44526,N_42155,N_41424);
or U44527 (N_44527,N_40058,N_40239);
nor U44528 (N_44528,N_42330,N_41832);
nor U44529 (N_44529,N_42209,N_40454);
xnor U44530 (N_44530,N_40985,N_40124);
nand U44531 (N_44531,N_40952,N_40087);
nand U44532 (N_44532,N_40202,N_40698);
nand U44533 (N_44533,N_41912,N_40488);
and U44534 (N_44534,N_40375,N_41441);
nor U44535 (N_44535,N_41000,N_41633);
xnor U44536 (N_44536,N_41445,N_41341);
nor U44537 (N_44537,N_42346,N_40410);
or U44538 (N_44538,N_41116,N_41746);
xnor U44539 (N_44539,N_40043,N_42270);
nor U44540 (N_44540,N_42375,N_41850);
nor U44541 (N_44541,N_41365,N_41412);
xor U44542 (N_44542,N_41281,N_42072);
nand U44543 (N_44543,N_41256,N_41590);
xnor U44544 (N_44544,N_42459,N_40618);
nor U44545 (N_44545,N_41818,N_41235);
and U44546 (N_44546,N_40364,N_42059);
or U44547 (N_44547,N_40153,N_41095);
nand U44548 (N_44548,N_41290,N_41615);
or U44549 (N_44549,N_41624,N_41956);
xor U44550 (N_44550,N_40800,N_41306);
or U44551 (N_44551,N_42284,N_41695);
nand U44552 (N_44552,N_41459,N_42486);
and U44553 (N_44553,N_40793,N_42341);
nor U44554 (N_44554,N_42309,N_41005);
and U44555 (N_44555,N_41025,N_40689);
xor U44556 (N_44556,N_42112,N_40956);
nand U44557 (N_44557,N_41199,N_40145);
xor U44558 (N_44558,N_41048,N_40100);
nand U44559 (N_44559,N_41017,N_41606);
nand U44560 (N_44560,N_40405,N_41801);
nor U44561 (N_44561,N_41510,N_42017);
xnor U44562 (N_44562,N_40746,N_41246);
nand U44563 (N_44563,N_42110,N_41922);
and U44564 (N_44564,N_40126,N_40485);
xor U44565 (N_44565,N_40729,N_41670);
nand U44566 (N_44566,N_42231,N_42421);
or U44567 (N_44567,N_41877,N_40927);
xnor U44568 (N_44568,N_42321,N_41907);
or U44569 (N_44569,N_40909,N_40453);
or U44570 (N_44570,N_40875,N_41121);
and U44571 (N_44571,N_42358,N_41728);
nor U44572 (N_44572,N_41921,N_42446);
and U44573 (N_44573,N_40277,N_40635);
xor U44574 (N_44574,N_40276,N_42138);
nand U44575 (N_44575,N_40366,N_40053);
nor U44576 (N_44576,N_40708,N_41586);
nor U44577 (N_44577,N_40713,N_40573);
or U44578 (N_44578,N_42434,N_42298);
xor U44579 (N_44579,N_41012,N_41787);
or U44580 (N_44580,N_40914,N_41129);
xnor U44581 (N_44581,N_41782,N_40463);
xor U44582 (N_44582,N_41122,N_42275);
and U44583 (N_44583,N_41250,N_40150);
nand U44584 (N_44584,N_40785,N_40064);
and U44585 (N_44585,N_42286,N_41019);
xnor U44586 (N_44586,N_40373,N_41951);
nor U44587 (N_44587,N_42309,N_40174);
xnor U44588 (N_44588,N_42415,N_41789);
xor U44589 (N_44589,N_41097,N_41004);
xor U44590 (N_44590,N_40761,N_41029);
xor U44591 (N_44591,N_41636,N_40861);
xnor U44592 (N_44592,N_40660,N_42146);
and U44593 (N_44593,N_41932,N_41198);
and U44594 (N_44594,N_41337,N_41503);
xnor U44595 (N_44595,N_41184,N_41632);
xnor U44596 (N_44596,N_40336,N_42237);
or U44597 (N_44597,N_41287,N_41872);
or U44598 (N_44598,N_41989,N_40631);
nand U44599 (N_44599,N_41684,N_42026);
or U44600 (N_44600,N_41956,N_42096);
and U44601 (N_44601,N_40229,N_42424);
nor U44602 (N_44602,N_41074,N_41776);
and U44603 (N_44603,N_40231,N_42090);
or U44604 (N_44604,N_42216,N_41398);
nand U44605 (N_44605,N_41629,N_40688);
or U44606 (N_44606,N_41196,N_40758);
xnor U44607 (N_44607,N_40726,N_40737);
nand U44608 (N_44608,N_40395,N_41678);
nor U44609 (N_44609,N_41018,N_41934);
xor U44610 (N_44610,N_42407,N_41296);
xor U44611 (N_44611,N_40668,N_42360);
xnor U44612 (N_44612,N_42249,N_42119);
nor U44613 (N_44613,N_41605,N_41358);
nor U44614 (N_44614,N_41788,N_40912);
nor U44615 (N_44615,N_41899,N_40945);
nand U44616 (N_44616,N_41464,N_41387);
and U44617 (N_44617,N_42230,N_40128);
or U44618 (N_44618,N_40543,N_41274);
nor U44619 (N_44619,N_40957,N_41071);
or U44620 (N_44620,N_42439,N_41882);
and U44621 (N_44621,N_40526,N_41841);
xnor U44622 (N_44622,N_41820,N_41548);
and U44623 (N_44623,N_42222,N_41286);
xor U44624 (N_44624,N_41690,N_42196);
or U44625 (N_44625,N_40091,N_41504);
and U44626 (N_44626,N_41732,N_41251);
xor U44627 (N_44627,N_40936,N_40015);
and U44628 (N_44628,N_40873,N_40302);
nor U44629 (N_44629,N_41433,N_41343);
or U44630 (N_44630,N_41122,N_40457);
nand U44631 (N_44631,N_41774,N_40510);
nand U44632 (N_44632,N_41246,N_42218);
or U44633 (N_44633,N_41296,N_40620);
and U44634 (N_44634,N_40981,N_42292);
nand U44635 (N_44635,N_41194,N_42266);
or U44636 (N_44636,N_41265,N_40678);
nand U44637 (N_44637,N_42138,N_41838);
or U44638 (N_44638,N_42457,N_41664);
nand U44639 (N_44639,N_42355,N_42311);
nor U44640 (N_44640,N_40672,N_40928);
and U44641 (N_44641,N_41768,N_40275);
nand U44642 (N_44642,N_42451,N_41036);
nor U44643 (N_44643,N_41079,N_41228);
xor U44644 (N_44644,N_42145,N_42195);
nor U44645 (N_44645,N_40362,N_41360);
or U44646 (N_44646,N_42316,N_42164);
nand U44647 (N_44647,N_41553,N_40525);
nand U44648 (N_44648,N_42290,N_40856);
nor U44649 (N_44649,N_40913,N_40326);
nand U44650 (N_44650,N_41859,N_40846);
or U44651 (N_44651,N_41687,N_40228);
and U44652 (N_44652,N_41109,N_40779);
xor U44653 (N_44653,N_42070,N_42168);
or U44654 (N_44654,N_40712,N_40734);
nand U44655 (N_44655,N_40980,N_42455);
and U44656 (N_44656,N_41361,N_41134);
and U44657 (N_44657,N_41016,N_41291);
nor U44658 (N_44658,N_42306,N_42195);
and U44659 (N_44659,N_42024,N_40139);
nand U44660 (N_44660,N_41438,N_40340);
and U44661 (N_44661,N_40831,N_40979);
nand U44662 (N_44662,N_40249,N_40309);
or U44663 (N_44663,N_42002,N_41028);
nand U44664 (N_44664,N_40846,N_40604);
xnor U44665 (N_44665,N_40064,N_40774);
xor U44666 (N_44666,N_42344,N_41384);
xnor U44667 (N_44667,N_41081,N_40142);
xor U44668 (N_44668,N_41762,N_41545);
nor U44669 (N_44669,N_42098,N_41063);
xnor U44670 (N_44670,N_40252,N_42410);
nand U44671 (N_44671,N_40608,N_40282);
xor U44672 (N_44672,N_40983,N_40938);
nor U44673 (N_44673,N_41100,N_41860);
and U44674 (N_44674,N_40357,N_42323);
nand U44675 (N_44675,N_41174,N_42100);
xnor U44676 (N_44676,N_40112,N_40876);
nand U44677 (N_44677,N_41773,N_40392);
or U44678 (N_44678,N_40811,N_41235);
or U44679 (N_44679,N_40685,N_42458);
nor U44680 (N_44680,N_42147,N_42295);
and U44681 (N_44681,N_42149,N_41470);
nand U44682 (N_44682,N_40307,N_42219);
nand U44683 (N_44683,N_41270,N_41737);
and U44684 (N_44684,N_41994,N_40103);
nand U44685 (N_44685,N_40221,N_40550);
and U44686 (N_44686,N_40559,N_41879);
and U44687 (N_44687,N_41770,N_41456);
nor U44688 (N_44688,N_42392,N_41200);
nor U44689 (N_44689,N_41509,N_42051);
or U44690 (N_44690,N_40219,N_41192);
xnor U44691 (N_44691,N_40350,N_41284);
and U44692 (N_44692,N_41564,N_41720);
or U44693 (N_44693,N_40373,N_40028);
xor U44694 (N_44694,N_41705,N_40844);
and U44695 (N_44695,N_41355,N_40746);
nor U44696 (N_44696,N_42257,N_41858);
or U44697 (N_44697,N_40028,N_40755);
nor U44698 (N_44698,N_40281,N_40573);
and U44699 (N_44699,N_42202,N_41865);
or U44700 (N_44700,N_42171,N_42418);
nand U44701 (N_44701,N_41864,N_41536);
xnor U44702 (N_44702,N_41597,N_41461);
nor U44703 (N_44703,N_40537,N_41092);
and U44704 (N_44704,N_41587,N_41554);
or U44705 (N_44705,N_40235,N_42042);
nand U44706 (N_44706,N_42047,N_40413);
or U44707 (N_44707,N_40010,N_42197);
or U44708 (N_44708,N_40560,N_40125);
and U44709 (N_44709,N_41097,N_40200);
or U44710 (N_44710,N_40070,N_40407);
nand U44711 (N_44711,N_42419,N_41053);
xnor U44712 (N_44712,N_40429,N_41190);
or U44713 (N_44713,N_40796,N_42067);
and U44714 (N_44714,N_41952,N_42390);
nor U44715 (N_44715,N_41407,N_41745);
nand U44716 (N_44716,N_41980,N_41052);
nand U44717 (N_44717,N_42495,N_41866);
and U44718 (N_44718,N_41905,N_41105);
or U44719 (N_44719,N_42401,N_40703);
nor U44720 (N_44720,N_40371,N_40415);
nand U44721 (N_44721,N_41309,N_40201);
or U44722 (N_44722,N_42433,N_42430);
xor U44723 (N_44723,N_41776,N_40322);
and U44724 (N_44724,N_41125,N_40032);
nor U44725 (N_44725,N_42236,N_41266);
or U44726 (N_44726,N_42416,N_40910);
and U44727 (N_44727,N_41227,N_40568);
and U44728 (N_44728,N_41001,N_40067);
xor U44729 (N_44729,N_40964,N_40769);
xor U44730 (N_44730,N_40599,N_41450);
nor U44731 (N_44731,N_41670,N_41256);
and U44732 (N_44732,N_40163,N_41163);
and U44733 (N_44733,N_41938,N_40793);
and U44734 (N_44734,N_41312,N_40839);
or U44735 (N_44735,N_41893,N_41762);
nand U44736 (N_44736,N_42082,N_41852);
and U44737 (N_44737,N_41784,N_41288);
or U44738 (N_44738,N_41569,N_40155);
nand U44739 (N_44739,N_40456,N_41495);
nand U44740 (N_44740,N_40711,N_40403);
nand U44741 (N_44741,N_41436,N_40739);
xor U44742 (N_44742,N_40398,N_40538);
and U44743 (N_44743,N_40127,N_41245);
xor U44744 (N_44744,N_40286,N_40121);
or U44745 (N_44745,N_40594,N_42131);
nand U44746 (N_44746,N_41182,N_42452);
xnor U44747 (N_44747,N_42452,N_42252);
nand U44748 (N_44748,N_41714,N_41544);
or U44749 (N_44749,N_41421,N_41535);
xor U44750 (N_44750,N_42406,N_42125);
nand U44751 (N_44751,N_41314,N_41588);
nand U44752 (N_44752,N_40120,N_41599);
nand U44753 (N_44753,N_40407,N_42072);
xor U44754 (N_44754,N_42324,N_40701);
or U44755 (N_44755,N_40950,N_42259);
and U44756 (N_44756,N_40378,N_41077);
and U44757 (N_44757,N_42122,N_41662);
and U44758 (N_44758,N_40116,N_40404);
or U44759 (N_44759,N_42375,N_41667);
and U44760 (N_44760,N_42442,N_41559);
or U44761 (N_44761,N_40289,N_40956);
nor U44762 (N_44762,N_41996,N_40779);
and U44763 (N_44763,N_41138,N_40180);
or U44764 (N_44764,N_41848,N_40530);
or U44765 (N_44765,N_41692,N_40767);
nor U44766 (N_44766,N_40760,N_41620);
nor U44767 (N_44767,N_41750,N_40454);
nor U44768 (N_44768,N_41967,N_40462);
and U44769 (N_44769,N_42313,N_41397);
or U44770 (N_44770,N_42269,N_40631);
nor U44771 (N_44771,N_41914,N_41942);
nand U44772 (N_44772,N_40872,N_40930);
nor U44773 (N_44773,N_41464,N_42231);
or U44774 (N_44774,N_40098,N_40414);
xnor U44775 (N_44775,N_40702,N_40690);
or U44776 (N_44776,N_40894,N_40502);
nand U44777 (N_44777,N_42117,N_42440);
xnor U44778 (N_44778,N_41986,N_40767);
nand U44779 (N_44779,N_41831,N_40481);
xnor U44780 (N_44780,N_41668,N_42001);
nor U44781 (N_44781,N_40804,N_41903);
or U44782 (N_44782,N_40804,N_41765);
nand U44783 (N_44783,N_41276,N_41640);
or U44784 (N_44784,N_40463,N_40186);
xor U44785 (N_44785,N_41441,N_42152);
and U44786 (N_44786,N_42234,N_40323);
nor U44787 (N_44787,N_40025,N_40144);
nand U44788 (N_44788,N_42308,N_42075);
or U44789 (N_44789,N_42418,N_41746);
nand U44790 (N_44790,N_40671,N_41704);
or U44791 (N_44791,N_41750,N_40559);
and U44792 (N_44792,N_41662,N_42061);
or U44793 (N_44793,N_42398,N_42372);
or U44794 (N_44794,N_41362,N_40264);
xor U44795 (N_44795,N_41422,N_41848);
xnor U44796 (N_44796,N_41133,N_41934);
xnor U44797 (N_44797,N_41117,N_41035);
nor U44798 (N_44798,N_40089,N_42193);
nor U44799 (N_44799,N_42211,N_40494);
nor U44800 (N_44800,N_41619,N_42256);
nor U44801 (N_44801,N_41231,N_40253);
nor U44802 (N_44802,N_40201,N_41763);
nand U44803 (N_44803,N_40732,N_42170);
nand U44804 (N_44804,N_40024,N_40520);
xor U44805 (N_44805,N_42099,N_42475);
nor U44806 (N_44806,N_41749,N_41695);
xor U44807 (N_44807,N_40772,N_40506);
nor U44808 (N_44808,N_40154,N_40027);
nor U44809 (N_44809,N_41612,N_42001);
or U44810 (N_44810,N_40221,N_42475);
or U44811 (N_44811,N_41197,N_40825);
and U44812 (N_44812,N_40728,N_42004);
xnor U44813 (N_44813,N_41687,N_41445);
xnor U44814 (N_44814,N_40238,N_40888);
nand U44815 (N_44815,N_40860,N_41508);
nand U44816 (N_44816,N_41283,N_42423);
xnor U44817 (N_44817,N_41120,N_42371);
xnor U44818 (N_44818,N_40227,N_40856);
and U44819 (N_44819,N_41197,N_41499);
nor U44820 (N_44820,N_41591,N_41676);
xnor U44821 (N_44821,N_42036,N_40236);
xor U44822 (N_44822,N_40508,N_42193);
and U44823 (N_44823,N_41352,N_41312);
nor U44824 (N_44824,N_42463,N_41431);
nor U44825 (N_44825,N_41306,N_41744);
nand U44826 (N_44826,N_41294,N_40264);
nand U44827 (N_44827,N_41499,N_41748);
nor U44828 (N_44828,N_42376,N_40527);
nor U44829 (N_44829,N_40445,N_41607);
xnor U44830 (N_44830,N_40584,N_40204);
xor U44831 (N_44831,N_41495,N_40401);
xnor U44832 (N_44832,N_40290,N_42148);
or U44833 (N_44833,N_40326,N_40509);
nand U44834 (N_44834,N_41631,N_41819);
nand U44835 (N_44835,N_41896,N_40191);
and U44836 (N_44836,N_40069,N_40675);
or U44837 (N_44837,N_40948,N_40803);
or U44838 (N_44838,N_41381,N_40372);
nand U44839 (N_44839,N_40569,N_40141);
and U44840 (N_44840,N_41465,N_42166);
and U44841 (N_44841,N_42072,N_41692);
and U44842 (N_44842,N_41069,N_40428);
or U44843 (N_44843,N_40004,N_40635);
xnor U44844 (N_44844,N_41432,N_42397);
or U44845 (N_44845,N_40113,N_40392);
nand U44846 (N_44846,N_42301,N_40699);
and U44847 (N_44847,N_41550,N_40853);
nand U44848 (N_44848,N_40321,N_40373);
nor U44849 (N_44849,N_42203,N_40665);
and U44850 (N_44850,N_41263,N_40412);
or U44851 (N_44851,N_42255,N_40600);
or U44852 (N_44852,N_41197,N_42042);
nand U44853 (N_44853,N_42248,N_41377);
and U44854 (N_44854,N_40427,N_41141);
or U44855 (N_44855,N_42376,N_42163);
nand U44856 (N_44856,N_41099,N_41861);
nor U44857 (N_44857,N_40167,N_40620);
nor U44858 (N_44858,N_42377,N_41778);
nand U44859 (N_44859,N_40114,N_42170);
or U44860 (N_44860,N_41832,N_41245);
xnor U44861 (N_44861,N_41954,N_42058);
nand U44862 (N_44862,N_41461,N_42178);
or U44863 (N_44863,N_40288,N_42003);
nor U44864 (N_44864,N_40297,N_41784);
or U44865 (N_44865,N_40079,N_41409);
or U44866 (N_44866,N_42353,N_40750);
and U44867 (N_44867,N_41384,N_41618);
and U44868 (N_44868,N_41148,N_41969);
nand U44869 (N_44869,N_41892,N_42423);
or U44870 (N_44870,N_40773,N_40785);
nor U44871 (N_44871,N_41673,N_40963);
nor U44872 (N_44872,N_40780,N_41141);
xnor U44873 (N_44873,N_40373,N_40435);
nand U44874 (N_44874,N_41692,N_41087);
or U44875 (N_44875,N_41112,N_40776);
nor U44876 (N_44876,N_40868,N_41665);
and U44877 (N_44877,N_41136,N_40279);
nor U44878 (N_44878,N_42346,N_42476);
and U44879 (N_44879,N_40894,N_41588);
nand U44880 (N_44880,N_41999,N_40431);
xor U44881 (N_44881,N_40120,N_40572);
xnor U44882 (N_44882,N_41309,N_41446);
nand U44883 (N_44883,N_41391,N_40135);
or U44884 (N_44884,N_41865,N_41609);
nand U44885 (N_44885,N_41933,N_41196);
nand U44886 (N_44886,N_41660,N_41967);
xor U44887 (N_44887,N_41604,N_40055);
nand U44888 (N_44888,N_40458,N_40611);
and U44889 (N_44889,N_41287,N_42383);
nor U44890 (N_44890,N_40778,N_40703);
or U44891 (N_44891,N_42033,N_41144);
nand U44892 (N_44892,N_40066,N_40531);
nor U44893 (N_44893,N_41662,N_41740);
and U44894 (N_44894,N_40613,N_42058);
or U44895 (N_44895,N_40694,N_40963);
and U44896 (N_44896,N_42392,N_41353);
and U44897 (N_44897,N_41327,N_41257);
xor U44898 (N_44898,N_41483,N_41085);
or U44899 (N_44899,N_41272,N_40160);
nand U44900 (N_44900,N_41469,N_42193);
nand U44901 (N_44901,N_40165,N_41269);
or U44902 (N_44902,N_42066,N_40761);
nor U44903 (N_44903,N_40187,N_40986);
or U44904 (N_44904,N_41526,N_42296);
nand U44905 (N_44905,N_41250,N_41121);
nand U44906 (N_44906,N_42000,N_40842);
nor U44907 (N_44907,N_40452,N_40171);
nand U44908 (N_44908,N_42257,N_42336);
and U44909 (N_44909,N_40214,N_41985);
xnor U44910 (N_44910,N_40611,N_42359);
and U44911 (N_44911,N_40043,N_40761);
xor U44912 (N_44912,N_41705,N_40992);
nand U44913 (N_44913,N_41900,N_40393);
and U44914 (N_44914,N_40273,N_40474);
or U44915 (N_44915,N_42492,N_42003);
nand U44916 (N_44916,N_40304,N_40596);
nand U44917 (N_44917,N_41813,N_40230);
or U44918 (N_44918,N_41757,N_41995);
nand U44919 (N_44919,N_42047,N_41889);
nor U44920 (N_44920,N_42438,N_40562);
xor U44921 (N_44921,N_40568,N_40686);
and U44922 (N_44922,N_40864,N_40566);
xnor U44923 (N_44923,N_40964,N_41435);
xor U44924 (N_44924,N_41277,N_42401);
nand U44925 (N_44925,N_41985,N_40656);
nor U44926 (N_44926,N_41841,N_41589);
nand U44927 (N_44927,N_40354,N_41473);
xnor U44928 (N_44928,N_41149,N_42048);
or U44929 (N_44929,N_40003,N_40654);
nor U44930 (N_44930,N_40939,N_42116);
and U44931 (N_44931,N_40935,N_40503);
nand U44932 (N_44932,N_40610,N_42419);
xor U44933 (N_44933,N_42354,N_41549);
nand U44934 (N_44934,N_42205,N_40531);
and U44935 (N_44935,N_41079,N_40472);
and U44936 (N_44936,N_41828,N_41643);
xor U44937 (N_44937,N_42005,N_40473);
nand U44938 (N_44938,N_41338,N_40530);
nand U44939 (N_44939,N_41475,N_41770);
or U44940 (N_44940,N_41005,N_40657);
nand U44941 (N_44941,N_41563,N_42325);
or U44942 (N_44942,N_40627,N_40065);
xor U44943 (N_44943,N_40598,N_40418);
nor U44944 (N_44944,N_40915,N_40929);
nand U44945 (N_44945,N_40894,N_40839);
or U44946 (N_44946,N_42110,N_41173);
or U44947 (N_44947,N_41986,N_40276);
or U44948 (N_44948,N_40861,N_41772);
nand U44949 (N_44949,N_42303,N_40164);
nor U44950 (N_44950,N_40894,N_40164);
xor U44951 (N_44951,N_40684,N_41393);
nor U44952 (N_44952,N_40503,N_41567);
and U44953 (N_44953,N_40178,N_41395);
nor U44954 (N_44954,N_40733,N_42323);
and U44955 (N_44955,N_40950,N_41977);
nor U44956 (N_44956,N_40135,N_42244);
nand U44957 (N_44957,N_40413,N_40855);
or U44958 (N_44958,N_42127,N_41677);
nand U44959 (N_44959,N_42053,N_42241);
nor U44960 (N_44960,N_42205,N_40058);
xor U44961 (N_44961,N_42018,N_41316);
and U44962 (N_44962,N_40726,N_42211);
or U44963 (N_44963,N_40146,N_40572);
nor U44964 (N_44964,N_40761,N_40456);
and U44965 (N_44965,N_41748,N_42126);
nor U44966 (N_44966,N_42350,N_40862);
nand U44967 (N_44967,N_41455,N_40994);
nand U44968 (N_44968,N_41711,N_41619);
nor U44969 (N_44969,N_42209,N_41565);
nand U44970 (N_44970,N_42383,N_40188);
or U44971 (N_44971,N_40082,N_41830);
nor U44972 (N_44972,N_40518,N_40388);
nand U44973 (N_44973,N_41212,N_41086);
nand U44974 (N_44974,N_40079,N_41338);
nor U44975 (N_44975,N_42233,N_40379);
nor U44976 (N_44976,N_41465,N_41228);
or U44977 (N_44977,N_40416,N_40247);
xnor U44978 (N_44978,N_40106,N_41278);
nand U44979 (N_44979,N_40519,N_41228);
xor U44980 (N_44980,N_41833,N_40472);
xnor U44981 (N_44981,N_41638,N_41929);
nor U44982 (N_44982,N_41075,N_41339);
nor U44983 (N_44983,N_42046,N_40619);
and U44984 (N_44984,N_42056,N_42033);
xor U44985 (N_44985,N_42280,N_41327);
and U44986 (N_44986,N_41708,N_41966);
or U44987 (N_44987,N_41562,N_41498);
and U44988 (N_44988,N_41653,N_40541);
nand U44989 (N_44989,N_41421,N_41291);
nand U44990 (N_44990,N_40372,N_41256);
or U44991 (N_44991,N_42348,N_40848);
nand U44992 (N_44992,N_42448,N_40047);
or U44993 (N_44993,N_40922,N_42042);
nand U44994 (N_44994,N_42461,N_40925);
nand U44995 (N_44995,N_40248,N_40465);
or U44996 (N_44996,N_40061,N_40552);
nor U44997 (N_44997,N_40233,N_42444);
xnor U44998 (N_44998,N_40784,N_41784);
xnor U44999 (N_44999,N_42148,N_41414);
xnor U45000 (N_45000,N_42873,N_44953);
nand U45001 (N_45001,N_44357,N_42992);
and U45002 (N_45002,N_44886,N_44916);
nand U45003 (N_45003,N_44042,N_44547);
and U45004 (N_45004,N_44118,N_43472);
xor U45005 (N_45005,N_43008,N_44555);
and U45006 (N_45006,N_44675,N_44749);
xor U45007 (N_45007,N_42773,N_43526);
or U45008 (N_45008,N_44963,N_44764);
and U45009 (N_45009,N_43805,N_43389);
xnor U45010 (N_45010,N_44709,N_43801);
nor U45011 (N_45011,N_44058,N_44591);
nor U45012 (N_45012,N_44854,N_43005);
and U45013 (N_45013,N_42807,N_43942);
and U45014 (N_45014,N_42579,N_44029);
xnor U45015 (N_45015,N_44410,N_43384);
or U45016 (N_45016,N_42821,N_42916);
or U45017 (N_45017,N_43042,N_43230);
xnor U45018 (N_45018,N_44853,N_43438);
nor U45019 (N_45019,N_44965,N_42869);
nor U45020 (N_45020,N_43348,N_44394);
xnor U45021 (N_45021,N_43945,N_44829);
and U45022 (N_45022,N_43475,N_43811);
nor U45023 (N_45023,N_43433,N_44380);
nand U45024 (N_45024,N_44710,N_43048);
xor U45025 (N_45025,N_43113,N_43376);
xnor U45026 (N_45026,N_42845,N_44503);
nand U45027 (N_45027,N_44570,N_44735);
or U45028 (N_45028,N_42888,N_44657);
or U45029 (N_45029,N_43779,N_43101);
xnor U45030 (N_45030,N_44177,N_43634);
nand U45031 (N_45031,N_43186,N_43733);
and U45032 (N_45032,N_43934,N_43986);
or U45033 (N_45033,N_42609,N_44383);
nor U45034 (N_45034,N_44768,N_43280);
or U45035 (N_45035,N_44517,N_43612);
and U45036 (N_45036,N_43855,N_43735);
nand U45037 (N_45037,N_44573,N_43254);
nor U45038 (N_45038,N_44337,N_43350);
nand U45039 (N_45039,N_43137,N_42859);
or U45040 (N_45040,N_43993,N_44722);
nor U45041 (N_45041,N_42720,N_42668);
nor U45042 (N_45042,N_43754,N_43912);
and U45043 (N_45043,N_43950,N_43498);
and U45044 (N_45044,N_44101,N_44344);
nor U45045 (N_45045,N_42870,N_44393);
nand U45046 (N_45046,N_44435,N_43512);
and U45047 (N_45047,N_44439,N_42721);
nor U45048 (N_45048,N_43323,N_43247);
and U45049 (N_45049,N_43164,N_44149);
nor U45050 (N_45050,N_44103,N_43667);
and U45051 (N_45051,N_42538,N_43202);
nor U45052 (N_45052,N_42717,N_43062);
or U45053 (N_45053,N_44355,N_44524);
or U45054 (N_45054,N_43253,N_44745);
nor U45055 (N_45055,N_44976,N_42800);
or U45056 (N_45056,N_43629,N_43252);
nand U45057 (N_45057,N_44179,N_43771);
nor U45058 (N_45058,N_42600,N_42833);
and U45059 (N_45059,N_44703,N_43145);
nand U45060 (N_45060,N_43259,N_43183);
xor U45061 (N_45061,N_43979,N_44719);
xnor U45062 (N_45062,N_43168,N_42852);
xor U45063 (N_45063,N_43120,N_42585);
xnor U45064 (N_45064,N_42557,N_44212);
and U45065 (N_45065,N_42589,N_44125);
or U45066 (N_45066,N_44673,N_44618);
and U45067 (N_45067,N_44512,N_44197);
and U45068 (N_45068,N_43958,N_44023);
nand U45069 (N_45069,N_44210,N_43239);
xnor U45070 (N_45070,N_44091,N_44952);
nand U45071 (N_45071,N_43535,N_42811);
nand U45072 (N_45072,N_43829,N_43665);
nor U45073 (N_45073,N_42687,N_44548);
nor U45074 (N_45074,N_44040,N_44924);
nor U45075 (N_45075,N_44985,N_44767);
xor U45076 (N_45076,N_42883,N_42723);
nor U45077 (N_45077,N_42655,N_42828);
xnor U45078 (N_45078,N_44265,N_43790);
and U45079 (N_45079,N_42536,N_42549);
xnor U45080 (N_45080,N_42694,N_44217);
nand U45081 (N_45081,N_42994,N_44990);
and U45082 (N_45082,N_43558,N_43234);
xor U45083 (N_45083,N_44496,N_44106);
nor U45084 (N_45084,N_43762,N_44651);
or U45085 (N_45085,N_42565,N_42970);
nor U45086 (N_45086,N_44987,N_44658);
and U45087 (N_45087,N_43179,N_42971);
and U45088 (N_45088,N_43840,N_43166);
nand U45089 (N_45089,N_44504,N_43410);
nor U45090 (N_45090,N_43293,N_42608);
nor U45091 (N_45091,N_42537,N_43455);
xor U45092 (N_45092,N_42508,N_43007);
or U45093 (N_45093,N_43887,N_42896);
or U45094 (N_45094,N_43387,N_43031);
nand U45095 (N_45095,N_44869,N_43814);
nand U45096 (N_45096,N_43714,N_43868);
or U45097 (N_45097,N_44870,N_43778);
or U45098 (N_45098,N_43998,N_44239);
xnor U45099 (N_45099,N_44546,N_43672);
or U45100 (N_45100,N_43644,N_43327);
and U45101 (N_45101,N_43268,N_43631);
or U45102 (N_45102,N_44331,N_44538);
nand U45103 (N_45103,N_44535,N_44529);
nor U45104 (N_45104,N_44689,N_43431);
and U45105 (N_45105,N_43209,N_44053);
or U45106 (N_45106,N_43370,N_43555);
nand U45107 (N_45107,N_44035,N_43205);
nand U45108 (N_45108,N_43755,N_43639);
xnor U45109 (N_45109,N_43622,N_44260);
xnor U45110 (N_45110,N_44859,N_43963);
nor U45111 (N_45111,N_43095,N_43425);
or U45112 (N_45112,N_43161,N_42599);
or U45113 (N_45113,N_44761,N_43856);
nand U45114 (N_45114,N_44758,N_44434);
xor U45115 (N_45115,N_42958,N_42804);
nand U45116 (N_45116,N_43572,N_43484);
and U45117 (N_45117,N_44259,N_42984);
or U45118 (N_45118,N_42552,N_43721);
nor U45119 (N_45119,N_43745,N_44848);
and U45120 (N_45120,N_42766,N_43686);
xnor U45121 (N_45121,N_44222,N_44114);
xnor U45122 (N_45122,N_43310,N_43541);
nor U45123 (N_45123,N_44637,N_44858);
and U45124 (N_45124,N_42707,N_43818);
and U45125 (N_45125,N_44949,N_43724);
and U45126 (N_45126,N_43107,N_44964);
xnor U45127 (N_45127,N_43016,N_44437);
nor U45128 (N_45128,N_43730,N_42654);
or U45129 (N_45129,N_44227,N_44313);
or U45130 (N_45130,N_42629,N_42698);
xnor U45131 (N_45131,N_43808,N_43025);
and U45132 (N_45132,N_43510,N_43369);
xor U45133 (N_45133,N_43079,N_43276);
and U45134 (N_45134,N_42582,N_43028);
or U45135 (N_45135,N_43368,N_44052);
nand U45136 (N_45136,N_44830,N_44624);
and U45137 (N_45137,N_42882,N_42685);
nand U45138 (N_45138,N_42851,N_43791);
xor U45139 (N_45139,N_44702,N_43412);
and U45140 (N_45140,N_43199,N_44378);
or U45141 (N_45141,N_44528,N_43203);
nand U45142 (N_45142,N_44010,N_44839);
or U45143 (N_45143,N_43121,N_44770);
nand U45144 (N_45144,N_44261,N_44065);
nor U45145 (N_45145,N_42729,N_43657);
nor U45146 (N_45146,N_42667,N_42808);
nand U45147 (N_45147,N_42843,N_43722);
and U45148 (N_45148,N_43608,N_43561);
xnor U45149 (N_45149,N_42719,N_42841);
xor U45150 (N_45150,N_42893,N_44801);
nand U45151 (N_45151,N_43875,N_42592);
and U45152 (N_45152,N_42554,N_44384);
and U45153 (N_45153,N_42682,N_43737);
nor U45154 (N_45154,N_44252,N_42510);
nand U45155 (N_45155,N_43692,N_44293);
nand U45156 (N_45156,N_42929,N_44283);
nor U45157 (N_45157,N_44073,N_44055);
xnor U45158 (N_45158,N_43898,N_42849);
nor U45159 (N_45159,N_44865,N_43590);
nand U45160 (N_45160,N_42948,N_43528);
or U45161 (N_45161,N_43816,N_44138);
nand U45162 (N_45162,N_43317,N_43577);
or U45163 (N_45163,N_44194,N_43351);
and U45164 (N_45164,N_42786,N_43479);
xnor U45165 (N_45165,N_43652,N_42923);
nor U45166 (N_45166,N_42933,N_44802);
nor U45167 (N_45167,N_43749,N_44559);
and U45168 (N_45168,N_44979,N_44287);
or U45169 (N_45169,N_43006,N_44959);
and U45170 (N_45170,N_44905,N_44778);
nand U45171 (N_45171,N_44751,N_43428);
and U45172 (N_45172,N_43797,N_43379);
nand U45173 (N_45173,N_42708,N_43493);
or U45174 (N_45174,N_43573,N_42605);
nor U45175 (N_45175,N_42699,N_43229);
or U45176 (N_45176,N_44338,N_43491);
xnor U45177 (N_45177,N_43576,N_44697);
and U45178 (N_45178,N_44968,N_43090);
nand U45179 (N_45179,N_44068,N_44551);
xor U45180 (N_45180,N_43078,N_42574);
or U45181 (N_45181,N_42922,N_43309);
nor U45182 (N_45182,N_42817,N_42701);
nor U45183 (N_45183,N_43546,N_44809);
nand U45184 (N_45184,N_44345,N_44371);
xnor U45185 (N_45185,N_44404,N_43262);
and U45186 (N_45186,N_44954,N_42691);
and U45187 (N_45187,N_43523,N_44774);
nor U45188 (N_45188,N_43878,N_43073);
nor U45189 (N_45189,N_43143,N_43093);
nand U45190 (N_45190,N_44124,N_43655);
nor U45191 (N_45191,N_43609,N_44526);
nand U45192 (N_45192,N_43944,N_42753);
nand U45193 (N_45193,N_43045,N_44539);
nand U45194 (N_45194,N_44776,N_44097);
nor U45195 (N_45195,N_44860,N_44593);
nor U45196 (N_45196,N_43699,N_43513);
nand U45197 (N_45197,N_42546,N_44084);
nor U45198 (N_45198,N_43988,N_44022);
xnor U45199 (N_45199,N_43138,N_43727);
xor U45200 (N_45200,N_44942,N_44291);
nand U45201 (N_45201,N_44113,N_44933);
nand U45202 (N_45202,N_43163,N_44013);
and U45203 (N_45203,N_42656,N_43751);
xor U45204 (N_45204,N_43647,N_43236);
and U45205 (N_45205,N_43420,N_44186);
nor U45206 (N_45206,N_42938,N_44137);
xor U45207 (N_45207,N_43447,N_43874);
or U45208 (N_45208,N_44929,N_43424);
or U45209 (N_45209,N_44750,N_42521);
xnor U45210 (N_45210,N_44468,N_44765);
nor U45211 (N_45211,N_44604,N_43244);
nand U45212 (N_45212,N_42799,N_44007);
nor U45213 (N_45213,N_44671,N_43112);
nand U45214 (N_45214,N_44203,N_44397);
xor U45215 (N_45215,N_42530,N_43683);
or U45216 (N_45216,N_43863,N_44989);
nand U45217 (N_45217,N_42746,N_44821);
and U45218 (N_45218,N_42739,N_43966);
or U45219 (N_45219,N_44707,N_43810);
and U45220 (N_45220,N_44188,N_43845);
xnor U45221 (N_45221,N_44237,N_44004);
nor U45222 (N_45222,N_42829,N_43905);
or U45223 (N_45223,N_44405,N_44098);
nand U45224 (N_45224,N_42714,N_43195);
xnor U45225 (N_45225,N_44320,N_44567);
and U45226 (N_45226,N_43766,N_44067);
or U45227 (N_45227,N_44921,N_43036);
nor U45228 (N_45228,N_44588,N_44134);
nor U45229 (N_45229,N_44792,N_44285);
or U45230 (N_45230,N_44824,N_44835);
xnor U45231 (N_45231,N_42596,N_43128);
and U45232 (N_45232,N_44896,N_44248);
nand U45233 (N_45233,N_42594,N_44466);
and U45234 (N_45234,N_44389,N_42503);
and U45235 (N_45235,N_43442,N_43058);
nor U45236 (N_45236,N_42881,N_43292);
nor U45237 (N_45237,N_43613,N_43518);
and U45238 (N_45238,N_44318,N_43047);
nor U45239 (N_45239,N_44780,N_42597);
and U45240 (N_45240,N_43775,N_42620);
nor U45241 (N_45241,N_42632,N_44174);
xnor U45242 (N_45242,N_43106,N_44568);
nand U45243 (N_45243,N_42640,N_42975);
nor U45244 (N_45244,N_42662,N_43592);
nor U45245 (N_45245,N_44928,N_44935);
nor U45246 (N_45246,N_44109,N_43467);
nand U45247 (N_45247,N_43499,N_43357);
nor U45248 (N_45248,N_42617,N_42903);
nand U45249 (N_45249,N_44864,N_44872);
or U45250 (N_45250,N_43663,N_44643);
or U45251 (N_45251,N_44172,N_43345);
xnor U45252 (N_45252,N_43397,N_43710);
or U45253 (N_45253,N_42778,N_44790);
nor U45254 (N_45254,N_44223,N_43802);
nand U45255 (N_45255,N_44043,N_43873);
nor U45256 (N_45256,N_44594,N_44514);
or U45257 (N_45257,N_44336,N_43536);
or U45258 (N_45258,N_42658,N_44322);
nand U45259 (N_45259,N_42688,N_42755);
xnor U45260 (N_45260,N_43275,N_43360);
nor U45261 (N_45261,N_44471,N_43642);
nand U45262 (N_45262,N_44253,N_42835);
and U45263 (N_45263,N_42587,N_43094);
or U45264 (N_45264,N_43598,N_44540);
and U45265 (N_45265,N_44522,N_43928);
or U45266 (N_45266,N_44730,N_43325);
nor U45267 (N_45267,N_42732,N_44789);
nor U45268 (N_45268,N_42533,N_42615);
nand U45269 (N_45269,N_43872,N_44332);
nor U45270 (N_45270,N_44421,N_43606);
nand U45271 (N_45271,N_44569,N_43153);
nand U45272 (N_45272,N_43921,N_44906);
nand U45273 (N_45273,N_43626,N_44925);
xor U45274 (N_45274,N_43838,N_42637);
or U45275 (N_45275,N_43474,N_43593);
xor U45276 (N_45276,N_44837,N_43911);
nor U45277 (N_45277,N_43313,N_44202);
or U45278 (N_45278,N_42718,N_42974);
or U45279 (N_45279,N_42818,N_44465);
nor U45280 (N_45280,N_42993,N_44305);
or U45281 (N_45281,N_43251,N_44717);
and U45282 (N_45282,N_43466,N_43198);
nand U45283 (N_45283,N_43933,N_44088);
nor U45284 (N_45284,N_44836,N_43955);
or U45285 (N_45285,N_42805,N_42567);
and U45286 (N_45286,N_44324,N_43901);
and U45287 (N_45287,N_43406,N_44883);
xor U45288 (N_45288,N_44492,N_44489);
nand U45289 (N_45289,N_43366,N_43653);
nand U45290 (N_45290,N_43991,N_44160);
nand U45291 (N_45291,N_43638,N_44303);
xnor U45292 (N_45292,N_43256,N_44585);
xnor U45293 (N_45293,N_43200,N_43689);
or U45294 (N_45294,N_44525,N_44556);
nand U45295 (N_45295,N_44108,N_43937);
xnor U45296 (N_45296,N_42797,N_44783);
nand U45297 (N_45297,N_43527,N_43462);
or U45298 (N_45298,N_43372,N_42623);
and U45299 (N_45299,N_42936,N_44294);
nand U45300 (N_45300,N_43483,N_44826);
nor U45301 (N_45301,N_43820,N_42751);
or U45302 (N_45302,N_43122,N_43516);
nand U45303 (N_45303,N_43550,N_44477);
or U45304 (N_45304,N_42966,N_43216);
or U45305 (N_45305,N_44028,N_44610);
and U45306 (N_45306,N_42782,N_43312);
nor U45307 (N_45307,N_43448,N_44617);
nand U45308 (N_45308,N_43114,N_44037);
and U45309 (N_45309,N_42573,N_43271);
nor U45310 (N_45310,N_43437,N_44667);
nor U45311 (N_45311,N_44796,N_42507);
xor U45312 (N_45312,N_43329,N_44150);
xor U45313 (N_45313,N_43789,N_44449);
nand U45314 (N_45314,N_43731,N_43570);
xnor U45315 (N_45315,N_43578,N_43990);
and U45316 (N_45316,N_43450,N_43929);
nor U45317 (N_45317,N_42969,N_43495);
xor U45318 (N_45318,N_42722,N_43426);
nor U45319 (N_45319,N_44025,N_44999);
or U45320 (N_45320,N_44629,N_43037);
nor U45321 (N_45321,N_43783,N_43883);
nor U45322 (N_45322,N_44143,N_44934);
nand U45323 (N_45323,N_44133,N_42924);
and U45324 (N_45324,N_44481,N_43060);
and U45325 (N_45325,N_42611,N_44470);
nand U45326 (N_45326,N_43897,N_43010);
nand U45327 (N_45327,N_44360,N_44572);
and U45328 (N_45328,N_42988,N_43242);
xnor U45329 (N_45329,N_44507,N_42560);
nor U45330 (N_45330,N_43481,N_43920);
nand U45331 (N_45331,N_43063,N_43110);
or U45332 (N_45332,N_44005,N_44152);
nor U45333 (N_45333,N_44206,N_42506);
and U45334 (N_45334,N_42648,N_43116);
nand U45335 (N_45335,N_44480,N_43674);
nand U45336 (N_45336,N_42990,N_44092);
and U45337 (N_45337,N_42520,N_44180);
xor U45338 (N_45338,N_43068,N_44533);
nor U45339 (N_45339,N_44048,N_43049);
and U45340 (N_45340,N_44416,N_44582);
xnor U45341 (N_45341,N_44662,N_44157);
and U45342 (N_45342,N_42928,N_43477);
xnor U45343 (N_45343,N_43334,N_42588);
nand U45344 (N_45344,N_44445,N_43651);
and U45345 (N_45345,N_43824,N_44427);
xnor U45346 (N_45346,N_42539,N_43524);
nand U45347 (N_45347,N_43458,N_43566);
or U45348 (N_45348,N_43908,N_44376);
nor U45349 (N_45349,N_43785,N_44856);
xnor U45350 (N_45350,N_44940,N_43235);
and U45351 (N_45351,N_43147,N_42680);
and U45352 (N_45352,N_43358,N_42514);
or U45353 (N_45353,N_42518,N_42952);
nand U45354 (N_45354,N_44482,N_43947);
or U45355 (N_45355,N_43548,N_44611);
nand U45356 (N_45356,N_43972,N_43764);
or U45357 (N_45357,N_43926,N_42932);
nor U45358 (N_45358,N_43021,N_44945);
and U45359 (N_45359,N_43086,N_42709);
xnor U45360 (N_45360,N_43607,N_42953);
nand U45361 (N_45361,N_43852,N_43050);
or U45362 (N_45362,N_44096,N_43034);
or U45363 (N_45363,N_44415,N_42505);
or U45364 (N_45364,N_43540,N_44142);
nand U45365 (N_45365,N_42855,N_43580);
xor U45366 (N_45366,N_43587,N_44557);
nor U45367 (N_45367,N_44909,N_43890);
xnor U45368 (N_45368,N_43715,N_44105);
xnor U45369 (N_45369,N_43338,N_42591);
nor U45370 (N_45370,N_42734,N_42889);
or U45371 (N_45371,N_42775,N_44061);
nor U45372 (N_45372,N_44904,N_42525);
or U45373 (N_45373,N_43367,N_44669);
nand U45374 (N_45374,N_42780,N_44732);
nand U45375 (N_45375,N_44050,N_44725);
or U45376 (N_45376,N_44456,N_43359);
and U45377 (N_45377,N_42972,N_43018);
and U45378 (N_45378,N_43851,N_43858);
xor U45379 (N_45379,N_43173,N_44930);
nor U45380 (N_45380,N_44807,N_43825);
nor U45381 (N_45381,N_44027,N_42747);
nor U45382 (N_45382,N_44325,N_43502);
xor U45383 (N_45383,N_42523,N_44230);
xnor U45384 (N_45384,N_44104,N_44740);
or U45385 (N_45385,N_42858,N_42765);
xnor U45386 (N_45386,N_42572,N_44431);
and U45387 (N_45387,N_43083,N_43889);
or U45388 (N_45388,N_43115,N_42693);
nor U45389 (N_45389,N_43418,N_43720);
xor U45390 (N_45390,N_44957,N_43579);
nor U45391 (N_45391,N_43102,N_43411);
nand U45392 (N_45392,N_44419,N_44799);
nor U45393 (N_45393,N_43954,N_43632);
or U45394 (N_45394,N_43662,N_43181);
xnor U45395 (N_45395,N_42850,N_43640);
or U45396 (N_45396,N_43286,N_44918);
or U45397 (N_45397,N_44135,N_43306);
nand U45398 (N_45398,N_44340,N_42844);
xnor U45399 (N_45399,N_43969,N_43193);
nand U45400 (N_45400,N_43105,N_42862);
nand U45401 (N_45401,N_43817,N_42559);
nor U45402 (N_45402,N_44739,N_43222);
nor U45403 (N_45403,N_43196,N_43178);
or U45404 (N_45404,N_43245,N_44314);
xor U45405 (N_45405,N_44298,N_42659);
nand U45406 (N_45406,N_43054,N_44011);
nor U45407 (N_45407,N_43213,N_44654);
nand U45408 (N_45408,N_43935,N_43756);
and U45409 (N_45409,N_42853,N_42622);
nand U45410 (N_45410,N_43999,N_44008);
xor U45411 (N_45411,N_43206,N_44286);
and U45412 (N_45412,N_43815,N_44012);
nor U45413 (N_45413,N_44615,N_43364);
xnor U45414 (N_45414,N_43487,N_42663);
nor U45415 (N_45415,N_43670,N_43780);
or U45416 (N_45416,N_43291,N_43353);
and U45417 (N_45417,N_42827,N_43882);
or U45418 (N_45418,N_44939,N_44351);
and U45419 (N_45419,N_43604,N_43959);
or U45420 (N_45420,N_43347,N_42957);
xor U45421 (N_45421,N_44199,N_43597);
and U45422 (N_45422,N_43332,N_44763);
or U45423 (N_45423,N_43223,N_42540);
xor U45424 (N_45424,N_44505,N_42743);
and U45425 (N_45425,N_43980,N_44882);
nor U45426 (N_45426,N_42583,N_43461);
and U45427 (N_45427,N_42907,N_44605);
nor U45428 (N_45428,N_43671,N_44851);
nor U45429 (N_45429,N_44912,N_43500);
xnor U45430 (N_45430,N_43123,N_44692);
xnor U45431 (N_45431,N_43281,N_44256);
xnor U45432 (N_45432,N_43261,N_44531);
nor U45433 (N_45433,N_42534,N_43155);
nand U45434 (N_45434,N_43501,N_43396);
and U45435 (N_45435,N_44146,N_42555);
xor U45436 (N_45436,N_42737,N_43250);
nand U45437 (N_45437,N_43563,N_43556);
xor U45438 (N_45438,N_44258,N_43097);
nand U45439 (N_45439,N_44122,N_44843);
nand U45440 (N_45440,N_42898,N_42606);
and U45441 (N_45441,N_43430,N_42779);
xor U45442 (N_45442,N_43243,N_43881);
nand U45443 (N_45443,N_42711,N_44576);
nand U45444 (N_45444,N_44874,N_44762);
xor U45445 (N_45445,N_42959,N_43706);
nor U45446 (N_45446,N_44867,N_42905);
nand U45447 (N_45447,N_43521,N_43956);
xor U45448 (N_45448,N_43591,N_42660);
nor U45449 (N_45449,N_44245,N_43488);
and U45450 (N_45450,N_44166,N_44509);
xor U45451 (N_45451,N_44094,N_43772);
and U45452 (N_45452,N_44386,N_43071);
xnor U45453 (N_45453,N_42946,N_44238);
or U45454 (N_45454,N_44664,N_44232);
nor U45455 (N_45455,N_43641,N_44897);
nand U45456 (N_45456,N_44603,N_44564);
and U45457 (N_45457,N_44759,N_44804);
and U45458 (N_45458,N_43554,N_42621);
and U45459 (N_45459,N_43207,N_42749);
nand U45460 (N_45460,N_44246,N_42806);
and U45461 (N_45461,N_43361,N_43057);
nor U45462 (N_45462,N_43322,N_43221);
nand U45463 (N_45463,N_43392,N_44808);
xor U45464 (N_45464,N_42877,N_44006);
or U45465 (N_45465,N_44661,N_44625);
or U45466 (N_45466,N_43103,N_44970);
nand U45467 (N_45467,N_44417,N_42677);
and U45468 (N_45468,N_44877,N_44969);
xnor U45469 (N_45469,N_42774,N_44626);
nand U45470 (N_45470,N_43408,N_44242);
nand U45471 (N_45471,N_43575,N_43489);
xnor U45472 (N_45472,N_44960,N_44892);
nand U45473 (N_45473,N_43543,N_44534);
and U45474 (N_45474,N_44737,N_43932);
and U45475 (N_45475,N_44448,N_43473);
or U45476 (N_45476,N_44558,N_44634);
xor U45477 (N_45477,N_43434,N_44411);
nor U45478 (N_45478,N_44296,N_44711);
or U45479 (N_45479,N_42967,N_44147);
xnor U45480 (N_45480,N_43834,N_44962);
or U45481 (N_45481,N_44353,N_42748);
or U45482 (N_45482,N_42684,N_42736);
nand U45483 (N_45483,N_43871,N_44346);
nand U45484 (N_45484,N_42979,N_44323);
or U45485 (N_45485,N_43660,N_44395);
nor U45486 (N_45486,N_42991,N_43380);
xor U45487 (N_45487,N_43398,N_43973);
or U45488 (N_45488,N_43821,N_43844);
xor U45489 (N_45489,N_42910,N_44024);
or U45490 (N_45490,N_44599,N_43189);
nor U45491 (N_45491,N_43174,N_44129);
nand U45492 (N_45492,N_43080,N_44579);
nor U45493 (N_45493,N_44335,N_42511);
nor U45494 (N_45494,N_42801,N_43864);
nand U45495 (N_45495,N_44064,N_44342);
or U45496 (N_45496,N_44871,N_43069);
or U45497 (N_45497,N_44880,N_42603);
or U45498 (N_45498,N_44312,N_44900);
and U45499 (N_45499,N_43589,N_43055);
nor U45500 (N_45500,N_44363,N_43318);
nand U45501 (N_45501,N_44844,N_43656);
nand U45502 (N_45502,N_43072,N_42716);
nor U45503 (N_45503,N_44060,N_44855);
nand U45504 (N_45504,N_43454,N_43204);
nand U45505 (N_45505,N_42604,N_43316);
nor U45506 (N_45506,N_42816,N_44267);
and U45507 (N_45507,N_44973,N_44045);
nand U45508 (N_45508,N_44898,N_43004);
nand U45509 (N_45509,N_44816,N_44278);
nor U45510 (N_45510,N_42781,N_44781);
nand U45511 (N_45511,N_44527,N_44814);
and U45512 (N_45512,N_42762,N_43218);
or U45513 (N_45513,N_43635,N_42683);
and U45514 (N_45514,N_44823,N_43266);
or U45515 (N_45515,N_44229,N_43070);
nor U45516 (N_45516,N_43661,N_43040);
nand U45517 (N_45517,N_43951,N_43354);
nand U45518 (N_45518,N_42931,N_43977);
or U45519 (N_45519,N_44670,N_44701);
xor U45520 (N_45520,N_44099,N_44329);
or U45521 (N_45521,N_43098,N_42543);
nand U45522 (N_45522,N_43038,N_43377);
or U45523 (N_45523,N_43127,N_44414);
xor U45524 (N_45524,N_43065,N_43767);
or U45525 (N_45525,N_43650,N_43300);
and U45526 (N_45526,N_44473,N_44330);
xnor U45527 (N_45527,N_43212,N_43630);
nor U45528 (N_45528,N_43586,N_44163);
and U45529 (N_45529,N_43141,N_43809);
and U45530 (N_45530,N_44676,N_44650);
nand U45531 (N_45531,N_44875,N_44630);
nor U45532 (N_45532,N_42704,N_43403);
nand U45533 (N_45533,N_42619,N_42876);
xor U45534 (N_45534,N_44075,N_43939);
xnor U45535 (N_45535,N_44300,N_44521);
nand U45536 (N_45536,N_42618,N_43492);
nor U45537 (N_45537,N_44966,N_43981);
or U45538 (N_45538,N_43533,N_44015);
or U45539 (N_45539,N_44622,N_43728);
nor U45540 (N_45540,N_44200,N_43227);
nor U45541 (N_45541,N_42879,N_43806);
nor U45542 (N_45542,N_43758,N_44991);
nor U45543 (N_45543,N_44447,N_43509);
nor U45544 (N_45544,N_43248,N_43659);
nor U45545 (N_45545,N_43719,N_44698);
xor U45546 (N_45546,N_43995,N_42965);
nand U45547 (N_45547,N_44696,N_42638);
and U45548 (N_45548,N_43539,N_44167);
nor U45549 (N_45549,N_43615,N_44619);
nor U45550 (N_45550,N_44406,N_42909);
or U45551 (N_45551,N_42919,N_44491);
nand U45552 (N_45552,N_42783,N_42954);
nor U45553 (N_45553,N_42942,N_43588);
or U45554 (N_45554,N_44276,N_43305);
and U45555 (N_45555,N_43320,N_44116);
xnor U45556 (N_45556,N_44888,N_44943);
or U45557 (N_45557,N_44545,N_43026);
and U45558 (N_45558,N_43628,N_44641);
and U45559 (N_45559,N_44047,N_43382);
nand U45560 (N_45560,N_44430,N_44056);
nor U45561 (N_45561,N_44811,N_43508);
and U45562 (N_45562,N_43023,N_43765);
xnor U45563 (N_45563,N_42790,N_42610);
or U45564 (N_45564,N_43800,N_42627);
xor U45565 (N_45565,N_43033,N_44082);
or U45566 (N_45566,N_42545,N_44178);
and U45567 (N_45567,N_44370,N_44034);
nand U45568 (N_45568,N_43167,N_43804);
or U45569 (N_45569,N_44021,N_44429);
or U45570 (N_45570,N_44714,N_43614);
and U45571 (N_45571,N_43032,N_43043);
nor U45572 (N_45572,N_42625,N_44306);
nand U45573 (N_45573,N_42689,N_43443);
and U45574 (N_45574,N_44895,N_42575);
nand U45575 (N_45575,N_42894,N_44126);
and U45576 (N_45576,N_42669,N_44828);
nor U45577 (N_45577,N_44998,N_43859);
or U45578 (N_45578,N_43549,N_43108);
and U45579 (N_45579,N_42927,N_43562);
nand U45580 (N_45580,N_44317,N_44753);
nor U45581 (N_45581,N_44805,N_44716);
or U45582 (N_45582,N_43303,N_44636);
nor U45583 (N_45583,N_44787,N_44341);
and U45584 (N_45584,N_43342,N_43409);
nand U45585 (N_45585,N_43744,N_44734);
or U45586 (N_45586,N_43910,N_42628);
xor U45587 (N_45587,N_43417,N_44986);
xor U45588 (N_45588,N_44086,N_43485);
xor U45589 (N_45589,N_43246,N_43399);
nor U45590 (N_45590,N_44520,N_44284);
nor U45591 (N_45591,N_42784,N_43716);
and U45592 (N_45592,N_43111,N_43970);
and U45593 (N_45593,N_42921,N_43344);
or U45594 (N_45594,N_43289,N_44852);
xnor U45595 (N_45595,N_44391,N_44530);
xnor U45596 (N_45596,N_44659,N_43341);
xor U45597 (N_45597,N_44295,N_44274);
or U45598 (N_45598,N_42802,N_43265);
or U45599 (N_45599,N_44182,N_42524);
and U45600 (N_45600,N_43228,N_44412);
xnor U45601 (N_45601,N_43441,N_42580);
and U45602 (N_45602,N_42908,N_43020);
nor U45603 (N_45603,N_42760,N_43807);
xnor U45604 (N_45604,N_42745,N_42744);
and U45605 (N_45605,N_43130,N_43717);
nand U45606 (N_45606,N_42769,N_43150);
xor U45607 (N_45607,N_44782,N_44656);
nand U45608 (N_45608,N_44089,N_44127);
or U45609 (N_45609,N_43676,N_43819);
xor U45610 (N_45610,N_42650,N_44117);
xnor U45611 (N_45611,N_43077,N_43769);
nand U45612 (N_45612,N_43846,N_42529);
nor U45613 (N_45613,N_44102,N_43279);
and U45614 (N_45614,N_43238,N_44159);
and U45615 (N_45615,N_42839,N_44361);
nand U45616 (N_45616,N_44155,N_44894);
nor U45617 (N_45617,N_43449,N_44899);
and U45618 (N_45618,N_44668,N_43696);
or U45619 (N_45619,N_44153,N_42768);
xor U45620 (N_45620,N_44077,N_43506);
xor U45621 (N_45621,N_43961,N_43994);
nand U45622 (N_45622,N_43964,N_42874);
and U45623 (N_45623,N_43511,N_42750);
nor U45624 (N_45624,N_43909,N_43948);
nand U45625 (N_45625,N_43432,N_43328);
xor U45626 (N_45626,N_44794,N_44185);
xor U45627 (N_45627,N_42985,N_44250);
nand U45628 (N_45628,N_44409,N_43451);
nor U45629 (N_45629,N_43708,N_43085);
nor U45630 (N_45630,N_43215,N_42836);
or U45631 (N_45631,N_42528,N_44078);
nand U45632 (N_45632,N_44218,N_42884);
and U45633 (N_45633,N_43784,N_43260);
nor U45634 (N_45634,N_44822,N_44192);
xor U45635 (N_45635,N_43984,N_42798);
and U45636 (N_45636,N_44868,N_44176);
nor U45637 (N_45637,N_43126,N_42725);
or U45638 (N_45638,N_43997,N_44700);
or U45639 (N_45639,N_44786,N_43974);
xor U45640 (N_45640,N_44690,N_43053);
nand U45641 (N_45641,N_43148,N_43585);
and U45642 (N_45642,N_43637,N_42551);
or U45643 (N_45643,N_43700,N_43552);
and U45644 (N_45644,N_43940,N_42885);
or U45645 (N_45645,N_44665,N_44565);
xnor U45646 (N_45646,N_42566,N_42724);
xnor U45647 (N_45647,N_44262,N_42643);
xnor U45648 (N_45648,N_42764,N_43918);
or U45649 (N_45649,N_43832,N_43666);
nor U45650 (N_45650,N_43738,N_44403);
or U45651 (N_45651,N_43378,N_44271);
nand U45652 (N_45652,N_44738,N_42631);
xnor U45653 (N_45653,N_43046,N_42501);
nor U45654 (N_45654,N_42978,N_43916);
nor U45655 (N_45655,N_43210,N_42875);
or U45656 (N_45656,N_44561,N_42848);
xor U45657 (N_45657,N_44461,N_44587);
xor U45658 (N_45658,N_43225,N_43680);
or U45659 (N_45659,N_44213,N_43930);
xnor U45660 (N_45660,N_42598,N_44866);
nand U45661 (N_45661,N_44623,N_43362);
or U45662 (N_45662,N_42767,N_42624);
or U45663 (N_45663,N_43761,N_44100);
nor U45664 (N_45664,N_44920,N_43600);
nor U45665 (N_45665,N_43893,N_44399);
and U45666 (N_45666,N_43854,N_43695);
nor U45667 (N_45667,N_44402,N_44820);
nor U45668 (N_45668,N_44847,N_44059);
or U45669 (N_45669,N_44779,N_42847);
or U45670 (N_45670,N_43645,N_44915);
nor U45671 (N_45671,N_43278,N_42860);
and U45672 (N_45672,N_43544,N_42541);
nor U45673 (N_45673,N_43365,N_43480);
nor U45674 (N_45674,N_44139,N_44597);
nand U45675 (N_45675,N_44297,N_42581);
nand U45676 (N_45676,N_43886,N_44132);
or U45677 (N_45677,N_44876,N_44066);
or U45678 (N_45678,N_43673,N_43701);
nor U45679 (N_45679,N_42980,N_44479);
nand U45680 (N_45680,N_42616,N_42854);
nand U45681 (N_45681,N_44518,N_43975);
or U45682 (N_45682,N_43843,N_44574);
xnor U45683 (N_45683,N_44884,N_42703);
and U45684 (N_45684,N_42666,N_44975);
xor U45685 (N_45685,N_43401,N_42920);
xnor U45686 (N_45686,N_43763,N_43240);
or U45687 (N_45687,N_42586,N_42825);
and U45688 (N_45688,N_43092,N_44677);
xor U45689 (N_45689,N_44946,N_43496);
xor U45690 (N_45690,N_42866,N_42785);
nor U45691 (N_45691,N_43336,N_44502);
nor U45692 (N_45692,N_44922,N_43985);
xor U45693 (N_45693,N_43837,N_43847);
or U45694 (N_45694,N_42633,N_42890);
xnor U45695 (N_45695,N_44878,N_42613);
nand U45696 (N_45696,N_42842,N_43452);
and U45697 (N_45697,N_43989,N_44598);
and U45698 (N_45698,N_44846,N_43171);
xor U45699 (N_45699,N_43601,N_43505);
or U45700 (N_45700,N_44343,N_43390);
xor U45701 (N_45701,N_43453,N_42700);
and U45702 (N_45702,N_43132,N_43056);
xor U45703 (N_45703,N_44085,N_42532);
or U45704 (N_45704,N_44356,N_43117);
nor U45705 (N_45705,N_44464,N_43142);
and U45706 (N_45706,N_43233,N_44679);
nand U45707 (N_45707,N_44632,N_44813);
nand U45708 (N_45708,N_44289,N_43159);
or U45709 (N_45709,N_43734,N_44196);
nor U45710 (N_45710,N_43009,N_43795);
or U45711 (N_45711,N_43664,N_44352);
nand U45712 (N_45712,N_42726,N_43707);
nor U45713 (N_45713,N_44220,N_44506);
or U45714 (N_45714,N_44074,N_42809);
nand U45715 (N_45715,N_43220,N_44368);
or U45716 (N_45716,N_43217,N_44683);
and U45717 (N_45717,N_43182,N_43041);
or U45718 (N_45718,N_42939,N_44956);
and U45719 (N_45719,N_44713,N_42796);
and U45720 (N_45720,N_42602,N_44553);
xnor U45721 (N_45721,N_43002,N_44319);
xnor U45722 (N_45722,N_43427,N_43232);
nand U45723 (N_45723,N_44207,N_44638);
xor U45724 (N_45724,N_44862,N_43760);
nand U45725 (N_45725,N_43781,N_44460);
nor U45726 (N_45726,N_43627,N_42897);
and U45727 (N_45727,N_43605,N_43074);
nor U45728 (N_45728,N_44401,N_43465);
nor U45729 (N_45729,N_43559,N_44684);
nand U45730 (N_45730,N_44081,N_43402);
xnor U45731 (N_45731,N_44771,N_42943);
nor U45732 (N_45732,N_44168,N_43743);
nand U45733 (N_45733,N_44408,N_44981);
xnor U45734 (N_45734,N_44057,N_43776);
and U45735 (N_45735,N_43992,N_43100);
nor U45736 (N_45736,N_43726,N_44542);
xnor U45737 (N_45737,N_44648,N_44704);
nor U45738 (N_45738,N_42526,N_42961);
xnor U45739 (N_45739,N_42856,N_42872);
xor U45740 (N_45740,N_42824,N_44112);
xnor U45741 (N_45741,N_42956,N_43169);
and U45742 (N_45742,N_44387,N_44812);
xor U45743 (N_45743,N_43698,N_43324);
and U45744 (N_45744,N_44815,N_43436);
nand U45745 (N_45745,N_43917,N_44381);
nor U45746 (N_45746,N_43862,N_43374);
or U45747 (N_45747,N_44901,N_44014);
and U45748 (N_45748,N_44349,N_44311);
xnor U45749 (N_45749,N_44845,N_43035);
nor U45750 (N_45750,N_42789,N_42675);
nor U45751 (N_45751,N_43165,N_44649);
and U45752 (N_45752,N_43064,N_44631);
or U45753 (N_45753,N_43191,N_43295);
nand U45754 (N_45754,N_42901,N_44307);
nand U45755 (N_45755,N_43914,N_44728);
or U45756 (N_45756,N_43214,N_42867);
xor U45757 (N_45757,N_43624,N_43445);
nand U45758 (N_45758,N_43617,N_43219);
and U45759 (N_45759,N_42676,N_43383);
xor U45760 (N_45760,N_42934,N_43407);
nand U45761 (N_45761,N_43768,N_42819);
or U45762 (N_45762,N_42519,N_43965);
or U45763 (N_45763,N_43793,N_44201);
nor U45764 (N_45764,N_42595,N_43162);
xnor U45765 (N_45765,N_44944,N_43534);
or U45766 (N_45766,N_44827,N_42820);
nor U45767 (N_45767,N_44422,N_42563);
xnor U45768 (N_45768,N_44020,N_44093);
nor U45769 (N_45769,N_44187,N_44685);
xor U45770 (N_45770,N_44236,N_42577);
nor U45771 (N_45771,N_43902,N_42823);
or U45772 (N_45772,N_43668,N_44993);
or U45773 (N_45773,N_44881,N_42962);
or U45774 (N_45774,N_44442,N_43439);
nand U45775 (N_45775,N_43542,N_42641);
or U45776 (N_45776,N_44241,N_43391);
and U45777 (N_45777,N_42727,N_44819);
nand U45778 (N_45778,N_44366,N_44003);
and U45779 (N_45779,N_42715,N_42642);
nand U45780 (N_45780,N_44500,N_44797);
or U45781 (N_45781,N_43519,N_44926);
xnor U45782 (N_45782,N_44240,N_42830);
or U45783 (N_45783,N_43786,N_43619);
nor U45784 (N_45784,N_44288,N_44727);
or U45785 (N_45785,N_44493,N_43015);
nor U45786 (N_45786,N_43388,N_44273);
nor U45787 (N_45787,N_44189,N_43339);
nand U45788 (N_45788,N_43770,N_43013);
nand U45789 (N_45789,N_42731,N_44919);
xor U45790 (N_45790,N_43773,N_43713);
xnor U45791 (N_45791,N_43867,N_44418);
nor U45792 (N_45792,N_43712,N_44388);
or U45793 (N_45793,N_43081,N_44832);
xnor U45794 (N_45794,N_42892,N_44686);
and U45795 (N_45795,N_42999,N_44729);
nor U45796 (N_45796,N_44902,N_44907);
nand U45797 (N_45797,N_43557,N_43827);
or U45798 (N_45798,N_44083,N_42679);
or U45799 (N_45799,N_44947,N_44861);
and U45800 (N_45800,N_43284,N_42738);
nand U45801 (N_45801,N_42647,N_43679);
or U45802 (N_45802,N_44984,N_43812);
xor U45803 (N_45803,N_44425,N_43799);
or U45804 (N_45804,N_42900,N_44609);
nor U45805 (N_45805,N_44645,N_44879);
or U45806 (N_45806,N_44798,N_43314);
xnor U45807 (N_45807,N_44169,N_44646);
xnor U45808 (N_45808,N_44937,N_43648);
nor U45809 (N_45809,N_44090,N_43899);
xnor U45810 (N_45810,N_44508,N_43517);
or U45811 (N_45811,N_44708,N_43294);
or U45812 (N_45812,N_44723,N_44120);
nand U45813 (N_45813,N_44760,N_43274);
nor U45814 (N_45814,N_44499,N_42742);
nor U45815 (N_45815,N_44908,N_43611);
nand U45816 (N_45816,N_44562,N_44148);
xor U45817 (N_45817,N_44581,N_43822);
nand U45818 (N_45818,N_44519,N_43001);
or U45819 (N_45819,N_44249,N_43030);
xor U45820 (N_45820,N_43571,N_44002);
xnor U45821 (N_45821,N_44486,N_42553);
nor U45822 (N_45822,N_43839,N_44678);
nand U45823 (N_45823,N_43677,N_44272);
nand U45824 (N_45824,N_43690,N_42926);
and U45825 (N_45825,N_44279,N_44369);
xor U45826 (N_45826,N_43860,N_43962);
xor U45827 (N_45827,N_44699,N_42614);
and U45828 (N_45828,N_44071,N_44941);
xor U45829 (N_45829,N_43149,N_43616);
nor U45830 (N_45830,N_43302,N_44251);
nand U45831 (N_45831,N_44205,N_43894);
xor U45832 (N_45832,N_42904,N_43423);
and U45833 (N_45833,N_43866,N_42791);
nor U45834 (N_45834,N_43177,N_42770);
nor U45835 (N_45835,N_44903,N_42815);
nand U45836 (N_45836,N_44691,N_42945);
nor U45837 (N_45837,N_42645,N_42692);
xor U45838 (N_45838,N_44961,N_42652);
nand U45839 (N_45839,N_42590,N_44644);
nor U45840 (N_45840,N_42516,N_44544);
nor U45841 (N_45841,N_42502,N_44566);
nor U45842 (N_45842,N_43904,N_43375);
nand U45843 (N_45843,N_44038,N_42561);
or U45844 (N_45844,N_42713,N_43363);
nand U45845 (N_45845,N_43283,N_44863);
or U45846 (N_45846,N_42960,N_43319);
and U45847 (N_45847,N_42644,N_43044);
nor U45848 (N_45848,N_43742,N_42576);
or U45849 (N_45849,N_43356,N_42803);
and U45850 (N_45850,N_43190,N_43750);
or U45851 (N_45851,N_42556,N_43440);
nand U45852 (N_45852,N_43330,N_44270);
nand U45853 (N_45853,N_42989,N_43014);
nand U45854 (N_45854,N_43346,N_43788);
or U45855 (N_45855,N_43538,N_44144);
or U45856 (N_45856,N_43277,N_43315);
nor U45857 (N_45857,N_44736,N_44304);
nor U45858 (N_45858,N_43446,N_43272);
and U45859 (N_45859,N_42899,N_43983);
nor U45860 (N_45860,N_43088,N_42902);
or U45861 (N_45861,N_43188,N_44825);
or U45862 (N_45862,N_44000,N_43869);
and U45863 (N_45863,N_44487,N_43746);
and U45864 (N_45864,N_44474,N_42880);
or U45865 (N_45865,N_43925,N_43307);
and U45866 (N_45866,N_43584,N_44483);
and U45867 (N_45867,N_42728,N_44472);
and U45868 (N_45868,N_44026,N_44087);
xnor U45869 (N_45869,N_42846,N_42944);
and U45870 (N_45870,N_43603,N_43681);
and U45871 (N_45871,N_44672,N_42674);
nor U45872 (N_45872,N_42813,N_43594);
nand U45873 (N_45873,N_42982,N_42626);
nor U45874 (N_45874,N_43915,N_44282);
nor U45875 (N_45875,N_43285,N_42983);
nor U45876 (N_45876,N_42690,N_44743);
nor U45877 (N_45877,N_43118,N_42741);
nor U45878 (N_45878,N_43478,N_43718);
or U45879 (N_45879,N_44140,N_44254);
and U45880 (N_45880,N_42695,N_43922);
xnor U45881 (N_45881,N_44584,N_44498);
and U45882 (N_45882,N_42995,N_44136);
nand U45883 (N_45883,N_42864,N_44062);
xnor U45884 (N_45884,N_43022,N_44214);
nand U45885 (N_45885,N_44347,N_44181);
and U45886 (N_45886,N_44420,N_44243);
and U45887 (N_45887,N_43208,N_44454);
and U45888 (N_45888,N_42702,N_44396);
nor U45889 (N_45889,N_42895,N_42788);
nand U45890 (N_45890,N_44385,N_44459);
nor U45891 (N_45891,N_43842,N_43620);
nor U45892 (N_45892,N_43996,N_42752);
nor U45893 (N_45893,N_44490,N_44688);
nand U45894 (N_45894,N_43175,N_42865);
xor U45895 (N_45895,N_44433,N_44079);
nand U45896 (N_45896,N_44110,N_43192);
xnor U45897 (N_45897,N_43136,N_43971);
xnor U45898 (N_45898,N_43705,N_44580);
nand U45899 (N_45899,N_44290,N_44788);
or U45900 (N_45900,N_42822,N_43119);
and U45901 (N_45901,N_43290,N_42840);
nand U45902 (N_45902,N_42792,N_44301);
xor U45903 (N_45903,N_43051,N_44932);
nor U45904 (N_45904,N_42673,N_44269);
nand U45905 (N_45905,N_44426,N_44621);
and U45906 (N_45906,N_43547,N_43831);
nand U45907 (N_45907,N_44592,N_44549);
nand U45908 (N_45908,N_42947,N_43059);
nand U45909 (N_45909,N_44806,N_43870);
or U45910 (N_45910,N_44161,N_42735);
xnor U45911 (N_45911,N_44151,N_43139);
xor U45912 (N_45912,N_44706,N_42756);
and U45913 (N_45913,N_43952,N_42955);
xnor U45914 (N_45914,N_44076,N_44156);
xor U45915 (N_45915,N_44639,N_44681);
nor U45916 (N_45916,N_43752,N_42544);
nand U45917 (N_45917,N_44983,N_44850);
nand U45918 (N_45918,N_43241,N_44444);
nor U45919 (N_45919,N_43355,N_43405);
nor U45920 (N_45920,N_43264,N_43187);
and U45921 (N_45921,N_43636,N_43296);
and U45922 (N_45922,N_43497,N_42730);
nor U45923 (N_45923,N_43340,N_43796);
and U45924 (N_45924,N_44978,N_44721);
or U45925 (N_45925,N_43067,N_44358);
nor U45926 (N_45926,N_42664,N_42776);
and U45927 (N_45927,N_44190,N_43156);
and U45928 (N_45928,N_43678,N_44247);
or U45929 (N_45929,N_43282,N_42986);
or U45930 (N_45930,N_44958,N_44742);
nand U45931 (N_45931,N_44215,N_44818);
xor U45932 (N_45932,N_42838,N_43160);
and U45933 (N_45933,N_44513,N_42509);
nor U45934 (N_45934,N_44911,N_42996);
xor U45935 (N_45935,N_42795,N_44575);
or U45936 (N_45936,N_42571,N_43560);
xnor U45937 (N_45937,N_43515,N_43471);
xnor U45938 (N_45938,N_44731,N_44613);
nand U45939 (N_45939,N_43936,N_43146);
xnor U45940 (N_45940,N_42777,N_42998);
nor U45941 (N_45941,N_43694,N_42547);
nand U45942 (N_45942,N_44754,N_44398);
nand U45943 (N_45943,N_44292,N_44497);
xor U45944 (N_45944,N_43896,N_44328);
nor U45945 (N_45945,N_43753,N_44955);
and U45946 (N_45946,N_43568,N_42757);
and U45947 (N_45947,N_44453,N_44316);
nor U45948 (N_45948,N_44141,N_42584);
nor U45949 (N_45949,N_43900,N_44054);
or U45950 (N_45950,N_44365,N_43089);
nor U45951 (N_45951,N_42686,N_42670);
xnor U45952 (N_45952,N_43421,N_43335);
xor U45953 (N_45953,N_44715,N_42794);
or U45954 (N_45954,N_43270,N_43599);
nor U45955 (N_45955,N_42886,N_44044);
nor U45956 (N_45956,N_43884,N_44032);
xnor U45957 (N_45957,N_44655,N_43267);
xor U45958 (N_45958,N_44327,N_43287);
xor U45959 (N_45959,N_44838,N_43151);
nand U45960 (N_45960,N_44800,N_44452);
xnor U45961 (N_45961,N_44211,N_43903);
and U45962 (N_45962,N_44164,N_43091);
nand U45963 (N_45963,N_42678,N_44170);
xor U45964 (N_45964,N_43551,N_43415);
and U45965 (N_45965,N_43140,N_44733);
and U45966 (N_45966,N_42878,N_44674);
and U45967 (N_45967,N_42548,N_42657);
nand U45968 (N_45968,N_42930,N_42911);
xnor U45969 (N_45969,N_44145,N_44457);
nor U45970 (N_45970,N_44578,N_42891);
nand U45971 (N_45971,N_44424,N_44165);
or U45972 (N_45972,N_44642,N_43237);
and U45973 (N_45973,N_43596,N_44873);
nor U45974 (N_45974,N_43257,N_44515);
nor U45975 (N_45975,N_43946,N_44184);
or U45976 (N_45976,N_43927,N_43545);
nand U45977 (N_45977,N_42761,N_43457);
and U45978 (N_45978,N_44123,N_43787);
nor U45979 (N_45979,N_43877,N_43012);
or U45980 (N_45980,N_42832,N_44154);
nor U45981 (N_45981,N_44606,N_43231);
nand U45982 (N_45982,N_43565,N_43595);
nand U45983 (N_45983,N_44030,N_44890);
nor U45984 (N_45984,N_44231,N_43429);
or U45985 (N_45985,N_42635,N_44451);
and U45986 (N_45986,N_43949,N_44746);
or U45987 (N_45987,N_44810,N_44033);
nand U45988 (N_45988,N_44917,N_44992);
nor U45989 (N_45989,N_44923,N_42987);
and U45990 (N_45990,N_44131,N_43569);
and U45991 (N_45991,N_44198,N_43027);
xnor U45992 (N_45992,N_43583,N_44620);
nor U45993 (N_45993,N_43185,N_43333);
and U45994 (N_45994,N_42810,N_43729);
nor U45995 (N_45995,N_43953,N_42564);
nor U45996 (N_45996,N_43337,N_44255);
xnor U45997 (N_45997,N_42857,N_43486);
nand U45998 (N_45998,N_42661,N_43813);
nor U45999 (N_45999,N_44607,N_43172);
xor U46000 (N_46000,N_44009,N_44333);
xnor U46001 (N_46001,N_44803,N_43326);
and U46002 (N_46002,N_42812,N_44280);
or U46003 (N_46003,N_43836,N_43052);
nor U46004 (N_46004,N_43621,N_44049);
nand U46005 (N_46005,N_44791,N_44095);
nor U46006 (N_46006,N_43777,N_42831);
xnor U46007 (N_46007,N_43931,N_44831);
or U46008 (N_46008,N_42705,N_44552);
or U46009 (N_46009,N_44162,N_43654);
xor U46010 (N_46010,N_42578,N_43308);
or U46011 (N_46011,N_42651,N_43957);
and U46012 (N_46012,N_43226,N_42787);
or U46013 (N_46013,N_44536,N_44612);
and U46014 (N_46014,N_44315,N_43741);
nand U46015 (N_46015,N_44663,N_42940);
xor U46016 (N_46016,N_42834,N_44495);
xor U46017 (N_46017,N_43688,N_43865);
or U46018 (N_46018,N_42915,N_42630);
nand U46019 (N_46019,N_43157,N_44016);
nand U46020 (N_46020,N_44595,N_42771);
nor U46021 (N_46021,N_44375,N_44577);
and U46022 (N_46022,N_44121,N_43567);
or U46023 (N_46023,N_44069,N_44478);
nor U46024 (N_46024,N_44972,N_44436);
nor U46025 (N_46025,N_43135,N_42759);
nand U46026 (N_46026,N_43792,N_44158);
or U46027 (N_46027,N_44485,N_44602);
or U46028 (N_46028,N_43794,N_44718);
nand U46029 (N_46029,N_44571,N_44308);
nor U46030 (N_46030,N_43386,N_43373);
nand U46031 (N_46031,N_43711,N_43066);
nor U46032 (N_46032,N_44350,N_44281);
and U46033 (N_46033,N_42754,N_44233);
and U46034 (N_46034,N_44275,N_44438);
xnor U46035 (N_46035,N_43194,N_44910);
or U46036 (N_46036,N_44590,N_44379);
nor U46037 (N_46037,N_44889,N_43919);
xor U46038 (N_46038,N_44446,N_44017);
xnor U46039 (N_46039,N_42593,N_43697);
nor U46040 (N_46040,N_43747,N_43757);
nand U46041 (N_46041,N_43381,N_43633);
nor U46042 (N_46042,N_42515,N_43404);
nand U46043 (N_46043,N_44950,N_43880);
nor U46044 (N_46044,N_44840,N_42837);
xnor U46045 (N_46045,N_43740,N_43099);
nand U46046 (N_46046,N_42504,N_44268);
xor U46047 (N_46047,N_44367,N_44257);
and U46048 (N_46048,N_43255,N_44467);
or U46049 (N_46049,N_44653,N_43468);
or U46050 (N_46050,N_44119,N_43861);
nor U46051 (N_46051,N_43304,N_43352);
nor U46052 (N_46052,N_42912,N_44785);
nand U46053 (N_46053,N_43180,N_43941);
xor U46054 (N_46054,N_42570,N_42814);
nor U46055 (N_46055,N_44769,N_44475);
and U46056 (N_46056,N_42527,N_42941);
nand U46057 (N_46057,N_44693,N_43618);
nor U46058 (N_46058,N_42672,N_44382);
and U46059 (N_46059,N_44842,N_44377);
nand U46060 (N_46060,N_44392,N_42671);
nand U46061 (N_46061,N_43416,N_44080);
xnor U46062 (N_46062,N_44747,N_42826);
or U46063 (N_46063,N_43835,N_43967);
and U46064 (N_46064,N_43906,N_44755);
nand U46065 (N_46065,N_44407,N_43987);
or U46066 (N_46066,N_43885,N_44072);
nor U46067 (N_46067,N_43841,N_44752);
nand U46068 (N_46068,N_44373,N_42918);
xor U46069 (N_46069,N_43803,N_44938);
and U46070 (N_46070,N_43395,N_43084);
nor U46071 (N_46071,N_44277,N_44885);
nand U46072 (N_46072,N_43643,N_42951);
nand U46073 (N_46073,N_43176,N_44628);
or U46074 (N_46074,N_44226,N_43422);
or U46075 (N_46075,N_44348,N_43000);
nor U46076 (N_46076,N_44775,N_44756);
xnor U46077 (N_46077,N_42512,N_43564);
xnor U46078 (N_46078,N_44772,N_42601);
and U46079 (N_46079,N_44586,N_43685);
xor U46080 (N_46080,N_43459,N_44633);
xnor U46081 (N_46081,N_44948,N_44554);
nor U46082 (N_46082,N_44046,N_44171);
nor U46083 (N_46083,N_43938,N_44833);
xnor U46084 (N_46084,N_43739,N_44773);
or U46085 (N_46085,N_43087,N_44455);
xnor U46086 (N_46086,N_43723,N_43076);
nand U46087 (N_46087,N_42763,N_42968);
and U46088 (N_46088,N_43269,N_42871);
and U46089 (N_46089,N_44228,N_44635);
nand U46090 (N_46090,N_44682,N_44757);
nand U46091 (N_46091,N_44777,N_44589);
nor U46092 (N_46092,N_44130,N_44400);
nand U46093 (N_46093,N_42913,N_43853);
nor U46094 (N_46094,N_44608,N_44680);
and U46095 (N_46095,N_44652,N_43299);
and U46096 (N_46096,N_43249,N_43197);
xnor U46097 (N_46097,N_43400,N_42935);
or U46098 (N_46098,N_44463,N_43124);
nand U46099 (N_46099,N_44488,N_43774);
xnor U46100 (N_46100,N_42733,N_42963);
nand U46101 (N_46101,N_44627,N_43514);
and U46102 (N_46102,N_42710,N_44225);
xor U46103 (N_46103,N_44532,N_43273);
xnor U46104 (N_46104,N_42887,N_43943);
or U46105 (N_46105,N_42950,N_43288);
or U46106 (N_46106,N_44516,N_44018);
nor U46107 (N_46107,N_44600,N_44362);
xnor U46108 (N_46108,N_44440,N_43444);
and U46109 (N_46109,N_43976,N_43019);
and U46110 (N_46110,N_44476,N_42868);
and U46111 (N_46111,N_42906,N_44563);
or U46112 (N_46112,N_43343,N_44019);
nand U46113 (N_46113,N_42964,N_43469);
and U46114 (N_46114,N_44263,N_43982);
xor U46115 (N_46115,N_42696,N_44913);
or U46116 (N_46116,N_44705,N_43531);
nand U46117 (N_46117,N_43895,N_43158);
nor U46118 (N_46118,N_43456,N_43133);
nor U46119 (N_46119,N_42917,N_44321);
xnor U46120 (N_46120,N_43675,N_44450);
xnor U46121 (N_46121,N_43888,N_43435);
xnor U46122 (N_46122,N_42607,N_43201);
xnor U46123 (N_46123,N_44204,N_44051);
xnor U46124 (N_46124,N_44462,N_42562);
or U46125 (N_46125,N_43144,N_44841);
xnor U46126 (N_46126,N_44795,N_44616);
or U46127 (N_46127,N_43907,N_42949);
or U46128 (N_46128,N_43646,N_43892);
and U46129 (N_46129,N_44660,N_43258);
or U46130 (N_46130,N_42500,N_42636);
nand U46131 (N_46131,N_43024,N_42758);
nor U46132 (N_46132,N_42542,N_44175);
nor U46133 (N_46133,N_42649,N_43553);
and U46134 (N_46134,N_44266,N_43104);
nor U46135 (N_46135,N_44712,N_42513);
xor U46136 (N_46136,N_43503,N_42568);
nor U46137 (N_46137,N_44748,N_43684);
nor U46138 (N_46138,N_44041,N_44817);
nor U46139 (N_46139,N_44364,N_44784);
and U46140 (N_46140,N_43520,N_43537);
and U46141 (N_46141,N_43736,N_43833);
and U46142 (N_46142,N_44596,N_43298);
nor U46143 (N_46143,N_42612,N_42977);
nor U46144 (N_46144,N_44036,N_44647);
xor U46145 (N_46145,N_43574,N_44209);
nor U46146 (N_46146,N_42517,N_43525);
and U46147 (N_46147,N_43464,N_44977);
nor U46148 (N_46148,N_43782,N_44931);
nand U46149 (N_46149,N_44354,N_44235);
xor U46150 (N_46150,N_43798,N_44887);
and U46151 (N_46151,N_44183,N_43385);
and U46152 (N_46152,N_43134,N_43687);
and U46153 (N_46153,N_44640,N_44720);
nand U46154 (N_46154,N_43891,N_43504);
or U46155 (N_46155,N_43625,N_44550);
xnor U46156 (N_46156,N_43748,N_44927);
and U46157 (N_46157,N_43691,N_43476);
or U46158 (N_46158,N_42976,N_43610);
or U46159 (N_46159,N_43830,N_44128);
and U46160 (N_46160,N_44974,N_44914);
and U46161 (N_46161,N_43669,N_44849);
nor U46162 (N_46162,N_43029,N_43702);
and U46163 (N_46163,N_42772,N_43154);
nand U46164 (N_46164,N_43828,N_44107);
or U46165 (N_46165,N_43331,N_43876);
or U46166 (N_46166,N_44988,N_42712);
and U46167 (N_46167,N_42914,N_43394);
or U46168 (N_46168,N_44432,N_44443);
xnor U46169 (N_46169,N_42646,N_43460);
nor U46170 (N_46170,N_42522,N_42861);
and U46171 (N_46171,N_43623,N_42997);
and U46172 (N_46172,N_44219,N_43857);
or U46173 (N_46173,N_44224,N_44302);
nor U46174 (N_46174,N_43490,N_44193);
or U46175 (N_46175,N_43170,N_43879);
or U46176 (N_46176,N_43759,N_43482);
xnor U46177 (N_46177,N_43913,N_43039);
nand U46178 (N_46178,N_42925,N_44339);
nor U46179 (N_46179,N_43297,N_43129);
nand U46180 (N_46180,N_42634,N_43082);
and U46181 (N_46181,N_42981,N_44793);
xor U46182 (N_46182,N_44441,N_44390);
xor U46183 (N_46183,N_44744,N_44541);
or U46184 (N_46184,N_43349,N_44413);
xnor U46185 (N_46185,N_43850,N_44766);
nor U46186 (N_46186,N_44695,N_44583);
nor U46187 (N_46187,N_43184,N_43849);
or U46188 (N_46188,N_44173,N_44063);
and U46189 (N_46189,N_44936,N_43017);
and U46190 (N_46190,N_42697,N_44971);
or U46191 (N_46191,N_43152,N_44834);
or U46192 (N_46192,N_44374,N_44031);
nor U46193 (N_46193,N_44982,N_44494);
nand U46194 (N_46194,N_42706,N_43371);
nor U46195 (N_46195,N_44997,N_43131);
and U46196 (N_46196,N_42558,N_44428);
nor U46197 (N_46197,N_44694,N_44234);
xnor U46198 (N_46198,N_43125,N_44299);
nand U46199 (N_46199,N_44741,N_43693);
and U46200 (N_46200,N_42681,N_44523);
or U46201 (N_46201,N_43532,N_43530);
and U46202 (N_46202,N_42639,N_42653);
and U46203 (N_46203,N_42973,N_44264);
nor U46204 (N_46204,N_43582,N_44666);
xnor U46205 (N_46205,N_44111,N_44891);
or U46206 (N_46206,N_43924,N_42665);
xor U46207 (N_46207,N_43414,N_43109);
nand U46208 (N_46208,N_44359,N_44309);
or U46209 (N_46209,N_44614,N_44469);
xor U46210 (N_46210,N_43263,N_43075);
xnor U46211 (N_46211,N_44039,N_43649);
nand U46212 (N_46212,N_43826,N_44726);
nor U46213 (N_46213,N_43703,N_43658);
nand U46214 (N_46214,N_43003,N_43823);
or U46215 (N_46215,N_42550,N_42793);
and U46216 (N_46216,N_43011,N_44484);
or U46217 (N_46217,N_43321,N_44537);
nor U46218 (N_46218,N_44216,N_44195);
nor U46219 (N_46219,N_44893,N_43061);
nor U46220 (N_46220,N_44372,N_43725);
xnor U46221 (N_46221,N_44191,N_44857);
xnor U46222 (N_46222,N_43413,N_44980);
xor U46223 (N_46223,N_44687,N_44543);
nor U46224 (N_46224,N_43581,N_44326);
nor U46225 (N_46225,N_43978,N_43494);
nand U46226 (N_46226,N_43682,N_44996);
and U46227 (N_46227,N_42937,N_44244);
xor U46228 (N_46228,N_42531,N_44967);
or U46229 (N_46229,N_44511,N_43848);
and U46230 (N_46230,N_44208,N_43522);
and U46231 (N_46231,N_42535,N_43311);
nor U46232 (N_46232,N_44334,N_43960);
nand U46233 (N_46233,N_44951,N_44560);
or U46234 (N_46234,N_43529,N_43709);
nor U46235 (N_46235,N_44458,N_43968);
nor U46236 (N_46236,N_44115,N_44423);
nand U46237 (N_46237,N_43211,N_44601);
nand U46238 (N_46238,N_42569,N_42740);
and U46239 (N_46239,N_43463,N_44995);
nand U46240 (N_46240,N_44501,N_44994);
nor U46241 (N_46241,N_42863,N_43301);
xnor U46242 (N_46242,N_44221,N_43096);
and U46243 (N_46243,N_43704,N_43224);
or U46244 (N_46244,N_44070,N_44510);
nor U46245 (N_46245,N_43732,N_43419);
xor U46246 (N_46246,N_43923,N_44724);
or U46247 (N_46247,N_43602,N_43470);
and U46248 (N_46248,N_43507,N_44001);
nor U46249 (N_46249,N_43393,N_44310);
xor U46250 (N_46250,N_43272,N_43241);
nor U46251 (N_46251,N_43450,N_42746);
xnor U46252 (N_46252,N_42766,N_43819);
nor U46253 (N_46253,N_43789,N_44035);
nand U46254 (N_46254,N_43962,N_43358);
and U46255 (N_46255,N_44887,N_44452);
nor U46256 (N_46256,N_43296,N_42599);
and U46257 (N_46257,N_44699,N_42779);
or U46258 (N_46258,N_43295,N_43230);
xnor U46259 (N_46259,N_42542,N_42963);
and U46260 (N_46260,N_44250,N_42826);
nand U46261 (N_46261,N_44426,N_42621);
or U46262 (N_46262,N_44363,N_43139);
xnor U46263 (N_46263,N_42761,N_42776);
or U46264 (N_46264,N_43494,N_44829);
nor U46265 (N_46265,N_42536,N_44442);
and U46266 (N_46266,N_43451,N_43165);
nor U46267 (N_46267,N_43514,N_43231);
nor U46268 (N_46268,N_43157,N_43282);
nor U46269 (N_46269,N_42505,N_44574);
nor U46270 (N_46270,N_43147,N_44030);
and U46271 (N_46271,N_43774,N_44838);
xnor U46272 (N_46272,N_43490,N_44459);
and U46273 (N_46273,N_42569,N_43503);
nor U46274 (N_46274,N_42608,N_44820);
or U46275 (N_46275,N_43188,N_44321);
xor U46276 (N_46276,N_43897,N_42970);
or U46277 (N_46277,N_42885,N_44290);
xor U46278 (N_46278,N_44833,N_43029);
or U46279 (N_46279,N_44581,N_43631);
xnor U46280 (N_46280,N_43704,N_44575);
or U46281 (N_46281,N_44908,N_43428);
nand U46282 (N_46282,N_44307,N_43820);
and U46283 (N_46283,N_43123,N_42596);
and U46284 (N_46284,N_43722,N_43356);
and U46285 (N_46285,N_44457,N_43664);
nor U46286 (N_46286,N_44242,N_44664);
xnor U46287 (N_46287,N_43675,N_44846);
nor U46288 (N_46288,N_42593,N_44520);
nor U46289 (N_46289,N_43803,N_44996);
nor U46290 (N_46290,N_43074,N_44590);
xnor U46291 (N_46291,N_43566,N_43467);
or U46292 (N_46292,N_43702,N_44116);
nand U46293 (N_46293,N_43248,N_43246);
xor U46294 (N_46294,N_43706,N_44283);
nor U46295 (N_46295,N_43913,N_42914);
and U46296 (N_46296,N_44530,N_44833);
nand U46297 (N_46297,N_44520,N_44060);
nor U46298 (N_46298,N_43852,N_44845);
or U46299 (N_46299,N_44526,N_44995);
nor U46300 (N_46300,N_44886,N_44941);
xnor U46301 (N_46301,N_43860,N_42851);
xor U46302 (N_46302,N_43059,N_43406);
nand U46303 (N_46303,N_44720,N_42511);
or U46304 (N_46304,N_43908,N_43506);
and U46305 (N_46305,N_44966,N_42560);
nand U46306 (N_46306,N_43450,N_42817);
xnor U46307 (N_46307,N_43916,N_44537);
xnor U46308 (N_46308,N_43367,N_43003);
or U46309 (N_46309,N_44382,N_43686);
and U46310 (N_46310,N_43530,N_44530);
and U46311 (N_46311,N_43941,N_44676);
nor U46312 (N_46312,N_43659,N_44417);
and U46313 (N_46313,N_42590,N_44390);
nor U46314 (N_46314,N_43522,N_42828);
xnor U46315 (N_46315,N_42766,N_43234);
xnor U46316 (N_46316,N_44515,N_43293);
nor U46317 (N_46317,N_44637,N_44162);
or U46318 (N_46318,N_43379,N_43426);
or U46319 (N_46319,N_44140,N_43810);
xor U46320 (N_46320,N_44250,N_43831);
or U46321 (N_46321,N_43217,N_44620);
xor U46322 (N_46322,N_43975,N_44313);
nand U46323 (N_46323,N_43891,N_43722);
xnor U46324 (N_46324,N_43474,N_43750);
and U46325 (N_46325,N_42788,N_43544);
nor U46326 (N_46326,N_42539,N_43774);
nand U46327 (N_46327,N_43914,N_43691);
xor U46328 (N_46328,N_44263,N_44107);
xnor U46329 (N_46329,N_44958,N_42940);
nand U46330 (N_46330,N_42657,N_43418);
and U46331 (N_46331,N_42781,N_44626);
nand U46332 (N_46332,N_43134,N_44691);
and U46333 (N_46333,N_43669,N_43676);
and U46334 (N_46334,N_44414,N_43119);
nor U46335 (N_46335,N_42534,N_44397);
xor U46336 (N_46336,N_43990,N_43120);
and U46337 (N_46337,N_44696,N_44994);
nor U46338 (N_46338,N_43552,N_44834);
or U46339 (N_46339,N_44416,N_43438);
nor U46340 (N_46340,N_43157,N_44950);
nor U46341 (N_46341,N_43466,N_43814);
and U46342 (N_46342,N_44155,N_44846);
nor U46343 (N_46343,N_42655,N_43157);
xor U46344 (N_46344,N_43664,N_43169);
nand U46345 (N_46345,N_44540,N_42623);
nor U46346 (N_46346,N_42849,N_44738);
nor U46347 (N_46347,N_43828,N_44927);
nor U46348 (N_46348,N_42604,N_44652);
xnor U46349 (N_46349,N_42914,N_44046);
nor U46350 (N_46350,N_42620,N_43719);
nand U46351 (N_46351,N_42509,N_43251);
and U46352 (N_46352,N_44951,N_43429);
and U46353 (N_46353,N_44590,N_44346);
nor U46354 (N_46354,N_43700,N_43984);
nor U46355 (N_46355,N_42883,N_44392);
and U46356 (N_46356,N_44020,N_42554);
or U46357 (N_46357,N_44120,N_43317);
xnor U46358 (N_46358,N_42702,N_43619);
xnor U46359 (N_46359,N_42573,N_44624);
xnor U46360 (N_46360,N_44688,N_43332);
and U46361 (N_46361,N_44823,N_44155);
nor U46362 (N_46362,N_44277,N_43904);
and U46363 (N_46363,N_43117,N_43743);
xnor U46364 (N_46364,N_44068,N_43624);
nand U46365 (N_46365,N_44302,N_44880);
nor U46366 (N_46366,N_43352,N_43184);
xnor U46367 (N_46367,N_44232,N_43279);
nand U46368 (N_46368,N_44862,N_43432);
or U46369 (N_46369,N_44409,N_42850);
or U46370 (N_46370,N_43601,N_44742);
nand U46371 (N_46371,N_44714,N_44072);
nand U46372 (N_46372,N_43085,N_43292);
xor U46373 (N_46373,N_42957,N_44134);
and U46374 (N_46374,N_42730,N_44245);
nand U46375 (N_46375,N_43684,N_44800);
nor U46376 (N_46376,N_43033,N_43979);
nor U46377 (N_46377,N_42999,N_42685);
and U46378 (N_46378,N_42679,N_42639);
nor U46379 (N_46379,N_44198,N_42508);
xnor U46380 (N_46380,N_43163,N_44136);
and U46381 (N_46381,N_43222,N_42833);
xor U46382 (N_46382,N_44107,N_43407);
xor U46383 (N_46383,N_44238,N_43081);
xor U46384 (N_46384,N_44405,N_42538);
nand U46385 (N_46385,N_42597,N_44570);
xor U46386 (N_46386,N_44581,N_44784);
xor U46387 (N_46387,N_42889,N_44617);
nor U46388 (N_46388,N_44814,N_43311);
nand U46389 (N_46389,N_42967,N_43260);
and U46390 (N_46390,N_44044,N_43902);
or U46391 (N_46391,N_43498,N_44853);
xnor U46392 (N_46392,N_44684,N_44470);
or U46393 (N_46393,N_43655,N_44859);
xnor U46394 (N_46394,N_43005,N_43214);
and U46395 (N_46395,N_43661,N_43667);
xnor U46396 (N_46396,N_44080,N_43613);
and U46397 (N_46397,N_43517,N_44940);
nor U46398 (N_46398,N_44017,N_44948);
or U46399 (N_46399,N_44667,N_43593);
nand U46400 (N_46400,N_43524,N_43926);
and U46401 (N_46401,N_42627,N_44566);
and U46402 (N_46402,N_42702,N_42996);
xor U46403 (N_46403,N_44770,N_42878);
and U46404 (N_46404,N_44630,N_44297);
nand U46405 (N_46405,N_43563,N_42513);
or U46406 (N_46406,N_43669,N_44614);
nor U46407 (N_46407,N_44589,N_42692);
or U46408 (N_46408,N_44067,N_43100);
nor U46409 (N_46409,N_42688,N_44593);
xnor U46410 (N_46410,N_43331,N_44695);
and U46411 (N_46411,N_43665,N_43422);
and U46412 (N_46412,N_43917,N_43020);
nor U46413 (N_46413,N_44302,N_44757);
or U46414 (N_46414,N_43972,N_44462);
or U46415 (N_46415,N_44803,N_42955);
xnor U46416 (N_46416,N_43877,N_44508);
or U46417 (N_46417,N_44224,N_44195);
nand U46418 (N_46418,N_43419,N_43170);
and U46419 (N_46419,N_43103,N_43446);
nand U46420 (N_46420,N_44744,N_43214);
or U46421 (N_46421,N_44495,N_44601);
nand U46422 (N_46422,N_44356,N_44667);
nor U46423 (N_46423,N_42765,N_42655);
nand U46424 (N_46424,N_43151,N_43206);
xnor U46425 (N_46425,N_43170,N_43678);
nand U46426 (N_46426,N_44842,N_44008);
xor U46427 (N_46427,N_42884,N_44507);
and U46428 (N_46428,N_42632,N_44129);
or U46429 (N_46429,N_44621,N_43681);
xnor U46430 (N_46430,N_43050,N_42532);
nand U46431 (N_46431,N_43957,N_44407);
xor U46432 (N_46432,N_42918,N_43973);
nor U46433 (N_46433,N_43767,N_44102);
and U46434 (N_46434,N_44721,N_43128);
xor U46435 (N_46435,N_42592,N_44282);
or U46436 (N_46436,N_44371,N_44019);
xor U46437 (N_46437,N_44379,N_44621);
or U46438 (N_46438,N_44005,N_44730);
nand U46439 (N_46439,N_42507,N_43615);
and U46440 (N_46440,N_44543,N_43964);
xor U46441 (N_46441,N_43241,N_43059);
or U46442 (N_46442,N_42819,N_42560);
and U46443 (N_46443,N_44196,N_44931);
nand U46444 (N_46444,N_44356,N_44270);
nor U46445 (N_46445,N_43223,N_43375);
nor U46446 (N_46446,N_44694,N_44912);
or U46447 (N_46447,N_44126,N_43785);
nor U46448 (N_46448,N_43343,N_44017);
nand U46449 (N_46449,N_43765,N_42572);
and U46450 (N_46450,N_43128,N_44196);
xor U46451 (N_46451,N_44031,N_44924);
and U46452 (N_46452,N_44004,N_43167);
nand U46453 (N_46453,N_43546,N_43623);
nor U46454 (N_46454,N_44996,N_43318);
nor U46455 (N_46455,N_44963,N_43776);
or U46456 (N_46456,N_43944,N_42554);
xnor U46457 (N_46457,N_44716,N_44721);
nand U46458 (N_46458,N_42661,N_44196);
and U46459 (N_46459,N_44675,N_44358);
nand U46460 (N_46460,N_42566,N_43939);
or U46461 (N_46461,N_44478,N_44397);
nand U46462 (N_46462,N_44669,N_44615);
or U46463 (N_46463,N_44125,N_43272);
or U46464 (N_46464,N_42864,N_43807);
or U46465 (N_46465,N_43719,N_43850);
and U46466 (N_46466,N_44053,N_43898);
xor U46467 (N_46467,N_43858,N_44931);
and U46468 (N_46468,N_42573,N_44390);
xor U46469 (N_46469,N_43156,N_44853);
nor U46470 (N_46470,N_44313,N_42681);
nor U46471 (N_46471,N_43704,N_44662);
and U46472 (N_46472,N_43963,N_43253);
or U46473 (N_46473,N_43645,N_43507);
nor U46474 (N_46474,N_44282,N_42624);
or U46475 (N_46475,N_43679,N_44637);
nand U46476 (N_46476,N_44456,N_44846);
or U46477 (N_46477,N_42951,N_42585);
or U46478 (N_46478,N_43753,N_44178);
xor U46479 (N_46479,N_44077,N_44162);
nor U46480 (N_46480,N_44625,N_42693);
or U46481 (N_46481,N_42955,N_43006);
nand U46482 (N_46482,N_43508,N_44406);
xnor U46483 (N_46483,N_44535,N_44544);
nand U46484 (N_46484,N_42756,N_42545);
and U46485 (N_46485,N_42955,N_43788);
and U46486 (N_46486,N_43817,N_44558);
nor U46487 (N_46487,N_43328,N_43076);
nand U46488 (N_46488,N_42658,N_42659);
and U46489 (N_46489,N_43019,N_43708);
nor U46490 (N_46490,N_42561,N_43588);
or U46491 (N_46491,N_43118,N_43863);
or U46492 (N_46492,N_43594,N_42978);
nor U46493 (N_46493,N_42781,N_43179);
and U46494 (N_46494,N_43003,N_43918);
nor U46495 (N_46495,N_44462,N_44263);
nor U46496 (N_46496,N_43807,N_43928);
or U46497 (N_46497,N_43887,N_44222);
xor U46498 (N_46498,N_43324,N_43596);
nand U46499 (N_46499,N_43882,N_42973);
nand U46500 (N_46500,N_42957,N_43593);
or U46501 (N_46501,N_43610,N_42587);
and U46502 (N_46502,N_43796,N_42890);
and U46503 (N_46503,N_43177,N_42902);
or U46504 (N_46504,N_44946,N_44298);
xor U46505 (N_46505,N_42807,N_43632);
and U46506 (N_46506,N_43107,N_42588);
nand U46507 (N_46507,N_44180,N_43622);
or U46508 (N_46508,N_42555,N_42693);
xor U46509 (N_46509,N_43785,N_44580);
and U46510 (N_46510,N_43798,N_43434);
xnor U46511 (N_46511,N_44361,N_43655);
xor U46512 (N_46512,N_43168,N_43709);
nor U46513 (N_46513,N_44367,N_44485);
nor U46514 (N_46514,N_43315,N_43938);
xnor U46515 (N_46515,N_43179,N_44862);
xor U46516 (N_46516,N_42510,N_44502);
nand U46517 (N_46517,N_43866,N_44018);
or U46518 (N_46518,N_42733,N_44180);
xor U46519 (N_46519,N_44323,N_42827);
xor U46520 (N_46520,N_43066,N_42775);
nand U46521 (N_46521,N_42556,N_43472);
or U46522 (N_46522,N_44993,N_43748);
and U46523 (N_46523,N_43827,N_43697);
nand U46524 (N_46524,N_43963,N_44812);
nand U46525 (N_46525,N_42571,N_43632);
xnor U46526 (N_46526,N_44467,N_44804);
nand U46527 (N_46527,N_44919,N_42789);
nand U46528 (N_46528,N_44221,N_42599);
and U46529 (N_46529,N_42812,N_44777);
nand U46530 (N_46530,N_43102,N_42992);
and U46531 (N_46531,N_43298,N_44086);
and U46532 (N_46532,N_42840,N_43425);
or U46533 (N_46533,N_44273,N_43654);
nand U46534 (N_46534,N_44748,N_42770);
nor U46535 (N_46535,N_43687,N_44566);
xor U46536 (N_46536,N_44750,N_42809);
xnor U46537 (N_46537,N_42748,N_44645);
nor U46538 (N_46538,N_43770,N_44021);
and U46539 (N_46539,N_42700,N_43437);
and U46540 (N_46540,N_42553,N_42755);
nand U46541 (N_46541,N_42890,N_43312);
nor U46542 (N_46542,N_44494,N_44904);
xnor U46543 (N_46543,N_44914,N_44367);
nand U46544 (N_46544,N_42626,N_43464);
nor U46545 (N_46545,N_44059,N_43609);
xor U46546 (N_46546,N_43122,N_43041);
xor U46547 (N_46547,N_43450,N_44047);
xor U46548 (N_46548,N_44683,N_43606);
or U46549 (N_46549,N_42704,N_42530);
xor U46550 (N_46550,N_43429,N_44430);
or U46551 (N_46551,N_42829,N_44460);
and U46552 (N_46552,N_44255,N_43061);
or U46553 (N_46553,N_43503,N_43658);
and U46554 (N_46554,N_43900,N_44339);
nand U46555 (N_46555,N_42748,N_43653);
and U46556 (N_46556,N_42954,N_44652);
nand U46557 (N_46557,N_43185,N_43694);
xnor U46558 (N_46558,N_43635,N_43655);
xnor U46559 (N_46559,N_43047,N_44783);
nor U46560 (N_46560,N_44943,N_43604);
xor U46561 (N_46561,N_44158,N_43250);
nor U46562 (N_46562,N_42702,N_44108);
xor U46563 (N_46563,N_43611,N_44127);
nor U46564 (N_46564,N_43099,N_44800);
and U46565 (N_46565,N_43932,N_42644);
and U46566 (N_46566,N_44259,N_42624);
nor U46567 (N_46567,N_44605,N_44657);
nand U46568 (N_46568,N_43583,N_42899);
nand U46569 (N_46569,N_44753,N_42763);
and U46570 (N_46570,N_43636,N_42984);
and U46571 (N_46571,N_44898,N_43127);
xor U46572 (N_46572,N_44817,N_43870);
and U46573 (N_46573,N_44884,N_42542);
and U46574 (N_46574,N_44559,N_44412);
xnor U46575 (N_46575,N_42644,N_43278);
nand U46576 (N_46576,N_44318,N_44356);
nand U46577 (N_46577,N_43512,N_43246);
and U46578 (N_46578,N_42502,N_44043);
or U46579 (N_46579,N_44710,N_44450);
nand U46580 (N_46580,N_43175,N_44855);
xor U46581 (N_46581,N_43380,N_43090);
nor U46582 (N_46582,N_42866,N_43206);
nor U46583 (N_46583,N_44698,N_44322);
or U46584 (N_46584,N_42907,N_44823);
or U46585 (N_46585,N_43969,N_43931);
and U46586 (N_46586,N_42997,N_44578);
and U46587 (N_46587,N_44743,N_43099);
and U46588 (N_46588,N_44326,N_42948);
nand U46589 (N_46589,N_44671,N_43697);
and U46590 (N_46590,N_43163,N_42807);
nand U46591 (N_46591,N_43325,N_44624);
and U46592 (N_46592,N_42974,N_42811);
nor U46593 (N_46593,N_43777,N_43299);
nand U46594 (N_46594,N_43983,N_42744);
and U46595 (N_46595,N_44634,N_44877);
nor U46596 (N_46596,N_43810,N_42836);
and U46597 (N_46597,N_43090,N_44689);
or U46598 (N_46598,N_44916,N_42743);
xor U46599 (N_46599,N_43528,N_43727);
xnor U46600 (N_46600,N_42624,N_44344);
and U46601 (N_46601,N_44404,N_43902);
xnor U46602 (N_46602,N_42678,N_43433);
nand U46603 (N_46603,N_44731,N_44300);
or U46604 (N_46604,N_44182,N_42710);
nand U46605 (N_46605,N_44086,N_43366);
and U46606 (N_46606,N_44712,N_43629);
and U46607 (N_46607,N_44719,N_44437);
or U46608 (N_46608,N_43096,N_44100);
nand U46609 (N_46609,N_43094,N_44743);
or U46610 (N_46610,N_44944,N_43075);
nand U46611 (N_46611,N_43318,N_43544);
and U46612 (N_46612,N_44892,N_43650);
and U46613 (N_46613,N_43641,N_44349);
nor U46614 (N_46614,N_42592,N_43395);
or U46615 (N_46615,N_42723,N_44943);
nor U46616 (N_46616,N_43314,N_42935);
or U46617 (N_46617,N_44459,N_43818);
xor U46618 (N_46618,N_43076,N_44947);
nand U46619 (N_46619,N_43063,N_44827);
nor U46620 (N_46620,N_42979,N_44657);
or U46621 (N_46621,N_43521,N_44431);
xor U46622 (N_46622,N_42708,N_43655);
nand U46623 (N_46623,N_44944,N_42518);
or U46624 (N_46624,N_43260,N_42975);
or U46625 (N_46625,N_43762,N_44454);
nor U46626 (N_46626,N_43877,N_42817);
or U46627 (N_46627,N_43890,N_42914);
nand U46628 (N_46628,N_43618,N_42911);
xor U46629 (N_46629,N_44516,N_42737);
nor U46630 (N_46630,N_44760,N_43748);
xnor U46631 (N_46631,N_42548,N_44601);
nand U46632 (N_46632,N_43875,N_43937);
xnor U46633 (N_46633,N_43259,N_43877);
or U46634 (N_46634,N_43914,N_44330);
and U46635 (N_46635,N_43417,N_44644);
xnor U46636 (N_46636,N_44056,N_42979);
or U46637 (N_46637,N_44053,N_43013);
or U46638 (N_46638,N_42958,N_43458);
nor U46639 (N_46639,N_44668,N_42709);
or U46640 (N_46640,N_44835,N_43211);
xnor U46641 (N_46641,N_44259,N_44919);
nand U46642 (N_46642,N_42959,N_42524);
and U46643 (N_46643,N_42888,N_44192);
nand U46644 (N_46644,N_44807,N_44484);
and U46645 (N_46645,N_42958,N_43599);
or U46646 (N_46646,N_43478,N_44277);
nor U46647 (N_46647,N_42748,N_42674);
or U46648 (N_46648,N_42795,N_44670);
nor U46649 (N_46649,N_43499,N_44577);
xnor U46650 (N_46650,N_43425,N_42769);
and U46651 (N_46651,N_44399,N_44450);
nand U46652 (N_46652,N_44987,N_44962);
xnor U46653 (N_46653,N_42731,N_44076);
or U46654 (N_46654,N_44916,N_43591);
nand U46655 (N_46655,N_44878,N_44970);
nor U46656 (N_46656,N_42823,N_43552);
nor U46657 (N_46657,N_43373,N_44904);
or U46658 (N_46658,N_43253,N_42623);
xor U46659 (N_46659,N_42827,N_43370);
nand U46660 (N_46660,N_42811,N_43182);
nor U46661 (N_46661,N_44591,N_43836);
xnor U46662 (N_46662,N_43970,N_44274);
xnor U46663 (N_46663,N_42808,N_43724);
and U46664 (N_46664,N_43583,N_44679);
xor U46665 (N_46665,N_44364,N_44397);
nand U46666 (N_46666,N_44123,N_42832);
and U46667 (N_46667,N_43280,N_42868);
or U46668 (N_46668,N_43115,N_43119);
nand U46669 (N_46669,N_44785,N_43247);
nand U46670 (N_46670,N_43162,N_43122);
xor U46671 (N_46671,N_44961,N_43803);
nor U46672 (N_46672,N_43543,N_43051);
or U46673 (N_46673,N_43769,N_44803);
nand U46674 (N_46674,N_43902,N_43333);
or U46675 (N_46675,N_43110,N_44031);
nor U46676 (N_46676,N_44011,N_43286);
xnor U46677 (N_46677,N_44441,N_44672);
nor U46678 (N_46678,N_44668,N_43115);
or U46679 (N_46679,N_43368,N_42572);
nand U46680 (N_46680,N_43670,N_42953);
and U46681 (N_46681,N_44226,N_43821);
nor U46682 (N_46682,N_42654,N_43557);
nand U46683 (N_46683,N_43291,N_43584);
xnor U46684 (N_46684,N_44864,N_43289);
nor U46685 (N_46685,N_43317,N_42934);
xor U46686 (N_46686,N_42629,N_43102);
nor U46687 (N_46687,N_44464,N_44802);
or U46688 (N_46688,N_44396,N_43245);
or U46689 (N_46689,N_43481,N_44860);
nand U46690 (N_46690,N_44326,N_44699);
xor U46691 (N_46691,N_43404,N_42615);
nand U46692 (N_46692,N_44801,N_44877);
nand U46693 (N_46693,N_43860,N_43768);
or U46694 (N_46694,N_43719,N_44344);
nand U46695 (N_46695,N_44539,N_42657);
nand U46696 (N_46696,N_42698,N_44132);
nand U46697 (N_46697,N_43325,N_44487);
nor U46698 (N_46698,N_44112,N_44973);
nor U46699 (N_46699,N_44781,N_43384);
xnor U46700 (N_46700,N_43864,N_42609);
and U46701 (N_46701,N_44163,N_43485);
nor U46702 (N_46702,N_43960,N_44342);
xnor U46703 (N_46703,N_42629,N_43273);
and U46704 (N_46704,N_43132,N_43382);
or U46705 (N_46705,N_44426,N_44644);
and U46706 (N_46706,N_42849,N_44281);
xor U46707 (N_46707,N_44594,N_44531);
nand U46708 (N_46708,N_44147,N_42748);
xor U46709 (N_46709,N_43013,N_43368);
and U46710 (N_46710,N_43538,N_44473);
or U46711 (N_46711,N_43413,N_44829);
xor U46712 (N_46712,N_43569,N_43438);
nand U46713 (N_46713,N_43631,N_43107);
nand U46714 (N_46714,N_43508,N_44790);
nand U46715 (N_46715,N_44421,N_43380);
or U46716 (N_46716,N_43330,N_44623);
nor U46717 (N_46717,N_43186,N_42697);
xor U46718 (N_46718,N_42653,N_44626);
nand U46719 (N_46719,N_44607,N_43494);
nor U46720 (N_46720,N_43465,N_43374);
and U46721 (N_46721,N_43769,N_43485);
nor U46722 (N_46722,N_42816,N_43215);
nand U46723 (N_46723,N_43520,N_43782);
nor U46724 (N_46724,N_43503,N_44449);
and U46725 (N_46725,N_43816,N_44678);
nand U46726 (N_46726,N_44059,N_43563);
nor U46727 (N_46727,N_44606,N_43800);
xor U46728 (N_46728,N_44014,N_43037);
nor U46729 (N_46729,N_42699,N_44020);
and U46730 (N_46730,N_43854,N_44712);
xor U46731 (N_46731,N_43436,N_44218);
or U46732 (N_46732,N_43932,N_43515);
nor U46733 (N_46733,N_44919,N_44758);
nand U46734 (N_46734,N_44758,N_44356);
nand U46735 (N_46735,N_44841,N_42692);
and U46736 (N_46736,N_44366,N_43249);
xor U46737 (N_46737,N_43860,N_44261);
nand U46738 (N_46738,N_44779,N_42942);
nand U46739 (N_46739,N_43338,N_44380);
and U46740 (N_46740,N_42532,N_44260);
nand U46741 (N_46741,N_44880,N_44676);
xor U46742 (N_46742,N_42784,N_43173);
and U46743 (N_46743,N_42986,N_43710);
and U46744 (N_46744,N_43400,N_43615);
nand U46745 (N_46745,N_43194,N_42530);
xnor U46746 (N_46746,N_44246,N_44252);
xor U46747 (N_46747,N_43833,N_44215);
nor U46748 (N_46748,N_43694,N_44692);
xor U46749 (N_46749,N_42702,N_44289);
nand U46750 (N_46750,N_44125,N_44184);
and U46751 (N_46751,N_42661,N_43338);
nand U46752 (N_46752,N_44560,N_43076);
nand U46753 (N_46753,N_42715,N_43914);
nor U46754 (N_46754,N_44846,N_43360);
xnor U46755 (N_46755,N_43135,N_43158);
and U46756 (N_46756,N_42618,N_43713);
nor U46757 (N_46757,N_44665,N_42813);
nor U46758 (N_46758,N_43215,N_43575);
nor U46759 (N_46759,N_44549,N_43066);
or U46760 (N_46760,N_43363,N_43734);
and U46761 (N_46761,N_44018,N_42915);
nand U46762 (N_46762,N_43337,N_44235);
and U46763 (N_46763,N_43648,N_43472);
xor U46764 (N_46764,N_43780,N_44252);
and U46765 (N_46765,N_43254,N_43408);
and U46766 (N_46766,N_44574,N_44348);
and U46767 (N_46767,N_43238,N_44519);
nor U46768 (N_46768,N_43562,N_42957);
and U46769 (N_46769,N_43471,N_43138);
or U46770 (N_46770,N_42794,N_42844);
nor U46771 (N_46771,N_44270,N_44726);
nor U46772 (N_46772,N_44285,N_44444);
or U46773 (N_46773,N_42832,N_43360);
or U46774 (N_46774,N_43761,N_44673);
or U46775 (N_46775,N_44681,N_42555);
nand U46776 (N_46776,N_44765,N_42996);
or U46777 (N_46777,N_44997,N_43922);
nor U46778 (N_46778,N_44439,N_44434);
xor U46779 (N_46779,N_44530,N_42583);
and U46780 (N_46780,N_44530,N_44061);
xnor U46781 (N_46781,N_43479,N_44412);
and U46782 (N_46782,N_44827,N_42992);
and U46783 (N_46783,N_44728,N_44638);
nand U46784 (N_46784,N_43203,N_42823);
xor U46785 (N_46785,N_43936,N_44017);
nor U46786 (N_46786,N_43168,N_43529);
or U46787 (N_46787,N_43315,N_43448);
or U46788 (N_46788,N_44694,N_43475);
nand U46789 (N_46789,N_42953,N_44523);
and U46790 (N_46790,N_43834,N_43922);
and U46791 (N_46791,N_44640,N_44932);
or U46792 (N_46792,N_43164,N_43207);
or U46793 (N_46793,N_43723,N_42973);
or U46794 (N_46794,N_44230,N_42554);
and U46795 (N_46795,N_44616,N_43643);
nand U46796 (N_46796,N_43471,N_42601);
nand U46797 (N_46797,N_44934,N_44692);
xnor U46798 (N_46798,N_44872,N_43560);
nand U46799 (N_46799,N_44121,N_44043);
or U46800 (N_46800,N_43980,N_43027);
and U46801 (N_46801,N_44610,N_43829);
or U46802 (N_46802,N_42766,N_44599);
or U46803 (N_46803,N_44709,N_42569);
or U46804 (N_46804,N_44815,N_43445);
or U46805 (N_46805,N_44781,N_42543);
xnor U46806 (N_46806,N_43545,N_43998);
or U46807 (N_46807,N_43353,N_43115);
xnor U46808 (N_46808,N_43943,N_43760);
nor U46809 (N_46809,N_43424,N_44202);
and U46810 (N_46810,N_43418,N_44054);
or U46811 (N_46811,N_44658,N_42637);
nor U46812 (N_46812,N_43336,N_42924);
and U46813 (N_46813,N_44879,N_42789);
nor U46814 (N_46814,N_43094,N_44169);
xor U46815 (N_46815,N_44472,N_43176);
nor U46816 (N_46816,N_44250,N_43928);
nand U46817 (N_46817,N_44618,N_43247);
nor U46818 (N_46818,N_44375,N_42977);
xnor U46819 (N_46819,N_42864,N_43754);
and U46820 (N_46820,N_44481,N_42750);
nand U46821 (N_46821,N_43635,N_42786);
and U46822 (N_46822,N_44873,N_44995);
xnor U46823 (N_46823,N_42771,N_42925);
xnor U46824 (N_46824,N_44058,N_44550);
xor U46825 (N_46825,N_42871,N_42830);
nor U46826 (N_46826,N_43827,N_44538);
nor U46827 (N_46827,N_44738,N_43190);
xor U46828 (N_46828,N_44051,N_43995);
or U46829 (N_46829,N_44484,N_43610);
or U46830 (N_46830,N_44481,N_43902);
and U46831 (N_46831,N_42795,N_44136);
xor U46832 (N_46832,N_42651,N_44338);
or U46833 (N_46833,N_44070,N_42828);
or U46834 (N_46834,N_43483,N_43925);
xor U46835 (N_46835,N_42634,N_42675);
or U46836 (N_46836,N_43488,N_42759);
nand U46837 (N_46837,N_44343,N_44530);
and U46838 (N_46838,N_44903,N_43795);
or U46839 (N_46839,N_44981,N_43600);
nand U46840 (N_46840,N_42535,N_44166);
nor U46841 (N_46841,N_43547,N_43199);
nor U46842 (N_46842,N_43864,N_43756);
and U46843 (N_46843,N_43960,N_44917);
nand U46844 (N_46844,N_44060,N_44778);
and U46845 (N_46845,N_44132,N_44266);
or U46846 (N_46846,N_44726,N_44372);
nor U46847 (N_46847,N_42733,N_44332);
nand U46848 (N_46848,N_42963,N_44985);
or U46849 (N_46849,N_42569,N_43849);
nor U46850 (N_46850,N_44490,N_44503);
nand U46851 (N_46851,N_43105,N_43014);
or U46852 (N_46852,N_44940,N_43480);
nand U46853 (N_46853,N_43718,N_43207);
nor U46854 (N_46854,N_43389,N_44929);
or U46855 (N_46855,N_44032,N_44733);
xor U46856 (N_46856,N_44547,N_44459);
or U46857 (N_46857,N_43152,N_43162);
and U46858 (N_46858,N_44161,N_42788);
nand U46859 (N_46859,N_43177,N_43423);
and U46860 (N_46860,N_43951,N_43549);
and U46861 (N_46861,N_44793,N_44949);
or U46862 (N_46862,N_44165,N_44091);
nor U46863 (N_46863,N_43012,N_42728);
nor U46864 (N_46864,N_42802,N_43719);
and U46865 (N_46865,N_43280,N_44312);
xnor U46866 (N_46866,N_43654,N_44612);
and U46867 (N_46867,N_42930,N_43561);
xor U46868 (N_46868,N_42588,N_43215);
or U46869 (N_46869,N_44528,N_43383);
xnor U46870 (N_46870,N_44314,N_43386);
and U46871 (N_46871,N_42944,N_43175);
xor U46872 (N_46872,N_42910,N_43860);
xnor U46873 (N_46873,N_42726,N_44913);
xnor U46874 (N_46874,N_42754,N_43038);
and U46875 (N_46875,N_44827,N_44248);
xnor U46876 (N_46876,N_43722,N_43224);
xor U46877 (N_46877,N_42549,N_43451);
nand U46878 (N_46878,N_42580,N_44062);
nand U46879 (N_46879,N_42563,N_44873);
xor U46880 (N_46880,N_43875,N_43227);
nor U46881 (N_46881,N_44701,N_44496);
nor U46882 (N_46882,N_42773,N_44107);
nor U46883 (N_46883,N_44124,N_44939);
or U46884 (N_46884,N_42637,N_43261);
and U46885 (N_46885,N_43874,N_42923);
nand U46886 (N_46886,N_44941,N_44792);
and U46887 (N_46887,N_43652,N_43470);
and U46888 (N_46888,N_43749,N_44823);
nand U46889 (N_46889,N_43961,N_43943);
or U46890 (N_46890,N_44014,N_44397);
or U46891 (N_46891,N_44688,N_42868);
nor U46892 (N_46892,N_42748,N_43554);
xnor U46893 (N_46893,N_43232,N_43886);
nand U46894 (N_46894,N_43928,N_43936);
nand U46895 (N_46895,N_43433,N_43915);
nand U46896 (N_46896,N_43658,N_44238);
and U46897 (N_46897,N_44972,N_44467);
nor U46898 (N_46898,N_43401,N_43658);
nor U46899 (N_46899,N_44155,N_44154);
xnor U46900 (N_46900,N_44079,N_43605);
nand U46901 (N_46901,N_44639,N_43443);
xor U46902 (N_46902,N_43451,N_42545);
xnor U46903 (N_46903,N_43451,N_44941);
nand U46904 (N_46904,N_44027,N_44253);
xnor U46905 (N_46905,N_43202,N_43156);
nor U46906 (N_46906,N_43181,N_44770);
nand U46907 (N_46907,N_42991,N_44192);
or U46908 (N_46908,N_42835,N_44534);
xor U46909 (N_46909,N_44271,N_43910);
or U46910 (N_46910,N_43119,N_44362);
nand U46911 (N_46911,N_44620,N_44849);
xor U46912 (N_46912,N_42590,N_43672);
and U46913 (N_46913,N_43858,N_44667);
or U46914 (N_46914,N_42705,N_42539);
nor U46915 (N_46915,N_43070,N_43239);
nor U46916 (N_46916,N_43642,N_43990);
xor U46917 (N_46917,N_42777,N_44923);
nor U46918 (N_46918,N_42845,N_44375);
nand U46919 (N_46919,N_42865,N_44116);
or U46920 (N_46920,N_42591,N_43469);
nor U46921 (N_46921,N_43340,N_44505);
nor U46922 (N_46922,N_44417,N_43936);
and U46923 (N_46923,N_43338,N_43589);
or U46924 (N_46924,N_43742,N_42836);
nand U46925 (N_46925,N_42561,N_43335);
nand U46926 (N_46926,N_43646,N_43426);
or U46927 (N_46927,N_43058,N_42894);
and U46928 (N_46928,N_43241,N_43833);
or U46929 (N_46929,N_44037,N_43733);
nor U46930 (N_46930,N_44430,N_43479);
nand U46931 (N_46931,N_44573,N_44977);
nor U46932 (N_46932,N_43481,N_43964);
nand U46933 (N_46933,N_42655,N_43352);
xnor U46934 (N_46934,N_42930,N_43152);
and U46935 (N_46935,N_44654,N_44523);
or U46936 (N_46936,N_43349,N_43100);
xnor U46937 (N_46937,N_42727,N_42675);
nand U46938 (N_46938,N_44552,N_42906);
or U46939 (N_46939,N_43496,N_44954);
xnor U46940 (N_46940,N_43427,N_42649);
and U46941 (N_46941,N_44733,N_43233);
and U46942 (N_46942,N_42563,N_43053);
and U46943 (N_46943,N_43341,N_44567);
nor U46944 (N_46944,N_42803,N_43827);
nor U46945 (N_46945,N_44033,N_44376);
and U46946 (N_46946,N_43759,N_43361);
or U46947 (N_46947,N_44766,N_44207);
and U46948 (N_46948,N_43976,N_43660);
nor U46949 (N_46949,N_42564,N_44190);
xor U46950 (N_46950,N_42789,N_42764);
nand U46951 (N_46951,N_43969,N_42694);
and U46952 (N_46952,N_44314,N_43299);
nand U46953 (N_46953,N_44398,N_43962);
xnor U46954 (N_46954,N_43602,N_42641);
or U46955 (N_46955,N_42920,N_44175);
nor U46956 (N_46956,N_43432,N_42877);
and U46957 (N_46957,N_44786,N_43647);
nand U46958 (N_46958,N_44085,N_43937);
or U46959 (N_46959,N_44962,N_44508);
xnor U46960 (N_46960,N_42563,N_42616);
xor U46961 (N_46961,N_42581,N_43859);
or U46962 (N_46962,N_44880,N_43270);
or U46963 (N_46963,N_42848,N_44765);
xnor U46964 (N_46964,N_44648,N_42945);
nand U46965 (N_46965,N_44976,N_44141);
nand U46966 (N_46966,N_44246,N_43787);
nor U46967 (N_46967,N_42807,N_43386);
xor U46968 (N_46968,N_43368,N_44348);
xor U46969 (N_46969,N_44034,N_44060);
and U46970 (N_46970,N_42587,N_43795);
and U46971 (N_46971,N_44429,N_44914);
nand U46972 (N_46972,N_44058,N_43147);
or U46973 (N_46973,N_43574,N_43040);
nor U46974 (N_46974,N_44886,N_43899);
nor U46975 (N_46975,N_44099,N_42519);
or U46976 (N_46976,N_44438,N_44588);
nand U46977 (N_46977,N_44030,N_44532);
xnor U46978 (N_46978,N_44628,N_44459);
nor U46979 (N_46979,N_43426,N_44121);
xor U46980 (N_46980,N_44892,N_44645);
or U46981 (N_46981,N_44339,N_43846);
nand U46982 (N_46982,N_44604,N_42689);
xor U46983 (N_46983,N_43516,N_44438);
or U46984 (N_46984,N_44069,N_43763);
and U46985 (N_46985,N_43583,N_43389);
nor U46986 (N_46986,N_43231,N_42862);
xor U46987 (N_46987,N_42503,N_44239);
nor U46988 (N_46988,N_44843,N_42707);
nand U46989 (N_46989,N_42897,N_42874);
nand U46990 (N_46990,N_44312,N_43796);
or U46991 (N_46991,N_44585,N_44945);
nor U46992 (N_46992,N_43777,N_44043);
and U46993 (N_46993,N_43406,N_44965);
and U46994 (N_46994,N_42876,N_44476);
and U46995 (N_46995,N_42686,N_44099);
nand U46996 (N_46996,N_44851,N_44479);
nor U46997 (N_46997,N_43481,N_44190);
nor U46998 (N_46998,N_43458,N_44036);
and U46999 (N_46999,N_42927,N_43009);
nor U47000 (N_47000,N_43408,N_44422);
xor U47001 (N_47001,N_43437,N_43489);
nand U47002 (N_47002,N_42819,N_44790);
nand U47003 (N_47003,N_44797,N_43321);
and U47004 (N_47004,N_44557,N_43014);
or U47005 (N_47005,N_43518,N_44988);
nand U47006 (N_47006,N_44051,N_44016);
nor U47007 (N_47007,N_43795,N_43366);
or U47008 (N_47008,N_43277,N_43869);
xnor U47009 (N_47009,N_44875,N_42934);
nor U47010 (N_47010,N_42991,N_42800);
nand U47011 (N_47011,N_42556,N_42503);
xor U47012 (N_47012,N_44579,N_44995);
and U47013 (N_47013,N_43830,N_44877);
or U47014 (N_47014,N_43045,N_44408);
xnor U47015 (N_47015,N_43090,N_44751);
xor U47016 (N_47016,N_43550,N_42958);
nand U47017 (N_47017,N_44240,N_44724);
nand U47018 (N_47018,N_42845,N_43083);
nand U47019 (N_47019,N_44355,N_43966);
or U47020 (N_47020,N_43595,N_44288);
nand U47021 (N_47021,N_43995,N_44249);
nand U47022 (N_47022,N_44184,N_44680);
nand U47023 (N_47023,N_43207,N_44399);
xor U47024 (N_47024,N_43515,N_44493);
or U47025 (N_47025,N_42597,N_42885);
xor U47026 (N_47026,N_43302,N_43452);
or U47027 (N_47027,N_43370,N_44902);
nand U47028 (N_47028,N_42585,N_44116);
nor U47029 (N_47029,N_43704,N_43129);
or U47030 (N_47030,N_43203,N_43297);
nand U47031 (N_47031,N_43084,N_42637);
and U47032 (N_47032,N_43901,N_42989);
and U47033 (N_47033,N_42550,N_44317);
or U47034 (N_47034,N_43351,N_44095);
xor U47035 (N_47035,N_43142,N_43671);
xor U47036 (N_47036,N_43849,N_42782);
and U47037 (N_47037,N_43223,N_42536);
or U47038 (N_47038,N_43168,N_44420);
or U47039 (N_47039,N_44593,N_44965);
xnor U47040 (N_47040,N_43094,N_42818);
and U47041 (N_47041,N_42816,N_43051);
or U47042 (N_47042,N_44789,N_44422);
and U47043 (N_47043,N_42920,N_42916);
xnor U47044 (N_47044,N_43774,N_43636);
and U47045 (N_47045,N_44085,N_43318);
and U47046 (N_47046,N_43773,N_42982);
or U47047 (N_47047,N_43485,N_42767);
nor U47048 (N_47048,N_42721,N_44554);
nand U47049 (N_47049,N_42723,N_43220);
or U47050 (N_47050,N_42670,N_42568);
nor U47051 (N_47051,N_44005,N_43174);
and U47052 (N_47052,N_43596,N_44282);
or U47053 (N_47053,N_43116,N_42507);
nor U47054 (N_47054,N_42635,N_43917);
xnor U47055 (N_47055,N_43661,N_43717);
nand U47056 (N_47056,N_42716,N_42754);
nor U47057 (N_47057,N_44336,N_42897);
nand U47058 (N_47058,N_43243,N_44375);
nor U47059 (N_47059,N_44939,N_43239);
and U47060 (N_47060,N_43421,N_43049);
xor U47061 (N_47061,N_42974,N_43038);
or U47062 (N_47062,N_44331,N_43221);
nor U47063 (N_47063,N_43877,N_42545);
nand U47064 (N_47064,N_43916,N_44225);
nor U47065 (N_47065,N_43023,N_42735);
nor U47066 (N_47066,N_43661,N_42833);
and U47067 (N_47067,N_43495,N_43360);
xor U47068 (N_47068,N_42667,N_44457);
nor U47069 (N_47069,N_44575,N_42619);
or U47070 (N_47070,N_43798,N_42651);
nor U47071 (N_47071,N_43350,N_43591);
and U47072 (N_47072,N_42592,N_43148);
nand U47073 (N_47073,N_44320,N_43663);
xor U47074 (N_47074,N_43816,N_43641);
nand U47075 (N_47075,N_44551,N_44790);
or U47076 (N_47076,N_42549,N_44640);
nand U47077 (N_47077,N_44081,N_44307);
xor U47078 (N_47078,N_43868,N_43244);
or U47079 (N_47079,N_43417,N_43152);
nor U47080 (N_47080,N_43941,N_43580);
and U47081 (N_47081,N_44766,N_43600);
xor U47082 (N_47082,N_44265,N_43007);
xor U47083 (N_47083,N_44132,N_43266);
or U47084 (N_47084,N_44386,N_44351);
nor U47085 (N_47085,N_43497,N_43415);
nand U47086 (N_47086,N_43497,N_43525);
nor U47087 (N_47087,N_44775,N_44878);
and U47088 (N_47088,N_43871,N_43505);
or U47089 (N_47089,N_44427,N_43785);
and U47090 (N_47090,N_43437,N_42897);
or U47091 (N_47091,N_44494,N_43979);
nor U47092 (N_47092,N_42947,N_44431);
nor U47093 (N_47093,N_44968,N_43070);
xor U47094 (N_47094,N_44048,N_43483);
and U47095 (N_47095,N_44588,N_42713);
or U47096 (N_47096,N_43414,N_44102);
or U47097 (N_47097,N_44851,N_43937);
or U47098 (N_47098,N_43228,N_44990);
or U47099 (N_47099,N_44257,N_44681);
or U47100 (N_47100,N_43688,N_44068);
nor U47101 (N_47101,N_43125,N_44355);
nand U47102 (N_47102,N_43513,N_43673);
or U47103 (N_47103,N_43042,N_44037);
nor U47104 (N_47104,N_44670,N_44103);
or U47105 (N_47105,N_44413,N_44764);
nor U47106 (N_47106,N_43903,N_44748);
and U47107 (N_47107,N_42582,N_44948);
nand U47108 (N_47108,N_43375,N_43482);
and U47109 (N_47109,N_43875,N_43206);
nand U47110 (N_47110,N_43945,N_42501);
nand U47111 (N_47111,N_43435,N_43050);
or U47112 (N_47112,N_43629,N_43355);
and U47113 (N_47113,N_42863,N_44066);
or U47114 (N_47114,N_42832,N_44203);
xnor U47115 (N_47115,N_43212,N_42654);
and U47116 (N_47116,N_44086,N_43378);
or U47117 (N_47117,N_42579,N_43081);
xor U47118 (N_47118,N_42657,N_43486);
xnor U47119 (N_47119,N_42706,N_43198);
or U47120 (N_47120,N_43780,N_43704);
and U47121 (N_47121,N_42877,N_44889);
and U47122 (N_47122,N_42654,N_44135);
or U47123 (N_47123,N_42771,N_44202);
xor U47124 (N_47124,N_43417,N_44228);
and U47125 (N_47125,N_44261,N_44689);
nor U47126 (N_47126,N_44859,N_43529);
nor U47127 (N_47127,N_44011,N_42591);
and U47128 (N_47128,N_42910,N_44881);
and U47129 (N_47129,N_43272,N_43145);
nand U47130 (N_47130,N_43938,N_42696);
and U47131 (N_47131,N_42885,N_43487);
and U47132 (N_47132,N_43425,N_44425);
nor U47133 (N_47133,N_43200,N_43465);
nand U47134 (N_47134,N_42715,N_42896);
nand U47135 (N_47135,N_44240,N_44663);
or U47136 (N_47136,N_42646,N_43394);
or U47137 (N_47137,N_44964,N_43504);
and U47138 (N_47138,N_43051,N_42639);
nand U47139 (N_47139,N_44098,N_44572);
or U47140 (N_47140,N_43257,N_44736);
and U47141 (N_47141,N_44378,N_44329);
and U47142 (N_47142,N_42857,N_43816);
xor U47143 (N_47143,N_43742,N_43692);
xnor U47144 (N_47144,N_44816,N_44836);
and U47145 (N_47145,N_44492,N_44462);
xor U47146 (N_47146,N_44686,N_44361);
or U47147 (N_47147,N_43195,N_44950);
and U47148 (N_47148,N_44013,N_44680);
and U47149 (N_47149,N_44858,N_43444);
and U47150 (N_47150,N_42885,N_43213);
or U47151 (N_47151,N_43041,N_43558);
and U47152 (N_47152,N_43061,N_43856);
nand U47153 (N_47153,N_42651,N_44227);
nor U47154 (N_47154,N_44734,N_44524);
xnor U47155 (N_47155,N_44671,N_43288);
and U47156 (N_47156,N_43061,N_43696);
or U47157 (N_47157,N_43971,N_43928);
nand U47158 (N_47158,N_43988,N_44609);
xnor U47159 (N_47159,N_43506,N_42628);
xnor U47160 (N_47160,N_43314,N_44412);
nor U47161 (N_47161,N_44390,N_44654);
xnor U47162 (N_47162,N_43459,N_44401);
nor U47163 (N_47163,N_43922,N_44222);
and U47164 (N_47164,N_43872,N_44559);
or U47165 (N_47165,N_44882,N_43235);
nor U47166 (N_47166,N_44470,N_44728);
xnor U47167 (N_47167,N_42527,N_44370);
xnor U47168 (N_47168,N_44737,N_42810);
and U47169 (N_47169,N_43074,N_44517);
and U47170 (N_47170,N_44015,N_43742);
and U47171 (N_47171,N_44721,N_43366);
nand U47172 (N_47172,N_44004,N_43906);
nand U47173 (N_47173,N_44673,N_44936);
nand U47174 (N_47174,N_43631,N_43716);
nor U47175 (N_47175,N_43410,N_43337);
nand U47176 (N_47176,N_44197,N_44326);
xnor U47177 (N_47177,N_44486,N_44271);
and U47178 (N_47178,N_44049,N_43224);
xnor U47179 (N_47179,N_44216,N_44471);
or U47180 (N_47180,N_44265,N_43214);
or U47181 (N_47181,N_42652,N_44616);
and U47182 (N_47182,N_43987,N_43888);
nor U47183 (N_47183,N_43969,N_43668);
nand U47184 (N_47184,N_44673,N_44443);
nand U47185 (N_47185,N_44311,N_42520);
nor U47186 (N_47186,N_44651,N_43786);
xor U47187 (N_47187,N_43418,N_43714);
nand U47188 (N_47188,N_44313,N_42600);
xnor U47189 (N_47189,N_44488,N_44627);
and U47190 (N_47190,N_42808,N_44178);
nor U47191 (N_47191,N_43170,N_43897);
and U47192 (N_47192,N_44482,N_43914);
xnor U47193 (N_47193,N_43187,N_44609);
nor U47194 (N_47194,N_44331,N_43716);
nor U47195 (N_47195,N_43625,N_43193);
nand U47196 (N_47196,N_43342,N_43697);
nand U47197 (N_47197,N_44698,N_42888);
and U47198 (N_47198,N_44887,N_44287);
nand U47199 (N_47199,N_43151,N_43621);
xor U47200 (N_47200,N_43589,N_44667);
nor U47201 (N_47201,N_43076,N_43631);
nor U47202 (N_47202,N_43028,N_44362);
and U47203 (N_47203,N_42786,N_43306);
nand U47204 (N_47204,N_44568,N_43128);
nor U47205 (N_47205,N_43205,N_44556);
xnor U47206 (N_47206,N_44046,N_44082);
nor U47207 (N_47207,N_44874,N_44997);
nor U47208 (N_47208,N_43576,N_43929);
xnor U47209 (N_47209,N_43039,N_43176);
and U47210 (N_47210,N_44278,N_43986);
nand U47211 (N_47211,N_43370,N_44807);
and U47212 (N_47212,N_43042,N_42768);
nor U47213 (N_47213,N_43782,N_43273);
xnor U47214 (N_47214,N_43931,N_43107);
xor U47215 (N_47215,N_44092,N_43106);
nor U47216 (N_47216,N_44694,N_43900);
nand U47217 (N_47217,N_43931,N_44213);
or U47218 (N_47218,N_43132,N_43433);
nor U47219 (N_47219,N_44024,N_44568);
nor U47220 (N_47220,N_44645,N_43349);
and U47221 (N_47221,N_43483,N_43308);
and U47222 (N_47222,N_43765,N_42689);
or U47223 (N_47223,N_44833,N_43003);
nand U47224 (N_47224,N_43731,N_43658);
nand U47225 (N_47225,N_44028,N_44227);
nand U47226 (N_47226,N_42580,N_44258);
or U47227 (N_47227,N_44491,N_43713);
nor U47228 (N_47228,N_42706,N_44656);
xor U47229 (N_47229,N_43741,N_42919);
nand U47230 (N_47230,N_42865,N_42616);
nand U47231 (N_47231,N_44140,N_44247);
nor U47232 (N_47232,N_44953,N_42606);
and U47233 (N_47233,N_43004,N_43775);
nor U47234 (N_47234,N_43945,N_43999);
and U47235 (N_47235,N_44108,N_43631);
nor U47236 (N_47236,N_43466,N_43066);
xnor U47237 (N_47237,N_43458,N_43357);
and U47238 (N_47238,N_44519,N_43812);
or U47239 (N_47239,N_42681,N_43512);
nand U47240 (N_47240,N_44686,N_44231);
nand U47241 (N_47241,N_44081,N_44701);
nand U47242 (N_47242,N_43348,N_44997);
nand U47243 (N_47243,N_43034,N_44574);
and U47244 (N_47244,N_43327,N_43551);
or U47245 (N_47245,N_43343,N_44824);
nand U47246 (N_47246,N_44622,N_42630);
xor U47247 (N_47247,N_44469,N_43238);
xnor U47248 (N_47248,N_43629,N_43772);
nor U47249 (N_47249,N_43532,N_43657);
or U47250 (N_47250,N_43592,N_44774);
and U47251 (N_47251,N_44847,N_43667);
nand U47252 (N_47252,N_44350,N_43567);
xnor U47253 (N_47253,N_43217,N_43351);
xor U47254 (N_47254,N_43403,N_43130);
and U47255 (N_47255,N_42874,N_43560);
nand U47256 (N_47256,N_43754,N_43399);
xnor U47257 (N_47257,N_43595,N_44283);
nor U47258 (N_47258,N_43189,N_44582);
xnor U47259 (N_47259,N_43533,N_43854);
nand U47260 (N_47260,N_43514,N_44655);
and U47261 (N_47261,N_43405,N_43446);
and U47262 (N_47262,N_42575,N_42787);
xnor U47263 (N_47263,N_44745,N_43935);
nand U47264 (N_47264,N_44593,N_44586);
nor U47265 (N_47265,N_44402,N_43587);
nor U47266 (N_47266,N_43815,N_44852);
and U47267 (N_47267,N_43890,N_42916);
xor U47268 (N_47268,N_43116,N_44335);
nand U47269 (N_47269,N_42932,N_44033);
nand U47270 (N_47270,N_42926,N_42562);
nand U47271 (N_47271,N_44181,N_44401);
nand U47272 (N_47272,N_43049,N_44927);
and U47273 (N_47273,N_43553,N_42919);
or U47274 (N_47274,N_44175,N_43154);
or U47275 (N_47275,N_44272,N_43519);
xnor U47276 (N_47276,N_43500,N_43302);
nand U47277 (N_47277,N_44832,N_44158);
nor U47278 (N_47278,N_44644,N_44737);
nand U47279 (N_47279,N_44121,N_42882);
nor U47280 (N_47280,N_44461,N_44593);
and U47281 (N_47281,N_43714,N_43376);
nor U47282 (N_47282,N_44770,N_42993);
or U47283 (N_47283,N_42586,N_43073);
or U47284 (N_47284,N_44929,N_43244);
nor U47285 (N_47285,N_43041,N_43505);
and U47286 (N_47286,N_44991,N_44411);
nand U47287 (N_47287,N_43179,N_43892);
nand U47288 (N_47288,N_43042,N_43861);
nor U47289 (N_47289,N_43904,N_44387);
nor U47290 (N_47290,N_43472,N_43403);
and U47291 (N_47291,N_43827,N_42534);
nand U47292 (N_47292,N_44679,N_44697);
and U47293 (N_47293,N_43999,N_42783);
nand U47294 (N_47294,N_43797,N_42811);
xor U47295 (N_47295,N_44381,N_44701);
nand U47296 (N_47296,N_43727,N_44826);
xor U47297 (N_47297,N_43001,N_44313);
nor U47298 (N_47298,N_43465,N_43044);
xnor U47299 (N_47299,N_43895,N_42767);
and U47300 (N_47300,N_42920,N_43178);
or U47301 (N_47301,N_42546,N_43271);
and U47302 (N_47302,N_42565,N_44164);
or U47303 (N_47303,N_44401,N_44238);
xnor U47304 (N_47304,N_43365,N_42510);
nand U47305 (N_47305,N_43767,N_44838);
nand U47306 (N_47306,N_44926,N_42647);
nor U47307 (N_47307,N_43252,N_44585);
or U47308 (N_47308,N_43626,N_44413);
and U47309 (N_47309,N_43680,N_43003);
or U47310 (N_47310,N_43145,N_42947);
and U47311 (N_47311,N_43008,N_44085);
or U47312 (N_47312,N_44755,N_43215);
xnor U47313 (N_47313,N_43165,N_43195);
xor U47314 (N_47314,N_44807,N_44808);
nand U47315 (N_47315,N_44812,N_43473);
nor U47316 (N_47316,N_43526,N_43889);
and U47317 (N_47317,N_43921,N_43815);
and U47318 (N_47318,N_43764,N_44816);
xnor U47319 (N_47319,N_43227,N_44685);
nand U47320 (N_47320,N_44537,N_44990);
and U47321 (N_47321,N_43260,N_42612);
nand U47322 (N_47322,N_43382,N_43639);
and U47323 (N_47323,N_44245,N_42681);
xnor U47324 (N_47324,N_42683,N_42730);
or U47325 (N_47325,N_44471,N_43426);
xnor U47326 (N_47326,N_42947,N_44270);
xor U47327 (N_47327,N_43171,N_43685);
nor U47328 (N_47328,N_44426,N_43767);
and U47329 (N_47329,N_44263,N_44989);
nor U47330 (N_47330,N_42607,N_43226);
nand U47331 (N_47331,N_44018,N_44492);
nor U47332 (N_47332,N_42984,N_42981);
or U47333 (N_47333,N_44367,N_43233);
xor U47334 (N_47334,N_42903,N_44146);
xor U47335 (N_47335,N_44619,N_43357);
and U47336 (N_47336,N_44392,N_42800);
nor U47337 (N_47337,N_43569,N_43597);
or U47338 (N_47338,N_44670,N_43740);
or U47339 (N_47339,N_43007,N_43976);
nand U47340 (N_47340,N_43869,N_42891);
xnor U47341 (N_47341,N_44135,N_42979);
and U47342 (N_47342,N_42508,N_44653);
xor U47343 (N_47343,N_44352,N_44129);
and U47344 (N_47344,N_43458,N_42778);
nor U47345 (N_47345,N_44845,N_44292);
xnor U47346 (N_47346,N_42664,N_44540);
nand U47347 (N_47347,N_43067,N_43236);
xnor U47348 (N_47348,N_42922,N_42674);
nand U47349 (N_47349,N_43350,N_44956);
nand U47350 (N_47350,N_43078,N_42878);
and U47351 (N_47351,N_44074,N_44351);
xnor U47352 (N_47352,N_42517,N_44565);
and U47353 (N_47353,N_44956,N_43067);
or U47354 (N_47354,N_44484,N_44550);
and U47355 (N_47355,N_43430,N_43670);
or U47356 (N_47356,N_44357,N_44806);
or U47357 (N_47357,N_43078,N_42752);
and U47358 (N_47358,N_44890,N_43203);
xnor U47359 (N_47359,N_44762,N_44498);
nand U47360 (N_47360,N_42644,N_43923);
or U47361 (N_47361,N_43208,N_44526);
nand U47362 (N_47362,N_42707,N_42588);
and U47363 (N_47363,N_42934,N_43080);
nand U47364 (N_47364,N_44506,N_44646);
xor U47365 (N_47365,N_43950,N_43873);
or U47366 (N_47366,N_44602,N_44434);
nor U47367 (N_47367,N_43322,N_43362);
and U47368 (N_47368,N_42885,N_44078);
nor U47369 (N_47369,N_43306,N_42552);
or U47370 (N_47370,N_43989,N_44014);
xor U47371 (N_47371,N_43665,N_43865);
or U47372 (N_47372,N_42871,N_44888);
or U47373 (N_47373,N_44955,N_44992);
nand U47374 (N_47374,N_42973,N_44869);
and U47375 (N_47375,N_43780,N_42621);
xor U47376 (N_47376,N_42716,N_43661);
nor U47377 (N_47377,N_42892,N_43586);
xnor U47378 (N_47378,N_44709,N_44111);
nand U47379 (N_47379,N_43501,N_43016);
or U47380 (N_47380,N_43125,N_43824);
or U47381 (N_47381,N_44040,N_43857);
and U47382 (N_47382,N_42936,N_43433);
nand U47383 (N_47383,N_43897,N_42563);
nand U47384 (N_47384,N_44095,N_43533);
xor U47385 (N_47385,N_42549,N_44480);
xor U47386 (N_47386,N_43863,N_44490);
and U47387 (N_47387,N_43087,N_42728);
and U47388 (N_47388,N_43754,N_44762);
nand U47389 (N_47389,N_44217,N_42631);
and U47390 (N_47390,N_44711,N_43218);
nand U47391 (N_47391,N_43880,N_44553);
xnor U47392 (N_47392,N_42924,N_44025);
nor U47393 (N_47393,N_43576,N_43751);
nor U47394 (N_47394,N_44319,N_43476);
nand U47395 (N_47395,N_43010,N_42906);
nor U47396 (N_47396,N_42841,N_44867);
nand U47397 (N_47397,N_44007,N_42614);
or U47398 (N_47398,N_44286,N_43965);
xor U47399 (N_47399,N_44367,N_44219);
xor U47400 (N_47400,N_43637,N_44582);
and U47401 (N_47401,N_43207,N_44733);
nand U47402 (N_47402,N_42891,N_43590);
nand U47403 (N_47403,N_44985,N_43056);
xor U47404 (N_47404,N_42806,N_43854);
nor U47405 (N_47405,N_42565,N_43627);
nor U47406 (N_47406,N_44862,N_42847);
and U47407 (N_47407,N_43252,N_44658);
xor U47408 (N_47408,N_42753,N_43748);
xnor U47409 (N_47409,N_44667,N_42505);
nand U47410 (N_47410,N_43332,N_44683);
or U47411 (N_47411,N_43166,N_43941);
and U47412 (N_47412,N_44953,N_43017);
xnor U47413 (N_47413,N_43664,N_43271);
or U47414 (N_47414,N_44595,N_43691);
nand U47415 (N_47415,N_43388,N_44239);
xnor U47416 (N_47416,N_43764,N_43451);
or U47417 (N_47417,N_44873,N_44986);
xnor U47418 (N_47418,N_44678,N_44424);
nand U47419 (N_47419,N_44619,N_44567);
nand U47420 (N_47420,N_42570,N_42898);
or U47421 (N_47421,N_44084,N_43631);
xnor U47422 (N_47422,N_44315,N_43029);
or U47423 (N_47423,N_44196,N_43219);
or U47424 (N_47424,N_42517,N_43869);
and U47425 (N_47425,N_44383,N_44504);
nand U47426 (N_47426,N_43984,N_44030);
xnor U47427 (N_47427,N_44612,N_44636);
xor U47428 (N_47428,N_44317,N_43593);
nor U47429 (N_47429,N_43939,N_43386);
or U47430 (N_47430,N_42714,N_44916);
xnor U47431 (N_47431,N_43253,N_43203);
nor U47432 (N_47432,N_43107,N_44789);
or U47433 (N_47433,N_43250,N_43364);
nand U47434 (N_47434,N_43871,N_43740);
and U47435 (N_47435,N_43648,N_43757);
nor U47436 (N_47436,N_43172,N_42921);
xor U47437 (N_47437,N_43501,N_43993);
and U47438 (N_47438,N_43930,N_44740);
xnor U47439 (N_47439,N_43200,N_42633);
nor U47440 (N_47440,N_43140,N_44974);
xor U47441 (N_47441,N_43929,N_44068);
nand U47442 (N_47442,N_42828,N_43354);
nand U47443 (N_47443,N_43838,N_42794);
nor U47444 (N_47444,N_42674,N_43493);
nand U47445 (N_47445,N_43999,N_42640);
nor U47446 (N_47446,N_44067,N_42843);
nor U47447 (N_47447,N_44213,N_43377);
xor U47448 (N_47448,N_42629,N_42971);
nand U47449 (N_47449,N_42681,N_43188);
xor U47450 (N_47450,N_43909,N_42791);
nand U47451 (N_47451,N_44181,N_42961);
or U47452 (N_47452,N_44546,N_43609);
nand U47453 (N_47453,N_43535,N_44135);
nand U47454 (N_47454,N_43149,N_42525);
xnor U47455 (N_47455,N_44192,N_43273);
nor U47456 (N_47456,N_42947,N_42661);
nor U47457 (N_47457,N_42941,N_44522);
or U47458 (N_47458,N_42602,N_43465);
nor U47459 (N_47459,N_43864,N_44613);
and U47460 (N_47460,N_43136,N_42868);
nor U47461 (N_47461,N_43610,N_43882);
nor U47462 (N_47462,N_44683,N_43506);
nor U47463 (N_47463,N_44009,N_44143);
nand U47464 (N_47464,N_42816,N_43492);
or U47465 (N_47465,N_43904,N_43709);
and U47466 (N_47466,N_42802,N_43580);
nand U47467 (N_47467,N_44312,N_42952);
or U47468 (N_47468,N_42764,N_43355);
nand U47469 (N_47469,N_43256,N_43908);
or U47470 (N_47470,N_42688,N_42912);
or U47471 (N_47471,N_44369,N_44690);
nor U47472 (N_47472,N_43677,N_44871);
and U47473 (N_47473,N_43312,N_44908);
nor U47474 (N_47474,N_43808,N_43570);
nor U47475 (N_47475,N_43645,N_43764);
nor U47476 (N_47476,N_44202,N_43606);
or U47477 (N_47477,N_44214,N_42689);
nand U47478 (N_47478,N_44606,N_43229);
or U47479 (N_47479,N_44499,N_43067);
and U47480 (N_47480,N_44293,N_43595);
or U47481 (N_47481,N_43873,N_44041);
nand U47482 (N_47482,N_43498,N_42937);
nor U47483 (N_47483,N_43956,N_43331);
nand U47484 (N_47484,N_44707,N_44518);
and U47485 (N_47485,N_44034,N_43239);
nand U47486 (N_47486,N_43731,N_44484);
nand U47487 (N_47487,N_42916,N_43776);
nand U47488 (N_47488,N_43184,N_44638);
or U47489 (N_47489,N_43506,N_43494);
and U47490 (N_47490,N_44408,N_42615);
xnor U47491 (N_47491,N_44716,N_44942);
and U47492 (N_47492,N_44767,N_44193);
or U47493 (N_47493,N_44248,N_44356);
and U47494 (N_47494,N_43541,N_44476);
nand U47495 (N_47495,N_44214,N_43566);
nor U47496 (N_47496,N_44205,N_42931);
nor U47497 (N_47497,N_42859,N_44436);
nand U47498 (N_47498,N_43921,N_43705);
nor U47499 (N_47499,N_42795,N_43830);
nor U47500 (N_47500,N_46094,N_47232);
nor U47501 (N_47501,N_47083,N_46662);
or U47502 (N_47502,N_45258,N_45407);
and U47503 (N_47503,N_46404,N_46116);
or U47504 (N_47504,N_46356,N_45664);
xnor U47505 (N_47505,N_45637,N_45220);
and U47506 (N_47506,N_45232,N_47064);
or U47507 (N_47507,N_46810,N_46566);
or U47508 (N_47508,N_45816,N_45646);
nand U47509 (N_47509,N_46440,N_47352);
and U47510 (N_47510,N_46861,N_47192);
and U47511 (N_47511,N_46848,N_47123);
nand U47512 (N_47512,N_46748,N_46881);
and U47513 (N_47513,N_46273,N_47166);
nand U47514 (N_47514,N_45808,N_45033);
nor U47515 (N_47515,N_45070,N_47258);
or U47516 (N_47516,N_46767,N_45050);
nand U47517 (N_47517,N_46766,N_46056);
and U47518 (N_47518,N_47145,N_45511);
nand U47519 (N_47519,N_45910,N_46971);
nor U47520 (N_47520,N_46202,N_46612);
and U47521 (N_47521,N_47372,N_47280);
and U47522 (N_47522,N_46235,N_45079);
xnor U47523 (N_47523,N_46561,N_46913);
nor U47524 (N_47524,N_45672,N_47117);
nor U47525 (N_47525,N_46554,N_46629);
nand U47526 (N_47526,N_45130,N_47034);
or U47527 (N_47527,N_47468,N_45777);
nand U47528 (N_47528,N_46528,N_46306);
xnor U47529 (N_47529,N_46258,N_47311);
nor U47530 (N_47530,N_46482,N_46130);
nand U47531 (N_47531,N_46802,N_47025);
xnor U47532 (N_47532,N_47479,N_45110);
and U47533 (N_47533,N_45668,N_47475);
and U47534 (N_47534,N_45817,N_46979);
or U47535 (N_47535,N_46840,N_45676);
nor U47536 (N_47536,N_45785,N_45820);
and U47537 (N_47537,N_45411,N_45546);
xnor U47538 (N_47538,N_47320,N_47128);
nand U47539 (N_47539,N_45206,N_45751);
xor U47540 (N_47540,N_46497,N_45889);
nand U47541 (N_47541,N_46206,N_46428);
nor U47542 (N_47542,N_47499,N_45291);
xor U47543 (N_47543,N_45461,N_46049);
nor U47544 (N_47544,N_45918,N_46562);
nor U47545 (N_47545,N_45954,N_46185);
nand U47546 (N_47546,N_47251,N_46184);
or U47547 (N_47547,N_46026,N_46289);
and U47548 (N_47548,N_46208,N_46768);
nor U47549 (N_47549,N_47329,N_45832);
xnor U47550 (N_47550,N_47336,N_46032);
or U47551 (N_47551,N_46901,N_45199);
and U47552 (N_47552,N_45690,N_46010);
xnor U47553 (N_47553,N_47481,N_45240);
xor U47554 (N_47554,N_46285,N_47409);
xor U47555 (N_47555,N_46892,N_46795);
xnor U47556 (N_47556,N_46695,N_45748);
nand U47557 (N_47557,N_47387,N_47045);
nor U47558 (N_47558,N_46948,N_47066);
xor U47559 (N_47559,N_47164,N_47285);
xnor U47560 (N_47560,N_45192,N_45457);
or U47561 (N_47561,N_46283,N_45340);
nand U47562 (N_47562,N_46376,N_46336);
nor U47563 (N_47563,N_47440,N_46242);
or U47564 (N_47564,N_46666,N_46035);
nand U47565 (N_47565,N_45562,N_46016);
or U47566 (N_47566,N_45567,N_46656);
xnor U47567 (N_47567,N_45024,N_45115);
and U47568 (N_47568,N_45507,N_45286);
or U47569 (N_47569,N_45011,N_47035);
nand U47570 (N_47570,N_46197,N_47058);
or U47571 (N_47571,N_45824,N_46655);
nand U47572 (N_47572,N_45594,N_45884);
nor U47573 (N_47573,N_45685,N_46251);
nor U47574 (N_47574,N_45492,N_45547);
nand U47575 (N_47575,N_47350,N_47093);
nand U47576 (N_47576,N_46292,N_46792);
or U47577 (N_47577,N_46644,N_46316);
nor U47578 (N_47578,N_46300,N_46790);
and U47579 (N_47579,N_46583,N_46863);
xnor U47580 (N_47580,N_46218,N_47428);
xnor U47581 (N_47581,N_47340,N_45093);
nand U47582 (N_47582,N_47410,N_46159);
or U47583 (N_47583,N_45628,N_45166);
or U47584 (N_47584,N_46494,N_46951);
or U47585 (N_47585,N_46024,N_46875);
nor U47586 (N_47586,N_47013,N_45607);
and U47587 (N_47587,N_45553,N_46133);
or U47588 (N_47588,N_46651,N_45635);
nand U47589 (N_47589,N_45727,N_47491);
xnor U47590 (N_47590,N_47161,N_47363);
nand U47591 (N_47591,N_45657,N_46304);
or U47592 (N_47592,N_46363,N_46592);
nand U47593 (N_47593,N_46013,N_46581);
xor U47594 (N_47594,N_47224,N_45439);
nand U47595 (N_47595,N_47016,N_46335);
nand U47596 (N_47596,N_47489,N_46775);
nor U47597 (N_47597,N_46163,N_47429);
and U47598 (N_47598,N_46081,N_46385);
and U47599 (N_47599,N_47373,N_46569);
and U47600 (N_47600,N_46837,N_47385);
xnor U47601 (N_47601,N_46752,N_45688);
and U47602 (N_47602,N_47388,N_46457);
or U47603 (N_47603,N_47426,N_45906);
nand U47604 (N_47604,N_46697,N_46037);
and U47605 (N_47605,N_45069,N_47143);
nor U47606 (N_47606,N_47355,N_46513);
xor U47607 (N_47607,N_46143,N_46772);
nor U47608 (N_47608,N_47114,N_47298);
nand U47609 (N_47609,N_45491,N_46483);
and U47610 (N_47610,N_45801,N_45670);
and U47611 (N_47611,N_45842,N_46800);
nor U47612 (N_47612,N_46698,N_47070);
nand U47613 (N_47613,N_47274,N_47076);
and U47614 (N_47614,N_45465,N_45054);
and U47615 (N_47615,N_45470,N_47495);
nand U47616 (N_47616,N_45004,N_47180);
or U47617 (N_47617,N_47130,N_45281);
or U47618 (N_47618,N_46212,N_45974);
or U47619 (N_47619,N_46641,N_47179);
or U47620 (N_47620,N_46076,N_46637);
nand U47621 (N_47621,N_46463,N_47225);
nand U47622 (N_47622,N_45843,N_47431);
nor U47623 (N_47623,N_45162,N_47235);
xor U47624 (N_47624,N_45396,N_46727);
xor U47625 (N_47625,N_46671,N_45821);
nor U47626 (N_47626,N_45473,N_45375);
nor U47627 (N_47627,N_45762,N_45418);
nor U47628 (N_47628,N_47208,N_45188);
or U47629 (N_47629,N_47250,N_46726);
nor U47630 (N_47630,N_46704,N_46370);
nand U47631 (N_47631,N_45988,N_45203);
nor U47632 (N_47632,N_47172,N_45888);
nor U47633 (N_47633,N_45154,N_45261);
and U47634 (N_47634,N_45689,N_46320);
nor U47635 (N_47635,N_46393,N_46495);
nor U47636 (N_47636,N_45613,N_45380);
xor U47637 (N_47637,N_46102,N_45433);
or U47638 (N_47638,N_46965,N_46147);
nor U47639 (N_47639,N_47343,N_46822);
xor U47640 (N_47640,N_46278,N_45969);
and U47641 (N_47641,N_45839,N_46128);
xor U47642 (N_47642,N_45043,N_45125);
nor U47643 (N_47643,N_45680,N_46362);
xnor U47644 (N_47644,N_45005,N_45981);
or U47645 (N_47645,N_47141,N_45662);
and U47646 (N_47646,N_47001,N_46958);
and U47647 (N_47647,N_46492,N_45106);
or U47648 (N_47648,N_47096,N_45268);
and U47649 (N_47649,N_45183,N_46509);
xor U47650 (N_47650,N_46557,N_46085);
and U47651 (N_47651,N_46676,N_47111);
nor U47652 (N_47652,N_47075,N_46524);
and U47653 (N_47653,N_45129,N_45373);
xor U47654 (N_47654,N_46559,N_47147);
or U47655 (N_47655,N_46932,N_46448);
nand U47656 (N_47656,N_46868,N_47450);
nand U47657 (N_47657,N_46911,N_45132);
xnor U47658 (N_47658,N_46976,N_47438);
and U47659 (N_47659,N_46589,N_47486);
or U47660 (N_47660,N_45939,N_46687);
and U47661 (N_47661,N_45951,N_46928);
xor U47662 (N_47662,N_46991,N_46753);
or U47663 (N_47663,N_45768,N_47073);
nand U47664 (N_47664,N_46160,N_47029);
xnor U47665 (N_47665,N_46804,N_46397);
nand U47666 (N_47666,N_46999,N_46801);
or U47667 (N_47667,N_45137,N_46952);
nand U47668 (N_47668,N_47344,N_45085);
nand U47669 (N_47669,N_45351,N_46731);
nor U47670 (N_47670,N_45847,N_45958);
xor U47671 (N_47671,N_47476,N_47318);
nand U47672 (N_47672,N_46023,N_46439);
and U47673 (N_47673,N_45128,N_47193);
nor U47674 (N_47674,N_45061,N_46152);
xor U47675 (N_47675,N_46438,N_46062);
and U47676 (N_47676,N_45798,N_47441);
xnor U47677 (N_47677,N_46445,N_47133);
nand U47678 (N_47678,N_45737,N_45828);
and U47679 (N_47679,N_47284,N_46433);
and U47680 (N_47680,N_46734,N_46180);
nand U47681 (N_47681,N_47047,N_47038);
or U47682 (N_47682,N_46073,N_47217);
or U47683 (N_47683,N_45500,N_45862);
nor U47684 (N_47684,N_45311,N_47214);
nor U47685 (N_47685,N_45378,N_47273);
and U47686 (N_47686,N_45257,N_47319);
nor U47687 (N_47687,N_45527,N_46904);
or U47688 (N_47688,N_46743,N_45479);
nor U47689 (N_47689,N_46137,N_47156);
xnor U47690 (N_47690,N_47050,N_45522);
nand U47691 (N_47691,N_46127,N_47202);
nor U47692 (N_47692,N_47167,N_46601);
and U47693 (N_47693,N_47240,N_45784);
and U47694 (N_47694,N_46856,N_46344);
nor U47695 (N_47695,N_45352,N_46898);
nor U47696 (N_47696,N_45113,N_46005);
nor U47697 (N_47697,N_45697,N_47322);
xnor U47698 (N_47698,N_46327,N_47149);
nand U47699 (N_47699,N_45467,N_45964);
and U47700 (N_47700,N_45791,N_47176);
nand U47701 (N_47701,N_46972,N_47213);
nor U47702 (N_47702,N_45708,N_47321);
nand U47703 (N_47703,N_46353,N_46926);
or U47704 (N_47704,N_45840,N_45363);
nor U47705 (N_47705,N_45770,N_45165);
nand U47706 (N_47706,N_46784,N_46294);
and U47707 (N_47707,N_45348,N_45018);
nor U47708 (N_47708,N_46339,N_46217);
xor U47709 (N_47709,N_46814,N_45437);
nand U47710 (N_47710,N_46452,N_46621);
nand U47711 (N_47711,N_46262,N_46201);
or U47712 (N_47712,N_47222,N_45691);
and U47713 (N_47713,N_45221,N_47412);
nand U47714 (N_47714,N_45793,N_45285);
xor U47715 (N_47715,N_47313,N_45645);
or U47716 (N_47716,N_47126,N_46269);
xnor U47717 (N_47717,N_47146,N_45992);
xnor U47718 (N_47718,N_45545,N_45436);
or U47719 (N_47719,N_46831,N_47371);
or U47720 (N_47720,N_46714,N_46069);
and U47721 (N_47721,N_46375,N_45075);
xnor U47722 (N_47722,N_45118,N_45323);
xor U47723 (N_47723,N_45283,N_46993);
and U47724 (N_47724,N_45759,N_45514);
nor U47725 (N_47725,N_45194,N_46603);
and U47726 (N_47726,N_45196,N_46434);
xnor U47727 (N_47727,N_45214,N_47245);
nand U47728 (N_47728,N_45742,N_46377);
or U47729 (N_47729,N_46626,N_45725);
or U47730 (N_47730,N_46883,N_47453);
nor U47731 (N_47731,N_47405,N_46732);
xor U47732 (N_47732,N_46711,N_46052);
and U47733 (N_47733,N_46110,N_46246);
or U47734 (N_47734,N_46144,N_46680);
nand U47735 (N_47735,N_45001,N_46834);
xnor U47736 (N_47736,N_45081,N_46650);
xor U47737 (N_47737,N_47369,N_45372);
nand U47738 (N_47738,N_46078,N_47366);
or U47739 (N_47739,N_47415,N_45153);
xor U47740 (N_47740,N_47090,N_46365);
nand U47741 (N_47741,N_45656,N_45448);
nor U47742 (N_47742,N_45528,N_46191);
nor U47743 (N_47743,N_46573,N_45468);
and U47744 (N_47744,N_45265,N_46717);
xnor U47745 (N_47745,N_46466,N_45779);
or U47746 (N_47746,N_47402,N_47042);
nand U47747 (N_47747,N_45937,N_46500);
and U47748 (N_47748,N_47353,N_47270);
xnor U47749 (N_47749,N_47332,N_45202);
nand U47750 (N_47750,N_47041,N_46855);
nor U47751 (N_47751,N_45661,N_45414);
or U47752 (N_47752,N_46040,N_45346);
and U47753 (N_47753,N_46488,N_45179);
nor U47754 (N_47754,N_45366,N_45702);
nor U47755 (N_47755,N_47471,N_46223);
nand U47756 (N_47756,N_46465,N_46813);
or U47757 (N_47757,N_45811,N_46550);
nor U47758 (N_47758,N_45101,N_46408);
nand U47759 (N_47759,N_45090,N_45634);
or U47760 (N_47760,N_46476,N_47478);
xor U47761 (N_47761,N_46888,N_47354);
or U47762 (N_47762,N_46759,N_45475);
xor U47763 (N_47763,N_46332,N_45250);
xnor U47764 (N_47764,N_46266,N_47361);
nor U47765 (N_47765,N_46899,N_46745);
nand U47766 (N_47766,N_46908,N_45191);
nor U47767 (N_47767,N_45699,N_46437);
and U47768 (N_47768,N_46876,N_45186);
nor U47769 (N_47769,N_47055,N_47155);
or U47770 (N_47770,N_46406,N_45819);
nand U47771 (N_47771,N_45388,N_45279);
or U47772 (N_47772,N_46877,N_45654);
nand U47773 (N_47773,N_45248,N_46693);
or U47774 (N_47774,N_45776,N_47238);
or U47775 (N_47775,N_45270,N_47323);
nand U47776 (N_47776,N_45216,N_45290);
xor U47777 (N_47777,N_45943,N_45082);
xor U47778 (N_47778,N_47234,N_45160);
nor U47779 (N_47779,N_46835,N_46471);
or U47780 (N_47780,N_45335,N_46526);
or U47781 (N_47781,N_45272,N_45289);
or U47782 (N_47782,N_46165,N_46473);
nand U47783 (N_47783,N_45857,N_46523);
and U47784 (N_47784,N_46022,N_45512);
and U47785 (N_47785,N_45723,N_45028);
nand U47786 (N_47786,N_45200,N_46134);
and U47787 (N_47787,N_45089,N_46394);
and U47788 (N_47788,N_47359,N_47456);
nand U47789 (N_47789,N_45629,N_45977);
or U47790 (N_47790,N_46967,N_45803);
and U47791 (N_47791,N_47472,N_46878);
xnor U47792 (N_47792,N_47307,N_46111);
xnor U47793 (N_47793,N_46087,N_46244);
nand U47794 (N_47794,N_46461,N_47434);
nand U47795 (N_47795,N_45995,N_46938);
nor U47796 (N_47796,N_47349,N_45576);
nand U47797 (N_47797,N_45837,N_45738);
nand U47798 (N_47798,N_47008,N_47315);
nor U47799 (N_47799,N_45136,N_47493);
nand U47800 (N_47800,N_46668,N_45387);
nor U47801 (N_47801,N_45157,N_46008);
xnor U47802 (N_47802,N_46516,N_45159);
or U47803 (N_47803,N_45073,N_46553);
nor U47804 (N_47804,N_45141,N_45934);
nand U47805 (N_47805,N_45956,N_47216);
nand U47806 (N_47806,N_45271,N_47305);
xor U47807 (N_47807,N_47086,N_46862);
and U47808 (N_47808,N_46120,N_45395);
and U47809 (N_47809,N_45239,N_46506);
and U47810 (N_47810,N_47432,N_46193);
xor U47811 (N_47811,N_46301,N_45155);
xnor U47812 (N_47812,N_46673,N_46199);
and U47813 (N_47813,N_46182,N_45584);
nor U47814 (N_47814,N_45880,N_46196);
nor U47815 (N_47815,N_46093,N_46885);
or U47816 (N_47816,N_47106,N_46916);
or U47817 (N_47817,N_45453,N_45487);
xnor U47818 (N_47818,N_46549,N_45423);
or U47819 (N_47819,N_45451,N_45369);
or U47820 (N_47820,N_47287,N_46207);
nand U47821 (N_47821,N_45480,N_47296);
nand U47822 (N_47822,N_47183,N_47324);
nand U47823 (N_47823,N_45682,N_45789);
or U47824 (N_47824,N_46275,N_45897);
nand U47825 (N_47825,N_45462,N_46994);
nand U47826 (N_47826,N_45959,N_45429);
xor U47827 (N_47827,N_46505,N_45556);
nand U47828 (N_47828,N_45703,N_45773);
or U47829 (N_47829,N_46805,N_45218);
and U47830 (N_47830,N_45790,N_46364);
and U47831 (N_47831,N_45059,N_47187);
nor U47832 (N_47832,N_47460,N_45151);
nand U47833 (N_47833,N_46934,N_46851);
or U47834 (N_47834,N_45318,N_45032);
nor U47835 (N_47835,N_47069,N_45663);
xnor U47836 (N_47836,N_45592,N_46762);
and U47837 (N_47837,N_45297,N_46011);
or U47838 (N_47838,N_46529,N_45651);
nor U47839 (N_47839,N_45447,N_45714);
or U47840 (N_47840,N_47443,N_45698);
nor U47841 (N_47841,N_46678,N_45313);
xor U47842 (N_47842,N_46226,N_46256);
nor U47843 (N_47843,N_45858,N_45961);
or U47844 (N_47844,N_45504,N_46215);
nand U47845 (N_47845,N_46340,N_46280);
nand U47846 (N_47846,N_45747,N_45097);
xnor U47847 (N_47847,N_46773,N_46351);
xor U47848 (N_47848,N_46691,N_45985);
nor U47849 (N_47849,N_46260,N_45523);
xnor U47850 (N_47850,N_45696,N_45275);
xor U47851 (N_47851,N_45940,N_46742);
nor U47852 (N_47852,N_45104,N_45339);
and U47853 (N_47853,N_47113,N_47089);
xor U47854 (N_47854,N_46902,N_46515);
and U47855 (N_47855,N_47162,N_45945);
nand U47856 (N_47856,N_45152,N_45397);
xor U47857 (N_47857,N_47046,N_46287);
and U47858 (N_47858,N_45901,N_47399);
nand U47859 (N_47859,N_45360,N_47056);
or U47860 (N_47860,N_46305,N_45233);
xnor U47861 (N_47861,N_45302,N_46540);
xor U47862 (N_47862,N_45677,N_46389);
or U47863 (N_47863,N_46741,N_46444);
xnor U47864 (N_47864,N_46489,N_45659);
nand U47865 (N_47865,N_45124,N_45262);
nor U47866 (N_47866,N_46625,N_45123);
xnor U47867 (N_47867,N_45300,N_45006);
xor U47868 (N_47868,N_45833,N_47446);
or U47869 (N_47869,N_46624,N_46295);
xnor U47870 (N_47870,N_47457,N_46200);
nand U47871 (N_47871,N_45099,N_45802);
nor U47872 (N_47872,N_47269,N_46996);
or U47873 (N_47873,N_46257,N_46190);
and U47874 (N_47874,N_47380,N_45600);
nand U47875 (N_47875,N_46227,N_45797);
nor U47876 (N_47876,N_47205,N_46818);
and U47877 (N_47877,N_46643,N_45147);
xor U47878 (N_47878,N_46481,N_45169);
nand U47879 (N_47879,N_45930,N_46783);
or U47880 (N_47880,N_46857,N_45119);
nand U47881 (N_47881,N_45450,N_47455);
xor U47882 (N_47882,N_46517,N_45383);
xor U47883 (N_47883,N_46322,N_45385);
and U47884 (N_47884,N_45210,N_45850);
or U47885 (N_47885,N_45307,N_45881);
nor U47886 (N_47886,N_46388,N_45301);
nand U47887 (N_47887,N_46520,N_47498);
nand U47888 (N_47888,N_46084,N_45066);
nand U47889 (N_47889,N_47158,N_47278);
or U47890 (N_47890,N_45516,N_46718);
nand U47891 (N_47891,N_46373,N_47157);
or U47892 (N_47892,N_46462,N_45317);
xnor U47893 (N_47893,N_46684,N_45693);
or U47894 (N_47894,N_46121,N_45185);
and U47895 (N_47895,N_45319,N_46619);
nor U47896 (N_47896,N_47283,N_45976);
nor U47897 (N_47897,N_45970,N_47376);
nor U47898 (N_47898,N_46455,N_47221);
and U47899 (N_47899,N_46749,N_45384);
or U47900 (N_47900,N_45841,N_45550);
xor U47901 (N_47901,N_45587,N_45225);
and U47902 (N_47902,N_46176,N_45569);
and U47903 (N_47903,N_45359,N_46158);
xor U47904 (N_47904,N_46648,N_45065);
or U47905 (N_47905,N_46705,N_47139);
and U47906 (N_47906,N_46797,N_45243);
xor U47907 (N_47907,N_45460,N_45161);
xor U47908 (N_47908,N_46887,N_46386);
and U47909 (N_47909,N_46041,N_47483);
and U47910 (N_47910,N_46175,N_47362);
xor U47911 (N_47911,N_46949,N_45483);
nor U47912 (N_47912,N_46203,N_46521);
nand U47913 (N_47913,N_45941,N_46145);
and U47914 (N_47914,N_45944,N_45368);
or U47915 (N_47915,N_46556,N_45813);
or U47916 (N_47916,N_45195,N_45390);
or U47917 (N_47917,N_45331,N_45932);
or U47918 (N_47918,N_46004,N_46108);
and U47919 (N_47919,N_46003,N_46507);
xor U47920 (N_47920,N_45076,N_46613);
nor U47921 (N_47921,N_45612,N_45253);
nand U47922 (N_47922,N_46681,N_45973);
nor U47923 (N_47923,N_45209,N_45679);
nor U47924 (N_47924,N_45394,N_45519);
and U47925 (N_47925,N_45260,N_46341);
xnor U47926 (N_47926,N_45478,N_45845);
nor U47927 (N_47927,N_45506,N_45795);
and U47928 (N_47928,N_46432,N_46347);
or U47929 (N_47929,N_45000,N_47033);
xnor U47930 (N_47930,N_47071,N_46995);
and U47931 (N_47931,N_45706,N_45484);
nand U47932 (N_47932,N_47062,N_46910);
nor U47933 (N_47933,N_45357,N_45362);
and U47934 (N_47934,N_45911,N_46115);
and U47935 (N_47935,N_45950,N_46006);
nand U47936 (N_47936,N_45533,N_47247);
nand U47937 (N_47937,N_46014,N_45347);
nand U47938 (N_47938,N_45649,N_45477);
nand U47939 (N_47939,N_45540,N_46148);
nand U47940 (N_47940,N_46164,N_47057);
nand U47941 (N_47941,N_46774,N_46844);
and U47942 (N_47942,N_46836,N_47254);
nor U47943 (N_47943,N_45534,N_47484);
nand U47944 (N_47944,N_47215,N_45139);
nand U47945 (N_47945,N_45343,N_46729);
nand U47946 (N_47946,N_45879,N_45055);
nor U47947 (N_47947,N_46962,N_47427);
nand U47948 (N_47948,N_47226,N_46334);
nand U47949 (N_47949,N_46532,N_46826);
and U47950 (N_47950,N_45120,N_46044);
xor U47951 (N_47951,N_46138,N_46400);
or U47952 (N_47952,N_45176,N_46874);
xnor U47953 (N_47953,N_45720,N_47473);
nand U47954 (N_47954,N_46527,N_46485);
nor U47955 (N_47955,N_45921,N_47236);
xnor U47956 (N_47956,N_46872,N_47011);
and U47957 (N_47957,N_47281,N_45716);
xor U47958 (N_47958,N_45783,N_46982);
nor U47959 (N_47959,N_47347,N_45598);
xor U47960 (N_47960,N_45909,N_45608);
nor U47961 (N_47961,N_46746,N_45227);
nor U47962 (N_47962,N_45952,N_47246);
nand U47963 (N_47963,N_46422,N_47346);
nor U47964 (N_47964,N_46931,N_47195);
nand U47965 (N_47965,N_46679,N_46618);
nor U47966 (N_47966,N_45715,N_45398);
and U47967 (N_47967,N_45367,N_46608);
xnor U47968 (N_47968,N_46204,N_46615);
nand U47969 (N_47969,N_45848,N_47068);
xor U47970 (N_47970,N_46418,N_46858);
or U47971 (N_47971,N_46059,N_46414);
nand U47972 (N_47972,N_45602,N_46989);
nand U47973 (N_47973,N_45400,N_46330);
nand U47974 (N_47974,N_45482,N_45681);
and U47975 (N_47975,N_47109,N_45652);
or U47976 (N_47976,N_45875,N_46906);
nor U47977 (N_47977,N_47403,N_47252);
nand U47978 (N_47978,N_45012,N_46025);
nand U47979 (N_47979,N_45560,N_46209);
and U47980 (N_47980,N_47459,N_46978);
or U47981 (N_47981,N_45008,N_45426);
or U47982 (N_47982,N_46066,N_46380);
xor U47983 (N_47983,N_46833,N_45409);
nand U47984 (N_47984,N_47014,N_45094);
xnor U47985 (N_47985,N_45276,N_45834);
xnor U47986 (N_47986,N_46828,N_46029);
nand U47987 (N_47987,N_46829,N_45805);
nand U47988 (N_47988,N_47101,N_45226);
or U47989 (N_47989,N_45083,N_45030);
xnor U47990 (N_47990,N_46538,N_46293);
or U47991 (N_47991,N_46788,N_45579);
xnor U47992 (N_47992,N_47060,N_46853);
and U47993 (N_47993,N_46969,N_45167);
and U47994 (N_47994,N_45886,N_45135);
nor U47995 (N_47995,N_45341,N_45316);
xor U47996 (N_47996,N_45107,N_45810);
or U47997 (N_47997,N_46270,N_45643);
nor U47998 (N_47998,N_47367,N_47003);
or U47999 (N_47999,N_46131,N_45566);
nor U48000 (N_48000,N_45029,N_45771);
xnor U48001 (N_48001,N_46942,N_45274);
nand U48002 (N_48002,N_45891,N_46054);
nor U48003 (N_48003,N_47301,N_47230);
xnor U48004 (N_48004,N_46083,N_45490);
nand U48005 (N_48005,N_46924,N_46597);
or U48006 (N_48006,N_45434,N_46747);
nor U48007 (N_48007,N_45168,N_46764);
xor U48008 (N_48008,N_46548,N_46017);
nand U48009 (N_48009,N_45053,N_47386);
xor U48010 (N_48010,N_45105,N_46761);
or U48011 (N_48011,N_45144,N_47439);
nor U48012 (N_48012,N_46068,N_47282);
and U48013 (N_48013,N_46825,N_47198);
xor U48014 (N_48014,N_45855,N_47077);
nand U48015 (N_48015,N_46161,N_45269);
xnor U48016 (N_48016,N_46395,N_46909);
or U48017 (N_48017,N_45709,N_46725);
nand U48018 (N_48018,N_47059,N_46470);
and U48019 (N_48019,N_46543,N_46900);
xor U48020 (N_48020,N_47078,N_46518);
nand U48021 (N_48021,N_45047,N_45023);
nor U48022 (N_48022,N_45249,N_45427);
xnor U48023 (N_48023,N_45374,N_45324);
and U48024 (N_48024,N_46645,N_45638);
nand U48025 (N_48025,N_46474,N_47242);
nor U48026 (N_48026,N_47088,N_45596);
and U48027 (N_48027,N_46346,N_46355);
or U48028 (N_48028,N_45904,N_45382);
nor U48029 (N_48029,N_45336,N_45349);
nor U48030 (N_48030,N_46359,N_46812);
and U48031 (N_48031,N_45887,N_45442);
and U48032 (N_48032,N_45539,N_46261);
nor U48033 (N_48033,N_46796,N_45966);
nand U48034 (N_48034,N_45876,N_46939);
xor U48035 (N_48035,N_46917,N_46970);
and U48036 (N_48036,N_46033,N_47334);
nand U48037 (N_48037,N_46968,N_46157);
or U48038 (N_48038,N_46091,N_46186);
xnor U48039 (N_48039,N_47173,N_46667);
or U48040 (N_48040,N_45846,N_46504);
xnor U48041 (N_48041,N_46806,N_47465);
or U48042 (N_48042,N_45224,N_45430);
xnor U48043 (N_48043,N_45215,N_46699);
nand U48044 (N_48044,N_45998,N_46415);
nand U48045 (N_48045,N_47206,N_45298);
nand U48046 (N_48046,N_46220,N_46129);
and U48047 (N_48047,N_45256,N_47186);
or U48048 (N_48048,N_47333,N_46379);
or U48049 (N_48049,N_46343,N_45780);
nor U48050 (N_48050,N_45717,N_46162);
nor U48051 (N_48051,N_47480,N_46750);
nor U48052 (N_48052,N_45700,N_46135);
xnor U48053 (N_48053,N_47189,N_45870);
nor U48054 (N_48054,N_47374,N_45775);
nand U48055 (N_48055,N_45361,N_46484);
xnor U48056 (N_48056,N_47150,N_45095);
nand U48057 (N_48057,N_47448,N_46089);
xnor U48058 (N_48058,N_45198,N_46689);
and U48059 (N_48059,N_45174,N_46250);
nand U48060 (N_48060,N_45744,N_46503);
nor U48061 (N_48061,N_46567,N_46021);
xnor U48062 (N_48062,N_46631,N_45619);
nor U48063 (N_48063,N_45530,N_45417);
nor U48064 (N_48064,N_46398,N_45822);
and U48065 (N_48065,N_45710,N_45864);
xor U48066 (N_48066,N_46591,N_46889);
xor U48067 (N_48067,N_46634,N_45752);
or U48068 (N_48068,N_47132,N_47048);
xnor U48069 (N_48069,N_45851,N_47419);
and U48070 (N_48070,N_46584,N_46382);
or U48071 (N_48071,N_46617,N_47009);
and U48072 (N_48072,N_46348,N_45309);
and U48073 (N_48073,N_45379,N_45595);
or U48074 (N_48074,N_46169,N_45518);
and U48075 (N_48075,N_45084,N_46151);
nand U48076 (N_48076,N_46823,N_46421);
and U48077 (N_48077,N_46113,N_46907);
nor U48078 (N_48078,N_47051,N_46990);
xnor U48079 (N_48079,N_47462,N_47308);
nand U48080 (N_48080,N_46297,N_46943);
nor U48081 (N_48081,N_46150,N_46281);
nand U48082 (N_48082,N_45282,N_46047);
xnor U48083 (N_48083,N_45912,N_47466);
nand U48084 (N_48084,N_45639,N_47067);
nand U48085 (N_48085,N_46058,N_45799);
xnor U48086 (N_48086,N_45838,N_45072);
or U48087 (N_48087,N_45068,N_46702);
or U48088 (N_48088,N_46233,N_47072);
nand U48089 (N_48089,N_45080,N_45893);
and U48090 (N_48090,N_45568,N_46696);
nor U48091 (N_48091,N_46112,N_46061);
xnor U48092 (N_48092,N_45815,N_46585);
nand U48093 (N_48093,N_45204,N_45365);
and U48094 (N_48094,N_45338,N_46633);
and U48095 (N_48095,N_46443,N_47030);
nor U48096 (N_48096,N_45278,N_46616);
nand U48097 (N_48097,N_46708,N_45295);
and U48098 (N_48098,N_45606,N_45178);
or U48099 (N_48099,N_46564,N_46819);
xnor U48100 (N_48100,N_45386,N_46237);
or U48101 (N_48101,N_45408,N_47125);
or U48102 (N_48102,N_46064,N_45989);
xnor U48103 (N_48103,N_45320,N_46787);
nor U48104 (N_48104,N_47134,N_46240);
nand U48105 (N_48105,N_47018,N_45117);
nor U48106 (N_48106,N_45878,N_45683);
nor U48107 (N_48107,N_47108,N_46399);
nor U48108 (N_48108,N_45403,N_45406);
or U48109 (N_48109,N_47211,N_45980);
or U48110 (N_48110,N_47017,N_46587);
or U48111 (N_48111,N_46168,N_46580);
xnor U48112 (N_48112,N_45647,N_45471);
and U48113 (N_48113,N_45108,N_45807);
nor U48114 (N_48114,N_45655,N_46771);
nand U48115 (N_48115,N_46265,N_45007);
xnor U48116 (N_48116,N_45003,N_47223);
nor U48117 (N_48117,N_45605,N_46477);
or U48118 (N_48118,N_46614,N_46665);
xnor U48119 (N_48119,N_46436,N_46722);
and U48120 (N_48120,N_46396,N_47023);
xnor U48121 (N_48121,N_45424,N_46225);
xnor U48122 (N_48122,N_46241,N_45149);
nand U48123 (N_48123,N_46785,N_46595);
xnor U48124 (N_48124,N_46019,N_46623);
nand U48125 (N_48125,N_46602,N_45449);
and U48126 (N_48126,N_45892,N_46230);
or U48127 (N_48127,N_47168,N_46622);
and U48128 (N_48128,N_47256,N_45525);
nand U48129 (N_48129,N_45133,N_45695);
nor U48130 (N_48130,N_46469,N_46053);
xor U48131 (N_48131,N_47260,N_45955);
xor U48132 (N_48132,N_47297,N_45488);
and U48133 (N_48133,N_45713,N_46658);
and U48134 (N_48134,N_46317,N_45990);
xor U48135 (N_48135,N_47259,N_45753);
nor U48136 (N_48136,N_46366,N_46213);
xnor U48137 (N_48137,N_46579,N_46001);
nor U48138 (N_48138,N_45578,N_46192);
nand U48139 (N_48139,N_47210,N_46922);
and U48140 (N_48140,N_45163,N_47171);
xnor U48141 (N_48141,N_47317,N_45495);
nand U48142 (N_48142,N_46211,N_47227);
nor U48143 (N_48143,N_45733,N_46036);
nand U48144 (N_48144,N_46728,N_47122);
xor U48145 (N_48145,N_45267,N_46803);
nand U48146 (N_48146,N_45583,N_47420);
nand U48147 (N_48147,N_46170,N_47474);
or U48148 (N_48148,N_47267,N_47095);
nand U48149 (N_48149,N_47378,N_45393);
and U48150 (N_48150,N_47110,N_45580);
and U48151 (N_48151,N_47194,N_46519);
and U48152 (N_48152,N_47174,N_45756);
nor U48153 (N_48153,N_46086,N_45321);
and U48154 (N_48154,N_45245,N_45074);
xor U48155 (N_48155,N_45907,N_46568);
nor U48156 (N_48156,N_47237,N_45520);
xnor U48157 (N_48157,N_47049,N_46815);
nor U48158 (N_48158,N_47435,N_47339);
xor U48159 (N_48159,N_46663,N_45381);
nor U48160 (N_48160,N_45729,N_46070);
nor U48161 (N_48161,N_47348,N_47181);
nand U48162 (N_48162,N_46007,N_46456);
xor U48163 (N_48163,N_45158,N_45509);
or U48164 (N_48164,N_45885,N_45920);
nand U48165 (N_48165,N_46720,N_47082);
nand U48166 (N_48166,N_45236,N_45922);
nor U48167 (N_48167,N_45062,N_45505);
xor U48168 (N_48168,N_45957,N_45122);
nor U48169 (N_48169,N_45098,N_45631);
nor U48170 (N_48170,N_47477,N_45919);
nand U48171 (N_48171,N_46546,N_46105);
or U48172 (N_48172,N_45057,N_45337);
or U48173 (N_48173,N_46933,N_47019);
nor U48174 (N_48174,N_46288,N_46838);
or U48175 (N_48175,N_46045,N_46832);
nand U48176 (N_48176,N_46530,N_46930);
and U48177 (N_48177,N_45814,N_47368);
nor U48178 (N_48178,N_46491,N_46048);
nand U48179 (N_48179,N_45705,N_45804);
and U48180 (N_48180,N_45678,N_45786);
xnor U48181 (N_48181,N_46154,N_45399);
or U48182 (N_48182,N_46416,N_46963);
or U48183 (N_48183,N_47451,N_45630);
nand U48184 (N_48184,N_46811,N_45284);
nor U48185 (N_48185,N_45035,N_45499);
xnor U48186 (N_48186,N_46172,N_47026);
nor U48187 (N_48187,N_47398,N_46117);
or U48188 (N_48188,N_47043,N_47007);
or U48189 (N_48189,N_47218,N_46555);
nor U48190 (N_48190,N_45831,N_46539);
nor U48191 (N_48191,N_45806,N_45558);
nand U48192 (N_48192,N_47081,N_46426);
or U48193 (N_48193,N_47401,N_46228);
xor U48194 (N_48194,N_46871,N_46088);
nand U48195 (N_48195,N_45739,N_45537);
and U48196 (N_48196,N_45975,N_46074);
nor U48197 (N_48197,N_46423,N_46997);
and U48198 (N_48198,N_45048,N_45052);
nand U48199 (N_48199,N_47228,N_45542);
xor U48200 (N_48200,N_45740,N_45788);
and U48201 (N_48201,N_45997,N_45190);
or U48202 (N_48202,N_45287,N_45371);
xor U48203 (N_48203,N_45428,N_46809);
or U48204 (N_48204,N_46560,N_45734);
and U48205 (N_48205,N_47191,N_45766);
nor U48206 (N_48206,N_46610,N_46194);
and U48207 (N_48207,N_45077,N_47006);
nand U48208 (N_48208,N_46757,N_46827);
or U48209 (N_48209,N_46309,N_47079);
xnor U48210 (N_48210,N_45926,N_47291);
nor U48211 (N_48211,N_46988,N_47015);
nand U48212 (N_48212,N_45597,N_46973);
and U48213 (N_48213,N_45622,N_46042);
or U48214 (N_48214,N_46502,N_45627);
and U48215 (N_48215,N_47127,N_45987);
xnor U48216 (N_48216,N_46736,N_47357);
nor U48217 (N_48217,N_46123,N_46884);
or U48218 (N_48218,N_47492,N_45895);
and U48219 (N_48219,N_45929,N_46807);
nor U48220 (N_48220,N_46879,N_47306);
nor U48221 (N_48221,N_46535,N_45148);
or U48222 (N_48222,N_46371,N_46738);
xnor U48223 (N_48223,N_47053,N_45593);
nand U48224 (N_48224,N_45060,N_45481);
xnor U48225 (N_48225,N_45498,N_45150);
nor U48226 (N_48226,N_46572,N_46401);
nand U48227 (N_48227,N_45131,N_46733);
and U48228 (N_48228,N_45303,N_45633);
or U48229 (N_48229,N_46323,N_46570);
and U48230 (N_48230,N_45551,N_45914);
and U48231 (N_48231,N_47425,N_45874);
nand U48232 (N_48232,N_45241,N_46232);
or U48233 (N_48233,N_47120,N_46118);
or U48234 (N_48234,N_46744,N_46252);
xor U48235 (N_48235,N_47437,N_45621);
nand U48236 (N_48236,N_46031,N_45446);
or U48237 (N_48237,N_45704,N_47391);
or U48238 (N_48238,N_46890,N_45707);
xor U48239 (N_48239,N_45049,N_45016);
xor U48240 (N_48240,N_46331,N_46611);
xnor U48241 (N_48241,N_45757,N_47279);
nor U48242 (N_48242,N_47105,N_45164);
and U48243 (N_48243,N_45389,N_45982);
nor U48244 (N_48244,N_45761,N_45825);
xnor U48245 (N_48245,N_45686,N_47005);
or U48246 (N_48246,N_45936,N_46222);
or U48247 (N_48247,N_46864,N_45787);
nand U48248 (N_48248,N_46060,N_45999);
and U48249 (N_48249,N_45724,N_46106);
or U48250 (N_48250,N_46337,N_47175);
or U48251 (N_48251,N_47263,N_45501);
nand U48252 (N_48252,N_45315,N_45058);
xnor U48253 (N_48253,N_45749,N_45641);
nand U48254 (N_48254,N_45454,N_46403);
xor U48255 (N_48255,N_45103,N_47392);
or U48256 (N_48256,N_46715,N_45420);
and U48257 (N_48257,N_46234,N_46501);
or U48258 (N_48258,N_46153,N_45238);
or U48259 (N_48259,N_45173,N_46542);
xor U48260 (N_48260,N_46413,N_47024);
nand U48261 (N_48261,N_46277,N_46435);
or U48262 (N_48262,N_45140,N_45304);
nor U48263 (N_48263,N_45452,N_45296);
or U48264 (N_48264,N_46311,N_46302);
xor U48265 (N_48265,N_45532,N_46245);
and U48266 (N_48266,N_46381,N_46867);
and U48267 (N_48267,N_45404,N_45288);
nor U48268 (N_48268,N_45967,N_46854);
and U48269 (N_48269,N_47377,N_45355);
and U48270 (N_48270,N_46912,N_47394);
xnor U48271 (N_48271,N_46367,N_45096);
or U48272 (N_48272,N_46239,N_47295);
or U48273 (N_48273,N_46565,N_45247);
and U48274 (N_48274,N_46430,N_47092);
nor U48275 (N_48275,N_47239,N_46630);
nor U48276 (N_48276,N_46586,N_46850);
nand U48277 (N_48277,N_45735,N_46303);
or U48278 (N_48278,N_47207,N_46472);
xor U48279 (N_48279,N_47012,N_46487);
or U48280 (N_48280,N_46998,N_47037);
xnor U48281 (N_48281,N_46098,N_45416);
xnor U48282 (N_48282,N_46314,N_46646);
nand U48283 (N_48283,N_45544,N_45251);
or U48284 (N_48284,N_45358,N_46284);
nand U48285 (N_48285,N_45599,N_45549);
nand U48286 (N_48286,N_46358,N_45938);
or U48287 (N_48287,N_45925,N_45354);
or U48288 (N_48288,N_45644,N_47103);
nand U48289 (N_48289,N_46578,N_45344);
xnor U48290 (N_48290,N_45971,N_46961);
nor U48291 (N_48291,N_46142,N_45986);
nand U48292 (N_48292,N_46315,N_46268);
or U48293 (N_48293,N_46177,N_45615);
or U48294 (N_48294,N_45252,N_46271);
xnor U48295 (N_48295,N_46966,N_45601);
xnor U48296 (N_48296,N_46946,N_46839);
nand U48297 (N_48297,N_47470,N_46378);
xnor U48298 (N_48298,N_46983,N_46383);
or U48299 (N_48299,N_45590,N_45277);
nand U48300 (N_48300,N_46824,N_46405);
or U48301 (N_48301,N_45325,N_45356);
and U48302 (N_48302,N_45046,N_47454);
xnor U48303 (N_48303,N_45350,N_47325);
and U48304 (N_48304,N_45181,N_45626);
xnor U48305 (N_48305,N_47330,N_46941);
nor U48306 (N_48306,N_45623,N_45535);
nand U48307 (N_48307,N_46310,N_47121);
nand U48308 (N_48308,N_45743,N_47316);
and U48309 (N_48309,N_47107,N_45322);
nor U48310 (N_48310,N_46279,N_47257);
and U48311 (N_48311,N_46000,N_46449);
or U48312 (N_48312,N_46675,N_45965);
or U48313 (N_48313,N_46628,N_45508);
or U48314 (N_48314,N_45306,N_45013);
or U48315 (N_48315,N_46954,N_45719);
or U48316 (N_48316,N_46674,N_46588);
or U48317 (N_48317,N_45675,N_45574);
xor U48318 (N_48318,N_46627,N_46778);
xor U48319 (N_48319,N_47165,N_47244);
and U48320 (N_48320,N_45564,N_45687);
or U48321 (N_48321,N_45658,N_45497);
nor U48322 (N_48322,N_47356,N_46038);
or U48323 (N_48323,N_45616,N_45088);
nand U48324 (N_48324,N_46642,N_45254);
nor U48325 (N_48325,N_46582,N_46852);
and U48326 (N_48326,N_46107,N_46984);
xnor U48327 (N_48327,N_47370,N_45067);
xor U48328 (N_48328,N_46420,N_46140);
xnor U48329 (N_48329,N_45042,N_47275);
xor U48330 (N_48330,N_45588,N_46886);
and U48331 (N_48331,N_46703,N_47300);
nand U48332 (N_48332,N_45444,N_45555);
nand U48333 (N_48333,N_47337,N_45617);
and U48334 (N_48334,N_45746,N_45728);
and U48335 (N_48335,N_45310,N_47463);
and U48336 (N_48336,N_47482,N_45684);
xnor U48337 (N_48337,N_45563,N_45146);
xor U48338 (N_48338,N_47177,N_46735);
nor U48339 (N_48339,N_46847,N_45445);
nor U48340 (N_48340,N_47276,N_45334);
or U48341 (N_48341,N_45486,N_45100);
and U48342 (N_48342,N_46286,N_46299);
or U48343 (N_48343,N_46338,N_45800);
and U48344 (N_48344,N_45212,N_46357);
nor U48345 (N_48345,N_47487,N_46075);
nor U48346 (N_48346,N_46936,N_46870);
or U48347 (N_48347,N_46779,N_46126);
nor U48348 (N_48348,N_45207,N_47341);
and U48349 (N_48349,N_45370,N_46412);
nor U48350 (N_48350,N_47190,N_45949);
and U48351 (N_48351,N_46092,N_45758);
xnor U48352 (N_48352,N_46701,N_46905);
nand U48353 (N_48353,N_46959,N_46057);
or U48354 (N_48354,N_47433,N_46985);
nand U48355 (N_48355,N_45931,N_47148);
nor U48356 (N_48356,N_45228,N_47102);
and U48357 (N_48357,N_45760,N_46508);
and U48358 (N_48358,N_46368,N_45292);
and U48359 (N_48359,N_45859,N_45180);
xor U48360 (N_48360,N_46243,N_47382);
xor U48361 (N_48361,N_46055,N_45201);
xnor U48362 (N_48362,N_45900,N_46974);
xor U48363 (N_48363,N_46119,N_46183);
xor U48364 (N_48364,N_45237,N_47124);
nand U48365 (N_48365,N_45342,N_46141);
and U48366 (N_48366,N_45994,N_45765);
nand U48367 (N_48367,N_45625,N_47039);
or U48368 (N_48368,N_45246,N_46419);
nand U48369 (N_48369,N_47413,N_46953);
nor U48370 (N_48370,N_46574,N_45827);
and U48371 (N_48371,N_47396,N_47271);
nor U48372 (N_48372,N_47299,N_47490);
nor U48373 (N_48373,N_46793,N_46756);
nand U48374 (N_48374,N_45860,N_45111);
nand U48375 (N_48375,N_46125,N_45667);
xor U48376 (N_48376,N_47137,N_47229);
or U48377 (N_48377,N_46547,N_46325);
nor U48378 (N_48378,N_46893,N_45611);
or U48379 (N_48379,N_46575,N_45438);
or U48380 (N_48380,N_46263,N_45222);
or U48381 (N_48381,N_46786,N_45435);
nor U48382 (N_48382,N_45868,N_45730);
nand U48383 (N_48383,N_45037,N_46639);
nand U48384 (N_48384,N_45711,N_47140);
xnor U48385 (N_48385,N_45112,N_46427);
nor U48386 (N_48386,N_46955,N_47302);
xor U48387 (N_48387,N_45573,N_46475);
or U48388 (N_48388,N_46981,N_47201);
nor U48389 (N_48389,N_46155,N_46224);
nor U48390 (N_48390,N_46605,N_45138);
or U48391 (N_48391,N_46424,N_46755);
nand U48392 (N_48392,N_46781,N_47400);
nor U48393 (N_48393,N_45223,N_46326);
and U48394 (N_48394,N_46975,N_45721);
and U48395 (N_48395,N_45856,N_46298);
nor U48396 (N_48396,N_47154,N_46345);
xor U48397 (N_48397,N_46740,N_45193);
or U48398 (N_48398,N_45496,N_46897);
xnor U48399 (N_48399,N_46723,N_46390);
nand U48400 (N_48400,N_46493,N_45421);
or U48401 (N_48401,N_47408,N_45040);
xor U48402 (N_48402,N_47375,N_46249);
and U48403 (N_48403,N_45182,N_47144);
nand U48404 (N_48404,N_47406,N_47255);
nor U48405 (N_48405,N_46034,N_47084);
xnor U48406 (N_48406,N_45515,N_45305);
nor U48407 (N_48407,N_46002,N_46480);
or U48408 (N_48408,N_47288,N_45996);
and U48409 (N_48409,N_46620,N_47326);
and U48410 (N_48410,N_45412,N_45778);
and U48411 (N_48411,N_45650,N_46935);
and U48412 (N_48412,N_45455,N_45469);
or U48413 (N_48413,N_46512,N_45559);
nor U48414 (N_48414,N_46713,N_47458);
and U48415 (N_48415,N_45494,N_46915);
nor U48416 (N_48416,N_45642,N_45582);
nand U48417 (N_48417,N_46319,N_46820);
xnor U48418 (N_48418,N_46374,N_46903);
xnor U48419 (N_48419,N_45902,N_47136);
nand U48420 (N_48420,N_46050,N_47040);
and U48421 (N_48421,N_46944,N_47310);
nand U48422 (N_48422,N_46097,N_47219);
xor U48423 (N_48423,N_47292,N_47129);
nor U48424 (N_48424,N_47212,N_46478);
nand U48425 (N_48425,N_46195,N_46914);
and U48426 (N_48426,N_45036,N_45890);
or U48427 (N_48427,N_45962,N_47390);
and U48428 (N_48428,N_45538,N_46318);
and U48429 (N_48429,N_45933,N_45660);
nor U48430 (N_48430,N_46533,N_45812);
nand U48431 (N_48431,N_46046,N_45440);
nor U48432 (N_48432,N_46409,N_47080);
nor U48433 (N_48433,N_46894,N_45829);
or U48434 (N_48434,N_46441,N_45792);
nor U48435 (N_48435,N_45968,N_45392);
and U48436 (N_48436,N_47159,N_45330);
and U48437 (N_48437,N_45946,N_45014);
or U48438 (N_48438,N_45489,N_45835);
nand U48439 (N_48439,N_45521,N_45726);
nand U48440 (N_48440,N_47097,N_45022);
xor U48441 (N_48441,N_45280,N_46682);
nand U48442 (N_48442,N_46015,N_47469);
nor U48443 (N_48443,N_45541,N_45794);
and U48444 (N_48444,N_46649,N_46896);
xnor U48445 (N_48445,N_45610,N_45872);
nor U48446 (N_48446,N_47231,N_47327);
or U48447 (N_48447,N_47488,N_47365);
nor U48448 (N_48448,N_45561,N_47182);
xnor U48449 (N_48449,N_46776,N_46384);
xor U48450 (N_48450,N_45905,N_46454);
nand U48451 (N_48451,N_47393,N_46536);
xnor U48452 (N_48452,N_45589,N_45328);
nand U48453 (N_48453,N_46782,N_46799);
xnor U48454 (N_48454,N_45314,N_47328);
nand U48455 (N_48455,N_46431,N_45767);
nand U48456 (N_48456,N_46313,N_46352);
xnor U48457 (N_48457,N_46522,N_46429);
nand U48458 (N_48458,N_45091,N_46647);
nor U48459 (N_48459,N_47163,N_46986);
xor U48460 (N_48460,N_45493,N_45126);
nand U48461 (N_48461,N_47098,N_47261);
xnor U48462 (N_48462,N_46636,N_45882);
nor U48463 (N_48463,N_45823,N_45266);
nand U48464 (N_48464,N_45517,N_46349);
or U48465 (N_48465,N_45419,N_45415);
nand U48466 (N_48466,N_45665,N_45960);
xnor U48467 (N_48467,N_45377,N_47360);
xor U48468 (N_48468,N_45963,N_47397);
nand U48469 (N_48469,N_46843,N_47119);
nor U48470 (N_48470,N_46173,N_46496);
or U48471 (N_48471,N_45017,N_47004);
and U48472 (N_48472,N_45443,N_47000);
xor U48473 (N_48473,N_46737,N_46082);
xnor U48474 (N_48474,N_47395,N_46205);
or U48475 (N_48475,N_45463,N_46960);
or U48476 (N_48476,N_46830,N_47100);
nor U48477 (N_48477,N_46683,N_46090);
and U48478 (N_48478,N_46754,N_45019);
xor U48479 (N_48479,N_45134,N_47293);
nand U48480 (N_48480,N_45009,N_45034);
or U48481 (N_48481,N_47099,N_46918);
nor U48482 (N_48482,N_47294,N_47335);
xnor U48483 (N_48483,N_47253,N_46447);
nor U48484 (N_48484,N_45754,N_47036);
nand U48485 (N_48485,N_46688,N_45020);
nand U48486 (N_48486,N_45422,N_45543);
nand U48487 (N_48487,N_45869,N_45585);
nand U48488 (N_48488,N_46510,N_45554);
or U48489 (N_48489,N_45896,N_46980);
and U48490 (N_48490,N_45273,N_46758);
xnor U48491 (N_48491,N_47184,N_46604);
nand U48492 (N_48492,N_46342,N_46677);
or U48493 (N_48493,N_46598,N_45745);
nand U48494 (N_48494,N_45712,N_46920);
or U48495 (N_48495,N_46453,N_46114);
or U48496 (N_48496,N_45972,N_45026);
nand U48497 (N_48497,N_46149,N_47027);
nor U48498 (N_48498,N_46685,N_46402);
or U48499 (N_48499,N_45865,N_45513);
or U48500 (N_48500,N_46267,N_45458);
or U48501 (N_48501,N_46577,N_46221);
nand U48502 (N_48502,N_46464,N_47312);
xor U48503 (N_48503,N_45086,N_45299);
and U48504 (N_48504,N_47494,N_46187);
or U48505 (N_48505,N_47418,N_46817);
nor U48506 (N_48506,N_47142,N_47169);
nor U48507 (N_48507,N_45983,N_47138);
nand U48508 (N_48508,N_45476,N_45259);
xnor U48509 (N_48509,N_46264,N_45984);
nor U48510 (N_48510,N_46307,N_47233);
nand U48511 (N_48511,N_46124,N_45524);
nor U48512 (N_48512,N_46511,N_45570);
and U48513 (N_48513,N_46730,N_46558);
xor U48514 (N_48514,N_46869,N_46051);
or U48515 (N_48515,N_46020,N_46030);
or U48516 (N_48516,N_46296,N_45863);
and U48517 (N_48517,N_45326,N_47464);
nor U48518 (N_48518,N_46361,N_45769);
and U48519 (N_48519,N_45577,N_47497);
and U48520 (N_48520,N_46156,N_46460);
and U48521 (N_48521,N_47342,N_46525);
and U48522 (N_48522,N_46109,N_46919);
and U48523 (N_48523,N_45063,N_46328);
xnor U48524 (N_48524,N_47032,N_45722);
xnor U48525 (N_48525,N_45327,N_47021);
and U48526 (N_48526,N_46664,N_47094);
nor U48527 (N_48527,N_46700,N_46067);
xor U48528 (N_48528,N_45213,N_46600);
and U48529 (N_48529,N_46765,N_45170);
and U48530 (N_48530,N_47203,N_45391);
nor U48531 (N_48531,N_45041,N_45915);
nand U48532 (N_48532,N_46009,N_45866);
nand U48533 (N_48533,N_45572,N_45312);
or U48534 (N_48534,N_45187,N_46274);
or U48535 (N_48535,N_45459,N_45736);
or U48536 (N_48536,N_45565,N_47091);
nor U48537 (N_48537,N_47309,N_46808);
xor U48538 (N_48538,N_45640,N_47379);
and U48539 (N_48539,N_45694,N_47188);
or U48540 (N_48540,N_45051,N_47304);
xnor U48541 (N_48541,N_46391,N_46763);
xor U48542 (N_48542,N_46816,N_45666);
or U48543 (N_48543,N_46719,N_46607);
nand U48544 (N_48544,N_45333,N_46179);
xnor U48545 (N_48545,N_45591,N_46028);
and U48546 (N_48546,N_47199,N_46537);
or U48547 (N_48547,N_46467,N_45205);
and U48548 (N_48548,N_46657,N_46977);
nand U48549 (N_48549,N_47104,N_47452);
or U48550 (N_48550,N_46659,N_46925);
and U48551 (N_48551,N_45456,N_46545);
and U48552 (N_48552,N_46710,N_47467);
or U48553 (N_48553,N_47151,N_46103);
nor U48554 (N_48554,N_46669,N_47200);
nor U48555 (N_48555,N_46238,N_46712);
and U48556 (N_48556,N_46451,N_46780);
nor U48557 (N_48557,N_46333,N_46079);
and U48558 (N_48558,N_45464,N_47160);
and U48559 (N_48559,N_46214,N_46231);
and U48560 (N_48560,N_45401,N_47152);
and U48561 (N_48561,N_45731,N_45121);
xor U48562 (N_48562,N_45410,N_45294);
xnor U48563 (N_48563,N_46770,N_46236);
or U48564 (N_48564,N_47416,N_47442);
or U48565 (N_48565,N_46080,N_45618);
nor U48566 (N_48566,N_46417,N_45750);
xnor U48567 (N_48567,N_45913,N_45899);
or U48568 (N_48568,N_46450,N_46672);
nand U48569 (N_48569,N_47414,N_45871);
xor U48570 (N_48570,N_46247,N_45308);
nand U48571 (N_48571,N_45502,N_45244);
xor U48572 (N_48572,N_46308,N_46372);
or U48573 (N_48573,N_46446,N_45526);
nor U48574 (N_48574,N_46789,N_45332);
xnor U48575 (N_48575,N_45531,N_47449);
xnor U48576 (N_48576,N_45102,N_46259);
nor U48577 (N_48577,N_45852,N_46873);
or U48578 (N_48578,N_47135,N_45039);
and U48579 (N_48579,N_46694,N_45624);
and U48580 (N_48580,N_46248,N_45692);
and U48581 (N_48581,N_46095,N_45809);
xor U48582 (N_48582,N_45978,N_45836);
xnor U48583 (N_48583,N_45604,N_47241);
or U48584 (N_48584,N_46940,N_45636);
and U48585 (N_48585,N_46576,N_45263);
nand U48586 (N_48586,N_45064,N_45529);
nor U48587 (N_48587,N_47204,N_47131);
nor U48588 (N_48588,N_45510,N_47389);
and U48589 (N_48589,N_46594,N_46101);
xnor U48590 (N_48590,N_46534,N_46321);
nor U48591 (N_48591,N_45432,N_46146);
nand U48592 (N_48592,N_46690,N_47345);
nor U48593 (N_48593,N_45208,N_47383);
or U48594 (N_48594,N_47436,N_45948);
nand U48595 (N_48595,N_46312,N_45782);
xor U48596 (N_48596,N_46178,N_46541);
xor U48597 (N_48597,N_46410,N_46670);
nand U48598 (N_48598,N_46065,N_45031);
nor U48599 (N_48599,N_45175,N_46724);
and U48600 (N_48600,N_46992,N_46739);
nand U48601 (N_48601,N_46652,N_45402);
or U48602 (N_48602,N_46122,N_47338);
xor U48603 (N_48603,N_46571,N_46411);
nand U48604 (N_48604,N_45575,N_46139);
or U48605 (N_48605,N_46188,N_46760);
or U48606 (N_48606,N_45293,N_46769);
xnor U48607 (N_48607,N_46950,N_46821);
and U48608 (N_48608,N_47052,N_47116);
xnor U48609 (N_48609,N_46071,N_46219);
nand U48610 (N_48610,N_47407,N_46387);
xnor U48611 (N_48611,N_45177,N_45171);
xnor U48612 (N_48612,N_45620,N_47422);
nand U48613 (N_48613,N_47022,N_46072);
or U48614 (N_48614,N_47074,N_45142);
nand U48615 (N_48615,N_45197,N_47044);
nor U48616 (N_48616,N_47170,N_46593);
nand U48617 (N_48617,N_45092,N_45844);
or U48618 (N_48618,N_47421,N_45669);
and U48619 (N_48619,N_46181,N_45242);
or U48620 (N_48620,N_45917,N_45264);
and U48621 (N_48621,N_45425,N_45405);
and U48622 (N_48622,N_46635,N_45114);
and U48623 (N_48623,N_46798,N_46229);
xor U48624 (N_48624,N_46100,N_46947);
nor U48625 (N_48625,N_46692,N_46957);
and U48626 (N_48626,N_45536,N_46895);
nand U48627 (N_48627,N_45002,N_45991);
and U48628 (N_48628,N_46039,N_46354);
or U48629 (N_48629,N_45116,N_45189);
nand U48630 (N_48630,N_47031,N_47065);
and U48631 (N_48631,N_46276,N_45025);
xnor U48632 (N_48632,N_46632,N_46654);
or U48633 (N_48633,N_45571,N_47054);
nor U48634 (N_48634,N_45603,N_45109);
nand U48635 (N_48635,N_46661,N_47249);
xor U48636 (N_48636,N_46136,N_46964);
or U48637 (N_48637,N_45609,N_45830);
nor U48638 (N_48638,N_47085,N_45849);
nand U48639 (N_48639,N_47264,N_45235);
xnor U48640 (N_48640,N_45867,N_46104);
xor U48641 (N_48641,N_45045,N_46171);
and U48642 (N_48642,N_45229,N_47196);
nand U48643 (N_48643,N_46531,N_45143);
nor U48644 (N_48644,N_46458,N_47020);
or U48645 (N_48645,N_45903,N_45898);
nand U48646 (N_48646,N_46849,N_45353);
or U48647 (N_48647,N_46794,N_45234);
nand U48648 (N_48648,N_45671,N_47303);
nand U48649 (N_48649,N_46027,N_45586);
and U48650 (N_48650,N_45127,N_45145);
nand U48651 (N_48651,N_47444,N_46891);
nand U48652 (N_48652,N_45632,N_47485);
nand U48653 (N_48653,N_45796,N_46291);
and U48654 (N_48654,N_46063,N_47010);
nor U48655 (N_48655,N_46167,N_45883);
or U48656 (N_48656,N_45924,N_45230);
xor U48657 (N_48657,N_45873,N_45219);
or U48658 (N_48658,N_45466,N_47496);
xor U48659 (N_48659,N_46956,N_47290);
nand U48660 (N_48660,N_47358,N_45908);
nor U48661 (N_48661,N_46272,N_45718);
nor U48662 (N_48662,N_45413,N_46479);
xnor U48663 (N_48663,N_47314,N_47209);
xor U48664 (N_48664,N_47028,N_47061);
xor U48665 (N_48665,N_45979,N_46514);
xnor U48666 (N_48666,N_45877,N_46442);
and U48667 (N_48667,N_46921,N_46859);
xnor U48668 (N_48668,N_46590,N_47289);
and U48669 (N_48669,N_46324,N_46606);
and U48670 (N_48670,N_46707,N_46499);
nor U48671 (N_48671,N_45038,N_47277);
and U48672 (N_48672,N_45674,N_45826);
xor U48673 (N_48673,N_45916,N_46686);
nand U48674 (N_48674,N_47364,N_45942);
and U48675 (N_48675,N_45781,N_47447);
and U48676 (N_48676,N_47262,N_47351);
nand U48677 (N_48677,N_47445,N_46751);
nand U48678 (N_48678,N_46544,N_46099);
xnor U48679 (N_48679,N_45701,N_47423);
and U48680 (N_48680,N_45364,N_46865);
xor U48681 (N_48681,N_45614,N_46468);
nand U48682 (N_48682,N_47461,N_46660);
nor U48683 (N_48683,N_46486,N_45653);
or U48684 (N_48684,N_46329,N_45217);
xor U48685 (N_48685,N_47197,N_45329);
nand U48686 (N_48686,N_45673,N_45741);
or U48687 (N_48687,N_47268,N_46706);
or U48688 (N_48688,N_46166,N_46077);
or U48689 (N_48689,N_46210,N_46043);
nand U48690 (N_48690,N_46253,N_45772);
and U48691 (N_48691,N_46721,N_45763);
nand U48692 (N_48692,N_45021,N_47424);
or U48693 (N_48693,N_46282,N_46498);
xor U48694 (N_48694,N_45087,N_46255);
xnor U48695 (N_48695,N_45503,N_46290);
xor U48696 (N_48696,N_47384,N_47286);
nand U48697 (N_48697,N_45431,N_45923);
nor U48698 (N_48698,N_46945,N_45474);
xor U48699 (N_48699,N_47087,N_47153);
and U48700 (N_48700,N_47248,N_46254);
xnor U48701 (N_48701,N_46987,N_46551);
xor U48702 (N_48702,N_45935,N_45255);
nand U48703 (N_48703,N_45552,N_46360);
nor U48704 (N_48704,N_45947,N_45156);
nand U48705 (N_48705,N_45056,N_45441);
xnor U48706 (N_48706,N_46018,N_47115);
or U48707 (N_48707,N_47220,N_46929);
or U48708 (N_48708,N_46860,N_45774);
nand U48709 (N_48709,N_46369,N_45172);
nor U48710 (N_48710,N_45648,N_45927);
and U48711 (N_48711,N_45472,N_46927);
xor U48712 (N_48712,N_45010,N_45953);
nand U48713 (N_48713,N_45854,N_45894);
and U48714 (N_48714,N_46653,N_46640);
xnor U48715 (N_48715,N_45044,N_46596);
nand U48716 (N_48716,N_46880,N_45345);
nand U48717 (N_48717,N_47243,N_45211);
nor U48718 (N_48718,N_46882,N_46866);
xnor U48719 (N_48719,N_45732,N_45376);
and U48720 (N_48720,N_46552,N_47266);
or U48721 (N_48721,N_46198,N_46490);
nor U48722 (N_48722,N_45581,N_46842);
xnor U48723 (N_48723,N_46599,N_46777);
or U48724 (N_48724,N_47063,N_47112);
or U48725 (N_48725,N_45818,N_47002);
nand U48726 (N_48726,N_47331,N_46638);
and U48727 (N_48727,N_46923,N_45928);
and U48728 (N_48728,N_47118,N_47178);
nor U48729 (N_48729,N_45755,N_46350);
or U48730 (N_48730,N_46846,N_46425);
and U48731 (N_48731,N_46841,N_45853);
nor U48732 (N_48732,N_45078,N_46609);
or U48733 (N_48733,N_46189,N_45015);
nand U48734 (N_48734,N_46132,N_47185);
or U48735 (N_48735,N_45993,N_45231);
or U48736 (N_48736,N_47430,N_46791);
or U48737 (N_48737,N_46392,N_47265);
nor U48738 (N_48738,N_45861,N_46563);
and U48739 (N_48739,N_46845,N_47404);
xor U48740 (N_48740,N_46709,N_46216);
nor U48741 (N_48741,N_46096,N_45548);
or U48742 (N_48742,N_46174,N_47411);
and U48743 (N_48743,N_45027,N_45557);
and U48744 (N_48744,N_45184,N_47272);
nor U48745 (N_48745,N_45071,N_45485);
and U48746 (N_48746,N_46716,N_45764);
or U48747 (N_48747,N_46012,N_47417);
or U48748 (N_48748,N_46407,N_46459);
or U48749 (N_48749,N_46937,N_47381);
and U48750 (N_48750,N_46524,N_46387);
nor U48751 (N_48751,N_45703,N_46019);
nand U48752 (N_48752,N_47374,N_45643);
and U48753 (N_48753,N_46717,N_46739);
or U48754 (N_48754,N_46040,N_46063);
xor U48755 (N_48755,N_46800,N_46484);
and U48756 (N_48756,N_45127,N_45142);
xor U48757 (N_48757,N_46309,N_47485);
or U48758 (N_48758,N_46795,N_45387);
nand U48759 (N_48759,N_47465,N_47155);
xnor U48760 (N_48760,N_45723,N_46975);
nand U48761 (N_48761,N_45394,N_45647);
or U48762 (N_48762,N_47097,N_46362);
nand U48763 (N_48763,N_45604,N_47239);
and U48764 (N_48764,N_45448,N_45547);
and U48765 (N_48765,N_45935,N_46074);
or U48766 (N_48766,N_46493,N_47371);
and U48767 (N_48767,N_47270,N_45900);
xor U48768 (N_48768,N_46624,N_46065);
nor U48769 (N_48769,N_45804,N_46657);
nor U48770 (N_48770,N_47387,N_46399);
nor U48771 (N_48771,N_45555,N_47424);
xor U48772 (N_48772,N_46684,N_46159);
and U48773 (N_48773,N_47232,N_45709);
xor U48774 (N_48774,N_46614,N_45911);
or U48775 (N_48775,N_47420,N_47157);
nand U48776 (N_48776,N_45629,N_46408);
nand U48777 (N_48777,N_46144,N_45920);
or U48778 (N_48778,N_46010,N_45183);
nor U48779 (N_48779,N_45259,N_47060);
nor U48780 (N_48780,N_46878,N_47034);
and U48781 (N_48781,N_45655,N_46945);
xor U48782 (N_48782,N_45329,N_46036);
nor U48783 (N_48783,N_47199,N_45437);
or U48784 (N_48784,N_47131,N_46619);
xnor U48785 (N_48785,N_47284,N_46115);
and U48786 (N_48786,N_47436,N_45882);
and U48787 (N_48787,N_46687,N_46050);
or U48788 (N_48788,N_47411,N_45828);
or U48789 (N_48789,N_47167,N_46785);
and U48790 (N_48790,N_47038,N_46917);
and U48791 (N_48791,N_45353,N_46290);
nor U48792 (N_48792,N_47078,N_46768);
and U48793 (N_48793,N_45315,N_46648);
nand U48794 (N_48794,N_46977,N_46013);
nor U48795 (N_48795,N_45252,N_47253);
xor U48796 (N_48796,N_47213,N_45342);
and U48797 (N_48797,N_45703,N_46911);
nor U48798 (N_48798,N_45877,N_45077);
or U48799 (N_48799,N_46371,N_45236);
nand U48800 (N_48800,N_45844,N_46668);
xor U48801 (N_48801,N_46792,N_45940);
nand U48802 (N_48802,N_45247,N_47219);
and U48803 (N_48803,N_45322,N_45607);
and U48804 (N_48804,N_46777,N_46134);
and U48805 (N_48805,N_46177,N_45716);
and U48806 (N_48806,N_45744,N_47002);
xor U48807 (N_48807,N_46100,N_46926);
or U48808 (N_48808,N_47247,N_45395);
and U48809 (N_48809,N_46080,N_45298);
or U48810 (N_48810,N_47495,N_45019);
nor U48811 (N_48811,N_46801,N_45753);
and U48812 (N_48812,N_47041,N_47099);
or U48813 (N_48813,N_46204,N_47417);
nor U48814 (N_48814,N_46796,N_45318);
or U48815 (N_48815,N_45780,N_46297);
xor U48816 (N_48816,N_47021,N_47339);
nand U48817 (N_48817,N_45844,N_46362);
nor U48818 (N_48818,N_47422,N_45270);
nand U48819 (N_48819,N_46679,N_45951);
xnor U48820 (N_48820,N_46469,N_46254);
nor U48821 (N_48821,N_46301,N_45111);
nor U48822 (N_48822,N_46277,N_45558);
nand U48823 (N_48823,N_46025,N_45981);
nand U48824 (N_48824,N_45230,N_45641);
or U48825 (N_48825,N_46007,N_45132);
nand U48826 (N_48826,N_46622,N_46967);
xnor U48827 (N_48827,N_45124,N_45774);
nor U48828 (N_48828,N_46980,N_46586);
and U48829 (N_48829,N_46135,N_46026);
nand U48830 (N_48830,N_45448,N_45320);
nand U48831 (N_48831,N_46847,N_45921);
nor U48832 (N_48832,N_45299,N_47174);
and U48833 (N_48833,N_45486,N_46400);
and U48834 (N_48834,N_47425,N_46074);
nor U48835 (N_48835,N_45363,N_46216);
or U48836 (N_48836,N_46042,N_47114);
nor U48837 (N_48837,N_45744,N_46173);
nor U48838 (N_48838,N_45703,N_46215);
nand U48839 (N_48839,N_46223,N_46636);
nor U48840 (N_48840,N_46888,N_45071);
xnor U48841 (N_48841,N_45773,N_46054);
or U48842 (N_48842,N_46937,N_46986);
nand U48843 (N_48843,N_46005,N_46190);
nand U48844 (N_48844,N_46337,N_46513);
xor U48845 (N_48845,N_46660,N_45955);
or U48846 (N_48846,N_47306,N_46266);
or U48847 (N_48847,N_45472,N_45095);
or U48848 (N_48848,N_46349,N_45053);
and U48849 (N_48849,N_45806,N_45077);
and U48850 (N_48850,N_46282,N_46573);
or U48851 (N_48851,N_45722,N_45038);
nand U48852 (N_48852,N_45833,N_47480);
nor U48853 (N_48853,N_46180,N_45631);
xnor U48854 (N_48854,N_46310,N_47371);
or U48855 (N_48855,N_45372,N_46134);
and U48856 (N_48856,N_45249,N_47380);
nand U48857 (N_48857,N_47053,N_46309);
and U48858 (N_48858,N_47088,N_47342);
nand U48859 (N_48859,N_47470,N_45819);
nor U48860 (N_48860,N_47474,N_46162);
nor U48861 (N_48861,N_45467,N_47247);
and U48862 (N_48862,N_46560,N_45576);
or U48863 (N_48863,N_47219,N_45946);
nor U48864 (N_48864,N_46278,N_45617);
nor U48865 (N_48865,N_47321,N_47267);
nand U48866 (N_48866,N_46677,N_46626);
and U48867 (N_48867,N_46112,N_46034);
nand U48868 (N_48868,N_46691,N_46119);
nand U48869 (N_48869,N_46783,N_45335);
nand U48870 (N_48870,N_46936,N_47246);
or U48871 (N_48871,N_45921,N_47367);
or U48872 (N_48872,N_45259,N_47168);
nor U48873 (N_48873,N_46801,N_45526);
xnor U48874 (N_48874,N_47063,N_46718);
or U48875 (N_48875,N_46073,N_46896);
nand U48876 (N_48876,N_45743,N_47276);
nor U48877 (N_48877,N_45877,N_45930);
nor U48878 (N_48878,N_46853,N_45834);
nand U48879 (N_48879,N_46434,N_47455);
xnor U48880 (N_48880,N_45844,N_47088);
xor U48881 (N_48881,N_45241,N_45139);
or U48882 (N_48882,N_45438,N_46127);
nor U48883 (N_48883,N_46972,N_46954);
xor U48884 (N_48884,N_46866,N_45283);
or U48885 (N_48885,N_46416,N_45545);
nand U48886 (N_48886,N_46817,N_45833);
and U48887 (N_48887,N_45579,N_45024);
or U48888 (N_48888,N_47138,N_45432);
and U48889 (N_48889,N_45190,N_46172);
or U48890 (N_48890,N_47108,N_46484);
xnor U48891 (N_48891,N_45905,N_47269);
xor U48892 (N_48892,N_47247,N_46996);
nor U48893 (N_48893,N_46245,N_46244);
or U48894 (N_48894,N_46674,N_45213);
nand U48895 (N_48895,N_45195,N_46016);
xor U48896 (N_48896,N_46876,N_45776);
or U48897 (N_48897,N_46347,N_45596);
and U48898 (N_48898,N_46119,N_45524);
xnor U48899 (N_48899,N_46585,N_47409);
xor U48900 (N_48900,N_47208,N_46361);
or U48901 (N_48901,N_45129,N_47039);
or U48902 (N_48902,N_45974,N_45462);
or U48903 (N_48903,N_45875,N_46574);
or U48904 (N_48904,N_45399,N_45414);
nor U48905 (N_48905,N_47366,N_47300);
and U48906 (N_48906,N_46958,N_46588);
nor U48907 (N_48907,N_45517,N_45941);
or U48908 (N_48908,N_45357,N_45401);
or U48909 (N_48909,N_47011,N_45677);
or U48910 (N_48910,N_47318,N_45351);
or U48911 (N_48911,N_45312,N_46019);
or U48912 (N_48912,N_45897,N_47147);
and U48913 (N_48913,N_46005,N_46645);
and U48914 (N_48914,N_46567,N_46838);
and U48915 (N_48915,N_46282,N_46302);
nor U48916 (N_48916,N_47236,N_45640);
or U48917 (N_48917,N_45777,N_47188);
nor U48918 (N_48918,N_45042,N_46785);
xor U48919 (N_48919,N_46164,N_45276);
nor U48920 (N_48920,N_46751,N_46362);
nor U48921 (N_48921,N_46692,N_46152);
nand U48922 (N_48922,N_45882,N_45031);
or U48923 (N_48923,N_45989,N_46950);
xnor U48924 (N_48924,N_47244,N_45767);
or U48925 (N_48925,N_46175,N_46820);
nor U48926 (N_48926,N_46411,N_45506);
nand U48927 (N_48927,N_47429,N_46921);
and U48928 (N_48928,N_45999,N_45454);
nand U48929 (N_48929,N_47071,N_46510);
nor U48930 (N_48930,N_46694,N_45885);
nor U48931 (N_48931,N_45071,N_45039);
nand U48932 (N_48932,N_45620,N_45080);
and U48933 (N_48933,N_47285,N_45236);
nor U48934 (N_48934,N_45095,N_45627);
and U48935 (N_48935,N_45908,N_47445);
xor U48936 (N_48936,N_47271,N_45411);
nor U48937 (N_48937,N_47011,N_46126);
or U48938 (N_48938,N_46056,N_45209);
nand U48939 (N_48939,N_45203,N_46099);
nand U48940 (N_48940,N_45344,N_47245);
nor U48941 (N_48941,N_47041,N_47279);
and U48942 (N_48942,N_46687,N_46900);
nor U48943 (N_48943,N_46381,N_46251);
xor U48944 (N_48944,N_45054,N_46770);
nor U48945 (N_48945,N_46406,N_45101);
and U48946 (N_48946,N_46914,N_46151);
xnor U48947 (N_48947,N_46472,N_46757);
xnor U48948 (N_48948,N_46347,N_47114);
nor U48949 (N_48949,N_45577,N_46453);
and U48950 (N_48950,N_46534,N_47411);
nor U48951 (N_48951,N_46967,N_46377);
or U48952 (N_48952,N_45201,N_46909);
nand U48953 (N_48953,N_46071,N_45515);
or U48954 (N_48954,N_45341,N_45674);
nand U48955 (N_48955,N_47282,N_45807);
nor U48956 (N_48956,N_46587,N_46824);
xnor U48957 (N_48957,N_45617,N_45131);
or U48958 (N_48958,N_46614,N_45383);
xor U48959 (N_48959,N_47382,N_47274);
nand U48960 (N_48960,N_47412,N_45630);
or U48961 (N_48961,N_47456,N_46027);
nor U48962 (N_48962,N_45756,N_45624);
or U48963 (N_48963,N_45428,N_45509);
and U48964 (N_48964,N_47285,N_45933);
xor U48965 (N_48965,N_45978,N_45960);
nand U48966 (N_48966,N_45497,N_46465);
or U48967 (N_48967,N_46049,N_46919);
nand U48968 (N_48968,N_46386,N_47058);
nand U48969 (N_48969,N_45054,N_46360);
nand U48970 (N_48970,N_46986,N_46232);
nand U48971 (N_48971,N_46387,N_47079);
xor U48972 (N_48972,N_47236,N_45760);
nand U48973 (N_48973,N_45089,N_46518);
xor U48974 (N_48974,N_46541,N_47083);
nand U48975 (N_48975,N_45418,N_46482);
and U48976 (N_48976,N_45264,N_46985);
and U48977 (N_48977,N_46962,N_45393);
xor U48978 (N_48978,N_47485,N_45955);
xnor U48979 (N_48979,N_46215,N_45562);
nand U48980 (N_48980,N_45215,N_46548);
xnor U48981 (N_48981,N_45332,N_45797);
nor U48982 (N_48982,N_45862,N_47265);
nor U48983 (N_48983,N_46875,N_47082);
nand U48984 (N_48984,N_46007,N_47123);
nand U48985 (N_48985,N_46932,N_47233);
nor U48986 (N_48986,N_46137,N_45543);
xor U48987 (N_48987,N_45342,N_46804);
nor U48988 (N_48988,N_46564,N_47378);
or U48989 (N_48989,N_45826,N_46748);
xnor U48990 (N_48990,N_46109,N_46897);
and U48991 (N_48991,N_45697,N_45389);
or U48992 (N_48992,N_46726,N_45160);
nand U48993 (N_48993,N_45468,N_45855);
and U48994 (N_48994,N_46589,N_45710);
xnor U48995 (N_48995,N_45144,N_46734);
xor U48996 (N_48996,N_45884,N_46137);
nand U48997 (N_48997,N_45382,N_46799);
and U48998 (N_48998,N_45496,N_46575);
xnor U48999 (N_48999,N_45390,N_46987);
or U49000 (N_49000,N_46695,N_45915);
xnor U49001 (N_49001,N_46030,N_46350);
and U49002 (N_49002,N_45133,N_47458);
nor U49003 (N_49003,N_46713,N_46948);
xor U49004 (N_49004,N_46993,N_45107);
nand U49005 (N_49005,N_46671,N_47256);
nand U49006 (N_49006,N_46296,N_46962);
nor U49007 (N_49007,N_46473,N_45295);
or U49008 (N_49008,N_47346,N_45738);
xnor U49009 (N_49009,N_46325,N_45878);
and U49010 (N_49010,N_46959,N_47169);
nor U49011 (N_49011,N_45844,N_45881);
xor U49012 (N_49012,N_46793,N_45931);
xnor U49013 (N_49013,N_46204,N_46536);
and U49014 (N_49014,N_46481,N_45020);
xnor U49015 (N_49015,N_46662,N_46438);
nor U49016 (N_49016,N_45742,N_46926);
and U49017 (N_49017,N_46698,N_45081);
xor U49018 (N_49018,N_46033,N_45966);
or U49019 (N_49019,N_46659,N_45599);
and U49020 (N_49020,N_46120,N_45952);
or U49021 (N_49021,N_47413,N_46865);
and U49022 (N_49022,N_47289,N_46766);
or U49023 (N_49023,N_45127,N_46061);
xor U49024 (N_49024,N_45597,N_46279);
nor U49025 (N_49025,N_45385,N_47376);
and U49026 (N_49026,N_47310,N_46124);
and U49027 (N_49027,N_45850,N_45874);
nand U49028 (N_49028,N_46771,N_46090);
nand U49029 (N_49029,N_45808,N_47138);
or U49030 (N_49030,N_45029,N_45126);
or U49031 (N_49031,N_45817,N_47058);
nor U49032 (N_49032,N_45221,N_46757);
nand U49033 (N_49033,N_45547,N_45725);
and U49034 (N_49034,N_45065,N_45566);
xor U49035 (N_49035,N_46414,N_46805);
or U49036 (N_49036,N_46780,N_46777);
nor U49037 (N_49037,N_47343,N_46731);
nand U49038 (N_49038,N_45265,N_46527);
xor U49039 (N_49039,N_46278,N_45105);
nand U49040 (N_49040,N_46974,N_47097);
and U49041 (N_49041,N_45301,N_46586);
xor U49042 (N_49042,N_47085,N_46502);
nor U49043 (N_49043,N_45544,N_47424);
or U49044 (N_49044,N_46684,N_45331);
nor U49045 (N_49045,N_45778,N_46198);
nor U49046 (N_49046,N_46769,N_47391);
nor U49047 (N_49047,N_45015,N_45963);
or U49048 (N_49048,N_47278,N_45626);
or U49049 (N_49049,N_47339,N_47412);
nor U49050 (N_49050,N_47482,N_45543);
or U49051 (N_49051,N_46135,N_47078);
nor U49052 (N_49052,N_47026,N_45929);
and U49053 (N_49053,N_46446,N_46007);
nor U49054 (N_49054,N_46911,N_45244);
xor U49055 (N_49055,N_46691,N_46474);
or U49056 (N_49056,N_46087,N_47278);
xnor U49057 (N_49057,N_47479,N_45235);
xnor U49058 (N_49058,N_45007,N_46492);
and U49059 (N_49059,N_46080,N_47167);
or U49060 (N_49060,N_45735,N_45651);
nor U49061 (N_49061,N_45263,N_45798);
xnor U49062 (N_49062,N_45894,N_45135);
nand U49063 (N_49063,N_45285,N_45594);
or U49064 (N_49064,N_47431,N_45346);
and U49065 (N_49065,N_45954,N_46201);
and U49066 (N_49066,N_45411,N_45174);
nand U49067 (N_49067,N_46427,N_46393);
and U49068 (N_49068,N_45408,N_46714);
and U49069 (N_49069,N_47057,N_45537);
nand U49070 (N_49070,N_46604,N_47013);
or U49071 (N_49071,N_45811,N_45189);
nor U49072 (N_49072,N_45937,N_46943);
or U49073 (N_49073,N_46801,N_45513);
or U49074 (N_49074,N_45173,N_45709);
nand U49075 (N_49075,N_46364,N_46155);
xnor U49076 (N_49076,N_45924,N_45687);
and U49077 (N_49077,N_45169,N_47345);
and U49078 (N_49078,N_47384,N_47272);
nor U49079 (N_49079,N_45310,N_47283);
nor U49080 (N_49080,N_47381,N_46830);
and U49081 (N_49081,N_46070,N_45691);
xnor U49082 (N_49082,N_47305,N_45027);
and U49083 (N_49083,N_45563,N_45828);
nand U49084 (N_49084,N_47142,N_45785);
xor U49085 (N_49085,N_46517,N_45527);
xor U49086 (N_49086,N_46382,N_46574);
xnor U49087 (N_49087,N_47412,N_46139);
xnor U49088 (N_49088,N_45081,N_45085);
or U49089 (N_49089,N_45258,N_45368);
xnor U49090 (N_49090,N_45774,N_47213);
nor U49091 (N_49091,N_47311,N_47388);
xor U49092 (N_49092,N_45500,N_46109);
nand U49093 (N_49093,N_46055,N_46090);
nor U49094 (N_49094,N_45623,N_46272);
and U49095 (N_49095,N_46775,N_45838);
nand U49096 (N_49096,N_46456,N_47214);
xor U49097 (N_49097,N_45213,N_45145);
nand U49098 (N_49098,N_47089,N_45211);
and U49099 (N_49099,N_46423,N_46170);
nand U49100 (N_49100,N_47302,N_45734);
nor U49101 (N_49101,N_46454,N_46663);
xnor U49102 (N_49102,N_46566,N_46456);
nor U49103 (N_49103,N_46310,N_45297);
nor U49104 (N_49104,N_45399,N_46488);
nor U49105 (N_49105,N_45766,N_45878);
or U49106 (N_49106,N_46115,N_45463);
and U49107 (N_49107,N_45423,N_47031);
and U49108 (N_49108,N_45242,N_46974);
or U49109 (N_49109,N_45570,N_46405);
nand U49110 (N_49110,N_45020,N_47470);
and U49111 (N_49111,N_46470,N_46338);
xnor U49112 (N_49112,N_45186,N_46006);
or U49113 (N_49113,N_45252,N_47246);
nand U49114 (N_49114,N_45165,N_46456);
nand U49115 (N_49115,N_45119,N_45223);
and U49116 (N_49116,N_46232,N_47156);
xnor U49117 (N_49117,N_47008,N_47084);
and U49118 (N_49118,N_47033,N_46328);
nor U49119 (N_49119,N_45037,N_46852);
or U49120 (N_49120,N_45604,N_45589);
nand U49121 (N_49121,N_47120,N_45340);
xnor U49122 (N_49122,N_47229,N_45881);
xnor U49123 (N_49123,N_45714,N_45739);
or U49124 (N_49124,N_45892,N_45740);
and U49125 (N_49125,N_45849,N_46274);
xnor U49126 (N_49126,N_45566,N_46266);
or U49127 (N_49127,N_47068,N_45319);
or U49128 (N_49128,N_45202,N_46718);
xnor U49129 (N_49129,N_45229,N_47458);
or U49130 (N_49130,N_47487,N_45408);
or U49131 (N_49131,N_46886,N_46684);
or U49132 (N_49132,N_46109,N_46890);
or U49133 (N_49133,N_45588,N_47297);
and U49134 (N_49134,N_45483,N_47461);
xnor U49135 (N_49135,N_46688,N_46570);
nor U49136 (N_49136,N_47376,N_45204);
xnor U49137 (N_49137,N_47331,N_45873);
and U49138 (N_49138,N_47373,N_47270);
and U49139 (N_49139,N_46511,N_46953);
nor U49140 (N_49140,N_45491,N_46214);
and U49141 (N_49141,N_45700,N_46743);
or U49142 (N_49142,N_47249,N_45599);
and U49143 (N_49143,N_45887,N_45431);
nor U49144 (N_49144,N_46014,N_45274);
nor U49145 (N_49145,N_45050,N_46766);
xor U49146 (N_49146,N_46938,N_45819);
or U49147 (N_49147,N_47077,N_46821);
nor U49148 (N_49148,N_46661,N_45711);
or U49149 (N_49149,N_45472,N_47044);
nor U49150 (N_49150,N_47306,N_45595);
xnor U49151 (N_49151,N_46147,N_45488);
or U49152 (N_49152,N_47088,N_47170);
or U49153 (N_49153,N_47163,N_47235);
and U49154 (N_49154,N_46492,N_46892);
and U49155 (N_49155,N_46288,N_46963);
nand U49156 (N_49156,N_45458,N_47421);
xnor U49157 (N_49157,N_46617,N_46214);
or U49158 (N_49158,N_46085,N_47061);
nor U49159 (N_49159,N_45284,N_45358);
and U49160 (N_49160,N_47333,N_46143);
or U49161 (N_49161,N_45607,N_45663);
nand U49162 (N_49162,N_46703,N_46016);
xnor U49163 (N_49163,N_45057,N_47014);
nand U49164 (N_49164,N_45808,N_47097);
nor U49165 (N_49165,N_46927,N_47331);
xnor U49166 (N_49166,N_45890,N_46259);
nand U49167 (N_49167,N_45506,N_47058);
nor U49168 (N_49168,N_45933,N_46965);
and U49169 (N_49169,N_46506,N_47104);
and U49170 (N_49170,N_45823,N_45452);
nand U49171 (N_49171,N_45002,N_45675);
nor U49172 (N_49172,N_46917,N_46483);
and U49173 (N_49173,N_45327,N_46170);
and U49174 (N_49174,N_45893,N_46207);
xnor U49175 (N_49175,N_46121,N_45221);
xnor U49176 (N_49176,N_46341,N_45133);
nand U49177 (N_49177,N_46299,N_46494);
xor U49178 (N_49178,N_45731,N_46630);
nor U49179 (N_49179,N_45240,N_45468);
nand U49180 (N_49180,N_46863,N_45163);
or U49181 (N_49181,N_46916,N_46334);
or U49182 (N_49182,N_46332,N_45514);
xnor U49183 (N_49183,N_46189,N_45427);
nor U49184 (N_49184,N_47244,N_47086);
nand U49185 (N_49185,N_46720,N_46488);
xor U49186 (N_49186,N_46975,N_45653);
or U49187 (N_49187,N_45227,N_47045);
or U49188 (N_49188,N_45628,N_47326);
xor U49189 (N_49189,N_46292,N_45475);
xor U49190 (N_49190,N_47102,N_46425);
nor U49191 (N_49191,N_45858,N_46885);
or U49192 (N_49192,N_45749,N_46922);
or U49193 (N_49193,N_45256,N_45395);
nor U49194 (N_49194,N_46990,N_45682);
or U49195 (N_49195,N_46151,N_46228);
nor U49196 (N_49196,N_46412,N_46148);
nand U49197 (N_49197,N_47384,N_45473);
nand U49198 (N_49198,N_47399,N_46473);
xor U49199 (N_49199,N_45785,N_46626);
or U49200 (N_49200,N_45631,N_47030);
nand U49201 (N_49201,N_45141,N_46261);
or U49202 (N_49202,N_45647,N_46175);
nand U49203 (N_49203,N_45338,N_45993);
xnor U49204 (N_49204,N_46257,N_45444);
and U49205 (N_49205,N_47464,N_46841);
nor U49206 (N_49206,N_46481,N_45649);
xnor U49207 (N_49207,N_45790,N_46902);
nor U49208 (N_49208,N_46011,N_45639);
or U49209 (N_49209,N_46941,N_46081);
and U49210 (N_49210,N_45128,N_47441);
and U49211 (N_49211,N_46078,N_45227);
xnor U49212 (N_49212,N_46179,N_45231);
nand U49213 (N_49213,N_45045,N_47255);
or U49214 (N_49214,N_46014,N_46810);
nor U49215 (N_49215,N_46233,N_46455);
and U49216 (N_49216,N_47379,N_45658);
xnor U49217 (N_49217,N_45883,N_47270);
nor U49218 (N_49218,N_46283,N_46500);
and U49219 (N_49219,N_46192,N_46866);
and U49220 (N_49220,N_47459,N_45148);
xnor U49221 (N_49221,N_46820,N_46268);
or U49222 (N_49222,N_47075,N_45050);
nand U49223 (N_49223,N_45390,N_47235);
xnor U49224 (N_49224,N_45452,N_45029);
and U49225 (N_49225,N_46099,N_45343);
nand U49226 (N_49226,N_46952,N_45463);
or U49227 (N_49227,N_47333,N_46747);
nand U49228 (N_49228,N_45718,N_47110);
xor U49229 (N_49229,N_47418,N_45393);
xor U49230 (N_49230,N_46931,N_45571);
or U49231 (N_49231,N_45772,N_46669);
or U49232 (N_49232,N_46206,N_45238);
nand U49233 (N_49233,N_46275,N_46403);
nor U49234 (N_49234,N_47182,N_46225);
and U49235 (N_49235,N_45713,N_45080);
nor U49236 (N_49236,N_46626,N_45019);
nand U49237 (N_49237,N_47363,N_47099);
or U49238 (N_49238,N_47441,N_46092);
nand U49239 (N_49239,N_45025,N_47474);
nand U49240 (N_49240,N_46623,N_47092);
nor U49241 (N_49241,N_46092,N_46544);
or U49242 (N_49242,N_46508,N_45444);
xnor U49243 (N_49243,N_45368,N_46938);
xor U49244 (N_49244,N_45995,N_45303);
nor U49245 (N_49245,N_46568,N_45832);
xor U49246 (N_49246,N_46428,N_45652);
xor U49247 (N_49247,N_45766,N_45697);
or U49248 (N_49248,N_47004,N_45449);
nand U49249 (N_49249,N_45838,N_45973);
or U49250 (N_49250,N_45836,N_45342);
xor U49251 (N_49251,N_46675,N_47016);
xor U49252 (N_49252,N_45824,N_45390);
nand U49253 (N_49253,N_46379,N_46216);
nand U49254 (N_49254,N_47450,N_46058);
and U49255 (N_49255,N_45564,N_46746);
nor U49256 (N_49256,N_45991,N_46146);
and U49257 (N_49257,N_46370,N_47488);
and U49258 (N_49258,N_45558,N_45832);
or U49259 (N_49259,N_45573,N_47164);
xor U49260 (N_49260,N_45927,N_46923);
nand U49261 (N_49261,N_46646,N_46930);
and U49262 (N_49262,N_46978,N_46113);
or U49263 (N_49263,N_46983,N_45312);
nor U49264 (N_49264,N_45842,N_46873);
xnor U49265 (N_49265,N_46545,N_45347);
and U49266 (N_49266,N_45586,N_47238);
xor U49267 (N_49267,N_46339,N_47199);
xor U49268 (N_49268,N_45506,N_45641);
and U49269 (N_49269,N_45844,N_45151);
and U49270 (N_49270,N_45003,N_46784);
xor U49271 (N_49271,N_46039,N_45760);
and U49272 (N_49272,N_46426,N_46574);
nor U49273 (N_49273,N_47273,N_47476);
or U49274 (N_49274,N_46854,N_45624);
or U49275 (N_49275,N_45922,N_47079);
or U49276 (N_49276,N_45013,N_46715);
nand U49277 (N_49277,N_45080,N_45269);
nand U49278 (N_49278,N_47053,N_45745);
xnor U49279 (N_49279,N_47339,N_46347);
nand U49280 (N_49280,N_46927,N_46104);
and U49281 (N_49281,N_45187,N_47467);
nor U49282 (N_49282,N_47230,N_46981);
or U49283 (N_49283,N_46617,N_45954);
or U49284 (N_49284,N_46807,N_45969);
nand U49285 (N_49285,N_45538,N_47012);
nand U49286 (N_49286,N_46617,N_45141);
nand U49287 (N_49287,N_46993,N_46583);
or U49288 (N_49288,N_47118,N_45592);
nor U49289 (N_49289,N_46765,N_45898);
nor U49290 (N_49290,N_45935,N_47447);
xor U49291 (N_49291,N_45182,N_45350);
and U49292 (N_49292,N_46071,N_45925);
or U49293 (N_49293,N_46908,N_45673);
nand U49294 (N_49294,N_46347,N_47050);
nor U49295 (N_49295,N_46197,N_45568);
or U49296 (N_49296,N_47386,N_46346);
nand U49297 (N_49297,N_45005,N_47490);
nand U49298 (N_49298,N_45372,N_45364);
xor U49299 (N_49299,N_45906,N_46595);
xnor U49300 (N_49300,N_45283,N_46915);
and U49301 (N_49301,N_45624,N_46782);
xnor U49302 (N_49302,N_45100,N_45586);
nor U49303 (N_49303,N_47154,N_47139);
nand U49304 (N_49304,N_45535,N_46366);
xor U49305 (N_49305,N_45742,N_45085);
xnor U49306 (N_49306,N_45183,N_45053);
or U49307 (N_49307,N_45479,N_45159);
and U49308 (N_49308,N_45980,N_45197);
nand U49309 (N_49309,N_47161,N_45100);
and U49310 (N_49310,N_45659,N_45773);
nor U49311 (N_49311,N_46016,N_47366);
nand U49312 (N_49312,N_46748,N_45143);
xnor U49313 (N_49313,N_46137,N_47221);
xnor U49314 (N_49314,N_45406,N_45736);
and U49315 (N_49315,N_45671,N_46585);
and U49316 (N_49316,N_45064,N_47356);
and U49317 (N_49317,N_45182,N_45435);
or U49318 (N_49318,N_46291,N_47369);
and U49319 (N_49319,N_45131,N_45130);
xnor U49320 (N_49320,N_45748,N_46594);
nor U49321 (N_49321,N_45189,N_47314);
nor U49322 (N_49322,N_47409,N_45665);
or U49323 (N_49323,N_45169,N_46527);
and U49324 (N_49324,N_46073,N_46820);
and U49325 (N_49325,N_46908,N_46789);
xor U49326 (N_49326,N_46737,N_46980);
nand U49327 (N_49327,N_45731,N_46376);
or U49328 (N_49328,N_45035,N_46598);
and U49329 (N_49329,N_46633,N_46020);
nor U49330 (N_49330,N_45674,N_46226);
nor U49331 (N_49331,N_46352,N_46528);
nor U49332 (N_49332,N_45137,N_46457);
xor U49333 (N_49333,N_45923,N_45407);
and U49334 (N_49334,N_46822,N_46521);
nor U49335 (N_49335,N_45314,N_47129);
nand U49336 (N_49336,N_47233,N_47173);
nor U49337 (N_49337,N_47414,N_45256);
nor U49338 (N_49338,N_47405,N_45797);
and U49339 (N_49339,N_46733,N_46016);
and U49340 (N_49340,N_45354,N_47226);
or U49341 (N_49341,N_45024,N_46904);
nor U49342 (N_49342,N_46792,N_47154);
nand U49343 (N_49343,N_46472,N_46759);
nor U49344 (N_49344,N_45995,N_46071);
nor U49345 (N_49345,N_46682,N_47365);
nor U49346 (N_49346,N_45974,N_45137);
and U49347 (N_49347,N_46699,N_47094);
nor U49348 (N_49348,N_46538,N_46025);
or U49349 (N_49349,N_47246,N_46791);
or U49350 (N_49350,N_47163,N_45421);
or U49351 (N_49351,N_45279,N_47382);
and U49352 (N_49352,N_46039,N_47362);
xnor U49353 (N_49353,N_45623,N_45857);
nor U49354 (N_49354,N_46050,N_45446);
xor U49355 (N_49355,N_45634,N_45362);
nand U49356 (N_49356,N_46642,N_45630);
xor U49357 (N_49357,N_45927,N_47400);
or U49358 (N_49358,N_46591,N_45488);
or U49359 (N_49359,N_46675,N_45067);
xor U49360 (N_49360,N_45903,N_46486);
or U49361 (N_49361,N_47318,N_46667);
xnor U49362 (N_49362,N_46334,N_45359);
and U49363 (N_49363,N_46190,N_45143);
nand U49364 (N_49364,N_47203,N_45797);
and U49365 (N_49365,N_47239,N_47152);
and U49366 (N_49366,N_46661,N_46450);
nand U49367 (N_49367,N_45225,N_46838);
xnor U49368 (N_49368,N_45345,N_46251);
or U49369 (N_49369,N_46116,N_47428);
nor U49370 (N_49370,N_45589,N_45514);
or U49371 (N_49371,N_45800,N_46981);
and U49372 (N_49372,N_45299,N_46096);
xor U49373 (N_49373,N_46963,N_47035);
and U49374 (N_49374,N_47187,N_45614);
nand U49375 (N_49375,N_45322,N_47073);
nand U49376 (N_49376,N_45271,N_45249);
or U49377 (N_49377,N_46573,N_46286);
and U49378 (N_49378,N_46329,N_46146);
nand U49379 (N_49379,N_45812,N_45948);
nand U49380 (N_49380,N_46206,N_45154);
or U49381 (N_49381,N_45904,N_45428);
nor U49382 (N_49382,N_45499,N_47149);
or U49383 (N_49383,N_46403,N_45733);
nor U49384 (N_49384,N_45918,N_45898);
xnor U49385 (N_49385,N_45795,N_45202);
xor U49386 (N_49386,N_45097,N_45988);
and U49387 (N_49387,N_46832,N_45509);
nor U49388 (N_49388,N_47209,N_46141);
nor U49389 (N_49389,N_45378,N_45427);
xor U49390 (N_49390,N_47131,N_46674);
nor U49391 (N_49391,N_45960,N_45500);
xor U49392 (N_49392,N_47068,N_45656);
or U49393 (N_49393,N_47310,N_47237);
or U49394 (N_49394,N_46064,N_47443);
nor U49395 (N_49395,N_45820,N_45868);
nor U49396 (N_49396,N_46949,N_46605);
and U49397 (N_49397,N_47051,N_45796);
nor U49398 (N_49398,N_47123,N_46774);
xor U49399 (N_49399,N_46044,N_47436);
xnor U49400 (N_49400,N_45386,N_46694);
and U49401 (N_49401,N_46484,N_46963);
xor U49402 (N_49402,N_46588,N_47206);
or U49403 (N_49403,N_46406,N_46671);
nor U49404 (N_49404,N_47084,N_46653);
nand U49405 (N_49405,N_47080,N_46558);
and U49406 (N_49406,N_46981,N_46573);
or U49407 (N_49407,N_45606,N_45379);
nand U49408 (N_49408,N_46346,N_47111);
and U49409 (N_49409,N_46238,N_47028);
nand U49410 (N_49410,N_45868,N_46200);
and U49411 (N_49411,N_45047,N_45597);
or U49412 (N_49412,N_47323,N_45342);
nor U49413 (N_49413,N_45096,N_46514);
and U49414 (N_49414,N_47301,N_46715);
nor U49415 (N_49415,N_45811,N_45699);
or U49416 (N_49416,N_46527,N_45840);
nand U49417 (N_49417,N_47092,N_45534);
or U49418 (N_49418,N_46300,N_46839);
nor U49419 (N_49419,N_46672,N_45668);
and U49420 (N_49420,N_47136,N_47369);
nor U49421 (N_49421,N_45437,N_46164);
nor U49422 (N_49422,N_45041,N_47324);
xor U49423 (N_49423,N_46611,N_46210);
nand U49424 (N_49424,N_45192,N_46875);
or U49425 (N_49425,N_46880,N_45488);
nor U49426 (N_49426,N_45850,N_45713);
xor U49427 (N_49427,N_45640,N_46505);
nand U49428 (N_49428,N_45704,N_47072);
xor U49429 (N_49429,N_46620,N_45795);
nand U49430 (N_49430,N_46531,N_45696);
xnor U49431 (N_49431,N_45744,N_46225);
xor U49432 (N_49432,N_47371,N_46053);
xor U49433 (N_49433,N_45246,N_46734);
and U49434 (N_49434,N_45538,N_47250);
or U49435 (N_49435,N_45956,N_46843);
or U49436 (N_49436,N_46412,N_45671);
xor U49437 (N_49437,N_45544,N_45878);
and U49438 (N_49438,N_45828,N_46773);
xor U49439 (N_49439,N_46250,N_45281);
or U49440 (N_49440,N_45454,N_45810);
nor U49441 (N_49441,N_47340,N_46591);
and U49442 (N_49442,N_46700,N_46330);
xnor U49443 (N_49443,N_45750,N_46148);
xnor U49444 (N_49444,N_46752,N_46572);
nand U49445 (N_49445,N_47146,N_46547);
and U49446 (N_49446,N_46598,N_46553);
nand U49447 (N_49447,N_45474,N_46788);
or U49448 (N_49448,N_45634,N_45902);
nand U49449 (N_49449,N_46738,N_47212);
nor U49450 (N_49450,N_45025,N_45565);
nor U49451 (N_49451,N_46877,N_46108);
nor U49452 (N_49452,N_46065,N_46611);
or U49453 (N_49453,N_45211,N_45017);
nand U49454 (N_49454,N_45710,N_47425);
and U49455 (N_49455,N_45305,N_47006);
and U49456 (N_49456,N_47347,N_45035);
and U49457 (N_49457,N_45864,N_47248);
xnor U49458 (N_49458,N_45189,N_45930);
or U49459 (N_49459,N_47469,N_45946);
nor U49460 (N_49460,N_46799,N_45351);
nand U49461 (N_49461,N_46987,N_46948);
or U49462 (N_49462,N_46390,N_45404);
or U49463 (N_49463,N_46119,N_47383);
or U49464 (N_49464,N_46902,N_46802);
or U49465 (N_49465,N_45690,N_46260);
nor U49466 (N_49466,N_45623,N_45875);
nor U49467 (N_49467,N_47324,N_45749);
nor U49468 (N_49468,N_46527,N_47487);
nor U49469 (N_49469,N_45421,N_45424);
xor U49470 (N_49470,N_46551,N_46099);
xnor U49471 (N_49471,N_46595,N_46533);
or U49472 (N_49472,N_46218,N_46387);
nand U49473 (N_49473,N_45918,N_46580);
nand U49474 (N_49474,N_47395,N_45244);
or U49475 (N_49475,N_45480,N_46708);
nor U49476 (N_49476,N_46897,N_45680);
and U49477 (N_49477,N_46165,N_47244);
and U49478 (N_49478,N_46800,N_46521);
nand U49479 (N_49479,N_45766,N_46351);
or U49480 (N_49480,N_46300,N_46961);
nand U49481 (N_49481,N_45441,N_46264);
nand U49482 (N_49482,N_46027,N_46980);
nand U49483 (N_49483,N_46100,N_45922);
or U49484 (N_49484,N_45892,N_45249);
nand U49485 (N_49485,N_45669,N_46154);
xnor U49486 (N_49486,N_46144,N_46120);
nor U49487 (N_49487,N_45924,N_46771);
xnor U49488 (N_49488,N_47355,N_47175);
or U49489 (N_49489,N_45068,N_46890);
xnor U49490 (N_49490,N_45120,N_46530);
nand U49491 (N_49491,N_45235,N_46229);
or U49492 (N_49492,N_45522,N_46416);
nor U49493 (N_49493,N_45370,N_47452);
and U49494 (N_49494,N_45197,N_47170);
xor U49495 (N_49495,N_45875,N_46928);
xor U49496 (N_49496,N_45535,N_45169);
and U49497 (N_49497,N_46613,N_47452);
and U49498 (N_49498,N_45884,N_46665);
and U49499 (N_49499,N_47475,N_46184);
or U49500 (N_49500,N_45353,N_47086);
xnor U49501 (N_49501,N_46142,N_46964);
nor U49502 (N_49502,N_47311,N_45429);
xor U49503 (N_49503,N_45527,N_46888);
xor U49504 (N_49504,N_45291,N_46707);
or U49505 (N_49505,N_45291,N_46547);
nor U49506 (N_49506,N_46426,N_46608);
xor U49507 (N_49507,N_46962,N_46070);
xnor U49508 (N_49508,N_47014,N_45207);
and U49509 (N_49509,N_45876,N_47164);
and U49510 (N_49510,N_47429,N_45306);
and U49511 (N_49511,N_45857,N_45279);
nand U49512 (N_49512,N_47138,N_45839);
xnor U49513 (N_49513,N_47364,N_45651);
nor U49514 (N_49514,N_47431,N_46007);
xor U49515 (N_49515,N_46576,N_47419);
nor U49516 (N_49516,N_46910,N_46515);
nand U49517 (N_49517,N_45351,N_47077);
or U49518 (N_49518,N_46556,N_46752);
nand U49519 (N_49519,N_45276,N_46010);
xnor U49520 (N_49520,N_46296,N_45583);
nand U49521 (N_49521,N_45156,N_45791);
nand U49522 (N_49522,N_45890,N_46137);
xor U49523 (N_49523,N_46141,N_46294);
or U49524 (N_49524,N_47272,N_46236);
nand U49525 (N_49525,N_47407,N_47190);
nand U49526 (N_49526,N_45734,N_46789);
xnor U49527 (N_49527,N_45232,N_47422);
or U49528 (N_49528,N_45416,N_46265);
nor U49529 (N_49529,N_46986,N_46178);
xor U49530 (N_49530,N_46247,N_46799);
xnor U49531 (N_49531,N_47305,N_46255);
and U49532 (N_49532,N_46115,N_46891);
or U49533 (N_49533,N_46127,N_46001);
nand U49534 (N_49534,N_46030,N_45270);
or U49535 (N_49535,N_46558,N_46962);
nor U49536 (N_49536,N_47023,N_45188);
nor U49537 (N_49537,N_47068,N_47202);
nand U49538 (N_49538,N_46027,N_46637);
and U49539 (N_49539,N_47030,N_47012);
xnor U49540 (N_49540,N_46659,N_47435);
nor U49541 (N_49541,N_46054,N_45289);
or U49542 (N_49542,N_46084,N_46517);
nand U49543 (N_49543,N_46212,N_45439);
nand U49544 (N_49544,N_45509,N_45318);
nand U49545 (N_49545,N_45321,N_45300);
nor U49546 (N_49546,N_45884,N_45606);
nor U49547 (N_49547,N_45498,N_45969);
nor U49548 (N_49548,N_47160,N_46033);
xor U49549 (N_49549,N_47376,N_45835);
and U49550 (N_49550,N_45476,N_45652);
nor U49551 (N_49551,N_45316,N_46619);
nand U49552 (N_49552,N_45574,N_45209);
and U49553 (N_49553,N_47495,N_45013);
and U49554 (N_49554,N_46157,N_47399);
or U49555 (N_49555,N_45146,N_46533);
xnor U49556 (N_49556,N_46104,N_47295);
xor U49557 (N_49557,N_45590,N_46431);
and U49558 (N_49558,N_47259,N_46004);
and U49559 (N_49559,N_46653,N_47314);
nor U49560 (N_49560,N_46989,N_47389);
xnor U49561 (N_49561,N_46699,N_46703);
xnor U49562 (N_49562,N_45307,N_45355);
nand U49563 (N_49563,N_46072,N_45198);
and U49564 (N_49564,N_47221,N_45945);
nand U49565 (N_49565,N_46114,N_45018);
nor U49566 (N_49566,N_45374,N_45263);
nor U49567 (N_49567,N_46170,N_45462);
or U49568 (N_49568,N_45590,N_46684);
or U49569 (N_49569,N_45930,N_45007);
and U49570 (N_49570,N_45354,N_46065);
and U49571 (N_49571,N_45320,N_47485);
and U49572 (N_49572,N_45415,N_46994);
and U49573 (N_49573,N_45501,N_45928);
and U49574 (N_49574,N_46383,N_45741);
or U49575 (N_49575,N_46728,N_46488);
and U49576 (N_49576,N_47320,N_47337);
xnor U49577 (N_49577,N_47441,N_47287);
nor U49578 (N_49578,N_46255,N_47034);
nor U49579 (N_49579,N_45036,N_46188);
nor U49580 (N_49580,N_46565,N_46578);
nor U49581 (N_49581,N_46948,N_45360);
xnor U49582 (N_49582,N_47339,N_45623);
nor U49583 (N_49583,N_46269,N_45467);
xor U49584 (N_49584,N_45058,N_46522);
and U49585 (N_49585,N_47316,N_46572);
or U49586 (N_49586,N_45238,N_47238);
or U49587 (N_49587,N_45031,N_47283);
nor U49588 (N_49588,N_45734,N_46591);
or U49589 (N_49589,N_45776,N_45350);
nor U49590 (N_49590,N_45485,N_46989);
nor U49591 (N_49591,N_46313,N_47269);
and U49592 (N_49592,N_45728,N_46996);
and U49593 (N_49593,N_45372,N_45203);
and U49594 (N_49594,N_47316,N_45742);
nand U49595 (N_49595,N_46803,N_46413);
nor U49596 (N_49596,N_45518,N_46524);
nor U49597 (N_49597,N_45042,N_46611);
and U49598 (N_49598,N_47149,N_45281);
nand U49599 (N_49599,N_46065,N_45598);
and U49600 (N_49600,N_45187,N_46797);
and U49601 (N_49601,N_47219,N_46518);
xor U49602 (N_49602,N_46127,N_47206);
and U49603 (N_49603,N_45713,N_46021);
or U49604 (N_49604,N_45354,N_46270);
nor U49605 (N_49605,N_45052,N_46551);
and U49606 (N_49606,N_46758,N_45841);
and U49607 (N_49607,N_47165,N_46293);
nor U49608 (N_49608,N_47395,N_47094);
and U49609 (N_49609,N_45278,N_46240);
and U49610 (N_49610,N_45293,N_47143);
and U49611 (N_49611,N_46107,N_46848);
or U49612 (N_49612,N_46299,N_46070);
nand U49613 (N_49613,N_45120,N_47166);
nand U49614 (N_49614,N_45395,N_46432);
nor U49615 (N_49615,N_46276,N_46947);
or U49616 (N_49616,N_46869,N_46789);
nor U49617 (N_49617,N_45091,N_45184);
xor U49618 (N_49618,N_46603,N_47393);
and U49619 (N_49619,N_45109,N_46908);
nor U49620 (N_49620,N_47212,N_45966);
nand U49621 (N_49621,N_46700,N_47313);
nand U49622 (N_49622,N_45078,N_46963);
nor U49623 (N_49623,N_46902,N_46273);
xor U49624 (N_49624,N_45142,N_46837);
nand U49625 (N_49625,N_47427,N_45102);
nand U49626 (N_49626,N_45074,N_47378);
nor U49627 (N_49627,N_46842,N_46502);
or U49628 (N_49628,N_45644,N_45188);
xor U49629 (N_49629,N_45497,N_46570);
nor U49630 (N_49630,N_46567,N_45437);
xnor U49631 (N_49631,N_47494,N_47006);
xnor U49632 (N_49632,N_46126,N_46058);
xnor U49633 (N_49633,N_45278,N_46801);
or U49634 (N_49634,N_45049,N_45208);
nand U49635 (N_49635,N_46171,N_46584);
nand U49636 (N_49636,N_45715,N_45388);
xor U49637 (N_49637,N_46668,N_47038);
nor U49638 (N_49638,N_45821,N_46315);
and U49639 (N_49639,N_46054,N_46721);
and U49640 (N_49640,N_47216,N_45246);
nor U49641 (N_49641,N_47431,N_47378);
nand U49642 (N_49642,N_46736,N_45806);
nor U49643 (N_49643,N_46661,N_45454);
nor U49644 (N_49644,N_47011,N_47103);
nand U49645 (N_49645,N_46217,N_46609);
or U49646 (N_49646,N_45804,N_45932);
and U49647 (N_49647,N_45694,N_45366);
and U49648 (N_49648,N_46548,N_46838);
xnor U49649 (N_49649,N_45399,N_45823);
and U49650 (N_49650,N_47290,N_46921);
nand U49651 (N_49651,N_47460,N_47495);
nor U49652 (N_49652,N_46384,N_45117);
or U49653 (N_49653,N_47052,N_46872);
xnor U49654 (N_49654,N_47427,N_45359);
or U49655 (N_49655,N_46738,N_45278);
or U49656 (N_49656,N_46522,N_46384);
or U49657 (N_49657,N_45245,N_47335);
nand U49658 (N_49658,N_45346,N_45331);
and U49659 (N_49659,N_46399,N_45240);
and U49660 (N_49660,N_47320,N_45197);
nand U49661 (N_49661,N_45851,N_45196);
nor U49662 (N_49662,N_46960,N_45995);
nand U49663 (N_49663,N_45156,N_46789);
or U49664 (N_49664,N_45644,N_45234);
nor U49665 (N_49665,N_45176,N_47456);
nor U49666 (N_49666,N_46519,N_46107);
or U49667 (N_49667,N_46598,N_46826);
nor U49668 (N_49668,N_45390,N_46254);
nand U49669 (N_49669,N_46645,N_45632);
or U49670 (N_49670,N_45518,N_47420);
nor U49671 (N_49671,N_45097,N_46050);
nor U49672 (N_49672,N_46445,N_47068);
or U49673 (N_49673,N_46766,N_47457);
or U49674 (N_49674,N_46832,N_45302);
nor U49675 (N_49675,N_45996,N_46881);
nor U49676 (N_49676,N_46262,N_45790);
or U49677 (N_49677,N_46363,N_46198);
xnor U49678 (N_49678,N_45442,N_45194);
or U49679 (N_49679,N_45178,N_46161);
and U49680 (N_49680,N_45010,N_46524);
nand U49681 (N_49681,N_45452,N_47458);
xor U49682 (N_49682,N_46384,N_46006);
nand U49683 (N_49683,N_45913,N_45454);
nor U49684 (N_49684,N_47076,N_45271);
nand U49685 (N_49685,N_46033,N_45549);
xor U49686 (N_49686,N_47414,N_45026);
or U49687 (N_49687,N_45734,N_47441);
nor U49688 (N_49688,N_45673,N_45078);
and U49689 (N_49689,N_45105,N_46537);
nand U49690 (N_49690,N_46795,N_46066);
and U49691 (N_49691,N_45798,N_46770);
nor U49692 (N_49692,N_46092,N_47286);
nand U49693 (N_49693,N_46242,N_45118);
nor U49694 (N_49694,N_45827,N_45026);
and U49695 (N_49695,N_45565,N_47129);
and U49696 (N_49696,N_46838,N_46432);
and U49697 (N_49697,N_46356,N_46238);
nor U49698 (N_49698,N_46496,N_46742);
and U49699 (N_49699,N_46287,N_45524);
nor U49700 (N_49700,N_46949,N_46464);
xor U49701 (N_49701,N_47485,N_46116);
and U49702 (N_49702,N_46241,N_45390);
nor U49703 (N_49703,N_46129,N_45789);
and U49704 (N_49704,N_47391,N_45836);
nor U49705 (N_49705,N_45115,N_46821);
xnor U49706 (N_49706,N_45005,N_47288);
nand U49707 (N_49707,N_47227,N_46561);
or U49708 (N_49708,N_46354,N_46152);
or U49709 (N_49709,N_45204,N_46268);
or U49710 (N_49710,N_46879,N_46136);
or U49711 (N_49711,N_47277,N_45077);
nand U49712 (N_49712,N_46948,N_45866);
nand U49713 (N_49713,N_45385,N_47356);
xnor U49714 (N_49714,N_45251,N_46112);
nand U49715 (N_49715,N_46897,N_46267);
nand U49716 (N_49716,N_45900,N_45751);
and U49717 (N_49717,N_45276,N_45104);
or U49718 (N_49718,N_45008,N_45199);
and U49719 (N_49719,N_45683,N_46440);
nand U49720 (N_49720,N_45666,N_45768);
nor U49721 (N_49721,N_45040,N_46213);
or U49722 (N_49722,N_45248,N_47045);
nor U49723 (N_49723,N_46575,N_45828);
nand U49724 (N_49724,N_47428,N_45376);
nand U49725 (N_49725,N_45748,N_45046);
nor U49726 (N_49726,N_45657,N_46704);
nor U49727 (N_49727,N_46750,N_45579);
nand U49728 (N_49728,N_45633,N_47226);
nor U49729 (N_49729,N_45570,N_46923);
nor U49730 (N_49730,N_46287,N_45439);
xnor U49731 (N_49731,N_45496,N_47462);
nand U49732 (N_49732,N_47264,N_45859);
nand U49733 (N_49733,N_46879,N_45555);
or U49734 (N_49734,N_45125,N_45455);
and U49735 (N_49735,N_45068,N_46562);
or U49736 (N_49736,N_46692,N_47480);
or U49737 (N_49737,N_46758,N_46633);
nand U49738 (N_49738,N_45105,N_46149);
and U49739 (N_49739,N_46225,N_45821);
and U49740 (N_49740,N_45840,N_45431);
and U49741 (N_49741,N_46322,N_46832);
nor U49742 (N_49742,N_47316,N_45707);
xnor U49743 (N_49743,N_47021,N_47249);
xor U49744 (N_49744,N_46871,N_45722);
and U49745 (N_49745,N_46872,N_45957);
or U49746 (N_49746,N_45887,N_46506);
xnor U49747 (N_49747,N_46159,N_45715);
and U49748 (N_49748,N_46434,N_47203);
nand U49749 (N_49749,N_47087,N_46256);
and U49750 (N_49750,N_45633,N_45132);
nor U49751 (N_49751,N_45310,N_46641);
nand U49752 (N_49752,N_46174,N_45890);
or U49753 (N_49753,N_45963,N_45499);
or U49754 (N_49754,N_45250,N_47494);
nor U49755 (N_49755,N_45338,N_47425);
xor U49756 (N_49756,N_45946,N_45351);
and U49757 (N_49757,N_47069,N_46466);
or U49758 (N_49758,N_45672,N_45119);
and U49759 (N_49759,N_45289,N_46586);
nor U49760 (N_49760,N_45030,N_45638);
and U49761 (N_49761,N_45510,N_46842);
and U49762 (N_49762,N_45318,N_46961);
nor U49763 (N_49763,N_46238,N_46063);
nor U49764 (N_49764,N_45926,N_47032);
xor U49765 (N_49765,N_45593,N_45262);
nor U49766 (N_49766,N_47232,N_45960);
or U49767 (N_49767,N_47138,N_46553);
nor U49768 (N_49768,N_46814,N_45568);
or U49769 (N_49769,N_45145,N_47265);
nor U49770 (N_49770,N_47427,N_46647);
xor U49771 (N_49771,N_45751,N_46208);
and U49772 (N_49772,N_46676,N_47194);
and U49773 (N_49773,N_46547,N_47084);
and U49774 (N_49774,N_47479,N_45532);
nand U49775 (N_49775,N_45932,N_47432);
xor U49776 (N_49776,N_46957,N_45792);
or U49777 (N_49777,N_46817,N_45390);
nor U49778 (N_49778,N_47198,N_46293);
xor U49779 (N_49779,N_47416,N_46422);
nand U49780 (N_49780,N_46786,N_45095);
and U49781 (N_49781,N_46323,N_46000);
nand U49782 (N_49782,N_47090,N_46213);
xor U49783 (N_49783,N_46965,N_47418);
and U49784 (N_49784,N_45779,N_47197);
or U49785 (N_49785,N_45917,N_46438);
and U49786 (N_49786,N_45153,N_46844);
nand U49787 (N_49787,N_46769,N_45301);
or U49788 (N_49788,N_46906,N_46103);
xor U49789 (N_49789,N_45593,N_46437);
nand U49790 (N_49790,N_46296,N_47104);
nand U49791 (N_49791,N_45515,N_45711);
and U49792 (N_49792,N_45292,N_46124);
nor U49793 (N_49793,N_46937,N_46136);
and U49794 (N_49794,N_45332,N_47430);
xnor U49795 (N_49795,N_47483,N_45979);
or U49796 (N_49796,N_46359,N_45683);
nor U49797 (N_49797,N_45999,N_47278);
xnor U49798 (N_49798,N_46312,N_47328);
xor U49799 (N_49799,N_45656,N_46183);
nand U49800 (N_49800,N_45641,N_45832);
nor U49801 (N_49801,N_47017,N_46887);
or U49802 (N_49802,N_45918,N_47175);
nand U49803 (N_49803,N_47194,N_47411);
xor U49804 (N_49804,N_45852,N_46739);
nor U49805 (N_49805,N_46583,N_47336);
or U49806 (N_49806,N_46765,N_46166);
and U49807 (N_49807,N_45776,N_46231);
xnor U49808 (N_49808,N_47390,N_46352);
and U49809 (N_49809,N_46166,N_45777);
nor U49810 (N_49810,N_47112,N_46344);
and U49811 (N_49811,N_45361,N_45560);
xor U49812 (N_49812,N_45783,N_45539);
nor U49813 (N_49813,N_46222,N_46889);
and U49814 (N_49814,N_46302,N_46588);
and U49815 (N_49815,N_45678,N_45031);
xnor U49816 (N_49816,N_46874,N_46742);
or U49817 (N_49817,N_47214,N_45511);
nand U49818 (N_49818,N_45425,N_46922);
xor U49819 (N_49819,N_46380,N_47336);
nor U49820 (N_49820,N_47023,N_45243);
nand U49821 (N_49821,N_46898,N_47348);
nor U49822 (N_49822,N_45944,N_45313);
nor U49823 (N_49823,N_47379,N_46706);
xnor U49824 (N_49824,N_47062,N_45236);
nand U49825 (N_49825,N_47456,N_45303);
xnor U49826 (N_49826,N_46036,N_46014);
nor U49827 (N_49827,N_46744,N_46021);
xor U49828 (N_49828,N_46380,N_46593);
xor U49829 (N_49829,N_45939,N_45155);
nor U49830 (N_49830,N_46075,N_46899);
nor U49831 (N_49831,N_45718,N_45225);
nand U49832 (N_49832,N_45595,N_46191);
nand U49833 (N_49833,N_46228,N_45869);
xor U49834 (N_49834,N_46775,N_45734);
and U49835 (N_49835,N_47302,N_46323);
or U49836 (N_49836,N_45302,N_45738);
and U49837 (N_49837,N_45597,N_45256);
and U49838 (N_49838,N_46175,N_45685);
xor U49839 (N_49839,N_46523,N_45605);
nor U49840 (N_49840,N_45492,N_46056);
xor U49841 (N_49841,N_46051,N_46288);
nor U49842 (N_49842,N_45254,N_45368);
xor U49843 (N_49843,N_46804,N_45904);
xor U49844 (N_49844,N_45339,N_47369);
nor U49845 (N_49845,N_45991,N_45768);
and U49846 (N_49846,N_46471,N_47303);
nand U49847 (N_49847,N_46640,N_46525);
nand U49848 (N_49848,N_45842,N_46881);
and U49849 (N_49849,N_46601,N_45119);
xor U49850 (N_49850,N_45878,N_46179);
nor U49851 (N_49851,N_46065,N_45896);
or U49852 (N_49852,N_46664,N_45648);
and U49853 (N_49853,N_45218,N_47171);
nand U49854 (N_49854,N_46275,N_45198);
or U49855 (N_49855,N_46133,N_46885);
nand U49856 (N_49856,N_46363,N_45211);
nor U49857 (N_49857,N_45547,N_45319);
xnor U49858 (N_49858,N_47065,N_45333);
xor U49859 (N_49859,N_47462,N_47483);
nand U49860 (N_49860,N_46475,N_45266);
xnor U49861 (N_49861,N_46800,N_46940);
nor U49862 (N_49862,N_46072,N_45851);
and U49863 (N_49863,N_47392,N_47475);
or U49864 (N_49864,N_46141,N_46182);
nand U49865 (N_49865,N_47191,N_46179);
xnor U49866 (N_49866,N_46539,N_46097);
or U49867 (N_49867,N_46539,N_45798);
xnor U49868 (N_49868,N_45934,N_45640);
xor U49869 (N_49869,N_45157,N_46720);
nor U49870 (N_49870,N_46110,N_47332);
and U49871 (N_49871,N_47385,N_46963);
nand U49872 (N_49872,N_47286,N_46587);
nor U49873 (N_49873,N_46991,N_47370);
or U49874 (N_49874,N_45902,N_46091);
nand U49875 (N_49875,N_45157,N_46746);
and U49876 (N_49876,N_45872,N_45802);
and U49877 (N_49877,N_47004,N_46350);
and U49878 (N_49878,N_45042,N_46224);
nor U49879 (N_49879,N_45515,N_46278);
and U49880 (N_49880,N_47199,N_46022);
xnor U49881 (N_49881,N_46080,N_46412);
nand U49882 (N_49882,N_47351,N_46849);
xor U49883 (N_49883,N_46160,N_45331);
nand U49884 (N_49884,N_47374,N_47242);
nand U49885 (N_49885,N_46071,N_46075);
nor U49886 (N_49886,N_47296,N_46362);
or U49887 (N_49887,N_46932,N_47423);
xor U49888 (N_49888,N_47356,N_46443);
nor U49889 (N_49889,N_45733,N_45950);
and U49890 (N_49890,N_46609,N_46558);
and U49891 (N_49891,N_47086,N_47269);
or U49892 (N_49892,N_45816,N_45169);
or U49893 (N_49893,N_46222,N_45861);
nand U49894 (N_49894,N_45958,N_46829);
nor U49895 (N_49895,N_46844,N_46322);
xnor U49896 (N_49896,N_46520,N_45834);
nor U49897 (N_49897,N_45309,N_45341);
and U49898 (N_49898,N_46027,N_45339);
nor U49899 (N_49899,N_47495,N_47057);
nand U49900 (N_49900,N_46668,N_47447);
xnor U49901 (N_49901,N_46093,N_46511);
nor U49902 (N_49902,N_46774,N_45297);
xnor U49903 (N_49903,N_46422,N_46321);
nand U49904 (N_49904,N_45030,N_46290);
or U49905 (N_49905,N_46741,N_45828);
nor U49906 (N_49906,N_45817,N_45642);
and U49907 (N_49907,N_46489,N_46818);
nor U49908 (N_49908,N_46729,N_46774);
xor U49909 (N_49909,N_45309,N_46680);
or U49910 (N_49910,N_47423,N_45013);
nand U49911 (N_49911,N_47329,N_46760);
nor U49912 (N_49912,N_46414,N_46864);
nor U49913 (N_49913,N_46659,N_46071);
xor U49914 (N_49914,N_45611,N_45719);
nor U49915 (N_49915,N_45021,N_47471);
xnor U49916 (N_49916,N_46225,N_45005);
or U49917 (N_49917,N_45748,N_45692);
or U49918 (N_49918,N_47075,N_45812);
nor U49919 (N_49919,N_46434,N_46405);
nor U49920 (N_49920,N_45626,N_45899);
xor U49921 (N_49921,N_45383,N_46397);
nand U49922 (N_49922,N_46713,N_47496);
xor U49923 (N_49923,N_45629,N_46134);
nand U49924 (N_49924,N_47110,N_45007);
nor U49925 (N_49925,N_45401,N_46987);
xnor U49926 (N_49926,N_45934,N_45924);
nand U49927 (N_49927,N_45045,N_46783);
nand U49928 (N_49928,N_46165,N_46590);
nor U49929 (N_49929,N_45147,N_47317);
xnor U49930 (N_49930,N_46367,N_46521);
xor U49931 (N_49931,N_45323,N_45856);
nand U49932 (N_49932,N_47077,N_47405);
or U49933 (N_49933,N_47313,N_45021);
nor U49934 (N_49934,N_46064,N_47171);
nor U49935 (N_49935,N_46304,N_47087);
nor U49936 (N_49936,N_46782,N_46852);
xnor U49937 (N_49937,N_46520,N_45245);
and U49938 (N_49938,N_46254,N_47102);
or U49939 (N_49939,N_46476,N_47485);
nor U49940 (N_49940,N_46626,N_46459);
or U49941 (N_49941,N_45530,N_46603);
or U49942 (N_49942,N_45321,N_45027);
nand U49943 (N_49943,N_46427,N_46666);
xnor U49944 (N_49944,N_46216,N_46315);
nand U49945 (N_49945,N_45747,N_46931);
or U49946 (N_49946,N_46985,N_46138);
nand U49947 (N_49947,N_45273,N_47012);
and U49948 (N_49948,N_46690,N_45749);
and U49949 (N_49949,N_45489,N_45552);
xnor U49950 (N_49950,N_46193,N_46439);
xnor U49951 (N_49951,N_46268,N_45615);
nand U49952 (N_49952,N_47140,N_45734);
and U49953 (N_49953,N_46581,N_45420);
xnor U49954 (N_49954,N_47222,N_47088);
nand U49955 (N_49955,N_45408,N_46991);
or U49956 (N_49956,N_46379,N_45994);
and U49957 (N_49957,N_45946,N_47277);
nor U49958 (N_49958,N_46534,N_47425);
xnor U49959 (N_49959,N_46657,N_46163);
nand U49960 (N_49960,N_45877,N_46577);
or U49961 (N_49961,N_45451,N_47410);
xnor U49962 (N_49962,N_45069,N_46131);
and U49963 (N_49963,N_45819,N_47273);
xor U49964 (N_49964,N_46766,N_46564);
or U49965 (N_49965,N_45675,N_46737);
and U49966 (N_49966,N_45054,N_45105);
nor U49967 (N_49967,N_47245,N_46528);
and U49968 (N_49968,N_46430,N_46639);
xor U49969 (N_49969,N_47354,N_46942);
xor U49970 (N_49970,N_45036,N_46884);
nand U49971 (N_49971,N_45349,N_46615);
nand U49972 (N_49972,N_45387,N_46074);
and U49973 (N_49973,N_46758,N_45421);
or U49974 (N_49974,N_46597,N_47251);
nor U49975 (N_49975,N_45933,N_47055);
xor U49976 (N_49976,N_45578,N_45608);
or U49977 (N_49977,N_45071,N_46069);
and U49978 (N_49978,N_45917,N_46441);
nor U49979 (N_49979,N_45661,N_46625);
or U49980 (N_49980,N_46085,N_46896);
and U49981 (N_49981,N_46157,N_45264);
nand U49982 (N_49982,N_47198,N_45767);
or U49983 (N_49983,N_46052,N_45116);
nand U49984 (N_49984,N_46360,N_45335);
nand U49985 (N_49985,N_45885,N_46035);
or U49986 (N_49986,N_45499,N_47196);
or U49987 (N_49987,N_45345,N_47356);
xnor U49988 (N_49988,N_46563,N_45406);
nand U49989 (N_49989,N_46275,N_46531);
and U49990 (N_49990,N_46053,N_45956);
nor U49991 (N_49991,N_47210,N_47158);
or U49992 (N_49992,N_46608,N_46780);
or U49993 (N_49993,N_45873,N_47060);
nor U49994 (N_49994,N_46611,N_46123);
xnor U49995 (N_49995,N_46693,N_47463);
and U49996 (N_49996,N_45295,N_47238);
nor U49997 (N_49997,N_45115,N_47462);
nor U49998 (N_49998,N_46891,N_46989);
xnor U49999 (N_49999,N_45592,N_45284);
nand UO_0 (O_0,N_49435,N_47895);
nor UO_1 (O_1,N_48021,N_47631);
or UO_2 (O_2,N_48797,N_47643);
nand UO_3 (O_3,N_49897,N_49410);
nand UO_4 (O_4,N_49749,N_49629);
xnor UO_5 (O_5,N_49908,N_48512);
nand UO_6 (O_6,N_48206,N_48274);
xor UO_7 (O_7,N_48181,N_49670);
nand UO_8 (O_8,N_48649,N_48537);
xnor UO_9 (O_9,N_47970,N_49309);
xor UO_10 (O_10,N_49934,N_48524);
nand UO_11 (O_11,N_49449,N_47736);
xor UO_12 (O_12,N_48628,N_49927);
nor UO_13 (O_13,N_47977,N_48919);
and UO_14 (O_14,N_48927,N_49930);
and UO_15 (O_15,N_48024,N_49648);
or UO_16 (O_16,N_47755,N_49935);
xnor UO_17 (O_17,N_47764,N_48773);
or UO_18 (O_18,N_49282,N_49478);
or UO_19 (O_19,N_49948,N_47510);
nor UO_20 (O_20,N_48178,N_47839);
nor UO_21 (O_21,N_48627,N_47570);
nor UO_22 (O_22,N_48429,N_48017);
nor UO_23 (O_23,N_49769,N_48395);
or UO_24 (O_24,N_48025,N_48254);
or UO_25 (O_25,N_48172,N_48129);
nor UO_26 (O_26,N_48621,N_48258);
nor UO_27 (O_27,N_49466,N_48288);
nand UO_28 (O_28,N_48651,N_48584);
xnor UO_29 (O_29,N_48404,N_48626);
or UO_30 (O_30,N_48565,N_49365);
nand UO_31 (O_31,N_49151,N_49414);
nand UO_32 (O_32,N_48957,N_48353);
nand UO_33 (O_33,N_49078,N_49809);
and UO_34 (O_34,N_48569,N_49877);
and UO_35 (O_35,N_48606,N_49185);
or UO_36 (O_36,N_49924,N_47954);
xnor UO_37 (O_37,N_48022,N_48142);
or UO_38 (O_38,N_49024,N_48367);
or UO_39 (O_39,N_49967,N_48093);
xor UO_40 (O_40,N_49394,N_47518);
xor UO_41 (O_41,N_49689,N_48012);
and UO_42 (O_42,N_48096,N_49945);
or UO_43 (O_43,N_49440,N_47822);
nand UO_44 (O_44,N_49686,N_48414);
nand UO_45 (O_45,N_48387,N_48375);
nor UO_46 (O_46,N_48831,N_48819);
nor UO_47 (O_47,N_48771,N_49131);
nor UO_48 (O_48,N_48318,N_48098);
nor UO_49 (O_49,N_49687,N_48917);
xnor UO_50 (O_50,N_47703,N_49878);
or UO_51 (O_51,N_49933,N_47758);
xnor UO_52 (O_52,N_48668,N_49952);
nand UO_53 (O_53,N_48095,N_47765);
and UO_54 (O_54,N_48213,N_49541);
or UO_55 (O_55,N_47941,N_48370);
xor UO_56 (O_56,N_49103,N_49223);
and UO_57 (O_57,N_47516,N_48718);
xnor UO_58 (O_58,N_49326,N_49144);
nand UO_59 (O_59,N_48188,N_48184);
nand UO_60 (O_60,N_47918,N_49373);
xor UO_61 (O_61,N_49305,N_48862);
and UO_62 (O_62,N_48278,N_49795);
nor UO_63 (O_63,N_48466,N_49029);
or UO_64 (O_64,N_49545,N_49599);
nand UO_65 (O_65,N_48496,N_49148);
and UO_66 (O_66,N_49274,N_48008);
nand UO_67 (O_67,N_49882,N_49287);
nor UO_68 (O_68,N_49804,N_49358);
nor UO_69 (O_69,N_49928,N_48657);
nand UO_70 (O_70,N_49690,N_49829);
xor UO_71 (O_71,N_47932,N_49671);
nor UO_72 (O_72,N_48330,N_49441);
nand UO_73 (O_73,N_48492,N_47779);
xor UO_74 (O_74,N_49177,N_49846);
and UO_75 (O_75,N_48564,N_49985);
nand UO_76 (O_76,N_49790,N_49944);
nand UO_77 (O_77,N_48475,N_49354);
nor UO_78 (O_78,N_47921,N_48062);
nor UO_79 (O_79,N_49612,N_47744);
xor UO_80 (O_80,N_47863,N_49752);
nand UO_81 (O_81,N_49297,N_48337);
nor UO_82 (O_82,N_49322,N_48020);
or UO_83 (O_83,N_48754,N_48212);
xor UO_84 (O_84,N_49243,N_49107);
xnor UO_85 (O_85,N_48360,N_49861);
xor UO_86 (O_86,N_48167,N_48248);
nor UO_87 (O_87,N_49011,N_47590);
nor UO_88 (O_88,N_48854,N_49490);
xnor UO_89 (O_89,N_49813,N_48937);
nor UO_90 (O_90,N_49357,N_48638);
nand UO_91 (O_91,N_48694,N_49866);
xnor UO_92 (O_92,N_48063,N_49120);
or UO_93 (O_93,N_48764,N_47672);
and UO_94 (O_94,N_49815,N_49502);
xor UO_95 (O_95,N_47698,N_49579);
nand UO_96 (O_96,N_48958,N_48730);
or UO_97 (O_97,N_47547,N_49306);
xor UO_98 (O_98,N_47679,N_48637);
nand UO_99 (O_99,N_49471,N_48232);
nor UO_100 (O_100,N_49625,N_49097);
xnor UO_101 (O_101,N_48393,N_49841);
or UO_102 (O_102,N_47555,N_48320);
nor UO_103 (O_103,N_49539,N_49210);
xnor UO_104 (O_104,N_48572,N_49839);
nand UO_105 (O_105,N_48309,N_48364);
or UO_106 (O_106,N_49130,N_49637);
xor UO_107 (O_107,N_47794,N_48077);
and UO_108 (O_108,N_47811,N_48275);
nand UO_109 (O_109,N_47539,N_47580);
and UO_110 (O_110,N_48104,N_47842);
or UO_111 (O_111,N_49605,N_47599);
xor UO_112 (O_112,N_48186,N_48642);
or UO_113 (O_113,N_48590,N_49685);
xnor UO_114 (O_114,N_49404,N_49377);
nor UO_115 (O_115,N_49173,N_47857);
xnor UO_116 (O_116,N_49618,N_49255);
or UO_117 (O_117,N_49083,N_48090);
xnor UO_118 (O_118,N_49027,N_48298);
xor UO_119 (O_119,N_49562,N_48658);
xnor UO_120 (O_120,N_48160,N_49467);
and UO_121 (O_121,N_47520,N_47709);
xor UO_122 (O_122,N_49656,N_49868);
nor UO_123 (O_123,N_49634,N_49493);
nand UO_124 (O_124,N_48903,N_49482);
nor UO_125 (O_125,N_47629,N_49063);
nand UO_126 (O_126,N_49835,N_48978);
and UO_127 (O_127,N_47958,N_49273);
nand UO_128 (O_128,N_47912,N_49571);
xnor UO_129 (O_129,N_49267,N_49037);
and UO_130 (O_130,N_49742,N_49789);
and UO_131 (O_131,N_49724,N_47908);
or UO_132 (O_132,N_48749,N_47964);
nor UO_133 (O_133,N_47931,N_48949);
or UO_134 (O_134,N_47691,N_48257);
nor UO_135 (O_135,N_49094,N_49244);
or UO_136 (O_136,N_47620,N_49045);
nand UO_137 (O_137,N_48230,N_48951);
xnor UO_138 (O_138,N_48520,N_47846);
and UO_139 (O_139,N_48516,N_48366);
or UO_140 (O_140,N_48923,N_48980);
nor UO_141 (O_141,N_49258,N_48089);
and UO_142 (O_142,N_48117,N_48128);
and UO_143 (O_143,N_48305,N_48913);
nand UO_144 (O_144,N_49697,N_48945);
nand UO_145 (O_145,N_49484,N_48836);
and UO_146 (O_146,N_48264,N_49760);
xor UO_147 (O_147,N_49716,N_48681);
and UO_148 (O_148,N_48725,N_49201);
or UO_149 (O_149,N_47593,N_47852);
nor UO_150 (O_150,N_49225,N_47843);
and UO_151 (O_151,N_48620,N_49475);
or UO_152 (O_152,N_48780,N_48815);
and UO_153 (O_153,N_47609,N_47663);
nand UO_154 (O_154,N_49291,N_47572);
or UO_155 (O_155,N_48454,N_47925);
xnor UO_156 (O_156,N_47910,N_49891);
nand UO_157 (O_157,N_49238,N_47681);
xnor UO_158 (O_158,N_48632,N_47529);
nor UO_159 (O_159,N_49863,N_49737);
nor UO_160 (O_160,N_48374,N_48840);
nor UO_161 (O_161,N_49904,N_49628);
xnor UO_162 (O_162,N_48488,N_48449);
or UO_163 (O_163,N_47899,N_49822);
nand UO_164 (O_164,N_48165,N_48164);
xor UO_165 (O_165,N_48758,N_49668);
or UO_166 (O_166,N_48231,N_48607);
nand UO_167 (O_167,N_48436,N_47805);
xor UO_168 (O_168,N_48156,N_49343);
nor UO_169 (O_169,N_48721,N_49620);
and UO_170 (O_170,N_48333,N_48736);
nor UO_171 (O_171,N_47608,N_49818);
xor UO_172 (O_172,N_47583,N_48419);
and UO_173 (O_173,N_48245,N_49821);
nor UO_174 (O_174,N_48465,N_49270);
nand UO_175 (O_175,N_49033,N_47692);
nand UO_176 (O_176,N_49677,N_49926);
xnor UO_177 (O_177,N_48613,N_49438);
xnor UO_178 (O_178,N_49303,N_47731);
nor UO_179 (O_179,N_48445,N_48385);
and UO_180 (O_180,N_47951,N_49960);
nand UO_181 (O_181,N_49588,N_49591);
nand UO_182 (O_182,N_49346,N_48046);
nor UO_183 (O_183,N_47715,N_48768);
nand UO_184 (O_184,N_49575,N_48037);
nand UO_185 (O_185,N_48659,N_47773);
or UO_186 (O_186,N_48587,N_49044);
and UO_187 (O_187,N_49654,N_48265);
nand UO_188 (O_188,N_48940,N_49112);
or UO_189 (O_189,N_48479,N_49290);
xor UO_190 (O_190,N_48582,N_48125);
nand UO_191 (O_191,N_49920,N_49115);
or UO_192 (O_192,N_49419,N_49900);
xnor UO_193 (O_193,N_47659,N_49371);
xor UO_194 (O_194,N_48636,N_48507);
or UO_195 (O_195,N_49775,N_48676);
nand UO_196 (O_196,N_48571,N_48432);
xnor UO_197 (O_197,N_48502,N_49192);
nor UO_198 (O_198,N_47735,N_48625);
nand UO_199 (O_199,N_48542,N_49264);
nand UO_200 (O_200,N_47615,N_48224);
nand UO_201 (O_201,N_47834,N_48540);
or UO_202 (O_202,N_49307,N_49643);
or UO_203 (O_203,N_49778,N_48656);
xnor UO_204 (O_204,N_48312,N_49016);
nand UO_205 (O_205,N_48014,N_48050);
xor UO_206 (O_206,N_48556,N_48826);
xor UO_207 (O_207,N_49164,N_47651);
xnor UO_208 (O_208,N_48852,N_48757);
or UO_209 (O_209,N_48368,N_47640);
nor UO_210 (O_210,N_47861,N_49764);
or UO_211 (O_211,N_49046,N_47512);
xnor UO_212 (O_212,N_48929,N_49320);
and UO_213 (O_213,N_49401,N_48083);
or UO_214 (O_214,N_49222,N_48110);
or UO_215 (O_215,N_48990,N_48453);
nor UO_216 (O_216,N_48900,N_48292);
xnor UO_217 (O_217,N_49183,N_49785);
xor UO_218 (O_218,N_47678,N_49105);
and UO_219 (O_219,N_49771,N_49247);
and UO_220 (O_220,N_47553,N_49080);
xor UO_221 (O_221,N_48648,N_49108);
and UO_222 (O_222,N_47653,N_48591);
or UO_223 (O_223,N_49012,N_49568);
or UO_224 (O_224,N_48994,N_49970);
xor UO_225 (O_225,N_47716,N_49919);
or UO_226 (O_226,N_48873,N_48672);
and UO_227 (O_227,N_49458,N_49196);
and UO_228 (O_228,N_48661,N_49188);
xor UO_229 (O_229,N_48868,N_49992);
or UO_230 (O_230,N_48126,N_48055);
or UO_231 (O_231,N_47637,N_48944);
and UO_232 (O_232,N_48735,N_48772);
or UO_233 (O_233,N_48597,N_48839);
xor UO_234 (O_234,N_48127,N_49528);
nand UO_235 (O_235,N_48774,N_47563);
xor UO_236 (O_236,N_49036,N_47550);
or UO_237 (O_237,N_48443,N_48788);
or UO_238 (O_238,N_49205,N_48150);
nor UO_239 (O_239,N_49791,N_49199);
nor UO_240 (O_240,N_49334,N_48968);
nand UO_241 (O_241,N_47658,N_47819);
nor UO_242 (O_242,N_49405,N_48853);
nor UO_243 (O_243,N_49399,N_48697);
or UO_244 (O_244,N_48192,N_49022);
nand UO_245 (O_245,N_49598,N_47853);
or UO_246 (O_246,N_48609,N_49206);
nand UO_247 (O_247,N_49595,N_47976);
xnor UO_248 (O_248,N_48141,N_48881);
or UO_249 (O_249,N_48216,N_48557);
nor UO_250 (O_250,N_47638,N_48324);
or UO_251 (O_251,N_47519,N_48804);
or UO_252 (O_252,N_48252,N_49682);
nor UO_253 (O_253,N_49215,N_47848);
xor UO_254 (O_254,N_49460,N_47796);
nor UO_255 (O_255,N_49141,N_49503);
nor UO_256 (O_256,N_49086,N_49235);
nand UO_257 (O_257,N_47892,N_49540);
xor UO_258 (O_258,N_48904,N_49705);
and UO_259 (O_259,N_49720,N_49416);
nor UO_260 (O_260,N_49828,N_48781);
xnor UO_261 (O_261,N_49319,N_48568);
or UO_262 (O_262,N_49254,N_49982);
xor UO_263 (O_263,N_49234,N_49393);
xnor UO_264 (O_264,N_49492,N_47675);
and UO_265 (O_265,N_49481,N_49002);
or UO_266 (O_266,N_49756,N_47740);
and UO_267 (O_267,N_48936,N_48845);
nand UO_268 (O_268,N_47605,N_48247);
xnor UO_269 (O_269,N_47841,N_48468);
nand UO_270 (O_270,N_47575,N_49832);
nor UO_271 (O_271,N_49709,N_49125);
nor UO_272 (O_272,N_48218,N_49746);
and UO_273 (O_273,N_48974,N_49523);
xor UO_274 (O_274,N_48448,N_47567);
and UO_275 (O_275,N_48291,N_49759);
or UO_276 (O_276,N_49496,N_47614);
xnor UO_277 (O_277,N_48510,N_48876);
nor UO_278 (O_278,N_48846,N_49831);
xor UO_279 (O_279,N_49383,N_48808);
xnor UO_280 (O_280,N_49389,N_48041);
and UO_281 (O_281,N_47896,N_49614);
nand UO_282 (O_282,N_49413,N_47617);
nor UO_283 (O_283,N_49047,N_48194);
nor UO_284 (O_284,N_48146,N_47965);
or UO_285 (O_285,N_49655,N_47995);
and UO_286 (O_286,N_49772,N_48266);
xor UO_287 (O_287,N_47902,N_48240);
xor UO_288 (O_288,N_47780,N_47635);
and UO_289 (O_289,N_49691,N_48082);
nand UO_290 (O_290,N_49510,N_48560);
and UO_291 (O_291,N_48786,N_47699);
nand UO_292 (O_292,N_47726,N_49781);
nand UO_293 (O_293,N_49281,N_47771);
nor UO_294 (O_294,N_48158,N_47546);
or UO_295 (O_295,N_49814,N_49980);
xnor UO_296 (O_296,N_49547,N_49088);
xor UO_297 (O_297,N_48901,N_49896);
and UO_298 (O_298,N_48462,N_49996);
or UO_299 (O_299,N_49633,N_48065);
nor UO_300 (O_300,N_48261,N_47787);
xnor UO_301 (O_301,N_48902,N_49702);
and UO_302 (O_302,N_49607,N_49098);
or UO_303 (O_303,N_49852,N_48983);
nor UO_304 (O_304,N_47628,N_48838);
or UO_305 (O_305,N_48920,N_49888);
nand UO_306 (O_306,N_48982,N_49989);
or UO_307 (O_307,N_47752,N_48437);
xor UO_308 (O_308,N_49739,N_47751);
nand UO_309 (O_309,N_47850,N_48402);
and UO_310 (O_310,N_49061,N_49293);
nand UO_311 (O_311,N_48238,N_48227);
or UO_312 (O_312,N_48433,N_47756);
or UO_313 (O_313,N_48586,N_49727);
or UO_314 (O_314,N_48469,N_48807);
nor UO_315 (O_315,N_49239,N_49550);
or UO_316 (O_316,N_48262,N_49198);
or UO_317 (O_317,N_49143,N_48813);
xor UO_318 (O_318,N_47802,N_47793);
or UO_319 (O_319,N_49572,N_48765);
or UO_320 (O_320,N_49056,N_48283);
nand UO_321 (O_321,N_48480,N_48962);
and UO_322 (O_322,N_47810,N_48491);
and UO_323 (O_323,N_49251,N_47632);
nand UO_324 (O_324,N_47924,N_49608);
and UO_325 (O_325,N_48263,N_47530);
xor UO_326 (O_326,N_48744,N_49708);
nand UO_327 (O_327,N_49999,N_47923);
nand UO_328 (O_328,N_47586,N_49233);
xnor UO_329 (O_329,N_48267,N_49884);
xnor UO_330 (O_330,N_47565,N_48647);
and UO_331 (O_331,N_48223,N_48912);
and UO_332 (O_332,N_49096,N_49754);
xor UO_333 (O_333,N_48293,N_47634);
xor UO_334 (O_334,N_49736,N_49340);
nor UO_335 (O_335,N_47743,N_49990);
nand UO_336 (O_336,N_47992,N_48946);
xor UO_337 (O_337,N_49179,N_47683);
nor UO_338 (O_338,N_48755,N_49156);
or UO_339 (O_339,N_47584,N_49959);
nor UO_340 (O_340,N_49476,N_49623);
nor UO_341 (O_341,N_48769,N_48612);
and UO_342 (O_342,N_48376,N_49245);
or UO_343 (O_343,N_47619,N_48966);
or UO_344 (O_344,N_48600,N_48822);
nand UO_345 (O_345,N_48677,N_48378);
nand UO_346 (O_346,N_48099,N_48144);
xor UO_347 (O_347,N_49001,N_49892);
nand UO_348 (O_348,N_48134,N_47549);
and UO_349 (O_349,N_49963,N_47745);
nand UO_350 (O_350,N_48506,N_49583);
and UO_351 (O_351,N_48219,N_49956);
or UO_352 (O_352,N_48776,N_49338);
nor UO_353 (O_353,N_49780,N_48652);
and UO_354 (O_354,N_49717,N_49837);
nor UO_355 (O_355,N_49178,N_48828);
nor UO_356 (O_356,N_48517,N_49844);
or UO_357 (O_357,N_49909,N_47785);
or UO_358 (O_358,N_49248,N_47877);
and UO_359 (O_359,N_47621,N_48209);
or UO_360 (O_360,N_48728,N_47677);
or UO_361 (O_361,N_48019,N_49893);
or UO_362 (O_362,N_48015,N_48361);
xnor UO_363 (O_363,N_49228,N_48965);
xnor UO_364 (O_364,N_48031,N_47581);
or UO_365 (O_365,N_47666,N_49489);
and UO_366 (O_366,N_49402,N_47812);
xnor UO_367 (O_367,N_49847,N_49025);
or UO_368 (O_368,N_49069,N_48111);
xor UO_369 (O_369,N_48044,N_48422);
or UO_370 (O_370,N_49379,N_47646);
nor UO_371 (O_371,N_47823,N_48622);
and UO_372 (O_372,N_47509,N_49561);
xor UO_373 (O_373,N_48075,N_49220);
and UO_374 (O_374,N_49175,N_49856);
or UO_375 (O_375,N_48027,N_47737);
xnor UO_376 (O_376,N_49796,N_48185);
or UO_377 (O_377,N_47935,N_48703);
or UO_378 (O_378,N_49464,N_49000);
or UO_379 (O_379,N_49548,N_49227);
xor UO_380 (O_380,N_49745,N_47824);
nand UO_381 (O_381,N_48573,N_48752);
and UO_382 (O_382,N_49127,N_47858);
and UO_383 (O_383,N_48221,N_48601);
and UO_384 (O_384,N_49283,N_48120);
nand UO_385 (O_385,N_49741,N_48880);
nor UO_386 (O_386,N_49372,N_48335);
nand UO_387 (O_387,N_48973,N_47854);
nor UO_388 (O_388,N_47864,N_49819);
or UO_389 (O_389,N_49093,N_48325);
xor UO_390 (O_390,N_48269,N_48992);
nor UO_391 (O_391,N_49139,N_48887);
nand UO_392 (O_392,N_47955,N_48319);
and UO_393 (O_393,N_48855,N_48499);
nor UO_394 (O_394,N_48300,N_48394);
nor UO_395 (O_395,N_48566,N_48820);
and UO_396 (O_396,N_48714,N_49567);
nor UO_397 (O_397,N_49043,N_48430);
xor UO_398 (O_398,N_48030,N_49957);
nand UO_399 (O_399,N_49549,N_48236);
and UO_400 (O_400,N_47882,N_48745);
nand UO_401 (O_401,N_49816,N_48726);
nand UO_402 (O_402,N_49506,N_48210);
xnor UO_403 (O_403,N_49180,N_48425);
nor UO_404 (O_404,N_47574,N_47873);
xnor UO_405 (O_405,N_49437,N_47807);
nor UO_406 (O_406,N_49555,N_49894);
and UO_407 (O_407,N_48446,N_47952);
xnor UO_408 (O_408,N_49619,N_47832);
and UO_409 (O_409,N_48611,N_49327);
or UO_410 (O_410,N_47554,N_49104);
and UO_411 (O_411,N_49729,N_48787);
or UO_412 (O_412,N_49157,N_47985);
and UO_413 (O_413,N_47991,N_49678);
nor UO_414 (O_414,N_47792,N_48727);
or UO_415 (O_415,N_48123,N_49524);
and UO_416 (O_416,N_48960,N_48614);
nor UO_417 (O_417,N_47649,N_49278);
or UO_418 (O_418,N_47960,N_49838);
nor UO_419 (O_419,N_48369,N_47984);
nor UO_420 (O_420,N_49504,N_48934);
or UO_421 (O_421,N_49360,N_47983);
nor UO_422 (O_422,N_49289,N_48598);
or UO_423 (O_423,N_49145,N_47813);
xnor UO_424 (O_424,N_49627,N_48690);
nor UO_425 (O_425,N_48197,N_48190);
nor UO_426 (O_426,N_49895,N_48038);
xor UO_427 (O_427,N_48544,N_47871);
and UO_428 (O_428,N_48925,N_49182);
or UO_429 (O_429,N_49824,N_49129);
nand UO_430 (O_430,N_49323,N_47888);
xor UO_431 (O_431,N_48793,N_48058);
xor UO_432 (O_432,N_48678,N_48049);
nor UO_433 (O_433,N_49546,N_48938);
xnor UO_434 (O_434,N_48106,N_48629);
nor UO_435 (O_435,N_49172,N_47623);
nor UO_436 (O_436,N_49486,N_48977);
nand UO_437 (O_437,N_49596,N_48147);
xor UO_438 (O_438,N_47720,N_48006);
nand UO_439 (O_439,N_47898,N_48211);
nor UO_440 (O_440,N_49299,N_48102);
nand UO_441 (O_441,N_48316,N_48894);
or UO_442 (O_442,N_48961,N_49714);
nor UO_443 (O_443,N_49350,N_49738);
xor UO_444 (O_444,N_49911,N_49328);
nand UO_445 (O_445,N_47904,N_49774);
or UO_446 (O_446,N_48438,N_49973);
nor UO_447 (O_447,N_49301,N_49035);
xnor UO_448 (O_448,N_47835,N_48047);
nand UO_449 (O_449,N_47997,N_47930);
or UO_450 (O_450,N_49743,N_49966);
or UO_451 (O_451,N_47778,N_48034);
nor UO_452 (O_452,N_49565,N_47815);
and UO_453 (O_453,N_49191,N_47706);
or UO_454 (O_454,N_48578,N_48365);
nor UO_455 (O_455,N_48159,N_49994);
or UO_456 (O_456,N_49417,N_47685);
nand UO_457 (O_457,N_49519,N_48897);
nand UO_458 (O_458,N_48233,N_47790);
and UO_459 (O_459,N_47814,N_48545);
nor UO_460 (O_460,N_47561,N_48886);
or UO_461 (O_461,N_48170,N_47972);
or UO_462 (O_462,N_49298,N_49231);
xnor UO_463 (O_463,N_49190,N_49518);
nor UO_464 (O_464,N_49976,N_48281);
nand UO_465 (O_465,N_47502,N_49784);
and UO_466 (O_466,N_48381,N_49998);
nor UO_467 (O_467,N_48866,N_48051);
or UO_468 (O_468,N_48280,N_48931);
and UO_469 (O_469,N_47697,N_47601);
xor UO_470 (O_470,N_48187,N_47508);
xor UO_471 (O_471,N_48801,N_48798);
and UO_472 (O_472,N_49721,N_49110);
nand UO_473 (O_473,N_49805,N_47523);
and UO_474 (O_474,N_49390,N_48411);
xor UO_475 (O_475,N_49950,N_48554);
xnor UO_476 (O_476,N_47800,N_47630);
and UO_477 (O_477,N_48225,N_47624);
and UO_478 (O_478,N_49232,N_48883);
nor UO_479 (O_479,N_48914,N_48336);
and UO_480 (O_480,N_49874,N_48829);
and UO_481 (O_481,N_48205,N_48605);
xnor UO_482 (O_482,N_48687,N_47507);
or UO_483 (O_483,N_47934,N_49848);
and UO_484 (O_484,N_47782,N_47627);
or UO_485 (O_485,N_49257,N_49366);
nand UO_486 (O_486,N_49276,N_47939);
nand UO_487 (O_487,N_48701,N_48359);
or UO_488 (O_488,N_49733,N_49165);
nor UO_489 (O_489,N_48924,N_49060);
nor UO_490 (O_490,N_49403,N_47504);
and UO_491 (O_491,N_49463,N_48472);
or UO_492 (O_492,N_49520,N_48287);
or UO_493 (O_493,N_49246,N_48323);
or UO_494 (O_494,N_47937,N_47738);
and UO_495 (O_495,N_49770,N_48321);
or UO_496 (O_496,N_48011,N_47521);
nor UO_497 (O_497,N_49378,N_48279);
nand UO_498 (O_498,N_48410,N_48457);
nor UO_499 (O_499,N_47641,N_47710);
xnor UO_500 (O_500,N_49854,N_48229);
nor UO_501 (O_501,N_49237,N_48489);
and UO_502 (O_502,N_49421,N_49947);
nand UO_503 (O_503,N_48013,N_48713);
nor UO_504 (O_504,N_48139,N_49256);
nor UO_505 (O_505,N_49279,N_49324);
nand UO_506 (O_506,N_48532,N_48377);
or UO_507 (O_507,N_49376,N_49170);
or UO_508 (O_508,N_49138,N_48890);
nand UO_509 (O_509,N_49867,N_47999);
nor UO_510 (O_510,N_49858,N_47541);
nor UO_511 (O_511,N_49412,N_49452);
xnor UO_512 (O_512,N_48308,N_49300);
and UO_513 (O_513,N_47862,N_48149);
and UO_514 (O_514,N_48345,N_48342);
xnor UO_515 (O_515,N_48817,N_49474);
nand UO_516 (O_516,N_48138,N_49669);
nor UO_517 (O_517,N_48619,N_48553);
and UO_518 (O_518,N_47856,N_47500);
xor UO_519 (O_519,N_47543,N_49028);
xor UO_520 (O_520,N_48029,N_48947);
or UO_521 (O_521,N_49135,N_48097);
and UO_522 (O_522,N_48124,N_48969);
nand UO_523 (O_523,N_48487,N_48811);
and UO_524 (O_524,N_49054,N_48646);
or UO_525 (O_525,N_49755,N_48390);
nor UO_526 (O_526,N_47757,N_49385);
nand UO_527 (O_527,N_47585,N_48882);
or UO_528 (O_528,N_49154,N_48624);
and UO_529 (O_529,N_48250,N_48474);
or UO_530 (O_530,N_47990,N_47719);
xor UO_531 (O_531,N_49684,N_48284);
nor UO_532 (O_532,N_48864,N_49885);
nand UO_533 (O_533,N_48290,N_47531);
xor UO_534 (O_534,N_49375,N_48326);
xnor UO_535 (O_535,N_48220,N_48702);
nand UO_536 (O_536,N_48155,N_49594);
and UO_537 (O_537,N_49589,N_47943);
nand UO_538 (O_538,N_47540,N_49674);
or UO_539 (O_539,N_47616,N_48416);
nor UO_540 (O_540,N_49940,N_48533);
xor UO_541 (O_541,N_49498,N_47618);
nor UO_542 (O_542,N_48693,N_49101);
xor UO_543 (O_543,N_49681,N_48068);
xnor UO_544 (O_544,N_48354,N_49133);
xor UO_545 (O_545,N_47676,N_49075);
nand UO_546 (O_546,N_48711,N_47728);
xor UO_547 (O_547,N_48076,N_48892);
and UO_548 (O_548,N_48379,N_49337);
xor UO_549 (O_549,N_48666,N_49734);
or UO_550 (O_550,N_49286,N_48498);
nand UO_551 (O_551,N_47544,N_47747);
and UO_552 (O_552,N_48641,N_49032);
or UO_553 (O_553,N_48331,N_48157);
nand UO_554 (O_554,N_48592,N_48975);
and UO_555 (O_555,N_49398,N_48806);
nor UO_556 (O_556,N_49149,N_48870);
and UO_557 (O_557,N_48271,N_48515);
and UO_558 (O_558,N_48135,N_48692);
nand UO_559 (O_559,N_47696,N_48355);
and UO_560 (O_560,N_48567,N_49067);
or UO_561 (O_561,N_48760,N_48650);
and UO_562 (O_562,N_47535,N_48372);
nand UO_563 (O_563,N_47868,N_49483);
nor UO_564 (O_564,N_48576,N_47859);
and UO_565 (O_565,N_48163,N_49590);
or UO_566 (O_566,N_48905,N_49470);
and UO_567 (O_567,N_47922,N_49962);
xnor UO_568 (O_568,N_48273,N_49213);
nor UO_569 (O_569,N_49269,N_48101);
and UO_570 (O_570,N_48195,N_49650);
or UO_571 (O_571,N_48843,N_48338);
xnor UO_572 (O_572,N_49696,N_49925);
nand UO_573 (O_573,N_47573,N_47684);
nand UO_574 (O_574,N_49014,N_48717);
or UO_575 (O_575,N_48400,N_49429);
nor UO_576 (O_576,N_49204,N_49522);
nor UO_577 (O_577,N_47725,N_48151);
xnor UO_578 (O_578,N_49997,N_48954);
nor UO_579 (O_579,N_48086,N_49788);
and UO_580 (O_580,N_49763,N_47926);
and UO_581 (O_581,N_48918,N_49532);
or UO_582 (O_582,N_48667,N_48500);
nor UO_583 (O_583,N_49609,N_48534);
or UO_584 (O_584,N_47996,N_47956);
or UO_585 (O_585,N_49645,N_48204);
nand UO_586 (O_586,N_48669,N_49272);
nor UO_587 (O_587,N_49352,N_49160);
nand UO_588 (O_588,N_47712,N_48879);
nor UO_589 (O_589,N_47761,N_47947);
and UO_590 (O_590,N_48634,N_48546);
nand UO_591 (O_591,N_48130,N_48464);
nand UO_592 (O_592,N_48683,N_48893);
or UO_593 (O_593,N_47946,N_49526);
or UO_594 (O_594,N_48493,N_48176);
nor UO_595 (O_595,N_49631,N_48057);
nand UO_596 (O_596,N_48921,N_47526);
and UO_597 (O_597,N_48527,N_49560);
nor UO_598 (O_598,N_49049,N_49806);
xor UO_599 (O_599,N_49021,N_49638);
xnor UO_600 (O_600,N_49794,N_48481);
nand UO_601 (O_601,N_48915,N_47915);
or UO_602 (O_602,N_47671,N_47872);
nor UO_603 (O_603,N_49969,N_49516);
nor UO_604 (O_604,N_48835,N_48109);
nor UO_605 (O_605,N_49530,N_48173);
or UO_606 (O_606,N_49679,N_48816);
or UO_607 (O_607,N_47969,N_48989);
nand UO_608 (O_608,N_49381,N_48299);
xnor UO_609 (O_609,N_49345,N_49428);
and UO_610 (O_610,N_48964,N_47821);
nand UO_611 (O_611,N_48002,N_48698);
xnor UO_612 (O_612,N_47538,N_49296);
or UO_613 (O_613,N_49166,N_48574);
nand UO_614 (O_614,N_48583,N_48078);
and UO_615 (O_615,N_49517,N_48952);
nor UO_616 (O_616,N_47718,N_47905);
and UO_617 (O_617,N_49731,N_49744);
nand UO_618 (O_618,N_48132,N_48955);
nand UO_619 (O_619,N_49811,N_48237);
or UO_620 (O_620,N_49833,N_48070);
xor UO_621 (O_621,N_48743,N_48373);
and UO_622 (O_622,N_47766,N_47986);
nor UO_623 (O_623,N_49604,N_47639);
xor UO_624 (O_624,N_48789,N_49747);
nor UO_625 (O_625,N_48043,N_48802);
and UO_626 (O_626,N_49860,N_48630);
and UO_627 (O_627,N_48140,N_48891);
and UO_628 (O_628,N_49875,N_48148);
and UO_629 (O_629,N_47881,N_49751);
or UO_630 (O_630,N_49673,N_48451);
nand UO_631 (O_631,N_49573,N_47597);
nand UO_632 (O_632,N_48707,N_49265);
or UO_633 (O_633,N_49701,N_49587);
nand UO_634 (O_634,N_49117,N_49602);
nand UO_635 (O_635,N_48501,N_49013);
nor UO_636 (O_636,N_47594,N_47569);
xnor UO_637 (O_637,N_47749,N_49783);
and UO_638 (O_638,N_48536,N_48682);
nor UO_639 (O_639,N_48654,N_49451);
and UO_640 (O_640,N_48007,N_49341);
nor UO_641 (O_641,N_49842,N_48091);
nand UO_642 (O_642,N_49912,N_49941);
and UO_643 (O_643,N_47760,N_47971);
nand UO_644 (O_644,N_48950,N_48114);
xnor UO_645 (O_645,N_47748,N_49040);
nor UO_646 (O_646,N_49122,N_48052);
nand UO_647 (O_647,N_49004,N_49830);
or UO_648 (O_648,N_48551,N_48617);
nor UO_649 (O_649,N_49066,N_49800);
xor UO_650 (O_650,N_49750,N_48033);
nand UO_651 (O_651,N_49740,N_49675);
nand UO_652 (O_652,N_48009,N_47829);
and UO_653 (O_653,N_48972,N_49827);
and UO_654 (O_654,N_48971,N_49787);
or UO_655 (O_655,N_48710,N_49983);
xnor UO_656 (O_656,N_48984,N_49597);
xnor UO_657 (O_657,N_47633,N_49803);
nor UO_658 (O_658,N_48979,N_47998);
or UO_659 (O_659,N_49472,N_48304);
or UO_660 (O_660,N_47897,N_48018);
xnor UO_661 (O_661,N_49556,N_48001);
nand UO_662 (O_662,N_49889,N_49162);
nor UO_663 (O_663,N_48442,N_49748);
nor UO_664 (O_664,N_48426,N_48933);
nor UO_665 (O_665,N_48827,N_49621);
and UO_666 (O_666,N_48334,N_49706);
xnor UO_667 (O_667,N_48332,N_49817);
xor UO_668 (O_668,N_47528,N_49488);
xor UO_669 (O_669,N_48388,N_48531);
and UO_670 (O_670,N_49387,N_48242);
or UO_671 (O_671,N_48778,N_48674);
and UO_672 (O_672,N_48228,N_48403);
xor UO_673 (O_673,N_49348,N_48746);
and UO_674 (O_674,N_48133,N_47704);
xnor UO_675 (O_675,N_48100,N_47808);
or UO_676 (O_676,N_49534,N_48276);
or UO_677 (O_677,N_48460,N_49053);
and UO_678 (O_678,N_48671,N_47688);
nand UO_679 (O_679,N_49195,N_48664);
nor UO_680 (O_680,N_49719,N_47517);
or UO_681 (O_681,N_49121,N_48032);
and UO_682 (O_682,N_48633,N_49055);
nor UO_683 (O_683,N_48131,N_47913);
and UO_684 (O_684,N_49544,N_47917);
xor UO_685 (O_685,N_49444,N_49186);
and UO_686 (O_686,N_49664,N_49434);
nor UO_687 (O_687,N_48152,N_48296);
xor UO_688 (O_688,N_48039,N_48993);
or UO_689 (O_689,N_47506,N_49559);
xor UO_690 (O_690,N_49552,N_47536);
or UO_691 (O_691,N_48653,N_47789);
nand UO_692 (O_692,N_48358,N_49917);
or UO_693 (O_693,N_49042,N_49427);
nand UO_694 (O_694,N_49667,N_49006);
or UO_695 (O_695,N_48581,N_47665);
or UO_696 (O_696,N_47820,N_47588);
and UO_697 (O_697,N_48618,N_47514);
nor UO_698 (O_698,N_48663,N_48405);
nor UO_699 (O_699,N_48249,N_48311);
xnor UO_700 (O_700,N_49777,N_47603);
nor UO_701 (O_701,N_48616,N_47722);
or UO_702 (O_702,N_47929,N_48767);
nand UO_703 (O_703,N_49420,N_49132);
nand UO_704 (O_704,N_48171,N_48246);
nand UO_705 (O_705,N_49711,N_47566);
or UO_706 (O_706,N_49735,N_48759);
and UO_707 (O_707,N_49280,N_49840);
nand UO_708 (O_708,N_47532,N_49563);
nor UO_709 (O_709,N_47669,N_47524);
xnor UO_710 (O_710,N_47711,N_49038);
nand UO_711 (O_711,N_49657,N_49659);
xor UO_712 (O_712,N_49163,N_47648);
nor UO_713 (O_713,N_49361,N_49872);
xor UO_714 (O_714,N_48538,N_49161);
nand UO_715 (O_715,N_48175,N_49072);
or UO_716 (O_716,N_48241,N_49184);
xor UO_717 (O_717,N_49616,N_48777);
and UO_718 (O_718,N_48577,N_49007);
nand UO_719 (O_719,N_48907,N_47894);
or UO_720 (O_720,N_49136,N_47587);
nor UO_721 (O_721,N_47979,N_49302);
or UO_722 (O_722,N_48930,N_49447);
or UO_723 (O_723,N_49810,N_49635);
or UO_724 (O_724,N_49020,N_48753);
or UO_725 (O_725,N_47763,N_49142);
nand UO_726 (O_726,N_47741,N_49003);
nor UO_727 (O_727,N_48286,N_49836);
nor UO_728 (O_728,N_49501,N_49639);
nor UO_729 (O_729,N_48908,N_49986);
nor UO_730 (O_730,N_49181,N_49495);
and UO_731 (O_731,N_48409,N_48511);
nand UO_732 (O_732,N_49988,N_49491);
xor UO_733 (O_733,N_49356,N_48199);
nor UO_734 (O_734,N_48935,N_47909);
and UO_735 (O_735,N_49041,N_47564);
xnor UO_736 (O_736,N_49937,N_48715);
xor UO_737 (O_737,N_49531,N_49951);
and UO_738 (O_738,N_47714,N_49355);
and UO_739 (O_739,N_49423,N_49676);
or UO_740 (O_740,N_49432,N_48116);
nand UO_741 (O_741,N_48217,N_48196);
xor UO_742 (O_742,N_49092,N_47527);
and UO_743 (O_743,N_49666,N_48738);
nand UO_744 (O_744,N_49155,N_49624);
and UO_745 (O_745,N_49622,N_48795);
nor UO_746 (O_746,N_47886,N_48504);
nor UO_747 (O_747,N_47582,N_49446);
xor UO_748 (O_748,N_48356,N_49870);
xor UO_749 (O_749,N_49946,N_48732);
xor UO_750 (O_750,N_48085,N_49353);
and UO_751 (O_751,N_48483,N_49406);
or UO_752 (O_752,N_48963,N_49536);
and UO_753 (O_753,N_48575,N_48169);
nor UO_754 (O_754,N_48396,N_47717);
or UO_755 (O_755,N_47933,N_48685);
or UO_756 (O_756,N_49152,N_49415);
nor UO_757 (O_757,N_48328,N_49411);
xnor UO_758 (O_758,N_48635,N_48401);
xnor UO_759 (O_759,N_49261,N_49647);
and UO_760 (O_760,N_48244,N_48910);
xor UO_761 (O_761,N_48067,N_47993);
and UO_762 (O_762,N_48412,N_48851);
and UO_763 (O_763,N_47826,N_49134);
nand UO_764 (O_764,N_49901,N_48108);
or UO_765 (O_765,N_47795,N_49207);
and UO_766 (O_766,N_48036,N_49758);
nand UO_767 (O_767,N_48985,N_47739);
and UO_768 (O_768,N_49074,N_49242);
nor UO_769 (O_769,N_48561,N_48485);
and UO_770 (O_770,N_49344,N_47901);
and UO_771 (O_771,N_48799,N_49903);
or UO_772 (O_772,N_47533,N_47818);
nor UO_773 (O_773,N_48644,N_48307);
or UO_774 (O_774,N_47959,N_48662);
xnor UO_775 (O_775,N_47963,N_48215);
nand UO_776 (O_776,N_49543,N_48115);
nor UO_777 (O_777,N_47613,N_48987);
nor UO_778 (O_778,N_49230,N_49294);
xor UO_779 (O_779,N_48850,N_49663);
and UO_780 (O_780,N_47880,N_49396);
nand UO_781 (O_781,N_48074,N_49017);
nand UO_782 (O_782,N_48302,N_48408);
or UO_783 (O_783,N_47602,N_47768);
nor UO_784 (O_784,N_48023,N_49030);
or UO_785 (O_785,N_49408,N_49923);
nor UO_786 (O_786,N_48800,N_48858);
xnor UO_787 (O_787,N_49487,N_47838);
or UO_788 (O_788,N_49922,N_48756);
or UO_789 (O_789,N_48731,N_48847);
nor UO_790 (O_790,N_48783,N_48035);
and UO_791 (O_791,N_47890,N_48340);
nand UO_792 (O_792,N_49445,N_49918);
or UO_793 (O_793,N_49424,N_47962);
and UO_794 (O_794,N_49692,N_48832);
nand UO_795 (O_795,N_47828,N_49250);
or UO_796 (O_796,N_47883,N_48392);
nand UO_797 (O_797,N_49766,N_48825);
or UO_798 (O_798,N_49845,N_49525);
xnor UO_799 (O_799,N_48207,N_49574);
xnor UO_800 (O_800,N_48877,N_49140);
xor UO_801 (O_801,N_49553,N_48494);
xor UO_802 (O_802,N_47874,N_48967);
or UO_803 (O_803,N_49116,N_49958);
xnor UO_804 (O_804,N_48926,N_48471);
and UO_805 (O_805,N_49019,N_48785);
xor UO_806 (O_806,N_47576,N_49266);
xnor UO_807 (O_807,N_49641,N_48704);
and UO_808 (O_808,N_47844,N_48830);
nor UO_809 (O_809,N_47791,N_49167);
or UO_810 (O_810,N_47604,N_49465);
xnor UO_811 (O_811,N_47689,N_47690);
or UO_812 (O_812,N_49613,N_48686);
nand UO_813 (O_813,N_49216,N_48589);
or UO_814 (O_814,N_49277,N_47982);
or UO_815 (O_815,N_49802,N_48739);
xor UO_816 (O_816,N_48243,N_47799);
and UO_817 (O_817,N_49189,N_49582);
xnor UO_818 (O_818,N_49159,N_49932);
nand UO_819 (O_819,N_49584,N_49823);
xor UO_820 (O_820,N_47849,N_48234);
nand UO_821 (O_821,N_47837,N_48040);
and UO_822 (O_822,N_48282,N_47695);
nand UO_823 (O_823,N_48505,N_49325);
or UO_824 (O_824,N_48593,N_49249);
or UO_825 (O_825,N_48665,N_49529);
nor UO_826 (O_826,N_49494,N_49095);
and UO_827 (O_827,N_48081,N_48239);
and UO_828 (O_828,N_49214,N_48137);
and UO_829 (O_829,N_49812,N_49048);
nor UO_830 (O_830,N_47723,N_48053);
nand UO_831 (O_831,N_47562,N_49153);
or UO_832 (O_832,N_49626,N_48547);
xnor UO_833 (O_833,N_48878,N_49782);
and UO_834 (O_834,N_48675,N_47705);
nand UO_835 (O_835,N_49513,N_49336);
nand UO_836 (O_836,N_49695,N_47557);
nor UO_837 (O_837,N_48193,N_49704);
and UO_838 (O_838,N_48389,N_48497);
nand UO_839 (O_839,N_49859,N_49462);
and UO_840 (O_840,N_47957,N_48362);
and UO_841 (O_841,N_49712,N_49409);
nor UO_842 (O_842,N_49569,N_48486);
or UO_843 (O_843,N_49557,N_47801);
nor UO_844 (O_844,N_49975,N_49732);
and UO_845 (O_845,N_49068,N_49331);
xor UO_846 (O_846,N_49241,N_48708);
nor UO_847 (O_847,N_49793,N_48059);
or UO_848 (O_848,N_47967,N_48603);
or UO_849 (O_849,N_47702,N_47652);
nor UO_850 (O_850,N_48235,N_48595);
or UO_851 (O_851,N_48841,N_48720);
or UO_852 (O_852,N_48872,N_48867);
xor UO_853 (O_853,N_48253,N_49661);
nor UO_854 (O_854,N_47730,N_48885);
nor UO_855 (O_855,N_48997,N_49318);
nor UO_856 (O_856,N_49100,N_47713);
xnor UO_857 (O_857,N_49422,N_47707);
nand UO_858 (O_858,N_49615,N_48803);
xnor UO_859 (O_859,N_48303,N_48942);
and UO_860 (O_860,N_47515,N_48559);
and UO_861 (O_861,N_47578,N_48450);
nor UO_862 (O_862,N_48088,N_48860);
and UO_863 (O_863,N_49085,N_49187);
nand UO_864 (O_864,N_49776,N_47680);
nand UO_865 (O_865,N_47579,N_48072);
and UO_866 (O_866,N_49059,N_48723);
or UO_867 (O_867,N_47545,N_49694);
and UO_868 (O_868,N_47827,N_48999);
or UO_869 (O_869,N_47889,N_47855);
nand UO_870 (O_870,N_49535,N_48585);
nor UO_871 (O_871,N_48645,N_49473);
or UO_872 (O_872,N_48875,N_49586);
nand UO_873 (O_873,N_48154,N_48898);
and UO_874 (O_874,N_48255,N_48779);
and UO_875 (O_875,N_49984,N_47595);
and UO_876 (O_876,N_49109,N_49174);
xor UO_877 (O_877,N_48643,N_47978);
nor UO_878 (O_878,N_47729,N_48837);
nand UO_879 (O_879,N_48784,N_48529);
nand UO_880 (O_880,N_47980,N_47927);
xnor UO_881 (O_881,N_48610,N_48064);
and UO_882 (O_882,N_49570,N_48191);
xnor UO_883 (O_883,N_48514,N_49899);
or UO_884 (O_884,N_48640,N_49512);
nor UO_885 (O_885,N_48198,N_49538);
xor UO_886 (O_886,N_49707,N_49370);
xnor UO_887 (O_887,N_48884,N_48418);
nand UO_888 (O_888,N_48823,N_48639);
xor UO_889 (O_889,N_47598,N_48796);
or UO_890 (O_890,N_48094,N_48350);
nand UO_891 (O_891,N_49367,N_48660);
and UO_892 (O_892,N_48161,N_49857);
nor UO_893 (O_893,N_48673,N_49079);
and UO_894 (O_894,N_48004,N_48916);
nand UO_895 (O_895,N_48200,N_49585);
xnor UO_896 (O_896,N_48048,N_48528);
nand UO_897 (O_897,N_49580,N_48087);
nand UO_898 (O_898,N_47622,N_47875);
or UO_899 (O_899,N_48523,N_49688);
nand UO_900 (O_900,N_47840,N_48112);
xnor UO_901 (O_901,N_47987,N_49862);
nand UO_902 (O_902,N_49527,N_49315);
nand UO_903 (O_903,N_49137,N_49603);
or UO_904 (O_904,N_48742,N_49906);
xnor UO_905 (O_905,N_49577,N_48071);
and UO_906 (O_906,N_48397,N_49200);
nand UO_907 (O_907,N_48136,N_47907);
xnor UO_908 (O_908,N_49114,N_47750);
and UO_909 (O_909,N_49699,N_49057);
or UO_910 (O_910,N_49359,N_48363);
nand UO_911 (O_911,N_48821,N_47968);
and UO_912 (O_912,N_48346,N_49425);
nand UO_913 (O_913,N_49073,N_49902);
nor UO_914 (O_914,N_48766,N_48339);
xnor UO_915 (O_915,N_48084,N_49786);
and UO_916 (O_916,N_47953,N_48459);
nand UO_917 (O_917,N_49683,N_49119);
nand UO_918 (O_918,N_49268,N_48503);
or UO_919 (O_919,N_48444,N_48016);
and UO_920 (O_920,N_48079,N_49564);
nor UO_921 (O_921,N_49380,N_49147);
and UO_922 (O_922,N_47727,N_49218);
and UO_923 (O_923,N_47655,N_49508);
nor UO_924 (O_924,N_49194,N_49312);
or UO_925 (O_925,N_47988,N_48272);
nor UO_926 (O_926,N_47804,N_48709);
or UO_927 (O_927,N_48042,N_48810);
nand UO_928 (O_928,N_49977,N_48509);
or UO_929 (O_929,N_48526,N_48105);
xor UO_930 (O_930,N_48548,N_48427);
or UO_931 (O_931,N_49713,N_48382);
and UO_932 (O_932,N_49202,N_48301);
nor UO_933 (O_933,N_48179,N_49600);
xnor UO_934 (O_934,N_49349,N_49965);
or UO_935 (O_935,N_47974,N_47833);
and UO_936 (O_936,N_49384,N_49386);
and UO_937 (O_937,N_48734,N_49005);
or UO_938 (O_938,N_48182,N_48719);
and UO_939 (O_939,N_49168,N_49392);
nor UO_940 (O_940,N_48380,N_49855);
or UO_941 (O_941,N_49426,N_49039);
nand UO_942 (O_942,N_49369,N_49514);
nand UO_943 (O_943,N_49853,N_49362);
nand UO_944 (O_944,N_49128,N_47885);
nand UO_945 (O_945,N_49461,N_48762);
nor UO_946 (O_946,N_47942,N_48716);
or UO_947 (O_947,N_49652,N_49881);
and UO_948 (O_948,N_48424,N_48570);
xor UO_949 (O_949,N_48168,N_49873);
nor UO_950 (O_950,N_49456,N_48490);
xnor UO_951 (O_951,N_47797,N_49942);
xor UO_952 (O_952,N_47724,N_49453);
or UO_953 (O_953,N_49321,N_47577);
and UO_954 (O_954,N_48834,N_47571);
or UO_955 (O_955,N_49391,N_48270);
nor UO_956 (O_956,N_47591,N_47798);
nor UO_957 (O_957,N_49773,N_47803);
nor UO_958 (O_958,N_47625,N_48740);
xnor UO_959 (O_959,N_48696,N_49448);
nor UO_960 (O_960,N_48809,N_49665);
and UO_961 (O_961,N_47664,N_48431);
xnor UO_962 (O_962,N_48391,N_49578);
and UO_963 (O_963,N_49335,N_48045);
or UO_964 (O_964,N_49219,N_49710);
or UO_965 (O_965,N_48113,N_48588);
or UO_966 (O_966,N_49253,N_47611);
xor UO_967 (O_967,N_47700,N_49026);
xor UO_968 (O_968,N_47733,N_47626);
xnor UO_969 (O_969,N_48535,N_48222);
or UO_970 (O_970,N_49089,N_49090);
and UO_971 (O_971,N_49015,N_48495);
and UO_972 (O_972,N_49680,N_48107);
nor UO_973 (O_973,N_49480,N_48313);
or UO_974 (O_974,N_48423,N_48177);
or UO_975 (O_975,N_48162,N_49397);
or UO_976 (O_976,N_49850,N_47560);
nor UO_977 (O_977,N_48986,N_48413);
or UO_978 (O_978,N_49106,N_48259);
xor UO_979 (O_979,N_48899,N_49723);
xnor UO_980 (O_980,N_49052,N_48608);
xnor UO_981 (O_981,N_49649,N_48599);
nand UO_982 (O_982,N_48909,N_47775);
xnor UO_983 (O_983,N_49558,N_48343);
xor UO_984 (O_984,N_48814,N_49929);
nand UO_985 (O_985,N_48297,N_48751);
or UO_986 (O_986,N_48824,N_48763);
nand UO_987 (O_987,N_49768,N_48005);
nor UO_988 (O_988,N_48420,N_48202);
nand UO_989 (O_989,N_49864,N_47940);
xnor UO_990 (O_990,N_48470,N_48775);
nand UO_991 (O_991,N_49799,N_49158);
xnor UO_992 (O_992,N_47656,N_48277);
and UO_993 (O_993,N_47674,N_48737);
or UO_994 (O_994,N_48579,N_48699);
or UO_995 (O_995,N_47650,N_47936);
and UO_996 (O_996,N_47642,N_49395);
and UO_997 (O_997,N_49009,N_48513);
and UO_998 (O_998,N_47670,N_49820);
and UO_999 (O_999,N_48407,N_47701);
xnor UO_1000 (O_1000,N_49757,N_49521);
nand UO_1001 (O_1001,N_49064,N_48174);
nor UO_1002 (O_1002,N_49949,N_49418);
or UO_1003 (O_1003,N_48519,N_48289);
nor UO_1004 (O_1004,N_49779,N_49454);
or UO_1005 (O_1005,N_49347,N_49382);
or UO_1006 (O_1006,N_47537,N_48530);
nor UO_1007 (O_1007,N_49275,N_48791);
xor UO_1008 (O_1008,N_49761,N_48026);
xor UO_1009 (O_1009,N_49436,N_49077);
xnor UO_1010 (O_1010,N_49658,N_49450);
xor UO_1011 (O_1011,N_48294,N_48056);
or UO_1012 (O_1012,N_47687,N_49111);
nand UO_1013 (O_1013,N_47596,N_49808);
or UO_1014 (O_1014,N_48434,N_49798);
nor UO_1015 (O_1015,N_47654,N_49825);
and UO_1016 (O_1016,N_49203,N_49953);
nand UO_1017 (O_1017,N_47694,N_49430);
nor UO_1018 (O_1018,N_49879,N_49468);
and UO_1019 (O_1019,N_49915,N_47878);
and UO_1020 (O_1020,N_47961,N_49081);
xnor UO_1021 (O_1021,N_48415,N_49497);
xnor UO_1022 (O_1022,N_48439,N_48092);
or UO_1023 (O_1023,N_48440,N_49070);
nand UO_1024 (O_1024,N_49515,N_47845);
xnor UO_1025 (O_1025,N_49333,N_48080);
nor UO_1026 (O_1026,N_49511,N_49124);
nor UO_1027 (O_1027,N_48467,N_48145);
and UO_1028 (O_1028,N_49176,N_48463);
nand UO_1029 (O_1029,N_47830,N_47786);
xnor UO_1030 (O_1030,N_48000,N_49715);
and UO_1031 (O_1031,N_49974,N_48981);
nor UO_1032 (O_1032,N_49728,N_49632);
and UO_1033 (O_1033,N_48953,N_48722);
xor UO_1034 (O_1034,N_49993,N_49722);
nand UO_1035 (O_1035,N_47589,N_47708);
and UO_1036 (O_1036,N_48322,N_47542);
nor UO_1037 (O_1037,N_48317,N_48922);
and UO_1038 (O_1038,N_47772,N_47945);
nor UO_1039 (O_1039,N_49913,N_49592);
and UO_1040 (O_1040,N_48543,N_49968);
xor UO_1041 (O_1041,N_49653,N_49113);
nand UO_1042 (O_1042,N_47551,N_49102);
and UO_1043 (O_1043,N_49886,N_48623);
nor UO_1044 (O_1044,N_47783,N_48794);
and UO_1045 (O_1045,N_47847,N_49542);
or UO_1046 (O_1046,N_49698,N_47505);
or UO_1047 (O_1047,N_48386,N_48371);
xor UO_1048 (O_1048,N_49010,N_47774);
xor UO_1049 (O_1049,N_48741,N_47879);
nand UO_1050 (O_1050,N_49051,N_49505);
xnor UO_1051 (O_1051,N_49593,N_48552);
or UO_1052 (O_1052,N_48888,N_47686);
or UO_1053 (O_1053,N_48932,N_49050);
and UO_1054 (O_1054,N_49500,N_48615);
or UO_1055 (O_1055,N_47673,N_49726);
nand UO_1056 (O_1056,N_47893,N_48842);
nand UO_1057 (O_1057,N_49566,N_48874);
nand UO_1058 (O_1058,N_49284,N_49260);
and UO_1059 (O_1059,N_47876,N_48456);
nor UO_1060 (O_1060,N_48596,N_49252);
or UO_1061 (O_1061,N_49062,N_47645);
nor UO_1062 (O_1062,N_48435,N_47903);
nand UO_1063 (O_1063,N_48143,N_48691);
or UO_1064 (O_1064,N_49644,N_48555);
nor UO_1065 (O_1065,N_47831,N_48790);
and UO_1066 (O_1066,N_47657,N_49058);
nand UO_1067 (O_1067,N_49208,N_49955);
nor UO_1068 (O_1068,N_47809,N_47966);
nor UO_1069 (O_1069,N_47610,N_49762);
nor UO_1070 (O_1070,N_47559,N_48348);
xnor UO_1071 (O_1071,N_49031,N_49171);
and UO_1072 (O_1072,N_49939,N_48995);
and UO_1073 (O_1073,N_49601,N_47606);
and UO_1074 (O_1074,N_48003,N_49651);
xor UO_1075 (O_1075,N_49304,N_47556);
nor UO_1076 (O_1076,N_49954,N_48812);
nand UO_1077 (O_1077,N_48384,N_47836);
nor UO_1078 (O_1078,N_48563,N_48352);
xnor UO_1079 (O_1079,N_47884,N_49914);
and UO_1080 (O_1080,N_48906,N_48295);
nor UO_1081 (O_1081,N_49193,N_49317);
xor UO_1082 (O_1082,N_49271,N_48153);
nand UO_1083 (O_1083,N_48203,N_47776);
nor UO_1084 (O_1084,N_47742,N_49887);
or UO_1085 (O_1085,N_48180,N_47568);
nand UO_1086 (O_1086,N_49880,N_47975);
nand UO_1087 (O_1087,N_49099,N_49581);
xnor UO_1088 (O_1088,N_48344,N_47928);
and UO_1089 (O_1089,N_47753,N_49576);
xnor UO_1090 (O_1090,N_48349,N_48679);
xnor UO_1091 (O_1091,N_47644,N_48166);
or UO_1092 (O_1092,N_49065,N_49672);
xor UO_1093 (O_1093,N_49834,N_47900);
nand UO_1094 (O_1094,N_48478,N_49455);
nor UO_1095 (O_1095,N_47548,N_48189);
nor UO_1096 (O_1096,N_47511,N_48863);
or UO_1097 (O_1097,N_48122,N_47866);
and UO_1098 (O_1098,N_48201,N_49197);
xor UO_1099 (O_1099,N_48421,N_49646);
xnor UO_1100 (O_1100,N_47851,N_49551);
xnor UO_1101 (O_1101,N_48959,N_48118);
or UO_1102 (O_1102,N_47534,N_49224);
nor UO_1103 (O_1103,N_47732,N_48895);
xor UO_1104 (O_1104,N_48996,N_48580);
and UO_1105 (O_1105,N_48792,N_49226);
nor UO_1106 (O_1106,N_49660,N_47754);
xor UO_1107 (O_1107,N_49313,N_49342);
nor UO_1108 (O_1108,N_48670,N_48329);
nor UO_1109 (O_1109,N_48428,N_49087);
or UO_1110 (O_1110,N_49431,N_48518);
nand UO_1111 (O_1111,N_49961,N_49725);
nand UO_1112 (O_1112,N_48558,N_49662);
or UO_1113 (O_1113,N_48998,N_48010);
xnor UO_1114 (O_1114,N_49971,N_49843);
nor UO_1115 (O_1115,N_49801,N_48028);
and UO_1116 (O_1116,N_49765,N_48857);
nor UO_1117 (O_1117,N_49883,N_49240);
and UO_1118 (O_1118,N_48066,N_49459);
nand UO_1119 (O_1119,N_48314,N_49797);
nand UO_1120 (O_1120,N_48939,N_49995);
nor UO_1121 (O_1121,N_48310,N_49118);
xor UO_1122 (O_1122,N_47769,N_47950);
and UO_1123 (O_1123,N_48782,N_48069);
nand UO_1124 (O_1124,N_48761,N_49211);
or UO_1125 (O_1125,N_49851,N_48251);
and UO_1126 (O_1126,N_47693,N_49023);
and UO_1127 (O_1127,N_49479,N_48550);
nand UO_1128 (O_1128,N_48054,N_49554);
or UO_1129 (O_1129,N_47647,N_48208);
nor UO_1130 (O_1130,N_49263,N_49611);
nand UO_1131 (O_1131,N_48695,N_49991);
nand UO_1132 (O_1132,N_49767,N_48484);
xor UO_1133 (O_1133,N_48602,N_49979);
nand UO_1134 (O_1134,N_49295,N_49865);
and UO_1135 (O_1135,N_47522,N_47513);
or UO_1136 (O_1136,N_47825,N_48889);
or UO_1137 (O_1137,N_48818,N_49126);
xor UO_1138 (O_1138,N_49898,N_47870);
nand UO_1139 (O_1139,N_49630,N_49146);
or UO_1140 (O_1140,N_49407,N_48896);
and UO_1141 (O_1141,N_48183,N_48121);
xor UO_1142 (O_1142,N_49617,N_47784);
or UO_1143 (O_1143,N_47746,N_49329);
nand UO_1144 (O_1144,N_47914,N_49938);
nand UO_1145 (O_1145,N_49890,N_49978);
and UO_1146 (O_1146,N_48684,N_48406);
and UO_1147 (O_1147,N_49693,N_49792);
xor UO_1148 (O_1148,N_48268,N_49700);
or UO_1149 (O_1149,N_49351,N_47682);
or UO_1150 (O_1150,N_48991,N_48473);
or UO_1151 (O_1151,N_48103,N_49330);
or UO_1152 (O_1152,N_49071,N_48844);
and UO_1153 (O_1153,N_49292,N_49314);
or UO_1154 (O_1154,N_47788,N_47552);
nand UO_1155 (O_1155,N_49509,N_48476);
or UO_1156 (O_1156,N_49259,N_47919);
nand UO_1157 (O_1157,N_48461,N_49363);
nand UO_1158 (O_1158,N_48073,N_49169);
or UO_1159 (O_1159,N_47906,N_48833);
or UO_1160 (O_1160,N_49236,N_48805);
xnor UO_1161 (O_1161,N_49477,N_48327);
xor UO_1162 (O_1162,N_49642,N_48383);
nand UO_1163 (O_1163,N_49034,N_47887);
nor UO_1164 (O_1164,N_47911,N_47994);
nand UO_1165 (O_1165,N_48441,N_49610);
and UO_1166 (O_1166,N_47981,N_49285);
and UO_1167 (O_1167,N_49730,N_47501);
nand UO_1168 (O_1168,N_49753,N_47734);
nor UO_1169 (O_1169,N_49388,N_47762);
xnor UO_1170 (O_1170,N_49606,N_47891);
nand UO_1171 (O_1171,N_49084,N_49533);
and UO_1172 (O_1172,N_47860,N_49076);
nor UO_1173 (O_1173,N_47668,N_48447);
xor UO_1174 (O_1174,N_48315,N_47989);
or UO_1175 (O_1175,N_47944,N_48477);
nor UO_1176 (O_1176,N_48948,N_48976);
nand UO_1177 (O_1177,N_48541,N_47777);
nor UO_1178 (O_1178,N_48549,N_47770);
or UO_1179 (O_1179,N_47721,N_49457);
nand UO_1180 (O_1180,N_49972,N_47636);
nand UO_1181 (O_1181,N_49439,N_49332);
and UO_1182 (O_1182,N_49943,N_49905);
and UO_1183 (O_1183,N_47869,N_48941);
nor UO_1184 (O_1184,N_49400,N_48562);
nor UO_1185 (O_1185,N_47503,N_48688);
or UO_1186 (O_1186,N_49964,N_47920);
nor UO_1187 (O_1187,N_48119,N_49807);
or UO_1188 (O_1188,N_49229,N_48928);
and UO_1189 (O_1189,N_49008,N_48869);
nor UO_1190 (O_1190,N_49443,N_47767);
nand UO_1191 (O_1191,N_48849,N_49507);
or UO_1192 (O_1192,N_48214,N_48455);
nand UO_1193 (O_1193,N_49936,N_48226);
or UO_1194 (O_1194,N_47612,N_49916);
and UO_1195 (O_1195,N_49987,N_48285);
nor UO_1196 (O_1196,N_48865,N_48871);
and UO_1197 (O_1197,N_49907,N_48970);
nor UO_1198 (O_1198,N_48712,N_47525);
and UO_1199 (O_1199,N_48705,N_49311);
or UO_1200 (O_1200,N_47806,N_47759);
xnor UO_1201 (O_1201,N_49499,N_49981);
and UO_1202 (O_1202,N_49921,N_47865);
xor UO_1203 (O_1203,N_48452,N_49339);
or UO_1204 (O_1204,N_47558,N_49212);
nor UO_1205 (O_1205,N_47660,N_49123);
xnor UO_1206 (O_1206,N_49091,N_48256);
and UO_1207 (O_1207,N_48724,N_47661);
xor UO_1208 (O_1208,N_48770,N_48521);
and UO_1209 (O_1209,N_48417,N_49469);
nand UO_1210 (O_1210,N_49262,N_49209);
nor UO_1211 (O_1211,N_47973,N_48748);
nor UO_1212 (O_1212,N_49082,N_48594);
nand UO_1213 (O_1213,N_49221,N_48539);
or UO_1214 (O_1214,N_48341,N_48482);
xnor UO_1215 (O_1215,N_49910,N_48604);
xnor UO_1216 (O_1216,N_49931,N_47817);
xor UO_1217 (O_1217,N_48061,N_48689);
or UO_1218 (O_1218,N_48856,N_48522);
xnor UO_1219 (O_1219,N_49433,N_47592);
xnor UO_1220 (O_1220,N_49374,N_49368);
and UO_1221 (O_1221,N_48260,N_48655);
xor UO_1222 (O_1222,N_48399,N_49636);
nand UO_1223 (O_1223,N_48700,N_49364);
nor UO_1224 (O_1224,N_48750,N_49871);
nor UO_1225 (O_1225,N_47949,N_47816);
or UO_1226 (O_1226,N_49537,N_48306);
and UO_1227 (O_1227,N_49316,N_49442);
and UO_1228 (O_1228,N_48706,N_47607);
xnor UO_1229 (O_1229,N_48733,N_48458);
or UO_1230 (O_1230,N_49018,N_48861);
xor UO_1231 (O_1231,N_48347,N_49485);
xor UO_1232 (O_1232,N_47781,N_48351);
nand UO_1233 (O_1233,N_48680,N_48631);
nand UO_1234 (O_1234,N_47938,N_49876);
xnor UO_1235 (O_1235,N_48525,N_47667);
and UO_1236 (O_1236,N_48398,N_49718);
or UO_1237 (O_1237,N_48859,N_49150);
and UO_1238 (O_1238,N_49826,N_49849);
nand UO_1239 (O_1239,N_49308,N_49703);
and UO_1240 (O_1240,N_47916,N_49310);
or UO_1241 (O_1241,N_49640,N_47662);
nor UO_1242 (O_1242,N_48060,N_48988);
and UO_1243 (O_1243,N_48911,N_49288);
nor UO_1244 (O_1244,N_48943,N_48747);
nand UO_1245 (O_1245,N_47948,N_48956);
nand UO_1246 (O_1246,N_49869,N_48729);
xor UO_1247 (O_1247,N_48357,N_47600);
xor UO_1248 (O_1248,N_48848,N_48508);
or UO_1249 (O_1249,N_47867,N_49217);
nand UO_1250 (O_1250,N_49218,N_47865);
or UO_1251 (O_1251,N_49751,N_49793);
and UO_1252 (O_1252,N_49887,N_47662);
or UO_1253 (O_1253,N_49249,N_47917);
nor UO_1254 (O_1254,N_49805,N_47811);
nor UO_1255 (O_1255,N_49403,N_49526);
nand UO_1256 (O_1256,N_49389,N_47795);
nand UO_1257 (O_1257,N_48420,N_48066);
or UO_1258 (O_1258,N_49739,N_48613);
nand UO_1259 (O_1259,N_48341,N_48326);
nand UO_1260 (O_1260,N_48844,N_49935);
xnor UO_1261 (O_1261,N_49884,N_47523);
and UO_1262 (O_1262,N_48299,N_49486);
or UO_1263 (O_1263,N_48525,N_48050);
nand UO_1264 (O_1264,N_48500,N_48126);
or UO_1265 (O_1265,N_49856,N_47543);
and UO_1266 (O_1266,N_49411,N_48357);
or UO_1267 (O_1267,N_48167,N_47713);
or UO_1268 (O_1268,N_48631,N_49300);
or UO_1269 (O_1269,N_49894,N_48813);
xor UO_1270 (O_1270,N_48365,N_48384);
xor UO_1271 (O_1271,N_49945,N_47972);
nand UO_1272 (O_1272,N_47956,N_48088);
and UO_1273 (O_1273,N_49260,N_49018);
and UO_1274 (O_1274,N_49937,N_49953);
or UO_1275 (O_1275,N_48761,N_49193);
and UO_1276 (O_1276,N_48933,N_49629);
nand UO_1277 (O_1277,N_49290,N_49823);
or UO_1278 (O_1278,N_49572,N_47992);
and UO_1279 (O_1279,N_47650,N_47543);
xor UO_1280 (O_1280,N_48059,N_48036);
xor UO_1281 (O_1281,N_48898,N_48729);
nor UO_1282 (O_1282,N_47978,N_48478);
nand UO_1283 (O_1283,N_48635,N_49463);
or UO_1284 (O_1284,N_47781,N_47540);
nor UO_1285 (O_1285,N_47534,N_49727);
nor UO_1286 (O_1286,N_49481,N_48523);
or UO_1287 (O_1287,N_48474,N_48873);
and UO_1288 (O_1288,N_47916,N_49767);
or UO_1289 (O_1289,N_48986,N_48060);
nand UO_1290 (O_1290,N_49665,N_48119);
xnor UO_1291 (O_1291,N_48097,N_48558);
nand UO_1292 (O_1292,N_49609,N_49853);
nor UO_1293 (O_1293,N_48043,N_49284);
nor UO_1294 (O_1294,N_47864,N_49280);
or UO_1295 (O_1295,N_48017,N_48986);
xnor UO_1296 (O_1296,N_48427,N_48485);
nor UO_1297 (O_1297,N_48735,N_49302);
nor UO_1298 (O_1298,N_48346,N_49286);
nand UO_1299 (O_1299,N_48354,N_47710);
xor UO_1300 (O_1300,N_48483,N_49644);
or UO_1301 (O_1301,N_48263,N_47952);
or UO_1302 (O_1302,N_48833,N_48484);
nor UO_1303 (O_1303,N_47780,N_49506);
or UO_1304 (O_1304,N_48825,N_48593);
and UO_1305 (O_1305,N_48680,N_48628);
and UO_1306 (O_1306,N_49024,N_47531);
or UO_1307 (O_1307,N_48423,N_49761);
or UO_1308 (O_1308,N_49103,N_48983);
xor UO_1309 (O_1309,N_47698,N_49634);
and UO_1310 (O_1310,N_49394,N_48648);
or UO_1311 (O_1311,N_47552,N_48816);
nand UO_1312 (O_1312,N_48036,N_49623);
nor UO_1313 (O_1313,N_49268,N_49019);
or UO_1314 (O_1314,N_47891,N_48847);
nor UO_1315 (O_1315,N_47780,N_48333);
nor UO_1316 (O_1316,N_48007,N_48543);
nor UO_1317 (O_1317,N_49986,N_47500);
xnor UO_1318 (O_1318,N_47793,N_48246);
and UO_1319 (O_1319,N_49826,N_48233);
or UO_1320 (O_1320,N_48794,N_49463);
and UO_1321 (O_1321,N_48409,N_47523);
nand UO_1322 (O_1322,N_48354,N_47749);
or UO_1323 (O_1323,N_49098,N_47599);
or UO_1324 (O_1324,N_47803,N_48911);
xnor UO_1325 (O_1325,N_47822,N_49914);
nor UO_1326 (O_1326,N_49515,N_49601);
and UO_1327 (O_1327,N_48702,N_49381);
nand UO_1328 (O_1328,N_48661,N_49891);
and UO_1329 (O_1329,N_49201,N_47507);
or UO_1330 (O_1330,N_47961,N_49839);
nor UO_1331 (O_1331,N_49006,N_49916);
or UO_1332 (O_1332,N_49831,N_47545);
nor UO_1333 (O_1333,N_48458,N_47501);
or UO_1334 (O_1334,N_49489,N_49166);
xor UO_1335 (O_1335,N_48121,N_49166);
or UO_1336 (O_1336,N_48703,N_48580);
xnor UO_1337 (O_1337,N_48417,N_48896);
xor UO_1338 (O_1338,N_49034,N_48488);
or UO_1339 (O_1339,N_48764,N_49665);
or UO_1340 (O_1340,N_49413,N_49652);
and UO_1341 (O_1341,N_49900,N_48149);
and UO_1342 (O_1342,N_48427,N_49525);
or UO_1343 (O_1343,N_48756,N_49397);
nand UO_1344 (O_1344,N_48886,N_49243);
xor UO_1345 (O_1345,N_48531,N_49095);
and UO_1346 (O_1346,N_49760,N_49401);
and UO_1347 (O_1347,N_47559,N_48536);
nand UO_1348 (O_1348,N_47794,N_49111);
or UO_1349 (O_1349,N_49006,N_49720);
or UO_1350 (O_1350,N_48357,N_48408);
or UO_1351 (O_1351,N_49690,N_47672);
nor UO_1352 (O_1352,N_47801,N_48701);
xnor UO_1353 (O_1353,N_49586,N_48014);
xnor UO_1354 (O_1354,N_48969,N_48625);
nor UO_1355 (O_1355,N_49891,N_49926);
nand UO_1356 (O_1356,N_49731,N_48304);
xor UO_1357 (O_1357,N_48945,N_49673);
nor UO_1358 (O_1358,N_48415,N_49862);
nand UO_1359 (O_1359,N_48908,N_48124);
or UO_1360 (O_1360,N_49793,N_48797);
xor UO_1361 (O_1361,N_47740,N_48559);
xor UO_1362 (O_1362,N_49277,N_49278);
nor UO_1363 (O_1363,N_47868,N_49570);
or UO_1364 (O_1364,N_48919,N_49127);
xnor UO_1365 (O_1365,N_49239,N_48009);
nor UO_1366 (O_1366,N_48961,N_49748);
nand UO_1367 (O_1367,N_49367,N_48590);
or UO_1368 (O_1368,N_47584,N_48157);
or UO_1369 (O_1369,N_47854,N_49489);
and UO_1370 (O_1370,N_49371,N_48063);
nand UO_1371 (O_1371,N_49655,N_47745);
nor UO_1372 (O_1372,N_49105,N_47586);
or UO_1373 (O_1373,N_49773,N_49631);
and UO_1374 (O_1374,N_48443,N_49685);
xnor UO_1375 (O_1375,N_48727,N_48733);
or UO_1376 (O_1376,N_48818,N_49889);
and UO_1377 (O_1377,N_49124,N_48631);
and UO_1378 (O_1378,N_49792,N_49556);
or UO_1379 (O_1379,N_49712,N_48083);
xor UO_1380 (O_1380,N_49747,N_49508);
or UO_1381 (O_1381,N_47740,N_49687);
and UO_1382 (O_1382,N_49023,N_47868);
or UO_1383 (O_1383,N_49004,N_47984);
and UO_1384 (O_1384,N_48551,N_48944);
nand UO_1385 (O_1385,N_48855,N_48145);
and UO_1386 (O_1386,N_47801,N_48114);
nand UO_1387 (O_1387,N_49357,N_49178);
xnor UO_1388 (O_1388,N_48954,N_48432);
or UO_1389 (O_1389,N_48550,N_49914);
and UO_1390 (O_1390,N_49206,N_49189);
nor UO_1391 (O_1391,N_47993,N_49066);
nand UO_1392 (O_1392,N_49003,N_49019);
and UO_1393 (O_1393,N_48175,N_47786);
and UO_1394 (O_1394,N_47984,N_49924);
and UO_1395 (O_1395,N_47947,N_48722);
nor UO_1396 (O_1396,N_48273,N_47564);
nand UO_1397 (O_1397,N_47535,N_47966);
xnor UO_1398 (O_1398,N_49687,N_49024);
nor UO_1399 (O_1399,N_48235,N_49650);
and UO_1400 (O_1400,N_49376,N_49534);
or UO_1401 (O_1401,N_48624,N_49380);
and UO_1402 (O_1402,N_49521,N_47889);
and UO_1403 (O_1403,N_48842,N_49920);
nor UO_1404 (O_1404,N_47912,N_49986);
or UO_1405 (O_1405,N_48388,N_47666);
xor UO_1406 (O_1406,N_48241,N_48986);
xnor UO_1407 (O_1407,N_47511,N_48501);
or UO_1408 (O_1408,N_48970,N_48479);
and UO_1409 (O_1409,N_48282,N_48668);
and UO_1410 (O_1410,N_47764,N_48546);
nand UO_1411 (O_1411,N_49690,N_49941);
nor UO_1412 (O_1412,N_47867,N_48195);
and UO_1413 (O_1413,N_48236,N_49985);
xnor UO_1414 (O_1414,N_48984,N_48281);
xnor UO_1415 (O_1415,N_49802,N_47588);
nand UO_1416 (O_1416,N_48094,N_47974);
nand UO_1417 (O_1417,N_48970,N_48102);
or UO_1418 (O_1418,N_48037,N_49829);
nor UO_1419 (O_1419,N_49153,N_49477);
and UO_1420 (O_1420,N_48163,N_49475);
or UO_1421 (O_1421,N_48635,N_47566);
and UO_1422 (O_1422,N_47883,N_48979);
and UO_1423 (O_1423,N_47886,N_49901);
or UO_1424 (O_1424,N_49761,N_49009);
nor UO_1425 (O_1425,N_48654,N_47841);
nand UO_1426 (O_1426,N_48917,N_47744);
and UO_1427 (O_1427,N_48658,N_49027);
or UO_1428 (O_1428,N_48023,N_49168);
xnor UO_1429 (O_1429,N_48707,N_48133);
or UO_1430 (O_1430,N_47525,N_49031);
or UO_1431 (O_1431,N_49319,N_49248);
nand UO_1432 (O_1432,N_48758,N_48367);
nand UO_1433 (O_1433,N_47747,N_48433);
or UO_1434 (O_1434,N_48291,N_49861);
xor UO_1435 (O_1435,N_49711,N_48294);
and UO_1436 (O_1436,N_47665,N_48335);
nand UO_1437 (O_1437,N_49663,N_48926);
or UO_1438 (O_1438,N_49798,N_48246);
and UO_1439 (O_1439,N_48185,N_48905);
or UO_1440 (O_1440,N_48557,N_48582);
or UO_1441 (O_1441,N_49023,N_48675);
nand UO_1442 (O_1442,N_49814,N_48037);
nor UO_1443 (O_1443,N_48720,N_48781);
and UO_1444 (O_1444,N_47964,N_49803);
xnor UO_1445 (O_1445,N_49182,N_49424);
nand UO_1446 (O_1446,N_49590,N_49166);
nor UO_1447 (O_1447,N_49999,N_49522);
nand UO_1448 (O_1448,N_49273,N_48622);
and UO_1449 (O_1449,N_48061,N_49824);
and UO_1450 (O_1450,N_49443,N_48082);
or UO_1451 (O_1451,N_49530,N_49320);
nor UO_1452 (O_1452,N_48730,N_47607);
xnor UO_1453 (O_1453,N_49707,N_48006);
and UO_1454 (O_1454,N_49319,N_49002);
nand UO_1455 (O_1455,N_49800,N_48946);
nor UO_1456 (O_1456,N_47546,N_49310);
xnor UO_1457 (O_1457,N_47861,N_47900);
or UO_1458 (O_1458,N_49332,N_47965);
nor UO_1459 (O_1459,N_48784,N_48079);
nor UO_1460 (O_1460,N_49841,N_49117);
nor UO_1461 (O_1461,N_48660,N_49898);
and UO_1462 (O_1462,N_48818,N_48992);
xor UO_1463 (O_1463,N_49354,N_49660);
nor UO_1464 (O_1464,N_49317,N_47793);
and UO_1465 (O_1465,N_48465,N_48498);
and UO_1466 (O_1466,N_47920,N_49898);
nor UO_1467 (O_1467,N_49378,N_49387);
xnor UO_1468 (O_1468,N_48712,N_48884);
or UO_1469 (O_1469,N_48380,N_49674);
xnor UO_1470 (O_1470,N_49688,N_48933);
nand UO_1471 (O_1471,N_47985,N_49021);
or UO_1472 (O_1472,N_48237,N_47890);
and UO_1473 (O_1473,N_47628,N_49309);
or UO_1474 (O_1474,N_47739,N_48953);
xor UO_1475 (O_1475,N_48438,N_47891);
nor UO_1476 (O_1476,N_49422,N_47650);
and UO_1477 (O_1477,N_48293,N_47872);
xnor UO_1478 (O_1478,N_49445,N_49215);
or UO_1479 (O_1479,N_48686,N_48813);
nor UO_1480 (O_1480,N_47756,N_47752);
xor UO_1481 (O_1481,N_48712,N_49557);
or UO_1482 (O_1482,N_48548,N_48754);
xnor UO_1483 (O_1483,N_49710,N_47981);
or UO_1484 (O_1484,N_49775,N_48754);
nand UO_1485 (O_1485,N_49089,N_49254);
nor UO_1486 (O_1486,N_49791,N_48334);
or UO_1487 (O_1487,N_47639,N_48002);
nand UO_1488 (O_1488,N_49678,N_49796);
nand UO_1489 (O_1489,N_47644,N_48671);
xnor UO_1490 (O_1490,N_47523,N_49520);
nand UO_1491 (O_1491,N_49956,N_49441);
xnor UO_1492 (O_1492,N_49347,N_49499);
and UO_1493 (O_1493,N_48867,N_49078);
nand UO_1494 (O_1494,N_47930,N_47998);
and UO_1495 (O_1495,N_49880,N_49771);
or UO_1496 (O_1496,N_48311,N_48551);
and UO_1497 (O_1497,N_49344,N_47972);
xnor UO_1498 (O_1498,N_48223,N_49678);
nor UO_1499 (O_1499,N_48175,N_48192);
or UO_1500 (O_1500,N_48975,N_47920);
or UO_1501 (O_1501,N_47926,N_49619);
xnor UO_1502 (O_1502,N_48648,N_49183);
nor UO_1503 (O_1503,N_48842,N_49516);
xnor UO_1504 (O_1504,N_47681,N_49286);
nand UO_1505 (O_1505,N_48108,N_48495);
or UO_1506 (O_1506,N_47562,N_48465);
and UO_1507 (O_1507,N_48575,N_48509);
or UO_1508 (O_1508,N_48815,N_49044);
or UO_1509 (O_1509,N_48263,N_49278);
nand UO_1510 (O_1510,N_49309,N_47698);
nor UO_1511 (O_1511,N_48566,N_48021);
nand UO_1512 (O_1512,N_49470,N_47961);
nor UO_1513 (O_1513,N_48819,N_48990);
nor UO_1514 (O_1514,N_48561,N_47859);
or UO_1515 (O_1515,N_47999,N_49185);
nand UO_1516 (O_1516,N_49687,N_48232);
and UO_1517 (O_1517,N_49618,N_47732);
or UO_1518 (O_1518,N_48350,N_48076);
or UO_1519 (O_1519,N_47568,N_47958);
nor UO_1520 (O_1520,N_49321,N_47842);
nand UO_1521 (O_1521,N_49409,N_49901);
xnor UO_1522 (O_1522,N_48128,N_49322);
nor UO_1523 (O_1523,N_49959,N_49022);
or UO_1524 (O_1524,N_48110,N_49306);
or UO_1525 (O_1525,N_47854,N_49639);
xnor UO_1526 (O_1526,N_49257,N_49470);
xor UO_1527 (O_1527,N_49598,N_48112);
or UO_1528 (O_1528,N_49628,N_47942);
or UO_1529 (O_1529,N_49744,N_49486);
and UO_1530 (O_1530,N_49879,N_48197);
nand UO_1531 (O_1531,N_49866,N_47820);
nand UO_1532 (O_1532,N_49062,N_48395);
nand UO_1533 (O_1533,N_48823,N_47843);
nor UO_1534 (O_1534,N_47600,N_49321);
nand UO_1535 (O_1535,N_48251,N_48839);
and UO_1536 (O_1536,N_49986,N_48088);
nand UO_1537 (O_1537,N_49632,N_48099);
xnor UO_1538 (O_1538,N_48998,N_48462);
or UO_1539 (O_1539,N_48292,N_49412);
nand UO_1540 (O_1540,N_49469,N_48152);
nor UO_1541 (O_1541,N_48344,N_49139);
and UO_1542 (O_1542,N_49926,N_48187);
or UO_1543 (O_1543,N_48950,N_49760);
xnor UO_1544 (O_1544,N_49705,N_47585);
or UO_1545 (O_1545,N_49842,N_48097);
or UO_1546 (O_1546,N_49765,N_48283);
nand UO_1547 (O_1547,N_49781,N_48654);
xnor UO_1548 (O_1548,N_49230,N_48538);
xnor UO_1549 (O_1549,N_49358,N_49082);
and UO_1550 (O_1550,N_47782,N_49486);
nand UO_1551 (O_1551,N_48096,N_49384);
or UO_1552 (O_1552,N_49415,N_47905);
or UO_1553 (O_1553,N_49986,N_49527);
nand UO_1554 (O_1554,N_49170,N_49707);
nand UO_1555 (O_1555,N_49949,N_48195);
xor UO_1556 (O_1556,N_48447,N_48376);
or UO_1557 (O_1557,N_48313,N_49454);
xnor UO_1558 (O_1558,N_49359,N_48632);
nand UO_1559 (O_1559,N_49892,N_47937);
or UO_1560 (O_1560,N_49453,N_49502);
xor UO_1561 (O_1561,N_49388,N_48197);
xor UO_1562 (O_1562,N_48969,N_49786);
or UO_1563 (O_1563,N_47813,N_48623);
xor UO_1564 (O_1564,N_48734,N_48846);
and UO_1565 (O_1565,N_48381,N_49800);
nor UO_1566 (O_1566,N_48876,N_48836);
nor UO_1567 (O_1567,N_49311,N_49709);
xor UO_1568 (O_1568,N_49894,N_48733);
xor UO_1569 (O_1569,N_49807,N_49465);
nor UO_1570 (O_1570,N_49397,N_49196);
or UO_1571 (O_1571,N_48445,N_48852);
nor UO_1572 (O_1572,N_49023,N_48095);
and UO_1573 (O_1573,N_48120,N_48685);
nor UO_1574 (O_1574,N_48324,N_49905);
nor UO_1575 (O_1575,N_47583,N_49193);
or UO_1576 (O_1576,N_49975,N_49498);
nand UO_1577 (O_1577,N_47731,N_47682);
xor UO_1578 (O_1578,N_48637,N_48106);
nor UO_1579 (O_1579,N_48547,N_48494);
or UO_1580 (O_1580,N_49076,N_47832);
or UO_1581 (O_1581,N_48980,N_49767);
nand UO_1582 (O_1582,N_48441,N_49353);
nand UO_1583 (O_1583,N_49496,N_49416);
xnor UO_1584 (O_1584,N_49960,N_49686);
xnor UO_1585 (O_1585,N_48385,N_49201);
nor UO_1586 (O_1586,N_47938,N_49860);
xnor UO_1587 (O_1587,N_49125,N_49142);
and UO_1588 (O_1588,N_48130,N_49747);
nand UO_1589 (O_1589,N_49162,N_49243);
nand UO_1590 (O_1590,N_49148,N_48874);
nor UO_1591 (O_1591,N_47751,N_49256);
xnor UO_1592 (O_1592,N_48764,N_48043);
xor UO_1593 (O_1593,N_48731,N_48548);
nand UO_1594 (O_1594,N_48264,N_48136);
nor UO_1595 (O_1595,N_48080,N_47811);
and UO_1596 (O_1596,N_49679,N_49931);
nor UO_1597 (O_1597,N_49117,N_48178);
nor UO_1598 (O_1598,N_49324,N_48146);
nand UO_1599 (O_1599,N_49718,N_48736);
and UO_1600 (O_1600,N_49220,N_49395);
xnor UO_1601 (O_1601,N_48320,N_49757);
nor UO_1602 (O_1602,N_49813,N_47721);
nand UO_1603 (O_1603,N_48256,N_49389);
and UO_1604 (O_1604,N_47907,N_48602);
and UO_1605 (O_1605,N_49289,N_48641);
xnor UO_1606 (O_1606,N_49165,N_47522);
xor UO_1607 (O_1607,N_48438,N_47540);
or UO_1608 (O_1608,N_49709,N_49693);
xor UO_1609 (O_1609,N_48516,N_48391);
and UO_1610 (O_1610,N_49749,N_49761);
nor UO_1611 (O_1611,N_48724,N_48123);
and UO_1612 (O_1612,N_48129,N_48391);
and UO_1613 (O_1613,N_48029,N_47852);
xnor UO_1614 (O_1614,N_49058,N_49821);
and UO_1615 (O_1615,N_49415,N_48549);
nand UO_1616 (O_1616,N_49559,N_48077);
xor UO_1617 (O_1617,N_48616,N_47927);
and UO_1618 (O_1618,N_48292,N_48967);
nand UO_1619 (O_1619,N_47872,N_48453);
nand UO_1620 (O_1620,N_48855,N_48989);
and UO_1621 (O_1621,N_49945,N_48857);
nor UO_1622 (O_1622,N_48973,N_48828);
nor UO_1623 (O_1623,N_49638,N_48574);
nand UO_1624 (O_1624,N_49619,N_48555);
nor UO_1625 (O_1625,N_48014,N_49935);
nand UO_1626 (O_1626,N_48607,N_48974);
nor UO_1627 (O_1627,N_48084,N_48207);
xnor UO_1628 (O_1628,N_48455,N_47903);
nor UO_1629 (O_1629,N_49739,N_48614);
nor UO_1630 (O_1630,N_47804,N_48557);
xor UO_1631 (O_1631,N_49487,N_49233);
nor UO_1632 (O_1632,N_49663,N_48948);
or UO_1633 (O_1633,N_49653,N_48399);
nand UO_1634 (O_1634,N_48984,N_48448);
xor UO_1635 (O_1635,N_48046,N_48487);
xor UO_1636 (O_1636,N_47937,N_48201);
xnor UO_1637 (O_1637,N_49732,N_47542);
nand UO_1638 (O_1638,N_49837,N_48017);
or UO_1639 (O_1639,N_48515,N_49859);
and UO_1640 (O_1640,N_48861,N_48600);
or UO_1641 (O_1641,N_49359,N_48389);
nor UO_1642 (O_1642,N_48295,N_49423);
xor UO_1643 (O_1643,N_48400,N_47939);
and UO_1644 (O_1644,N_48772,N_47613);
or UO_1645 (O_1645,N_47945,N_49015);
nand UO_1646 (O_1646,N_49598,N_47674);
nand UO_1647 (O_1647,N_47801,N_48742);
or UO_1648 (O_1648,N_48007,N_48851);
nor UO_1649 (O_1649,N_49002,N_49231);
nand UO_1650 (O_1650,N_48097,N_48803);
and UO_1651 (O_1651,N_48902,N_47892);
nand UO_1652 (O_1652,N_48613,N_49277);
and UO_1653 (O_1653,N_48172,N_47868);
nand UO_1654 (O_1654,N_49417,N_48202);
xnor UO_1655 (O_1655,N_47604,N_49716);
and UO_1656 (O_1656,N_48155,N_49845);
xor UO_1657 (O_1657,N_48264,N_49415);
xnor UO_1658 (O_1658,N_49725,N_48891);
nand UO_1659 (O_1659,N_48170,N_48953);
nor UO_1660 (O_1660,N_49278,N_48677);
nand UO_1661 (O_1661,N_47731,N_48139);
nand UO_1662 (O_1662,N_48804,N_48523);
and UO_1663 (O_1663,N_49797,N_48192);
nand UO_1664 (O_1664,N_48004,N_47899);
and UO_1665 (O_1665,N_48094,N_48785);
xnor UO_1666 (O_1666,N_49243,N_49696);
nor UO_1667 (O_1667,N_49206,N_49080);
and UO_1668 (O_1668,N_48816,N_49225);
nand UO_1669 (O_1669,N_49084,N_47597);
and UO_1670 (O_1670,N_47525,N_49897);
nor UO_1671 (O_1671,N_47864,N_49208);
or UO_1672 (O_1672,N_47886,N_48016);
nor UO_1673 (O_1673,N_49179,N_48079);
nor UO_1674 (O_1674,N_47660,N_47978);
nor UO_1675 (O_1675,N_48870,N_49787);
xor UO_1676 (O_1676,N_47827,N_47656);
xnor UO_1677 (O_1677,N_49852,N_49432);
nor UO_1678 (O_1678,N_48847,N_49262);
nand UO_1679 (O_1679,N_47619,N_47990);
or UO_1680 (O_1680,N_48162,N_49706);
nand UO_1681 (O_1681,N_49359,N_48916);
xor UO_1682 (O_1682,N_47805,N_48224);
nor UO_1683 (O_1683,N_49257,N_48679);
and UO_1684 (O_1684,N_47727,N_48765);
or UO_1685 (O_1685,N_49161,N_48052);
nor UO_1686 (O_1686,N_47775,N_48405);
and UO_1687 (O_1687,N_49647,N_49248);
and UO_1688 (O_1688,N_49346,N_48741);
xnor UO_1689 (O_1689,N_49375,N_49805);
or UO_1690 (O_1690,N_49900,N_49060);
nand UO_1691 (O_1691,N_47772,N_49391);
or UO_1692 (O_1692,N_49235,N_47814);
nor UO_1693 (O_1693,N_48935,N_49396);
xnor UO_1694 (O_1694,N_49631,N_48047);
nor UO_1695 (O_1695,N_49007,N_47997);
nor UO_1696 (O_1696,N_48319,N_49088);
nor UO_1697 (O_1697,N_49776,N_49827);
xnor UO_1698 (O_1698,N_49549,N_49726);
xor UO_1699 (O_1699,N_49399,N_48847);
nor UO_1700 (O_1700,N_49270,N_48585);
nor UO_1701 (O_1701,N_48624,N_48547);
nand UO_1702 (O_1702,N_49825,N_49746);
or UO_1703 (O_1703,N_47891,N_48700);
xor UO_1704 (O_1704,N_48280,N_48063);
nor UO_1705 (O_1705,N_49853,N_48554);
or UO_1706 (O_1706,N_47895,N_48097);
xnor UO_1707 (O_1707,N_48771,N_49121);
xor UO_1708 (O_1708,N_49300,N_49938);
nor UO_1709 (O_1709,N_48951,N_49129);
xnor UO_1710 (O_1710,N_48801,N_48195);
xnor UO_1711 (O_1711,N_47647,N_49732);
xor UO_1712 (O_1712,N_49365,N_49198);
and UO_1713 (O_1713,N_48220,N_49146);
and UO_1714 (O_1714,N_49946,N_48498);
nand UO_1715 (O_1715,N_49430,N_47996);
nor UO_1716 (O_1716,N_48552,N_47947);
and UO_1717 (O_1717,N_49463,N_48459);
nor UO_1718 (O_1718,N_48726,N_48341);
nand UO_1719 (O_1719,N_48209,N_47749);
or UO_1720 (O_1720,N_49619,N_47725);
and UO_1721 (O_1721,N_48900,N_49894);
nor UO_1722 (O_1722,N_48107,N_47596);
xor UO_1723 (O_1723,N_49595,N_48871);
or UO_1724 (O_1724,N_47794,N_48748);
and UO_1725 (O_1725,N_49529,N_49571);
xnor UO_1726 (O_1726,N_48487,N_49009);
nor UO_1727 (O_1727,N_49739,N_48159);
and UO_1728 (O_1728,N_48324,N_49773);
and UO_1729 (O_1729,N_49488,N_48340);
xor UO_1730 (O_1730,N_47862,N_48875);
and UO_1731 (O_1731,N_48897,N_48823);
or UO_1732 (O_1732,N_48722,N_47834);
and UO_1733 (O_1733,N_49714,N_49671);
nor UO_1734 (O_1734,N_49831,N_49636);
and UO_1735 (O_1735,N_49094,N_49134);
nand UO_1736 (O_1736,N_49370,N_49385);
xnor UO_1737 (O_1737,N_49925,N_49642);
or UO_1738 (O_1738,N_48726,N_49641);
xor UO_1739 (O_1739,N_49140,N_49034);
nor UO_1740 (O_1740,N_47599,N_48673);
xor UO_1741 (O_1741,N_48584,N_48995);
xor UO_1742 (O_1742,N_48184,N_49167);
nand UO_1743 (O_1743,N_47693,N_49907);
or UO_1744 (O_1744,N_48463,N_48879);
nor UO_1745 (O_1745,N_47847,N_48610);
and UO_1746 (O_1746,N_49736,N_48716);
nand UO_1747 (O_1747,N_48383,N_48268);
nor UO_1748 (O_1748,N_47656,N_49531);
and UO_1749 (O_1749,N_49338,N_49218);
xor UO_1750 (O_1750,N_47962,N_47778);
or UO_1751 (O_1751,N_47645,N_49353);
xnor UO_1752 (O_1752,N_48653,N_47570);
xnor UO_1753 (O_1753,N_48659,N_47582);
and UO_1754 (O_1754,N_48512,N_49792);
or UO_1755 (O_1755,N_48044,N_47507);
or UO_1756 (O_1756,N_49750,N_49173);
and UO_1757 (O_1757,N_48931,N_49204);
xor UO_1758 (O_1758,N_47986,N_49482);
nand UO_1759 (O_1759,N_47981,N_48206);
xnor UO_1760 (O_1760,N_49082,N_48844);
nand UO_1761 (O_1761,N_48207,N_47564);
nand UO_1762 (O_1762,N_48731,N_47936);
xor UO_1763 (O_1763,N_49453,N_48887);
and UO_1764 (O_1764,N_49096,N_47620);
nor UO_1765 (O_1765,N_48510,N_47655);
xnor UO_1766 (O_1766,N_48264,N_47733);
nor UO_1767 (O_1767,N_49383,N_47697);
nand UO_1768 (O_1768,N_48187,N_48695);
and UO_1769 (O_1769,N_47969,N_48526);
nand UO_1770 (O_1770,N_48157,N_48346);
nand UO_1771 (O_1771,N_48714,N_49011);
or UO_1772 (O_1772,N_48425,N_47934);
and UO_1773 (O_1773,N_47652,N_49308);
or UO_1774 (O_1774,N_49904,N_48705);
nor UO_1775 (O_1775,N_49532,N_48068);
xor UO_1776 (O_1776,N_47634,N_49805);
or UO_1777 (O_1777,N_49211,N_49001);
xor UO_1778 (O_1778,N_48111,N_48719);
or UO_1779 (O_1779,N_48440,N_48591);
nor UO_1780 (O_1780,N_48059,N_49884);
xor UO_1781 (O_1781,N_47502,N_49887);
nand UO_1782 (O_1782,N_49375,N_49936);
nor UO_1783 (O_1783,N_49045,N_49774);
nand UO_1784 (O_1784,N_49715,N_48766);
or UO_1785 (O_1785,N_49486,N_48823);
and UO_1786 (O_1786,N_49588,N_49685);
xnor UO_1787 (O_1787,N_49059,N_49276);
or UO_1788 (O_1788,N_47773,N_48555);
or UO_1789 (O_1789,N_49888,N_49802);
and UO_1790 (O_1790,N_47901,N_48903);
nand UO_1791 (O_1791,N_49134,N_47875);
nor UO_1792 (O_1792,N_48575,N_48216);
nand UO_1793 (O_1793,N_47914,N_49746);
nor UO_1794 (O_1794,N_49522,N_49885);
and UO_1795 (O_1795,N_48011,N_49613);
nor UO_1796 (O_1796,N_49589,N_49270);
nor UO_1797 (O_1797,N_48369,N_48332);
nand UO_1798 (O_1798,N_49851,N_49665);
nand UO_1799 (O_1799,N_49767,N_47552);
or UO_1800 (O_1800,N_48578,N_49458);
nor UO_1801 (O_1801,N_48594,N_48276);
nor UO_1802 (O_1802,N_48438,N_48823);
or UO_1803 (O_1803,N_48904,N_48114);
and UO_1804 (O_1804,N_49824,N_49764);
nand UO_1805 (O_1805,N_47504,N_49108);
or UO_1806 (O_1806,N_47951,N_49117);
and UO_1807 (O_1807,N_48905,N_48128);
or UO_1808 (O_1808,N_49466,N_49251);
nand UO_1809 (O_1809,N_47593,N_48445);
and UO_1810 (O_1810,N_49147,N_49159);
nand UO_1811 (O_1811,N_49003,N_49450);
and UO_1812 (O_1812,N_49725,N_48798);
xnor UO_1813 (O_1813,N_49740,N_48264);
and UO_1814 (O_1814,N_48799,N_49432);
xor UO_1815 (O_1815,N_47927,N_48990);
and UO_1816 (O_1816,N_48660,N_49231);
or UO_1817 (O_1817,N_49377,N_48398);
xnor UO_1818 (O_1818,N_49384,N_49049);
xor UO_1819 (O_1819,N_47744,N_47521);
nor UO_1820 (O_1820,N_49848,N_47860);
and UO_1821 (O_1821,N_48165,N_49984);
and UO_1822 (O_1822,N_49499,N_48115);
nor UO_1823 (O_1823,N_49135,N_49070);
or UO_1824 (O_1824,N_48922,N_47671);
and UO_1825 (O_1825,N_47610,N_49013);
and UO_1826 (O_1826,N_47834,N_47543);
nor UO_1827 (O_1827,N_48599,N_49278);
and UO_1828 (O_1828,N_47788,N_49725);
or UO_1829 (O_1829,N_47827,N_49100);
nand UO_1830 (O_1830,N_48046,N_48590);
and UO_1831 (O_1831,N_49714,N_48723);
or UO_1832 (O_1832,N_48673,N_49941);
and UO_1833 (O_1833,N_48295,N_48098);
nand UO_1834 (O_1834,N_48069,N_49679);
nand UO_1835 (O_1835,N_48955,N_48153);
and UO_1836 (O_1836,N_47975,N_49546);
nand UO_1837 (O_1837,N_49614,N_48452);
nand UO_1838 (O_1838,N_49564,N_49300);
nand UO_1839 (O_1839,N_49669,N_49750);
nand UO_1840 (O_1840,N_48392,N_49316);
xor UO_1841 (O_1841,N_48048,N_48277);
nand UO_1842 (O_1842,N_48497,N_49732);
nand UO_1843 (O_1843,N_49619,N_48689);
nor UO_1844 (O_1844,N_49914,N_47744);
and UO_1845 (O_1845,N_47556,N_49442);
nand UO_1846 (O_1846,N_47690,N_49806);
xnor UO_1847 (O_1847,N_49285,N_49187);
and UO_1848 (O_1848,N_49027,N_47827);
nor UO_1849 (O_1849,N_49346,N_48255);
or UO_1850 (O_1850,N_47999,N_49769);
nor UO_1851 (O_1851,N_47813,N_49359);
or UO_1852 (O_1852,N_49735,N_49521);
and UO_1853 (O_1853,N_49747,N_48068);
nand UO_1854 (O_1854,N_48289,N_49237);
and UO_1855 (O_1855,N_48320,N_49466);
and UO_1856 (O_1856,N_47568,N_49351);
xor UO_1857 (O_1857,N_49915,N_49020);
nand UO_1858 (O_1858,N_47649,N_47889);
and UO_1859 (O_1859,N_49823,N_49119);
nor UO_1860 (O_1860,N_49386,N_48707);
xnor UO_1861 (O_1861,N_49466,N_49055);
nor UO_1862 (O_1862,N_48336,N_49404);
nand UO_1863 (O_1863,N_48636,N_49182);
and UO_1864 (O_1864,N_47646,N_48128);
nand UO_1865 (O_1865,N_47968,N_47925);
xnor UO_1866 (O_1866,N_47678,N_49478);
xor UO_1867 (O_1867,N_47527,N_48877);
or UO_1868 (O_1868,N_47706,N_49284);
xor UO_1869 (O_1869,N_49709,N_47855);
nand UO_1870 (O_1870,N_48044,N_48541);
or UO_1871 (O_1871,N_47725,N_49169);
xnor UO_1872 (O_1872,N_48629,N_48677);
xnor UO_1873 (O_1873,N_48116,N_49140);
nor UO_1874 (O_1874,N_49752,N_48996);
nand UO_1875 (O_1875,N_49643,N_48293);
or UO_1876 (O_1876,N_47757,N_49682);
and UO_1877 (O_1877,N_48696,N_48656);
xor UO_1878 (O_1878,N_49139,N_48574);
nor UO_1879 (O_1879,N_49039,N_49475);
nand UO_1880 (O_1880,N_47593,N_48830);
nand UO_1881 (O_1881,N_48116,N_47588);
xor UO_1882 (O_1882,N_47977,N_48196);
nor UO_1883 (O_1883,N_47880,N_48771);
nor UO_1884 (O_1884,N_47518,N_48016);
xnor UO_1885 (O_1885,N_49044,N_49289);
xor UO_1886 (O_1886,N_48506,N_48619);
or UO_1887 (O_1887,N_49657,N_47682);
and UO_1888 (O_1888,N_49510,N_49961);
xnor UO_1889 (O_1889,N_47988,N_48236);
xnor UO_1890 (O_1890,N_49963,N_49804);
and UO_1891 (O_1891,N_48764,N_48689);
xor UO_1892 (O_1892,N_48537,N_47825);
nor UO_1893 (O_1893,N_47734,N_48986);
xor UO_1894 (O_1894,N_49872,N_48499);
or UO_1895 (O_1895,N_49144,N_47992);
nor UO_1896 (O_1896,N_48365,N_49657);
and UO_1897 (O_1897,N_48587,N_48555);
and UO_1898 (O_1898,N_48969,N_48249);
nor UO_1899 (O_1899,N_48482,N_47952);
nor UO_1900 (O_1900,N_49135,N_48295);
or UO_1901 (O_1901,N_48514,N_48187);
or UO_1902 (O_1902,N_48623,N_47754);
and UO_1903 (O_1903,N_47889,N_48222);
and UO_1904 (O_1904,N_47766,N_49135);
nor UO_1905 (O_1905,N_47931,N_49899);
nor UO_1906 (O_1906,N_49683,N_47965);
or UO_1907 (O_1907,N_47668,N_48066);
nor UO_1908 (O_1908,N_47855,N_47521);
xor UO_1909 (O_1909,N_49163,N_48109);
xor UO_1910 (O_1910,N_48645,N_48823);
nor UO_1911 (O_1911,N_49645,N_49080);
or UO_1912 (O_1912,N_47954,N_49016);
and UO_1913 (O_1913,N_48014,N_49168);
and UO_1914 (O_1914,N_49673,N_48026);
and UO_1915 (O_1915,N_49978,N_48904);
or UO_1916 (O_1916,N_49451,N_48805);
nand UO_1917 (O_1917,N_49253,N_49958);
nand UO_1918 (O_1918,N_48188,N_47694);
nor UO_1919 (O_1919,N_49976,N_48597);
nand UO_1920 (O_1920,N_47520,N_49464);
or UO_1921 (O_1921,N_47730,N_49851);
and UO_1922 (O_1922,N_49505,N_48762);
xor UO_1923 (O_1923,N_49972,N_47887);
and UO_1924 (O_1924,N_48690,N_48198);
xor UO_1925 (O_1925,N_49937,N_49601);
nor UO_1926 (O_1926,N_48226,N_48738);
or UO_1927 (O_1927,N_47512,N_47887);
and UO_1928 (O_1928,N_47629,N_47915);
nor UO_1929 (O_1929,N_48950,N_49831);
nor UO_1930 (O_1930,N_48602,N_47959);
and UO_1931 (O_1931,N_49735,N_49195);
nor UO_1932 (O_1932,N_47502,N_49084);
or UO_1933 (O_1933,N_48470,N_48376);
or UO_1934 (O_1934,N_48030,N_49314);
nand UO_1935 (O_1935,N_49297,N_48855);
or UO_1936 (O_1936,N_49132,N_49010);
or UO_1937 (O_1937,N_48337,N_47583);
or UO_1938 (O_1938,N_48362,N_48020);
and UO_1939 (O_1939,N_49517,N_49951);
nor UO_1940 (O_1940,N_47571,N_48738);
or UO_1941 (O_1941,N_49462,N_49844);
xnor UO_1942 (O_1942,N_49856,N_49748);
nand UO_1943 (O_1943,N_49019,N_48719);
and UO_1944 (O_1944,N_48496,N_48616);
and UO_1945 (O_1945,N_47930,N_49637);
and UO_1946 (O_1946,N_48223,N_48618);
nor UO_1947 (O_1947,N_49735,N_48654);
and UO_1948 (O_1948,N_49648,N_47834);
nor UO_1949 (O_1949,N_47748,N_47816);
or UO_1950 (O_1950,N_47835,N_49877);
nand UO_1951 (O_1951,N_47781,N_49966);
or UO_1952 (O_1952,N_48033,N_48369);
xnor UO_1953 (O_1953,N_48396,N_48363);
nand UO_1954 (O_1954,N_48988,N_47588);
xnor UO_1955 (O_1955,N_48930,N_47988);
or UO_1956 (O_1956,N_47758,N_48473);
nand UO_1957 (O_1957,N_47720,N_48856);
nand UO_1958 (O_1958,N_49159,N_48314);
nor UO_1959 (O_1959,N_47772,N_49825);
nor UO_1960 (O_1960,N_48601,N_48692);
or UO_1961 (O_1961,N_49273,N_49356);
xnor UO_1962 (O_1962,N_48430,N_47905);
nor UO_1963 (O_1963,N_48417,N_47952);
xor UO_1964 (O_1964,N_48172,N_48975);
or UO_1965 (O_1965,N_47541,N_49434);
nand UO_1966 (O_1966,N_49384,N_48220);
and UO_1967 (O_1967,N_48137,N_47593);
and UO_1968 (O_1968,N_48929,N_49279);
or UO_1969 (O_1969,N_49781,N_48416);
or UO_1970 (O_1970,N_47612,N_49969);
xor UO_1971 (O_1971,N_48993,N_49880);
nor UO_1972 (O_1972,N_47952,N_49071);
nand UO_1973 (O_1973,N_48935,N_49815);
nor UO_1974 (O_1974,N_49317,N_48233);
nor UO_1975 (O_1975,N_48006,N_49469);
and UO_1976 (O_1976,N_48084,N_48066);
nand UO_1977 (O_1977,N_49858,N_49794);
xnor UO_1978 (O_1978,N_48926,N_49381);
and UO_1979 (O_1979,N_49610,N_47944);
nand UO_1980 (O_1980,N_49654,N_49875);
nand UO_1981 (O_1981,N_47784,N_48085);
nor UO_1982 (O_1982,N_49496,N_47907);
or UO_1983 (O_1983,N_47556,N_47810);
nand UO_1984 (O_1984,N_49056,N_48469);
and UO_1985 (O_1985,N_49040,N_49515);
nor UO_1986 (O_1986,N_48170,N_48240);
nand UO_1987 (O_1987,N_47960,N_49214);
nor UO_1988 (O_1988,N_48117,N_48839);
nor UO_1989 (O_1989,N_48847,N_48332);
and UO_1990 (O_1990,N_47713,N_49608);
and UO_1991 (O_1991,N_49816,N_49860);
xnor UO_1992 (O_1992,N_49464,N_48524);
or UO_1993 (O_1993,N_48866,N_49227);
and UO_1994 (O_1994,N_49858,N_48359);
or UO_1995 (O_1995,N_49235,N_47657);
and UO_1996 (O_1996,N_48147,N_49526);
and UO_1997 (O_1997,N_49788,N_49728);
xor UO_1998 (O_1998,N_48006,N_48378);
nand UO_1999 (O_1999,N_49313,N_48813);
and UO_2000 (O_2000,N_48890,N_49484);
nand UO_2001 (O_2001,N_48762,N_49242);
and UO_2002 (O_2002,N_49005,N_49009);
nor UO_2003 (O_2003,N_47965,N_49033);
and UO_2004 (O_2004,N_49050,N_47662);
and UO_2005 (O_2005,N_48286,N_48161);
or UO_2006 (O_2006,N_49800,N_48284);
nor UO_2007 (O_2007,N_48570,N_47536);
and UO_2008 (O_2008,N_48361,N_49682);
xnor UO_2009 (O_2009,N_49676,N_49036);
and UO_2010 (O_2010,N_47519,N_48908);
or UO_2011 (O_2011,N_47816,N_48651);
nand UO_2012 (O_2012,N_49521,N_48096);
nor UO_2013 (O_2013,N_48204,N_48691);
or UO_2014 (O_2014,N_48128,N_49583);
nand UO_2015 (O_2015,N_49170,N_48543);
xnor UO_2016 (O_2016,N_49485,N_49018);
nand UO_2017 (O_2017,N_48683,N_49669);
nand UO_2018 (O_2018,N_48911,N_49839);
nand UO_2019 (O_2019,N_48929,N_49588);
xor UO_2020 (O_2020,N_49767,N_47998);
or UO_2021 (O_2021,N_48007,N_48062);
nor UO_2022 (O_2022,N_49769,N_49264);
nor UO_2023 (O_2023,N_47768,N_48829);
or UO_2024 (O_2024,N_49617,N_48282);
and UO_2025 (O_2025,N_48974,N_48514);
nand UO_2026 (O_2026,N_49594,N_48249);
or UO_2027 (O_2027,N_47606,N_48443);
nor UO_2028 (O_2028,N_49197,N_48168);
nand UO_2029 (O_2029,N_47987,N_48299);
nand UO_2030 (O_2030,N_48376,N_49762);
or UO_2031 (O_2031,N_47968,N_49756);
and UO_2032 (O_2032,N_47816,N_48031);
nor UO_2033 (O_2033,N_49622,N_48634);
or UO_2034 (O_2034,N_47573,N_49941);
nor UO_2035 (O_2035,N_48812,N_49525);
xor UO_2036 (O_2036,N_48684,N_48186);
nor UO_2037 (O_2037,N_49540,N_48264);
nand UO_2038 (O_2038,N_48129,N_49589);
or UO_2039 (O_2039,N_48830,N_48148);
and UO_2040 (O_2040,N_48489,N_49009);
or UO_2041 (O_2041,N_49241,N_48842);
xnor UO_2042 (O_2042,N_48136,N_48781);
nand UO_2043 (O_2043,N_49856,N_49375);
xnor UO_2044 (O_2044,N_48289,N_49779);
xor UO_2045 (O_2045,N_49474,N_49311);
nor UO_2046 (O_2046,N_48176,N_47763);
xor UO_2047 (O_2047,N_49852,N_49039);
or UO_2048 (O_2048,N_48173,N_48261);
xor UO_2049 (O_2049,N_49975,N_48262);
nor UO_2050 (O_2050,N_48847,N_49863);
xnor UO_2051 (O_2051,N_49688,N_47504);
xnor UO_2052 (O_2052,N_49868,N_47928);
nand UO_2053 (O_2053,N_49266,N_49704);
or UO_2054 (O_2054,N_47992,N_47641);
nor UO_2055 (O_2055,N_48072,N_48078);
xor UO_2056 (O_2056,N_49411,N_49427);
or UO_2057 (O_2057,N_48451,N_49958);
or UO_2058 (O_2058,N_48859,N_49315);
nor UO_2059 (O_2059,N_49344,N_47526);
xor UO_2060 (O_2060,N_48820,N_47543);
xnor UO_2061 (O_2061,N_47718,N_48658);
nor UO_2062 (O_2062,N_48101,N_47767);
and UO_2063 (O_2063,N_48523,N_48298);
nand UO_2064 (O_2064,N_49715,N_48370);
or UO_2065 (O_2065,N_48053,N_47870);
xor UO_2066 (O_2066,N_49176,N_48916);
and UO_2067 (O_2067,N_49177,N_48566);
xnor UO_2068 (O_2068,N_48386,N_47660);
nor UO_2069 (O_2069,N_49506,N_47506);
and UO_2070 (O_2070,N_47682,N_47526);
or UO_2071 (O_2071,N_49680,N_48008);
nand UO_2072 (O_2072,N_49054,N_49531);
nor UO_2073 (O_2073,N_48189,N_48181);
or UO_2074 (O_2074,N_48357,N_47601);
and UO_2075 (O_2075,N_48927,N_49599);
xnor UO_2076 (O_2076,N_49057,N_47502);
xnor UO_2077 (O_2077,N_47823,N_47619);
or UO_2078 (O_2078,N_48591,N_47500);
or UO_2079 (O_2079,N_48589,N_48668);
nor UO_2080 (O_2080,N_48335,N_48771);
nor UO_2081 (O_2081,N_47637,N_47718);
nor UO_2082 (O_2082,N_47658,N_48016);
nor UO_2083 (O_2083,N_48137,N_48245);
nand UO_2084 (O_2084,N_47814,N_47663);
nand UO_2085 (O_2085,N_48691,N_47598);
nor UO_2086 (O_2086,N_47740,N_48308);
nand UO_2087 (O_2087,N_48709,N_48959);
xor UO_2088 (O_2088,N_47945,N_48961);
nor UO_2089 (O_2089,N_48577,N_47616);
xor UO_2090 (O_2090,N_49866,N_48350);
xor UO_2091 (O_2091,N_48731,N_49161);
or UO_2092 (O_2092,N_48567,N_49500);
nor UO_2093 (O_2093,N_48593,N_48712);
or UO_2094 (O_2094,N_49873,N_49191);
nand UO_2095 (O_2095,N_49704,N_49884);
or UO_2096 (O_2096,N_48596,N_48423);
or UO_2097 (O_2097,N_47615,N_48399);
nand UO_2098 (O_2098,N_47876,N_49775);
nor UO_2099 (O_2099,N_48918,N_48065);
or UO_2100 (O_2100,N_48322,N_48208);
or UO_2101 (O_2101,N_48589,N_48025);
nand UO_2102 (O_2102,N_48751,N_48028);
or UO_2103 (O_2103,N_48851,N_48505);
xor UO_2104 (O_2104,N_49721,N_48731);
nor UO_2105 (O_2105,N_49579,N_49871);
and UO_2106 (O_2106,N_49052,N_49041);
or UO_2107 (O_2107,N_48656,N_48626);
xor UO_2108 (O_2108,N_48328,N_48487);
nand UO_2109 (O_2109,N_48881,N_49067);
or UO_2110 (O_2110,N_48211,N_48214);
xnor UO_2111 (O_2111,N_47684,N_48603);
nand UO_2112 (O_2112,N_49745,N_49398);
xnor UO_2113 (O_2113,N_49691,N_47673);
nor UO_2114 (O_2114,N_48753,N_49410);
and UO_2115 (O_2115,N_49631,N_49371);
nand UO_2116 (O_2116,N_49329,N_48934);
xnor UO_2117 (O_2117,N_49353,N_48270);
and UO_2118 (O_2118,N_47977,N_49046);
or UO_2119 (O_2119,N_47854,N_48466);
and UO_2120 (O_2120,N_49600,N_48490);
xnor UO_2121 (O_2121,N_49592,N_49514);
nor UO_2122 (O_2122,N_48410,N_49076);
nand UO_2123 (O_2123,N_48950,N_47919);
and UO_2124 (O_2124,N_49569,N_49806);
and UO_2125 (O_2125,N_49609,N_48389);
and UO_2126 (O_2126,N_47516,N_48140);
nor UO_2127 (O_2127,N_48402,N_48529);
or UO_2128 (O_2128,N_47531,N_48140);
or UO_2129 (O_2129,N_49212,N_48738);
nor UO_2130 (O_2130,N_49384,N_48962);
and UO_2131 (O_2131,N_48417,N_49966);
or UO_2132 (O_2132,N_47736,N_49289);
nand UO_2133 (O_2133,N_49749,N_48476);
nand UO_2134 (O_2134,N_49732,N_47915);
xnor UO_2135 (O_2135,N_48940,N_47690);
xnor UO_2136 (O_2136,N_47853,N_48845);
nor UO_2137 (O_2137,N_49953,N_48292);
nor UO_2138 (O_2138,N_49350,N_48844);
xnor UO_2139 (O_2139,N_48210,N_49271);
nor UO_2140 (O_2140,N_49812,N_48223);
and UO_2141 (O_2141,N_47782,N_48355);
and UO_2142 (O_2142,N_49522,N_49410);
or UO_2143 (O_2143,N_48025,N_49287);
nand UO_2144 (O_2144,N_49076,N_49346);
nor UO_2145 (O_2145,N_49997,N_49256);
nand UO_2146 (O_2146,N_48308,N_49536);
xnor UO_2147 (O_2147,N_48038,N_47825);
and UO_2148 (O_2148,N_48463,N_48819);
or UO_2149 (O_2149,N_49295,N_48017);
and UO_2150 (O_2150,N_48949,N_48859);
and UO_2151 (O_2151,N_48723,N_49110);
and UO_2152 (O_2152,N_49355,N_48676);
and UO_2153 (O_2153,N_49619,N_47749);
xnor UO_2154 (O_2154,N_49603,N_48453);
or UO_2155 (O_2155,N_49325,N_48383);
and UO_2156 (O_2156,N_48485,N_47595);
nor UO_2157 (O_2157,N_49423,N_47854);
xor UO_2158 (O_2158,N_48308,N_48709);
xor UO_2159 (O_2159,N_48863,N_48547);
nand UO_2160 (O_2160,N_48093,N_47925);
nand UO_2161 (O_2161,N_49873,N_49842);
nor UO_2162 (O_2162,N_48288,N_48972);
or UO_2163 (O_2163,N_47522,N_48681);
and UO_2164 (O_2164,N_48013,N_49831);
nor UO_2165 (O_2165,N_49849,N_49547);
xor UO_2166 (O_2166,N_48240,N_48738);
or UO_2167 (O_2167,N_48139,N_48065);
or UO_2168 (O_2168,N_48278,N_49287);
xor UO_2169 (O_2169,N_49493,N_47967);
nor UO_2170 (O_2170,N_48486,N_49673);
nor UO_2171 (O_2171,N_48109,N_49293);
nand UO_2172 (O_2172,N_47864,N_48645);
nand UO_2173 (O_2173,N_49008,N_48401);
nand UO_2174 (O_2174,N_47713,N_48053);
xnor UO_2175 (O_2175,N_49176,N_49789);
xnor UO_2176 (O_2176,N_47667,N_49871);
xnor UO_2177 (O_2177,N_49487,N_48045);
nor UO_2178 (O_2178,N_49193,N_49422);
xnor UO_2179 (O_2179,N_48254,N_49617);
nor UO_2180 (O_2180,N_49126,N_48139);
nor UO_2181 (O_2181,N_49428,N_49490);
nor UO_2182 (O_2182,N_47717,N_49654);
nor UO_2183 (O_2183,N_49278,N_48761);
and UO_2184 (O_2184,N_49979,N_49534);
xor UO_2185 (O_2185,N_48964,N_49762);
and UO_2186 (O_2186,N_49478,N_49377);
and UO_2187 (O_2187,N_47974,N_49024);
xor UO_2188 (O_2188,N_48477,N_47651);
or UO_2189 (O_2189,N_48698,N_47987);
and UO_2190 (O_2190,N_49771,N_48888);
and UO_2191 (O_2191,N_48141,N_48771);
or UO_2192 (O_2192,N_49099,N_49531);
xnor UO_2193 (O_2193,N_48796,N_47892);
nand UO_2194 (O_2194,N_48043,N_48123);
xnor UO_2195 (O_2195,N_48689,N_49116);
nand UO_2196 (O_2196,N_47762,N_49385);
nor UO_2197 (O_2197,N_49880,N_47670);
nand UO_2198 (O_2198,N_49508,N_49568);
or UO_2199 (O_2199,N_48712,N_49252);
and UO_2200 (O_2200,N_48795,N_48599);
nand UO_2201 (O_2201,N_48436,N_48253);
or UO_2202 (O_2202,N_47664,N_47587);
xnor UO_2203 (O_2203,N_49442,N_47574);
nand UO_2204 (O_2204,N_49312,N_49410);
or UO_2205 (O_2205,N_48483,N_49833);
xnor UO_2206 (O_2206,N_47606,N_49231);
xor UO_2207 (O_2207,N_49537,N_48902);
nand UO_2208 (O_2208,N_49248,N_49330);
nor UO_2209 (O_2209,N_48542,N_47989);
nand UO_2210 (O_2210,N_49402,N_49750);
nor UO_2211 (O_2211,N_48257,N_49643);
nand UO_2212 (O_2212,N_48830,N_49364);
nand UO_2213 (O_2213,N_48076,N_48091);
nor UO_2214 (O_2214,N_47767,N_48727);
and UO_2215 (O_2215,N_48713,N_49569);
or UO_2216 (O_2216,N_49068,N_49401);
and UO_2217 (O_2217,N_47696,N_48814);
xnor UO_2218 (O_2218,N_49952,N_49696);
nor UO_2219 (O_2219,N_49644,N_49438);
nand UO_2220 (O_2220,N_48565,N_49954);
xnor UO_2221 (O_2221,N_49388,N_49743);
nor UO_2222 (O_2222,N_49795,N_49583);
or UO_2223 (O_2223,N_47649,N_48662);
and UO_2224 (O_2224,N_47931,N_48951);
and UO_2225 (O_2225,N_48268,N_48349);
nand UO_2226 (O_2226,N_48988,N_48123);
xnor UO_2227 (O_2227,N_49709,N_49350);
and UO_2228 (O_2228,N_48416,N_49762);
nor UO_2229 (O_2229,N_49366,N_49261);
or UO_2230 (O_2230,N_47771,N_49261);
nand UO_2231 (O_2231,N_49491,N_48780);
or UO_2232 (O_2232,N_48134,N_48500);
or UO_2233 (O_2233,N_48910,N_48015);
xnor UO_2234 (O_2234,N_49670,N_48202);
xor UO_2235 (O_2235,N_49326,N_47982);
xor UO_2236 (O_2236,N_49116,N_49288);
and UO_2237 (O_2237,N_48905,N_48285);
and UO_2238 (O_2238,N_47578,N_49700);
and UO_2239 (O_2239,N_48830,N_48815);
nor UO_2240 (O_2240,N_49993,N_47781);
nand UO_2241 (O_2241,N_48172,N_49437);
xor UO_2242 (O_2242,N_49801,N_49392);
nor UO_2243 (O_2243,N_48312,N_48896);
or UO_2244 (O_2244,N_48429,N_49581);
or UO_2245 (O_2245,N_47505,N_47770);
nand UO_2246 (O_2246,N_49577,N_47862);
and UO_2247 (O_2247,N_48878,N_47527);
and UO_2248 (O_2248,N_49390,N_48857);
nor UO_2249 (O_2249,N_48202,N_49885);
nor UO_2250 (O_2250,N_47652,N_48450);
or UO_2251 (O_2251,N_47892,N_48749);
and UO_2252 (O_2252,N_47842,N_48942);
nand UO_2253 (O_2253,N_47943,N_49139);
nand UO_2254 (O_2254,N_49675,N_48449);
and UO_2255 (O_2255,N_48083,N_48130);
nor UO_2256 (O_2256,N_48202,N_48587);
nor UO_2257 (O_2257,N_48658,N_48791);
nor UO_2258 (O_2258,N_49230,N_48347);
and UO_2259 (O_2259,N_49682,N_48949);
nand UO_2260 (O_2260,N_48308,N_49981);
nor UO_2261 (O_2261,N_49094,N_48354);
or UO_2262 (O_2262,N_48331,N_48953);
and UO_2263 (O_2263,N_47836,N_49150);
xnor UO_2264 (O_2264,N_48198,N_48775);
xnor UO_2265 (O_2265,N_48907,N_47536);
nand UO_2266 (O_2266,N_48503,N_48995);
xnor UO_2267 (O_2267,N_47852,N_48522);
and UO_2268 (O_2268,N_47979,N_49940);
or UO_2269 (O_2269,N_49990,N_47540);
nand UO_2270 (O_2270,N_48050,N_48171);
or UO_2271 (O_2271,N_47799,N_49001);
and UO_2272 (O_2272,N_49795,N_48216);
and UO_2273 (O_2273,N_47714,N_47973);
nand UO_2274 (O_2274,N_47940,N_49901);
and UO_2275 (O_2275,N_48389,N_48204);
nand UO_2276 (O_2276,N_47567,N_47766);
nand UO_2277 (O_2277,N_48334,N_48710);
and UO_2278 (O_2278,N_48306,N_48251);
xnor UO_2279 (O_2279,N_49288,N_49500);
nand UO_2280 (O_2280,N_49213,N_48751);
xor UO_2281 (O_2281,N_48545,N_49425);
xor UO_2282 (O_2282,N_49173,N_49866);
or UO_2283 (O_2283,N_47777,N_48629);
nor UO_2284 (O_2284,N_49116,N_48488);
and UO_2285 (O_2285,N_47840,N_47863);
nor UO_2286 (O_2286,N_48704,N_48609);
nor UO_2287 (O_2287,N_49830,N_49623);
nand UO_2288 (O_2288,N_47706,N_47794);
xor UO_2289 (O_2289,N_48155,N_47798);
nor UO_2290 (O_2290,N_49061,N_49986);
or UO_2291 (O_2291,N_49455,N_49024);
or UO_2292 (O_2292,N_47791,N_48276);
and UO_2293 (O_2293,N_48641,N_48076);
or UO_2294 (O_2294,N_49073,N_49230);
and UO_2295 (O_2295,N_48927,N_48090);
xnor UO_2296 (O_2296,N_49502,N_48157);
nor UO_2297 (O_2297,N_49521,N_49768);
and UO_2298 (O_2298,N_49554,N_47723);
and UO_2299 (O_2299,N_47807,N_47521);
or UO_2300 (O_2300,N_48788,N_48452);
or UO_2301 (O_2301,N_49279,N_49744);
nand UO_2302 (O_2302,N_49291,N_47901);
or UO_2303 (O_2303,N_47581,N_49034);
xnor UO_2304 (O_2304,N_48582,N_49759);
nor UO_2305 (O_2305,N_48320,N_48640);
and UO_2306 (O_2306,N_49437,N_48206);
or UO_2307 (O_2307,N_47743,N_49060);
nor UO_2308 (O_2308,N_48034,N_48306);
nand UO_2309 (O_2309,N_49681,N_47569);
and UO_2310 (O_2310,N_49631,N_48841);
xor UO_2311 (O_2311,N_48094,N_48510);
or UO_2312 (O_2312,N_48894,N_49709);
or UO_2313 (O_2313,N_48654,N_49068);
xor UO_2314 (O_2314,N_48617,N_47703);
or UO_2315 (O_2315,N_48205,N_47556);
or UO_2316 (O_2316,N_48742,N_48382);
nor UO_2317 (O_2317,N_47883,N_47848);
nand UO_2318 (O_2318,N_49986,N_47903);
or UO_2319 (O_2319,N_47919,N_47807);
nor UO_2320 (O_2320,N_48898,N_49149);
xor UO_2321 (O_2321,N_49396,N_48400);
nor UO_2322 (O_2322,N_49161,N_48532);
nand UO_2323 (O_2323,N_49704,N_48413);
nor UO_2324 (O_2324,N_49405,N_48721);
and UO_2325 (O_2325,N_48539,N_47916);
or UO_2326 (O_2326,N_48198,N_47949);
xor UO_2327 (O_2327,N_48206,N_47886);
xnor UO_2328 (O_2328,N_49480,N_47540);
and UO_2329 (O_2329,N_48083,N_48968);
or UO_2330 (O_2330,N_48906,N_48268);
nor UO_2331 (O_2331,N_48085,N_49292);
or UO_2332 (O_2332,N_49824,N_49453);
nand UO_2333 (O_2333,N_48816,N_49187);
nand UO_2334 (O_2334,N_49820,N_48564);
nor UO_2335 (O_2335,N_48954,N_47744);
nand UO_2336 (O_2336,N_48124,N_47822);
nor UO_2337 (O_2337,N_48440,N_47925);
nor UO_2338 (O_2338,N_49493,N_48729);
nor UO_2339 (O_2339,N_49919,N_48435);
nor UO_2340 (O_2340,N_48495,N_48042);
xnor UO_2341 (O_2341,N_49542,N_49933);
and UO_2342 (O_2342,N_48430,N_49610);
xnor UO_2343 (O_2343,N_48838,N_47856);
and UO_2344 (O_2344,N_48900,N_49445);
nand UO_2345 (O_2345,N_48679,N_49692);
nor UO_2346 (O_2346,N_48427,N_49824);
or UO_2347 (O_2347,N_48326,N_48829);
xor UO_2348 (O_2348,N_49709,N_49323);
or UO_2349 (O_2349,N_49929,N_48532);
nand UO_2350 (O_2350,N_49283,N_49499);
xnor UO_2351 (O_2351,N_47887,N_49086);
nand UO_2352 (O_2352,N_49572,N_48150);
nor UO_2353 (O_2353,N_47690,N_49407);
nand UO_2354 (O_2354,N_48696,N_49436);
nand UO_2355 (O_2355,N_47816,N_48145);
nand UO_2356 (O_2356,N_47797,N_49437);
and UO_2357 (O_2357,N_47650,N_47767);
xnor UO_2358 (O_2358,N_47837,N_47679);
xnor UO_2359 (O_2359,N_48926,N_48808);
nor UO_2360 (O_2360,N_49978,N_47563);
or UO_2361 (O_2361,N_48297,N_49088);
nor UO_2362 (O_2362,N_48859,N_48825);
xnor UO_2363 (O_2363,N_47572,N_48419);
or UO_2364 (O_2364,N_47690,N_48976);
or UO_2365 (O_2365,N_47556,N_49981);
xnor UO_2366 (O_2366,N_49355,N_48773);
xor UO_2367 (O_2367,N_48411,N_49516);
nand UO_2368 (O_2368,N_48631,N_47984);
nand UO_2369 (O_2369,N_48936,N_49059);
or UO_2370 (O_2370,N_47877,N_49561);
nand UO_2371 (O_2371,N_49143,N_49119);
nand UO_2372 (O_2372,N_48795,N_48279);
and UO_2373 (O_2373,N_47503,N_47573);
or UO_2374 (O_2374,N_48189,N_49940);
or UO_2375 (O_2375,N_49661,N_48219);
or UO_2376 (O_2376,N_47888,N_49158);
or UO_2377 (O_2377,N_49066,N_49192);
nand UO_2378 (O_2378,N_49084,N_49472);
xnor UO_2379 (O_2379,N_47975,N_48703);
nor UO_2380 (O_2380,N_47540,N_47747);
and UO_2381 (O_2381,N_49838,N_48245);
or UO_2382 (O_2382,N_48578,N_48797);
nor UO_2383 (O_2383,N_49393,N_49561);
nand UO_2384 (O_2384,N_49343,N_49446);
and UO_2385 (O_2385,N_49353,N_49009);
xor UO_2386 (O_2386,N_49588,N_47900);
and UO_2387 (O_2387,N_48104,N_49602);
xor UO_2388 (O_2388,N_49468,N_49133);
nor UO_2389 (O_2389,N_48014,N_48208);
and UO_2390 (O_2390,N_49464,N_48459);
nand UO_2391 (O_2391,N_48922,N_48555);
nor UO_2392 (O_2392,N_48424,N_49551);
and UO_2393 (O_2393,N_49340,N_48460);
or UO_2394 (O_2394,N_49670,N_48806);
or UO_2395 (O_2395,N_47938,N_49991);
nor UO_2396 (O_2396,N_47777,N_49265);
xnor UO_2397 (O_2397,N_49427,N_49287);
or UO_2398 (O_2398,N_49334,N_48085);
and UO_2399 (O_2399,N_49755,N_48796);
xor UO_2400 (O_2400,N_49367,N_48781);
and UO_2401 (O_2401,N_47573,N_49221);
xnor UO_2402 (O_2402,N_49216,N_47978);
xor UO_2403 (O_2403,N_48594,N_49076);
nand UO_2404 (O_2404,N_49494,N_49401);
nor UO_2405 (O_2405,N_48351,N_49393);
or UO_2406 (O_2406,N_47731,N_47671);
or UO_2407 (O_2407,N_48899,N_47961);
nor UO_2408 (O_2408,N_47617,N_48621);
or UO_2409 (O_2409,N_49139,N_48270);
nor UO_2410 (O_2410,N_49815,N_48127);
xor UO_2411 (O_2411,N_48911,N_47813);
xnor UO_2412 (O_2412,N_48535,N_48515);
xnor UO_2413 (O_2413,N_48823,N_49823);
nor UO_2414 (O_2414,N_49505,N_48430);
or UO_2415 (O_2415,N_48144,N_49390);
or UO_2416 (O_2416,N_48546,N_49108);
and UO_2417 (O_2417,N_49361,N_48544);
or UO_2418 (O_2418,N_48933,N_49193);
nand UO_2419 (O_2419,N_49139,N_49278);
nand UO_2420 (O_2420,N_49957,N_48778);
xor UO_2421 (O_2421,N_48319,N_48379);
nor UO_2422 (O_2422,N_47630,N_49987);
or UO_2423 (O_2423,N_47692,N_49448);
xor UO_2424 (O_2424,N_47894,N_48605);
nand UO_2425 (O_2425,N_48383,N_47606);
nand UO_2426 (O_2426,N_47924,N_48568);
and UO_2427 (O_2427,N_48378,N_48714);
xnor UO_2428 (O_2428,N_49455,N_49387);
or UO_2429 (O_2429,N_49849,N_49440);
xor UO_2430 (O_2430,N_49485,N_49227);
and UO_2431 (O_2431,N_47940,N_49557);
nand UO_2432 (O_2432,N_49967,N_47753);
nor UO_2433 (O_2433,N_47664,N_49437);
or UO_2434 (O_2434,N_49733,N_49090);
nand UO_2435 (O_2435,N_48505,N_47886);
nand UO_2436 (O_2436,N_47950,N_48274);
and UO_2437 (O_2437,N_49686,N_48694);
nor UO_2438 (O_2438,N_48762,N_47822);
xor UO_2439 (O_2439,N_47504,N_49983);
nor UO_2440 (O_2440,N_48637,N_48119);
and UO_2441 (O_2441,N_48351,N_49594);
nand UO_2442 (O_2442,N_49165,N_49507);
and UO_2443 (O_2443,N_47959,N_49564);
nor UO_2444 (O_2444,N_48438,N_49436);
and UO_2445 (O_2445,N_48169,N_49259);
and UO_2446 (O_2446,N_48370,N_49840);
nor UO_2447 (O_2447,N_48111,N_49579);
and UO_2448 (O_2448,N_48401,N_48674);
nand UO_2449 (O_2449,N_48124,N_48222);
and UO_2450 (O_2450,N_49028,N_47886);
xor UO_2451 (O_2451,N_48757,N_49830);
nand UO_2452 (O_2452,N_47955,N_49968);
nor UO_2453 (O_2453,N_48666,N_49410);
and UO_2454 (O_2454,N_49040,N_48592);
or UO_2455 (O_2455,N_49171,N_47922);
nand UO_2456 (O_2456,N_49735,N_49535);
and UO_2457 (O_2457,N_48920,N_48853);
or UO_2458 (O_2458,N_48814,N_49437);
nand UO_2459 (O_2459,N_49816,N_47764);
xnor UO_2460 (O_2460,N_48902,N_49679);
nand UO_2461 (O_2461,N_49960,N_49183);
xnor UO_2462 (O_2462,N_49053,N_48188);
nor UO_2463 (O_2463,N_47609,N_49514);
or UO_2464 (O_2464,N_48535,N_48946);
or UO_2465 (O_2465,N_48683,N_49962);
nand UO_2466 (O_2466,N_48559,N_49101);
nand UO_2467 (O_2467,N_47637,N_47764);
nor UO_2468 (O_2468,N_49607,N_49452);
nand UO_2469 (O_2469,N_49416,N_47861);
xor UO_2470 (O_2470,N_49591,N_48809);
nand UO_2471 (O_2471,N_47555,N_47865);
or UO_2472 (O_2472,N_48973,N_49833);
nand UO_2473 (O_2473,N_49368,N_49253);
or UO_2474 (O_2474,N_48725,N_48371);
xnor UO_2475 (O_2475,N_48193,N_47613);
xor UO_2476 (O_2476,N_48837,N_48797);
or UO_2477 (O_2477,N_47731,N_49505);
and UO_2478 (O_2478,N_48448,N_49493);
or UO_2479 (O_2479,N_48875,N_49629);
nor UO_2480 (O_2480,N_47581,N_49636);
xor UO_2481 (O_2481,N_48928,N_48429);
xnor UO_2482 (O_2482,N_47592,N_49657);
and UO_2483 (O_2483,N_49825,N_48446);
or UO_2484 (O_2484,N_47750,N_47685);
and UO_2485 (O_2485,N_47959,N_48052);
or UO_2486 (O_2486,N_49683,N_47969);
and UO_2487 (O_2487,N_47621,N_48876);
nor UO_2488 (O_2488,N_49856,N_48372);
nand UO_2489 (O_2489,N_48885,N_49639);
xnor UO_2490 (O_2490,N_48418,N_48832);
nand UO_2491 (O_2491,N_49520,N_48118);
or UO_2492 (O_2492,N_47939,N_48477);
and UO_2493 (O_2493,N_47639,N_49830);
xnor UO_2494 (O_2494,N_49474,N_48119);
xnor UO_2495 (O_2495,N_48601,N_49354);
xnor UO_2496 (O_2496,N_49085,N_48175);
or UO_2497 (O_2497,N_49384,N_49997);
and UO_2498 (O_2498,N_47577,N_47592);
and UO_2499 (O_2499,N_49271,N_48788);
or UO_2500 (O_2500,N_48760,N_48989);
and UO_2501 (O_2501,N_48237,N_48899);
and UO_2502 (O_2502,N_48188,N_49410);
nand UO_2503 (O_2503,N_48445,N_47626);
xnor UO_2504 (O_2504,N_49924,N_47709);
nor UO_2505 (O_2505,N_48178,N_48451);
nand UO_2506 (O_2506,N_49503,N_47900);
nor UO_2507 (O_2507,N_49578,N_48836);
or UO_2508 (O_2508,N_47821,N_49641);
and UO_2509 (O_2509,N_48281,N_49125);
and UO_2510 (O_2510,N_47755,N_49964);
nor UO_2511 (O_2511,N_47542,N_47766);
nand UO_2512 (O_2512,N_48777,N_49593);
xnor UO_2513 (O_2513,N_48592,N_49101);
or UO_2514 (O_2514,N_48879,N_49369);
or UO_2515 (O_2515,N_48524,N_48776);
or UO_2516 (O_2516,N_49630,N_48700);
and UO_2517 (O_2517,N_49116,N_48984);
and UO_2518 (O_2518,N_49251,N_48522);
xor UO_2519 (O_2519,N_47681,N_48982);
nor UO_2520 (O_2520,N_48960,N_47900);
nand UO_2521 (O_2521,N_48014,N_47864);
and UO_2522 (O_2522,N_48457,N_49354);
nor UO_2523 (O_2523,N_49472,N_49962);
nand UO_2524 (O_2524,N_49566,N_47849);
or UO_2525 (O_2525,N_48284,N_49797);
or UO_2526 (O_2526,N_48924,N_49308);
nor UO_2527 (O_2527,N_47867,N_48777);
nand UO_2528 (O_2528,N_48384,N_48915);
and UO_2529 (O_2529,N_49341,N_48726);
and UO_2530 (O_2530,N_49186,N_48820);
nand UO_2531 (O_2531,N_47710,N_47502);
nor UO_2532 (O_2532,N_49467,N_48286);
and UO_2533 (O_2533,N_48619,N_48051);
and UO_2534 (O_2534,N_49380,N_47524);
nand UO_2535 (O_2535,N_48498,N_48279);
and UO_2536 (O_2536,N_48674,N_47618);
nor UO_2537 (O_2537,N_48672,N_48682);
and UO_2538 (O_2538,N_48740,N_47868);
nor UO_2539 (O_2539,N_47614,N_48686);
and UO_2540 (O_2540,N_48079,N_48912);
nand UO_2541 (O_2541,N_49180,N_48382);
xor UO_2542 (O_2542,N_48690,N_49331);
or UO_2543 (O_2543,N_49976,N_49921);
xor UO_2544 (O_2544,N_48420,N_47547);
nand UO_2545 (O_2545,N_48013,N_49760);
nand UO_2546 (O_2546,N_47827,N_48604);
nor UO_2547 (O_2547,N_48468,N_47857);
and UO_2548 (O_2548,N_49056,N_49982);
or UO_2549 (O_2549,N_49612,N_49383);
or UO_2550 (O_2550,N_49566,N_47754);
or UO_2551 (O_2551,N_49696,N_49310);
and UO_2552 (O_2552,N_47552,N_48484);
nand UO_2553 (O_2553,N_48762,N_49167);
xor UO_2554 (O_2554,N_47683,N_47586);
nor UO_2555 (O_2555,N_49939,N_48041);
and UO_2556 (O_2556,N_49207,N_47549);
or UO_2557 (O_2557,N_49889,N_49929);
nand UO_2558 (O_2558,N_47855,N_49048);
xnor UO_2559 (O_2559,N_48815,N_49917);
nor UO_2560 (O_2560,N_48731,N_49666);
and UO_2561 (O_2561,N_49377,N_48649);
nand UO_2562 (O_2562,N_47618,N_49229);
xor UO_2563 (O_2563,N_49549,N_48699);
nor UO_2564 (O_2564,N_48532,N_49711);
or UO_2565 (O_2565,N_49759,N_49122);
nand UO_2566 (O_2566,N_48075,N_48524);
xnor UO_2567 (O_2567,N_48938,N_48466);
nor UO_2568 (O_2568,N_47556,N_48467);
xnor UO_2569 (O_2569,N_49979,N_48402);
or UO_2570 (O_2570,N_49935,N_49856);
nor UO_2571 (O_2571,N_49191,N_47770);
or UO_2572 (O_2572,N_48641,N_49063);
and UO_2573 (O_2573,N_49037,N_49142);
nand UO_2574 (O_2574,N_47768,N_48208);
xor UO_2575 (O_2575,N_48580,N_48257);
nor UO_2576 (O_2576,N_48045,N_49286);
nor UO_2577 (O_2577,N_49248,N_48466);
or UO_2578 (O_2578,N_48553,N_49630);
xor UO_2579 (O_2579,N_47891,N_47673);
or UO_2580 (O_2580,N_49357,N_49583);
xnor UO_2581 (O_2581,N_49080,N_49263);
and UO_2582 (O_2582,N_49828,N_48769);
nand UO_2583 (O_2583,N_48291,N_47622);
or UO_2584 (O_2584,N_47822,N_48472);
or UO_2585 (O_2585,N_49197,N_48205);
nor UO_2586 (O_2586,N_49101,N_48064);
nor UO_2587 (O_2587,N_48128,N_47664);
nand UO_2588 (O_2588,N_47730,N_48855);
xor UO_2589 (O_2589,N_48364,N_49628);
or UO_2590 (O_2590,N_47667,N_48588);
xnor UO_2591 (O_2591,N_49861,N_48968);
or UO_2592 (O_2592,N_48502,N_48260);
nor UO_2593 (O_2593,N_48476,N_49056);
nand UO_2594 (O_2594,N_47598,N_48993);
and UO_2595 (O_2595,N_47587,N_49303);
xnor UO_2596 (O_2596,N_48118,N_48465);
or UO_2597 (O_2597,N_47598,N_48970);
nand UO_2598 (O_2598,N_47555,N_48174);
or UO_2599 (O_2599,N_48156,N_49980);
or UO_2600 (O_2600,N_48362,N_49323);
or UO_2601 (O_2601,N_47715,N_49191);
nand UO_2602 (O_2602,N_48747,N_48366);
xnor UO_2603 (O_2603,N_49243,N_47588);
nand UO_2604 (O_2604,N_48196,N_48969);
and UO_2605 (O_2605,N_47951,N_48634);
and UO_2606 (O_2606,N_48150,N_49697);
and UO_2607 (O_2607,N_49044,N_49669);
or UO_2608 (O_2608,N_49874,N_49706);
nor UO_2609 (O_2609,N_49595,N_49044);
nand UO_2610 (O_2610,N_48312,N_48685);
nor UO_2611 (O_2611,N_49422,N_48178);
xnor UO_2612 (O_2612,N_47960,N_48192);
nand UO_2613 (O_2613,N_47699,N_47523);
nand UO_2614 (O_2614,N_49435,N_49305);
and UO_2615 (O_2615,N_49521,N_48918);
nor UO_2616 (O_2616,N_48344,N_48240);
or UO_2617 (O_2617,N_48321,N_49577);
nand UO_2618 (O_2618,N_48699,N_48266);
nor UO_2619 (O_2619,N_47577,N_47665);
or UO_2620 (O_2620,N_48228,N_49649);
xor UO_2621 (O_2621,N_47574,N_48911);
xnor UO_2622 (O_2622,N_48980,N_49476);
and UO_2623 (O_2623,N_48569,N_47852);
nand UO_2624 (O_2624,N_48151,N_48571);
nand UO_2625 (O_2625,N_49466,N_49071);
xor UO_2626 (O_2626,N_48895,N_49375);
xnor UO_2627 (O_2627,N_48346,N_49572);
xnor UO_2628 (O_2628,N_47524,N_48687);
xnor UO_2629 (O_2629,N_48679,N_48356);
or UO_2630 (O_2630,N_47771,N_48852);
and UO_2631 (O_2631,N_48916,N_48084);
nand UO_2632 (O_2632,N_47761,N_48607);
and UO_2633 (O_2633,N_49304,N_48937);
or UO_2634 (O_2634,N_48979,N_48644);
nand UO_2635 (O_2635,N_47960,N_49896);
nor UO_2636 (O_2636,N_48348,N_49545);
or UO_2637 (O_2637,N_49256,N_48378);
nand UO_2638 (O_2638,N_48529,N_47896);
nand UO_2639 (O_2639,N_47912,N_48272);
nand UO_2640 (O_2640,N_47745,N_49054);
and UO_2641 (O_2641,N_49785,N_48402);
xor UO_2642 (O_2642,N_48307,N_48542);
xor UO_2643 (O_2643,N_48815,N_47878);
and UO_2644 (O_2644,N_48961,N_49056);
and UO_2645 (O_2645,N_48225,N_48571);
or UO_2646 (O_2646,N_49482,N_47780);
nand UO_2647 (O_2647,N_47535,N_48201);
nor UO_2648 (O_2648,N_48757,N_49737);
xor UO_2649 (O_2649,N_48931,N_47998);
and UO_2650 (O_2650,N_49787,N_48248);
nor UO_2651 (O_2651,N_48310,N_48162);
nand UO_2652 (O_2652,N_49489,N_49160);
xnor UO_2653 (O_2653,N_47771,N_49185);
nor UO_2654 (O_2654,N_48983,N_49267);
nor UO_2655 (O_2655,N_49088,N_49157);
nor UO_2656 (O_2656,N_49452,N_48787);
or UO_2657 (O_2657,N_48140,N_47836);
and UO_2658 (O_2658,N_48386,N_49683);
nand UO_2659 (O_2659,N_49202,N_48563);
or UO_2660 (O_2660,N_47620,N_48049);
nor UO_2661 (O_2661,N_49023,N_48563);
and UO_2662 (O_2662,N_48549,N_48675);
nor UO_2663 (O_2663,N_49091,N_49018);
nor UO_2664 (O_2664,N_49828,N_48535);
or UO_2665 (O_2665,N_47799,N_47956);
and UO_2666 (O_2666,N_48088,N_49590);
or UO_2667 (O_2667,N_49157,N_47692);
or UO_2668 (O_2668,N_48485,N_47939);
and UO_2669 (O_2669,N_49755,N_48165);
xor UO_2670 (O_2670,N_48145,N_48291);
and UO_2671 (O_2671,N_47792,N_47689);
and UO_2672 (O_2672,N_48249,N_48197);
nor UO_2673 (O_2673,N_47836,N_49697);
nand UO_2674 (O_2674,N_49815,N_48378);
and UO_2675 (O_2675,N_48521,N_49526);
nand UO_2676 (O_2676,N_48316,N_49199);
or UO_2677 (O_2677,N_47591,N_48212);
and UO_2678 (O_2678,N_49195,N_49107);
nor UO_2679 (O_2679,N_49442,N_48651);
nand UO_2680 (O_2680,N_47680,N_47530);
or UO_2681 (O_2681,N_49762,N_48215);
and UO_2682 (O_2682,N_49344,N_48120);
and UO_2683 (O_2683,N_49287,N_49677);
xor UO_2684 (O_2684,N_48433,N_48906);
and UO_2685 (O_2685,N_48504,N_49244);
and UO_2686 (O_2686,N_49584,N_48483);
or UO_2687 (O_2687,N_48823,N_49960);
nor UO_2688 (O_2688,N_49841,N_49474);
xor UO_2689 (O_2689,N_48931,N_48794);
xnor UO_2690 (O_2690,N_47977,N_47985);
nand UO_2691 (O_2691,N_48544,N_49760);
and UO_2692 (O_2692,N_48143,N_48811);
nor UO_2693 (O_2693,N_49072,N_48196);
or UO_2694 (O_2694,N_49458,N_48061);
xnor UO_2695 (O_2695,N_48227,N_49400);
nand UO_2696 (O_2696,N_47672,N_48375);
or UO_2697 (O_2697,N_49579,N_49629);
and UO_2698 (O_2698,N_49218,N_49204);
xor UO_2699 (O_2699,N_47988,N_48845);
nand UO_2700 (O_2700,N_47715,N_48708);
xnor UO_2701 (O_2701,N_48410,N_49629);
nand UO_2702 (O_2702,N_48022,N_47777);
nor UO_2703 (O_2703,N_48237,N_48574);
xnor UO_2704 (O_2704,N_47696,N_49589);
nand UO_2705 (O_2705,N_48253,N_49789);
and UO_2706 (O_2706,N_49340,N_49169);
or UO_2707 (O_2707,N_49550,N_47949);
or UO_2708 (O_2708,N_48792,N_47670);
nand UO_2709 (O_2709,N_48138,N_48937);
and UO_2710 (O_2710,N_48190,N_48750);
nand UO_2711 (O_2711,N_47647,N_49766);
nand UO_2712 (O_2712,N_49163,N_49932);
xor UO_2713 (O_2713,N_48127,N_47836);
nand UO_2714 (O_2714,N_49299,N_49668);
nand UO_2715 (O_2715,N_49606,N_48323);
nor UO_2716 (O_2716,N_47981,N_48301);
nand UO_2717 (O_2717,N_49299,N_49450);
or UO_2718 (O_2718,N_48956,N_48763);
nor UO_2719 (O_2719,N_49465,N_48906);
xor UO_2720 (O_2720,N_47931,N_48883);
nor UO_2721 (O_2721,N_48346,N_47751);
xnor UO_2722 (O_2722,N_48996,N_48353);
and UO_2723 (O_2723,N_48244,N_47642);
nor UO_2724 (O_2724,N_49811,N_49674);
or UO_2725 (O_2725,N_49635,N_48224);
and UO_2726 (O_2726,N_49777,N_48349);
nand UO_2727 (O_2727,N_49051,N_49584);
or UO_2728 (O_2728,N_49351,N_48394);
or UO_2729 (O_2729,N_48890,N_48771);
xor UO_2730 (O_2730,N_48714,N_48669);
or UO_2731 (O_2731,N_48058,N_49654);
nand UO_2732 (O_2732,N_49548,N_48609);
nand UO_2733 (O_2733,N_48203,N_47673);
xor UO_2734 (O_2734,N_47604,N_49072);
nand UO_2735 (O_2735,N_48868,N_49606);
nand UO_2736 (O_2736,N_49801,N_49219);
nand UO_2737 (O_2737,N_48049,N_49261);
nand UO_2738 (O_2738,N_48787,N_49633);
xnor UO_2739 (O_2739,N_47538,N_49480);
nand UO_2740 (O_2740,N_48846,N_49063);
nand UO_2741 (O_2741,N_49915,N_49301);
or UO_2742 (O_2742,N_48036,N_48322);
xor UO_2743 (O_2743,N_49993,N_49216);
and UO_2744 (O_2744,N_47937,N_48169);
or UO_2745 (O_2745,N_49334,N_48485);
nor UO_2746 (O_2746,N_49473,N_48507);
nor UO_2747 (O_2747,N_47916,N_47522);
xor UO_2748 (O_2748,N_48687,N_48792);
xnor UO_2749 (O_2749,N_47625,N_48022);
nor UO_2750 (O_2750,N_49504,N_47844);
nor UO_2751 (O_2751,N_47791,N_48518);
xnor UO_2752 (O_2752,N_49994,N_49954);
or UO_2753 (O_2753,N_48487,N_48287);
xor UO_2754 (O_2754,N_48805,N_49527);
nand UO_2755 (O_2755,N_49629,N_49921);
or UO_2756 (O_2756,N_48751,N_48969);
nor UO_2757 (O_2757,N_48981,N_48673);
and UO_2758 (O_2758,N_49753,N_49137);
or UO_2759 (O_2759,N_49382,N_47598);
nand UO_2760 (O_2760,N_47529,N_49174);
nor UO_2761 (O_2761,N_49145,N_47917);
xnor UO_2762 (O_2762,N_48037,N_49356);
xor UO_2763 (O_2763,N_49301,N_48087);
nand UO_2764 (O_2764,N_49571,N_48924);
nand UO_2765 (O_2765,N_47845,N_48967);
xor UO_2766 (O_2766,N_49539,N_48669);
xor UO_2767 (O_2767,N_47612,N_47876);
xor UO_2768 (O_2768,N_49374,N_49670);
and UO_2769 (O_2769,N_47846,N_49199);
or UO_2770 (O_2770,N_48372,N_49566);
nor UO_2771 (O_2771,N_49615,N_49518);
nor UO_2772 (O_2772,N_47985,N_47627);
nand UO_2773 (O_2773,N_48426,N_48280);
and UO_2774 (O_2774,N_49476,N_49916);
xnor UO_2775 (O_2775,N_48555,N_49274);
or UO_2776 (O_2776,N_48485,N_48814);
and UO_2777 (O_2777,N_48082,N_48576);
and UO_2778 (O_2778,N_49174,N_47634);
nor UO_2779 (O_2779,N_48344,N_49142);
xnor UO_2780 (O_2780,N_49593,N_47728);
and UO_2781 (O_2781,N_47755,N_49992);
xor UO_2782 (O_2782,N_47693,N_48635);
nor UO_2783 (O_2783,N_49435,N_47853);
nor UO_2784 (O_2784,N_49311,N_49641);
nand UO_2785 (O_2785,N_49576,N_49697);
or UO_2786 (O_2786,N_49560,N_48649);
and UO_2787 (O_2787,N_49994,N_49951);
or UO_2788 (O_2788,N_48129,N_47684);
xnor UO_2789 (O_2789,N_47528,N_48888);
or UO_2790 (O_2790,N_48657,N_48803);
xor UO_2791 (O_2791,N_49106,N_48826);
xnor UO_2792 (O_2792,N_49593,N_49054);
or UO_2793 (O_2793,N_48879,N_48581);
or UO_2794 (O_2794,N_48712,N_47867);
nand UO_2795 (O_2795,N_49280,N_48586);
and UO_2796 (O_2796,N_47982,N_48168);
or UO_2797 (O_2797,N_48955,N_47565);
nand UO_2798 (O_2798,N_48931,N_49451);
or UO_2799 (O_2799,N_48858,N_49323);
and UO_2800 (O_2800,N_47734,N_49372);
xnor UO_2801 (O_2801,N_49342,N_48202);
or UO_2802 (O_2802,N_49708,N_49257);
or UO_2803 (O_2803,N_49683,N_48750);
nor UO_2804 (O_2804,N_49782,N_47699);
nor UO_2805 (O_2805,N_49679,N_48357);
nand UO_2806 (O_2806,N_48798,N_49446);
or UO_2807 (O_2807,N_49289,N_48415);
or UO_2808 (O_2808,N_49972,N_47721);
nand UO_2809 (O_2809,N_49662,N_48673);
nor UO_2810 (O_2810,N_49715,N_49893);
xnor UO_2811 (O_2811,N_48380,N_48675);
or UO_2812 (O_2812,N_48442,N_47906);
xnor UO_2813 (O_2813,N_49725,N_49682);
and UO_2814 (O_2814,N_48659,N_49214);
nand UO_2815 (O_2815,N_48120,N_48361);
and UO_2816 (O_2816,N_48178,N_49147);
and UO_2817 (O_2817,N_49860,N_48885);
nor UO_2818 (O_2818,N_47669,N_48193);
nand UO_2819 (O_2819,N_49661,N_49214);
and UO_2820 (O_2820,N_47717,N_48773);
nor UO_2821 (O_2821,N_49451,N_49905);
and UO_2822 (O_2822,N_47880,N_49013);
nand UO_2823 (O_2823,N_49022,N_47773);
nor UO_2824 (O_2824,N_48010,N_48310);
xor UO_2825 (O_2825,N_48738,N_49143);
nand UO_2826 (O_2826,N_49883,N_49663);
or UO_2827 (O_2827,N_49140,N_48940);
xnor UO_2828 (O_2828,N_49705,N_48058);
or UO_2829 (O_2829,N_47795,N_48723);
xnor UO_2830 (O_2830,N_49126,N_49283);
nand UO_2831 (O_2831,N_49275,N_49436);
xnor UO_2832 (O_2832,N_48027,N_48257);
xnor UO_2833 (O_2833,N_48288,N_48578);
nor UO_2834 (O_2834,N_49396,N_48530);
and UO_2835 (O_2835,N_48326,N_48062);
or UO_2836 (O_2836,N_48651,N_49119);
or UO_2837 (O_2837,N_49276,N_49553);
and UO_2838 (O_2838,N_48459,N_47747);
nand UO_2839 (O_2839,N_48765,N_49790);
and UO_2840 (O_2840,N_49366,N_48581);
nand UO_2841 (O_2841,N_48848,N_48902);
and UO_2842 (O_2842,N_48415,N_47698);
and UO_2843 (O_2843,N_48119,N_48535);
xor UO_2844 (O_2844,N_47990,N_48713);
or UO_2845 (O_2845,N_48348,N_48258);
nand UO_2846 (O_2846,N_49462,N_49516);
nand UO_2847 (O_2847,N_49527,N_48308);
or UO_2848 (O_2848,N_48474,N_48175);
nand UO_2849 (O_2849,N_48077,N_49956);
and UO_2850 (O_2850,N_49983,N_49869);
nand UO_2851 (O_2851,N_48875,N_47638);
nand UO_2852 (O_2852,N_49653,N_48920);
xnor UO_2853 (O_2853,N_49463,N_48478);
nand UO_2854 (O_2854,N_47571,N_47531);
xor UO_2855 (O_2855,N_49329,N_47520);
or UO_2856 (O_2856,N_48047,N_49067);
nor UO_2857 (O_2857,N_49777,N_49705);
xor UO_2858 (O_2858,N_48844,N_49484);
xor UO_2859 (O_2859,N_48780,N_48525);
or UO_2860 (O_2860,N_49583,N_49809);
or UO_2861 (O_2861,N_48343,N_49806);
and UO_2862 (O_2862,N_47965,N_48664);
nand UO_2863 (O_2863,N_49998,N_48995);
xor UO_2864 (O_2864,N_48002,N_49318);
or UO_2865 (O_2865,N_48742,N_48672);
and UO_2866 (O_2866,N_49314,N_49819);
nand UO_2867 (O_2867,N_48099,N_48327);
or UO_2868 (O_2868,N_47651,N_47713);
or UO_2869 (O_2869,N_49218,N_48075);
xnor UO_2870 (O_2870,N_47608,N_47834);
xnor UO_2871 (O_2871,N_48783,N_49131);
xor UO_2872 (O_2872,N_49660,N_49109);
nor UO_2873 (O_2873,N_47803,N_49291);
nor UO_2874 (O_2874,N_49122,N_47584);
or UO_2875 (O_2875,N_47630,N_48263);
and UO_2876 (O_2876,N_49447,N_48762);
or UO_2877 (O_2877,N_48099,N_47927);
nand UO_2878 (O_2878,N_47897,N_49010);
nand UO_2879 (O_2879,N_47573,N_48396);
nor UO_2880 (O_2880,N_49015,N_48220);
xnor UO_2881 (O_2881,N_48261,N_49856);
and UO_2882 (O_2882,N_48298,N_49620);
nand UO_2883 (O_2883,N_49255,N_47864);
nor UO_2884 (O_2884,N_48916,N_49161);
xor UO_2885 (O_2885,N_49644,N_48724);
nand UO_2886 (O_2886,N_47918,N_47510);
and UO_2887 (O_2887,N_49894,N_49063);
nand UO_2888 (O_2888,N_48846,N_49909);
nor UO_2889 (O_2889,N_49360,N_49663);
nor UO_2890 (O_2890,N_48769,N_49771);
nand UO_2891 (O_2891,N_48144,N_49927);
xor UO_2892 (O_2892,N_48558,N_49656);
nand UO_2893 (O_2893,N_47861,N_49625);
or UO_2894 (O_2894,N_47531,N_48046);
or UO_2895 (O_2895,N_47797,N_49233);
and UO_2896 (O_2896,N_49129,N_49144);
xnor UO_2897 (O_2897,N_47879,N_49634);
xnor UO_2898 (O_2898,N_47879,N_49446);
xnor UO_2899 (O_2899,N_47801,N_48898);
nand UO_2900 (O_2900,N_47813,N_49373);
xor UO_2901 (O_2901,N_48361,N_49102);
or UO_2902 (O_2902,N_48140,N_47744);
nor UO_2903 (O_2903,N_47770,N_49087);
nand UO_2904 (O_2904,N_49710,N_47930);
or UO_2905 (O_2905,N_47545,N_48004);
nand UO_2906 (O_2906,N_49049,N_48251);
nor UO_2907 (O_2907,N_48229,N_47543);
or UO_2908 (O_2908,N_49810,N_48945);
or UO_2909 (O_2909,N_48083,N_49379);
xor UO_2910 (O_2910,N_49616,N_48608);
and UO_2911 (O_2911,N_48056,N_48135);
and UO_2912 (O_2912,N_49942,N_47970);
nand UO_2913 (O_2913,N_49883,N_48039);
and UO_2914 (O_2914,N_47721,N_47648);
and UO_2915 (O_2915,N_49393,N_48979);
nand UO_2916 (O_2916,N_49124,N_49735);
or UO_2917 (O_2917,N_47844,N_48028);
or UO_2918 (O_2918,N_48295,N_47510);
xnor UO_2919 (O_2919,N_49887,N_49540);
and UO_2920 (O_2920,N_49529,N_49376);
nor UO_2921 (O_2921,N_48765,N_49001);
xor UO_2922 (O_2922,N_48470,N_48757);
or UO_2923 (O_2923,N_47604,N_48192);
nand UO_2924 (O_2924,N_49251,N_49913);
nand UO_2925 (O_2925,N_48682,N_48694);
xnor UO_2926 (O_2926,N_47974,N_49226);
nor UO_2927 (O_2927,N_48986,N_49071);
and UO_2928 (O_2928,N_48402,N_48757);
nor UO_2929 (O_2929,N_48318,N_49905);
nand UO_2930 (O_2930,N_49942,N_48957);
nand UO_2931 (O_2931,N_48435,N_48322);
xnor UO_2932 (O_2932,N_49303,N_49778);
nor UO_2933 (O_2933,N_49480,N_49244);
and UO_2934 (O_2934,N_47730,N_49645);
xor UO_2935 (O_2935,N_48255,N_48443);
and UO_2936 (O_2936,N_48765,N_49524);
nor UO_2937 (O_2937,N_48715,N_48570);
nor UO_2938 (O_2938,N_49689,N_48195);
or UO_2939 (O_2939,N_48392,N_49639);
nand UO_2940 (O_2940,N_49834,N_47743);
and UO_2941 (O_2941,N_49132,N_49004);
xor UO_2942 (O_2942,N_49763,N_49260);
xor UO_2943 (O_2943,N_48096,N_48446);
or UO_2944 (O_2944,N_49952,N_48762);
nor UO_2945 (O_2945,N_47878,N_48269);
and UO_2946 (O_2946,N_47861,N_47684);
nand UO_2947 (O_2947,N_49967,N_49858);
nor UO_2948 (O_2948,N_47880,N_49678);
or UO_2949 (O_2949,N_48302,N_48714);
nand UO_2950 (O_2950,N_49526,N_48844);
nand UO_2951 (O_2951,N_48689,N_49383);
nand UO_2952 (O_2952,N_47732,N_47904);
xnor UO_2953 (O_2953,N_47598,N_48169);
and UO_2954 (O_2954,N_49924,N_49717);
or UO_2955 (O_2955,N_47795,N_48913);
or UO_2956 (O_2956,N_48749,N_48974);
nand UO_2957 (O_2957,N_49892,N_48933);
nand UO_2958 (O_2958,N_49134,N_48751);
xnor UO_2959 (O_2959,N_48416,N_48017);
nor UO_2960 (O_2960,N_49611,N_48351);
xor UO_2961 (O_2961,N_47986,N_49941);
xnor UO_2962 (O_2962,N_48379,N_47995);
or UO_2963 (O_2963,N_47660,N_49003);
nor UO_2964 (O_2964,N_48674,N_48269);
nand UO_2965 (O_2965,N_47617,N_47763);
and UO_2966 (O_2966,N_49529,N_49591);
and UO_2967 (O_2967,N_49421,N_47870);
xnor UO_2968 (O_2968,N_48277,N_48599);
nand UO_2969 (O_2969,N_48305,N_48943);
xor UO_2970 (O_2970,N_49186,N_47929);
or UO_2971 (O_2971,N_49000,N_48058);
xor UO_2972 (O_2972,N_49833,N_48296);
nor UO_2973 (O_2973,N_47886,N_49474);
nor UO_2974 (O_2974,N_48996,N_49290);
nor UO_2975 (O_2975,N_48451,N_49678);
or UO_2976 (O_2976,N_48505,N_49397);
xnor UO_2977 (O_2977,N_49896,N_48998);
nand UO_2978 (O_2978,N_48994,N_48522);
xnor UO_2979 (O_2979,N_49829,N_49875);
or UO_2980 (O_2980,N_49583,N_48187);
or UO_2981 (O_2981,N_48904,N_49933);
xnor UO_2982 (O_2982,N_49926,N_49545);
nand UO_2983 (O_2983,N_48517,N_49310);
nand UO_2984 (O_2984,N_48574,N_49463);
nor UO_2985 (O_2985,N_48841,N_49615);
and UO_2986 (O_2986,N_48613,N_49345);
or UO_2987 (O_2987,N_48941,N_48454);
nand UO_2988 (O_2988,N_48992,N_49676);
nand UO_2989 (O_2989,N_49933,N_49760);
nand UO_2990 (O_2990,N_49341,N_49443);
nor UO_2991 (O_2991,N_49396,N_48026);
or UO_2992 (O_2992,N_49594,N_49234);
or UO_2993 (O_2993,N_47737,N_48276);
or UO_2994 (O_2994,N_49655,N_48536);
nor UO_2995 (O_2995,N_49798,N_49193);
or UO_2996 (O_2996,N_48729,N_49685);
nand UO_2997 (O_2997,N_48001,N_48131);
nor UO_2998 (O_2998,N_47829,N_49091);
nand UO_2999 (O_2999,N_48913,N_48848);
and UO_3000 (O_3000,N_49407,N_48028);
and UO_3001 (O_3001,N_47795,N_47572);
nor UO_3002 (O_3002,N_47836,N_49412);
xnor UO_3003 (O_3003,N_49615,N_48378);
or UO_3004 (O_3004,N_49820,N_49857);
or UO_3005 (O_3005,N_47730,N_47582);
nand UO_3006 (O_3006,N_49400,N_49517);
and UO_3007 (O_3007,N_49109,N_47952);
nor UO_3008 (O_3008,N_49179,N_47586);
xor UO_3009 (O_3009,N_48230,N_47823);
nor UO_3010 (O_3010,N_49844,N_49292);
or UO_3011 (O_3011,N_49060,N_47664);
xnor UO_3012 (O_3012,N_48474,N_48039);
and UO_3013 (O_3013,N_48216,N_49466);
nor UO_3014 (O_3014,N_48679,N_49060);
and UO_3015 (O_3015,N_49522,N_49501);
and UO_3016 (O_3016,N_48660,N_48348);
xnor UO_3017 (O_3017,N_48258,N_47815);
nand UO_3018 (O_3018,N_49865,N_49796);
and UO_3019 (O_3019,N_48747,N_49705);
nand UO_3020 (O_3020,N_49005,N_49355);
xnor UO_3021 (O_3021,N_48684,N_47543);
and UO_3022 (O_3022,N_47928,N_49167);
and UO_3023 (O_3023,N_49542,N_49457);
and UO_3024 (O_3024,N_49185,N_49497);
nor UO_3025 (O_3025,N_47979,N_49845);
and UO_3026 (O_3026,N_48321,N_49693);
nand UO_3027 (O_3027,N_49492,N_49076);
nand UO_3028 (O_3028,N_48937,N_48967);
and UO_3029 (O_3029,N_48479,N_49101);
and UO_3030 (O_3030,N_49268,N_48970);
nor UO_3031 (O_3031,N_49763,N_49342);
or UO_3032 (O_3032,N_48086,N_49058);
nand UO_3033 (O_3033,N_49995,N_48223);
nand UO_3034 (O_3034,N_47969,N_47939);
xnor UO_3035 (O_3035,N_48668,N_48755);
nand UO_3036 (O_3036,N_49606,N_48412);
nand UO_3037 (O_3037,N_47782,N_49633);
or UO_3038 (O_3038,N_49994,N_47855);
nand UO_3039 (O_3039,N_49053,N_49810);
nor UO_3040 (O_3040,N_49461,N_49096);
or UO_3041 (O_3041,N_48098,N_49088);
nor UO_3042 (O_3042,N_48430,N_49602);
nand UO_3043 (O_3043,N_48859,N_48579);
xor UO_3044 (O_3044,N_49977,N_49574);
or UO_3045 (O_3045,N_49554,N_49164);
nor UO_3046 (O_3046,N_48615,N_48499);
and UO_3047 (O_3047,N_49662,N_47554);
or UO_3048 (O_3048,N_49345,N_49639);
nor UO_3049 (O_3049,N_49297,N_48059);
nand UO_3050 (O_3050,N_48263,N_48600);
nand UO_3051 (O_3051,N_48237,N_49981);
or UO_3052 (O_3052,N_47502,N_49188);
xor UO_3053 (O_3053,N_49232,N_48417);
and UO_3054 (O_3054,N_49465,N_47846);
or UO_3055 (O_3055,N_49567,N_47589);
nor UO_3056 (O_3056,N_48646,N_49612);
nand UO_3057 (O_3057,N_47972,N_49860);
or UO_3058 (O_3058,N_48375,N_47568);
or UO_3059 (O_3059,N_47992,N_49193);
xnor UO_3060 (O_3060,N_49456,N_48148);
nor UO_3061 (O_3061,N_47622,N_48634);
nand UO_3062 (O_3062,N_47814,N_48946);
nand UO_3063 (O_3063,N_49328,N_48861);
or UO_3064 (O_3064,N_48689,N_48059);
or UO_3065 (O_3065,N_47518,N_47534);
and UO_3066 (O_3066,N_48414,N_47665);
nor UO_3067 (O_3067,N_48932,N_49830);
and UO_3068 (O_3068,N_48177,N_49700);
or UO_3069 (O_3069,N_48871,N_49462);
nor UO_3070 (O_3070,N_48902,N_49952);
or UO_3071 (O_3071,N_47735,N_49480);
xor UO_3072 (O_3072,N_48138,N_49765);
nand UO_3073 (O_3073,N_47870,N_48296);
xnor UO_3074 (O_3074,N_48176,N_48392);
nor UO_3075 (O_3075,N_49127,N_47528);
nand UO_3076 (O_3076,N_48202,N_47876);
and UO_3077 (O_3077,N_48450,N_47559);
xor UO_3078 (O_3078,N_48370,N_48248);
xor UO_3079 (O_3079,N_47889,N_48292);
nor UO_3080 (O_3080,N_49092,N_49074);
xor UO_3081 (O_3081,N_49277,N_49339);
and UO_3082 (O_3082,N_48433,N_48672);
nand UO_3083 (O_3083,N_47503,N_49875);
and UO_3084 (O_3084,N_49956,N_48120);
and UO_3085 (O_3085,N_48890,N_47568);
and UO_3086 (O_3086,N_48025,N_49625);
xnor UO_3087 (O_3087,N_47503,N_49031);
nor UO_3088 (O_3088,N_49641,N_49669);
nand UO_3089 (O_3089,N_48332,N_49714);
nor UO_3090 (O_3090,N_48221,N_49594);
nor UO_3091 (O_3091,N_47908,N_48919);
or UO_3092 (O_3092,N_48559,N_47558);
xor UO_3093 (O_3093,N_48001,N_49189);
or UO_3094 (O_3094,N_49845,N_48791);
xnor UO_3095 (O_3095,N_48383,N_47778);
and UO_3096 (O_3096,N_49233,N_48719);
nand UO_3097 (O_3097,N_48723,N_49369);
and UO_3098 (O_3098,N_48525,N_48927);
and UO_3099 (O_3099,N_47881,N_48450);
xnor UO_3100 (O_3100,N_47757,N_48387);
and UO_3101 (O_3101,N_49792,N_48411);
and UO_3102 (O_3102,N_48520,N_48576);
and UO_3103 (O_3103,N_49584,N_48741);
nor UO_3104 (O_3104,N_49094,N_48554);
xor UO_3105 (O_3105,N_48072,N_48485);
and UO_3106 (O_3106,N_49806,N_48431);
nor UO_3107 (O_3107,N_48304,N_49225);
nand UO_3108 (O_3108,N_48040,N_48892);
or UO_3109 (O_3109,N_48745,N_47650);
nand UO_3110 (O_3110,N_47788,N_47641);
and UO_3111 (O_3111,N_48897,N_48812);
xor UO_3112 (O_3112,N_47546,N_48368);
and UO_3113 (O_3113,N_49984,N_49194);
and UO_3114 (O_3114,N_49247,N_48753);
and UO_3115 (O_3115,N_48754,N_49016);
or UO_3116 (O_3116,N_48485,N_48889);
nand UO_3117 (O_3117,N_48676,N_48678);
xnor UO_3118 (O_3118,N_48598,N_47710);
xnor UO_3119 (O_3119,N_49531,N_48016);
nor UO_3120 (O_3120,N_47609,N_47599);
xor UO_3121 (O_3121,N_49735,N_48477);
or UO_3122 (O_3122,N_49410,N_48579);
nand UO_3123 (O_3123,N_47786,N_48155);
or UO_3124 (O_3124,N_49496,N_49877);
nand UO_3125 (O_3125,N_49864,N_49582);
or UO_3126 (O_3126,N_48489,N_49592);
nor UO_3127 (O_3127,N_49059,N_49866);
or UO_3128 (O_3128,N_49272,N_48637);
and UO_3129 (O_3129,N_48739,N_48032);
or UO_3130 (O_3130,N_48149,N_47655);
or UO_3131 (O_3131,N_48777,N_47743);
and UO_3132 (O_3132,N_48481,N_47923);
and UO_3133 (O_3133,N_49836,N_49937);
and UO_3134 (O_3134,N_48534,N_47688);
xor UO_3135 (O_3135,N_48071,N_49260);
and UO_3136 (O_3136,N_48440,N_49555);
or UO_3137 (O_3137,N_49195,N_48289);
nor UO_3138 (O_3138,N_48541,N_47945);
or UO_3139 (O_3139,N_48676,N_49525);
nor UO_3140 (O_3140,N_48380,N_49682);
or UO_3141 (O_3141,N_48987,N_48275);
and UO_3142 (O_3142,N_47806,N_48100);
xnor UO_3143 (O_3143,N_49452,N_49823);
nor UO_3144 (O_3144,N_48671,N_49028);
xnor UO_3145 (O_3145,N_48215,N_49004);
nand UO_3146 (O_3146,N_49255,N_47506);
nand UO_3147 (O_3147,N_49955,N_49922);
xor UO_3148 (O_3148,N_49113,N_47903);
nor UO_3149 (O_3149,N_49306,N_48029);
nor UO_3150 (O_3150,N_49791,N_48162);
nor UO_3151 (O_3151,N_47901,N_47868);
nand UO_3152 (O_3152,N_48604,N_48737);
nand UO_3153 (O_3153,N_49228,N_48823);
nand UO_3154 (O_3154,N_47666,N_48240);
and UO_3155 (O_3155,N_48278,N_48040);
and UO_3156 (O_3156,N_48698,N_48899);
nand UO_3157 (O_3157,N_48996,N_49172);
nand UO_3158 (O_3158,N_47580,N_48011);
nor UO_3159 (O_3159,N_49513,N_48674);
xnor UO_3160 (O_3160,N_47568,N_48561);
xnor UO_3161 (O_3161,N_49828,N_49033);
nand UO_3162 (O_3162,N_48173,N_47594);
and UO_3163 (O_3163,N_47960,N_48520);
nand UO_3164 (O_3164,N_49633,N_47627);
xor UO_3165 (O_3165,N_48785,N_47949);
xnor UO_3166 (O_3166,N_48266,N_48371);
nand UO_3167 (O_3167,N_49875,N_47893);
xnor UO_3168 (O_3168,N_48701,N_48386);
xnor UO_3169 (O_3169,N_48225,N_48308);
and UO_3170 (O_3170,N_48663,N_48320);
xnor UO_3171 (O_3171,N_48785,N_49710);
or UO_3172 (O_3172,N_48804,N_47667);
nor UO_3173 (O_3173,N_47531,N_49657);
nand UO_3174 (O_3174,N_48216,N_49797);
nor UO_3175 (O_3175,N_48715,N_48311);
nor UO_3176 (O_3176,N_47800,N_48882);
or UO_3177 (O_3177,N_48198,N_47552);
or UO_3178 (O_3178,N_49189,N_49153);
xor UO_3179 (O_3179,N_48620,N_47539);
and UO_3180 (O_3180,N_49599,N_47754);
xor UO_3181 (O_3181,N_49515,N_49607);
and UO_3182 (O_3182,N_48750,N_49909);
nand UO_3183 (O_3183,N_47760,N_49904);
nor UO_3184 (O_3184,N_49217,N_49274);
nor UO_3185 (O_3185,N_49563,N_49904);
or UO_3186 (O_3186,N_49641,N_48486);
or UO_3187 (O_3187,N_49141,N_49669);
or UO_3188 (O_3188,N_49269,N_48245);
or UO_3189 (O_3189,N_49232,N_48838);
xor UO_3190 (O_3190,N_49788,N_47587);
nor UO_3191 (O_3191,N_48858,N_48523);
nor UO_3192 (O_3192,N_49649,N_49147);
or UO_3193 (O_3193,N_48773,N_49853);
or UO_3194 (O_3194,N_48111,N_48380);
and UO_3195 (O_3195,N_49004,N_48762);
nand UO_3196 (O_3196,N_48523,N_49133);
or UO_3197 (O_3197,N_47987,N_47717);
or UO_3198 (O_3198,N_49261,N_49062);
or UO_3199 (O_3199,N_48181,N_47836);
nand UO_3200 (O_3200,N_48405,N_47993);
and UO_3201 (O_3201,N_49021,N_48478);
nor UO_3202 (O_3202,N_48428,N_48409);
xor UO_3203 (O_3203,N_49085,N_49706);
or UO_3204 (O_3204,N_49249,N_48022);
and UO_3205 (O_3205,N_48994,N_47531);
and UO_3206 (O_3206,N_49061,N_49409);
xor UO_3207 (O_3207,N_48941,N_48142);
or UO_3208 (O_3208,N_48581,N_48395);
xor UO_3209 (O_3209,N_49000,N_48382);
and UO_3210 (O_3210,N_49344,N_49972);
and UO_3211 (O_3211,N_47951,N_47572);
nand UO_3212 (O_3212,N_49216,N_48397);
nor UO_3213 (O_3213,N_48337,N_48998);
nand UO_3214 (O_3214,N_48228,N_49142);
nor UO_3215 (O_3215,N_49442,N_48588);
xor UO_3216 (O_3216,N_47706,N_49679);
nand UO_3217 (O_3217,N_47978,N_49237);
xnor UO_3218 (O_3218,N_48102,N_48845);
nor UO_3219 (O_3219,N_48173,N_49283);
xnor UO_3220 (O_3220,N_49064,N_48430);
or UO_3221 (O_3221,N_49267,N_48756);
xnor UO_3222 (O_3222,N_48920,N_49473);
nor UO_3223 (O_3223,N_49443,N_49626);
or UO_3224 (O_3224,N_49702,N_48999);
nor UO_3225 (O_3225,N_48385,N_49963);
or UO_3226 (O_3226,N_49229,N_48726);
nand UO_3227 (O_3227,N_48734,N_48881);
xor UO_3228 (O_3228,N_47856,N_47901);
nor UO_3229 (O_3229,N_47652,N_47737);
nor UO_3230 (O_3230,N_48194,N_49742);
nor UO_3231 (O_3231,N_49866,N_49039);
nor UO_3232 (O_3232,N_48549,N_47801);
nor UO_3233 (O_3233,N_49211,N_48378);
nor UO_3234 (O_3234,N_48322,N_48095);
nor UO_3235 (O_3235,N_47902,N_49134);
nand UO_3236 (O_3236,N_48408,N_47530);
nor UO_3237 (O_3237,N_48490,N_49133);
nand UO_3238 (O_3238,N_49922,N_49985);
or UO_3239 (O_3239,N_49100,N_49794);
xor UO_3240 (O_3240,N_47606,N_49483);
and UO_3241 (O_3241,N_48774,N_48342);
nor UO_3242 (O_3242,N_48214,N_48873);
xnor UO_3243 (O_3243,N_49175,N_49990);
nor UO_3244 (O_3244,N_47878,N_49576);
nor UO_3245 (O_3245,N_49032,N_49540);
nand UO_3246 (O_3246,N_47550,N_48427);
nor UO_3247 (O_3247,N_49221,N_49805);
xor UO_3248 (O_3248,N_48928,N_48559);
and UO_3249 (O_3249,N_49300,N_48848);
xnor UO_3250 (O_3250,N_47621,N_48248);
nand UO_3251 (O_3251,N_48003,N_48002);
nor UO_3252 (O_3252,N_49851,N_47986);
nor UO_3253 (O_3253,N_48818,N_49684);
or UO_3254 (O_3254,N_47688,N_49826);
xor UO_3255 (O_3255,N_48177,N_49703);
nand UO_3256 (O_3256,N_49407,N_49598);
nand UO_3257 (O_3257,N_48014,N_49259);
nor UO_3258 (O_3258,N_49621,N_48784);
xnor UO_3259 (O_3259,N_47635,N_49963);
xnor UO_3260 (O_3260,N_49794,N_47671);
nor UO_3261 (O_3261,N_49135,N_48199);
or UO_3262 (O_3262,N_48669,N_48463);
nor UO_3263 (O_3263,N_49324,N_49194);
or UO_3264 (O_3264,N_49589,N_48845);
or UO_3265 (O_3265,N_49271,N_49478);
and UO_3266 (O_3266,N_48508,N_48715);
and UO_3267 (O_3267,N_48629,N_49037);
or UO_3268 (O_3268,N_47727,N_49897);
xnor UO_3269 (O_3269,N_49792,N_49320);
and UO_3270 (O_3270,N_47610,N_47966);
nor UO_3271 (O_3271,N_48151,N_49717);
nand UO_3272 (O_3272,N_49483,N_49812);
and UO_3273 (O_3273,N_48563,N_47628);
nor UO_3274 (O_3274,N_47792,N_49671);
and UO_3275 (O_3275,N_49534,N_49549);
and UO_3276 (O_3276,N_49406,N_48162);
nand UO_3277 (O_3277,N_49447,N_49574);
nand UO_3278 (O_3278,N_47681,N_49852);
or UO_3279 (O_3279,N_48106,N_49176);
xor UO_3280 (O_3280,N_48829,N_49201);
or UO_3281 (O_3281,N_49955,N_49859);
xnor UO_3282 (O_3282,N_49638,N_49172);
or UO_3283 (O_3283,N_48917,N_49094);
nand UO_3284 (O_3284,N_47807,N_48940);
or UO_3285 (O_3285,N_47848,N_48864);
nand UO_3286 (O_3286,N_49033,N_48977);
or UO_3287 (O_3287,N_49487,N_48366);
and UO_3288 (O_3288,N_48425,N_48410);
or UO_3289 (O_3289,N_47932,N_49354);
or UO_3290 (O_3290,N_48244,N_48901);
or UO_3291 (O_3291,N_48591,N_47742);
or UO_3292 (O_3292,N_49945,N_47930);
xnor UO_3293 (O_3293,N_49498,N_48157);
nand UO_3294 (O_3294,N_47604,N_48926);
nand UO_3295 (O_3295,N_49857,N_49626);
or UO_3296 (O_3296,N_49146,N_49079);
xor UO_3297 (O_3297,N_49809,N_48484);
and UO_3298 (O_3298,N_48858,N_49784);
and UO_3299 (O_3299,N_49799,N_48631);
or UO_3300 (O_3300,N_49831,N_47779);
nand UO_3301 (O_3301,N_47915,N_49564);
or UO_3302 (O_3302,N_47501,N_48657);
nand UO_3303 (O_3303,N_49094,N_48910);
and UO_3304 (O_3304,N_48873,N_48994);
nand UO_3305 (O_3305,N_49345,N_49333);
nand UO_3306 (O_3306,N_47785,N_47531);
and UO_3307 (O_3307,N_49648,N_48790);
nand UO_3308 (O_3308,N_48852,N_48497);
xor UO_3309 (O_3309,N_48071,N_48211);
nor UO_3310 (O_3310,N_48821,N_48445);
and UO_3311 (O_3311,N_48430,N_47826);
nand UO_3312 (O_3312,N_47607,N_48319);
xnor UO_3313 (O_3313,N_49438,N_48147);
and UO_3314 (O_3314,N_49525,N_49911);
and UO_3315 (O_3315,N_49165,N_47738);
and UO_3316 (O_3316,N_49506,N_47913);
and UO_3317 (O_3317,N_49669,N_48021);
or UO_3318 (O_3318,N_49957,N_48533);
xnor UO_3319 (O_3319,N_49146,N_48189);
and UO_3320 (O_3320,N_48655,N_48543);
or UO_3321 (O_3321,N_48625,N_48083);
and UO_3322 (O_3322,N_47560,N_48776);
and UO_3323 (O_3323,N_48337,N_49108);
nor UO_3324 (O_3324,N_48206,N_48017);
nor UO_3325 (O_3325,N_48792,N_47557);
nand UO_3326 (O_3326,N_49116,N_49984);
nor UO_3327 (O_3327,N_48316,N_49221);
nand UO_3328 (O_3328,N_48571,N_48218);
nor UO_3329 (O_3329,N_49263,N_49036);
nand UO_3330 (O_3330,N_49728,N_49249);
or UO_3331 (O_3331,N_48618,N_49395);
nor UO_3332 (O_3332,N_49992,N_49485);
nor UO_3333 (O_3333,N_49759,N_49091);
nor UO_3334 (O_3334,N_48497,N_49627);
nand UO_3335 (O_3335,N_49922,N_47869);
and UO_3336 (O_3336,N_47639,N_49917);
nand UO_3337 (O_3337,N_49374,N_47636);
nor UO_3338 (O_3338,N_49230,N_47510);
and UO_3339 (O_3339,N_47656,N_48534);
and UO_3340 (O_3340,N_49894,N_49110);
and UO_3341 (O_3341,N_49969,N_49370);
nor UO_3342 (O_3342,N_48665,N_49059);
nor UO_3343 (O_3343,N_48928,N_48891);
and UO_3344 (O_3344,N_48496,N_47667);
xnor UO_3345 (O_3345,N_48993,N_48000);
or UO_3346 (O_3346,N_47891,N_47872);
xnor UO_3347 (O_3347,N_48445,N_48800);
nor UO_3348 (O_3348,N_48501,N_48355);
xor UO_3349 (O_3349,N_49617,N_48148);
or UO_3350 (O_3350,N_49687,N_48581);
xnor UO_3351 (O_3351,N_49914,N_49877);
xor UO_3352 (O_3352,N_48233,N_48504);
xnor UO_3353 (O_3353,N_49729,N_47558);
xnor UO_3354 (O_3354,N_47641,N_49798);
and UO_3355 (O_3355,N_48767,N_49916);
or UO_3356 (O_3356,N_49049,N_49469);
and UO_3357 (O_3357,N_47891,N_47954);
xor UO_3358 (O_3358,N_47647,N_49301);
nor UO_3359 (O_3359,N_47810,N_49173);
and UO_3360 (O_3360,N_47672,N_49006);
nor UO_3361 (O_3361,N_49396,N_48653);
nor UO_3362 (O_3362,N_47829,N_49603);
nand UO_3363 (O_3363,N_48309,N_48746);
and UO_3364 (O_3364,N_49877,N_49431);
or UO_3365 (O_3365,N_49414,N_49141);
xor UO_3366 (O_3366,N_48085,N_48862);
or UO_3367 (O_3367,N_49490,N_48259);
or UO_3368 (O_3368,N_48029,N_48671);
xor UO_3369 (O_3369,N_49581,N_48849);
xnor UO_3370 (O_3370,N_49208,N_49639);
xnor UO_3371 (O_3371,N_49829,N_47843);
xnor UO_3372 (O_3372,N_47702,N_48542);
nand UO_3373 (O_3373,N_49667,N_49566);
xnor UO_3374 (O_3374,N_48428,N_48364);
or UO_3375 (O_3375,N_47514,N_48204);
nor UO_3376 (O_3376,N_49676,N_48684);
or UO_3377 (O_3377,N_48402,N_47791);
and UO_3378 (O_3378,N_49145,N_48914);
xnor UO_3379 (O_3379,N_47500,N_47773);
xor UO_3380 (O_3380,N_47962,N_49307);
nand UO_3381 (O_3381,N_49907,N_48131);
and UO_3382 (O_3382,N_49598,N_49491);
or UO_3383 (O_3383,N_48074,N_48964);
nand UO_3384 (O_3384,N_47786,N_47968);
nor UO_3385 (O_3385,N_47732,N_49648);
and UO_3386 (O_3386,N_48623,N_48796);
xnor UO_3387 (O_3387,N_48925,N_47539);
nand UO_3388 (O_3388,N_47802,N_49516);
xnor UO_3389 (O_3389,N_48219,N_48850);
xnor UO_3390 (O_3390,N_47877,N_49783);
and UO_3391 (O_3391,N_49783,N_47717);
or UO_3392 (O_3392,N_48862,N_48155);
nor UO_3393 (O_3393,N_48245,N_49813);
and UO_3394 (O_3394,N_49330,N_49428);
nand UO_3395 (O_3395,N_47643,N_48450);
xnor UO_3396 (O_3396,N_48316,N_48533);
or UO_3397 (O_3397,N_49181,N_47715);
nor UO_3398 (O_3398,N_49950,N_48626);
xor UO_3399 (O_3399,N_49174,N_49805);
and UO_3400 (O_3400,N_49038,N_48339);
nor UO_3401 (O_3401,N_49092,N_48270);
nor UO_3402 (O_3402,N_47660,N_48596);
xor UO_3403 (O_3403,N_48289,N_47908);
nor UO_3404 (O_3404,N_47848,N_48905);
nor UO_3405 (O_3405,N_48498,N_47650);
and UO_3406 (O_3406,N_48321,N_49229);
or UO_3407 (O_3407,N_49459,N_47652);
or UO_3408 (O_3408,N_49532,N_48382);
nor UO_3409 (O_3409,N_49634,N_48037);
xor UO_3410 (O_3410,N_49073,N_49072);
or UO_3411 (O_3411,N_47898,N_49106);
or UO_3412 (O_3412,N_47798,N_47545);
xor UO_3413 (O_3413,N_48519,N_47824);
nand UO_3414 (O_3414,N_47680,N_48918);
nor UO_3415 (O_3415,N_49275,N_48008);
nor UO_3416 (O_3416,N_48459,N_48849);
and UO_3417 (O_3417,N_49519,N_49738);
or UO_3418 (O_3418,N_49625,N_48669);
and UO_3419 (O_3419,N_49760,N_47584);
nor UO_3420 (O_3420,N_48009,N_49929);
and UO_3421 (O_3421,N_47569,N_48437);
nor UO_3422 (O_3422,N_48510,N_49096);
and UO_3423 (O_3423,N_49970,N_47513);
or UO_3424 (O_3424,N_47742,N_48207);
nor UO_3425 (O_3425,N_47857,N_47699);
nand UO_3426 (O_3426,N_48498,N_49128);
and UO_3427 (O_3427,N_47997,N_49773);
nor UO_3428 (O_3428,N_49849,N_49641);
xnor UO_3429 (O_3429,N_48180,N_47740);
nand UO_3430 (O_3430,N_48226,N_48419);
nand UO_3431 (O_3431,N_48479,N_48354);
xnor UO_3432 (O_3432,N_49756,N_48778);
or UO_3433 (O_3433,N_49196,N_47730);
xnor UO_3434 (O_3434,N_48102,N_49624);
and UO_3435 (O_3435,N_47951,N_49777);
nand UO_3436 (O_3436,N_49597,N_49843);
nor UO_3437 (O_3437,N_48421,N_47796);
xor UO_3438 (O_3438,N_48898,N_47850);
and UO_3439 (O_3439,N_49927,N_47750);
nand UO_3440 (O_3440,N_47607,N_49663);
or UO_3441 (O_3441,N_48167,N_49288);
or UO_3442 (O_3442,N_47931,N_49709);
nand UO_3443 (O_3443,N_48015,N_48685);
or UO_3444 (O_3444,N_49666,N_49164);
and UO_3445 (O_3445,N_48155,N_49621);
xor UO_3446 (O_3446,N_49819,N_48369);
and UO_3447 (O_3447,N_47985,N_47722);
xnor UO_3448 (O_3448,N_48553,N_48376);
xor UO_3449 (O_3449,N_49838,N_49968);
nand UO_3450 (O_3450,N_48317,N_49354);
and UO_3451 (O_3451,N_48064,N_49277);
or UO_3452 (O_3452,N_48803,N_49843);
or UO_3453 (O_3453,N_47829,N_49234);
nand UO_3454 (O_3454,N_48765,N_48533);
xor UO_3455 (O_3455,N_49734,N_49108);
nor UO_3456 (O_3456,N_49665,N_47685);
xor UO_3457 (O_3457,N_47583,N_49893);
nand UO_3458 (O_3458,N_49027,N_49099);
nand UO_3459 (O_3459,N_48962,N_47759);
or UO_3460 (O_3460,N_48304,N_49801);
or UO_3461 (O_3461,N_48755,N_48850);
and UO_3462 (O_3462,N_49796,N_47761);
xor UO_3463 (O_3463,N_47893,N_49344);
or UO_3464 (O_3464,N_47929,N_47513);
and UO_3465 (O_3465,N_48746,N_49380);
nand UO_3466 (O_3466,N_49958,N_48559);
and UO_3467 (O_3467,N_49759,N_49745);
nor UO_3468 (O_3468,N_49770,N_47985);
and UO_3469 (O_3469,N_49711,N_48598);
or UO_3470 (O_3470,N_49228,N_48009);
nor UO_3471 (O_3471,N_48246,N_47585);
or UO_3472 (O_3472,N_47786,N_48674);
and UO_3473 (O_3473,N_49693,N_47510);
or UO_3474 (O_3474,N_48464,N_48061);
xnor UO_3475 (O_3475,N_49319,N_49964);
nor UO_3476 (O_3476,N_48332,N_48761);
nor UO_3477 (O_3477,N_48403,N_48198);
nand UO_3478 (O_3478,N_49315,N_49561);
or UO_3479 (O_3479,N_49496,N_49320);
nor UO_3480 (O_3480,N_48577,N_49241);
and UO_3481 (O_3481,N_49758,N_48878);
nor UO_3482 (O_3482,N_49817,N_47934);
and UO_3483 (O_3483,N_49799,N_47735);
and UO_3484 (O_3484,N_47529,N_49413);
xnor UO_3485 (O_3485,N_49363,N_49703);
and UO_3486 (O_3486,N_47879,N_48729);
nand UO_3487 (O_3487,N_49651,N_49478);
or UO_3488 (O_3488,N_47735,N_48473);
and UO_3489 (O_3489,N_49623,N_47568);
nand UO_3490 (O_3490,N_48158,N_48936);
nand UO_3491 (O_3491,N_47764,N_47977);
or UO_3492 (O_3492,N_47704,N_48495);
nand UO_3493 (O_3493,N_48933,N_47800);
and UO_3494 (O_3494,N_48474,N_47728);
and UO_3495 (O_3495,N_49112,N_49121);
nor UO_3496 (O_3496,N_49630,N_48579);
and UO_3497 (O_3497,N_48211,N_49491);
nor UO_3498 (O_3498,N_49980,N_48833);
nand UO_3499 (O_3499,N_48498,N_49824);
nand UO_3500 (O_3500,N_48571,N_49517);
or UO_3501 (O_3501,N_48027,N_48200);
and UO_3502 (O_3502,N_47895,N_49309);
or UO_3503 (O_3503,N_47708,N_48066);
xor UO_3504 (O_3504,N_47680,N_48171);
nor UO_3505 (O_3505,N_49736,N_48742);
or UO_3506 (O_3506,N_48283,N_48891);
nand UO_3507 (O_3507,N_47980,N_47625);
nand UO_3508 (O_3508,N_47878,N_47891);
xor UO_3509 (O_3509,N_49072,N_48588);
nand UO_3510 (O_3510,N_48311,N_49305);
xnor UO_3511 (O_3511,N_48379,N_48466);
and UO_3512 (O_3512,N_48801,N_49488);
nand UO_3513 (O_3513,N_47570,N_49337);
or UO_3514 (O_3514,N_48695,N_49904);
xor UO_3515 (O_3515,N_48187,N_48130);
and UO_3516 (O_3516,N_48234,N_48480);
or UO_3517 (O_3517,N_48950,N_48032);
or UO_3518 (O_3518,N_49019,N_48271);
nor UO_3519 (O_3519,N_47556,N_49077);
and UO_3520 (O_3520,N_47615,N_49503);
nand UO_3521 (O_3521,N_47972,N_49783);
or UO_3522 (O_3522,N_47884,N_48403);
xor UO_3523 (O_3523,N_49191,N_47522);
xor UO_3524 (O_3524,N_48654,N_48836);
or UO_3525 (O_3525,N_49827,N_47903);
xnor UO_3526 (O_3526,N_49583,N_48885);
and UO_3527 (O_3527,N_49968,N_48304);
nand UO_3528 (O_3528,N_48272,N_48286);
xnor UO_3529 (O_3529,N_48182,N_49345);
nor UO_3530 (O_3530,N_48973,N_47569);
and UO_3531 (O_3531,N_49962,N_47973);
nand UO_3532 (O_3532,N_49995,N_49791);
xor UO_3533 (O_3533,N_47570,N_48876);
and UO_3534 (O_3534,N_47543,N_47937);
nand UO_3535 (O_3535,N_47887,N_47745);
and UO_3536 (O_3536,N_48345,N_48683);
nor UO_3537 (O_3537,N_47822,N_48512);
xor UO_3538 (O_3538,N_47673,N_49819);
xnor UO_3539 (O_3539,N_48914,N_48055);
nor UO_3540 (O_3540,N_48711,N_47554);
and UO_3541 (O_3541,N_47945,N_49685);
nand UO_3542 (O_3542,N_49921,N_47867);
nand UO_3543 (O_3543,N_49829,N_48174);
nand UO_3544 (O_3544,N_48708,N_48364);
and UO_3545 (O_3545,N_47701,N_49903);
or UO_3546 (O_3546,N_49302,N_49744);
or UO_3547 (O_3547,N_49891,N_47603);
or UO_3548 (O_3548,N_48685,N_48248);
nand UO_3549 (O_3549,N_49648,N_49841);
xor UO_3550 (O_3550,N_48223,N_48020);
nand UO_3551 (O_3551,N_47869,N_49557);
nand UO_3552 (O_3552,N_49508,N_47708);
nor UO_3553 (O_3553,N_49070,N_49060);
or UO_3554 (O_3554,N_47890,N_49251);
or UO_3555 (O_3555,N_48600,N_49510);
xor UO_3556 (O_3556,N_49414,N_49692);
nand UO_3557 (O_3557,N_47909,N_49535);
or UO_3558 (O_3558,N_47947,N_48101);
and UO_3559 (O_3559,N_49225,N_48059);
nor UO_3560 (O_3560,N_48934,N_49800);
nor UO_3561 (O_3561,N_48018,N_48686);
and UO_3562 (O_3562,N_47662,N_48791);
nor UO_3563 (O_3563,N_49621,N_49242);
xor UO_3564 (O_3564,N_48837,N_47985);
nor UO_3565 (O_3565,N_49730,N_47979);
nand UO_3566 (O_3566,N_48049,N_47693);
and UO_3567 (O_3567,N_48379,N_48515);
nand UO_3568 (O_3568,N_49518,N_49569);
nand UO_3569 (O_3569,N_49860,N_47790);
or UO_3570 (O_3570,N_49368,N_47602);
nand UO_3571 (O_3571,N_48133,N_47887);
or UO_3572 (O_3572,N_48953,N_47797);
and UO_3573 (O_3573,N_49717,N_48202);
and UO_3574 (O_3574,N_47940,N_49815);
nand UO_3575 (O_3575,N_47972,N_48540);
xnor UO_3576 (O_3576,N_48801,N_49995);
xor UO_3577 (O_3577,N_48730,N_48296);
nor UO_3578 (O_3578,N_48116,N_47632);
nand UO_3579 (O_3579,N_48273,N_49488);
nor UO_3580 (O_3580,N_48521,N_48272);
and UO_3581 (O_3581,N_49733,N_48958);
nor UO_3582 (O_3582,N_48904,N_49266);
or UO_3583 (O_3583,N_47785,N_47621);
and UO_3584 (O_3584,N_47979,N_48579);
nand UO_3585 (O_3585,N_47794,N_49792);
or UO_3586 (O_3586,N_49036,N_47642);
nor UO_3587 (O_3587,N_49424,N_48708);
nor UO_3588 (O_3588,N_48289,N_47712);
or UO_3589 (O_3589,N_47824,N_49027);
or UO_3590 (O_3590,N_49505,N_48746);
nand UO_3591 (O_3591,N_47790,N_49601);
xnor UO_3592 (O_3592,N_47656,N_49381);
xor UO_3593 (O_3593,N_48165,N_48542);
or UO_3594 (O_3594,N_49628,N_48955);
nand UO_3595 (O_3595,N_48975,N_49748);
nand UO_3596 (O_3596,N_48945,N_49184);
and UO_3597 (O_3597,N_48499,N_49763);
nor UO_3598 (O_3598,N_48336,N_49390);
and UO_3599 (O_3599,N_48495,N_49492);
or UO_3600 (O_3600,N_48532,N_48978);
or UO_3601 (O_3601,N_48192,N_48188);
nand UO_3602 (O_3602,N_49556,N_48858);
or UO_3603 (O_3603,N_48679,N_49314);
xnor UO_3604 (O_3604,N_48897,N_48961);
nand UO_3605 (O_3605,N_48169,N_49589);
or UO_3606 (O_3606,N_47781,N_48890);
or UO_3607 (O_3607,N_49607,N_48278);
xnor UO_3608 (O_3608,N_49156,N_47990);
nand UO_3609 (O_3609,N_47675,N_49182);
or UO_3610 (O_3610,N_48945,N_47685);
nand UO_3611 (O_3611,N_48980,N_49247);
nand UO_3612 (O_3612,N_48892,N_47603);
or UO_3613 (O_3613,N_47586,N_48285);
or UO_3614 (O_3614,N_48018,N_48418);
nand UO_3615 (O_3615,N_48572,N_48155);
or UO_3616 (O_3616,N_49385,N_47681);
nand UO_3617 (O_3617,N_48426,N_48990);
or UO_3618 (O_3618,N_47509,N_49838);
nor UO_3619 (O_3619,N_49697,N_48480);
and UO_3620 (O_3620,N_49587,N_48879);
and UO_3621 (O_3621,N_49648,N_47632);
nand UO_3622 (O_3622,N_48457,N_47574);
xnor UO_3623 (O_3623,N_49754,N_49815);
nor UO_3624 (O_3624,N_47862,N_47553);
and UO_3625 (O_3625,N_49750,N_47598);
and UO_3626 (O_3626,N_48626,N_48385);
nand UO_3627 (O_3627,N_48868,N_48798);
and UO_3628 (O_3628,N_48148,N_49387);
or UO_3629 (O_3629,N_47693,N_49499);
nor UO_3630 (O_3630,N_47810,N_48073);
or UO_3631 (O_3631,N_48333,N_48277);
and UO_3632 (O_3632,N_49367,N_49364);
nand UO_3633 (O_3633,N_48072,N_48774);
nand UO_3634 (O_3634,N_49498,N_49193);
nand UO_3635 (O_3635,N_49611,N_48649);
nor UO_3636 (O_3636,N_49966,N_47739);
nor UO_3637 (O_3637,N_47705,N_47769);
nand UO_3638 (O_3638,N_48428,N_48795);
and UO_3639 (O_3639,N_47808,N_48244);
xnor UO_3640 (O_3640,N_49434,N_49378);
or UO_3641 (O_3641,N_49678,N_48763);
and UO_3642 (O_3642,N_49555,N_49372);
or UO_3643 (O_3643,N_48558,N_49181);
nand UO_3644 (O_3644,N_48373,N_48186);
or UO_3645 (O_3645,N_47623,N_49952);
nand UO_3646 (O_3646,N_48729,N_48756);
xor UO_3647 (O_3647,N_49186,N_48341);
nand UO_3648 (O_3648,N_49413,N_49285);
or UO_3649 (O_3649,N_48747,N_49527);
and UO_3650 (O_3650,N_49119,N_48198);
nor UO_3651 (O_3651,N_47830,N_49287);
xor UO_3652 (O_3652,N_49483,N_48971);
nand UO_3653 (O_3653,N_48569,N_47517);
and UO_3654 (O_3654,N_47524,N_48409);
nor UO_3655 (O_3655,N_48372,N_49432);
xor UO_3656 (O_3656,N_48274,N_47992);
and UO_3657 (O_3657,N_48662,N_49643);
xnor UO_3658 (O_3658,N_49686,N_47646);
or UO_3659 (O_3659,N_49070,N_48052);
nor UO_3660 (O_3660,N_49073,N_47896);
or UO_3661 (O_3661,N_48588,N_49368);
or UO_3662 (O_3662,N_48707,N_49398);
or UO_3663 (O_3663,N_47549,N_47853);
nand UO_3664 (O_3664,N_48149,N_49858);
and UO_3665 (O_3665,N_48481,N_48029);
nand UO_3666 (O_3666,N_48530,N_48216);
and UO_3667 (O_3667,N_49133,N_47986);
and UO_3668 (O_3668,N_48245,N_49868);
or UO_3669 (O_3669,N_48255,N_48519);
nor UO_3670 (O_3670,N_47904,N_47768);
nor UO_3671 (O_3671,N_48826,N_49662);
and UO_3672 (O_3672,N_47821,N_49692);
nand UO_3673 (O_3673,N_48734,N_47977);
and UO_3674 (O_3674,N_49449,N_48917);
or UO_3675 (O_3675,N_49162,N_47988);
nor UO_3676 (O_3676,N_48169,N_49788);
and UO_3677 (O_3677,N_48995,N_49704);
and UO_3678 (O_3678,N_47878,N_49167);
or UO_3679 (O_3679,N_49347,N_49655);
and UO_3680 (O_3680,N_49075,N_49021);
or UO_3681 (O_3681,N_48430,N_48092);
or UO_3682 (O_3682,N_48160,N_48502);
and UO_3683 (O_3683,N_49950,N_49795);
and UO_3684 (O_3684,N_48462,N_48314);
nor UO_3685 (O_3685,N_47764,N_47934);
nand UO_3686 (O_3686,N_47628,N_48104);
nand UO_3687 (O_3687,N_47925,N_48465);
or UO_3688 (O_3688,N_49382,N_49799);
nand UO_3689 (O_3689,N_48518,N_49216);
xnor UO_3690 (O_3690,N_48364,N_49840);
or UO_3691 (O_3691,N_48755,N_49280);
or UO_3692 (O_3692,N_49460,N_48817);
and UO_3693 (O_3693,N_49694,N_47610);
nand UO_3694 (O_3694,N_48676,N_49975);
nor UO_3695 (O_3695,N_48404,N_47568);
nand UO_3696 (O_3696,N_47592,N_48170);
nand UO_3697 (O_3697,N_49475,N_48938);
nor UO_3698 (O_3698,N_49711,N_47763);
and UO_3699 (O_3699,N_47639,N_47850);
nor UO_3700 (O_3700,N_48232,N_48612);
nand UO_3701 (O_3701,N_49760,N_49845);
nor UO_3702 (O_3702,N_48350,N_47642);
nand UO_3703 (O_3703,N_47897,N_49180);
and UO_3704 (O_3704,N_47790,N_49993);
nor UO_3705 (O_3705,N_49321,N_48381);
and UO_3706 (O_3706,N_49437,N_49361);
and UO_3707 (O_3707,N_49073,N_48620);
xor UO_3708 (O_3708,N_48248,N_48755);
nand UO_3709 (O_3709,N_49680,N_48453);
or UO_3710 (O_3710,N_49323,N_47763);
xnor UO_3711 (O_3711,N_48761,N_49385);
nand UO_3712 (O_3712,N_48877,N_48016);
or UO_3713 (O_3713,N_48461,N_49849);
nor UO_3714 (O_3714,N_48423,N_49081);
or UO_3715 (O_3715,N_47644,N_49334);
and UO_3716 (O_3716,N_49830,N_49477);
nand UO_3717 (O_3717,N_49768,N_48053);
xnor UO_3718 (O_3718,N_48674,N_48145);
nor UO_3719 (O_3719,N_48786,N_49354);
or UO_3720 (O_3720,N_49565,N_49068);
nor UO_3721 (O_3721,N_49259,N_49091);
nor UO_3722 (O_3722,N_48067,N_48819);
nor UO_3723 (O_3723,N_48041,N_49037);
xor UO_3724 (O_3724,N_49479,N_48901);
nor UO_3725 (O_3725,N_48957,N_49818);
nand UO_3726 (O_3726,N_47792,N_48828);
and UO_3727 (O_3727,N_48450,N_49479);
xor UO_3728 (O_3728,N_49819,N_49180);
nand UO_3729 (O_3729,N_48815,N_48197);
and UO_3730 (O_3730,N_49222,N_49545);
nor UO_3731 (O_3731,N_48659,N_49652);
and UO_3732 (O_3732,N_49108,N_49899);
nor UO_3733 (O_3733,N_48624,N_47736);
or UO_3734 (O_3734,N_49331,N_47949);
nand UO_3735 (O_3735,N_49477,N_49185);
xor UO_3736 (O_3736,N_49603,N_49449);
and UO_3737 (O_3737,N_49293,N_49122);
and UO_3738 (O_3738,N_48201,N_47516);
or UO_3739 (O_3739,N_48140,N_47549);
nor UO_3740 (O_3740,N_47814,N_47541);
nor UO_3741 (O_3741,N_48212,N_48048);
or UO_3742 (O_3742,N_49839,N_48151);
xnor UO_3743 (O_3743,N_49747,N_49035);
xor UO_3744 (O_3744,N_49997,N_49472);
nand UO_3745 (O_3745,N_49460,N_49051);
nor UO_3746 (O_3746,N_47949,N_48820);
or UO_3747 (O_3747,N_48194,N_49936);
xnor UO_3748 (O_3748,N_48088,N_49907);
nor UO_3749 (O_3749,N_48856,N_49980);
xnor UO_3750 (O_3750,N_48241,N_48835);
nor UO_3751 (O_3751,N_48233,N_47962);
nand UO_3752 (O_3752,N_49684,N_47782);
nor UO_3753 (O_3753,N_48099,N_49131);
nand UO_3754 (O_3754,N_47728,N_49952);
xor UO_3755 (O_3755,N_48133,N_48236);
nand UO_3756 (O_3756,N_48730,N_49671);
nand UO_3757 (O_3757,N_49725,N_49316);
nor UO_3758 (O_3758,N_48632,N_47533);
nor UO_3759 (O_3759,N_47521,N_47694);
nand UO_3760 (O_3760,N_48782,N_49055);
nor UO_3761 (O_3761,N_48471,N_48610);
xor UO_3762 (O_3762,N_49260,N_47594);
or UO_3763 (O_3763,N_48771,N_48893);
xor UO_3764 (O_3764,N_48428,N_47858);
or UO_3765 (O_3765,N_49916,N_49269);
xor UO_3766 (O_3766,N_47596,N_49327);
nor UO_3767 (O_3767,N_47703,N_48602);
nor UO_3768 (O_3768,N_47818,N_49054);
and UO_3769 (O_3769,N_48170,N_49366);
and UO_3770 (O_3770,N_49157,N_48629);
nand UO_3771 (O_3771,N_47704,N_48449);
and UO_3772 (O_3772,N_48028,N_47960);
or UO_3773 (O_3773,N_49816,N_47540);
and UO_3774 (O_3774,N_49959,N_47790);
nand UO_3775 (O_3775,N_48356,N_47990);
xnor UO_3776 (O_3776,N_49146,N_48024);
nor UO_3777 (O_3777,N_47685,N_49374);
xor UO_3778 (O_3778,N_48154,N_47850);
nor UO_3779 (O_3779,N_49001,N_49536);
nor UO_3780 (O_3780,N_48246,N_48841);
and UO_3781 (O_3781,N_49038,N_49039);
and UO_3782 (O_3782,N_49779,N_49180);
xor UO_3783 (O_3783,N_49975,N_48296);
xor UO_3784 (O_3784,N_48967,N_48019);
nor UO_3785 (O_3785,N_49267,N_47520);
and UO_3786 (O_3786,N_48448,N_49144);
or UO_3787 (O_3787,N_48834,N_49828);
nand UO_3788 (O_3788,N_47849,N_47823);
nand UO_3789 (O_3789,N_47974,N_49196);
nand UO_3790 (O_3790,N_48462,N_47958);
nor UO_3791 (O_3791,N_49466,N_49607);
or UO_3792 (O_3792,N_49548,N_48674);
and UO_3793 (O_3793,N_47518,N_49934);
and UO_3794 (O_3794,N_49737,N_49623);
nor UO_3795 (O_3795,N_48145,N_48582);
and UO_3796 (O_3796,N_48323,N_49674);
nor UO_3797 (O_3797,N_47857,N_47507);
nand UO_3798 (O_3798,N_47919,N_47782);
nor UO_3799 (O_3799,N_47935,N_48177);
or UO_3800 (O_3800,N_47664,N_49530);
nor UO_3801 (O_3801,N_49566,N_48290);
nor UO_3802 (O_3802,N_47984,N_48047);
nor UO_3803 (O_3803,N_48480,N_48366);
nand UO_3804 (O_3804,N_48776,N_48183);
and UO_3805 (O_3805,N_47822,N_48461);
and UO_3806 (O_3806,N_48369,N_49967);
nor UO_3807 (O_3807,N_49581,N_48312);
xor UO_3808 (O_3808,N_49934,N_48857);
nor UO_3809 (O_3809,N_49622,N_47996);
nand UO_3810 (O_3810,N_47903,N_47558);
nand UO_3811 (O_3811,N_49248,N_49795);
or UO_3812 (O_3812,N_47831,N_47979);
and UO_3813 (O_3813,N_48471,N_47776);
xnor UO_3814 (O_3814,N_49177,N_48278);
or UO_3815 (O_3815,N_49593,N_48718);
and UO_3816 (O_3816,N_49586,N_48407);
nor UO_3817 (O_3817,N_49722,N_49540);
xnor UO_3818 (O_3818,N_49238,N_48561);
nor UO_3819 (O_3819,N_49167,N_48706);
xor UO_3820 (O_3820,N_49954,N_48642);
or UO_3821 (O_3821,N_48819,N_48648);
or UO_3822 (O_3822,N_49093,N_49592);
nor UO_3823 (O_3823,N_48774,N_49493);
and UO_3824 (O_3824,N_48931,N_49587);
and UO_3825 (O_3825,N_49798,N_47818);
nor UO_3826 (O_3826,N_49409,N_47689);
or UO_3827 (O_3827,N_48937,N_48925);
and UO_3828 (O_3828,N_47665,N_48513);
nand UO_3829 (O_3829,N_49023,N_48403);
xnor UO_3830 (O_3830,N_47933,N_48602);
and UO_3831 (O_3831,N_49299,N_48455);
nor UO_3832 (O_3832,N_49790,N_49663);
xor UO_3833 (O_3833,N_48255,N_49905);
nor UO_3834 (O_3834,N_49542,N_48490);
and UO_3835 (O_3835,N_47554,N_48065);
xnor UO_3836 (O_3836,N_49001,N_49594);
nand UO_3837 (O_3837,N_49219,N_49896);
xnor UO_3838 (O_3838,N_48944,N_48870);
nor UO_3839 (O_3839,N_49756,N_48791);
and UO_3840 (O_3840,N_47697,N_48291);
xor UO_3841 (O_3841,N_49272,N_49194);
xnor UO_3842 (O_3842,N_49071,N_49741);
xor UO_3843 (O_3843,N_48128,N_48865);
or UO_3844 (O_3844,N_48478,N_48441);
or UO_3845 (O_3845,N_49299,N_47561);
or UO_3846 (O_3846,N_47607,N_47893);
nand UO_3847 (O_3847,N_49230,N_49239);
nand UO_3848 (O_3848,N_49180,N_49755);
nand UO_3849 (O_3849,N_48620,N_48455);
nand UO_3850 (O_3850,N_48796,N_47693);
nand UO_3851 (O_3851,N_49259,N_47896);
nand UO_3852 (O_3852,N_48032,N_49705);
nor UO_3853 (O_3853,N_48800,N_48207);
and UO_3854 (O_3854,N_49389,N_48794);
nand UO_3855 (O_3855,N_47585,N_49689);
nand UO_3856 (O_3856,N_48505,N_49918);
or UO_3857 (O_3857,N_48487,N_49200);
or UO_3858 (O_3858,N_48632,N_48372);
xnor UO_3859 (O_3859,N_48074,N_49818);
xnor UO_3860 (O_3860,N_48615,N_49964);
xnor UO_3861 (O_3861,N_49167,N_48580);
and UO_3862 (O_3862,N_49504,N_49025);
or UO_3863 (O_3863,N_49794,N_48293);
or UO_3864 (O_3864,N_49929,N_47718);
or UO_3865 (O_3865,N_47978,N_49952);
or UO_3866 (O_3866,N_47614,N_48708);
xor UO_3867 (O_3867,N_49056,N_49512);
or UO_3868 (O_3868,N_47743,N_49571);
xor UO_3869 (O_3869,N_47787,N_49788);
nor UO_3870 (O_3870,N_48743,N_48204);
or UO_3871 (O_3871,N_49842,N_49085);
xnor UO_3872 (O_3872,N_47762,N_47662);
nand UO_3873 (O_3873,N_48814,N_48968);
nor UO_3874 (O_3874,N_47743,N_49707);
and UO_3875 (O_3875,N_47794,N_47572);
or UO_3876 (O_3876,N_49372,N_49445);
and UO_3877 (O_3877,N_48121,N_47572);
nand UO_3878 (O_3878,N_49405,N_48888);
nand UO_3879 (O_3879,N_48438,N_48873);
nand UO_3880 (O_3880,N_49490,N_48822);
or UO_3881 (O_3881,N_48439,N_47572);
nand UO_3882 (O_3882,N_49197,N_48206);
or UO_3883 (O_3883,N_48971,N_49347);
and UO_3884 (O_3884,N_48404,N_48569);
nand UO_3885 (O_3885,N_48252,N_49274);
or UO_3886 (O_3886,N_49720,N_48808);
nor UO_3887 (O_3887,N_49856,N_49406);
and UO_3888 (O_3888,N_49451,N_49589);
nor UO_3889 (O_3889,N_48488,N_47515);
nand UO_3890 (O_3890,N_48999,N_49521);
xnor UO_3891 (O_3891,N_48362,N_49331);
nand UO_3892 (O_3892,N_47763,N_47667);
nand UO_3893 (O_3893,N_47936,N_48345);
nor UO_3894 (O_3894,N_47966,N_48728);
nand UO_3895 (O_3895,N_49170,N_49118);
xor UO_3896 (O_3896,N_47665,N_49717);
or UO_3897 (O_3897,N_48009,N_47773);
or UO_3898 (O_3898,N_48304,N_49994);
xnor UO_3899 (O_3899,N_49732,N_47947);
or UO_3900 (O_3900,N_49435,N_48289);
xor UO_3901 (O_3901,N_48147,N_49366);
xnor UO_3902 (O_3902,N_47504,N_49653);
xnor UO_3903 (O_3903,N_48303,N_49025);
and UO_3904 (O_3904,N_49054,N_48804);
and UO_3905 (O_3905,N_49772,N_49442);
nand UO_3906 (O_3906,N_48583,N_48395);
and UO_3907 (O_3907,N_48194,N_49121);
or UO_3908 (O_3908,N_48191,N_49392);
nor UO_3909 (O_3909,N_48747,N_49335);
and UO_3910 (O_3910,N_48769,N_49535);
and UO_3911 (O_3911,N_48969,N_47816);
nor UO_3912 (O_3912,N_48879,N_48645);
and UO_3913 (O_3913,N_49034,N_47974);
and UO_3914 (O_3914,N_49138,N_48421);
and UO_3915 (O_3915,N_47903,N_48965);
nand UO_3916 (O_3916,N_48525,N_49477);
and UO_3917 (O_3917,N_47803,N_48625);
and UO_3918 (O_3918,N_49545,N_47860);
xnor UO_3919 (O_3919,N_49522,N_48480);
and UO_3920 (O_3920,N_47649,N_48138);
or UO_3921 (O_3921,N_48533,N_48698);
xor UO_3922 (O_3922,N_47737,N_48401);
and UO_3923 (O_3923,N_49871,N_48570);
or UO_3924 (O_3924,N_48754,N_49686);
nand UO_3925 (O_3925,N_47865,N_49130);
nand UO_3926 (O_3926,N_48520,N_47893);
xnor UO_3927 (O_3927,N_47528,N_47548);
and UO_3928 (O_3928,N_47527,N_48445);
and UO_3929 (O_3929,N_48726,N_49661);
xnor UO_3930 (O_3930,N_48714,N_48383);
or UO_3931 (O_3931,N_48737,N_47970);
xor UO_3932 (O_3932,N_49362,N_47612);
and UO_3933 (O_3933,N_48535,N_49393);
xor UO_3934 (O_3934,N_48384,N_47527);
and UO_3935 (O_3935,N_49526,N_49023);
or UO_3936 (O_3936,N_49282,N_48036);
and UO_3937 (O_3937,N_48489,N_49705);
nand UO_3938 (O_3938,N_47577,N_48571);
nor UO_3939 (O_3939,N_47803,N_48564);
xnor UO_3940 (O_3940,N_47567,N_48033);
nand UO_3941 (O_3941,N_47663,N_48002);
xor UO_3942 (O_3942,N_49886,N_47787);
or UO_3943 (O_3943,N_49232,N_49386);
nor UO_3944 (O_3944,N_49689,N_49157);
or UO_3945 (O_3945,N_48076,N_49065);
xor UO_3946 (O_3946,N_49931,N_48059);
or UO_3947 (O_3947,N_48205,N_47984);
nor UO_3948 (O_3948,N_47895,N_48861);
xor UO_3949 (O_3949,N_49668,N_47566);
nor UO_3950 (O_3950,N_47662,N_47857);
nor UO_3951 (O_3951,N_48933,N_49299);
nor UO_3952 (O_3952,N_48918,N_48319);
or UO_3953 (O_3953,N_47892,N_48690);
nor UO_3954 (O_3954,N_49695,N_48054);
xor UO_3955 (O_3955,N_48384,N_48164);
or UO_3956 (O_3956,N_48762,N_49756);
or UO_3957 (O_3957,N_49475,N_48736);
nand UO_3958 (O_3958,N_48435,N_49024);
nand UO_3959 (O_3959,N_48041,N_48626);
and UO_3960 (O_3960,N_49945,N_48285);
and UO_3961 (O_3961,N_49886,N_49572);
nor UO_3962 (O_3962,N_48179,N_48623);
and UO_3963 (O_3963,N_49442,N_48440);
nor UO_3964 (O_3964,N_47555,N_49138);
nand UO_3965 (O_3965,N_48126,N_48996);
xnor UO_3966 (O_3966,N_49621,N_48852);
xor UO_3967 (O_3967,N_49873,N_47708);
or UO_3968 (O_3968,N_48532,N_48855);
and UO_3969 (O_3969,N_48556,N_47655);
or UO_3970 (O_3970,N_48488,N_49939);
xor UO_3971 (O_3971,N_49135,N_49433);
xor UO_3972 (O_3972,N_49383,N_49340);
nand UO_3973 (O_3973,N_49549,N_49514);
nand UO_3974 (O_3974,N_49839,N_48618);
or UO_3975 (O_3975,N_48503,N_47811);
nand UO_3976 (O_3976,N_47929,N_49609);
nor UO_3977 (O_3977,N_49062,N_49754);
nand UO_3978 (O_3978,N_48340,N_49012);
and UO_3979 (O_3979,N_49724,N_49149);
xor UO_3980 (O_3980,N_47846,N_48983);
nand UO_3981 (O_3981,N_48501,N_48006);
or UO_3982 (O_3982,N_47971,N_49401);
nor UO_3983 (O_3983,N_49101,N_48843);
xnor UO_3984 (O_3984,N_49689,N_48990);
or UO_3985 (O_3985,N_48229,N_49781);
nor UO_3986 (O_3986,N_48684,N_48614);
xor UO_3987 (O_3987,N_47985,N_49928);
nand UO_3988 (O_3988,N_48484,N_48498);
or UO_3989 (O_3989,N_47535,N_48459);
xor UO_3990 (O_3990,N_49377,N_48569);
nor UO_3991 (O_3991,N_49391,N_47604);
xor UO_3992 (O_3992,N_47573,N_47677);
xor UO_3993 (O_3993,N_47890,N_49041);
xnor UO_3994 (O_3994,N_47867,N_48222);
nor UO_3995 (O_3995,N_49402,N_48322);
nand UO_3996 (O_3996,N_48657,N_48848);
and UO_3997 (O_3997,N_48466,N_47930);
and UO_3998 (O_3998,N_48973,N_49516);
and UO_3999 (O_3999,N_47634,N_47775);
nor UO_4000 (O_4000,N_48565,N_49017);
or UO_4001 (O_4001,N_48550,N_49546);
and UO_4002 (O_4002,N_48878,N_48721);
nand UO_4003 (O_4003,N_47592,N_49705);
nor UO_4004 (O_4004,N_48158,N_48971);
xor UO_4005 (O_4005,N_48059,N_49731);
xor UO_4006 (O_4006,N_47570,N_48168);
or UO_4007 (O_4007,N_47711,N_47551);
nand UO_4008 (O_4008,N_48187,N_48315);
xnor UO_4009 (O_4009,N_49055,N_49807);
and UO_4010 (O_4010,N_49916,N_49164);
nand UO_4011 (O_4011,N_48524,N_49582);
xnor UO_4012 (O_4012,N_49419,N_49392);
or UO_4013 (O_4013,N_49255,N_47563);
nor UO_4014 (O_4014,N_48004,N_49427);
and UO_4015 (O_4015,N_49322,N_48935);
nand UO_4016 (O_4016,N_48769,N_48678);
nor UO_4017 (O_4017,N_49366,N_48382);
or UO_4018 (O_4018,N_48287,N_49246);
or UO_4019 (O_4019,N_47705,N_48321);
nor UO_4020 (O_4020,N_47628,N_48552);
or UO_4021 (O_4021,N_49341,N_48073);
nand UO_4022 (O_4022,N_49271,N_47911);
or UO_4023 (O_4023,N_47635,N_49124);
and UO_4024 (O_4024,N_48178,N_47862);
nand UO_4025 (O_4025,N_48299,N_48101);
nor UO_4026 (O_4026,N_49596,N_47882);
nand UO_4027 (O_4027,N_48909,N_49621);
or UO_4028 (O_4028,N_48370,N_49311);
or UO_4029 (O_4029,N_49334,N_48607);
nor UO_4030 (O_4030,N_48430,N_49758);
or UO_4031 (O_4031,N_49641,N_48326);
or UO_4032 (O_4032,N_48550,N_49897);
nor UO_4033 (O_4033,N_48116,N_48157);
nand UO_4034 (O_4034,N_49582,N_49847);
xnor UO_4035 (O_4035,N_47516,N_48558);
nand UO_4036 (O_4036,N_48403,N_48609);
nor UO_4037 (O_4037,N_48267,N_49691);
xor UO_4038 (O_4038,N_49140,N_48240);
xor UO_4039 (O_4039,N_48778,N_48134);
xor UO_4040 (O_4040,N_48830,N_48222);
or UO_4041 (O_4041,N_48881,N_49362);
xnor UO_4042 (O_4042,N_48732,N_48856);
nor UO_4043 (O_4043,N_47590,N_48752);
nand UO_4044 (O_4044,N_48723,N_49431);
nor UO_4045 (O_4045,N_48039,N_47799);
or UO_4046 (O_4046,N_48621,N_48867);
nand UO_4047 (O_4047,N_49293,N_49336);
or UO_4048 (O_4048,N_48441,N_47659);
nor UO_4049 (O_4049,N_48813,N_49196);
xnor UO_4050 (O_4050,N_49371,N_49156);
or UO_4051 (O_4051,N_49955,N_48477);
or UO_4052 (O_4052,N_48008,N_49723);
xnor UO_4053 (O_4053,N_49855,N_48914);
or UO_4054 (O_4054,N_49685,N_49816);
xor UO_4055 (O_4055,N_48792,N_48501);
and UO_4056 (O_4056,N_48814,N_47972);
nand UO_4057 (O_4057,N_49643,N_48444);
nor UO_4058 (O_4058,N_48475,N_48847);
and UO_4059 (O_4059,N_48751,N_48914);
nor UO_4060 (O_4060,N_49810,N_48075);
and UO_4061 (O_4061,N_47986,N_49436);
or UO_4062 (O_4062,N_49539,N_49341);
xnor UO_4063 (O_4063,N_49235,N_49933);
xnor UO_4064 (O_4064,N_48633,N_47972);
nand UO_4065 (O_4065,N_48819,N_49920);
or UO_4066 (O_4066,N_49683,N_48527);
nand UO_4067 (O_4067,N_48252,N_49162);
nor UO_4068 (O_4068,N_47816,N_48481);
nor UO_4069 (O_4069,N_49844,N_49043);
xor UO_4070 (O_4070,N_49324,N_48449);
or UO_4071 (O_4071,N_49726,N_48898);
nand UO_4072 (O_4072,N_49754,N_48198);
nor UO_4073 (O_4073,N_48672,N_49557);
nand UO_4074 (O_4074,N_48549,N_47629);
xnor UO_4075 (O_4075,N_48999,N_49849);
nor UO_4076 (O_4076,N_49419,N_47771);
xor UO_4077 (O_4077,N_48075,N_49178);
nand UO_4078 (O_4078,N_49663,N_48361);
nor UO_4079 (O_4079,N_48319,N_47625);
and UO_4080 (O_4080,N_48272,N_49980);
xor UO_4081 (O_4081,N_49738,N_48866);
or UO_4082 (O_4082,N_49530,N_49873);
or UO_4083 (O_4083,N_48067,N_47796);
or UO_4084 (O_4084,N_47558,N_48220);
or UO_4085 (O_4085,N_49470,N_47649);
nor UO_4086 (O_4086,N_48521,N_47913);
nor UO_4087 (O_4087,N_49264,N_49091);
nor UO_4088 (O_4088,N_49478,N_49210);
nor UO_4089 (O_4089,N_49543,N_48877);
xor UO_4090 (O_4090,N_48397,N_48907);
and UO_4091 (O_4091,N_48996,N_49542);
and UO_4092 (O_4092,N_49633,N_48058);
and UO_4093 (O_4093,N_49950,N_49624);
or UO_4094 (O_4094,N_48950,N_47580);
xnor UO_4095 (O_4095,N_48530,N_48146);
or UO_4096 (O_4096,N_48717,N_49338);
xnor UO_4097 (O_4097,N_48945,N_49043);
nand UO_4098 (O_4098,N_48577,N_47823);
and UO_4099 (O_4099,N_48971,N_49924);
nor UO_4100 (O_4100,N_48680,N_49203);
nand UO_4101 (O_4101,N_48436,N_49664);
nor UO_4102 (O_4102,N_49911,N_49965);
nor UO_4103 (O_4103,N_48176,N_48775);
xnor UO_4104 (O_4104,N_48654,N_48974);
nand UO_4105 (O_4105,N_49372,N_49461);
nand UO_4106 (O_4106,N_47819,N_49258);
xor UO_4107 (O_4107,N_47741,N_48533);
nand UO_4108 (O_4108,N_48111,N_48436);
nand UO_4109 (O_4109,N_48752,N_47929);
xnor UO_4110 (O_4110,N_47546,N_47989);
and UO_4111 (O_4111,N_48238,N_49069);
or UO_4112 (O_4112,N_48817,N_48837);
or UO_4113 (O_4113,N_49681,N_49223);
and UO_4114 (O_4114,N_49413,N_49815);
nand UO_4115 (O_4115,N_49187,N_49078);
and UO_4116 (O_4116,N_47987,N_47510);
xor UO_4117 (O_4117,N_49582,N_49179);
and UO_4118 (O_4118,N_47978,N_49001);
or UO_4119 (O_4119,N_47963,N_49568);
or UO_4120 (O_4120,N_48162,N_48173);
nand UO_4121 (O_4121,N_49351,N_48421);
and UO_4122 (O_4122,N_49507,N_48948);
xor UO_4123 (O_4123,N_47698,N_49996);
xnor UO_4124 (O_4124,N_49807,N_48757);
or UO_4125 (O_4125,N_48625,N_49139);
nor UO_4126 (O_4126,N_48766,N_49926);
and UO_4127 (O_4127,N_47796,N_48936);
nand UO_4128 (O_4128,N_47968,N_48205);
xnor UO_4129 (O_4129,N_47537,N_47849);
or UO_4130 (O_4130,N_48542,N_49065);
xnor UO_4131 (O_4131,N_48331,N_49874);
or UO_4132 (O_4132,N_47597,N_47573);
nor UO_4133 (O_4133,N_49278,N_49094);
xnor UO_4134 (O_4134,N_47827,N_47698);
xnor UO_4135 (O_4135,N_49296,N_48757);
and UO_4136 (O_4136,N_48833,N_48132);
or UO_4137 (O_4137,N_48906,N_49177);
nor UO_4138 (O_4138,N_49479,N_47690);
xnor UO_4139 (O_4139,N_49719,N_48800);
nand UO_4140 (O_4140,N_49819,N_48184);
or UO_4141 (O_4141,N_47881,N_48317);
or UO_4142 (O_4142,N_49009,N_47670);
xnor UO_4143 (O_4143,N_48413,N_48806);
or UO_4144 (O_4144,N_49529,N_49204);
nor UO_4145 (O_4145,N_47923,N_47785);
xnor UO_4146 (O_4146,N_47759,N_48939);
and UO_4147 (O_4147,N_48001,N_48989);
nand UO_4148 (O_4148,N_48153,N_47968);
nand UO_4149 (O_4149,N_48686,N_49504);
xnor UO_4150 (O_4150,N_48318,N_48359);
and UO_4151 (O_4151,N_49093,N_49627);
nand UO_4152 (O_4152,N_49155,N_47606);
xnor UO_4153 (O_4153,N_48611,N_49750);
xor UO_4154 (O_4154,N_48336,N_47949);
xor UO_4155 (O_4155,N_48528,N_49372);
or UO_4156 (O_4156,N_49465,N_48591);
and UO_4157 (O_4157,N_48086,N_47659);
nand UO_4158 (O_4158,N_47862,N_47797);
or UO_4159 (O_4159,N_48183,N_49849);
and UO_4160 (O_4160,N_47844,N_48066);
or UO_4161 (O_4161,N_47638,N_48623);
xnor UO_4162 (O_4162,N_47619,N_48004);
or UO_4163 (O_4163,N_49195,N_47873);
and UO_4164 (O_4164,N_49108,N_47847);
or UO_4165 (O_4165,N_48855,N_49109);
xor UO_4166 (O_4166,N_49367,N_48986);
nor UO_4167 (O_4167,N_48586,N_47980);
nor UO_4168 (O_4168,N_48140,N_48381);
or UO_4169 (O_4169,N_48286,N_49342);
xor UO_4170 (O_4170,N_48223,N_49527);
nand UO_4171 (O_4171,N_48293,N_48671);
and UO_4172 (O_4172,N_47687,N_49369);
nor UO_4173 (O_4173,N_47880,N_48890);
nand UO_4174 (O_4174,N_49002,N_48412);
xor UO_4175 (O_4175,N_49727,N_48690);
and UO_4176 (O_4176,N_49707,N_47789);
nand UO_4177 (O_4177,N_47599,N_49860);
and UO_4178 (O_4178,N_49475,N_47853);
nand UO_4179 (O_4179,N_48830,N_48092);
or UO_4180 (O_4180,N_49854,N_47868);
nand UO_4181 (O_4181,N_47836,N_48477);
or UO_4182 (O_4182,N_48721,N_48014);
nor UO_4183 (O_4183,N_48210,N_48122);
xor UO_4184 (O_4184,N_49332,N_48507);
nor UO_4185 (O_4185,N_49442,N_47975);
or UO_4186 (O_4186,N_48901,N_47811);
nand UO_4187 (O_4187,N_47813,N_49044);
xor UO_4188 (O_4188,N_48105,N_48482);
xor UO_4189 (O_4189,N_47509,N_49510);
and UO_4190 (O_4190,N_49420,N_49871);
nand UO_4191 (O_4191,N_48808,N_49114);
and UO_4192 (O_4192,N_48484,N_48058);
nor UO_4193 (O_4193,N_49030,N_49678);
nor UO_4194 (O_4194,N_48077,N_48137);
xnor UO_4195 (O_4195,N_49048,N_47638);
and UO_4196 (O_4196,N_49573,N_48421);
and UO_4197 (O_4197,N_47910,N_49340);
xnor UO_4198 (O_4198,N_48789,N_47904);
or UO_4199 (O_4199,N_49442,N_48897);
nor UO_4200 (O_4200,N_48202,N_47550);
or UO_4201 (O_4201,N_48682,N_48189);
xor UO_4202 (O_4202,N_48035,N_49957);
or UO_4203 (O_4203,N_49999,N_49577);
nor UO_4204 (O_4204,N_48937,N_49308);
or UO_4205 (O_4205,N_49469,N_48670);
and UO_4206 (O_4206,N_48568,N_49447);
and UO_4207 (O_4207,N_48549,N_49910);
nand UO_4208 (O_4208,N_49367,N_48305);
or UO_4209 (O_4209,N_48863,N_49748);
and UO_4210 (O_4210,N_49546,N_49412);
and UO_4211 (O_4211,N_47591,N_49487);
and UO_4212 (O_4212,N_48358,N_49418);
and UO_4213 (O_4213,N_47786,N_49193);
and UO_4214 (O_4214,N_47896,N_49501);
nand UO_4215 (O_4215,N_48746,N_49110);
nor UO_4216 (O_4216,N_49840,N_49914);
xor UO_4217 (O_4217,N_49030,N_47601);
nor UO_4218 (O_4218,N_48941,N_49495);
or UO_4219 (O_4219,N_48986,N_49081);
nor UO_4220 (O_4220,N_47747,N_49387);
xor UO_4221 (O_4221,N_47622,N_47806);
nand UO_4222 (O_4222,N_48774,N_49067);
nand UO_4223 (O_4223,N_49607,N_48469);
or UO_4224 (O_4224,N_47859,N_49828);
xnor UO_4225 (O_4225,N_48955,N_48156);
nand UO_4226 (O_4226,N_49952,N_49607);
xor UO_4227 (O_4227,N_48364,N_49162);
xnor UO_4228 (O_4228,N_47572,N_48511);
nor UO_4229 (O_4229,N_47727,N_48791);
nor UO_4230 (O_4230,N_48710,N_48630);
or UO_4231 (O_4231,N_49923,N_49522);
nor UO_4232 (O_4232,N_49756,N_49207);
and UO_4233 (O_4233,N_49358,N_48284);
nand UO_4234 (O_4234,N_49077,N_48580);
nor UO_4235 (O_4235,N_48190,N_47706);
or UO_4236 (O_4236,N_48971,N_49336);
or UO_4237 (O_4237,N_49722,N_48360);
nor UO_4238 (O_4238,N_49029,N_49336);
and UO_4239 (O_4239,N_49487,N_48033);
and UO_4240 (O_4240,N_47885,N_48272);
xnor UO_4241 (O_4241,N_48465,N_47573);
xnor UO_4242 (O_4242,N_49685,N_48224);
or UO_4243 (O_4243,N_48563,N_48839);
and UO_4244 (O_4244,N_49191,N_47656);
nor UO_4245 (O_4245,N_47731,N_47747);
xor UO_4246 (O_4246,N_48306,N_48845);
nor UO_4247 (O_4247,N_49344,N_49174);
and UO_4248 (O_4248,N_48009,N_48264);
nor UO_4249 (O_4249,N_49126,N_49044);
nand UO_4250 (O_4250,N_49647,N_49886);
xnor UO_4251 (O_4251,N_49624,N_48457);
nand UO_4252 (O_4252,N_49949,N_48884);
xor UO_4253 (O_4253,N_47632,N_48635);
or UO_4254 (O_4254,N_48903,N_48486);
nor UO_4255 (O_4255,N_48416,N_48459);
nor UO_4256 (O_4256,N_49245,N_47794);
or UO_4257 (O_4257,N_47795,N_48198);
nand UO_4258 (O_4258,N_48846,N_49352);
nand UO_4259 (O_4259,N_48007,N_49325);
or UO_4260 (O_4260,N_48597,N_49482);
nand UO_4261 (O_4261,N_48311,N_48607);
xor UO_4262 (O_4262,N_47601,N_48322);
nor UO_4263 (O_4263,N_49827,N_48651);
or UO_4264 (O_4264,N_49901,N_49955);
xor UO_4265 (O_4265,N_48414,N_47843);
or UO_4266 (O_4266,N_48586,N_47788);
and UO_4267 (O_4267,N_49182,N_47710);
nand UO_4268 (O_4268,N_48855,N_48582);
and UO_4269 (O_4269,N_48364,N_47977);
and UO_4270 (O_4270,N_48533,N_49917);
nand UO_4271 (O_4271,N_49454,N_48586);
xor UO_4272 (O_4272,N_49595,N_47652);
nand UO_4273 (O_4273,N_49152,N_49176);
and UO_4274 (O_4274,N_48506,N_48994);
nor UO_4275 (O_4275,N_48533,N_49474);
nor UO_4276 (O_4276,N_49070,N_49466);
and UO_4277 (O_4277,N_49209,N_48169);
or UO_4278 (O_4278,N_49011,N_47912);
nor UO_4279 (O_4279,N_48088,N_49144);
or UO_4280 (O_4280,N_48991,N_48898);
or UO_4281 (O_4281,N_49223,N_49129);
and UO_4282 (O_4282,N_49679,N_48770);
xor UO_4283 (O_4283,N_49024,N_48315);
or UO_4284 (O_4284,N_49923,N_49773);
and UO_4285 (O_4285,N_48468,N_48338);
or UO_4286 (O_4286,N_47672,N_49059);
nand UO_4287 (O_4287,N_47795,N_48318);
and UO_4288 (O_4288,N_49792,N_49528);
xnor UO_4289 (O_4289,N_49571,N_49520);
nor UO_4290 (O_4290,N_48283,N_47951);
nand UO_4291 (O_4291,N_49165,N_48969);
nand UO_4292 (O_4292,N_49381,N_48598);
and UO_4293 (O_4293,N_48929,N_47630);
and UO_4294 (O_4294,N_48092,N_49773);
xnor UO_4295 (O_4295,N_47580,N_49439);
nand UO_4296 (O_4296,N_48604,N_47769);
nor UO_4297 (O_4297,N_49563,N_47511);
xor UO_4298 (O_4298,N_48194,N_49389);
xnor UO_4299 (O_4299,N_49370,N_49161);
nand UO_4300 (O_4300,N_48425,N_49109);
xor UO_4301 (O_4301,N_48150,N_47719);
xnor UO_4302 (O_4302,N_47734,N_47639);
nand UO_4303 (O_4303,N_49917,N_49352);
or UO_4304 (O_4304,N_48636,N_48471);
xnor UO_4305 (O_4305,N_48480,N_49850);
and UO_4306 (O_4306,N_47721,N_49111);
xor UO_4307 (O_4307,N_47501,N_47745);
nand UO_4308 (O_4308,N_49651,N_47822);
and UO_4309 (O_4309,N_49720,N_47967);
and UO_4310 (O_4310,N_47789,N_48396);
nor UO_4311 (O_4311,N_49089,N_48543);
nand UO_4312 (O_4312,N_49760,N_48738);
nor UO_4313 (O_4313,N_47933,N_47984);
nand UO_4314 (O_4314,N_49770,N_49829);
nor UO_4315 (O_4315,N_47888,N_49219);
nor UO_4316 (O_4316,N_49458,N_49091);
xor UO_4317 (O_4317,N_48633,N_47620);
nand UO_4318 (O_4318,N_48134,N_49140);
nor UO_4319 (O_4319,N_48559,N_47760);
nor UO_4320 (O_4320,N_48977,N_48107);
nand UO_4321 (O_4321,N_48884,N_49940);
nand UO_4322 (O_4322,N_49746,N_48832);
and UO_4323 (O_4323,N_49884,N_49233);
xnor UO_4324 (O_4324,N_48439,N_48990);
or UO_4325 (O_4325,N_49687,N_49440);
xor UO_4326 (O_4326,N_49124,N_47546);
xor UO_4327 (O_4327,N_49757,N_49375);
xnor UO_4328 (O_4328,N_49195,N_49864);
or UO_4329 (O_4329,N_48863,N_47522);
nor UO_4330 (O_4330,N_47964,N_49369);
nor UO_4331 (O_4331,N_48316,N_49776);
and UO_4332 (O_4332,N_49459,N_48300);
or UO_4333 (O_4333,N_49480,N_47786);
and UO_4334 (O_4334,N_47618,N_49445);
xor UO_4335 (O_4335,N_48020,N_47692);
xor UO_4336 (O_4336,N_49809,N_49656);
xnor UO_4337 (O_4337,N_47711,N_47957);
xnor UO_4338 (O_4338,N_48313,N_49670);
or UO_4339 (O_4339,N_48065,N_49223);
nor UO_4340 (O_4340,N_49984,N_49826);
nor UO_4341 (O_4341,N_49369,N_49231);
xnor UO_4342 (O_4342,N_48514,N_49786);
nand UO_4343 (O_4343,N_49200,N_49758);
xor UO_4344 (O_4344,N_47544,N_49221);
or UO_4345 (O_4345,N_49301,N_49562);
nand UO_4346 (O_4346,N_49175,N_48414);
and UO_4347 (O_4347,N_48044,N_48379);
nand UO_4348 (O_4348,N_47646,N_49440);
nor UO_4349 (O_4349,N_48658,N_48862);
xor UO_4350 (O_4350,N_48757,N_47717);
or UO_4351 (O_4351,N_48754,N_48193);
or UO_4352 (O_4352,N_48333,N_49208);
and UO_4353 (O_4353,N_49485,N_49636);
xnor UO_4354 (O_4354,N_48844,N_49869);
nor UO_4355 (O_4355,N_47931,N_49676);
and UO_4356 (O_4356,N_48208,N_48412);
and UO_4357 (O_4357,N_48823,N_49802);
nor UO_4358 (O_4358,N_49053,N_48450);
or UO_4359 (O_4359,N_49551,N_48046);
or UO_4360 (O_4360,N_47583,N_48535);
or UO_4361 (O_4361,N_49943,N_49978);
nand UO_4362 (O_4362,N_49240,N_49553);
nor UO_4363 (O_4363,N_49983,N_49206);
and UO_4364 (O_4364,N_48721,N_48195);
and UO_4365 (O_4365,N_48829,N_47705);
and UO_4366 (O_4366,N_48726,N_49385);
and UO_4367 (O_4367,N_49580,N_49505);
nor UO_4368 (O_4368,N_49586,N_48832);
and UO_4369 (O_4369,N_48357,N_48403);
xnor UO_4370 (O_4370,N_49934,N_49593);
xnor UO_4371 (O_4371,N_48389,N_48538);
nand UO_4372 (O_4372,N_48135,N_49406);
nor UO_4373 (O_4373,N_49239,N_49101);
xnor UO_4374 (O_4374,N_47525,N_49277);
nand UO_4375 (O_4375,N_48718,N_47748);
nor UO_4376 (O_4376,N_47703,N_48350);
nand UO_4377 (O_4377,N_49809,N_48460);
nand UO_4378 (O_4378,N_48058,N_47914);
and UO_4379 (O_4379,N_47503,N_48095);
and UO_4380 (O_4380,N_47767,N_48554);
nor UO_4381 (O_4381,N_48343,N_49442);
and UO_4382 (O_4382,N_49319,N_48245);
nand UO_4383 (O_4383,N_49908,N_48381);
or UO_4384 (O_4384,N_47972,N_48541);
nor UO_4385 (O_4385,N_48779,N_49853);
or UO_4386 (O_4386,N_48376,N_47791);
and UO_4387 (O_4387,N_49317,N_48216);
or UO_4388 (O_4388,N_49805,N_49759);
and UO_4389 (O_4389,N_48273,N_49330);
nand UO_4390 (O_4390,N_48878,N_49119);
nor UO_4391 (O_4391,N_49450,N_48398);
nor UO_4392 (O_4392,N_48907,N_49383);
nand UO_4393 (O_4393,N_47528,N_47504);
nor UO_4394 (O_4394,N_49132,N_47796);
nand UO_4395 (O_4395,N_47653,N_49416);
nor UO_4396 (O_4396,N_49680,N_48922);
or UO_4397 (O_4397,N_48060,N_48623);
nor UO_4398 (O_4398,N_49775,N_47665);
or UO_4399 (O_4399,N_49809,N_49356);
nand UO_4400 (O_4400,N_49747,N_47865);
nand UO_4401 (O_4401,N_49913,N_49590);
nand UO_4402 (O_4402,N_49621,N_49857);
xor UO_4403 (O_4403,N_49794,N_49777);
or UO_4404 (O_4404,N_47616,N_49312);
nor UO_4405 (O_4405,N_49848,N_47998);
nor UO_4406 (O_4406,N_48962,N_48318);
and UO_4407 (O_4407,N_49308,N_48405);
nor UO_4408 (O_4408,N_49897,N_49347);
xor UO_4409 (O_4409,N_49513,N_48881);
xnor UO_4410 (O_4410,N_49447,N_49551);
nand UO_4411 (O_4411,N_48554,N_47577);
and UO_4412 (O_4412,N_47777,N_48895);
nor UO_4413 (O_4413,N_49426,N_49113);
nor UO_4414 (O_4414,N_47995,N_48165);
nand UO_4415 (O_4415,N_48502,N_49042);
xnor UO_4416 (O_4416,N_49282,N_48143);
or UO_4417 (O_4417,N_48840,N_49192);
and UO_4418 (O_4418,N_48658,N_49304);
and UO_4419 (O_4419,N_48609,N_48045);
and UO_4420 (O_4420,N_49068,N_47906);
nor UO_4421 (O_4421,N_48377,N_48022);
and UO_4422 (O_4422,N_49286,N_49678);
xor UO_4423 (O_4423,N_48608,N_49304);
xor UO_4424 (O_4424,N_48554,N_47750);
nand UO_4425 (O_4425,N_48987,N_48532);
or UO_4426 (O_4426,N_49956,N_49394);
and UO_4427 (O_4427,N_49980,N_48354);
nor UO_4428 (O_4428,N_48825,N_48324);
xor UO_4429 (O_4429,N_47966,N_49425);
nand UO_4430 (O_4430,N_47975,N_48810);
xnor UO_4431 (O_4431,N_49331,N_47745);
nor UO_4432 (O_4432,N_48896,N_49747);
xor UO_4433 (O_4433,N_47515,N_49158);
and UO_4434 (O_4434,N_48985,N_49035);
nand UO_4435 (O_4435,N_48331,N_48894);
nor UO_4436 (O_4436,N_47652,N_47918);
nand UO_4437 (O_4437,N_47610,N_48593);
and UO_4438 (O_4438,N_49039,N_49997);
or UO_4439 (O_4439,N_47775,N_48098);
or UO_4440 (O_4440,N_47530,N_47528);
nor UO_4441 (O_4441,N_48873,N_49659);
nand UO_4442 (O_4442,N_49892,N_48048);
xor UO_4443 (O_4443,N_48303,N_48713);
and UO_4444 (O_4444,N_47828,N_49872);
and UO_4445 (O_4445,N_49813,N_49587);
or UO_4446 (O_4446,N_49163,N_48408);
xnor UO_4447 (O_4447,N_48904,N_49005);
or UO_4448 (O_4448,N_49602,N_48804);
nor UO_4449 (O_4449,N_49582,N_48151);
or UO_4450 (O_4450,N_47970,N_49806);
nand UO_4451 (O_4451,N_48273,N_49918);
nor UO_4452 (O_4452,N_48759,N_49934);
or UO_4453 (O_4453,N_49372,N_48115);
xor UO_4454 (O_4454,N_49879,N_49804);
or UO_4455 (O_4455,N_49941,N_48293);
and UO_4456 (O_4456,N_48625,N_49167);
and UO_4457 (O_4457,N_48989,N_49008);
or UO_4458 (O_4458,N_49229,N_48362);
or UO_4459 (O_4459,N_49766,N_48251);
and UO_4460 (O_4460,N_47666,N_48119);
xor UO_4461 (O_4461,N_48825,N_47836);
nor UO_4462 (O_4462,N_47996,N_49424);
and UO_4463 (O_4463,N_49325,N_48134);
and UO_4464 (O_4464,N_48045,N_47502);
nand UO_4465 (O_4465,N_48707,N_48028);
or UO_4466 (O_4466,N_49355,N_47928);
nor UO_4467 (O_4467,N_49884,N_49926);
xor UO_4468 (O_4468,N_48415,N_49773);
or UO_4469 (O_4469,N_47541,N_47735);
and UO_4470 (O_4470,N_48631,N_47513);
nor UO_4471 (O_4471,N_48820,N_48973);
nor UO_4472 (O_4472,N_49404,N_48262);
nand UO_4473 (O_4473,N_47516,N_48753);
or UO_4474 (O_4474,N_48247,N_49183);
nor UO_4475 (O_4475,N_49865,N_48142);
nor UO_4476 (O_4476,N_47848,N_47524);
or UO_4477 (O_4477,N_49247,N_49378);
xnor UO_4478 (O_4478,N_49845,N_49519);
and UO_4479 (O_4479,N_48285,N_48423);
nand UO_4480 (O_4480,N_47798,N_48768);
xor UO_4481 (O_4481,N_49282,N_47618);
and UO_4482 (O_4482,N_47515,N_47526);
nand UO_4483 (O_4483,N_49967,N_49094);
or UO_4484 (O_4484,N_48615,N_47759);
and UO_4485 (O_4485,N_48554,N_49014);
or UO_4486 (O_4486,N_47884,N_48418);
xor UO_4487 (O_4487,N_48653,N_49946);
and UO_4488 (O_4488,N_49885,N_49265);
or UO_4489 (O_4489,N_49328,N_49865);
nand UO_4490 (O_4490,N_48562,N_49606);
xor UO_4491 (O_4491,N_48325,N_49114);
or UO_4492 (O_4492,N_49103,N_49351);
nor UO_4493 (O_4493,N_49788,N_48250);
nor UO_4494 (O_4494,N_48118,N_49536);
xnor UO_4495 (O_4495,N_49522,N_48186);
and UO_4496 (O_4496,N_47892,N_48531);
nand UO_4497 (O_4497,N_49703,N_48908);
and UO_4498 (O_4498,N_48901,N_48974);
and UO_4499 (O_4499,N_49497,N_49099);
nor UO_4500 (O_4500,N_48482,N_48658);
or UO_4501 (O_4501,N_49475,N_48688);
and UO_4502 (O_4502,N_48048,N_49331);
or UO_4503 (O_4503,N_48855,N_49134);
or UO_4504 (O_4504,N_49893,N_48203);
nor UO_4505 (O_4505,N_49479,N_47599);
or UO_4506 (O_4506,N_47948,N_47738);
nand UO_4507 (O_4507,N_48965,N_49595);
nor UO_4508 (O_4508,N_47949,N_48632);
xnor UO_4509 (O_4509,N_47994,N_49225);
or UO_4510 (O_4510,N_49727,N_48240);
or UO_4511 (O_4511,N_48036,N_49038);
nand UO_4512 (O_4512,N_48396,N_47952);
or UO_4513 (O_4513,N_49282,N_47999);
nor UO_4514 (O_4514,N_48609,N_47642);
or UO_4515 (O_4515,N_48902,N_48273);
xor UO_4516 (O_4516,N_47835,N_47729);
xor UO_4517 (O_4517,N_49055,N_48321);
nor UO_4518 (O_4518,N_49557,N_49040);
and UO_4519 (O_4519,N_49660,N_47763);
and UO_4520 (O_4520,N_49395,N_48531);
xor UO_4521 (O_4521,N_48127,N_47813);
nor UO_4522 (O_4522,N_48330,N_48840);
xor UO_4523 (O_4523,N_48917,N_48476);
or UO_4524 (O_4524,N_49096,N_48925);
xor UO_4525 (O_4525,N_48063,N_47799);
and UO_4526 (O_4526,N_49766,N_48643);
xor UO_4527 (O_4527,N_49889,N_47948);
nor UO_4528 (O_4528,N_48777,N_48573);
nand UO_4529 (O_4529,N_48911,N_49402);
nand UO_4530 (O_4530,N_49183,N_48274);
xnor UO_4531 (O_4531,N_49090,N_48456);
nor UO_4532 (O_4532,N_49590,N_49002);
xnor UO_4533 (O_4533,N_49793,N_47904);
or UO_4534 (O_4534,N_47845,N_48216);
nor UO_4535 (O_4535,N_47629,N_48565);
nor UO_4536 (O_4536,N_48764,N_48772);
nor UO_4537 (O_4537,N_47661,N_49887);
xor UO_4538 (O_4538,N_48342,N_47936);
or UO_4539 (O_4539,N_49749,N_48003);
or UO_4540 (O_4540,N_48535,N_48524);
nor UO_4541 (O_4541,N_48743,N_48849);
xnor UO_4542 (O_4542,N_47874,N_47893);
nand UO_4543 (O_4543,N_47848,N_48915);
nand UO_4544 (O_4544,N_49613,N_49443);
nor UO_4545 (O_4545,N_47972,N_47585);
nor UO_4546 (O_4546,N_47937,N_49407);
or UO_4547 (O_4547,N_48056,N_48446);
and UO_4548 (O_4548,N_49825,N_48456);
and UO_4549 (O_4549,N_48122,N_48568);
nand UO_4550 (O_4550,N_48766,N_47611);
nand UO_4551 (O_4551,N_47556,N_49443);
or UO_4552 (O_4552,N_48489,N_49455);
and UO_4553 (O_4553,N_47635,N_48694);
nand UO_4554 (O_4554,N_49607,N_48247);
and UO_4555 (O_4555,N_48050,N_49040);
or UO_4556 (O_4556,N_49133,N_48133);
nand UO_4557 (O_4557,N_49107,N_49683);
and UO_4558 (O_4558,N_47528,N_48003);
xor UO_4559 (O_4559,N_48249,N_48727);
nand UO_4560 (O_4560,N_49486,N_47938);
or UO_4561 (O_4561,N_48293,N_48595);
or UO_4562 (O_4562,N_47834,N_48108);
xor UO_4563 (O_4563,N_48074,N_49443);
or UO_4564 (O_4564,N_49625,N_47984);
xnor UO_4565 (O_4565,N_48129,N_48320);
or UO_4566 (O_4566,N_49600,N_48908);
xor UO_4567 (O_4567,N_47686,N_48073);
nand UO_4568 (O_4568,N_48026,N_49058);
or UO_4569 (O_4569,N_47586,N_49928);
xor UO_4570 (O_4570,N_49524,N_47895);
nor UO_4571 (O_4571,N_48143,N_48155);
nor UO_4572 (O_4572,N_47759,N_49235);
or UO_4573 (O_4573,N_49565,N_47863);
or UO_4574 (O_4574,N_49965,N_49281);
xnor UO_4575 (O_4575,N_49249,N_49696);
nand UO_4576 (O_4576,N_49993,N_49988);
or UO_4577 (O_4577,N_49190,N_49794);
nor UO_4578 (O_4578,N_49982,N_48318);
xnor UO_4579 (O_4579,N_48173,N_47976);
nand UO_4580 (O_4580,N_49263,N_49043);
xor UO_4581 (O_4581,N_47843,N_48653);
or UO_4582 (O_4582,N_49812,N_48170);
nand UO_4583 (O_4583,N_47562,N_48340);
nand UO_4584 (O_4584,N_49578,N_48792);
nand UO_4585 (O_4585,N_49156,N_49738);
nand UO_4586 (O_4586,N_48656,N_48919);
nor UO_4587 (O_4587,N_47973,N_47540);
or UO_4588 (O_4588,N_47711,N_48027);
nand UO_4589 (O_4589,N_48008,N_48059);
xor UO_4590 (O_4590,N_49838,N_48087);
or UO_4591 (O_4591,N_48484,N_47713);
nand UO_4592 (O_4592,N_48385,N_48774);
xnor UO_4593 (O_4593,N_48595,N_48603);
nand UO_4594 (O_4594,N_48455,N_47715);
or UO_4595 (O_4595,N_48713,N_49783);
xor UO_4596 (O_4596,N_48684,N_49990);
or UO_4597 (O_4597,N_49676,N_48591);
nand UO_4598 (O_4598,N_49212,N_48363);
nand UO_4599 (O_4599,N_49756,N_47574);
or UO_4600 (O_4600,N_49305,N_48472);
or UO_4601 (O_4601,N_49004,N_48478);
nand UO_4602 (O_4602,N_48849,N_48087);
nand UO_4603 (O_4603,N_49789,N_49268);
nor UO_4604 (O_4604,N_49377,N_49192);
nand UO_4605 (O_4605,N_48421,N_49886);
xor UO_4606 (O_4606,N_47800,N_49176);
nor UO_4607 (O_4607,N_48390,N_47534);
nand UO_4608 (O_4608,N_47549,N_48567);
or UO_4609 (O_4609,N_49861,N_48123);
nand UO_4610 (O_4610,N_47697,N_49392);
nand UO_4611 (O_4611,N_47781,N_48406);
nor UO_4612 (O_4612,N_47770,N_48865);
and UO_4613 (O_4613,N_47538,N_48952);
or UO_4614 (O_4614,N_49551,N_48185);
nor UO_4615 (O_4615,N_49872,N_49288);
or UO_4616 (O_4616,N_49959,N_47514);
nor UO_4617 (O_4617,N_48497,N_48296);
xnor UO_4618 (O_4618,N_48293,N_49029);
nor UO_4619 (O_4619,N_49541,N_48823);
nand UO_4620 (O_4620,N_49392,N_49420);
and UO_4621 (O_4621,N_49087,N_48400);
nor UO_4622 (O_4622,N_47540,N_48329);
or UO_4623 (O_4623,N_49926,N_48150);
nor UO_4624 (O_4624,N_48856,N_48458);
xnor UO_4625 (O_4625,N_48021,N_48192);
or UO_4626 (O_4626,N_48432,N_48076);
or UO_4627 (O_4627,N_48962,N_48686);
and UO_4628 (O_4628,N_48435,N_48118);
nor UO_4629 (O_4629,N_49640,N_49926);
nand UO_4630 (O_4630,N_49049,N_49275);
nor UO_4631 (O_4631,N_49636,N_47937);
or UO_4632 (O_4632,N_48848,N_49165);
and UO_4633 (O_4633,N_49426,N_48704);
nand UO_4634 (O_4634,N_49816,N_48973);
nor UO_4635 (O_4635,N_48298,N_48222);
xnor UO_4636 (O_4636,N_49875,N_48522);
xor UO_4637 (O_4637,N_47650,N_49042);
nand UO_4638 (O_4638,N_49433,N_49305);
nor UO_4639 (O_4639,N_48038,N_48927);
nand UO_4640 (O_4640,N_49410,N_48639);
or UO_4641 (O_4641,N_49830,N_47784);
xor UO_4642 (O_4642,N_48443,N_48614);
and UO_4643 (O_4643,N_49160,N_47784);
nand UO_4644 (O_4644,N_47706,N_47756);
xnor UO_4645 (O_4645,N_49033,N_49740);
xnor UO_4646 (O_4646,N_48838,N_48522);
or UO_4647 (O_4647,N_47573,N_48820);
xnor UO_4648 (O_4648,N_47935,N_48917);
xnor UO_4649 (O_4649,N_48442,N_47566);
or UO_4650 (O_4650,N_48810,N_47837);
nand UO_4651 (O_4651,N_49735,N_47787);
or UO_4652 (O_4652,N_48935,N_48265);
xor UO_4653 (O_4653,N_47845,N_49035);
nor UO_4654 (O_4654,N_49850,N_47511);
xnor UO_4655 (O_4655,N_48301,N_49757);
nor UO_4656 (O_4656,N_49799,N_47591);
nand UO_4657 (O_4657,N_47968,N_48009);
and UO_4658 (O_4658,N_48523,N_47607);
or UO_4659 (O_4659,N_48535,N_48907);
nor UO_4660 (O_4660,N_47866,N_48403);
nor UO_4661 (O_4661,N_49731,N_49461);
nor UO_4662 (O_4662,N_49636,N_48221);
nor UO_4663 (O_4663,N_48095,N_49150);
nor UO_4664 (O_4664,N_47630,N_49627);
xnor UO_4665 (O_4665,N_49671,N_49522);
nand UO_4666 (O_4666,N_49551,N_48496);
or UO_4667 (O_4667,N_48944,N_49980);
or UO_4668 (O_4668,N_49184,N_48189);
or UO_4669 (O_4669,N_49423,N_48517);
or UO_4670 (O_4670,N_49637,N_48033);
and UO_4671 (O_4671,N_48531,N_47815);
xor UO_4672 (O_4672,N_49533,N_49264);
nand UO_4673 (O_4673,N_48814,N_49190);
nand UO_4674 (O_4674,N_49617,N_48644);
nor UO_4675 (O_4675,N_47970,N_48265);
nand UO_4676 (O_4676,N_49736,N_49602);
nand UO_4677 (O_4677,N_48491,N_49747);
or UO_4678 (O_4678,N_47777,N_48060);
nor UO_4679 (O_4679,N_47822,N_49285);
nand UO_4680 (O_4680,N_48864,N_49350);
or UO_4681 (O_4681,N_48290,N_47650);
nor UO_4682 (O_4682,N_49863,N_49066);
or UO_4683 (O_4683,N_48538,N_47695);
or UO_4684 (O_4684,N_48718,N_47930);
or UO_4685 (O_4685,N_48693,N_47725);
and UO_4686 (O_4686,N_47611,N_49400);
nand UO_4687 (O_4687,N_49440,N_48458);
xnor UO_4688 (O_4688,N_47637,N_48557);
xor UO_4689 (O_4689,N_49164,N_47541);
nor UO_4690 (O_4690,N_49889,N_49267);
or UO_4691 (O_4691,N_47778,N_48181);
xnor UO_4692 (O_4692,N_48419,N_48093);
or UO_4693 (O_4693,N_47876,N_47792);
nand UO_4694 (O_4694,N_47681,N_48133);
nor UO_4695 (O_4695,N_47695,N_48899);
nor UO_4696 (O_4696,N_47790,N_49262);
and UO_4697 (O_4697,N_48695,N_48446);
or UO_4698 (O_4698,N_48676,N_48419);
and UO_4699 (O_4699,N_48556,N_49502);
or UO_4700 (O_4700,N_48883,N_47794);
nor UO_4701 (O_4701,N_48803,N_48428);
or UO_4702 (O_4702,N_49981,N_48024);
xor UO_4703 (O_4703,N_49354,N_48741);
nor UO_4704 (O_4704,N_49026,N_49864);
or UO_4705 (O_4705,N_49321,N_49906);
or UO_4706 (O_4706,N_49610,N_49278);
and UO_4707 (O_4707,N_48901,N_48031);
and UO_4708 (O_4708,N_47706,N_48259);
xor UO_4709 (O_4709,N_49244,N_47544);
nor UO_4710 (O_4710,N_49987,N_48071);
or UO_4711 (O_4711,N_49233,N_48559);
xnor UO_4712 (O_4712,N_49528,N_47779);
nand UO_4713 (O_4713,N_47992,N_49310);
or UO_4714 (O_4714,N_48443,N_48276);
and UO_4715 (O_4715,N_49283,N_49131);
nand UO_4716 (O_4716,N_49048,N_48125);
or UO_4717 (O_4717,N_47799,N_47692);
or UO_4718 (O_4718,N_49590,N_48840);
xor UO_4719 (O_4719,N_48831,N_49638);
or UO_4720 (O_4720,N_48404,N_49390);
and UO_4721 (O_4721,N_48793,N_47669);
nand UO_4722 (O_4722,N_48195,N_47694);
or UO_4723 (O_4723,N_49857,N_48345);
nor UO_4724 (O_4724,N_49043,N_49287);
or UO_4725 (O_4725,N_48203,N_47824);
nor UO_4726 (O_4726,N_49258,N_48668);
xor UO_4727 (O_4727,N_49909,N_48594);
nand UO_4728 (O_4728,N_49367,N_49865);
or UO_4729 (O_4729,N_48026,N_48139);
or UO_4730 (O_4730,N_48148,N_48340);
xnor UO_4731 (O_4731,N_48921,N_47904);
or UO_4732 (O_4732,N_48586,N_48681);
and UO_4733 (O_4733,N_48877,N_47715);
nand UO_4734 (O_4734,N_49556,N_49498);
xor UO_4735 (O_4735,N_48563,N_49914);
nor UO_4736 (O_4736,N_48349,N_47786);
or UO_4737 (O_4737,N_48502,N_49968);
or UO_4738 (O_4738,N_48292,N_49068);
nor UO_4739 (O_4739,N_49381,N_48955);
nand UO_4740 (O_4740,N_48373,N_48830);
and UO_4741 (O_4741,N_49092,N_48522);
or UO_4742 (O_4742,N_48948,N_49535);
and UO_4743 (O_4743,N_49408,N_48535);
nand UO_4744 (O_4744,N_49402,N_48263);
nand UO_4745 (O_4745,N_49880,N_48758);
and UO_4746 (O_4746,N_48852,N_47501);
or UO_4747 (O_4747,N_49001,N_48031);
xnor UO_4748 (O_4748,N_48147,N_48552);
nand UO_4749 (O_4749,N_47665,N_48230);
and UO_4750 (O_4750,N_48947,N_49516);
nand UO_4751 (O_4751,N_48756,N_49741);
nor UO_4752 (O_4752,N_49073,N_48300);
or UO_4753 (O_4753,N_48114,N_48477);
or UO_4754 (O_4754,N_48232,N_48011);
nor UO_4755 (O_4755,N_48448,N_48709);
and UO_4756 (O_4756,N_49834,N_48401);
xnor UO_4757 (O_4757,N_48023,N_47640);
xor UO_4758 (O_4758,N_49405,N_48238);
nor UO_4759 (O_4759,N_49415,N_48212);
xor UO_4760 (O_4760,N_47916,N_49225);
nor UO_4761 (O_4761,N_48856,N_48066);
nand UO_4762 (O_4762,N_49335,N_49770);
nor UO_4763 (O_4763,N_49332,N_49581);
nand UO_4764 (O_4764,N_49349,N_48554);
and UO_4765 (O_4765,N_48136,N_48571);
nand UO_4766 (O_4766,N_47965,N_47755);
and UO_4767 (O_4767,N_49584,N_48812);
or UO_4768 (O_4768,N_48460,N_48217);
or UO_4769 (O_4769,N_49074,N_47938);
or UO_4770 (O_4770,N_49170,N_49513);
or UO_4771 (O_4771,N_48043,N_49232);
xnor UO_4772 (O_4772,N_48553,N_49774);
nor UO_4773 (O_4773,N_49487,N_49050);
xor UO_4774 (O_4774,N_48109,N_49651);
nor UO_4775 (O_4775,N_49824,N_49669);
xor UO_4776 (O_4776,N_49498,N_49427);
nand UO_4777 (O_4777,N_49356,N_47587);
and UO_4778 (O_4778,N_49997,N_47889);
or UO_4779 (O_4779,N_48159,N_49648);
or UO_4780 (O_4780,N_48913,N_49354);
and UO_4781 (O_4781,N_49989,N_47728);
and UO_4782 (O_4782,N_49163,N_47824);
nand UO_4783 (O_4783,N_49215,N_49734);
and UO_4784 (O_4784,N_48755,N_48691);
xnor UO_4785 (O_4785,N_48818,N_49216);
nor UO_4786 (O_4786,N_48203,N_48376);
or UO_4787 (O_4787,N_48928,N_49553);
or UO_4788 (O_4788,N_48488,N_47942);
and UO_4789 (O_4789,N_49272,N_48954);
nand UO_4790 (O_4790,N_47743,N_49976);
or UO_4791 (O_4791,N_47724,N_48469);
or UO_4792 (O_4792,N_47522,N_47572);
and UO_4793 (O_4793,N_48943,N_49908);
nand UO_4794 (O_4794,N_48055,N_49888);
and UO_4795 (O_4795,N_48156,N_49763);
and UO_4796 (O_4796,N_48615,N_48438);
xor UO_4797 (O_4797,N_49846,N_49617);
and UO_4798 (O_4798,N_49577,N_49833);
and UO_4799 (O_4799,N_49176,N_49029);
nand UO_4800 (O_4800,N_48155,N_48978);
nor UO_4801 (O_4801,N_49094,N_49128);
or UO_4802 (O_4802,N_48272,N_49282);
or UO_4803 (O_4803,N_48802,N_48151);
and UO_4804 (O_4804,N_47810,N_48197);
or UO_4805 (O_4805,N_48458,N_48807);
nor UO_4806 (O_4806,N_49106,N_48557);
or UO_4807 (O_4807,N_47652,N_49677);
nor UO_4808 (O_4808,N_49716,N_47538);
xor UO_4809 (O_4809,N_48608,N_48540);
and UO_4810 (O_4810,N_49718,N_48777);
and UO_4811 (O_4811,N_48401,N_48301);
or UO_4812 (O_4812,N_48985,N_49164);
nand UO_4813 (O_4813,N_48011,N_49120);
or UO_4814 (O_4814,N_47982,N_48073);
or UO_4815 (O_4815,N_49312,N_48642);
nor UO_4816 (O_4816,N_49047,N_48263);
or UO_4817 (O_4817,N_49972,N_49028);
nor UO_4818 (O_4818,N_48080,N_48296);
xor UO_4819 (O_4819,N_49425,N_49172);
nand UO_4820 (O_4820,N_47634,N_48115);
nor UO_4821 (O_4821,N_49923,N_49741);
nand UO_4822 (O_4822,N_49832,N_49992);
nand UO_4823 (O_4823,N_48038,N_47870);
nor UO_4824 (O_4824,N_47539,N_49423);
or UO_4825 (O_4825,N_47755,N_48052);
or UO_4826 (O_4826,N_47570,N_49924);
or UO_4827 (O_4827,N_48703,N_49547);
nor UO_4828 (O_4828,N_49167,N_49052);
xor UO_4829 (O_4829,N_49043,N_49473);
xor UO_4830 (O_4830,N_49172,N_47636);
nor UO_4831 (O_4831,N_48177,N_48599);
nor UO_4832 (O_4832,N_49004,N_49141);
nand UO_4833 (O_4833,N_47857,N_49034);
nor UO_4834 (O_4834,N_47778,N_47654);
nor UO_4835 (O_4835,N_48436,N_47800);
xnor UO_4836 (O_4836,N_48327,N_47547);
or UO_4837 (O_4837,N_49010,N_48461);
nor UO_4838 (O_4838,N_48262,N_47517);
xnor UO_4839 (O_4839,N_47747,N_49831);
xor UO_4840 (O_4840,N_49800,N_49445);
nor UO_4841 (O_4841,N_48497,N_49599);
nand UO_4842 (O_4842,N_47856,N_47946);
nand UO_4843 (O_4843,N_47866,N_49356);
and UO_4844 (O_4844,N_49844,N_49926);
and UO_4845 (O_4845,N_48206,N_47548);
nand UO_4846 (O_4846,N_49893,N_47569);
xor UO_4847 (O_4847,N_48987,N_47583);
nand UO_4848 (O_4848,N_49252,N_48983);
xnor UO_4849 (O_4849,N_49073,N_49976);
xnor UO_4850 (O_4850,N_49180,N_49371);
or UO_4851 (O_4851,N_49639,N_49390);
xor UO_4852 (O_4852,N_49951,N_48205);
xnor UO_4853 (O_4853,N_49716,N_48566);
xnor UO_4854 (O_4854,N_48600,N_49531);
nand UO_4855 (O_4855,N_49554,N_47941);
nand UO_4856 (O_4856,N_48093,N_47636);
or UO_4857 (O_4857,N_48274,N_48803);
nor UO_4858 (O_4858,N_48790,N_49982);
nor UO_4859 (O_4859,N_49484,N_49447);
or UO_4860 (O_4860,N_49471,N_48091);
xor UO_4861 (O_4861,N_47722,N_49081);
and UO_4862 (O_4862,N_49369,N_47753);
nand UO_4863 (O_4863,N_49238,N_48501);
or UO_4864 (O_4864,N_48726,N_49105);
and UO_4865 (O_4865,N_48571,N_48896);
and UO_4866 (O_4866,N_48412,N_47532);
and UO_4867 (O_4867,N_47510,N_48729);
and UO_4868 (O_4868,N_48044,N_49619);
xnor UO_4869 (O_4869,N_48141,N_49441);
nor UO_4870 (O_4870,N_48431,N_48187);
and UO_4871 (O_4871,N_48620,N_47879);
and UO_4872 (O_4872,N_49057,N_48352);
nor UO_4873 (O_4873,N_48291,N_48874);
and UO_4874 (O_4874,N_48146,N_49059);
or UO_4875 (O_4875,N_47956,N_47852);
or UO_4876 (O_4876,N_49889,N_48858);
nor UO_4877 (O_4877,N_48074,N_48571);
nand UO_4878 (O_4878,N_48236,N_48500);
or UO_4879 (O_4879,N_47883,N_49675);
nand UO_4880 (O_4880,N_48363,N_47680);
xnor UO_4881 (O_4881,N_49916,N_48680);
xor UO_4882 (O_4882,N_48226,N_49311);
nor UO_4883 (O_4883,N_48204,N_48326);
nor UO_4884 (O_4884,N_49740,N_49562);
and UO_4885 (O_4885,N_47612,N_47816);
or UO_4886 (O_4886,N_48627,N_47914);
nor UO_4887 (O_4887,N_48438,N_47734);
and UO_4888 (O_4888,N_49362,N_48629);
nand UO_4889 (O_4889,N_49742,N_47537);
and UO_4890 (O_4890,N_48073,N_49448);
xnor UO_4891 (O_4891,N_47957,N_48755);
nor UO_4892 (O_4892,N_48051,N_48510);
xor UO_4893 (O_4893,N_48780,N_48328);
nand UO_4894 (O_4894,N_49137,N_48385);
nor UO_4895 (O_4895,N_47685,N_49535);
nand UO_4896 (O_4896,N_47896,N_47515);
nand UO_4897 (O_4897,N_47748,N_48326);
nand UO_4898 (O_4898,N_48086,N_48473);
xnor UO_4899 (O_4899,N_49283,N_49124);
xor UO_4900 (O_4900,N_48762,N_47888);
nand UO_4901 (O_4901,N_48380,N_48701);
xnor UO_4902 (O_4902,N_48509,N_47760);
nand UO_4903 (O_4903,N_49933,N_48533);
nand UO_4904 (O_4904,N_49649,N_48509);
nand UO_4905 (O_4905,N_48105,N_47885);
xnor UO_4906 (O_4906,N_48387,N_48805);
nor UO_4907 (O_4907,N_49139,N_49526);
and UO_4908 (O_4908,N_48096,N_49834);
nand UO_4909 (O_4909,N_49271,N_48690);
nor UO_4910 (O_4910,N_48612,N_47585);
and UO_4911 (O_4911,N_49708,N_49006);
xnor UO_4912 (O_4912,N_48187,N_48620);
nand UO_4913 (O_4913,N_48918,N_48770);
xor UO_4914 (O_4914,N_49549,N_49912);
nand UO_4915 (O_4915,N_49452,N_48235);
xor UO_4916 (O_4916,N_49931,N_47694);
and UO_4917 (O_4917,N_48731,N_47858);
or UO_4918 (O_4918,N_47996,N_48719);
or UO_4919 (O_4919,N_49131,N_48681);
nor UO_4920 (O_4920,N_49833,N_48553);
nand UO_4921 (O_4921,N_48191,N_48894);
nand UO_4922 (O_4922,N_47560,N_49379);
and UO_4923 (O_4923,N_47784,N_47790);
xor UO_4924 (O_4924,N_49342,N_48292);
or UO_4925 (O_4925,N_48287,N_49189);
nand UO_4926 (O_4926,N_47926,N_49455);
nor UO_4927 (O_4927,N_48081,N_48253);
or UO_4928 (O_4928,N_48553,N_48420);
or UO_4929 (O_4929,N_48784,N_47715);
xor UO_4930 (O_4930,N_47574,N_48115);
and UO_4931 (O_4931,N_47632,N_49424);
nand UO_4932 (O_4932,N_47713,N_49771);
nor UO_4933 (O_4933,N_49654,N_48559);
nor UO_4934 (O_4934,N_49037,N_49354);
xor UO_4935 (O_4935,N_48356,N_48580);
and UO_4936 (O_4936,N_49434,N_48135);
nand UO_4937 (O_4937,N_47509,N_48939);
nand UO_4938 (O_4938,N_48347,N_49642);
nor UO_4939 (O_4939,N_48141,N_47793);
or UO_4940 (O_4940,N_48929,N_49743);
nand UO_4941 (O_4941,N_47554,N_49029);
and UO_4942 (O_4942,N_48302,N_48148);
xor UO_4943 (O_4943,N_49877,N_47529);
xnor UO_4944 (O_4944,N_49245,N_49836);
or UO_4945 (O_4945,N_49310,N_47976);
and UO_4946 (O_4946,N_49313,N_48962);
nand UO_4947 (O_4947,N_49721,N_47729);
xor UO_4948 (O_4948,N_48696,N_49732);
nor UO_4949 (O_4949,N_48802,N_49998);
or UO_4950 (O_4950,N_49370,N_47836);
nor UO_4951 (O_4951,N_48923,N_48996);
and UO_4952 (O_4952,N_48256,N_49856);
xor UO_4953 (O_4953,N_48301,N_47884);
nand UO_4954 (O_4954,N_47949,N_48104);
xor UO_4955 (O_4955,N_48328,N_48741);
nand UO_4956 (O_4956,N_47971,N_48612);
nand UO_4957 (O_4957,N_47788,N_48013);
nand UO_4958 (O_4958,N_49295,N_49346);
nand UO_4959 (O_4959,N_48990,N_49805);
nand UO_4960 (O_4960,N_47761,N_47674);
and UO_4961 (O_4961,N_47834,N_47852);
nor UO_4962 (O_4962,N_48842,N_48475);
nor UO_4963 (O_4963,N_47646,N_47945);
or UO_4964 (O_4964,N_47907,N_47925);
nor UO_4965 (O_4965,N_49411,N_49229);
nor UO_4966 (O_4966,N_49446,N_47578);
nor UO_4967 (O_4967,N_48907,N_49713);
nor UO_4968 (O_4968,N_49143,N_48402);
nand UO_4969 (O_4969,N_49491,N_47851);
nand UO_4970 (O_4970,N_48256,N_49726);
or UO_4971 (O_4971,N_48576,N_47686);
or UO_4972 (O_4972,N_48727,N_47942);
xnor UO_4973 (O_4973,N_47540,N_49763);
xor UO_4974 (O_4974,N_49316,N_49824);
xnor UO_4975 (O_4975,N_49851,N_49782);
or UO_4976 (O_4976,N_49312,N_48620);
xnor UO_4977 (O_4977,N_47958,N_49551);
nor UO_4978 (O_4978,N_48244,N_47523);
xnor UO_4979 (O_4979,N_48854,N_48251);
and UO_4980 (O_4980,N_49372,N_48219);
and UO_4981 (O_4981,N_49081,N_48432);
nand UO_4982 (O_4982,N_48920,N_49975);
and UO_4983 (O_4983,N_49478,N_47773);
nand UO_4984 (O_4984,N_48586,N_47946);
and UO_4985 (O_4985,N_48969,N_48076);
or UO_4986 (O_4986,N_48668,N_48080);
nor UO_4987 (O_4987,N_49791,N_48217);
or UO_4988 (O_4988,N_47840,N_47911);
and UO_4989 (O_4989,N_48976,N_49139);
and UO_4990 (O_4990,N_48490,N_48879);
or UO_4991 (O_4991,N_49715,N_48060);
xnor UO_4992 (O_4992,N_48158,N_48743);
xor UO_4993 (O_4993,N_49425,N_48174);
and UO_4994 (O_4994,N_47638,N_49192);
nand UO_4995 (O_4995,N_48099,N_47958);
xnor UO_4996 (O_4996,N_49150,N_48937);
and UO_4997 (O_4997,N_47802,N_49282);
xor UO_4998 (O_4998,N_49183,N_49655);
xnor UO_4999 (O_4999,N_47893,N_49842);
endmodule