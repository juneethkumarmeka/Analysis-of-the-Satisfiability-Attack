module basic_750_5000_1000_2_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2503,N_2504,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2541,N_2542,N_2543,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2555,N_2556,N_2557,N_2558,N_2559,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2570,N_2571,N_2572,N_2573,N_2575,N_2576,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2599,N_2600,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2612,N_2614,N_2615,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2630,N_2633,N_2634,N_2635,N_2636,N_2637,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2651,N_2652,N_2653,N_2655,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2684,N_2685,N_2687,N_2688,N_2690,N_2691,N_2692,N_2693,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2724,N_2725,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2747,N_2748,N_2749,N_2750,N_2751,N_2753,N_2754,N_2755,N_2757,N_2758,N_2759,N_2760,N_2761,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2787,N_2788,N_2789,N_2790,N_2791,N_2793,N_2795,N_2797,N_2798,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2817,N_2818,N_2819,N_2820,N_2821,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2846,N_2847,N_2848,N_2849,N_2850,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2862,N_2865,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2887,N_2888,N_2889,N_2890,N_2892,N_2893,N_2894,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2904,N_2905,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2925,N_2928,N_2930,N_2931,N_2933,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2967,N_2969,N_2970,N_2973,N_2974,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2985,N_2986,N_2987,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3005,N_3008,N_3009,N_3010,N_3012,N_3013,N_3014,N_3016,N_3017,N_3019,N_3020,N_3021,N_3022,N_3024,N_3026,N_3027,N_3030,N_3031,N_3032,N_3033,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3050,N_3051,N_3052,N_3055,N_3056,N_3057,N_3059,N_3060,N_3061,N_3062,N_3063,N_3065,N_3066,N_3068,N_3071,N_3072,N_3074,N_3075,N_3077,N_3078,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3090,N_3091,N_3092,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3103,N_3105,N_3106,N_3107,N_3111,N_3112,N_3113,N_3114,N_3115,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3128,N_3129,N_3130,N_3131,N_3132,N_3134,N_3137,N_3139,N_3142,N_3143,N_3144,N_3148,N_3149,N_3151,N_3152,N_3153,N_3154,N_3155,N_3157,N_3158,N_3159,N_3161,N_3162,N_3163,N_3164,N_3165,N_3167,N_3169,N_3172,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3182,N_3183,N_3185,N_3187,N_3188,N_3190,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3200,N_3201,N_3202,N_3203,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3230,N_3234,N_3236,N_3238,N_3239,N_3240,N_3241,N_3244,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3254,N_3255,N_3256,N_3258,N_3259,N_3260,N_3261,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3271,N_3272,N_3273,N_3274,N_3276,N_3277,N_3278,N_3280,N_3281,N_3282,N_3283,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3303,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3317,N_3319,N_3320,N_3321,N_3322,N_3325,N_3326,N_3327,N_3329,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3348,N_3349,N_3350,N_3352,N_3353,N_3355,N_3356,N_3357,N_3360,N_3361,N_3362,N_3363,N_3365,N_3366,N_3367,N_3368,N_3369,N_3371,N_3373,N_3374,N_3375,N_3376,N_3377,N_3380,N_3381,N_3382,N_3383,N_3386,N_3388,N_3389,N_3390,N_3391,N_3393,N_3396,N_3398,N_3399,N_3402,N_3403,N_3404,N_3407,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3416,N_3418,N_3419,N_3420,N_3421,N_3422,N_3424,N_3426,N_3428,N_3429,N_3430,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3440,N_3442,N_3443,N_3444,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3457,N_3458,N_3459,N_3460,N_3461,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3473,N_3474,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3483,N_3484,N_3486,N_3487,N_3488,N_3491,N_3492,N_3494,N_3495,N_3496,N_3498,N_3499,N_3500,N_3501,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3520,N_3521,N_3522,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3555,N_3556,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3571,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3586,N_3587,N_3590,N_3592,N_3594,N_3595,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3609,N_3611,N_3612,N_3613,N_3614,N_3615,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3656,N_3658,N_3659,N_3660,N_3661,N_3663,N_3664,N_3665,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3675,N_3676,N_3677,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3729,N_3731,N_3732,N_3733,N_3735,N_3736,N_3737,N_3739,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3750,N_3751,N_3754,N_3756,N_3757,N_3759,N_3760,N_3761,N_3762,N_3763,N_3765,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3777,N_3778,N_3779,N_3781,N_3782,N_3784,N_3785,N_3787,N_3789,N_3790,N_3792,N_3793,N_3796,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3805,N_3806,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3825,N_3826,N_3828,N_3830,N_3832,N_3833,N_3834,N_3836,N_3837,N_3838,N_3839,N_3841,N_3842,N_3843,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3873,N_3874,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3883,N_3884,N_3885,N_3887,N_3888,N_3889,N_3890,N_3891,N_3893,N_3894,N_3895,N_3896,N_3898,N_3899,N_3900,N_3902,N_3903,N_3904,N_3905,N_3907,N_3909,N_3910,N_3911,N_3913,N_3914,N_3915,N_3917,N_3918,N_3919,N_3921,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3940,N_3941,N_3942,N_3943,N_3945,N_3946,N_3947,N_3949,N_3950,N_3951,N_3952,N_3953,N_3957,N_3958,N_3959,N_3961,N_3962,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3982,N_3983,N_3984,N_3986,N_3987,N_3989,N_3990,N_3991,N_3992,N_3993,N_3996,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4026,N_4027,N_4029,N_4030,N_4032,N_4033,N_4034,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4057,N_4059,N_4060,N_4062,N_4063,N_4065,N_4067,N_4068,N_4069,N_4071,N_4072,N_4073,N_4074,N_4076,N_4078,N_4079,N_4080,N_4081,N_4082,N_4084,N_4085,N_4088,N_4089,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4098,N_4099,N_4100,N_4102,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4145,N_4147,N_4149,N_4150,N_4152,N_4153,N_4154,N_4155,N_4157,N_4158,N_4159,N_4160,N_4161,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4187,N_4188,N_4190,N_4191,N_4194,N_4196,N_4197,N_4198,N_4199,N_4200,N_4202,N_4204,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4274,N_4275,N_4276,N_4278,N_4279,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4296,N_4297,N_4298,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4317,N_4319,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4347,N_4348,N_4350,N_4351,N_4355,N_4356,N_4357,N_4358,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4367,N_4368,N_4369,N_4370,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4379,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4409,N_4410,N_4411,N_4412,N_4413,N_4415,N_4416,N_4417,N_4420,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4444,N_4445,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4472,N_4473,N_4474,N_4475,N_4476,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4496,N_4497,N_4498,N_4499,N_4500,N_4503,N_4504,N_4505,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4517,N_4518,N_4519,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4541,N_4542,N_4544,N_4545,N_4546,N_4547,N_4549,N_4550,N_4551,N_4552,N_4554,N_4555,N_4557,N_4558,N_4559,N_4560,N_4561,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4594,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4606,N_4607,N_4608,N_4609,N_4610,N_4612,N_4613,N_4614,N_4616,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4628,N_4629,N_4630,N_4631,N_4632,N_4634,N_4635,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4658,N_4659,N_4660,N_4661,N_4662,N_4664,N_4665,N_4666,N_4667,N_4669,N_4670,N_4672,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4683,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4728,N_4730,N_4732,N_4733,N_4734,N_4735,N_4736,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4766,N_4767,N_4768,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4777,N_4778,N_4779,N_4780,N_4781,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4803,N_4804,N_4805,N_4806,N_4807,N_4809,N_4810,N_4811,N_4812,N_4814,N_4815,N_4816,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4860,N_4861,N_4862,N_4863,N_4866,N_4867,N_4868,N_4869,N_4870,N_4872,N_4873,N_4874,N_4875,N_4877,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4915,N_4916,N_4917,N_4918,N_4919,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4932,N_4933,N_4934,N_4935,N_4937,N_4938,N_4939,N_4941,N_4942,N_4944,N_4945,N_4946,N_4947,N_4949,N_4950,N_4951,N_4953,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4986,N_4987,N_4988,N_4989,N_4990,N_4992,N_4993,N_4994,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_318,In_300);
or U1 (N_1,In_477,In_743);
and U2 (N_2,In_92,In_462);
nor U3 (N_3,In_431,In_668);
and U4 (N_4,In_536,In_369);
nand U5 (N_5,In_238,In_191);
or U6 (N_6,In_732,In_167);
nor U7 (N_7,In_727,In_235);
nand U8 (N_8,In_19,In_210);
nor U9 (N_9,In_422,In_733);
or U10 (N_10,In_298,In_365);
and U11 (N_11,In_691,In_411);
or U12 (N_12,In_159,In_450);
nand U13 (N_13,In_185,In_680);
nor U14 (N_14,In_35,In_56);
nor U15 (N_15,In_270,In_43);
or U16 (N_16,In_459,In_98);
and U17 (N_17,In_272,In_460);
nor U18 (N_18,In_227,In_513);
nand U19 (N_19,In_657,In_271);
nand U20 (N_20,In_340,In_47);
nor U21 (N_21,In_140,In_664);
or U22 (N_22,In_722,In_103);
nand U23 (N_23,In_430,In_223);
nor U24 (N_24,In_403,In_489);
or U25 (N_25,In_586,In_22);
nand U26 (N_26,In_330,In_237);
or U27 (N_27,In_281,In_372);
or U28 (N_28,In_173,In_111);
and U29 (N_29,In_120,In_518);
nor U30 (N_30,In_453,In_714);
nor U31 (N_31,In_410,In_452);
or U32 (N_32,In_283,In_163);
or U33 (N_33,In_1,In_472);
or U34 (N_34,In_537,In_8);
or U35 (N_35,In_746,In_89);
or U36 (N_36,In_707,In_323);
nor U37 (N_37,In_614,In_484);
or U38 (N_38,In_418,In_224);
and U39 (N_39,In_735,In_48);
and U40 (N_40,In_348,In_646);
and U41 (N_41,In_189,In_730);
and U42 (N_42,In_661,In_608);
or U43 (N_43,In_294,In_108);
nand U44 (N_44,In_442,In_692);
nand U45 (N_45,In_389,In_675);
or U46 (N_46,In_391,In_617);
and U47 (N_47,In_506,In_571);
and U48 (N_48,In_166,In_558);
nand U49 (N_49,In_457,In_343);
nor U50 (N_50,In_219,In_665);
nor U51 (N_51,In_704,In_151);
nor U52 (N_52,In_543,In_468);
or U53 (N_53,In_458,In_307);
or U54 (N_54,In_611,In_44);
and U55 (N_55,In_154,In_544);
and U56 (N_56,In_473,In_639);
or U57 (N_57,In_315,In_624);
or U58 (N_58,In_427,In_125);
nor U59 (N_59,In_501,In_240);
or U60 (N_60,In_16,In_115);
nand U61 (N_61,In_350,In_697);
nand U62 (N_62,In_532,In_612);
and U63 (N_63,In_726,In_244);
or U64 (N_64,In_336,In_126);
nor U65 (N_65,In_519,In_723);
nand U66 (N_66,In_717,In_200);
or U67 (N_67,In_41,In_696);
or U68 (N_68,In_289,In_647);
or U69 (N_69,In_160,In_408);
and U70 (N_70,In_316,In_604);
nand U71 (N_71,In_677,In_362);
nor U72 (N_72,In_253,In_64);
or U73 (N_73,In_539,In_375);
nand U74 (N_74,In_358,In_526);
nand U75 (N_75,In_404,In_74);
nand U76 (N_76,In_494,In_119);
and U77 (N_77,In_203,In_280);
or U78 (N_78,In_613,In_88);
or U79 (N_79,In_168,In_734);
or U80 (N_80,In_371,In_585);
nor U81 (N_81,In_602,In_80);
nand U82 (N_82,In_226,In_748);
or U83 (N_83,In_708,In_291);
nor U84 (N_84,In_352,In_21);
and U85 (N_85,In_498,In_106);
nor U86 (N_86,In_178,In_40);
nor U87 (N_87,In_693,In_250);
nor U88 (N_88,In_478,In_215);
nand U89 (N_89,In_355,In_123);
nor U90 (N_90,In_268,In_58);
nand U91 (N_91,In_738,In_86);
and U92 (N_92,In_533,In_45);
nand U93 (N_93,In_405,In_231);
or U94 (N_94,In_229,In_275);
or U95 (N_95,In_715,In_520);
and U96 (N_96,In_170,In_700);
and U97 (N_97,In_82,In_214);
nand U98 (N_98,In_188,In_491);
and U99 (N_99,In_562,In_671);
nand U100 (N_100,In_525,In_322);
and U101 (N_101,In_161,In_186);
or U102 (N_102,In_469,In_312);
and U103 (N_103,In_694,In_504);
nor U104 (N_104,In_552,In_256);
or U105 (N_105,In_625,In_242);
nor U106 (N_106,In_699,In_334);
nor U107 (N_107,In_95,In_445);
nand U108 (N_108,In_156,In_337);
and U109 (N_109,In_407,In_678);
and U110 (N_110,In_109,In_690);
nor U111 (N_111,In_338,In_740);
and U112 (N_112,In_20,In_703);
or U113 (N_113,In_12,In_616);
nand U114 (N_114,In_172,In_202);
or U115 (N_115,In_667,In_297);
or U116 (N_116,In_666,In_341);
nand U117 (N_117,In_252,In_509);
or U118 (N_118,In_580,In_654);
or U119 (N_119,In_197,In_364);
and U120 (N_120,In_42,In_397);
nand U121 (N_121,In_447,In_4);
nor U122 (N_122,In_248,In_61);
and U123 (N_123,In_195,In_465);
nor U124 (N_124,In_183,In_480);
nor U125 (N_125,In_32,In_205);
and U126 (N_126,In_635,In_236);
nand U127 (N_127,In_531,In_288);
and U128 (N_128,In_598,In_425);
nand U129 (N_129,In_642,In_475);
or U130 (N_130,In_524,In_438);
nand U131 (N_131,In_9,In_510);
and U132 (N_132,In_116,In_607);
nand U133 (N_133,In_303,In_204);
and U134 (N_134,In_36,In_637);
or U135 (N_135,In_541,In_326);
and U136 (N_136,In_424,In_545);
and U137 (N_137,In_634,In_486);
nand U138 (N_138,In_241,In_650);
nand U139 (N_139,In_588,In_104);
or U140 (N_140,In_534,In_739);
or U141 (N_141,In_29,In_681);
and U142 (N_142,In_349,In_266);
and U143 (N_143,In_550,In_101);
nor U144 (N_144,In_555,In_409);
and U145 (N_145,In_132,In_744);
or U146 (N_146,In_594,In_522);
and U147 (N_147,In_557,In_622);
nor U148 (N_148,In_228,In_609);
nor U149 (N_149,In_345,In_648);
or U150 (N_150,In_426,In_451);
nor U151 (N_151,In_630,In_702);
nand U152 (N_152,In_179,In_652);
or U153 (N_153,In_387,In_245);
or U154 (N_154,In_31,In_261);
or U155 (N_155,In_146,In_276);
or U156 (N_156,In_333,In_466);
nor U157 (N_157,In_716,In_379);
and U158 (N_158,In_269,In_570);
or U159 (N_159,In_134,In_90);
nor U160 (N_160,In_600,In_34);
nand U161 (N_161,In_496,In_569);
and U162 (N_162,In_311,In_279);
or U163 (N_163,In_512,In_328);
or U164 (N_164,In_249,In_376);
nor U165 (N_165,In_164,In_470);
nor U166 (N_166,In_314,In_105);
or U167 (N_167,In_626,In_147);
nor U168 (N_168,In_467,In_685);
and U169 (N_169,In_382,In_290);
or U170 (N_170,In_412,In_107);
or U171 (N_171,In_720,In_413);
nand U172 (N_172,In_117,In_402);
nor U173 (N_173,In_464,In_361);
nor U174 (N_174,In_479,In_623);
nand U175 (N_175,In_24,In_69);
nand U176 (N_176,In_595,In_566);
and U177 (N_177,In_251,In_267);
and U178 (N_178,In_420,In_527);
nor U179 (N_179,In_419,In_25);
and U180 (N_180,In_71,In_517);
nor U181 (N_181,In_423,In_388);
nor U182 (N_182,In_535,In_313);
or U183 (N_183,In_15,In_142);
and U184 (N_184,In_296,In_653);
nand U185 (N_185,In_135,In_414);
nor U186 (N_186,In_670,In_574);
and U187 (N_187,In_96,In_706);
and U188 (N_188,In_332,In_278);
or U189 (N_189,In_390,In_674);
nor U190 (N_190,In_564,In_719);
or U191 (N_191,In_136,In_736);
and U192 (N_192,In_193,In_57);
or U193 (N_193,In_91,In_621);
nor U194 (N_194,In_579,In_474);
nand U195 (N_195,In_218,In_201);
nor U196 (N_196,In_53,In_139);
nand U197 (N_197,In_2,In_721);
nor U198 (N_198,In_503,In_73);
nor U199 (N_199,In_13,In_689);
nand U200 (N_200,In_78,In_380);
or U201 (N_201,In_663,In_428);
nor U202 (N_202,In_745,In_565);
nand U203 (N_203,In_177,In_437);
and U204 (N_204,In_645,In_711);
or U205 (N_205,In_317,In_605);
nor U206 (N_206,In_575,In_687);
or U207 (N_207,In_23,In_577);
and U208 (N_208,In_488,In_187);
nor U209 (N_209,In_180,In_599);
nand U210 (N_210,In_93,In_737);
nor U211 (N_211,In_399,In_302);
or U212 (N_212,In_521,In_357);
nand U213 (N_213,In_384,In_265);
or U214 (N_214,In_137,In_698);
nor U215 (N_215,In_640,In_686);
and U216 (N_216,In_370,In_655);
nor U217 (N_217,In_455,In_556);
or U218 (N_218,In_293,In_432);
and U219 (N_219,In_208,In_401);
nand U220 (N_220,In_295,In_439);
nand U221 (N_221,In_55,In_216);
nand U222 (N_222,In_331,In_217);
nor U223 (N_223,In_99,In_514);
or U224 (N_224,In_485,In_483);
nand U225 (N_225,In_672,In_644);
and U226 (N_226,In_335,In_502);
or U227 (N_227,In_162,In_259);
nand U228 (N_228,In_153,In_84);
and U229 (N_229,In_695,In_615);
or U230 (N_230,In_500,In_587);
and U231 (N_231,In_392,In_14);
nor U232 (N_232,In_567,In_277);
nand U233 (N_233,In_286,In_239);
and U234 (N_234,In_515,In_339);
nor U235 (N_235,In_551,In_393);
and U236 (N_236,In_433,In_589);
and U237 (N_237,In_68,In_461);
and U238 (N_238,In_150,In_148);
and U239 (N_239,In_492,In_100);
and U240 (N_240,In_346,In_274);
and U241 (N_241,In_597,In_70);
nor U242 (N_242,In_516,In_495);
and U243 (N_243,In_220,In_122);
and U244 (N_244,In_308,In_523);
nand U245 (N_245,In_128,In_581);
and U246 (N_246,In_66,In_131);
or U247 (N_247,In_596,In_378);
or U248 (N_248,In_232,In_287);
and U249 (N_249,In_206,In_631);
or U250 (N_250,In_17,In_454);
nor U251 (N_251,In_542,In_385);
nor U252 (N_252,In_742,In_285);
nor U253 (N_253,In_27,In_212);
nand U254 (N_254,In_560,In_610);
nor U255 (N_255,In_138,In_747);
nand U256 (N_256,In_124,In_234);
or U257 (N_257,In_563,In_310);
or U258 (N_258,In_87,In_366);
nor U259 (N_259,In_632,In_656);
nor U260 (N_260,In_52,In_729);
nand U261 (N_261,In_76,In_324);
nor U262 (N_262,In_304,In_230);
nor U263 (N_263,In_582,In_222);
nand U264 (N_264,In_712,In_353);
or U265 (N_265,In_559,In_264);
nor U266 (N_266,In_673,In_505);
nand U267 (N_267,In_568,In_499);
or U268 (N_268,In_493,In_171);
nand U269 (N_269,In_415,In_368);
or U270 (N_270,In_471,In_643);
or U271 (N_271,In_476,In_155);
nor U272 (N_272,In_174,In_627);
or U273 (N_273,In_254,In_97);
or U274 (N_274,In_50,In_37);
or U275 (N_275,In_143,In_416);
nand U276 (N_276,In_243,In_725);
nor U277 (N_277,In_434,In_59);
or U278 (N_278,In_446,In_246);
nand U279 (N_279,In_396,In_121);
nand U280 (N_280,In_114,In_709);
or U281 (N_281,In_731,In_741);
and U282 (N_282,In_75,In_309);
nor U283 (N_283,In_628,In_110);
or U284 (N_284,In_33,In_481);
nor U285 (N_285,In_629,In_60);
nand U286 (N_286,In_342,In_169);
nor U287 (N_287,In_530,In_327);
or U288 (N_288,In_603,In_7);
and U289 (N_289,In_3,In_18);
nand U290 (N_290,In_28,In_94);
or U291 (N_291,In_320,In_129);
nand U292 (N_292,In_38,In_344);
nor U293 (N_293,In_688,In_54);
or U294 (N_294,In_260,In_436);
nor U295 (N_295,In_386,In_62);
or U296 (N_296,In_30,In_705);
and U297 (N_297,In_659,In_724);
or U298 (N_298,In_507,In_490);
or U299 (N_299,In_394,In_576);
or U300 (N_300,In_181,In_618);
nor U301 (N_301,In_540,In_429);
nor U302 (N_302,In_440,In_676);
and U303 (N_303,In_118,In_39);
nand U304 (N_304,In_553,In_435);
or U305 (N_305,In_158,In_301);
nand U306 (N_306,In_196,In_548);
or U307 (N_307,In_549,In_601);
and U308 (N_308,In_133,In_593);
nor U309 (N_309,In_347,In_583);
or U310 (N_310,In_620,In_207);
nor U311 (N_311,In_710,In_669);
and U312 (N_312,In_547,In_46);
xor U313 (N_313,In_511,In_329);
nand U314 (N_314,In_592,In_590);
nor U315 (N_315,In_157,In_65);
nor U316 (N_316,In_658,In_141);
or U317 (N_317,In_258,In_211);
or U318 (N_318,In_395,In_374);
and U319 (N_319,In_529,In_263);
nor U320 (N_320,In_79,In_194);
and U321 (N_321,In_11,In_354);
nand U322 (N_322,In_373,In_561);
nand U323 (N_323,In_359,In_292);
nor U324 (N_324,In_255,In_538);
and U325 (N_325,In_152,In_381);
or U326 (N_326,In_83,In_528);
and U327 (N_327,In_701,In_456);
nor U328 (N_328,In_262,In_26);
or U329 (N_329,In_619,In_554);
nor U330 (N_330,In_463,In_367);
nor U331 (N_331,In_398,In_85);
nand U332 (N_332,In_72,In_572);
nand U333 (N_333,In_225,In_5);
nand U334 (N_334,In_683,In_273);
and U335 (N_335,In_377,In_10);
nor U336 (N_336,In_417,In_321);
or U337 (N_337,In_6,In_351);
and U338 (N_338,In_546,In_641);
and U339 (N_339,In_728,In_448);
nor U340 (N_340,In_282,In_406);
nand U341 (N_341,In_299,In_130);
or U342 (N_342,In_176,In_198);
and U343 (N_343,In_199,In_578);
nor U344 (N_344,In_182,In_636);
and U345 (N_345,In_144,In_508);
and U346 (N_346,In_660,In_441);
nor U347 (N_347,In_81,In_684);
and U348 (N_348,In_584,In_233);
nor U349 (N_349,In_319,In_0);
and U350 (N_350,In_487,In_165);
or U351 (N_351,In_606,In_257);
or U352 (N_352,In_591,In_306);
and U353 (N_353,In_444,In_184);
nor U354 (N_354,In_325,In_209);
and U355 (N_355,In_113,In_284);
nand U356 (N_356,In_305,In_77);
nand U357 (N_357,In_497,In_718);
or U358 (N_358,In_63,In_679);
nand U359 (N_359,In_400,In_102);
and U360 (N_360,In_149,In_482);
nand U361 (N_361,In_175,In_192);
nor U362 (N_362,In_221,In_443);
and U363 (N_363,In_682,In_749);
nand U364 (N_364,In_247,In_662);
or U365 (N_365,In_213,In_356);
nand U366 (N_366,In_145,In_633);
or U367 (N_367,In_421,In_713);
or U368 (N_368,In_651,In_67);
nor U369 (N_369,In_363,In_190);
nor U370 (N_370,In_383,In_127);
nand U371 (N_371,In_649,In_49);
and U372 (N_372,In_112,In_360);
nand U373 (N_373,In_449,In_51);
nand U374 (N_374,In_573,In_638);
or U375 (N_375,In_184,In_76);
nor U376 (N_376,In_385,In_140);
or U377 (N_377,In_467,In_694);
nor U378 (N_378,In_85,In_244);
and U379 (N_379,In_443,In_556);
nand U380 (N_380,In_459,In_389);
nor U381 (N_381,In_227,In_21);
nor U382 (N_382,In_451,In_187);
xor U383 (N_383,In_202,In_226);
nor U384 (N_384,In_737,In_274);
or U385 (N_385,In_293,In_568);
nand U386 (N_386,In_59,In_417);
nand U387 (N_387,In_195,In_462);
or U388 (N_388,In_658,In_347);
nand U389 (N_389,In_555,In_10);
nor U390 (N_390,In_522,In_388);
or U391 (N_391,In_128,In_428);
and U392 (N_392,In_696,In_508);
and U393 (N_393,In_307,In_728);
nand U394 (N_394,In_442,In_402);
and U395 (N_395,In_555,In_1);
and U396 (N_396,In_643,In_389);
nand U397 (N_397,In_257,In_603);
nor U398 (N_398,In_475,In_267);
and U399 (N_399,In_216,In_683);
nor U400 (N_400,In_706,In_452);
or U401 (N_401,In_111,In_126);
and U402 (N_402,In_709,In_614);
and U403 (N_403,In_123,In_617);
nand U404 (N_404,In_316,In_315);
and U405 (N_405,In_30,In_531);
nor U406 (N_406,In_285,In_184);
and U407 (N_407,In_446,In_685);
nand U408 (N_408,In_179,In_609);
or U409 (N_409,In_700,In_74);
or U410 (N_410,In_214,In_455);
or U411 (N_411,In_295,In_547);
nand U412 (N_412,In_411,In_461);
nand U413 (N_413,In_389,In_410);
nand U414 (N_414,In_378,In_663);
nand U415 (N_415,In_418,In_424);
xnor U416 (N_416,In_218,In_232);
nand U417 (N_417,In_44,In_528);
and U418 (N_418,In_613,In_76);
nor U419 (N_419,In_236,In_195);
nand U420 (N_420,In_514,In_116);
or U421 (N_421,In_284,In_602);
or U422 (N_422,In_565,In_363);
and U423 (N_423,In_410,In_439);
nand U424 (N_424,In_424,In_710);
nor U425 (N_425,In_259,In_45);
or U426 (N_426,In_82,In_304);
or U427 (N_427,In_585,In_273);
nor U428 (N_428,In_715,In_295);
or U429 (N_429,In_634,In_115);
and U430 (N_430,In_25,In_631);
nor U431 (N_431,In_143,In_534);
or U432 (N_432,In_239,In_362);
nor U433 (N_433,In_139,In_164);
and U434 (N_434,In_326,In_0);
nand U435 (N_435,In_489,In_473);
nand U436 (N_436,In_142,In_561);
and U437 (N_437,In_410,In_531);
nand U438 (N_438,In_245,In_187);
or U439 (N_439,In_244,In_651);
nor U440 (N_440,In_382,In_381);
and U441 (N_441,In_29,In_390);
and U442 (N_442,In_451,In_730);
nor U443 (N_443,In_654,In_342);
nand U444 (N_444,In_92,In_747);
nand U445 (N_445,In_666,In_673);
or U446 (N_446,In_696,In_541);
and U447 (N_447,In_607,In_695);
nand U448 (N_448,In_125,In_101);
nor U449 (N_449,In_98,In_17);
nand U450 (N_450,In_722,In_446);
and U451 (N_451,In_363,In_202);
nor U452 (N_452,In_256,In_429);
or U453 (N_453,In_212,In_86);
and U454 (N_454,In_718,In_414);
nand U455 (N_455,In_37,In_482);
and U456 (N_456,In_58,In_376);
nand U457 (N_457,In_604,In_112);
nand U458 (N_458,In_459,In_123);
nand U459 (N_459,In_577,In_634);
or U460 (N_460,In_547,In_575);
nand U461 (N_461,In_708,In_35);
or U462 (N_462,In_238,In_463);
or U463 (N_463,In_1,In_340);
and U464 (N_464,In_464,In_206);
nand U465 (N_465,In_140,In_609);
nor U466 (N_466,In_204,In_495);
or U467 (N_467,In_629,In_329);
or U468 (N_468,In_509,In_423);
nand U469 (N_469,In_502,In_301);
nor U470 (N_470,In_604,In_530);
xor U471 (N_471,In_54,In_504);
nand U472 (N_472,In_377,In_709);
nand U473 (N_473,In_124,In_462);
nor U474 (N_474,In_500,In_693);
and U475 (N_475,In_269,In_582);
nand U476 (N_476,In_560,In_646);
nor U477 (N_477,In_88,In_694);
nand U478 (N_478,In_82,In_326);
nor U479 (N_479,In_81,In_46);
or U480 (N_480,In_345,In_93);
and U481 (N_481,In_398,In_4);
nand U482 (N_482,In_8,In_307);
and U483 (N_483,In_516,In_445);
and U484 (N_484,In_670,In_524);
and U485 (N_485,In_250,In_384);
nand U486 (N_486,In_21,In_236);
and U487 (N_487,In_179,In_695);
or U488 (N_488,In_41,In_626);
and U489 (N_489,In_749,In_673);
or U490 (N_490,In_251,In_469);
nand U491 (N_491,In_128,In_199);
nor U492 (N_492,In_326,In_530);
and U493 (N_493,In_251,In_688);
or U494 (N_494,In_260,In_406);
and U495 (N_495,In_601,In_529);
and U496 (N_496,In_536,In_450);
or U497 (N_497,In_717,In_256);
or U498 (N_498,In_634,In_225);
nor U499 (N_499,In_317,In_284);
nor U500 (N_500,In_720,In_529);
and U501 (N_501,In_214,In_374);
or U502 (N_502,In_655,In_310);
and U503 (N_503,In_743,In_335);
or U504 (N_504,In_498,In_126);
or U505 (N_505,In_313,In_693);
and U506 (N_506,In_188,In_271);
nand U507 (N_507,In_460,In_655);
nor U508 (N_508,In_115,In_385);
nor U509 (N_509,In_659,In_251);
nand U510 (N_510,In_658,In_655);
and U511 (N_511,In_220,In_733);
and U512 (N_512,In_709,In_136);
nor U513 (N_513,In_39,In_544);
and U514 (N_514,In_461,In_745);
nand U515 (N_515,In_349,In_699);
or U516 (N_516,In_671,In_104);
nor U517 (N_517,In_659,In_459);
and U518 (N_518,In_379,In_702);
or U519 (N_519,In_219,In_207);
nor U520 (N_520,In_177,In_382);
nand U521 (N_521,In_469,In_696);
nand U522 (N_522,In_9,In_408);
and U523 (N_523,In_341,In_327);
nand U524 (N_524,In_523,In_433);
and U525 (N_525,In_142,In_182);
and U526 (N_526,In_711,In_346);
nor U527 (N_527,In_0,In_180);
nor U528 (N_528,In_555,In_559);
or U529 (N_529,In_720,In_112);
nor U530 (N_530,In_439,In_320);
nor U531 (N_531,In_300,In_23);
nor U532 (N_532,In_353,In_675);
nand U533 (N_533,In_631,In_558);
or U534 (N_534,In_555,In_231);
nor U535 (N_535,In_739,In_106);
or U536 (N_536,In_709,In_714);
or U537 (N_537,In_416,In_498);
or U538 (N_538,In_460,In_357);
or U539 (N_539,In_480,In_203);
nand U540 (N_540,In_173,In_311);
nand U541 (N_541,In_72,In_318);
or U542 (N_542,In_244,In_71);
and U543 (N_543,In_377,In_167);
or U544 (N_544,In_118,In_451);
and U545 (N_545,In_50,In_546);
and U546 (N_546,In_279,In_614);
nor U547 (N_547,In_264,In_665);
and U548 (N_548,In_613,In_676);
nand U549 (N_549,In_471,In_136);
and U550 (N_550,In_69,In_327);
and U551 (N_551,In_602,In_724);
nand U552 (N_552,In_570,In_169);
nand U553 (N_553,In_367,In_115);
nor U554 (N_554,In_390,In_115);
nand U555 (N_555,In_332,In_217);
or U556 (N_556,In_220,In_420);
nand U557 (N_557,In_442,In_691);
nor U558 (N_558,In_461,In_147);
nor U559 (N_559,In_36,In_732);
nor U560 (N_560,In_68,In_592);
nand U561 (N_561,In_713,In_431);
nor U562 (N_562,In_637,In_86);
or U563 (N_563,In_599,In_650);
or U564 (N_564,In_711,In_102);
and U565 (N_565,In_337,In_271);
and U566 (N_566,In_634,In_285);
and U567 (N_567,In_490,In_99);
or U568 (N_568,In_623,In_188);
and U569 (N_569,In_626,In_155);
or U570 (N_570,In_653,In_265);
or U571 (N_571,In_46,In_664);
or U572 (N_572,In_481,In_115);
or U573 (N_573,In_67,In_518);
nand U574 (N_574,In_332,In_468);
nand U575 (N_575,In_444,In_485);
nand U576 (N_576,In_294,In_187);
nor U577 (N_577,In_738,In_27);
and U578 (N_578,In_431,In_0);
nor U579 (N_579,In_186,In_204);
and U580 (N_580,In_672,In_5);
and U581 (N_581,In_320,In_63);
or U582 (N_582,In_150,In_63);
and U583 (N_583,In_307,In_467);
nand U584 (N_584,In_268,In_551);
or U585 (N_585,In_190,In_125);
nand U586 (N_586,In_736,In_596);
and U587 (N_587,In_287,In_43);
or U588 (N_588,In_248,In_579);
or U589 (N_589,In_661,In_429);
nand U590 (N_590,In_662,In_334);
nand U591 (N_591,In_289,In_604);
nor U592 (N_592,In_118,In_321);
or U593 (N_593,In_376,In_404);
nand U594 (N_594,In_356,In_223);
and U595 (N_595,In_710,In_146);
or U596 (N_596,In_280,In_540);
and U597 (N_597,In_479,In_589);
nand U598 (N_598,In_460,In_81);
nor U599 (N_599,In_149,In_421);
and U600 (N_600,In_38,In_167);
xnor U601 (N_601,In_565,In_699);
or U602 (N_602,In_412,In_121);
nor U603 (N_603,In_166,In_636);
and U604 (N_604,In_414,In_130);
or U605 (N_605,In_263,In_376);
nor U606 (N_606,In_69,In_96);
nor U607 (N_607,In_326,In_470);
nand U608 (N_608,In_647,In_619);
nand U609 (N_609,In_580,In_358);
nor U610 (N_610,In_123,In_47);
and U611 (N_611,In_553,In_286);
and U612 (N_612,In_230,In_637);
nor U613 (N_613,In_247,In_265);
nor U614 (N_614,In_141,In_108);
nand U615 (N_615,In_413,In_28);
nor U616 (N_616,In_558,In_720);
nor U617 (N_617,In_312,In_36);
nand U618 (N_618,In_525,In_618);
nor U619 (N_619,In_310,In_558);
or U620 (N_620,In_275,In_293);
and U621 (N_621,In_335,In_224);
or U622 (N_622,In_535,In_151);
nor U623 (N_623,In_401,In_684);
nand U624 (N_624,In_194,In_567);
nor U625 (N_625,In_313,In_482);
nand U626 (N_626,In_711,In_343);
nand U627 (N_627,In_128,In_332);
nor U628 (N_628,In_73,In_399);
and U629 (N_629,In_746,In_71);
nor U630 (N_630,In_403,In_320);
nand U631 (N_631,In_184,In_435);
nand U632 (N_632,In_320,In_417);
and U633 (N_633,In_178,In_158);
and U634 (N_634,In_242,In_118);
and U635 (N_635,In_148,In_375);
or U636 (N_636,In_617,In_37);
and U637 (N_637,In_289,In_710);
nor U638 (N_638,In_627,In_596);
and U639 (N_639,In_83,In_647);
nor U640 (N_640,In_735,In_362);
nor U641 (N_641,In_723,In_426);
and U642 (N_642,In_345,In_163);
or U643 (N_643,In_640,In_96);
nor U644 (N_644,In_321,In_613);
nand U645 (N_645,In_377,In_714);
nor U646 (N_646,In_296,In_137);
nor U647 (N_647,In_566,In_99);
or U648 (N_648,In_616,In_265);
nand U649 (N_649,In_637,In_49);
and U650 (N_650,In_553,In_244);
nor U651 (N_651,In_487,In_462);
or U652 (N_652,In_291,In_3);
and U653 (N_653,In_105,In_674);
and U654 (N_654,In_714,In_678);
nor U655 (N_655,In_678,In_42);
nor U656 (N_656,In_160,In_484);
nor U657 (N_657,In_742,In_506);
nand U658 (N_658,In_198,In_110);
or U659 (N_659,In_695,In_588);
or U660 (N_660,In_365,In_417);
nor U661 (N_661,In_199,In_418);
nand U662 (N_662,In_524,In_487);
nor U663 (N_663,In_186,In_582);
or U664 (N_664,In_706,In_671);
and U665 (N_665,In_640,In_625);
and U666 (N_666,In_521,In_293);
or U667 (N_667,In_320,In_237);
xnor U668 (N_668,In_189,In_574);
and U669 (N_669,In_245,In_314);
or U670 (N_670,In_653,In_336);
nand U671 (N_671,In_230,In_680);
nand U672 (N_672,In_254,In_52);
nor U673 (N_673,In_398,In_660);
or U674 (N_674,In_276,In_272);
or U675 (N_675,In_650,In_614);
nand U676 (N_676,In_422,In_356);
nand U677 (N_677,In_105,In_441);
and U678 (N_678,In_21,In_455);
and U679 (N_679,In_739,In_121);
and U680 (N_680,In_228,In_540);
nor U681 (N_681,In_136,In_399);
or U682 (N_682,In_103,In_148);
and U683 (N_683,In_21,In_556);
nor U684 (N_684,In_634,In_585);
nor U685 (N_685,In_666,In_436);
xnor U686 (N_686,In_147,In_141);
or U687 (N_687,In_339,In_233);
or U688 (N_688,In_495,In_388);
or U689 (N_689,In_680,In_172);
nor U690 (N_690,In_676,In_567);
nor U691 (N_691,In_387,In_556);
or U692 (N_692,In_426,In_492);
and U693 (N_693,In_614,In_326);
or U694 (N_694,In_421,In_201);
nand U695 (N_695,In_98,In_530);
or U696 (N_696,In_691,In_464);
and U697 (N_697,In_748,In_5);
nor U698 (N_698,In_96,In_543);
and U699 (N_699,In_207,In_589);
nand U700 (N_700,In_29,In_242);
nor U701 (N_701,In_299,In_421);
nor U702 (N_702,In_743,In_681);
and U703 (N_703,In_400,In_6);
or U704 (N_704,In_378,In_244);
or U705 (N_705,In_296,In_132);
nand U706 (N_706,In_713,In_142);
or U707 (N_707,In_343,In_239);
nor U708 (N_708,In_400,In_512);
nor U709 (N_709,In_291,In_304);
or U710 (N_710,In_349,In_222);
or U711 (N_711,In_374,In_335);
nor U712 (N_712,In_376,In_415);
nor U713 (N_713,In_269,In_720);
nor U714 (N_714,In_690,In_334);
or U715 (N_715,In_83,In_361);
or U716 (N_716,In_92,In_691);
nor U717 (N_717,In_318,In_409);
nor U718 (N_718,In_179,In_687);
and U719 (N_719,In_46,In_383);
nand U720 (N_720,In_645,In_732);
nor U721 (N_721,In_501,In_535);
and U722 (N_722,In_428,In_203);
and U723 (N_723,In_515,In_27);
nor U724 (N_724,In_60,In_182);
nand U725 (N_725,In_706,In_141);
and U726 (N_726,In_430,In_427);
or U727 (N_727,In_275,In_645);
nand U728 (N_728,In_60,In_418);
nor U729 (N_729,In_390,In_150);
and U730 (N_730,In_368,In_113);
or U731 (N_731,In_318,In_236);
nand U732 (N_732,In_229,In_288);
and U733 (N_733,In_0,In_685);
or U734 (N_734,In_232,In_640);
nor U735 (N_735,In_671,In_236);
nor U736 (N_736,In_218,In_730);
nand U737 (N_737,In_612,In_340);
nor U738 (N_738,In_16,In_320);
nor U739 (N_739,In_70,In_21);
nand U740 (N_740,In_309,In_111);
and U741 (N_741,In_582,In_67);
nor U742 (N_742,In_110,In_555);
nand U743 (N_743,In_441,In_632);
nor U744 (N_744,In_12,In_397);
and U745 (N_745,In_699,In_643);
nor U746 (N_746,In_2,In_249);
nor U747 (N_747,In_47,In_183);
nand U748 (N_748,In_349,In_198);
or U749 (N_749,In_657,In_656);
nand U750 (N_750,In_141,In_86);
or U751 (N_751,In_661,In_537);
and U752 (N_752,In_53,In_458);
and U753 (N_753,In_242,In_398);
and U754 (N_754,In_186,In_431);
and U755 (N_755,In_12,In_517);
nand U756 (N_756,In_145,In_626);
nor U757 (N_757,In_144,In_285);
nor U758 (N_758,In_324,In_677);
nor U759 (N_759,In_405,In_12);
nor U760 (N_760,In_303,In_119);
nor U761 (N_761,In_323,In_170);
and U762 (N_762,In_231,In_371);
nor U763 (N_763,In_624,In_261);
nor U764 (N_764,In_685,In_84);
or U765 (N_765,In_358,In_178);
and U766 (N_766,In_409,In_603);
nand U767 (N_767,In_474,In_555);
and U768 (N_768,In_570,In_49);
and U769 (N_769,In_697,In_655);
or U770 (N_770,In_64,In_199);
or U771 (N_771,In_705,In_64);
nor U772 (N_772,In_101,In_249);
and U773 (N_773,In_541,In_161);
nor U774 (N_774,In_662,In_657);
and U775 (N_775,In_659,In_693);
nor U776 (N_776,In_34,In_532);
nand U777 (N_777,In_429,In_650);
nand U778 (N_778,In_500,In_642);
nor U779 (N_779,In_122,In_656);
or U780 (N_780,In_233,In_470);
nor U781 (N_781,In_548,In_367);
and U782 (N_782,In_491,In_416);
or U783 (N_783,In_177,In_392);
and U784 (N_784,In_561,In_705);
or U785 (N_785,In_195,In_261);
nand U786 (N_786,In_414,In_676);
nand U787 (N_787,In_234,In_617);
or U788 (N_788,In_345,In_177);
and U789 (N_789,In_375,In_236);
nor U790 (N_790,In_103,In_118);
or U791 (N_791,In_382,In_327);
or U792 (N_792,In_727,In_26);
and U793 (N_793,In_125,In_324);
and U794 (N_794,In_637,In_131);
nor U795 (N_795,In_400,In_699);
and U796 (N_796,In_77,In_609);
nand U797 (N_797,In_381,In_206);
or U798 (N_798,In_692,In_607);
nand U799 (N_799,In_526,In_455);
nand U800 (N_800,In_123,In_178);
nor U801 (N_801,In_464,In_422);
or U802 (N_802,In_445,In_194);
and U803 (N_803,In_113,In_628);
nor U804 (N_804,In_613,In_423);
and U805 (N_805,In_425,In_204);
nor U806 (N_806,In_439,In_525);
nand U807 (N_807,In_639,In_51);
nand U808 (N_808,In_312,In_506);
or U809 (N_809,In_729,In_415);
or U810 (N_810,In_62,In_211);
or U811 (N_811,In_562,In_501);
or U812 (N_812,In_101,In_389);
nor U813 (N_813,In_637,In_648);
or U814 (N_814,In_153,In_308);
nor U815 (N_815,In_298,In_511);
nor U816 (N_816,In_0,In_722);
nor U817 (N_817,In_165,In_335);
nand U818 (N_818,In_674,In_5);
nor U819 (N_819,In_45,In_375);
or U820 (N_820,In_315,In_456);
nand U821 (N_821,In_430,In_166);
nor U822 (N_822,In_453,In_603);
nor U823 (N_823,In_677,In_649);
or U824 (N_824,In_361,In_542);
nand U825 (N_825,In_336,In_711);
and U826 (N_826,In_236,In_530);
or U827 (N_827,In_429,In_136);
and U828 (N_828,In_127,In_310);
or U829 (N_829,In_669,In_82);
nand U830 (N_830,In_312,In_552);
nand U831 (N_831,In_408,In_484);
or U832 (N_832,In_402,In_465);
nor U833 (N_833,In_407,In_467);
and U834 (N_834,In_54,In_479);
nor U835 (N_835,In_268,In_521);
nand U836 (N_836,In_270,In_171);
nor U837 (N_837,In_171,In_227);
or U838 (N_838,In_323,In_477);
and U839 (N_839,In_380,In_240);
nor U840 (N_840,In_275,In_223);
nand U841 (N_841,In_302,In_628);
or U842 (N_842,In_400,In_324);
nor U843 (N_843,In_727,In_157);
or U844 (N_844,In_537,In_117);
and U845 (N_845,In_275,In_40);
nor U846 (N_846,In_494,In_390);
nor U847 (N_847,In_541,In_419);
nand U848 (N_848,In_165,In_548);
and U849 (N_849,In_333,In_219);
nor U850 (N_850,In_426,In_265);
and U851 (N_851,In_417,In_663);
nor U852 (N_852,In_56,In_291);
nand U853 (N_853,In_458,In_463);
and U854 (N_854,In_170,In_528);
nor U855 (N_855,In_647,In_251);
nor U856 (N_856,In_681,In_289);
and U857 (N_857,In_97,In_736);
nand U858 (N_858,In_587,In_367);
or U859 (N_859,In_318,In_185);
nor U860 (N_860,In_335,In_56);
or U861 (N_861,In_318,In_712);
nor U862 (N_862,In_356,In_439);
and U863 (N_863,In_578,In_527);
and U864 (N_864,In_62,In_53);
nand U865 (N_865,In_114,In_587);
or U866 (N_866,In_517,In_575);
or U867 (N_867,In_577,In_584);
nor U868 (N_868,In_237,In_20);
and U869 (N_869,In_305,In_640);
nor U870 (N_870,In_639,In_83);
and U871 (N_871,In_443,In_236);
or U872 (N_872,In_616,In_491);
and U873 (N_873,In_37,In_696);
or U874 (N_874,In_530,In_40);
nor U875 (N_875,In_477,In_338);
nor U876 (N_876,In_334,In_449);
or U877 (N_877,In_663,In_629);
nand U878 (N_878,In_145,In_704);
or U879 (N_879,In_701,In_450);
or U880 (N_880,In_164,In_224);
nand U881 (N_881,In_46,In_103);
or U882 (N_882,In_216,In_733);
nand U883 (N_883,In_730,In_231);
or U884 (N_884,In_522,In_369);
or U885 (N_885,In_328,In_412);
nand U886 (N_886,In_20,In_376);
or U887 (N_887,In_641,In_477);
and U888 (N_888,In_717,In_419);
nand U889 (N_889,In_640,In_218);
nand U890 (N_890,In_146,In_10);
or U891 (N_891,In_723,In_79);
nand U892 (N_892,In_476,In_349);
nand U893 (N_893,In_359,In_296);
or U894 (N_894,In_122,In_361);
nand U895 (N_895,In_733,In_59);
nor U896 (N_896,In_158,In_268);
nand U897 (N_897,In_261,In_502);
nor U898 (N_898,In_102,In_749);
nor U899 (N_899,In_673,In_445);
or U900 (N_900,In_518,In_459);
or U901 (N_901,In_66,In_38);
nor U902 (N_902,In_46,In_270);
or U903 (N_903,In_80,In_331);
nor U904 (N_904,In_444,In_560);
or U905 (N_905,In_74,In_517);
nor U906 (N_906,In_100,In_320);
nand U907 (N_907,In_450,In_177);
or U908 (N_908,In_47,In_706);
nor U909 (N_909,In_263,In_272);
nor U910 (N_910,In_90,In_696);
nor U911 (N_911,In_410,In_139);
or U912 (N_912,In_344,In_538);
and U913 (N_913,In_434,In_659);
nand U914 (N_914,In_220,In_363);
nor U915 (N_915,In_576,In_56);
nand U916 (N_916,In_482,In_278);
and U917 (N_917,In_96,In_1);
nor U918 (N_918,In_586,In_65);
or U919 (N_919,In_81,In_276);
or U920 (N_920,In_170,In_415);
nand U921 (N_921,In_260,In_292);
nor U922 (N_922,In_660,In_410);
nor U923 (N_923,In_391,In_711);
nor U924 (N_924,In_665,In_565);
nor U925 (N_925,In_446,In_160);
and U926 (N_926,In_112,In_734);
nor U927 (N_927,In_465,In_428);
nor U928 (N_928,In_23,In_198);
and U929 (N_929,In_482,In_595);
nor U930 (N_930,In_331,In_155);
and U931 (N_931,In_328,In_181);
or U932 (N_932,In_297,In_484);
and U933 (N_933,In_705,In_595);
nor U934 (N_934,In_544,In_679);
and U935 (N_935,In_12,In_288);
and U936 (N_936,In_239,In_515);
nand U937 (N_937,In_130,In_273);
or U938 (N_938,In_153,In_643);
nor U939 (N_939,In_365,In_411);
nand U940 (N_940,In_726,In_259);
nor U941 (N_941,In_278,In_568);
nor U942 (N_942,In_336,In_392);
nor U943 (N_943,In_67,In_445);
or U944 (N_944,In_254,In_234);
and U945 (N_945,In_491,In_215);
nand U946 (N_946,In_156,In_242);
nor U947 (N_947,In_49,In_740);
nor U948 (N_948,In_186,In_462);
and U949 (N_949,In_301,In_345);
or U950 (N_950,In_84,In_159);
nand U951 (N_951,In_328,In_255);
or U952 (N_952,In_176,In_253);
and U953 (N_953,In_270,In_564);
or U954 (N_954,In_573,In_590);
and U955 (N_955,In_99,In_633);
nand U956 (N_956,In_695,In_605);
and U957 (N_957,In_732,In_589);
and U958 (N_958,In_35,In_471);
nand U959 (N_959,In_620,In_321);
nor U960 (N_960,In_69,In_741);
nand U961 (N_961,In_639,In_8);
or U962 (N_962,In_505,In_577);
or U963 (N_963,In_326,In_301);
nand U964 (N_964,In_712,In_96);
nor U965 (N_965,In_674,In_345);
or U966 (N_966,In_197,In_614);
nor U967 (N_967,In_229,In_61);
or U968 (N_968,In_662,In_626);
or U969 (N_969,In_6,In_31);
nor U970 (N_970,In_648,In_98);
nor U971 (N_971,In_506,In_475);
nand U972 (N_972,In_342,In_74);
nor U973 (N_973,In_363,In_631);
or U974 (N_974,In_504,In_34);
nand U975 (N_975,In_421,In_725);
or U976 (N_976,In_449,In_208);
and U977 (N_977,In_441,In_594);
and U978 (N_978,In_535,In_541);
nor U979 (N_979,In_247,In_290);
and U980 (N_980,In_517,In_68);
or U981 (N_981,In_590,In_194);
nor U982 (N_982,In_549,In_635);
nor U983 (N_983,In_738,In_592);
and U984 (N_984,In_554,In_349);
nor U985 (N_985,In_187,In_566);
nor U986 (N_986,In_733,In_87);
nor U987 (N_987,In_304,In_29);
or U988 (N_988,In_253,In_332);
nor U989 (N_989,In_377,In_99);
and U990 (N_990,In_424,In_15);
and U991 (N_991,In_211,In_668);
and U992 (N_992,In_502,In_61);
or U993 (N_993,In_258,In_514);
and U994 (N_994,In_329,In_205);
nor U995 (N_995,In_79,In_44);
xnor U996 (N_996,In_512,In_468);
nor U997 (N_997,In_72,In_305);
nand U998 (N_998,In_112,In_565);
nand U999 (N_999,In_448,In_475);
nand U1000 (N_1000,In_457,In_488);
nor U1001 (N_1001,In_61,In_464);
nand U1002 (N_1002,In_453,In_645);
or U1003 (N_1003,In_665,In_500);
nor U1004 (N_1004,In_28,In_329);
or U1005 (N_1005,In_173,In_495);
nor U1006 (N_1006,In_264,In_429);
and U1007 (N_1007,In_293,In_70);
and U1008 (N_1008,In_153,In_162);
and U1009 (N_1009,In_427,In_275);
or U1010 (N_1010,In_27,In_462);
nor U1011 (N_1011,In_372,In_698);
and U1012 (N_1012,In_375,In_168);
nand U1013 (N_1013,In_199,In_485);
or U1014 (N_1014,In_569,In_12);
nor U1015 (N_1015,In_711,In_688);
nor U1016 (N_1016,In_444,In_1);
or U1017 (N_1017,In_534,In_22);
or U1018 (N_1018,In_215,In_251);
nor U1019 (N_1019,In_74,In_96);
or U1020 (N_1020,In_253,In_223);
and U1021 (N_1021,In_576,In_714);
and U1022 (N_1022,In_384,In_502);
nand U1023 (N_1023,In_28,In_35);
nor U1024 (N_1024,In_597,In_539);
and U1025 (N_1025,In_7,In_86);
nand U1026 (N_1026,In_157,In_108);
and U1027 (N_1027,In_666,In_126);
nor U1028 (N_1028,In_277,In_580);
and U1029 (N_1029,In_482,In_387);
and U1030 (N_1030,In_504,In_291);
nand U1031 (N_1031,In_238,In_147);
or U1032 (N_1032,In_155,In_367);
or U1033 (N_1033,In_401,In_160);
nand U1034 (N_1034,In_208,In_606);
and U1035 (N_1035,In_733,In_256);
nand U1036 (N_1036,In_557,In_607);
and U1037 (N_1037,In_360,In_416);
nor U1038 (N_1038,In_638,In_412);
nand U1039 (N_1039,In_71,In_632);
nand U1040 (N_1040,In_527,In_599);
or U1041 (N_1041,In_239,In_575);
nor U1042 (N_1042,In_566,In_729);
nor U1043 (N_1043,In_123,In_52);
or U1044 (N_1044,In_531,In_275);
nand U1045 (N_1045,In_31,In_406);
nor U1046 (N_1046,In_239,In_32);
nor U1047 (N_1047,In_512,In_394);
or U1048 (N_1048,In_645,In_527);
xor U1049 (N_1049,In_361,In_565);
or U1050 (N_1050,In_738,In_517);
or U1051 (N_1051,In_345,In_129);
and U1052 (N_1052,In_505,In_176);
nand U1053 (N_1053,In_728,In_72);
or U1054 (N_1054,In_363,In_457);
xor U1055 (N_1055,In_332,In_624);
nand U1056 (N_1056,In_307,In_706);
nand U1057 (N_1057,In_540,In_259);
or U1058 (N_1058,In_490,In_234);
and U1059 (N_1059,In_368,In_695);
and U1060 (N_1060,In_162,In_113);
nor U1061 (N_1061,In_440,In_202);
or U1062 (N_1062,In_519,In_69);
and U1063 (N_1063,In_689,In_738);
or U1064 (N_1064,In_32,In_613);
nor U1065 (N_1065,In_422,In_506);
or U1066 (N_1066,In_299,In_674);
and U1067 (N_1067,In_414,In_418);
or U1068 (N_1068,In_623,In_114);
nor U1069 (N_1069,In_156,In_198);
and U1070 (N_1070,In_650,In_8);
and U1071 (N_1071,In_442,In_660);
and U1072 (N_1072,In_655,In_705);
nor U1073 (N_1073,In_300,In_549);
or U1074 (N_1074,In_636,In_119);
nor U1075 (N_1075,In_624,In_476);
nor U1076 (N_1076,In_649,In_246);
and U1077 (N_1077,In_390,In_32);
xnor U1078 (N_1078,In_421,In_476);
nand U1079 (N_1079,In_117,In_613);
nand U1080 (N_1080,In_376,In_3);
xnor U1081 (N_1081,In_484,In_601);
or U1082 (N_1082,In_497,In_437);
and U1083 (N_1083,In_34,In_250);
or U1084 (N_1084,In_477,In_494);
and U1085 (N_1085,In_708,In_466);
nand U1086 (N_1086,In_489,In_303);
or U1087 (N_1087,In_673,In_130);
xor U1088 (N_1088,In_717,In_441);
nor U1089 (N_1089,In_565,In_304);
and U1090 (N_1090,In_732,In_328);
or U1091 (N_1091,In_567,In_692);
nor U1092 (N_1092,In_267,In_654);
nand U1093 (N_1093,In_554,In_55);
nand U1094 (N_1094,In_417,In_387);
or U1095 (N_1095,In_513,In_46);
xnor U1096 (N_1096,In_124,In_548);
and U1097 (N_1097,In_251,In_316);
nor U1098 (N_1098,In_411,In_644);
or U1099 (N_1099,In_424,In_626);
and U1100 (N_1100,In_374,In_94);
nor U1101 (N_1101,In_613,In_427);
nand U1102 (N_1102,In_748,In_521);
and U1103 (N_1103,In_736,In_674);
nor U1104 (N_1104,In_302,In_283);
nor U1105 (N_1105,In_98,In_474);
nor U1106 (N_1106,In_490,In_719);
nor U1107 (N_1107,In_747,In_377);
or U1108 (N_1108,In_691,In_20);
nand U1109 (N_1109,In_663,In_687);
nor U1110 (N_1110,In_697,In_143);
or U1111 (N_1111,In_546,In_610);
or U1112 (N_1112,In_741,In_333);
and U1113 (N_1113,In_76,In_80);
and U1114 (N_1114,In_380,In_292);
and U1115 (N_1115,In_614,In_727);
nand U1116 (N_1116,In_157,In_189);
and U1117 (N_1117,In_84,In_10);
and U1118 (N_1118,In_249,In_248);
or U1119 (N_1119,In_480,In_448);
nand U1120 (N_1120,In_718,In_697);
and U1121 (N_1121,In_66,In_161);
or U1122 (N_1122,In_468,In_553);
nor U1123 (N_1123,In_1,In_727);
nand U1124 (N_1124,In_639,In_474);
nor U1125 (N_1125,In_599,In_544);
nand U1126 (N_1126,In_321,In_411);
or U1127 (N_1127,In_482,In_461);
nand U1128 (N_1128,In_542,In_172);
or U1129 (N_1129,In_340,In_694);
nand U1130 (N_1130,In_194,In_46);
and U1131 (N_1131,In_165,In_134);
or U1132 (N_1132,In_468,In_260);
xor U1133 (N_1133,In_180,In_207);
nor U1134 (N_1134,In_54,In_177);
nand U1135 (N_1135,In_299,In_368);
and U1136 (N_1136,In_147,In_564);
nand U1137 (N_1137,In_659,In_586);
and U1138 (N_1138,In_122,In_574);
nor U1139 (N_1139,In_173,In_515);
and U1140 (N_1140,In_61,In_276);
nor U1141 (N_1141,In_652,In_359);
nand U1142 (N_1142,In_599,In_267);
nand U1143 (N_1143,In_596,In_107);
or U1144 (N_1144,In_232,In_186);
nand U1145 (N_1145,In_708,In_341);
nor U1146 (N_1146,In_635,In_256);
and U1147 (N_1147,In_719,In_589);
or U1148 (N_1148,In_22,In_643);
or U1149 (N_1149,In_588,In_639);
nand U1150 (N_1150,In_115,In_717);
or U1151 (N_1151,In_519,In_748);
and U1152 (N_1152,In_176,In_188);
or U1153 (N_1153,In_456,In_698);
and U1154 (N_1154,In_536,In_349);
nor U1155 (N_1155,In_635,In_620);
nor U1156 (N_1156,In_178,In_281);
and U1157 (N_1157,In_293,In_449);
and U1158 (N_1158,In_159,In_46);
or U1159 (N_1159,In_555,In_449);
and U1160 (N_1160,In_175,In_710);
or U1161 (N_1161,In_595,In_82);
and U1162 (N_1162,In_84,In_359);
and U1163 (N_1163,In_417,In_689);
and U1164 (N_1164,In_97,In_249);
or U1165 (N_1165,In_48,In_230);
or U1166 (N_1166,In_343,In_529);
nand U1167 (N_1167,In_694,In_660);
nand U1168 (N_1168,In_706,In_146);
nor U1169 (N_1169,In_265,In_690);
nor U1170 (N_1170,In_260,In_481);
and U1171 (N_1171,In_464,In_45);
and U1172 (N_1172,In_28,In_538);
nor U1173 (N_1173,In_316,In_490);
and U1174 (N_1174,In_695,In_485);
nand U1175 (N_1175,In_206,In_459);
or U1176 (N_1176,In_540,In_376);
nor U1177 (N_1177,In_379,In_738);
nand U1178 (N_1178,In_729,In_119);
nand U1179 (N_1179,In_645,In_550);
or U1180 (N_1180,In_488,In_344);
nor U1181 (N_1181,In_132,In_665);
and U1182 (N_1182,In_195,In_323);
or U1183 (N_1183,In_306,In_488);
and U1184 (N_1184,In_398,In_148);
nor U1185 (N_1185,In_254,In_85);
nand U1186 (N_1186,In_95,In_265);
and U1187 (N_1187,In_518,In_420);
nor U1188 (N_1188,In_659,In_497);
and U1189 (N_1189,In_536,In_183);
nand U1190 (N_1190,In_123,In_183);
nor U1191 (N_1191,In_551,In_491);
nand U1192 (N_1192,In_228,In_350);
or U1193 (N_1193,In_62,In_19);
nand U1194 (N_1194,In_352,In_287);
nor U1195 (N_1195,In_203,In_711);
or U1196 (N_1196,In_334,In_88);
or U1197 (N_1197,In_486,In_690);
or U1198 (N_1198,In_675,In_682);
nor U1199 (N_1199,In_704,In_592);
nor U1200 (N_1200,In_482,In_303);
and U1201 (N_1201,In_535,In_620);
nand U1202 (N_1202,In_368,In_495);
and U1203 (N_1203,In_284,In_124);
nor U1204 (N_1204,In_496,In_179);
nor U1205 (N_1205,In_38,In_701);
and U1206 (N_1206,In_560,In_283);
and U1207 (N_1207,In_397,In_475);
nand U1208 (N_1208,In_248,In_719);
and U1209 (N_1209,In_38,In_210);
or U1210 (N_1210,In_26,In_111);
nor U1211 (N_1211,In_75,In_304);
nand U1212 (N_1212,In_147,In_222);
nand U1213 (N_1213,In_471,In_320);
nand U1214 (N_1214,In_229,In_94);
or U1215 (N_1215,In_105,In_398);
and U1216 (N_1216,In_269,In_155);
nand U1217 (N_1217,In_725,In_231);
nor U1218 (N_1218,In_540,In_119);
and U1219 (N_1219,In_190,In_140);
and U1220 (N_1220,In_722,In_167);
and U1221 (N_1221,In_733,In_510);
nand U1222 (N_1222,In_404,In_304);
nor U1223 (N_1223,In_700,In_354);
nand U1224 (N_1224,In_541,In_493);
and U1225 (N_1225,In_23,In_146);
nand U1226 (N_1226,In_600,In_563);
nand U1227 (N_1227,In_217,In_60);
and U1228 (N_1228,In_124,In_83);
nor U1229 (N_1229,In_11,In_341);
or U1230 (N_1230,In_244,In_199);
or U1231 (N_1231,In_631,In_257);
nor U1232 (N_1232,In_26,In_721);
or U1233 (N_1233,In_523,In_530);
and U1234 (N_1234,In_205,In_462);
nand U1235 (N_1235,In_528,In_107);
or U1236 (N_1236,In_696,In_706);
nand U1237 (N_1237,In_517,In_164);
and U1238 (N_1238,In_15,In_410);
nand U1239 (N_1239,In_82,In_678);
nor U1240 (N_1240,In_595,In_742);
nor U1241 (N_1241,In_259,In_583);
and U1242 (N_1242,In_135,In_293);
or U1243 (N_1243,In_221,In_46);
or U1244 (N_1244,In_672,In_195);
nand U1245 (N_1245,In_721,In_528);
nor U1246 (N_1246,In_80,In_388);
or U1247 (N_1247,In_591,In_140);
nor U1248 (N_1248,In_654,In_684);
nand U1249 (N_1249,In_120,In_328);
and U1250 (N_1250,In_349,In_210);
or U1251 (N_1251,In_308,In_316);
and U1252 (N_1252,In_180,In_181);
nand U1253 (N_1253,In_332,In_709);
and U1254 (N_1254,In_77,In_317);
and U1255 (N_1255,In_696,In_152);
or U1256 (N_1256,In_685,In_27);
nand U1257 (N_1257,In_0,In_90);
and U1258 (N_1258,In_391,In_748);
nand U1259 (N_1259,In_651,In_124);
nand U1260 (N_1260,In_736,In_549);
nor U1261 (N_1261,In_171,In_430);
nand U1262 (N_1262,In_416,In_409);
and U1263 (N_1263,In_196,In_37);
or U1264 (N_1264,In_546,In_575);
and U1265 (N_1265,In_620,In_655);
and U1266 (N_1266,In_425,In_521);
and U1267 (N_1267,In_498,In_678);
and U1268 (N_1268,In_112,In_724);
or U1269 (N_1269,In_677,In_659);
and U1270 (N_1270,In_554,In_697);
nor U1271 (N_1271,In_728,In_108);
and U1272 (N_1272,In_365,In_201);
and U1273 (N_1273,In_292,In_490);
or U1274 (N_1274,In_225,In_594);
nand U1275 (N_1275,In_443,In_724);
or U1276 (N_1276,In_415,In_497);
and U1277 (N_1277,In_578,In_40);
and U1278 (N_1278,In_168,In_48);
nor U1279 (N_1279,In_539,In_642);
xor U1280 (N_1280,In_697,In_126);
nand U1281 (N_1281,In_252,In_337);
nor U1282 (N_1282,In_79,In_278);
or U1283 (N_1283,In_99,In_120);
nand U1284 (N_1284,In_299,In_598);
and U1285 (N_1285,In_305,In_587);
or U1286 (N_1286,In_85,In_542);
nand U1287 (N_1287,In_744,In_582);
nor U1288 (N_1288,In_677,In_19);
nand U1289 (N_1289,In_317,In_293);
and U1290 (N_1290,In_342,In_614);
nand U1291 (N_1291,In_316,In_449);
nand U1292 (N_1292,In_58,In_609);
nor U1293 (N_1293,In_338,In_585);
nand U1294 (N_1294,In_376,In_520);
and U1295 (N_1295,In_579,In_550);
nor U1296 (N_1296,In_24,In_270);
and U1297 (N_1297,In_402,In_160);
nor U1298 (N_1298,In_313,In_573);
and U1299 (N_1299,In_254,In_511);
nor U1300 (N_1300,In_629,In_4);
nor U1301 (N_1301,In_496,In_234);
or U1302 (N_1302,In_554,In_476);
nand U1303 (N_1303,In_657,In_535);
or U1304 (N_1304,In_152,In_166);
nor U1305 (N_1305,In_197,In_271);
xor U1306 (N_1306,In_524,In_167);
nand U1307 (N_1307,In_308,In_254);
nand U1308 (N_1308,In_736,In_228);
nor U1309 (N_1309,In_431,In_721);
nor U1310 (N_1310,In_321,In_481);
or U1311 (N_1311,In_30,In_409);
nor U1312 (N_1312,In_417,In_739);
nor U1313 (N_1313,In_207,In_497);
or U1314 (N_1314,In_45,In_486);
nand U1315 (N_1315,In_241,In_228);
nor U1316 (N_1316,In_636,In_342);
and U1317 (N_1317,In_370,In_573);
nand U1318 (N_1318,In_253,In_602);
nand U1319 (N_1319,In_329,In_497);
and U1320 (N_1320,In_523,In_693);
nand U1321 (N_1321,In_577,In_416);
or U1322 (N_1322,In_682,In_619);
nand U1323 (N_1323,In_620,In_9);
and U1324 (N_1324,In_75,In_58);
nand U1325 (N_1325,In_592,In_354);
or U1326 (N_1326,In_49,In_560);
nand U1327 (N_1327,In_47,In_658);
nand U1328 (N_1328,In_567,In_749);
nand U1329 (N_1329,In_739,In_322);
nand U1330 (N_1330,In_538,In_75);
nand U1331 (N_1331,In_653,In_60);
and U1332 (N_1332,In_626,In_231);
or U1333 (N_1333,In_169,In_318);
nand U1334 (N_1334,In_742,In_55);
nor U1335 (N_1335,In_603,In_631);
nand U1336 (N_1336,In_74,In_191);
nor U1337 (N_1337,In_275,In_538);
or U1338 (N_1338,In_694,In_589);
or U1339 (N_1339,In_699,In_148);
or U1340 (N_1340,In_534,In_368);
and U1341 (N_1341,In_601,In_507);
nand U1342 (N_1342,In_113,In_222);
nor U1343 (N_1343,In_233,In_345);
nand U1344 (N_1344,In_328,In_243);
nand U1345 (N_1345,In_604,In_600);
or U1346 (N_1346,In_200,In_599);
nand U1347 (N_1347,In_370,In_665);
nor U1348 (N_1348,In_701,In_74);
nor U1349 (N_1349,In_15,In_343);
nor U1350 (N_1350,In_130,In_258);
nand U1351 (N_1351,In_11,In_433);
and U1352 (N_1352,In_45,In_179);
and U1353 (N_1353,In_457,In_713);
nor U1354 (N_1354,In_391,In_724);
nand U1355 (N_1355,In_62,In_165);
and U1356 (N_1356,In_709,In_107);
nand U1357 (N_1357,In_711,In_1);
and U1358 (N_1358,In_134,In_675);
nand U1359 (N_1359,In_68,In_175);
and U1360 (N_1360,In_237,In_645);
or U1361 (N_1361,In_117,In_583);
or U1362 (N_1362,In_685,In_22);
or U1363 (N_1363,In_18,In_335);
nor U1364 (N_1364,In_272,In_564);
nor U1365 (N_1365,In_91,In_602);
nand U1366 (N_1366,In_79,In_336);
nor U1367 (N_1367,In_579,In_204);
and U1368 (N_1368,In_57,In_497);
or U1369 (N_1369,In_440,In_401);
nor U1370 (N_1370,In_707,In_119);
or U1371 (N_1371,In_592,In_190);
nand U1372 (N_1372,In_247,In_523);
nand U1373 (N_1373,In_221,In_584);
nor U1374 (N_1374,In_123,In_728);
nand U1375 (N_1375,In_568,In_77);
and U1376 (N_1376,In_672,In_186);
nor U1377 (N_1377,In_749,In_45);
nor U1378 (N_1378,In_521,In_743);
or U1379 (N_1379,In_161,In_724);
nor U1380 (N_1380,In_556,In_113);
nor U1381 (N_1381,In_46,In_541);
nor U1382 (N_1382,In_89,In_578);
and U1383 (N_1383,In_141,In_638);
nor U1384 (N_1384,In_641,In_490);
nand U1385 (N_1385,In_99,In_740);
xnor U1386 (N_1386,In_627,In_161);
nor U1387 (N_1387,In_245,In_55);
nand U1388 (N_1388,In_183,In_580);
and U1389 (N_1389,In_441,In_98);
and U1390 (N_1390,In_61,In_360);
nand U1391 (N_1391,In_71,In_547);
nor U1392 (N_1392,In_565,In_90);
nor U1393 (N_1393,In_329,In_177);
nand U1394 (N_1394,In_630,In_728);
or U1395 (N_1395,In_724,In_433);
nand U1396 (N_1396,In_721,In_494);
or U1397 (N_1397,In_19,In_36);
nor U1398 (N_1398,In_266,In_563);
nand U1399 (N_1399,In_131,In_233);
nand U1400 (N_1400,In_673,In_691);
nand U1401 (N_1401,In_465,In_184);
and U1402 (N_1402,In_596,In_225);
nand U1403 (N_1403,In_250,In_307);
nor U1404 (N_1404,In_243,In_424);
or U1405 (N_1405,In_396,In_536);
nand U1406 (N_1406,In_475,In_491);
or U1407 (N_1407,In_136,In_641);
and U1408 (N_1408,In_678,In_106);
nand U1409 (N_1409,In_79,In_157);
or U1410 (N_1410,In_550,In_85);
or U1411 (N_1411,In_412,In_52);
nand U1412 (N_1412,In_603,In_680);
or U1413 (N_1413,In_591,In_270);
or U1414 (N_1414,In_183,In_524);
and U1415 (N_1415,In_642,In_104);
nand U1416 (N_1416,In_390,In_13);
or U1417 (N_1417,In_212,In_633);
or U1418 (N_1418,In_406,In_157);
or U1419 (N_1419,In_647,In_487);
nand U1420 (N_1420,In_586,In_460);
and U1421 (N_1421,In_348,In_240);
nor U1422 (N_1422,In_741,In_542);
and U1423 (N_1423,In_666,In_59);
and U1424 (N_1424,In_623,In_707);
nand U1425 (N_1425,In_593,In_194);
nor U1426 (N_1426,In_110,In_576);
or U1427 (N_1427,In_108,In_189);
or U1428 (N_1428,In_157,In_288);
and U1429 (N_1429,In_322,In_333);
xnor U1430 (N_1430,In_416,In_295);
and U1431 (N_1431,In_458,In_34);
and U1432 (N_1432,In_76,In_676);
nor U1433 (N_1433,In_713,In_62);
and U1434 (N_1434,In_54,In_18);
or U1435 (N_1435,In_356,In_191);
nor U1436 (N_1436,In_460,In_23);
or U1437 (N_1437,In_501,In_464);
nand U1438 (N_1438,In_362,In_155);
nor U1439 (N_1439,In_476,In_220);
nand U1440 (N_1440,In_372,In_622);
nand U1441 (N_1441,In_198,In_534);
and U1442 (N_1442,In_162,In_635);
nand U1443 (N_1443,In_617,In_417);
nor U1444 (N_1444,In_368,In_658);
nor U1445 (N_1445,In_110,In_501);
nand U1446 (N_1446,In_128,In_61);
or U1447 (N_1447,In_582,In_480);
and U1448 (N_1448,In_540,In_144);
and U1449 (N_1449,In_544,In_197);
or U1450 (N_1450,In_145,In_81);
and U1451 (N_1451,In_539,In_139);
nand U1452 (N_1452,In_550,In_267);
and U1453 (N_1453,In_502,In_493);
and U1454 (N_1454,In_387,In_497);
or U1455 (N_1455,In_352,In_693);
or U1456 (N_1456,In_642,In_142);
or U1457 (N_1457,In_588,In_333);
nor U1458 (N_1458,In_279,In_157);
and U1459 (N_1459,In_126,In_443);
or U1460 (N_1460,In_732,In_741);
and U1461 (N_1461,In_465,In_728);
nor U1462 (N_1462,In_9,In_245);
nand U1463 (N_1463,In_464,In_352);
or U1464 (N_1464,In_638,In_189);
and U1465 (N_1465,In_481,In_726);
nor U1466 (N_1466,In_160,In_145);
nor U1467 (N_1467,In_674,In_451);
nand U1468 (N_1468,In_467,In_532);
or U1469 (N_1469,In_164,In_708);
or U1470 (N_1470,In_741,In_711);
and U1471 (N_1471,In_389,In_358);
or U1472 (N_1472,In_164,In_65);
or U1473 (N_1473,In_719,In_562);
nor U1474 (N_1474,In_518,In_515);
or U1475 (N_1475,In_192,In_216);
nor U1476 (N_1476,In_684,In_21);
nor U1477 (N_1477,In_747,In_351);
nand U1478 (N_1478,In_4,In_599);
nand U1479 (N_1479,In_135,In_384);
nor U1480 (N_1480,In_412,In_379);
or U1481 (N_1481,In_213,In_68);
and U1482 (N_1482,In_120,In_736);
or U1483 (N_1483,In_186,In_419);
nand U1484 (N_1484,In_276,In_100);
or U1485 (N_1485,In_720,In_414);
and U1486 (N_1486,In_668,In_490);
and U1487 (N_1487,In_13,In_337);
and U1488 (N_1488,In_298,In_143);
nand U1489 (N_1489,In_68,In_149);
xor U1490 (N_1490,In_693,In_273);
or U1491 (N_1491,In_604,In_554);
nand U1492 (N_1492,In_409,In_432);
and U1493 (N_1493,In_308,In_259);
nor U1494 (N_1494,In_140,In_586);
or U1495 (N_1495,In_188,In_629);
or U1496 (N_1496,In_162,In_394);
and U1497 (N_1497,In_328,In_358);
nand U1498 (N_1498,In_138,In_433);
nand U1499 (N_1499,In_520,In_727);
nand U1500 (N_1500,In_239,In_20);
or U1501 (N_1501,In_713,In_10);
and U1502 (N_1502,In_677,In_351);
nand U1503 (N_1503,In_85,In_10);
or U1504 (N_1504,In_127,In_629);
nand U1505 (N_1505,In_52,In_36);
or U1506 (N_1506,In_432,In_162);
nor U1507 (N_1507,In_55,In_528);
nor U1508 (N_1508,In_110,In_56);
nor U1509 (N_1509,In_210,In_438);
nor U1510 (N_1510,In_176,In_30);
nand U1511 (N_1511,In_743,In_558);
nor U1512 (N_1512,In_5,In_141);
nor U1513 (N_1513,In_384,In_230);
and U1514 (N_1514,In_333,In_456);
nand U1515 (N_1515,In_677,In_387);
nand U1516 (N_1516,In_105,In_419);
and U1517 (N_1517,In_571,In_593);
and U1518 (N_1518,In_348,In_298);
nor U1519 (N_1519,In_79,In_674);
or U1520 (N_1520,In_741,In_409);
nor U1521 (N_1521,In_224,In_262);
and U1522 (N_1522,In_185,In_295);
or U1523 (N_1523,In_286,In_521);
nor U1524 (N_1524,In_134,In_367);
nor U1525 (N_1525,In_655,In_332);
nand U1526 (N_1526,In_733,In_552);
nor U1527 (N_1527,In_654,In_291);
nand U1528 (N_1528,In_629,In_530);
or U1529 (N_1529,In_719,In_349);
nand U1530 (N_1530,In_231,In_717);
and U1531 (N_1531,In_25,In_400);
nand U1532 (N_1532,In_576,In_335);
or U1533 (N_1533,In_717,In_531);
or U1534 (N_1534,In_586,In_519);
and U1535 (N_1535,In_112,In_695);
nand U1536 (N_1536,In_630,In_207);
xor U1537 (N_1537,In_316,In_258);
nand U1538 (N_1538,In_395,In_649);
nand U1539 (N_1539,In_203,In_517);
nand U1540 (N_1540,In_30,In_296);
nand U1541 (N_1541,In_377,In_686);
nand U1542 (N_1542,In_336,In_736);
or U1543 (N_1543,In_593,In_294);
nor U1544 (N_1544,In_362,In_673);
nand U1545 (N_1545,In_481,In_178);
or U1546 (N_1546,In_568,In_506);
nand U1547 (N_1547,In_174,In_390);
or U1548 (N_1548,In_375,In_503);
nor U1549 (N_1549,In_658,In_181);
nand U1550 (N_1550,In_426,In_707);
nand U1551 (N_1551,In_329,In_590);
or U1552 (N_1552,In_131,In_161);
nand U1553 (N_1553,In_582,In_409);
nand U1554 (N_1554,In_202,In_682);
or U1555 (N_1555,In_499,In_13);
nand U1556 (N_1556,In_579,In_591);
nand U1557 (N_1557,In_206,In_377);
or U1558 (N_1558,In_396,In_606);
nand U1559 (N_1559,In_33,In_363);
and U1560 (N_1560,In_724,In_655);
nor U1561 (N_1561,In_682,In_529);
and U1562 (N_1562,In_536,In_461);
nand U1563 (N_1563,In_728,In_204);
and U1564 (N_1564,In_391,In_566);
nand U1565 (N_1565,In_452,In_54);
nand U1566 (N_1566,In_567,In_38);
nor U1567 (N_1567,In_95,In_419);
nor U1568 (N_1568,In_200,In_171);
xor U1569 (N_1569,In_482,In_498);
nand U1570 (N_1570,In_150,In_474);
nand U1571 (N_1571,In_178,In_562);
or U1572 (N_1572,In_665,In_708);
nor U1573 (N_1573,In_552,In_35);
or U1574 (N_1574,In_365,In_65);
nand U1575 (N_1575,In_630,In_164);
nor U1576 (N_1576,In_676,In_679);
nand U1577 (N_1577,In_305,In_528);
and U1578 (N_1578,In_324,In_520);
nor U1579 (N_1579,In_108,In_215);
nand U1580 (N_1580,In_302,In_385);
and U1581 (N_1581,In_279,In_275);
nor U1582 (N_1582,In_592,In_166);
nand U1583 (N_1583,In_279,In_76);
or U1584 (N_1584,In_270,In_164);
nand U1585 (N_1585,In_161,In_556);
or U1586 (N_1586,In_307,In_220);
nor U1587 (N_1587,In_232,In_360);
nor U1588 (N_1588,In_485,In_648);
and U1589 (N_1589,In_662,In_704);
nor U1590 (N_1590,In_349,In_292);
nand U1591 (N_1591,In_361,In_510);
and U1592 (N_1592,In_85,In_429);
or U1593 (N_1593,In_131,In_322);
nor U1594 (N_1594,In_284,In_230);
and U1595 (N_1595,In_562,In_600);
nor U1596 (N_1596,In_486,In_212);
and U1597 (N_1597,In_633,In_254);
nor U1598 (N_1598,In_260,In_95);
or U1599 (N_1599,In_84,In_741);
and U1600 (N_1600,In_648,In_605);
nor U1601 (N_1601,In_376,In_374);
and U1602 (N_1602,In_411,In_526);
nor U1603 (N_1603,In_303,In_558);
and U1604 (N_1604,In_284,In_224);
and U1605 (N_1605,In_193,In_411);
and U1606 (N_1606,In_203,In_622);
and U1607 (N_1607,In_108,In_740);
nor U1608 (N_1608,In_406,In_380);
and U1609 (N_1609,In_294,In_174);
nor U1610 (N_1610,In_117,In_72);
or U1611 (N_1611,In_437,In_547);
and U1612 (N_1612,In_528,In_222);
nand U1613 (N_1613,In_126,In_542);
and U1614 (N_1614,In_636,In_500);
nor U1615 (N_1615,In_245,In_433);
or U1616 (N_1616,In_210,In_297);
nor U1617 (N_1617,In_254,In_9);
or U1618 (N_1618,In_644,In_366);
or U1619 (N_1619,In_191,In_691);
nor U1620 (N_1620,In_616,In_355);
or U1621 (N_1621,In_210,In_151);
or U1622 (N_1622,In_525,In_84);
nor U1623 (N_1623,In_685,In_629);
nor U1624 (N_1624,In_376,In_233);
or U1625 (N_1625,In_266,In_574);
and U1626 (N_1626,In_457,In_484);
and U1627 (N_1627,In_527,In_398);
nor U1628 (N_1628,In_400,In_277);
nor U1629 (N_1629,In_205,In_225);
and U1630 (N_1630,In_528,In_284);
nand U1631 (N_1631,In_328,In_563);
nor U1632 (N_1632,In_200,In_109);
nor U1633 (N_1633,In_109,In_562);
and U1634 (N_1634,In_130,In_530);
nor U1635 (N_1635,In_457,In_628);
nor U1636 (N_1636,In_46,In_19);
and U1637 (N_1637,In_57,In_237);
nand U1638 (N_1638,In_340,In_287);
and U1639 (N_1639,In_679,In_538);
or U1640 (N_1640,In_249,In_556);
or U1641 (N_1641,In_81,In_94);
and U1642 (N_1642,In_468,In_432);
or U1643 (N_1643,In_587,In_111);
and U1644 (N_1644,In_82,In_204);
and U1645 (N_1645,In_89,In_67);
xor U1646 (N_1646,In_170,In_533);
and U1647 (N_1647,In_563,In_21);
nand U1648 (N_1648,In_117,In_533);
or U1649 (N_1649,In_450,In_5);
or U1650 (N_1650,In_545,In_172);
nand U1651 (N_1651,In_624,In_236);
nand U1652 (N_1652,In_393,In_461);
or U1653 (N_1653,In_47,In_360);
nand U1654 (N_1654,In_386,In_200);
nand U1655 (N_1655,In_674,In_21);
nand U1656 (N_1656,In_127,In_618);
nor U1657 (N_1657,In_670,In_703);
or U1658 (N_1658,In_636,In_609);
and U1659 (N_1659,In_281,In_202);
nand U1660 (N_1660,In_240,In_259);
or U1661 (N_1661,In_562,In_236);
or U1662 (N_1662,In_608,In_626);
and U1663 (N_1663,In_114,In_492);
and U1664 (N_1664,In_493,In_16);
and U1665 (N_1665,In_56,In_726);
nand U1666 (N_1666,In_237,In_2);
nand U1667 (N_1667,In_127,In_347);
and U1668 (N_1668,In_710,In_480);
and U1669 (N_1669,In_380,In_166);
and U1670 (N_1670,In_257,In_305);
and U1671 (N_1671,In_378,In_695);
nor U1672 (N_1672,In_333,In_610);
nand U1673 (N_1673,In_301,In_440);
xor U1674 (N_1674,In_580,In_389);
or U1675 (N_1675,In_29,In_480);
nand U1676 (N_1676,In_20,In_414);
and U1677 (N_1677,In_74,In_726);
nand U1678 (N_1678,In_737,In_657);
and U1679 (N_1679,In_413,In_461);
and U1680 (N_1680,In_288,In_164);
and U1681 (N_1681,In_236,In_48);
or U1682 (N_1682,In_488,In_499);
nor U1683 (N_1683,In_66,In_683);
or U1684 (N_1684,In_486,In_354);
and U1685 (N_1685,In_135,In_745);
or U1686 (N_1686,In_99,In_259);
nor U1687 (N_1687,In_400,In_211);
and U1688 (N_1688,In_707,In_627);
or U1689 (N_1689,In_205,In_203);
and U1690 (N_1690,In_80,In_732);
nor U1691 (N_1691,In_282,In_430);
nand U1692 (N_1692,In_276,In_509);
nand U1693 (N_1693,In_157,In_320);
or U1694 (N_1694,In_343,In_26);
nor U1695 (N_1695,In_349,In_525);
nor U1696 (N_1696,In_635,In_647);
nor U1697 (N_1697,In_112,In_397);
or U1698 (N_1698,In_303,In_617);
and U1699 (N_1699,In_688,In_164);
nor U1700 (N_1700,In_407,In_651);
nor U1701 (N_1701,In_591,In_122);
nand U1702 (N_1702,In_649,In_209);
nand U1703 (N_1703,In_237,In_747);
and U1704 (N_1704,In_109,In_398);
nor U1705 (N_1705,In_364,In_34);
and U1706 (N_1706,In_38,In_164);
nand U1707 (N_1707,In_270,In_273);
nor U1708 (N_1708,In_42,In_366);
and U1709 (N_1709,In_638,In_679);
nand U1710 (N_1710,In_147,In_275);
nor U1711 (N_1711,In_748,In_380);
nor U1712 (N_1712,In_655,In_110);
and U1713 (N_1713,In_227,In_15);
nand U1714 (N_1714,In_740,In_515);
or U1715 (N_1715,In_126,In_665);
or U1716 (N_1716,In_267,In_360);
or U1717 (N_1717,In_434,In_656);
or U1718 (N_1718,In_229,In_658);
nor U1719 (N_1719,In_607,In_10);
and U1720 (N_1720,In_19,In_656);
nand U1721 (N_1721,In_14,In_205);
and U1722 (N_1722,In_493,In_28);
and U1723 (N_1723,In_368,In_699);
or U1724 (N_1724,In_498,In_516);
nor U1725 (N_1725,In_419,In_641);
and U1726 (N_1726,In_724,In_178);
nand U1727 (N_1727,In_374,In_669);
or U1728 (N_1728,In_288,In_250);
and U1729 (N_1729,In_308,In_662);
nor U1730 (N_1730,In_613,In_569);
or U1731 (N_1731,In_654,In_264);
nor U1732 (N_1732,In_272,In_528);
and U1733 (N_1733,In_322,In_724);
nor U1734 (N_1734,In_676,In_144);
nand U1735 (N_1735,In_530,In_35);
and U1736 (N_1736,In_295,In_323);
nand U1737 (N_1737,In_144,In_434);
nand U1738 (N_1738,In_32,In_509);
nor U1739 (N_1739,In_303,In_179);
and U1740 (N_1740,In_372,In_38);
nand U1741 (N_1741,In_555,In_430);
nand U1742 (N_1742,In_124,In_375);
and U1743 (N_1743,In_664,In_604);
or U1744 (N_1744,In_671,In_172);
nand U1745 (N_1745,In_601,In_589);
nor U1746 (N_1746,In_380,In_274);
nor U1747 (N_1747,In_592,In_342);
and U1748 (N_1748,In_411,In_611);
nor U1749 (N_1749,In_716,In_581);
nor U1750 (N_1750,In_244,In_456);
or U1751 (N_1751,In_724,In_402);
and U1752 (N_1752,In_345,In_327);
nand U1753 (N_1753,In_397,In_8);
nand U1754 (N_1754,In_239,In_706);
nor U1755 (N_1755,In_446,In_242);
nor U1756 (N_1756,In_676,In_499);
xnor U1757 (N_1757,In_437,In_224);
and U1758 (N_1758,In_516,In_124);
or U1759 (N_1759,In_85,In_500);
and U1760 (N_1760,In_720,In_133);
and U1761 (N_1761,In_216,In_398);
nor U1762 (N_1762,In_362,In_299);
xnor U1763 (N_1763,In_89,In_525);
and U1764 (N_1764,In_256,In_14);
and U1765 (N_1765,In_306,In_554);
and U1766 (N_1766,In_734,In_285);
and U1767 (N_1767,In_70,In_344);
nand U1768 (N_1768,In_439,In_196);
and U1769 (N_1769,In_539,In_86);
nand U1770 (N_1770,In_87,In_726);
nand U1771 (N_1771,In_715,In_178);
and U1772 (N_1772,In_430,In_374);
nand U1773 (N_1773,In_449,In_434);
and U1774 (N_1774,In_181,In_42);
or U1775 (N_1775,In_671,In_373);
nand U1776 (N_1776,In_572,In_223);
nand U1777 (N_1777,In_722,In_189);
or U1778 (N_1778,In_562,In_295);
nor U1779 (N_1779,In_196,In_204);
nor U1780 (N_1780,In_743,In_376);
xnor U1781 (N_1781,In_464,In_57);
and U1782 (N_1782,In_599,In_611);
nand U1783 (N_1783,In_510,In_535);
nand U1784 (N_1784,In_403,In_288);
and U1785 (N_1785,In_454,In_535);
or U1786 (N_1786,In_172,In_548);
nand U1787 (N_1787,In_403,In_137);
nor U1788 (N_1788,In_38,In_113);
nand U1789 (N_1789,In_669,In_195);
nor U1790 (N_1790,In_489,In_320);
nor U1791 (N_1791,In_216,In_291);
or U1792 (N_1792,In_250,In_274);
and U1793 (N_1793,In_275,In_247);
or U1794 (N_1794,In_468,In_124);
and U1795 (N_1795,In_266,In_424);
or U1796 (N_1796,In_415,In_734);
or U1797 (N_1797,In_384,In_458);
nand U1798 (N_1798,In_351,In_673);
and U1799 (N_1799,In_192,In_512);
nor U1800 (N_1800,In_674,In_584);
and U1801 (N_1801,In_561,In_613);
nor U1802 (N_1802,In_379,In_383);
nor U1803 (N_1803,In_362,In_371);
nor U1804 (N_1804,In_18,In_278);
and U1805 (N_1805,In_458,In_707);
or U1806 (N_1806,In_693,In_179);
nor U1807 (N_1807,In_636,In_249);
nand U1808 (N_1808,In_178,In_573);
or U1809 (N_1809,In_389,In_737);
or U1810 (N_1810,In_730,In_340);
nand U1811 (N_1811,In_127,In_563);
nor U1812 (N_1812,In_248,In_86);
or U1813 (N_1813,In_677,In_145);
nor U1814 (N_1814,In_740,In_653);
nor U1815 (N_1815,In_416,In_369);
or U1816 (N_1816,In_260,In_710);
or U1817 (N_1817,In_675,In_269);
nor U1818 (N_1818,In_113,In_206);
nor U1819 (N_1819,In_311,In_508);
nand U1820 (N_1820,In_261,In_702);
nand U1821 (N_1821,In_212,In_312);
and U1822 (N_1822,In_393,In_658);
or U1823 (N_1823,In_209,In_530);
or U1824 (N_1824,In_494,In_245);
or U1825 (N_1825,In_596,In_29);
nand U1826 (N_1826,In_598,In_342);
nor U1827 (N_1827,In_515,In_395);
nand U1828 (N_1828,In_430,In_674);
nand U1829 (N_1829,In_450,In_729);
and U1830 (N_1830,In_396,In_288);
nor U1831 (N_1831,In_102,In_724);
or U1832 (N_1832,In_489,In_592);
nand U1833 (N_1833,In_293,In_410);
nand U1834 (N_1834,In_385,In_551);
and U1835 (N_1835,In_142,In_184);
nor U1836 (N_1836,In_385,In_133);
or U1837 (N_1837,In_161,In_20);
or U1838 (N_1838,In_584,In_653);
nand U1839 (N_1839,In_279,In_139);
nand U1840 (N_1840,In_27,In_557);
or U1841 (N_1841,In_230,In_626);
nand U1842 (N_1842,In_273,In_193);
nor U1843 (N_1843,In_60,In_79);
nand U1844 (N_1844,In_592,In_695);
nand U1845 (N_1845,In_574,In_512);
nor U1846 (N_1846,In_409,In_269);
and U1847 (N_1847,In_712,In_742);
nor U1848 (N_1848,In_279,In_445);
nand U1849 (N_1849,In_347,In_459);
and U1850 (N_1850,In_65,In_14);
and U1851 (N_1851,In_548,In_637);
nor U1852 (N_1852,In_710,In_359);
and U1853 (N_1853,In_360,In_610);
nand U1854 (N_1854,In_179,In_312);
nor U1855 (N_1855,In_695,In_441);
nand U1856 (N_1856,In_324,In_232);
or U1857 (N_1857,In_225,In_715);
or U1858 (N_1858,In_252,In_295);
nand U1859 (N_1859,In_300,In_424);
and U1860 (N_1860,In_205,In_632);
nand U1861 (N_1861,In_170,In_316);
or U1862 (N_1862,In_376,In_687);
nand U1863 (N_1863,In_170,In_18);
nand U1864 (N_1864,In_4,In_693);
or U1865 (N_1865,In_142,In_277);
or U1866 (N_1866,In_186,In_456);
and U1867 (N_1867,In_74,In_280);
nand U1868 (N_1868,In_52,In_744);
nand U1869 (N_1869,In_576,In_601);
or U1870 (N_1870,In_424,In_405);
nand U1871 (N_1871,In_59,In_411);
nand U1872 (N_1872,In_230,In_727);
nor U1873 (N_1873,In_711,In_690);
or U1874 (N_1874,In_150,In_515);
nor U1875 (N_1875,In_307,In_684);
nor U1876 (N_1876,In_55,In_361);
and U1877 (N_1877,In_389,In_659);
xor U1878 (N_1878,In_411,In_475);
and U1879 (N_1879,In_60,In_336);
nor U1880 (N_1880,In_665,In_618);
and U1881 (N_1881,In_151,In_582);
nor U1882 (N_1882,In_645,In_67);
and U1883 (N_1883,In_493,In_142);
nor U1884 (N_1884,In_310,In_373);
or U1885 (N_1885,In_731,In_198);
nand U1886 (N_1886,In_550,In_233);
and U1887 (N_1887,In_452,In_217);
or U1888 (N_1888,In_644,In_208);
nor U1889 (N_1889,In_164,In_325);
nor U1890 (N_1890,In_556,In_720);
or U1891 (N_1891,In_337,In_634);
and U1892 (N_1892,In_40,In_323);
and U1893 (N_1893,In_11,In_154);
nor U1894 (N_1894,In_29,In_740);
and U1895 (N_1895,In_94,In_133);
nor U1896 (N_1896,In_547,In_334);
nand U1897 (N_1897,In_280,In_432);
nor U1898 (N_1898,In_385,In_507);
or U1899 (N_1899,In_465,In_590);
or U1900 (N_1900,In_690,In_75);
nand U1901 (N_1901,In_655,In_41);
and U1902 (N_1902,In_152,In_570);
and U1903 (N_1903,In_517,In_262);
nand U1904 (N_1904,In_154,In_167);
nand U1905 (N_1905,In_120,In_173);
nor U1906 (N_1906,In_87,In_495);
nor U1907 (N_1907,In_141,In_114);
nand U1908 (N_1908,In_84,In_287);
or U1909 (N_1909,In_370,In_50);
and U1910 (N_1910,In_645,In_583);
nand U1911 (N_1911,In_450,In_161);
or U1912 (N_1912,In_388,In_532);
or U1913 (N_1913,In_350,In_738);
and U1914 (N_1914,In_30,In_55);
and U1915 (N_1915,In_680,In_312);
nand U1916 (N_1916,In_221,In_412);
nand U1917 (N_1917,In_397,In_611);
and U1918 (N_1918,In_679,In_132);
and U1919 (N_1919,In_687,In_538);
nor U1920 (N_1920,In_459,In_263);
and U1921 (N_1921,In_521,In_343);
and U1922 (N_1922,In_673,In_157);
nor U1923 (N_1923,In_637,In_64);
nand U1924 (N_1924,In_485,In_573);
or U1925 (N_1925,In_601,In_480);
and U1926 (N_1926,In_638,In_552);
nor U1927 (N_1927,In_514,In_652);
or U1928 (N_1928,In_119,In_645);
and U1929 (N_1929,In_153,In_51);
or U1930 (N_1930,In_261,In_713);
nand U1931 (N_1931,In_718,In_651);
nand U1932 (N_1932,In_693,In_260);
and U1933 (N_1933,In_87,In_647);
nand U1934 (N_1934,In_322,In_411);
or U1935 (N_1935,In_388,In_657);
nand U1936 (N_1936,In_510,In_447);
and U1937 (N_1937,In_161,In_709);
nand U1938 (N_1938,In_503,In_58);
nor U1939 (N_1939,In_124,In_310);
nand U1940 (N_1940,In_727,In_150);
and U1941 (N_1941,In_493,In_114);
and U1942 (N_1942,In_676,In_434);
and U1943 (N_1943,In_689,In_2);
nand U1944 (N_1944,In_238,In_353);
nor U1945 (N_1945,In_122,In_311);
and U1946 (N_1946,In_512,In_542);
nor U1947 (N_1947,In_427,In_632);
nor U1948 (N_1948,In_82,In_598);
nand U1949 (N_1949,In_588,In_262);
or U1950 (N_1950,In_66,In_515);
nor U1951 (N_1951,In_224,In_357);
or U1952 (N_1952,In_715,In_294);
or U1953 (N_1953,In_278,In_272);
nand U1954 (N_1954,In_749,In_105);
nand U1955 (N_1955,In_165,In_295);
nor U1956 (N_1956,In_298,In_214);
nor U1957 (N_1957,In_152,In_223);
nor U1958 (N_1958,In_713,In_250);
nor U1959 (N_1959,In_276,In_706);
nor U1960 (N_1960,In_195,In_597);
or U1961 (N_1961,In_558,In_513);
or U1962 (N_1962,In_456,In_173);
nand U1963 (N_1963,In_505,In_278);
and U1964 (N_1964,In_708,In_253);
nor U1965 (N_1965,In_468,In_276);
or U1966 (N_1966,In_67,In_128);
nand U1967 (N_1967,In_417,In_286);
or U1968 (N_1968,In_682,In_729);
nand U1969 (N_1969,In_235,In_233);
nor U1970 (N_1970,In_195,In_80);
or U1971 (N_1971,In_266,In_284);
or U1972 (N_1972,In_500,In_7);
nand U1973 (N_1973,In_71,In_310);
or U1974 (N_1974,In_571,In_182);
and U1975 (N_1975,In_433,In_684);
or U1976 (N_1976,In_556,In_487);
nand U1977 (N_1977,In_442,In_431);
nor U1978 (N_1978,In_4,In_321);
and U1979 (N_1979,In_161,In_628);
nor U1980 (N_1980,In_465,In_601);
nor U1981 (N_1981,In_19,In_274);
nor U1982 (N_1982,In_215,In_463);
nor U1983 (N_1983,In_445,In_381);
nand U1984 (N_1984,In_82,In_375);
nor U1985 (N_1985,In_167,In_464);
and U1986 (N_1986,In_652,In_107);
or U1987 (N_1987,In_389,In_683);
nor U1988 (N_1988,In_601,In_101);
and U1989 (N_1989,In_158,In_266);
and U1990 (N_1990,In_394,In_566);
xnor U1991 (N_1991,In_473,In_450);
nand U1992 (N_1992,In_173,In_676);
nand U1993 (N_1993,In_82,In_741);
xor U1994 (N_1994,In_83,In_224);
nand U1995 (N_1995,In_318,In_262);
or U1996 (N_1996,In_715,In_468);
and U1997 (N_1997,In_90,In_229);
and U1998 (N_1998,In_92,In_339);
or U1999 (N_1999,In_339,In_634);
or U2000 (N_2000,In_288,In_384);
or U2001 (N_2001,In_12,In_258);
and U2002 (N_2002,In_360,In_414);
nand U2003 (N_2003,In_242,In_408);
nand U2004 (N_2004,In_246,In_551);
nand U2005 (N_2005,In_311,In_381);
nor U2006 (N_2006,In_501,In_16);
or U2007 (N_2007,In_590,In_657);
nand U2008 (N_2008,In_47,In_668);
nor U2009 (N_2009,In_220,In_736);
and U2010 (N_2010,In_603,In_199);
and U2011 (N_2011,In_486,In_556);
nand U2012 (N_2012,In_409,In_184);
or U2013 (N_2013,In_630,In_361);
nand U2014 (N_2014,In_636,In_535);
and U2015 (N_2015,In_30,In_128);
nor U2016 (N_2016,In_693,In_15);
and U2017 (N_2017,In_685,In_683);
and U2018 (N_2018,In_281,In_573);
and U2019 (N_2019,In_626,In_704);
nand U2020 (N_2020,In_296,In_297);
and U2021 (N_2021,In_36,In_176);
nand U2022 (N_2022,In_609,In_405);
or U2023 (N_2023,In_95,In_589);
nor U2024 (N_2024,In_727,In_348);
nand U2025 (N_2025,In_726,In_340);
and U2026 (N_2026,In_420,In_654);
and U2027 (N_2027,In_291,In_309);
nand U2028 (N_2028,In_437,In_211);
nor U2029 (N_2029,In_30,In_477);
and U2030 (N_2030,In_390,In_371);
nand U2031 (N_2031,In_716,In_334);
nand U2032 (N_2032,In_125,In_506);
nand U2033 (N_2033,In_20,In_692);
and U2034 (N_2034,In_472,In_539);
nand U2035 (N_2035,In_254,In_205);
nor U2036 (N_2036,In_126,In_328);
nand U2037 (N_2037,In_313,In_686);
nand U2038 (N_2038,In_288,In_360);
or U2039 (N_2039,In_399,In_323);
nor U2040 (N_2040,In_127,In_204);
or U2041 (N_2041,In_125,In_684);
nand U2042 (N_2042,In_116,In_688);
nand U2043 (N_2043,In_692,In_559);
and U2044 (N_2044,In_108,In_379);
nor U2045 (N_2045,In_330,In_553);
and U2046 (N_2046,In_573,In_155);
or U2047 (N_2047,In_710,In_391);
and U2048 (N_2048,In_517,In_224);
or U2049 (N_2049,In_565,In_345);
and U2050 (N_2050,In_459,In_221);
or U2051 (N_2051,In_82,In_39);
or U2052 (N_2052,In_180,In_428);
or U2053 (N_2053,In_690,In_77);
or U2054 (N_2054,In_262,In_445);
nor U2055 (N_2055,In_293,In_481);
and U2056 (N_2056,In_434,In_354);
and U2057 (N_2057,In_623,In_154);
and U2058 (N_2058,In_285,In_218);
nor U2059 (N_2059,In_259,In_88);
nand U2060 (N_2060,In_202,In_748);
and U2061 (N_2061,In_465,In_694);
and U2062 (N_2062,In_35,In_54);
and U2063 (N_2063,In_715,In_699);
nor U2064 (N_2064,In_411,In_490);
or U2065 (N_2065,In_322,In_260);
nor U2066 (N_2066,In_439,In_628);
or U2067 (N_2067,In_701,In_62);
or U2068 (N_2068,In_690,In_22);
or U2069 (N_2069,In_604,In_198);
nand U2070 (N_2070,In_709,In_10);
and U2071 (N_2071,In_3,In_280);
nor U2072 (N_2072,In_497,In_163);
or U2073 (N_2073,In_662,In_66);
nand U2074 (N_2074,In_641,In_308);
or U2075 (N_2075,In_542,In_137);
and U2076 (N_2076,In_546,In_289);
nor U2077 (N_2077,In_557,In_547);
nand U2078 (N_2078,In_22,In_305);
and U2079 (N_2079,In_498,In_739);
nand U2080 (N_2080,In_517,In_266);
and U2081 (N_2081,In_125,In_114);
and U2082 (N_2082,In_90,In_635);
nand U2083 (N_2083,In_22,In_483);
and U2084 (N_2084,In_182,In_347);
or U2085 (N_2085,In_1,In_191);
nor U2086 (N_2086,In_123,In_363);
and U2087 (N_2087,In_524,In_575);
nor U2088 (N_2088,In_236,In_528);
nor U2089 (N_2089,In_89,In_229);
nand U2090 (N_2090,In_377,In_178);
nand U2091 (N_2091,In_192,In_597);
or U2092 (N_2092,In_298,In_352);
or U2093 (N_2093,In_114,In_734);
nor U2094 (N_2094,In_90,In_447);
nand U2095 (N_2095,In_66,In_413);
and U2096 (N_2096,In_273,In_552);
nand U2097 (N_2097,In_436,In_566);
and U2098 (N_2098,In_57,In_583);
or U2099 (N_2099,In_739,In_653);
or U2100 (N_2100,In_468,In_652);
or U2101 (N_2101,In_683,In_695);
or U2102 (N_2102,In_155,In_130);
nand U2103 (N_2103,In_281,In_371);
and U2104 (N_2104,In_66,In_89);
nor U2105 (N_2105,In_236,In_68);
nor U2106 (N_2106,In_268,In_215);
nand U2107 (N_2107,In_78,In_425);
or U2108 (N_2108,In_427,In_272);
or U2109 (N_2109,In_399,In_305);
and U2110 (N_2110,In_679,In_644);
or U2111 (N_2111,In_499,In_380);
nand U2112 (N_2112,In_74,In_220);
nor U2113 (N_2113,In_536,In_747);
nor U2114 (N_2114,In_580,In_556);
or U2115 (N_2115,In_207,In_533);
nor U2116 (N_2116,In_16,In_219);
nor U2117 (N_2117,In_538,In_702);
nand U2118 (N_2118,In_541,In_131);
nor U2119 (N_2119,In_410,In_173);
or U2120 (N_2120,In_739,In_233);
and U2121 (N_2121,In_47,In_459);
or U2122 (N_2122,In_516,In_714);
nand U2123 (N_2123,In_639,In_640);
nand U2124 (N_2124,In_361,In_284);
or U2125 (N_2125,In_666,In_213);
or U2126 (N_2126,In_733,In_716);
and U2127 (N_2127,In_681,In_429);
and U2128 (N_2128,In_573,In_436);
and U2129 (N_2129,In_453,In_312);
nor U2130 (N_2130,In_95,In_117);
or U2131 (N_2131,In_194,In_200);
or U2132 (N_2132,In_675,In_64);
and U2133 (N_2133,In_487,In_720);
or U2134 (N_2134,In_139,In_9);
or U2135 (N_2135,In_433,In_428);
nand U2136 (N_2136,In_589,In_208);
nand U2137 (N_2137,In_615,In_159);
nor U2138 (N_2138,In_551,In_130);
and U2139 (N_2139,In_26,In_347);
nand U2140 (N_2140,In_432,In_396);
nor U2141 (N_2141,In_559,In_619);
nand U2142 (N_2142,In_686,In_395);
nor U2143 (N_2143,In_749,In_215);
or U2144 (N_2144,In_362,In_183);
nand U2145 (N_2145,In_163,In_510);
or U2146 (N_2146,In_616,In_48);
or U2147 (N_2147,In_27,In_601);
nand U2148 (N_2148,In_429,In_11);
nor U2149 (N_2149,In_100,In_604);
nand U2150 (N_2150,In_533,In_398);
nor U2151 (N_2151,In_184,In_54);
and U2152 (N_2152,In_81,In_221);
nand U2153 (N_2153,In_160,In_104);
nand U2154 (N_2154,In_593,In_500);
nor U2155 (N_2155,In_399,In_143);
nand U2156 (N_2156,In_466,In_560);
nand U2157 (N_2157,In_14,In_481);
nor U2158 (N_2158,In_657,In_650);
nor U2159 (N_2159,In_708,In_441);
and U2160 (N_2160,In_501,In_509);
or U2161 (N_2161,In_135,In_692);
or U2162 (N_2162,In_122,In_539);
nor U2163 (N_2163,In_571,In_73);
nor U2164 (N_2164,In_80,In_406);
nor U2165 (N_2165,In_308,In_110);
nor U2166 (N_2166,In_725,In_139);
nor U2167 (N_2167,In_387,In_723);
nand U2168 (N_2168,In_724,In_625);
nor U2169 (N_2169,In_663,In_699);
or U2170 (N_2170,In_504,In_380);
nor U2171 (N_2171,In_725,In_355);
or U2172 (N_2172,In_598,In_377);
or U2173 (N_2173,In_457,In_373);
nand U2174 (N_2174,In_203,In_598);
nand U2175 (N_2175,In_182,In_465);
nor U2176 (N_2176,In_437,In_742);
and U2177 (N_2177,In_533,In_566);
or U2178 (N_2178,In_637,In_719);
nor U2179 (N_2179,In_612,In_565);
nand U2180 (N_2180,In_24,In_314);
nor U2181 (N_2181,In_136,In_654);
nand U2182 (N_2182,In_667,In_550);
nand U2183 (N_2183,In_447,In_386);
or U2184 (N_2184,In_52,In_492);
or U2185 (N_2185,In_601,In_303);
xnor U2186 (N_2186,In_219,In_314);
and U2187 (N_2187,In_533,In_1);
nand U2188 (N_2188,In_21,In_28);
nor U2189 (N_2189,In_73,In_397);
and U2190 (N_2190,In_355,In_449);
nor U2191 (N_2191,In_55,In_105);
or U2192 (N_2192,In_503,In_4);
and U2193 (N_2193,In_722,In_486);
nor U2194 (N_2194,In_309,In_267);
and U2195 (N_2195,In_108,In_702);
and U2196 (N_2196,In_745,In_389);
nand U2197 (N_2197,In_513,In_677);
or U2198 (N_2198,In_665,In_29);
or U2199 (N_2199,In_103,In_296);
and U2200 (N_2200,In_134,In_588);
nor U2201 (N_2201,In_355,In_226);
xnor U2202 (N_2202,In_269,In_604);
or U2203 (N_2203,In_346,In_474);
nand U2204 (N_2204,In_83,In_57);
nor U2205 (N_2205,In_84,In_381);
or U2206 (N_2206,In_679,In_674);
nand U2207 (N_2207,In_419,In_573);
and U2208 (N_2208,In_408,In_641);
or U2209 (N_2209,In_17,In_435);
and U2210 (N_2210,In_102,In_84);
nor U2211 (N_2211,In_571,In_157);
and U2212 (N_2212,In_85,In_463);
nand U2213 (N_2213,In_337,In_521);
nor U2214 (N_2214,In_403,In_246);
or U2215 (N_2215,In_14,In_553);
or U2216 (N_2216,In_473,In_501);
or U2217 (N_2217,In_455,In_195);
and U2218 (N_2218,In_581,In_39);
nand U2219 (N_2219,In_517,In_377);
or U2220 (N_2220,In_101,In_647);
and U2221 (N_2221,In_695,In_722);
nor U2222 (N_2222,In_656,In_438);
or U2223 (N_2223,In_328,In_159);
and U2224 (N_2224,In_82,In_433);
and U2225 (N_2225,In_284,In_107);
xor U2226 (N_2226,In_273,In_86);
and U2227 (N_2227,In_542,In_701);
nand U2228 (N_2228,In_514,In_598);
or U2229 (N_2229,In_293,In_43);
or U2230 (N_2230,In_178,In_23);
nor U2231 (N_2231,In_609,In_104);
nor U2232 (N_2232,In_330,In_537);
nand U2233 (N_2233,In_285,In_636);
and U2234 (N_2234,In_393,In_80);
nor U2235 (N_2235,In_68,In_375);
and U2236 (N_2236,In_484,In_541);
nor U2237 (N_2237,In_484,In_453);
and U2238 (N_2238,In_122,In_524);
nor U2239 (N_2239,In_120,In_749);
nor U2240 (N_2240,In_559,In_338);
and U2241 (N_2241,In_139,In_382);
nor U2242 (N_2242,In_338,In_286);
nand U2243 (N_2243,In_342,In_291);
nor U2244 (N_2244,In_301,In_404);
nor U2245 (N_2245,In_481,In_199);
nand U2246 (N_2246,In_739,In_525);
or U2247 (N_2247,In_551,In_122);
nand U2248 (N_2248,In_24,In_385);
nand U2249 (N_2249,In_264,In_569);
and U2250 (N_2250,In_739,In_415);
and U2251 (N_2251,In_459,In_29);
nor U2252 (N_2252,In_546,In_168);
and U2253 (N_2253,In_647,In_581);
or U2254 (N_2254,In_509,In_283);
and U2255 (N_2255,In_666,In_530);
or U2256 (N_2256,In_173,In_433);
or U2257 (N_2257,In_654,In_372);
or U2258 (N_2258,In_721,In_700);
and U2259 (N_2259,In_65,In_73);
nand U2260 (N_2260,In_0,In_684);
nor U2261 (N_2261,In_615,In_598);
and U2262 (N_2262,In_269,In_458);
nand U2263 (N_2263,In_396,In_274);
or U2264 (N_2264,In_142,In_469);
and U2265 (N_2265,In_8,In_138);
nand U2266 (N_2266,In_438,In_321);
nand U2267 (N_2267,In_468,In_376);
nor U2268 (N_2268,In_142,In_408);
and U2269 (N_2269,In_358,In_543);
or U2270 (N_2270,In_88,In_211);
nand U2271 (N_2271,In_585,In_75);
and U2272 (N_2272,In_685,In_67);
and U2273 (N_2273,In_594,In_158);
nand U2274 (N_2274,In_54,In_458);
and U2275 (N_2275,In_472,In_392);
or U2276 (N_2276,In_34,In_520);
nor U2277 (N_2277,In_545,In_101);
and U2278 (N_2278,In_585,In_188);
and U2279 (N_2279,In_129,In_654);
nor U2280 (N_2280,In_663,In_591);
and U2281 (N_2281,In_719,In_609);
nand U2282 (N_2282,In_715,In_165);
or U2283 (N_2283,In_663,In_371);
or U2284 (N_2284,In_600,In_298);
or U2285 (N_2285,In_448,In_526);
and U2286 (N_2286,In_294,In_646);
nand U2287 (N_2287,In_36,In_579);
nor U2288 (N_2288,In_60,In_738);
or U2289 (N_2289,In_42,In_242);
nand U2290 (N_2290,In_473,In_317);
nand U2291 (N_2291,In_193,In_23);
and U2292 (N_2292,In_2,In_478);
nor U2293 (N_2293,In_152,In_92);
nor U2294 (N_2294,In_94,In_407);
nor U2295 (N_2295,In_716,In_46);
and U2296 (N_2296,In_330,In_414);
nor U2297 (N_2297,In_395,In_451);
or U2298 (N_2298,In_228,In_661);
nor U2299 (N_2299,In_455,In_232);
nor U2300 (N_2300,In_484,In_640);
and U2301 (N_2301,In_347,In_437);
nor U2302 (N_2302,In_307,In_523);
nor U2303 (N_2303,In_724,In_651);
and U2304 (N_2304,In_95,In_133);
and U2305 (N_2305,In_362,In_161);
nand U2306 (N_2306,In_641,In_91);
or U2307 (N_2307,In_586,In_257);
and U2308 (N_2308,In_461,In_483);
or U2309 (N_2309,In_65,In_158);
nand U2310 (N_2310,In_20,In_54);
and U2311 (N_2311,In_2,In_275);
or U2312 (N_2312,In_88,In_33);
nand U2313 (N_2313,In_217,In_39);
nor U2314 (N_2314,In_714,In_59);
or U2315 (N_2315,In_635,In_452);
and U2316 (N_2316,In_566,In_368);
nand U2317 (N_2317,In_120,In_449);
nor U2318 (N_2318,In_731,In_240);
and U2319 (N_2319,In_688,In_395);
nand U2320 (N_2320,In_296,In_639);
nor U2321 (N_2321,In_726,In_11);
nand U2322 (N_2322,In_562,In_438);
nor U2323 (N_2323,In_114,In_620);
nor U2324 (N_2324,In_713,In_116);
and U2325 (N_2325,In_308,In_712);
nor U2326 (N_2326,In_201,In_357);
and U2327 (N_2327,In_579,In_217);
and U2328 (N_2328,In_588,In_708);
nand U2329 (N_2329,In_683,In_433);
nand U2330 (N_2330,In_445,In_149);
nor U2331 (N_2331,In_422,In_72);
or U2332 (N_2332,In_44,In_377);
and U2333 (N_2333,In_213,In_497);
and U2334 (N_2334,In_245,In_516);
nand U2335 (N_2335,In_722,In_609);
or U2336 (N_2336,In_626,In_42);
or U2337 (N_2337,In_728,In_65);
nand U2338 (N_2338,In_461,In_367);
or U2339 (N_2339,In_656,In_76);
xnor U2340 (N_2340,In_132,In_489);
nor U2341 (N_2341,In_156,In_216);
or U2342 (N_2342,In_413,In_422);
or U2343 (N_2343,In_730,In_64);
and U2344 (N_2344,In_291,In_571);
and U2345 (N_2345,In_251,In_10);
and U2346 (N_2346,In_543,In_380);
nand U2347 (N_2347,In_277,In_267);
and U2348 (N_2348,In_376,In_49);
or U2349 (N_2349,In_151,In_526);
or U2350 (N_2350,In_599,In_609);
and U2351 (N_2351,In_282,In_596);
nor U2352 (N_2352,In_282,In_128);
nor U2353 (N_2353,In_358,In_50);
nor U2354 (N_2354,In_555,In_454);
nand U2355 (N_2355,In_522,In_188);
nand U2356 (N_2356,In_83,In_34);
nand U2357 (N_2357,In_729,In_511);
or U2358 (N_2358,In_486,In_134);
nand U2359 (N_2359,In_522,In_371);
and U2360 (N_2360,In_423,In_552);
or U2361 (N_2361,In_92,In_558);
nand U2362 (N_2362,In_0,In_667);
or U2363 (N_2363,In_345,In_156);
and U2364 (N_2364,In_725,In_719);
or U2365 (N_2365,In_568,In_545);
or U2366 (N_2366,In_111,In_554);
or U2367 (N_2367,In_320,In_113);
or U2368 (N_2368,In_15,In_163);
and U2369 (N_2369,In_516,In_276);
nor U2370 (N_2370,In_250,In_607);
nand U2371 (N_2371,In_409,In_423);
nor U2372 (N_2372,In_139,In_480);
nor U2373 (N_2373,In_489,In_156);
nor U2374 (N_2374,In_609,In_533);
nor U2375 (N_2375,In_449,In_614);
nor U2376 (N_2376,In_197,In_590);
nand U2377 (N_2377,In_57,In_591);
nand U2378 (N_2378,In_552,In_538);
nand U2379 (N_2379,In_448,In_609);
and U2380 (N_2380,In_279,In_691);
or U2381 (N_2381,In_608,In_471);
nand U2382 (N_2382,In_18,In_532);
nand U2383 (N_2383,In_708,In_46);
nand U2384 (N_2384,In_120,In_542);
nand U2385 (N_2385,In_368,In_581);
xor U2386 (N_2386,In_541,In_236);
and U2387 (N_2387,In_205,In_180);
or U2388 (N_2388,In_411,In_221);
nor U2389 (N_2389,In_283,In_23);
nand U2390 (N_2390,In_468,In_474);
and U2391 (N_2391,In_133,In_521);
nand U2392 (N_2392,In_402,In_588);
nor U2393 (N_2393,In_49,In_161);
and U2394 (N_2394,In_571,In_253);
and U2395 (N_2395,In_610,In_666);
or U2396 (N_2396,In_110,In_746);
nor U2397 (N_2397,In_313,In_702);
nor U2398 (N_2398,In_383,In_403);
or U2399 (N_2399,In_351,In_81);
or U2400 (N_2400,In_238,In_3);
or U2401 (N_2401,In_631,In_83);
or U2402 (N_2402,In_549,In_202);
or U2403 (N_2403,In_479,In_747);
nor U2404 (N_2404,In_267,In_291);
nor U2405 (N_2405,In_95,In_68);
nor U2406 (N_2406,In_209,In_299);
and U2407 (N_2407,In_232,In_727);
or U2408 (N_2408,In_708,In_447);
and U2409 (N_2409,In_261,In_95);
or U2410 (N_2410,In_668,In_692);
nand U2411 (N_2411,In_482,In_379);
nor U2412 (N_2412,In_157,In_253);
or U2413 (N_2413,In_746,In_50);
nor U2414 (N_2414,In_45,In_524);
nor U2415 (N_2415,In_673,In_35);
or U2416 (N_2416,In_700,In_392);
xor U2417 (N_2417,In_464,In_685);
nor U2418 (N_2418,In_426,In_27);
nand U2419 (N_2419,In_522,In_16);
or U2420 (N_2420,In_146,In_47);
nor U2421 (N_2421,In_428,In_199);
or U2422 (N_2422,In_509,In_714);
and U2423 (N_2423,In_138,In_636);
nor U2424 (N_2424,In_351,In_511);
or U2425 (N_2425,In_372,In_689);
or U2426 (N_2426,In_210,In_411);
xor U2427 (N_2427,In_543,In_334);
nor U2428 (N_2428,In_346,In_250);
xnor U2429 (N_2429,In_682,In_361);
nor U2430 (N_2430,In_445,In_739);
or U2431 (N_2431,In_341,In_212);
nor U2432 (N_2432,In_483,In_651);
nor U2433 (N_2433,In_605,In_536);
and U2434 (N_2434,In_60,In_737);
nand U2435 (N_2435,In_89,In_157);
and U2436 (N_2436,In_651,In_97);
nor U2437 (N_2437,In_570,In_400);
and U2438 (N_2438,In_641,In_464);
or U2439 (N_2439,In_518,In_432);
nand U2440 (N_2440,In_268,In_652);
or U2441 (N_2441,In_129,In_158);
nand U2442 (N_2442,In_396,In_213);
nand U2443 (N_2443,In_14,In_212);
nand U2444 (N_2444,In_185,In_144);
xor U2445 (N_2445,In_56,In_288);
nor U2446 (N_2446,In_91,In_716);
nand U2447 (N_2447,In_17,In_419);
and U2448 (N_2448,In_446,In_665);
and U2449 (N_2449,In_164,In_682);
nand U2450 (N_2450,In_632,In_77);
nand U2451 (N_2451,In_551,In_284);
or U2452 (N_2452,In_400,In_299);
nor U2453 (N_2453,In_276,In_125);
nor U2454 (N_2454,In_525,In_389);
nand U2455 (N_2455,In_152,In_630);
or U2456 (N_2456,In_67,In_169);
or U2457 (N_2457,In_499,In_535);
nand U2458 (N_2458,In_411,In_78);
or U2459 (N_2459,In_707,In_347);
nor U2460 (N_2460,In_160,In_517);
nor U2461 (N_2461,In_718,In_72);
and U2462 (N_2462,In_729,In_338);
or U2463 (N_2463,In_95,In_136);
nor U2464 (N_2464,In_13,In_82);
nor U2465 (N_2465,In_96,In_260);
nor U2466 (N_2466,In_392,In_522);
nand U2467 (N_2467,In_718,In_748);
or U2468 (N_2468,In_573,In_138);
nor U2469 (N_2469,In_186,In_106);
or U2470 (N_2470,In_84,In_75);
or U2471 (N_2471,In_273,In_45);
nand U2472 (N_2472,In_388,In_287);
or U2473 (N_2473,In_135,In_576);
nor U2474 (N_2474,In_424,In_108);
and U2475 (N_2475,In_103,In_330);
or U2476 (N_2476,In_514,In_140);
or U2477 (N_2477,In_188,In_391);
nand U2478 (N_2478,In_585,In_14);
nand U2479 (N_2479,In_747,In_180);
or U2480 (N_2480,In_261,In_654);
nand U2481 (N_2481,In_234,In_189);
or U2482 (N_2482,In_494,In_351);
or U2483 (N_2483,In_706,In_127);
nand U2484 (N_2484,In_483,In_700);
nor U2485 (N_2485,In_420,In_628);
or U2486 (N_2486,In_668,In_437);
nor U2487 (N_2487,In_140,In_101);
or U2488 (N_2488,In_684,In_34);
nand U2489 (N_2489,In_299,In_487);
or U2490 (N_2490,In_177,In_648);
and U2491 (N_2491,In_457,In_587);
or U2492 (N_2492,In_592,In_27);
nand U2493 (N_2493,In_242,In_170);
nand U2494 (N_2494,In_123,In_591);
nor U2495 (N_2495,In_657,In_542);
nor U2496 (N_2496,In_720,In_113);
or U2497 (N_2497,In_630,In_535);
or U2498 (N_2498,In_112,In_551);
and U2499 (N_2499,In_472,In_559);
and U2500 (N_2500,N_376,N_2469);
and U2501 (N_2501,N_218,N_698);
or U2502 (N_2502,N_295,N_236);
and U2503 (N_2503,N_1776,N_597);
nand U2504 (N_2504,N_1399,N_2483);
or U2505 (N_2505,N_2373,N_9);
nor U2506 (N_2506,N_1611,N_2247);
nand U2507 (N_2507,N_503,N_2147);
nor U2508 (N_2508,N_851,N_1267);
and U2509 (N_2509,N_1457,N_1720);
or U2510 (N_2510,N_1264,N_379);
nor U2511 (N_2511,N_2108,N_2401);
nand U2512 (N_2512,N_2279,N_1243);
and U2513 (N_2513,N_791,N_1225);
or U2514 (N_2514,N_1578,N_2417);
nand U2515 (N_2515,N_1566,N_373);
or U2516 (N_2516,N_102,N_2257);
nand U2517 (N_2517,N_30,N_1051);
nor U2518 (N_2518,N_954,N_2087);
nor U2519 (N_2519,N_1966,N_2062);
nand U2520 (N_2520,N_2213,N_43);
nor U2521 (N_2521,N_1734,N_465);
nor U2522 (N_2522,N_1618,N_1178);
nor U2523 (N_2523,N_1534,N_1949);
or U2524 (N_2524,N_1275,N_1749);
or U2525 (N_2525,N_805,N_1510);
nor U2526 (N_2526,N_470,N_1222);
nor U2527 (N_2527,N_1440,N_456);
and U2528 (N_2528,N_2329,N_1011);
or U2529 (N_2529,N_1296,N_1960);
or U2530 (N_2530,N_1147,N_2333);
nand U2531 (N_2531,N_1093,N_1013);
or U2532 (N_2532,N_2038,N_2080);
xor U2533 (N_2533,N_335,N_1294);
nor U2534 (N_2534,N_63,N_1366);
and U2535 (N_2535,N_2015,N_2260);
nand U2536 (N_2536,N_2176,N_427);
nor U2537 (N_2537,N_2236,N_1560);
xnor U2538 (N_2538,N_23,N_765);
nand U2539 (N_2539,N_641,N_1829);
nand U2540 (N_2540,N_1281,N_1493);
nor U2541 (N_2541,N_919,N_88);
nand U2542 (N_2542,N_561,N_1922);
nor U2543 (N_2543,N_254,N_2351);
nand U2544 (N_2544,N_200,N_1079);
or U2545 (N_2545,N_1809,N_1754);
or U2546 (N_2546,N_211,N_2061);
and U2547 (N_2547,N_1814,N_1488);
nor U2548 (N_2548,N_183,N_1811);
or U2549 (N_2549,N_2241,N_408);
nor U2550 (N_2550,N_391,N_2453);
nand U2551 (N_2551,N_1165,N_125);
nor U2552 (N_2552,N_595,N_1444);
or U2553 (N_2553,N_1634,N_1047);
or U2554 (N_2554,N_915,N_545);
and U2555 (N_2555,N_1956,N_1072);
and U2556 (N_2556,N_725,N_1097);
and U2557 (N_2557,N_126,N_823);
nand U2558 (N_2558,N_1610,N_1442);
nor U2559 (N_2559,N_1102,N_1323);
nor U2560 (N_2560,N_850,N_913);
nand U2561 (N_2561,N_2227,N_675);
nor U2562 (N_2562,N_1141,N_1739);
nand U2563 (N_2563,N_2299,N_885);
and U2564 (N_2564,N_318,N_1827);
or U2565 (N_2565,N_2078,N_1530);
nor U2566 (N_2566,N_681,N_941);
nand U2567 (N_2567,N_1128,N_238);
nor U2568 (N_2568,N_294,N_2394);
and U2569 (N_2569,N_1825,N_1792);
and U2570 (N_2570,N_1240,N_2322);
and U2571 (N_2571,N_600,N_161);
nand U2572 (N_2572,N_2271,N_1631);
or U2573 (N_2573,N_1887,N_2146);
nor U2574 (N_2574,N_644,N_1723);
or U2575 (N_2575,N_2337,N_1398);
nand U2576 (N_2576,N_1682,N_1726);
nor U2577 (N_2577,N_1220,N_1637);
nand U2578 (N_2578,N_627,N_1121);
or U2579 (N_2579,N_235,N_1248);
nand U2580 (N_2580,N_889,N_1905);
nand U2581 (N_2581,N_2250,N_224);
nor U2582 (N_2582,N_1623,N_193);
and U2583 (N_2583,N_1049,N_2255);
or U2584 (N_2584,N_769,N_744);
or U2585 (N_2585,N_2452,N_486);
or U2586 (N_2586,N_60,N_2274);
or U2587 (N_2587,N_479,N_1095);
nor U2588 (N_2588,N_735,N_970);
or U2589 (N_2589,N_2419,N_20);
or U2590 (N_2590,N_383,N_1064);
nand U2591 (N_2591,N_279,N_421);
and U2592 (N_2592,N_336,N_369);
and U2593 (N_2593,N_50,N_1235);
nor U2594 (N_2594,N_2184,N_2223);
or U2595 (N_2595,N_59,N_655);
or U2596 (N_2596,N_149,N_1461);
nand U2597 (N_2597,N_1777,N_1783);
and U2598 (N_2598,N_782,N_340);
xor U2599 (N_2599,N_273,N_1098);
or U2600 (N_2600,N_801,N_2211);
or U2601 (N_2601,N_718,N_1718);
nor U2602 (N_2602,N_1940,N_720);
nor U2603 (N_2603,N_1443,N_1840);
nand U2604 (N_2604,N_1210,N_1632);
nor U2605 (N_2605,N_1062,N_1801);
and U2606 (N_2606,N_1424,N_819);
nand U2607 (N_2607,N_118,N_35);
nand U2608 (N_2608,N_972,N_1429);
nor U2609 (N_2609,N_1286,N_83);
nand U2610 (N_2610,N_745,N_2066);
xnor U2611 (N_2611,N_2347,N_2064);
nor U2612 (N_2612,N_438,N_308);
nor U2613 (N_2613,N_99,N_1375);
nor U2614 (N_2614,N_1498,N_1885);
nand U2615 (N_2615,N_300,N_1168);
or U2616 (N_2616,N_420,N_522);
and U2617 (N_2617,N_1224,N_122);
nand U2618 (N_2618,N_1755,N_1061);
nor U2619 (N_2619,N_2306,N_394);
and U2620 (N_2620,N_1668,N_1545);
nor U2621 (N_2621,N_800,N_1138);
or U2622 (N_2622,N_616,N_808);
nand U2623 (N_2623,N_1988,N_743);
nand U2624 (N_2624,N_239,N_2043);
and U2625 (N_2625,N_1023,N_2293);
nand U2626 (N_2626,N_1149,N_1687);
nor U2627 (N_2627,N_906,N_528);
and U2628 (N_2628,N_1336,N_1886);
nand U2629 (N_2629,N_1343,N_966);
or U2630 (N_2630,N_2242,N_943);
nand U2631 (N_2631,N_480,N_724);
and U2632 (N_2632,N_1122,N_554);
nand U2633 (N_2633,N_843,N_2178);
nor U2634 (N_2634,N_2138,N_275);
and U2635 (N_2635,N_794,N_1470);
or U2636 (N_2636,N_1549,N_1181);
nor U2637 (N_2637,N_414,N_1691);
nand U2638 (N_2638,N_1502,N_1215);
nor U2639 (N_2639,N_1474,N_307);
and U2640 (N_2640,N_2130,N_1939);
nand U2641 (N_2641,N_1743,N_2209);
nor U2642 (N_2642,N_1028,N_2323);
nor U2643 (N_2643,N_305,N_1480);
and U2644 (N_2644,N_1793,N_1692);
and U2645 (N_2645,N_1035,N_2234);
nand U2646 (N_2646,N_136,N_1009);
or U2647 (N_2647,N_75,N_1606);
xnor U2648 (N_2648,N_1347,N_276);
and U2649 (N_2649,N_2370,N_1937);
or U2650 (N_2650,N_1857,N_1781);
and U2651 (N_2651,N_260,N_19);
and U2652 (N_2652,N_2177,N_291);
nand U2653 (N_2653,N_1362,N_2238);
nor U2654 (N_2654,N_678,N_581);
or U2655 (N_2655,N_527,N_34);
and U2656 (N_2656,N_304,N_731);
xnor U2657 (N_2657,N_1308,N_1889);
or U2658 (N_2658,N_1931,N_1831);
or U2659 (N_2659,N_1383,N_609);
or U2660 (N_2660,N_2189,N_497);
and U2661 (N_2661,N_1033,N_1305);
xnor U2662 (N_2662,N_213,N_2326);
or U2663 (N_2663,N_980,N_1561);
nor U2664 (N_2664,N_810,N_1499);
nand U2665 (N_2665,N_1242,N_1883);
nand U2666 (N_2666,N_1678,N_194);
or U2667 (N_2667,N_2024,N_2450);
or U2668 (N_2668,N_952,N_706);
or U2669 (N_2669,N_1202,N_1650);
or U2670 (N_2670,N_1538,N_2389);
nand U2671 (N_2671,N_1293,N_1869);
or U2672 (N_2672,N_1915,N_778);
nor U2673 (N_2673,N_2208,N_483);
nor U2674 (N_2674,N_338,N_1845);
nor U2675 (N_2675,N_2127,N_2346);
xnor U2676 (N_2676,N_1920,N_1213);
and U2677 (N_2677,N_1559,N_2265);
or U2678 (N_2678,N_2449,N_494);
and U2679 (N_2679,N_297,N_1015);
xor U2680 (N_2680,N_385,N_790);
or U2681 (N_2681,N_1688,N_2245);
xor U2682 (N_2682,N_2280,N_842);
nand U2683 (N_2683,N_2479,N_2133);
or U2684 (N_2684,N_968,N_1856);
xor U2685 (N_2685,N_2153,N_1891);
nand U2686 (N_2686,N_3,N_74);
nand U2687 (N_2687,N_1640,N_64);
nand U2688 (N_2688,N_1513,N_371);
nand U2689 (N_2689,N_2020,N_1415);
nor U2690 (N_2690,N_57,N_84);
or U2691 (N_2691,N_645,N_799);
nor U2692 (N_2692,N_2399,N_729);
and U2693 (N_2693,N_524,N_1842);
nand U2694 (N_2694,N_631,N_855);
or U2695 (N_2695,N_667,N_1875);
nor U2696 (N_2696,N_1106,N_1802);
or U2697 (N_2697,N_1914,N_2287);
nand U2698 (N_2698,N_253,N_1170);
nor U2699 (N_2699,N_2413,N_424);
nand U2700 (N_2700,N_197,N_1164);
nand U2701 (N_2701,N_339,N_1198);
and U2702 (N_2702,N_478,N_2438);
nand U2703 (N_2703,N_2318,N_1974);
nand U2704 (N_2704,N_432,N_848);
nor U2705 (N_2705,N_2458,N_47);
nor U2706 (N_2706,N_1604,N_500);
and U2707 (N_2707,N_257,N_1785);
and U2708 (N_2708,N_1774,N_1896);
or U2709 (N_2709,N_1773,N_1854);
or U2710 (N_2710,N_2217,N_1277);
and U2711 (N_2711,N_484,N_632);
nor U2712 (N_2712,N_1467,N_159);
or U2713 (N_2713,N_2140,N_1395);
nand U2714 (N_2714,N_1163,N_1975);
or U2715 (N_2715,N_2385,N_1420);
or U2716 (N_2716,N_891,N_2122);
nand U2717 (N_2717,N_113,N_490);
nand U2718 (N_2718,N_415,N_1481);
or U2719 (N_2719,N_1259,N_2277);
nor U2720 (N_2720,N_455,N_1083);
nor U2721 (N_2721,N_180,N_608);
and U2722 (N_2722,N_162,N_1263);
nor U2723 (N_2723,N_1482,N_961);
and U2724 (N_2724,N_2447,N_1673);
nand U2725 (N_2725,N_2395,N_271);
and U2726 (N_2726,N_986,N_523);
and U2727 (N_2727,N_2074,N_2120);
or U2728 (N_2728,N_2044,N_911);
nor U2729 (N_2729,N_418,N_2484);
nor U2730 (N_2730,N_2405,N_2065);
nand U2731 (N_2731,N_1309,N_2359);
and U2732 (N_2732,N_18,N_775);
nor U2733 (N_2733,N_1600,N_1594);
and U2734 (N_2734,N_1616,N_2488);
nand U2735 (N_2735,N_158,N_298);
and U2736 (N_2736,N_1455,N_1929);
and U2737 (N_2737,N_142,N_838);
or U2738 (N_2738,N_2009,N_959);
nor U2739 (N_2739,N_1888,N_1719);
and U2740 (N_2740,N_2056,N_502);
or U2741 (N_2741,N_894,N_240);
nor U2742 (N_2742,N_1821,N_1663);
or U2743 (N_2743,N_2314,N_1676);
nor U2744 (N_2744,N_2124,N_137);
nand U2745 (N_2745,N_825,N_1464);
and U2746 (N_2746,N_929,N_1058);
or U2747 (N_2747,N_1377,N_1855);
nand U2748 (N_2748,N_1982,N_732);
nor U2749 (N_2749,N_127,N_449);
nor U2750 (N_2750,N_1471,N_649);
or U2751 (N_2751,N_1846,N_560);
or U2752 (N_2752,N_314,N_1318);
and U2753 (N_2753,N_1588,N_1491);
nand U2754 (N_2754,N_2243,N_2426);
nor U2755 (N_2755,N_1830,N_2069);
and U2756 (N_2756,N_873,N_2305);
nand U2757 (N_2757,N_1119,N_2186);
and U2758 (N_2758,N_1331,N_1867);
or U2759 (N_2759,N_967,N_989);
or U2760 (N_2760,N_1782,N_835);
or U2761 (N_2761,N_826,N_256);
or U2762 (N_2762,N_387,N_100);
nand U2763 (N_2763,N_2276,N_1237);
nand U2764 (N_2764,N_2028,N_2202);
and U2765 (N_2765,N_2349,N_343);
nor U2766 (N_2766,N_673,N_2266);
and U2767 (N_2767,N_1099,N_936);
nand U2768 (N_2768,N_987,N_2170);
or U2769 (N_2769,N_766,N_199);
or U2770 (N_2770,N_2014,N_1298);
nor U2771 (N_2771,N_1657,N_144);
nand U2772 (N_2772,N_1463,N_2156);
nor U2773 (N_2773,N_365,N_507);
nor U2774 (N_2774,N_1849,N_1156);
nand U2775 (N_2775,N_1112,N_606);
nand U2776 (N_2776,N_772,N_1570);
or U2777 (N_2777,N_1451,N_1134);
nor U2778 (N_2778,N_1936,N_1189);
nor U2779 (N_2779,N_901,N_2088);
nand U2780 (N_2780,N_1828,N_2248);
nor U2781 (N_2781,N_1086,N_1052);
and U2782 (N_2782,N_2075,N_1357);
nand U2783 (N_2783,N_2407,N_2475);
nand U2784 (N_2784,N_173,N_388);
and U2785 (N_2785,N_883,N_1492);
nor U2786 (N_2786,N_2316,N_53);
and U2787 (N_2787,N_82,N_405);
or U2788 (N_2788,N_2461,N_1658);
nor U2789 (N_2789,N_374,N_979);
nor U2790 (N_2790,N_1786,N_2391);
nor U2791 (N_2791,N_2165,N_512);
nand U2792 (N_2792,N_1656,N_730);
nor U2793 (N_2793,N_2376,N_2378);
and U2794 (N_2794,N_2083,N_1667);
and U2795 (N_2795,N_1812,N_1662);
and U2796 (N_2796,N_313,N_111);
and U2797 (N_2797,N_402,N_2112);
and U2798 (N_2798,N_1185,N_1008);
or U2799 (N_2799,N_68,N_1322);
nor U2800 (N_2800,N_133,N_1154);
and U2801 (N_2801,N_1567,N_1535);
nor U2802 (N_2802,N_1552,N_1972);
nand U2803 (N_2803,N_764,N_1496);
and U2804 (N_2804,N_328,N_624);
nor U2805 (N_2805,N_139,N_1543);
nor U2806 (N_2806,N_822,N_2336);
and U2807 (N_2807,N_441,N_1495);
or U2808 (N_2808,N_1234,N_1071);
and U2809 (N_2809,N_106,N_1020);
nor U2810 (N_2810,N_853,N_1878);
or U2811 (N_2811,N_2442,N_531);
and U2812 (N_2812,N_400,N_1577);
nor U2813 (N_2813,N_1026,N_114);
nand U2814 (N_2814,N_2012,N_1376);
or U2815 (N_2815,N_1256,N_1761);
and U2816 (N_2816,N_658,N_2325);
and U2817 (N_2817,N_1971,N_1705);
or U2818 (N_2818,N_1211,N_1823);
and U2819 (N_2819,N_1188,N_1077);
nor U2820 (N_2820,N_1116,N_1289);
and U2821 (N_2821,N_2155,N_1239);
nor U2822 (N_2822,N_591,N_1943);
or U2823 (N_2823,N_1737,N_1813);
or U2824 (N_2824,N_960,N_1268);
or U2825 (N_2825,N_1852,N_92);
or U2826 (N_2826,N_897,N_1146);
nor U2827 (N_2827,N_2459,N_109);
nand U2828 (N_2828,N_820,N_1465);
and U2829 (N_2829,N_2036,N_1417);
or U2830 (N_2830,N_1032,N_869);
and U2831 (N_2831,N_1806,N_601);
and U2832 (N_2832,N_2215,N_1350);
and U2833 (N_2833,N_195,N_501);
nand U2834 (N_2834,N_1452,N_2082);
or U2835 (N_2835,N_2411,N_435);
nor U2836 (N_2836,N_1626,N_975);
nand U2837 (N_2837,N_46,N_419);
and U2838 (N_2838,N_48,N_1664);
and U2839 (N_2839,N_1503,N_1574);
and U2840 (N_2840,N_1693,N_157);
and U2841 (N_2841,N_80,N_2200);
nor U2842 (N_2842,N_2431,N_491);
nor U2843 (N_2843,N_2197,N_153);
nand U2844 (N_2844,N_895,N_36);
nor U2845 (N_2845,N_806,N_2101);
and U2846 (N_2846,N_1969,N_1174);
or U2847 (N_2847,N_2151,N_1329);
nor U2848 (N_2848,N_108,N_1150);
and U2849 (N_2849,N_728,N_2171);
and U2850 (N_2850,N_622,N_1873);
or U2851 (N_2851,N_1906,N_2296);
nand U2852 (N_2852,N_2079,N_1344);
nor U2853 (N_2853,N_450,N_995);
nand U2854 (N_2854,N_1391,N_178);
and U2855 (N_2855,N_1476,N_79);
nand U2856 (N_2856,N_2353,N_585);
and U2857 (N_2857,N_288,N_2408);
or U2858 (N_2858,N_2262,N_1991);
xnor U2859 (N_2859,N_676,N_813);
and U2860 (N_2860,N_1591,N_1511);
nand U2861 (N_2861,N_603,N_546);
or U2862 (N_2862,N_549,N_1125);
or U2863 (N_2863,N_1388,N_492);
nor U2864 (N_2864,N_942,N_2383);
nand U2865 (N_2865,N_377,N_1708);
nand U2866 (N_2866,N_693,N_1458);
nor U2867 (N_2867,N_2201,N_1901);
nand U2868 (N_2868,N_1907,N_1370);
and U2869 (N_2869,N_52,N_221);
nor U2870 (N_2870,N_1069,N_662);
nand U2871 (N_2871,N_505,N_1368);
or U2872 (N_2872,N_1103,N_1520);
or U2873 (N_2873,N_443,N_973);
and U2874 (N_2874,N_977,N_788);
and U2875 (N_2875,N_1933,N_1460);
nor U2876 (N_2876,N_1540,N_749);
nand U2877 (N_2877,N_2253,N_2086);
or U2878 (N_2878,N_154,N_2194);
nand U2879 (N_2879,N_2398,N_1515);
nand U2880 (N_2880,N_1759,N_1012);
nor U2881 (N_2881,N_837,N_2244);
nor U2882 (N_2882,N_926,N_780);
nor U2883 (N_2883,N_1136,N_1921);
or U2884 (N_2884,N_1382,N_2456);
nand U2885 (N_2885,N_1596,N_551);
nor U2886 (N_2886,N_177,N_1054);
nand U2887 (N_2887,N_2016,N_733);
nor U2888 (N_2888,N_2228,N_1844);
nor U2889 (N_2889,N_1927,N_1807);
nand U2890 (N_2890,N_2139,N_740);
nor U2891 (N_2891,N_1251,N_54);
nor U2892 (N_2892,N_208,N_2181);
nor U2893 (N_2893,N_1393,N_584);
or U2894 (N_2894,N_1579,N_858);
and U2895 (N_2895,N_839,N_642);
and U2896 (N_2896,N_1731,N_2188);
nor U2897 (N_2897,N_1006,N_768);
and U2898 (N_2898,N_1249,N_242);
nor U2899 (N_2899,N_882,N_1446);
xnor U2900 (N_2900,N_789,N_1639);
and U2901 (N_2901,N_1760,N_2448);
nor U2902 (N_2902,N_2481,N_955);
or U2903 (N_2903,N_2115,N_1182);
nand U2904 (N_2904,N_1021,N_1041);
nor U2905 (N_2905,N_326,N_925);
nor U2906 (N_2906,N_992,N_781);
and U2907 (N_2907,N_1968,N_1405);
nand U2908 (N_2908,N_1763,N_736);
or U2909 (N_2909,N_917,N_2099);
and U2910 (N_2910,N_2286,N_2141);
and U2911 (N_2911,N_2167,N_1517);
nand U2912 (N_2912,N_504,N_511);
nor U2913 (N_2913,N_1724,N_1419);
or U2914 (N_2914,N_1,N_544);
nand U2915 (N_2915,N_1367,N_1647);
nor U2916 (N_2916,N_1868,N_357);
or U2917 (N_2917,N_1302,N_1837);
or U2918 (N_2918,N_1158,N_1555);
nand U2919 (N_2919,N_1372,N_459);
or U2920 (N_2920,N_533,N_2477);
or U2921 (N_2921,N_2090,N_1483);
nand U2922 (N_2922,N_2142,N_1582);
nor U2923 (N_2923,N_940,N_1865);
and U2924 (N_2924,N_14,N_2392);
and U2925 (N_2925,N_2386,N_2117);
and U2926 (N_2926,N_91,N_2034);
or U2927 (N_2927,N_1757,N_1528);
and U2928 (N_2928,N_1356,N_956);
and U2929 (N_2929,N_286,N_1653);
nor U2930 (N_2930,N_252,N_1038);
and U2931 (N_2931,N_1416,N_2008);
or U2932 (N_2932,N_1109,N_694);
nor U2933 (N_2933,N_2397,N_2463);
nand U2934 (N_2934,N_1217,N_1722);
or U2935 (N_2935,N_844,N_124);
nand U2936 (N_2936,N_396,N_1478);
or U2937 (N_2937,N_690,N_2103);
nand U2938 (N_2938,N_974,N_39);
nand U2939 (N_2939,N_2482,N_814);
nand U2940 (N_2940,N_121,N_1714);
and U2941 (N_2941,N_738,N_1941);
or U2942 (N_2942,N_2031,N_1747);
and U2943 (N_2943,N_508,N_22);
nor U2944 (N_2944,N_119,N_933);
xor U2945 (N_2945,N_888,N_1410);
nand U2946 (N_2946,N_1817,N_42);
and U2947 (N_2947,N_1151,N_1646);
or U2948 (N_2948,N_881,N_1177);
or U2949 (N_2949,N_802,N_991);
nor U2950 (N_2950,N_2451,N_1598);
nor U2951 (N_2951,N_2169,N_132);
nand U2952 (N_2952,N_1554,N_207);
and U2953 (N_2953,N_700,N_1270);
nand U2954 (N_2954,N_2429,N_1565);
nand U2955 (N_2955,N_1732,N_303);
or U2956 (N_2956,N_555,N_854);
and U2957 (N_2957,N_2272,N_903);
or U2958 (N_2958,N_1649,N_31);
nand U2959 (N_2959,N_181,N_1583);
and U2960 (N_2960,N_1950,N_939);
or U2961 (N_2961,N_2288,N_2134);
nand U2962 (N_2962,N_971,N_2308);
nor U2963 (N_2963,N_2252,N_1986);
xor U2964 (N_2964,N_721,N_2317);
xnor U2965 (N_2965,N_2123,N_2363);
and U2966 (N_2966,N_1192,N_1190);
nor U2967 (N_2967,N_1660,N_1385);
and U2968 (N_2968,N_1703,N_2304);
xnor U2969 (N_2969,N_1386,N_1274);
or U2970 (N_2970,N_309,N_417);
and U2971 (N_2971,N_187,N_1669);
nor U2972 (N_2972,N_186,N_1406);
nand U2973 (N_2973,N_2343,N_1683);
and U2974 (N_2974,N_1186,N_1862);
nand U2975 (N_2975,N_1314,N_1278);
nor U2976 (N_2976,N_107,N_1412);
or U2977 (N_2977,N_2093,N_1615);
or U2978 (N_2978,N_117,N_2290);
or U2979 (N_2979,N_1300,N_871);
and U2980 (N_2980,N_1898,N_1529);
nor U2981 (N_2981,N_2106,N_776);
and U2982 (N_2982,N_251,N_845);
nor U2983 (N_2983,N_1129,N_2284);
xnor U2984 (N_2984,N_847,N_1381);
and U2985 (N_2985,N_1387,N_821);
or U2986 (N_2986,N_630,N_1500);
or U2987 (N_2987,N_2145,N_337);
and U2988 (N_2988,N_701,N_677);
or U2989 (N_2989,N_1522,N_543);
nor U2990 (N_2990,N_1518,N_341);
nor U2991 (N_2991,N_1628,N_2113);
and U2992 (N_2992,N_1354,N_1983);
or U2993 (N_2993,N_754,N_1789);
and U2994 (N_2994,N_824,N_1519);
nor U2995 (N_2995,N_445,N_472);
nand U2996 (N_2996,N_2434,N_2050);
nor U2997 (N_2997,N_1307,N_130);
or U2998 (N_2998,N_583,N_37);
nand U2999 (N_2999,N_702,N_1433);
or U3000 (N_3000,N_547,N_1355);
or U3001 (N_3001,N_2158,N_171);
or U3002 (N_3002,N_784,N_2059);
nand U3003 (N_3003,N_717,N_1568);
nor U3004 (N_3004,N_269,N_1715);
or U3005 (N_3005,N_1486,N_1908);
nor U3006 (N_3006,N_4,N_1310);
and U3007 (N_3007,N_638,N_466);
and U3008 (N_3008,N_1401,N_49);
nor U3009 (N_3009,N_953,N_1374);
nand U3010 (N_3010,N_16,N_281);
nand U3011 (N_3011,N_2289,N_2068);
nand U3012 (N_3012,N_617,N_1685);
nor U3013 (N_3013,N_1411,N_112);
nand U3014 (N_3014,N_1919,N_1358);
and U3015 (N_3015,N_349,N_216);
nand U3016 (N_3016,N_1609,N_671);
and U3017 (N_3017,N_2216,N_1748);
nand U3018 (N_3018,N_12,N_1053);
and U3019 (N_3019,N_864,N_870);
or U3020 (N_3020,N_829,N_1184);
nand U3021 (N_3021,N_1414,N_918);
nand U3022 (N_3022,N_963,N_1324);
and U3023 (N_3023,N_2076,N_2052);
or U3024 (N_3024,N_190,N_1979);
nand U3025 (N_3025,N_1874,N_1132);
nand U3026 (N_3026,N_2467,N_1835);
and U3027 (N_3027,N_1612,N_636);
nor U3028 (N_3028,N_1040,N_1764);
and U3029 (N_3029,N_2400,N_2182);
nand U3030 (N_3030,N_774,N_734);
or U3031 (N_3031,N_2421,N_2275);
and U3032 (N_3032,N_1964,N_2410);
or U3033 (N_3033,N_5,N_1524);
nand U3034 (N_3034,N_1283,N_381);
nand U3035 (N_3035,N_1729,N_244);
nand U3036 (N_3036,N_912,N_368);
or U3037 (N_3037,N_202,N_237);
nand U3038 (N_3038,N_1349,N_468);
and U3039 (N_3039,N_1359,N_1730);
nand U3040 (N_3040,N_2381,N_1209);
nand U3041 (N_3041,N_1576,N_1917);
and U3042 (N_3042,N_232,N_579);
nor U3043 (N_3043,N_1996,N_625);
or U3044 (N_3044,N_2022,N_712);
nand U3045 (N_3045,N_1961,N_348);
nand U3046 (N_3046,N_1059,N_397);
nor U3047 (N_3047,N_796,N_1162);
or U3048 (N_3048,N_2470,N_2478);
and U3049 (N_3049,N_947,N_1475);
or U3050 (N_3050,N_2473,N_32);
nand U3051 (N_3051,N_2443,N_1090);
or U3052 (N_3052,N_1456,N_1903);
and U3053 (N_3053,N_2319,N_233);
nand U3054 (N_3054,N_1843,N_664);
and U3055 (N_3055,N_1228,N_1721);
and U3056 (N_3056,N_884,N_423);
or U3057 (N_3057,N_2309,N_168);
nor U3058 (N_3058,N_1851,N_1173);
or U3059 (N_3059,N_2406,N_103);
nand U3060 (N_3060,N_1531,N_612);
nor U3061 (N_3061,N_1810,N_1425);
nor U3062 (N_3062,N_2091,N_351);
nand U3063 (N_3063,N_230,N_1870);
nor U3064 (N_3064,N_1580,N_2204);
nand U3065 (N_3065,N_762,N_2269);
or U3066 (N_3066,N_1273,N_761);
nand U3067 (N_3067,N_1621,N_1504);
and U3068 (N_3068,N_1166,N_1959);
nand U3069 (N_3069,N_1369,N_1342);
nor U3070 (N_3070,N_2497,N_2047);
nor U3071 (N_3071,N_619,N_865);
nand U3072 (N_3072,N_1625,N_1784);
nor U3073 (N_3073,N_680,N_2254);
and U3074 (N_3074,N_586,N_265);
nor U3075 (N_3075,N_811,N_556);
nor U3076 (N_3076,N_493,N_1970);
nor U3077 (N_3077,N_1031,N_1586);
nor U3078 (N_3078,N_2235,N_1665);
and U3079 (N_3079,N_15,N_2312);
nand U3080 (N_3080,N_1326,N_607);
nand U3081 (N_3081,N_518,N_510);
or U3082 (N_3082,N_1644,N_1379);
and U3083 (N_3083,N_29,N_1584);
or U3084 (N_3084,N_1445,N_2154);
and U3085 (N_3085,N_1624,N_1018);
and U3086 (N_3086,N_1882,N_258);
or U3087 (N_3087,N_1076,N_131);
and U3088 (N_3088,N_1765,N_1378);
nor U3089 (N_3089,N_880,N_785);
and U3090 (N_3090,N_1602,N_220);
or U3091 (N_3091,N_747,N_1295);
nand U3092 (N_3092,N_430,N_2023);
nand U3093 (N_3093,N_831,N_1108);
nand U3094 (N_3094,N_559,N_1297);
nor U3095 (N_3095,N_552,N_2046);
and U3096 (N_3096,N_392,N_1952);
nor U3097 (N_3097,N_2057,N_104);
nand U3098 (N_3098,N_590,N_146);
and U3099 (N_3099,N_1214,N_1536);
or U3100 (N_3100,N_247,N_1153);
and U3101 (N_3101,N_1257,N_558);
or U3102 (N_3102,N_1571,N_1506);
and U3103 (N_3103,N_1321,N_1587);
nor U3104 (N_3104,N_134,N_428);
nand U3105 (N_3105,N_1562,N_1233);
nor U3106 (N_3106,N_2382,N_1934);
nand U3107 (N_3107,N_442,N_2116);
or U3108 (N_3108,N_726,N_1622);
nand U3109 (N_3109,N_40,N_2166);
and U3110 (N_3110,N_378,N_1365);
and U3111 (N_3111,N_1595,N_1101);
or U3112 (N_3112,N_347,N_564);
or U3113 (N_3113,N_1306,N_1771);
and U3114 (N_3114,N_2361,N_2330);
or U3115 (N_3115,N_2092,N_1160);
nor U3116 (N_3116,N_691,N_2073);
nor U3117 (N_3117,N_1155,N_203);
nor U3118 (N_3118,N_1316,N_38);
and U3119 (N_3119,N_147,N_930);
or U3120 (N_3120,N_1778,N_452);
nand U3121 (N_3121,N_302,N_1636);
nor U3122 (N_3122,N_1384,N_978);
nor U3123 (N_3123,N_1861,N_2297);
and U3124 (N_3124,N_1453,N_914);
or U3125 (N_3125,N_346,N_2077);
nor U3126 (N_3126,N_105,N_51);
and U3127 (N_3127,N_1913,N_2035);
nor U3128 (N_3128,N_267,N_1046);
nor U3129 (N_3129,N_562,N_1951);
and U3130 (N_3130,N_626,N_569);
nor U3131 (N_3131,N_329,N_1060);
nand U3132 (N_3132,N_1219,N_462);
nor U3133 (N_3133,N_2480,N_469);
nor U3134 (N_3134,N_1766,N_684);
nor U3135 (N_3135,N_167,N_2393);
nor U3136 (N_3136,N_90,N_2230);
or U3137 (N_3137,N_436,N_758);
nor U3138 (N_3138,N_2298,N_2307);
or U3139 (N_3139,N_1717,N_21);
or U3140 (N_3140,N_922,N_928);
nand U3141 (N_3141,N_2164,N_2131);
and U3142 (N_3142,N_2367,N_1699);
and U3143 (N_3143,N_176,N_2198);
nor U3144 (N_3144,N_861,N_656);
nand U3145 (N_3145,N_1548,N_1208);
and U3146 (N_3146,N_2415,N_2163);
nor U3147 (N_3147,N_156,N_2160);
and U3148 (N_3148,N_1547,N_1911);
or U3149 (N_3149,N_17,N_1716);
or U3150 (N_3150,N_1527,N_757);
or U3151 (N_3151,N_1638,N_249);
and U3152 (N_3152,N_2006,N_716);
and U3153 (N_3153,N_1820,N_990);
nor U3154 (N_3154,N_375,N_1993);
nor U3155 (N_3155,N_1945,N_663);
or U3156 (N_3156,N_786,N_266);
and U3157 (N_3157,N_2104,N_2179);
or U3158 (N_3158,N_1203,N_1123);
nor U3159 (N_3159,N_598,N_1947);
and U3160 (N_3160,N_1066,N_705);
and U3161 (N_3161,N_78,N_1836);
nand U3162 (N_3162,N_1659,N_605);
xor U3163 (N_3163,N_1803,N_1942);
and U3164 (N_3164,N_877,N_708);
or U3165 (N_3165,N_592,N_1328);
nand U3166 (N_3166,N_760,N_1311);
and U3167 (N_3167,N_2085,N_1334);
or U3168 (N_3168,N_2030,N_818);
or U3169 (N_3169,N_481,N_403);
nor U3170 (N_3170,N_1977,N_94);
or U3171 (N_3171,N_2355,N_2185);
and U3172 (N_3172,N_2402,N_1756);
or U3173 (N_3173,N_407,N_301);
nand U3174 (N_3174,N_661,N_138);
and U3175 (N_3175,N_2425,N_945);
nor U3176 (N_3176,N_447,N_2058);
nor U3177 (N_3177,N_2472,N_234);
and U3178 (N_3178,N_334,N_1981);
or U3179 (N_3179,N_429,N_2246);
or U3180 (N_3180,N_214,N_2377);
nand U3181 (N_3181,N_367,N_1137);
or U3182 (N_3182,N_70,N_1702);
nor U3183 (N_3183,N_317,N_172);
or U3184 (N_3184,N_285,N_931);
nor U3185 (N_3185,N_2029,N_682);
or U3186 (N_3186,N_2264,N_2424);
nand U3187 (N_3187,N_152,N_25);
nand U3188 (N_3188,N_859,N_1258);
or U3189 (N_3189,N_1016,N_1193);
or U3190 (N_3190,N_2476,N_2191);
nand U3191 (N_3191,N_353,N_910);
and U3192 (N_3192,N_1126,N_1327);
nor U3193 (N_3193,N_1082,N_1516);
nand U3194 (N_3194,N_841,N_2143);
or U3195 (N_3195,N_1271,N_1436);
or U3196 (N_3196,N_1614,N_2422);
and U3197 (N_3197,N_11,N_393);
nor U3198 (N_3198,N_689,N_1978);
and U3199 (N_3199,N_860,N_529);
or U3200 (N_3200,N_1751,N_434);
nand U3201 (N_3201,N_615,N_695);
and U3202 (N_3202,N_927,N_1532);
and U3203 (N_3203,N_653,N_1044);
and U3204 (N_3204,N_1575,N_61);
or U3205 (N_3205,N_2432,N_999);
nand U3206 (N_3206,N_2493,N_513);
nor U3207 (N_3207,N_902,N_1984);
or U3208 (N_3208,N_1753,N_1345);
nor U3209 (N_3209,N_2071,N_1484);
nor U3210 (N_3210,N_1866,N_2435);
and U3211 (N_3211,N_188,N_589);
nor U3212 (N_3212,N_1468,N_2129);
nand U3213 (N_3213,N_1247,N_1438);
nor U3214 (N_3214,N_2486,N_1161);
nor U3215 (N_3215,N_325,N_2240);
and U3216 (N_3216,N_1994,N_1435);
nand U3217 (N_3217,N_1490,N_1055);
or U3218 (N_3218,N_283,N_282);
nand U3219 (N_3219,N_809,N_1092);
nor U3220 (N_3220,N_2315,N_1838);
nor U3221 (N_3221,N_1312,N_1505);
nor U3222 (N_3222,N_2187,N_333);
nand U3223 (N_3223,N_666,N_582);
or U3224 (N_3224,N_1212,N_2135);
and U3225 (N_3225,N_1740,N_2372);
and U3226 (N_3226,N_1364,N_965);
or U3227 (N_3227,N_1938,N_1916);
or U3228 (N_3228,N_1253,N_643);
nor U3229 (N_3229,N_874,N_2460);
and U3230 (N_3230,N_1796,N_1131);
nor U3231 (N_3231,N_1361,N_201);
and U3232 (N_3232,N_1551,N_45);
and U3233 (N_3233,N_1973,N_1613);
and U3234 (N_3234,N_1172,N_548);
and U3235 (N_3235,N_129,N_2041);
and U3236 (N_3236,N_2371,N_1340);
and U3237 (N_3237,N_1169,N_227);
and U3238 (N_3238,N_1130,N_2331);
xor U3239 (N_3239,N_1254,N_1680);
and U3240 (N_3240,N_2100,N_135);
nor U3241 (N_3241,N_1805,N_150);
and U3242 (N_3242,N_1403,N_453);
or U3243 (N_3243,N_2390,N_1244);
nand U3244 (N_3244,N_1900,N_1695);
nor U3245 (N_3245,N_1205,N_1432);
nand U3246 (N_3246,N_2000,N_2471);
nand U3247 (N_3247,N_205,N_2152);
nor U3248 (N_3248,N_1111,N_55);
and U3249 (N_3249,N_360,N_2466);
or U3250 (N_3250,N_44,N_697);
nor U3251 (N_3251,N_1206,N_997);
and U3252 (N_3252,N_2225,N_862);
nand U3253 (N_3253,N_1423,N_1822);
and U3254 (N_3254,N_1133,N_1081);
or U3255 (N_3255,N_2295,N_1201);
nor U3256 (N_3256,N_1422,N_1078);
or U3257 (N_3257,N_1681,N_1932);
or U3258 (N_3258,N_354,N_1003);
nand U3259 (N_3259,N_983,N_2251);
or U3260 (N_3260,N_834,N_1946);
and U3261 (N_3261,N_1317,N_433);
nand U3262 (N_3262,N_1087,N_1573);
nor U3263 (N_3263,N_2212,N_246);
and U3264 (N_3264,N_1544,N_1767);
nand U3265 (N_3265,N_1619,N_867);
or U3266 (N_3266,N_1672,N_1989);
and U3267 (N_3267,N_1280,N_2445);
and U3268 (N_3268,N_1426,N_259);
xor U3269 (N_3269,N_935,N_1091);
or U3270 (N_3270,N_1677,N_1255);
or U3271 (N_3271,N_413,N_566);
nor U3272 (N_3272,N_567,N_2021);
or U3273 (N_3273,N_165,N_2344);
nand U3274 (N_3274,N_537,N_2368);
and U3275 (N_3275,N_2278,N_166);
nand U3276 (N_3276,N_2001,N_623);
nand U3277 (N_3277,N_1877,N_2498);
and U3278 (N_3278,N_1057,N_1962);
nor U3279 (N_3279,N_2321,N_2060);
nor U3280 (N_3280,N_1114,N_742);
xor U3281 (N_3281,N_1674,N_640);
and U3282 (N_3282,N_312,N_628);
and U3283 (N_3283,N_1226,N_570);
nand U3284 (N_3284,N_2172,N_1341);
and U3285 (N_3285,N_565,N_148);
or U3286 (N_3286,N_2441,N_2348);
nor U3287 (N_3287,N_1462,N_1645);
or U3288 (N_3288,N_1034,N_422);
and U3289 (N_3289,N_832,N_1434);
nand U3290 (N_3290,N_920,N_1590);
and U3291 (N_3291,N_284,N_87);
and U3292 (N_3292,N_1265,N_425);
and U3293 (N_3293,N_2233,N_406);
and U3294 (N_3294,N_28,N_1671);
or U3295 (N_3295,N_849,N_225);
or U3296 (N_3296,N_2474,N_2327);
or U3297 (N_3297,N_66,N_398);
or U3298 (N_3298,N_2404,N_1145);
nor U3299 (N_3299,N_1601,N_140);
and U3300 (N_3300,N_356,N_243);
and U3301 (N_3301,N_1834,N_2222);
xnor U3302 (N_3302,N_1142,N_1935);
or U3303 (N_3303,N_798,N_2396);
or U3304 (N_3304,N_2045,N_1704);
xor U3305 (N_3305,N_710,N_1100);
nand U3306 (N_3306,N_2301,N_1871);
or U3307 (N_3307,N_1448,N_24);
or U3308 (N_3308,N_1279,N_2267);
and U3309 (N_3309,N_1526,N_1180);
or U3310 (N_3310,N_2258,N_1036);
nor U3311 (N_3311,N_290,N_1120);
nand U3312 (N_3312,N_2364,N_1080);
or U3313 (N_3313,N_58,N_274);
or U3314 (N_3314,N_1910,N_713);
nor U3315 (N_3315,N_2054,N_1779);
nor U3316 (N_3316,N_489,N_618);
and U3317 (N_3317,N_2273,N_1402);
nand U3318 (N_3318,N_2311,N_2350);
and U3319 (N_3319,N_840,N_2436);
or U3320 (N_3320,N_2128,N_1744);
and U3321 (N_3321,N_2097,N_1396);
and U3322 (N_3322,N_573,N_141);
or U3323 (N_3323,N_2125,N_516);
and U3324 (N_3324,N_1139,N_587);
nand U3325 (N_3325,N_1980,N_779);
nor U3326 (N_3326,N_517,N_1643);
nand U3327 (N_3327,N_1824,N_386);
nand U3328 (N_3328,N_1325,N_1276);
or U3329 (N_3329,N_1439,N_263);
and U3330 (N_3330,N_1319,N_306);
nand U3331 (N_3331,N_852,N_1320);
or U3332 (N_3332,N_81,N_2366);
and U3333 (N_3333,N_651,N_2320);
nor U3334 (N_3334,N_668,N_1728);
and U3335 (N_3335,N_1148,N_1346);
or U3336 (N_3336,N_1230,N_2002);
nor U3337 (N_3337,N_1958,N_1648);
or U3338 (N_3338,N_2263,N_1794);
and U3339 (N_3339,N_2499,N_1787);
nand U3340 (N_3340,N_2239,N_460);
nand U3341 (N_3341,N_2437,N_833);
nor U3342 (N_3342,N_1893,N_904);
and U3343 (N_3343,N_1404,N_1521);
nor U3344 (N_3344,N_981,N_907);
or U3345 (N_3345,N_1750,N_756);
and U3346 (N_3346,N_924,N_1339);
nand U3347 (N_3347,N_1159,N_1428);
or U3348 (N_3348,N_293,N_1696);
or U3349 (N_3349,N_359,N_635);
nor U3350 (N_3350,N_1797,N_198);
nor U3351 (N_3351,N_1666,N_685);
or U3352 (N_3352,N_2300,N_2446);
nand U3353 (N_3353,N_330,N_41);
nor U3354 (N_3354,N_898,N_2220);
and U3355 (N_3355,N_2193,N_1775);
nand U3356 (N_3356,N_245,N_262);
or U3357 (N_3357,N_709,N_1512);
nor U3358 (N_3358,N_2418,N_440);
and U3359 (N_3359,N_1110,N_1655);
nor U3360 (N_3360,N_451,N_65);
nand U3361 (N_3361,N_1000,N_1262);
nor U3362 (N_3362,N_993,N_890);
nand U3363 (N_3363,N_1990,N_1363);
and U3364 (N_3364,N_299,N_1603);
nand U3365 (N_3365,N_362,N_792);
or U3366 (N_3366,N_2063,N_1700);
and U3367 (N_3367,N_1608,N_637);
or U3368 (N_3368,N_674,N_621);
or U3369 (N_3369,N_538,N_272);
nand U3370 (N_3370,N_2256,N_1096);
and U3371 (N_3371,N_988,N_892);
nor U3372 (N_3372,N_473,N_1872);
nor U3373 (N_3373,N_827,N_969);
or U3374 (N_3374,N_686,N_2084);
nand U3375 (N_3375,N_412,N_364);
nor U3376 (N_3376,N_344,N_982);
nand U3377 (N_3377,N_410,N_1712);
nand U3378 (N_3378,N_1313,N_1075);
nand U3379 (N_3379,N_212,N_2207);
and U3380 (N_3380,N_575,N_223);
nor U3381 (N_3381,N_571,N_909);
or U3382 (N_3382,N_98,N_2102);
nand U3383 (N_3383,N_482,N_714);
nand U3384 (N_3384,N_1808,N_0);
and U3385 (N_3385,N_1985,N_2403);
and U3386 (N_3386,N_345,N_2494);
or U3387 (N_3387,N_2428,N_2352);
or U3388 (N_3388,N_596,N_1651);
nand U3389 (N_3389,N_1944,N_1074);
nor U3390 (N_3390,N_1848,N_1007);
and U3391 (N_3391,N_886,N_2096);
or U3392 (N_3392,N_795,N_1707);
nand U3393 (N_3393,N_1833,N_96);
and U3394 (N_3394,N_539,N_1741);
or U3395 (N_3395,N_2495,N_1599);
nor U3396 (N_3396,N_151,N_2292);
nand U3397 (N_3397,N_231,N_1437);
or U3398 (N_3398,N_2414,N_1963);
nand U3399 (N_3399,N_1738,N_692);
or U3400 (N_3400,N_1581,N_1019);
or U3401 (N_3401,N_577,N_1014);
and U3402 (N_3402,N_1501,N_1236);
or U3403 (N_3403,N_759,N_2192);
nand U3404 (N_3404,N_1135,N_226);
nor U3405 (N_3405,N_2025,N_1430);
and U3406 (N_3406,N_2492,N_476);
or U3407 (N_3407,N_278,N_1541);
and U3408 (N_3408,N_1459,N_657);
or U3409 (N_3409,N_2338,N_1918);
and U3410 (N_3410,N_2037,N_727);
or U3411 (N_3411,N_1207,N_77);
nand U3412 (N_3412,N_1143,N_2119);
nand U3413 (N_3413,N_777,N_2157);
or U3414 (N_3414,N_1839,N_2159);
or U3415 (N_3415,N_1250,N_1881);
nor U3416 (N_3416,N_2439,N_2221);
nor U3417 (N_3417,N_1926,N_310);
nor U3418 (N_3418,N_1617,N_175);
and U3419 (N_3419,N_1826,N_1758);
nor U3420 (N_3420,N_2455,N_1252);
nand U3421 (N_3421,N_669,N_812);
nor U3422 (N_3422,N_1925,N_2374);
and U3423 (N_3423,N_1304,N_2161);
and U3424 (N_3424,N_485,N_2042);
xnor U3425 (N_3425,N_530,N_593);
nor U3426 (N_3426,N_143,N_1954);
nand U3427 (N_3427,N_1995,N_155);
or U3428 (N_3428,N_2464,N_1204);
nand U3429 (N_3429,N_2282,N_363);
nand U3430 (N_3430,N_574,N_289);
nand U3431 (N_3431,N_1157,N_711);
and U3432 (N_3432,N_2137,N_62);
and U3433 (N_3433,N_1183,N_1115);
and U3434 (N_3434,N_120,N_264);
and U3435 (N_3435,N_836,N_962);
and U3436 (N_3436,N_830,N_2335);
and U3437 (N_3437,N_2126,N_487);
and U3438 (N_3438,N_495,N_578);
and U3439 (N_3439,N_1407,N_261);
or U3440 (N_3440,N_944,N_887);
and U3441 (N_3441,N_748,N_2196);
nor U3442 (N_3442,N_8,N_2053);
and U3443 (N_3443,N_1641,N_1675);
nand U3444 (N_3444,N_1373,N_1421);
nand U3445 (N_3445,N_1360,N_174);
nand U3446 (N_3446,N_350,N_985);
and U3447 (N_3447,N_866,N_1191);
nand U3448 (N_3448,N_1819,N_704);
nand U3449 (N_3449,N_217,N_1909);
nand U3450 (N_3450,N_604,N_938);
nand U3451 (N_3451,N_2427,N_1291);
nand U3452 (N_3452,N_629,N_1175);
nor U3453 (N_3453,N_467,N_206);
nor U3454 (N_3454,N_1348,N_1967);
or U3455 (N_3455,N_1029,N_1928);
nand U3456 (N_3456,N_679,N_2210);
xnor U3457 (N_3457,N_1024,N_659);
nor U3458 (N_3458,N_1408,N_1285);
and U3459 (N_3459,N_1303,N_519);
or U3460 (N_3460,N_2457,N_1238);
or U3461 (N_3461,N_210,N_1001);
and U3462 (N_3462,N_783,N_1930);
nand U3463 (N_3463,N_1380,N_1923);
nor U3464 (N_3464,N_2345,N_797);
nand U3465 (N_3465,N_1697,N_1400);
or U3466 (N_3466,N_2007,N_1431);
or U3467 (N_3467,N_2114,N_817);
nor U3468 (N_3468,N_509,N_1427);
and U3469 (N_3469,N_370,N_1022);
nand U3470 (N_3470,N_255,N_1144);
and U3471 (N_3471,N_56,N_2095);
and U3472 (N_3472,N_401,N_1698);
or U3473 (N_3473,N_355,N_793);
or U3474 (N_3474,N_1620,N_1880);
nand U3475 (N_3475,N_1627,N_2);
nor U3476 (N_3476,N_2107,N_934);
and U3477 (N_3477,N_1564,N_2303);
or U3478 (N_3478,N_399,N_816);
nor U3479 (N_3479,N_1333,N_660);
and U3480 (N_3480,N_1070,N_1832);
and U3481 (N_3481,N_160,N_477);
nor U3482 (N_3482,N_228,N_1710);
and U3483 (N_3483,N_2485,N_750);
nand U3484 (N_3484,N_67,N_532);
nand U3485 (N_3485,N_1800,N_2011);
and U3486 (N_3486,N_1113,N_647);
and U3487 (N_3487,N_457,N_1542);
or U3488 (N_3488,N_2268,N_1105);
nand U3489 (N_3489,N_128,N_1472);
and U3490 (N_3490,N_1088,N_803);
and U3491 (N_3491,N_72,N_2433);
or U3492 (N_3492,N_1642,N_1048);
and U3493 (N_3493,N_1245,N_182);
nand U3494 (N_3494,N_179,N_1798);
or U3495 (N_3495,N_1742,N_1487);
nand U3496 (N_3496,N_534,N_2219);
nor U3497 (N_3497,N_1999,N_1196);
nand U3498 (N_3498,N_1030,N_1965);
and U3499 (N_3499,N_1924,N_1746);
and U3500 (N_3500,N_2224,N_2358);
and U3501 (N_3501,N_634,N_170);
nand U3502 (N_3502,N_594,N_2072);
nand U3503 (N_3503,N_2203,N_324);
nor U3504 (N_3504,N_2328,N_1409);
nand U3505 (N_3505,N_957,N_949);
nand U3506 (N_3506,N_1002,N_204);
and U3507 (N_3507,N_439,N_1037);
or U3508 (N_3508,N_2049,N_1085);
or U3509 (N_3509,N_1194,N_1523);
and U3510 (N_3510,N_268,N_1332);
and U3511 (N_3511,N_2094,N_1569);
nor U3512 (N_3512,N_296,N_1514);
nand U3513 (N_3513,N_389,N_1799);
nand U3514 (N_3514,N_390,N_1390);
or U3515 (N_3515,N_2180,N_2040);
and U3516 (N_3516,N_1706,N_1353);
and U3517 (N_3517,N_1860,N_1454);
nor U3518 (N_3518,N_2136,N_639);
nand U3519 (N_3519,N_1117,N_1572);
nand U3520 (N_3520,N_332,N_876);
and U3521 (N_3521,N_958,N_2270);
and U3522 (N_3522,N_2462,N_1292);
and U3523 (N_3523,N_1630,N_1397);
or U3524 (N_3524,N_1790,N_2313);
nor U3525 (N_3525,N_164,N_751);
and U3526 (N_3526,N_857,N_1635);
or U3527 (N_3527,N_13,N_521);
xnor U3528 (N_3528,N_2465,N_2017);
and U3529 (N_3529,N_1269,N_1629);
nor U3530 (N_3530,N_1272,N_270);
nor U3531 (N_3531,N_2420,N_1473);
nand U3532 (N_3532,N_6,N_1684);
nor U3533 (N_3533,N_514,N_1895);
nand U3534 (N_3534,N_863,N_1546);
nand U3535 (N_3535,N_1899,N_722);
nand U3536 (N_3536,N_97,N_1127);
and U3537 (N_3537,N_2291,N_739);
and U3538 (N_3538,N_2081,N_568);
nor U3539 (N_3539,N_311,N_771);
or U3540 (N_3540,N_1389,N_319);
nor U3541 (N_3541,N_1413,N_899);
nor U3542 (N_3542,N_1745,N_446);
and U3543 (N_3543,N_7,N_2055);
nand U3544 (N_3544,N_846,N_1171);
and U3545 (N_3545,N_1508,N_1735);
and U3546 (N_3546,N_1231,N_1084);
nand U3547 (N_3547,N_316,N_2205);
nand U3548 (N_3548,N_948,N_905);
nor U3549 (N_3549,N_2334,N_650);
and U3550 (N_3550,N_633,N_1284);
nand U3551 (N_3551,N_2232,N_1736);
or U3552 (N_3552,N_1713,N_875);
and U3553 (N_3553,N_807,N_1027);
and U3554 (N_3554,N_2098,N_1897);
or U3555 (N_3555,N_2365,N_563);
nand U3556 (N_3556,N_1661,N_672);
and U3557 (N_3557,N_1094,N_1890);
or U3558 (N_3558,N_2259,N_1176);
nand U3559 (N_3559,N_2010,N_2237);
nor U3560 (N_3560,N_576,N_95);
nor U3561 (N_3561,N_1118,N_2118);
nand U3562 (N_3562,N_1067,N_2281);
and U3563 (N_3563,N_409,N_145);
and U3564 (N_3564,N_872,N_1863);
and U3565 (N_3565,N_526,N_1227);
and U3566 (N_3566,N_2004,N_1073);
or U3567 (N_3567,N_2490,N_27);
nand U3568 (N_3568,N_2150,N_2110);
or U3569 (N_3569,N_665,N_1068);
nor U3570 (N_3570,N_1815,N_654);
nor U3571 (N_3571,N_101,N_1654);
and U3572 (N_3572,N_209,N_1892);
nor U3573 (N_3573,N_2416,N_787);
and U3574 (N_3574,N_2226,N_2173);
or U3575 (N_3575,N_994,N_1553);
or U3576 (N_3576,N_395,N_1694);
nor U3577 (N_3577,N_1762,N_1287);
or U3578 (N_3578,N_1768,N_2356);
and U3579 (N_3579,N_361,N_384);
nand U3580 (N_3580,N_2310,N_1948);
or U3581 (N_3581,N_1853,N_652);
or U3582 (N_3582,N_536,N_1864);
and U3583 (N_3583,N_1795,N_292);
and U3584 (N_3584,N_1850,N_557);
nand U3585 (N_3585,N_2294,N_1352);
xor U3586 (N_3586,N_1752,N_1450);
nor U3587 (N_3587,N_646,N_2168);
or U3588 (N_3588,N_1633,N_916);
and U3589 (N_3589,N_1449,N_184);
or U3590 (N_3590,N_1772,N_1288);
and U3591 (N_3591,N_222,N_1197);
and U3592 (N_3592,N_737,N_2067);
nor U3593 (N_3593,N_372,N_241);
or U3594 (N_3594,N_431,N_1780);
nand U3595 (N_3595,N_1266,N_2468);
or U3596 (N_3596,N_416,N_542);
nand U3597 (N_3597,N_2149,N_1585);
nor U3598 (N_3598,N_1261,N_1525);
nor U3599 (N_3599,N_614,N_1709);
or U3600 (N_3600,N_1246,N_366);
or U3601 (N_3601,N_580,N_2380);
and U3602 (N_3602,N_1063,N_1241);
nor U3603 (N_3603,N_2388,N_753);
or U3604 (N_3604,N_315,N_2423);
or U3605 (N_3605,N_1065,N_219);
nor U3606 (N_3606,N_1179,N_506);
and U3607 (N_3607,N_1679,N_1043);
xnor U3608 (N_3608,N_461,N_1152);
and U3609 (N_3609,N_828,N_1957);
nor U3610 (N_3610,N_815,N_613);
or U3611 (N_3611,N_946,N_215);
nor U3612 (N_3612,N_553,N_755);
and U3613 (N_3613,N_196,N_900);
nand U3614 (N_3614,N_1733,N_2375);
or U3615 (N_3615,N_1140,N_1904);
or U3616 (N_3616,N_1727,N_893);
nand U3617 (N_3617,N_1818,N_1371);
nand U3618 (N_3618,N_1045,N_169);
or U3619 (N_3619,N_687,N_908);
and U3620 (N_3620,N_1912,N_426);
and U3621 (N_3621,N_1017,N_1441);
or U3622 (N_3622,N_535,N_2105);
nor U3623 (N_3623,N_248,N_1187);
or U3624 (N_3624,N_444,N_1689);
or U3625 (N_3625,N_1533,N_2111);
nand U3626 (N_3626,N_2357,N_1351);
nand U3627 (N_3627,N_525,N_1859);
or U3628 (N_3628,N_2132,N_33);
nand U3629 (N_3629,N_2354,N_572);
nand U3630 (N_3630,N_1607,N_1711);
nand U3631 (N_3631,N_2384,N_2144);
or U3632 (N_3632,N_380,N_352);
and U3633 (N_3633,N_683,N_404);
and U3634 (N_3634,N_2089,N_2285);
or U3635 (N_3635,N_588,N_2341);
and U3636 (N_3636,N_2454,N_498);
nor U3637 (N_3637,N_2199,N_923);
and U3638 (N_3638,N_320,N_2214);
nor U3639 (N_3639,N_2444,N_2206);
and U3640 (N_3640,N_1167,N_2027);
nor U3641 (N_3641,N_1690,N_1987);
and U3642 (N_3642,N_471,N_715);
and U3643 (N_3643,N_611,N_1605);
nor U3644 (N_3644,N_1953,N_85);
or U3645 (N_3645,N_1556,N_93);
xor U3646 (N_3646,N_1539,N_2005);
nand U3647 (N_3647,N_1788,N_964);
or U3648 (N_3648,N_2162,N_2491);
or U3649 (N_3649,N_767,N_1769);
nand U3650 (N_3650,N_1894,N_2033);
nand U3651 (N_3651,N_2340,N_382);
nand U3652 (N_3652,N_2013,N_71);
or U3653 (N_3653,N_723,N_1592);
or U3654 (N_3654,N_2183,N_1976);
nand U3655 (N_3655,N_2109,N_2342);
and U3656 (N_3656,N_1330,N_1010);
or U3657 (N_3657,N_719,N_996);
nand U3658 (N_3658,N_2195,N_2019);
nor U3659 (N_3659,N_475,N_2430);
and U3660 (N_3660,N_1260,N_1039);
or U3661 (N_3661,N_1557,N_1847);
and U3662 (N_3662,N_1394,N_115);
nor U3663 (N_3663,N_699,N_515);
or U3664 (N_3664,N_189,N_707);
nor U3665 (N_3665,N_192,N_1558);
nor U3666 (N_3666,N_1232,N_1218);
or U3667 (N_3667,N_741,N_1337);
and U3668 (N_3668,N_2249,N_1418);
or U3669 (N_3669,N_2324,N_540);
and U3670 (N_3670,N_951,N_2003);
and U3671 (N_3671,N_1290,N_998);
xnor U3672 (N_3672,N_1223,N_10);
nor U3673 (N_3673,N_1589,N_1497);
nand U3674 (N_3674,N_1199,N_1466);
and U3675 (N_3675,N_496,N_921);
nor U3676 (N_3676,N_1884,N_76);
or U3677 (N_3677,N_1992,N_937);
or U3678 (N_3678,N_1725,N_610);
nor U3679 (N_3679,N_163,N_1955);
and U3680 (N_3680,N_280,N_1902);
nand U3681 (N_3681,N_2039,N_322);
nor U3682 (N_3682,N_229,N_89);
nand U3683 (N_3683,N_1507,N_463);
nand U3684 (N_3684,N_763,N_1004);
nor U3685 (N_3685,N_1056,N_123);
and U3686 (N_3686,N_2175,N_1701);
or U3687 (N_3687,N_1200,N_1816);
and U3688 (N_3688,N_703,N_1652);
nor U3689 (N_3689,N_2302,N_464);
or U3690 (N_3690,N_950,N_116);
nand U3691 (N_3691,N_1804,N_773);
nand U3692 (N_3692,N_1299,N_342);
nor U3693 (N_3693,N_1005,N_550);
nand U3694 (N_3694,N_1104,N_488);
or U3695 (N_3695,N_1282,N_2026);
nand U3696 (N_3696,N_602,N_191);
or U3697 (N_3697,N_1301,N_2229);
and U3698 (N_3698,N_1876,N_1998);
or U3699 (N_3699,N_287,N_541);
nor U3700 (N_3700,N_2231,N_185);
nand U3701 (N_3701,N_1550,N_2218);
nand U3702 (N_3702,N_688,N_520);
or U3703 (N_3703,N_856,N_2070);
nor U3704 (N_3704,N_250,N_448);
nor U3705 (N_3705,N_2440,N_437);
or U3706 (N_3706,N_1335,N_1089);
or U3707 (N_3707,N_2048,N_458);
nor U3708 (N_3708,N_1195,N_2362);
nand U3709 (N_3709,N_69,N_752);
and U3710 (N_3710,N_2261,N_2332);
nand U3711 (N_3711,N_879,N_648);
nor U3712 (N_3712,N_1221,N_1485);
and U3713 (N_3713,N_599,N_1791);
nand U3714 (N_3714,N_2018,N_358);
and U3715 (N_3715,N_1229,N_932);
and U3716 (N_3716,N_670,N_878);
nor U3717 (N_3717,N_331,N_1477);
or U3718 (N_3718,N_1563,N_1392);
or U3719 (N_3719,N_1025,N_474);
or U3720 (N_3720,N_2339,N_1509);
nand U3721 (N_3721,N_2369,N_2032);
or U3722 (N_3722,N_2387,N_1858);
nor U3723 (N_3723,N_1841,N_1447);
and U3724 (N_3724,N_1479,N_2121);
or U3725 (N_3725,N_110,N_1107);
and U3726 (N_3726,N_2190,N_984);
nor U3727 (N_3727,N_1997,N_2489);
or U3728 (N_3728,N_411,N_499);
nor U3729 (N_3729,N_1216,N_746);
or U3730 (N_3730,N_2379,N_1042);
xor U3731 (N_3731,N_327,N_1494);
and U3732 (N_3732,N_2174,N_1469);
and U3733 (N_3733,N_1537,N_1124);
nor U3734 (N_3734,N_976,N_2412);
and U3735 (N_3735,N_1050,N_321);
nand U3736 (N_3736,N_770,N_2148);
or U3737 (N_3737,N_1593,N_2051);
and U3738 (N_3738,N_1686,N_620);
or U3739 (N_3739,N_1489,N_1770);
or U3740 (N_3740,N_696,N_804);
nor U3741 (N_3741,N_1879,N_26);
or U3742 (N_3742,N_1670,N_868);
nand U3743 (N_3743,N_86,N_2360);
nand U3744 (N_3744,N_454,N_1338);
nor U3745 (N_3745,N_73,N_2496);
or U3746 (N_3746,N_1597,N_323);
or U3747 (N_3747,N_2283,N_2409);
nor U3748 (N_3748,N_277,N_1315);
or U3749 (N_3749,N_2487,N_896);
and U3750 (N_3750,N_297,N_1342);
or U3751 (N_3751,N_803,N_681);
nor U3752 (N_3752,N_1459,N_1183);
and U3753 (N_3753,N_2205,N_1196);
and U3754 (N_3754,N_905,N_1516);
or U3755 (N_3755,N_1634,N_756);
and U3756 (N_3756,N_1625,N_1133);
nor U3757 (N_3757,N_1800,N_1798);
or U3758 (N_3758,N_2409,N_1904);
nand U3759 (N_3759,N_860,N_1607);
and U3760 (N_3760,N_1432,N_1237);
and U3761 (N_3761,N_111,N_343);
nand U3762 (N_3762,N_1423,N_927);
xnor U3763 (N_3763,N_1380,N_2448);
xnor U3764 (N_3764,N_1843,N_1897);
nor U3765 (N_3765,N_1983,N_1049);
or U3766 (N_3766,N_52,N_361);
nor U3767 (N_3767,N_1170,N_624);
nand U3768 (N_3768,N_58,N_1434);
and U3769 (N_3769,N_2226,N_2252);
and U3770 (N_3770,N_353,N_711);
nor U3771 (N_3771,N_213,N_167);
nand U3772 (N_3772,N_802,N_1009);
nor U3773 (N_3773,N_1022,N_475);
or U3774 (N_3774,N_2280,N_1533);
or U3775 (N_3775,N_1376,N_1225);
nor U3776 (N_3776,N_902,N_2006);
and U3777 (N_3777,N_1832,N_1778);
and U3778 (N_3778,N_1476,N_2345);
and U3779 (N_3779,N_402,N_410);
nor U3780 (N_3780,N_250,N_2033);
nor U3781 (N_3781,N_973,N_967);
and U3782 (N_3782,N_1423,N_2051);
nand U3783 (N_3783,N_302,N_132);
and U3784 (N_3784,N_2179,N_1581);
and U3785 (N_3785,N_1169,N_1271);
nor U3786 (N_3786,N_297,N_245);
or U3787 (N_3787,N_2041,N_938);
and U3788 (N_3788,N_2276,N_1580);
nor U3789 (N_3789,N_1200,N_1647);
nand U3790 (N_3790,N_1999,N_284);
nand U3791 (N_3791,N_115,N_1639);
and U3792 (N_3792,N_637,N_755);
and U3793 (N_3793,N_1467,N_707);
and U3794 (N_3794,N_653,N_2190);
or U3795 (N_3795,N_51,N_1175);
nand U3796 (N_3796,N_945,N_1430);
or U3797 (N_3797,N_2135,N_1419);
nor U3798 (N_3798,N_1036,N_1814);
nand U3799 (N_3799,N_426,N_1580);
nor U3800 (N_3800,N_1956,N_1662);
nand U3801 (N_3801,N_1282,N_1227);
nor U3802 (N_3802,N_1051,N_1932);
or U3803 (N_3803,N_606,N_1331);
or U3804 (N_3804,N_387,N_1643);
or U3805 (N_3805,N_2386,N_301);
nand U3806 (N_3806,N_147,N_665);
or U3807 (N_3807,N_1411,N_1059);
nor U3808 (N_3808,N_1292,N_1148);
or U3809 (N_3809,N_1349,N_153);
or U3810 (N_3810,N_2431,N_698);
nor U3811 (N_3811,N_1397,N_844);
and U3812 (N_3812,N_1910,N_1475);
nor U3813 (N_3813,N_2307,N_1309);
nand U3814 (N_3814,N_1033,N_1677);
nand U3815 (N_3815,N_357,N_1901);
or U3816 (N_3816,N_751,N_2384);
or U3817 (N_3817,N_2323,N_1484);
and U3818 (N_3818,N_271,N_1302);
nand U3819 (N_3819,N_64,N_1146);
and U3820 (N_3820,N_714,N_1171);
nand U3821 (N_3821,N_2370,N_1670);
or U3822 (N_3822,N_1337,N_877);
or U3823 (N_3823,N_281,N_631);
nor U3824 (N_3824,N_1969,N_1344);
nand U3825 (N_3825,N_1938,N_1357);
and U3826 (N_3826,N_2205,N_1412);
xnor U3827 (N_3827,N_1110,N_1439);
and U3828 (N_3828,N_208,N_1639);
or U3829 (N_3829,N_1777,N_1285);
or U3830 (N_3830,N_2037,N_2395);
and U3831 (N_3831,N_982,N_168);
or U3832 (N_3832,N_2421,N_2054);
and U3833 (N_3833,N_2065,N_2171);
nor U3834 (N_3834,N_539,N_1948);
and U3835 (N_3835,N_2300,N_913);
nand U3836 (N_3836,N_2068,N_1273);
nor U3837 (N_3837,N_2392,N_2127);
and U3838 (N_3838,N_1357,N_1824);
or U3839 (N_3839,N_203,N_1722);
and U3840 (N_3840,N_734,N_1405);
xnor U3841 (N_3841,N_238,N_450);
nor U3842 (N_3842,N_1006,N_456);
and U3843 (N_3843,N_1776,N_2485);
nand U3844 (N_3844,N_452,N_2441);
or U3845 (N_3845,N_2395,N_2384);
nand U3846 (N_3846,N_979,N_1288);
nand U3847 (N_3847,N_1980,N_33);
nand U3848 (N_3848,N_1919,N_2356);
nor U3849 (N_3849,N_1376,N_1784);
and U3850 (N_3850,N_1362,N_1370);
nor U3851 (N_3851,N_1291,N_1552);
nor U3852 (N_3852,N_413,N_373);
nand U3853 (N_3853,N_816,N_593);
and U3854 (N_3854,N_1605,N_1665);
or U3855 (N_3855,N_2005,N_1681);
nand U3856 (N_3856,N_2152,N_133);
and U3857 (N_3857,N_867,N_389);
nand U3858 (N_3858,N_1726,N_992);
or U3859 (N_3859,N_522,N_1322);
or U3860 (N_3860,N_1937,N_15);
nor U3861 (N_3861,N_1371,N_1941);
or U3862 (N_3862,N_402,N_246);
nand U3863 (N_3863,N_342,N_420);
nor U3864 (N_3864,N_2108,N_731);
nand U3865 (N_3865,N_2254,N_1142);
nand U3866 (N_3866,N_2256,N_811);
nor U3867 (N_3867,N_1848,N_9);
nor U3868 (N_3868,N_2126,N_1049);
xnor U3869 (N_3869,N_1474,N_154);
nor U3870 (N_3870,N_1511,N_2368);
or U3871 (N_3871,N_1680,N_2410);
nand U3872 (N_3872,N_2492,N_847);
nor U3873 (N_3873,N_1859,N_130);
nand U3874 (N_3874,N_2401,N_2244);
nor U3875 (N_3875,N_210,N_1206);
nand U3876 (N_3876,N_88,N_1564);
nand U3877 (N_3877,N_1773,N_15);
or U3878 (N_3878,N_1075,N_459);
and U3879 (N_3879,N_538,N_1012);
and U3880 (N_3880,N_1683,N_1810);
nor U3881 (N_3881,N_1527,N_737);
nor U3882 (N_3882,N_558,N_501);
and U3883 (N_3883,N_471,N_2329);
and U3884 (N_3884,N_1417,N_132);
nand U3885 (N_3885,N_1479,N_205);
nand U3886 (N_3886,N_2092,N_1123);
and U3887 (N_3887,N_120,N_978);
nor U3888 (N_3888,N_49,N_16);
or U3889 (N_3889,N_88,N_574);
or U3890 (N_3890,N_1680,N_1959);
or U3891 (N_3891,N_1803,N_2142);
and U3892 (N_3892,N_186,N_1104);
and U3893 (N_3893,N_831,N_1852);
nand U3894 (N_3894,N_360,N_2221);
and U3895 (N_3895,N_1035,N_1428);
nor U3896 (N_3896,N_75,N_1349);
nor U3897 (N_3897,N_2427,N_1002);
nand U3898 (N_3898,N_584,N_2307);
nor U3899 (N_3899,N_140,N_1085);
nor U3900 (N_3900,N_64,N_1861);
or U3901 (N_3901,N_741,N_2305);
and U3902 (N_3902,N_2143,N_1398);
and U3903 (N_3903,N_667,N_1037);
and U3904 (N_3904,N_1466,N_698);
and U3905 (N_3905,N_1753,N_5);
nand U3906 (N_3906,N_1351,N_517);
nor U3907 (N_3907,N_2096,N_978);
or U3908 (N_3908,N_1374,N_1193);
and U3909 (N_3909,N_2094,N_438);
and U3910 (N_3910,N_911,N_843);
nand U3911 (N_3911,N_2297,N_2231);
nand U3912 (N_3912,N_2120,N_172);
and U3913 (N_3913,N_34,N_601);
nand U3914 (N_3914,N_1956,N_1896);
nand U3915 (N_3915,N_2022,N_1603);
or U3916 (N_3916,N_1591,N_1302);
nand U3917 (N_3917,N_768,N_989);
nand U3918 (N_3918,N_904,N_2116);
nand U3919 (N_3919,N_994,N_1030);
nor U3920 (N_3920,N_1758,N_20);
or U3921 (N_3921,N_463,N_1494);
and U3922 (N_3922,N_1352,N_1151);
and U3923 (N_3923,N_1280,N_1189);
or U3924 (N_3924,N_372,N_339);
and U3925 (N_3925,N_1956,N_343);
and U3926 (N_3926,N_1478,N_2174);
nor U3927 (N_3927,N_2478,N_1565);
or U3928 (N_3928,N_802,N_2112);
nand U3929 (N_3929,N_1140,N_293);
nand U3930 (N_3930,N_557,N_2345);
nor U3931 (N_3931,N_1268,N_1227);
nor U3932 (N_3932,N_2368,N_1138);
and U3933 (N_3933,N_1635,N_1996);
and U3934 (N_3934,N_1506,N_41);
or U3935 (N_3935,N_2064,N_363);
and U3936 (N_3936,N_11,N_729);
nand U3937 (N_3937,N_1406,N_323);
and U3938 (N_3938,N_1705,N_84);
or U3939 (N_3939,N_998,N_229);
nor U3940 (N_3940,N_750,N_237);
or U3941 (N_3941,N_345,N_2237);
or U3942 (N_3942,N_1012,N_65);
nor U3943 (N_3943,N_6,N_1332);
or U3944 (N_3944,N_2335,N_897);
nor U3945 (N_3945,N_1018,N_1593);
nor U3946 (N_3946,N_491,N_63);
or U3947 (N_3947,N_1295,N_2372);
and U3948 (N_3948,N_464,N_2485);
and U3949 (N_3949,N_1146,N_204);
or U3950 (N_3950,N_201,N_1957);
nand U3951 (N_3951,N_1464,N_1022);
and U3952 (N_3952,N_2453,N_1489);
nand U3953 (N_3953,N_1389,N_935);
nand U3954 (N_3954,N_119,N_2305);
or U3955 (N_3955,N_1555,N_1914);
nor U3956 (N_3956,N_1968,N_1818);
nand U3957 (N_3957,N_1403,N_368);
or U3958 (N_3958,N_1129,N_2405);
and U3959 (N_3959,N_2213,N_696);
nor U3960 (N_3960,N_186,N_1964);
nor U3961 (N_3961,N_2084,N_592);
nor U3962 (N_3962,N_2037,N_1645);
or U3963 (N_3963,N_201,N_2253);
and U3964 (N_3964,N_536,N_1540);
nor U3965 (N_3965,N_648,N_1445);
nand U3966 (N_3966,N_1312,N_1563);
or U3967 (N_3967,N_1332,N_687);
and U3968 (N_3968,N_422,N_1243);
nand U3969 (N_3969,N_2170,N_452);
and U3970 (N_3970,N_1715,N_1614);
nand U3971 (N_3971,N_210,N_1384);
or U3972 (N_3972,N_1201,N_128);
or U3973 (N_3973,N_532,N_1973);
nor U3974 (N_3974,N_566,N_2299);
nand U3975 (N_3975,N_2273,N_1378);
nor U3976 (N_3976,N_1123,N_1016);
nand U3977 (N_3977,N_2221,N_331);
nand U3978 (N_3978,N_1983,N_2054);
nor U3979 (N_3979,N_393,N_2180);
and U3980 (N_3980,N_2156,N_141);
and U3981 (N_3981,N_204,N_1026);
nand U3982 (N_3982,N_1856,N_415);
nand U3983 (N_3983,N_1585,N_747);
or U3984 (N_3984,N_705,N_1904);
nand U3985 (N_3985,N_1837,N_1963);
nor U3986 (N_3986,N_1417,N_614);
or U3987 (N_3987,N_90,N_362);
nor U3988 (N_3988,N_982,N_1414);
or U3989 (N_3989,N_932,N_1787);
or U3990 (N_3990,N_1326,N_1011);
or U3991 (N_3991,N_1363,N_2142);
nor U3992 (N_3992,N_2422,N_1195);
and U3993 (N_3993,N_2082,N_1733);
or U3994 (N_3994,N_1206,N_346);
nand U3995 (N_3995,N_437,N_2293);
or U3996 (N_3996,N_2152,N_976);
nor U3997 (N_3997,N_1339,N_2010);
or U3998 (N_3998,N_899,N_2078);
nor U3999 (N_3999,N_2420,N_117);
nor U4000 (N_4000,N_2065,N_102);
nand U4001 (N_4001,N_2495,N_811);
nor U4002 (N_4002,N_955,N_1532);
nor U4003 (N_4003,N_281,N_829);
nand U4004 (N_4004,N_770,N_155);
nor U4005 (N_4005,N_684,N_2261);
or U4006 (N_4006,N_1071,N_1102);
nor U4007 (N_4007,N_1076,N_290);
nor U4008 (N_4008,N_292,N_1963);
or U4009 (N_4009,N_737,N_615);
nor U4010 (N_4010,N_16,N_1577);
or U4011 (N_4011,N_1109,N_2221);
and U4012 (N_4012,N_1744,N_1500);
or U4013 (N_4013,N_465,N_1945);
and U4014 (N_4014,N_2315,N_2350);
nand U4015 (N_4015,N_414,N_2087);
nand U4016 (N_4016,N_13,N_2178);
and U4017 (N_4017,N_2403,N_2346);
nand U4018 (N_4018,N_2465,N_156);
and U4019 (N_4019,N_1383,N_1182);
nand U4020 (N_4020,N_2309,N_2261);
nand U4021 (N_4021,N_1264,N_2404);
nand U4022 (N_4022,N_2399,N_667);
or U4023 (N_4023,N_1907,N_2490);
and U4024 (N_4024,N_415,N_1867);
or U4025 (N_4025,N_1379,N_789);
and U4026 (N_4026,N_388,N_515);
nand U4027 (N_4027,N_2435,N_2346);
or U4028 (N_4028,N_158,N_430);
or U4029 (N_4029,N_988,N_1820);
or U4030 (N_4030,N_281,N_1477);
or U4031 (N_4031,N_804,N_2239);
and U4032 (N_4032,N_165,N_2007);
or U4033 (N_4033,N_2388,N_888);
and U4034 (N_4034,N_395,N_2167);
nor U4035 (N_4035,N_1209,N_86);
xor U4036 (N_4036,N_739,N_287);
nor U4037 (N_4037,N_211,N_1764);
nor U4038 (N_4038,N_914,N_382);
nand U4039 (N_4039,N_1370,N_2216);
and U4040 (N_4040,N_1584,N_1297);
or U4041 (N_4041,N_2343,N_2052);
nand U4042 (N_4042,N_6,N_546);
or U4043 (N_4043,N_284,N_2404);
xor U4044 (N_4044,N_301,N_894);
or U4045 (N_4045,N_1515,N_148);
or U4046 (N_4046,N_1466,N_1157);
nor U4047 (N_4047,N_794,N_1707);
and U4048 (N_4048,N_2428,N_2380);
and U4049 (N_4049,N_153,N_915);
nand U4050 (N_4050,N_2263,N_880);
or U4051 (N_4051,N_2300,N_1196);
nand U4052 (N_4052,N_2407,N_2316);
or U4053 (N_4053,N_2152,N_1873);
and U4054 (N_4054,N_955,N_210);
nand U4055 (N_4055,N_890,N_662);
or U4056 (N_4056,N_205,N_2078);
nand U4057 (N_4057,N_1706,N_449);
nand U4058 (N_4058,N_384,N_2416);
or U4059 (N_4059,N_112,N_1121);
xor U4060 (N_4060,N_1031,N_1953);
and U4061 (N_4061,N_432,N_1415);
nor U4062 (N_4062,N_915,N_788);
and U4063 (N_4063,N_340,N_1159);
nand U4064 (N_4064,N_411,N_124);
nor U4065 (N_4065,N_2139,N_1364);
and U4066 (N_4066,N_2185,N_41);
or U4067 (N_4067,N_1302,N_2411);
and U4068 (N_4068,N_1525,N_892);
nor U4069 (N_4069,N_1278,N_1201);
or U4070 (N_4070,N_1436,N_2370);
nor U4071 (N_4071,N_2075,N_2435);
or U4072 (N_4072,N_612,N_346);
nand U4073 (N_4073,N_302,N_1185);
nor U4074 (N_4074,N_1057,N_635);
and U4075 (N_4075,N_980,N_2072);
nor U4076 (N_4076,N_2428,N_226);
or U4077 (N_4077,N_2269,N_1784);
nand U4078 (N_4078,N_320,N_66);
nand U4079 (N_4079,N_2117,N_970);
or U4080 (N_4080,N_2033,N_2037);
or U4081 (N_4081,N_1309,N_473);
and U4082 (N_4082,N_30,N_50);
xnor U4083 (N_4083,N_1353,N_1148);
or U4084 (N_4084,N_249,N_266);
and U4085 (N_4085,N_1272,N_1576);
and U4086 (N_4086,N_488,N_1332);
or U4087 (N_4087,N_1016,N_2165);
or U4088 (N_4088,N_1309,N_1369);
nor U4089 (N_4089,N_2145,N_2073);
or U4090 (N_4090,N_2220,N_518);
nor U4091 (N_4091,N_1793,N_1897);
and U4092 (N_4092,N_1147,N_1402);
nand U4093 (N_4093,N_1248,N_2342);
nor U4094 (N_4094,N_1651,N_677);
and U4095 (N_4095,N_1335,N_1911);
and U4096 (N_4096,N_279,N_1030);
or U4097 (N_4097,N_1513,N_44);
nor U4098 (N_4098,N_1918,N_1217);
nor U4099 (N_4099,N_2214,N_2093);
nand U4100 (N_4100,N_1384,N_329);
nor U4101 (N_4101,N_1524,N_2116);
nand U4102 (N_4102,N_1038,N_1652);
nor U4103 (N_4103,N_6,N_909);
and U4104 (N_4104,N_1918,N_360);
xnor U4105 (N_4105,N_146,N_856);
or U4106 (N_4106,N_881,N_310);
nor U4107 (N_4107,N_1533,N_1246);
nor U4108 (N_4108,N_1327,N_1127);
nor U4109 (N_4109,N_2268,N_370);
nor U4110 (N_4110,N_2439,N_246);
and U4111 (N_4111,N_2072,N_345);
nand U4112 (N_4112,N_2164,N_2003);
and U4113 (N_4113,N_1490,N_508);
and U4114 (N_4114,N_2082,N_638);
or U4115 (N_4115,N_2281,N_1299);
and U4116 (N_4116,N_859,N_264);
and U4117 (N_4117,N_2336,N_203);
nor U4118 (N_4118,N_185,N_333);
or U4119 (N_4119,N_1558,N_1801);
nand U4120 (N_4120,N_1282,N_1036);
nand U4121 (N_4121,N_738,N_1308);
nand U4122 (N_4122,N_860,N_989);
or U4123 (N_4123,N_963,N_624);
nand U4124 (N_4124,N_1466,N_1876);
and U4125 (N_4125,N_1738,N_1385);
and U4126 (N_4126,N_1614,N_110);
nand U4127 (N_4127,N_1621,N_2240);
and U4128 (N_4128,N_2452,N_2183);
and U4129 (N_4129,N_2237,N_1256);
nor U4130 (N_4130,N_1059,N_2048);
nor U4131 (N_4131,N_1625,N_1613);
and U4132 (N_4132,N_2131,N_940);
xnor U4133 (N_4133,N_12,N_44);
and U4134 (N_4134,N_1422,N_1738);
nor U4135 (N_4135,N_79,N_1595);
nand U4136 (N_4136,N_957,N_445);
or U4137 (N_4137,N_699,N_1988);
nand U4138 (N_4138,N_1814,N_1347);
nand U4139 (N_4139,N_1562,N_1622);
and U4140 (N_4140,N_2419,N_73);
nand U4141 (N_4141,N_2119,N_215);
nor U4142 (N_4142,N_650,N_2153);
and U4143 (N_4143,N_76,N_1566);
or U4144 (N_4144,N_294,N_1090);
nand U4145 (N_4145,N_2170,N_504);
nor U4146 (N_4146,N_2498,N_1830);
or U4147 (N_4147,N_258,N_1147);
nor U4148 (N_4148,N_2155,N_1192);
nand U4149 (N_4149,N_1753,N_1955);
and U4150 (N_4150,N_1546,N_1207);
nor U4151 (N_4151,N_1675,N_2429);
nor U4152 (N_4152,N_2200,N_2138);
and U4153 (N_4153,N_1409,N_1155);
nor U4154 (N_4154,N_2174,N_1237);
or U4155 (N_4155,N_1900,N_1623);
and U4156 (N_4156,N_23,N_1219);
nor U4157 (N_4157,N_171,N_676);
nor U4158 (N_4158,N_52,N_103);
or U4159 (N_4159,N_27,N_1314);
nand U4160 (N_4160,N_1804,N_1143);
nand U4161 (N_4161,N_649,N_439);
nor U4162 (N_4162,N_949,N_2491);
nand U4163 (N_4163,N_972,N_447);
or U4164 (N_4164,N_124,N_231);
or U4165 (N_4165,N_73,N_186);
or U4166 (N_4166,N_483,N_1958);
and U4167 (N_4167,N_2387,N_851);
and U4168 (N_4168,N_568,N_1041);
nor U4169 (N_4169,N_1807,N_132);
nand U4170 (N_4170,N_584,N_194);
nand U4171 (N_4171,N_73,N_588);
nand U4172 (N_4172,N_350,N_1523);
and U4173 (N_4173,N_1442,N_748);
or U4174 (N_4174,N_433,N_1686);
and U4175 (N_4175,N_1773,N_1273);
nor U4176 (N_4176,N_1375,N_122);
and U4177 (N_4177,N_315,N_632);
nand U4178 (N_4178,N_329,N_21);
or U4179 (N_4179,N_68,N_2106);
or U4180 (N_4180,N_105,N_56);
and U4181 (N_4181,N_838,N_230);
nand U4182 (N_4182,N_876,N_1872);
nand U4183 (N_4183,N_489,N_1803);
nand U4184 (N_4184,N_356,N_1586);
nand U4185 (N_4185,N_2386,N_1189);
xor U4186 (N_4186,N_1516,N_913);
or U4187 (N_4187,N_1586,N_292);
and U4188 (N_4188,N_226,N_1115);
nor U4189 (N_4189,N_1329,N_595);
and U4190 (N_4190,N_2473,N_49);
nand U4191 (N_4191,N_1220,N_511);
and U4192 (N_4192,N_361,N_808);
or U4193 (N_4193,N_43,N_959);
or U4194 (N_4194,N_1532,N_902);
or U4195 (N_4195,N_2084,N_2286);
nor U4196 (N_4196,N_1895,N_81);
nor U4197 (N_4197,N_1383,N_1246);
nor U4198 (N_4198,N_1971,N_1797);
and U4199 (N_4199,N_1932,N_1422);
nand U4200 (N_4200,N_931,N_1032);
nand U4201 (N_4201,N_1446,N_947);
or U4202 (N_4202,N_567,N_1119);
or U4203 (N_4203,N_1047,N_499);
or U4204 (N_4204,N_252,N_505);
nand U4205 (N_4205,N_2475,N_2361);
nor U4206 (N_4206,N_1351,N_2057);
and U4207 (N_4207,N_175,N_2029);
or U4208 (N_4208,N_2409,N_1346);
nor U4209 (N_4209,N_1573,N_1738);
or U4210 (N_4210,N_1062,N_1730);
nor U4211 (N_4211,N_2476,N_12);
nand U4212 (N_4212,N_365,N_1391);
nand U4213 (N_4213,N_1447,N_680);
or U4214 (N_4214,N_198,N_1238);
nand U4215 (N_4215,N_1703,N_2335);
and U4216 (N_4216,N_230,N_1297);
nand U4217 (N_4217,N_304,N_2062);
nand U4218 (N_4218,N_387,N_2415);
nor U4219 (N_4219,N_839,N_1427);
nor U4220 (N_4220,N_300,N_1300);
nand U4221 (N_4221,N_1223,N_1003);
and U4222 (N_4222,N_1371,N_1317);
nand U4223 (N_4223,N_82,N_715);
nor U4224 (N_4224,N_466,N_1079);
nand U4225 (N_4225,N_270,N_182);
and U4226 (N_4226,N_847,N_917);
or U4227 (N_4227,N_2321,N_1868);
and U4228 (N_4228,N_1129,N_1694);
or U4229 (N_4229,N_1979,N_823);
and U4230 (N_4230,N_2046,N_750);
and U4231 (N_4231,N_1643,N_1957);
nand U4232 (N_4232,N_478,N_1061);
nor U4233 (N_4233,N_1414,N_428);
nor U4234 (N_4234,N_615,N_1579);
nor U4235 (N_4235,N_1033,N_30);
nor U4236 (N_4236,N_1105,N_257);
and U4237 (N_4237,N_1405,N_1335);
nand U4238 (N_4238,N_1620,N_2427);
nand U4239 (N_4239,N_430,N_1816);
nor U4240 (N_4240,N_464,N_481);
or U4241 (N_4241,N_333,N_2298);
or U4242 (N_4242,N_1016,N_1462);
and U4243 (N_4243,N_146,N_1666);
and U4244 (N_4244,N_852,N_1434);
or U4245 (N_4245,N_934,N_2088);
or U4246 (N_4246,N_1632,N_2029);
and U4247 (N_4247,N_2432,N_1635);
and U4248 (N_4248,N_2195,N_2244);
and U4249 (N_4249,N_1342,N_1187);
and U4250 (N_4250,N_1824,N_1723);
nand U4251 (N_4251,N_373,N_1371);
nor U4252 (N_4252,N_2273,N_811);
nand U4253 (N_4253,N_170,N_549);
nand U4254 (N_4254,N_1217,N_761);
and U4255 (N_4255,N_1858,N_2274);
and U4256 (N_4256,N_1237,N_500);
and U4257 (N_4257,N_1014,N_2303);
nand U4258 (N_4258,N_684,N_1507);
or U4259 (N_4259,N_346,N_903);
or U4260 (N_4260,N_108,N_2399);
or U4261 (N_4261,N_847,N_279);
nor U4262 (N_4262,N_158,N_110);
nand U4263 (N_4263,N_2308,N_53);
nor U4264 (N_4264,N_272,N_657);
nand U4265 (N_4265,N_2267,N_1889);
or U4266 (N_4266,N_1695,N_191);
nor U4267 (N_4267,N_1392,N_1261);
and U4268 (N_4268,N_2312,N_805);
and U4269 (N_4269,N_2429,N_949);
and U4270 (N_4270,N_965,N_494);
nor U4271 (N_4271,N_2207,N_1681);
and U4272 (N_4272,N_1864,N_852);
nor U4273 (N_4273,N_800,N_1660);
nor U4274 (N_4274,N_2432,N_863);
nand U4275 (N_4275,N_1901,N_1267);
nor U4276 (N_4276,N_1736,N_2444);
nand U4277 (N_4277,N_1187,N_1114);
and U4278 (N_4278,N_400,N_952);
nor U4279 (N_4279,N_689,N_695);
or U4280 (N_4280,N_1185,N_564);
or U4281 (N_4281,N_636,N_135);
nand U4282 (N_4282,N_1892,N_2461);
and U4283 (N_4283,N_1329,N_2226);
nor U4284 (N_4284,N_267,N_1508);
and U4285 (N_4285,N_1486,N_1836);
and U4286 (N_4286,N_245,N_1240);
nor U4287 (N_4287,N_481,N_831);
or U4288 (N_4288,N_1769,N_1171);
and U4289 (N_4289,N_2109,N_512);
or U4290 (N_4290,N_1306,N_732);
and U4291 (N_4291,N_809,N_2082);
or U4292 (N_4292,N_1874,N_2250);
nor U4293 (N_4293,N_478,N_2294);
or U4294 (N_4294,N_600,N_19);
and U4295 (N_4295,N_1759,N_148);
nand U4296 (N_4296,N_1790,N_2019);
nor U4297 (N_4297,N_793,N_1946);
or U4298 (N_4298,N_1614,N_782);
and U4299 (N_4299,N_2442,N_592);
and U4300 (N_4300,N_242,N_1525);
nor U4301 (N_4301,N_790,N_2173);
and U4302 (N_4302,N_2266,N_231);
or U4303 (N_4303,N_1104,N_739);
nor U4304 (N_4304,N_609,N_208);
nand U4305 (N_4305,N_425,N_485);
and U4306 (N_4306,N_1214,N_997);
xnor U4307 (N_4307,N_1961,N_712);
nor U4308 (N_4308,N_954,N_1314);
or U4309 (N_4309,N_1297,N_1097);
and U4310 (N_4310,N_1233,N_949);
or U4311 (N_4311,N_1860,N_59);
nor U4312 (N_4312,N_2280,N_882);
nand U4313 (N_4313,N_2396,N_2108);
nand U4314 (N_4314,N_320,N_1156);
nor U4315 (N_4315,N_983,N_2019);
or U4316 (N_4316,N_326,N_1361);
or U4317 (N_4317,N_305,N_2105);
and U4318 (N_4318,N_2482,N_2119);
nand U4319 (N_4319,N_1119,N_1185);
nor U4320 (N_4320,N_1857,N_2173);
and U4321 (N_4321,N_2127,N_1420);
nand U4322 (N_4322,N_1396,N_1664);
or U4323 (N_4323,N_1521,N_1115);
or U4324 (N_4324,N_1402,N_787);
nor U4325 (N_4325,N_537,N_54);
nand U4326 (N_4326,N_1557,N_1867);
nor U4327 (N_4327,N_2200,N_296);
and U4328 (N_4328,N_356,N_671);
nor U4329 (N_4329,N_1285,N_1808);
nor U4330 (N_4330,N_1188,N_672);
nand U4331 (N_4331,N_1338,N_2227);
and U4332 (N_4332,N_2185,N_1573);
or U4333 (N_4333,N_722,N_1371);
nor U4334 (N_4334,N_22,N_905);
nand U4335 (N_4335,N_80,N_1231);
nor U4336 (N_4336,N_1665,N_1462);
xor U4337 (N_4337,N_1243,N_1748);
and U4338 (N_4338,N_1464,N_997);
and U4339 (N_4339,N_832,N_1333);
nor U4340 (N_4340,N_2097,N_713);
nor U4341 (N_4341,N_1608,N_1845);
nor U4342 (N_4342,N_470,N_1539);
nor U4343 (N_4343,N_213,N_2320);
and U4344 (N_4344,N_1409,N_1817);
and U4345 (N_4345,N_2170,N_624);
nand U4346 (N_4346,N_2043,N_1127);
or U4347 (N_4347,N_1136,N_2079);
or U4348 (N_4348,N_224,N_469);
or U4349 (N_4349,N_1310,N_94);
nand U4350 (N_4350,N_249,N_280);
nor U4351 (N_4351,N_816,N_623);
nor U4352 (N_4352,N_146,N_369);
and U4353 (N_4353,N_1048,N_1728);
or U4354 (N_4354,N_2241,N_753);
or U4355 (N_4355,N_216,N_1447);
or U4356 (N_4356,N_99,N_1116);
nand U4357 (N_4357,N_408,N_2208);
nor U4358 (N_4358,N_266,N_1828);
or U4359 (N_4359,N_552,N_1571);
or U4360 (N_4360,N_1855,N_62);
xnor U4361 (N_4361,N_689,N_1974);
and U4362 (N_4362,N_1744,N_500);
nand U4363 (N_4363,N_2150,N_406);
or U4364 (N_4364,N_577,N_154);
nand U4365 (N_4365,N_335,N_991);
and U4366 (N_4366,N_269,N_1224);
nand U4367 (N_4367,N_1000,N_1495);
nor U4368 (N_4368,N_2010,N_1013);
nor U4369 (N_4369,N_1475,N_124);
nand U4370 (N_4370,N_2046,N_1505);
or U4371 (N_4371,N_2116,N_1858);
nand U4372 (N_4372,N_689,N_768);
and U4373 (N_4373,N_158,N_860);
and U4374 (N_4374,N_2150,N_2071);
or U4375 (N_4375,N_2334,N_1548);
and U4376 (N_4376,N_1395,N_1265);
nand U4377 (N_4377,N_688,N_2010);
nor U4378 (N_4378,N_1486,N_1581);
nand U4379 (N_4379,N_1733,N_1800);
nor U4380 (N_4380,N_1719,N_2283);
nor U4381 (N_4381,N_1539,N_307);
nor U4382 (N_4382,N_213,N_1685);
and U4383 (N_4383,N_2158,N_991);
or U4384 (N_4384,N_56,N_2492);
or U4385 (N_4385,N_1280,N_1661);
nor U4386 (N_4386,N_1381,N_2223);
and U4387 (N_4387,N_1736,N_2215);
nor U4388 (N_4388,N_810,N_1074);
and U4389 (N_4389,N_1310,N_1115);
and U4390 (N_4390,N_1483,N_1879);
nor U4391 (N_4391,N_1966,N_1589);
nor U4392 (N_4392,N_1613,N_1496);
or U4393 (N_4393,N_2399,N_1869);
nor U4394 (N_4394,N_1610,N_249);
or U4395 (N_4395,N_113,N_1545);
nand U4396 (N_4396,N_1611,N_872);
and U4397 (N_4397,N_1368,N_1963);
or U4398 (N_4398,N_992,N_1896);
nand U4399 (N_4399,N_1052,N_2424);
nand U4400 (N_4400,N_422,N_2211);
nand U4401 (N_4401,N_146,N_536);
nor U4402 (N_4402,N_187,N_582);
and U4403 (N_4403,N_1136,N_2198);
nor U4404 (N_4404,N_639,N_1711);
and U4405 (N_4405,N_1505,N_2281);
nor U4406 (N_4406,N_296,N_1181);
xor U4407 (N_4407,N_1673,N_1967);
nand U4408 (N_4408,N_1156,N_2240);
or U4409 (N_4409,N_1168,N_364);
nor U4410 (N_4410,N_596,N_899);
or U4411 (N_4411,N_51,N_2110);
and U4412 (N_4412,N_778,N_2090);
nand U4413 (N_4413,N_1208,N_608);
or U4414 (N_4414,N_119,N_1729);
or U4415 (N_4415,N_767,N_2019);
or U4416 (N_4416,N_1579,N_1519);
nand U4417 (N_4417,N_1831,N_2222);
and U4418 (N_4418,N_495,N_1106);
nand U4419 (N_4419,N_897,N_1525);
nor U4420 (N_4420,N_1887,N_1729);
nor U4421 (N_4421,N_1023,N_1);
nand U4422 (N_4422,N_387,N_1180);
and U4423 (N_4423,N_1545,N_1248);
or U4424 (N_4424,N_505,N_2494);
nand U4425 (N_4425,N_2262,N_6);
and U4426 (N_4426,N_1106,N_785);
and U4427 (N_4427,N_1152,N_722);
nand U4428 (N_4428,N_1816,N_544);
or U4429 (N_4429,N_1453,N_1942);
nand U4430 (N_4430,N_2119,N_73);
or U4431 (N_4431,N_2381,N_1881);
or U4432 (N_4432,N_1998,N_1522);
nor U4433 (N_4433,N_190,N_1805);
and U4434 (N_4434,N_1120,N_907);
and U4435 (N_4435,N_523,N_681);
and U4436 (N_4436,N_2069,N_880);
and U4437 (N_4437,N_1177,N_2344);
and U4438 (N_4438,N_1868,N_561);
and U4439 (N_4439,N_2125,N_2305);
nor U4440 (N_4440,N_1323,N_1262);
or U4441 (N_4441,N_2092,N_793);
nor U4442 (N_4442,N_700,N_734);
or U4443 (N_4443,N_2418,N_589);
nor U4444 (N_4444,N_1564,N_1046);
and U4445 (N_4445,N_2382,N_1879);
nand U4446 (N_4446,N_197,N_9);
nand U4447 (N_4447,N_379,N_2017);
nand U4448 (N_4448,N_1312,N_476);
and U4449 (N_4449,N_487,N_1782);
nand U4450 (N_4450,N_38,N_1659);
nand U4451 (N_4451,N_1315,N_2315);
nand U4452 (N_4452,N_211,N_982);
nor U4453 (N_4453,N_1152,N_1428);
or U4454 (N_4454,N_2268,N_1631);
nor U4455 (N_4455,N_1546,N_730);
and U4456 (N_4456,N_2087,N_1591);
nand U4457 (N_4457,N_672,N_1559);
and U4458 (N_4458,N_1192,N_1240);
and U4459 (N_4459,N_2040,N_1774);
nand U4460 (N_4460,N_544,N_1401);
nor U4461 (N_4461,N_1632,N_2097);
and U4462 (N_4462,N_1130,N_2199);
nor U4463 (N_4463,N_1025,N_1075);
or U4464 (N_4464,N_92,N_2411);
and U4465 (N_4465,N_912,N_1959);
nand U4466 (N_4466,N_673,N_2400);
and U4467 (N_4467,N_1610,N_997);
nor U4468 (N_4468,N_2238,N_576);
and U4469 (N_4469,N_403,N_1474);
nor U4470 (N_4470,N_646,N_413);
nand U4471 (N_4471,N_199,N_998);
nand U4472 (N_4472,N_1146,N_924);
and U4473 (N_4473,N_1989,N_1168);
or U4474 (N_4474,N_466,N_811);
and U4475 (N_4475,N_681,N_1015);
nand U4476 (N_4476,N_2273,N_1916);
nand U4477 (N_4477,N_687,N_157);
nand U4478 (N_4478,N_1735,N_1846);
nand U4479 (N_4479,N_81,N_105);
or U4480 (N_4480,N_1808,N_882);
and U4481 (N_4481,N_1358,N_601);
and U4482 (N_4482,N_304,N_1404);
nor U4483 (N_4483,N_557,N_1004);
nor U4484 (N_4484,N_1406,N_367);
nor U4485 (N_4485,N_2223,N_1065);
nor U4486 (N_4486,N_2227,N_1529);
nand U4487 (N_4487,N_489,N_1192);
or U4488 (N_4488,N_1687,N_727);
nand U4489 (N_4489,N_2025,N_290);
nor U4490 (N_4490,N_1432,N_1593);
nor U4491 (N_4491,N_2486,N_1798);
nand U4492 (N_4492,N_274,N_952);
and U4493 (N_4493,N_1572,N_2482);
nand U4494 (N_4494,N_53,N_2251);
and U4495 (N_4495,N_2104,N_1014);
nand U4496 (N_4496,N_122,N_2051);
and U4497 (N_4497,N_1429,N_1794);
or U4498 (N_4498,N_1515,N_1246);
nor U4499 (N_4499,N_603,N_1374);
and U4500 (N_4500,N_200,N_404);
nand U4501 (N_4501,N_1892,N_1967);
or U4502 (N_4502,N_1074,N_587);
and U4503 (N_4503,N_2169,N_975);
or U4504 (N_4504,N_824,N_1037);
nor U4505 (N_4505,N_1263,N_392);
and U4506 (N_4506,N_2452,N_1597);
and U4507 (N_4507,N_1301,N_2453);
and U4508 (N_4508,N_1864,N_369);
and U4509 (N_4509,N_144,N_675);
nand U4510 (N_4510,N_2263,N_1112);
nor U4511 (N_4511,N_1712,N_1118);
and U4512 (N_4512,N_1362,N_305);
nor U4513 (N_4513,N_170,N_2491);
nor U4514 (N_4514,N_297,N_1211);
nor U4515 (N_4515,N_2399,N_141);
nor U4516 (N_4516,N_2209,N_989);
nor U4517 (N_4517,N_403,N_2299);
or U4518 (N_4518,N_1383,N_936);
or U4519 (N_4519,N_1092,N_950);
or U4520 (N_4520,N_1917,N_1388);
or U4521 (N_4521,N_1257,N_691);
and U4522 (N_4522,N_1839,N_501);
nor U4523 (N_4523,N_642,N_1088);
nand U4524 (N_4524,N_444,N_975);
nor U4525 (N_4525,N_1033,N_855);
and U4526 (N_4526,N_1605,N_1133);
and U4527 (N_4527,N_1220,N_1341);
and U4528 (N_4528,N_179,N_2196);
nand U4529 (N_4529,N_1296,N_1242);
nor U4530 (N_4530,N_1049,N_1295);
or U4531 (N_4531,N_648,N_1254);
nor U4532 (N_4532,N_2434,N_2450);
or U4533 (N_4533,N_380,N_1785);
and U4534 (N_4534,N_458,N_761);
nor U4535 (N_4535,N_802,N_1440);
nor U4536 (N_4536,N_479,N_505);
or U4537 (N_4537,N_2402,N_1966);
nand U4538 (N_4538,N_884,N_1921);
and U4539 (N_4539,N_168,N_2385);
nand U4540 (N_4540,N_1737,N_1274);
or U4541 (N_4541,N_334,N_1718);
nand U4542 (N_4542,N_2032,N_607);
and U4543 (N_4543,N_639,N_1507);
and U4544 (N_4544,N_2207,N_2095);
or U4545 (N_4545,N_2163,N_850);
and U4546 (N_4546,N_1410,N_868);
nand U4547 (N_4547,N_1837,N_1129);
or U4548 (N_4548,N_343,N_172);
nand U4549 (N_4549,N_151,N_2295);
nand U4550 (N_4550,N_794,N_2400);
nand U4551 (N_4551,N_915,N_1849);
and U4552 (N_4552,N_356,N_1700);
nor U4553 (N_4553,N_1815,N_2345);
or U4554 (N_4554,N_1320,N_282);
and U4555 (N_4555,N_1211,N_2491);
nand U4556 (N_4556,N_919,N_1582);
nor U4557 (N_4557,N_1427,N_1248);
nand U4558 (N_4558,N_990,N_1090);
nand U4559 (N_4559,N_1525,N_39);
or U4560 (N_4560,N_1166,N_588);
or U4561 (N_4561,N_1769,N_652);
and U4562 (N_4562,N_1318,N_1456);
and U4563 (N_4563,N_1547,N_939);
or U4564 (N_4564,N_163,N_1378);
nor U4565 (N_4565,N_997,N_2333);
and U4566 (N_4566,N_712,N_2160);
and U4567 (N_4567,N_437,N_1350);
nor U4568 (N_4568,N_2076,N_1920);
and U4569 (N_4569,N_2418,N_449);
or U4570 (N_4570,N_804,N_994);
or U4571 (N_4571,N_2444,N_409);
and U4572 (N_4572,N_487,N_1938);
nand U4573 (N_4573,N_808,N_1670);
and U4574 (N_4574,N_109,N_4);
nand U4575 (N_4575,N_1653,N_1798);
or U4576 (N_4576,N_1199,N_76);
and U4577 (N_4577,N_211,N_877);
and U4578 (N_4578,N_1849,N_192);
nand U4579 (N_4579,N_2031,N_1854);
nor U4580 (N_4580,N_2479,N_1493);
and U4581 (N_4581,N_1604,N_1229);
and U4582 (N_4582,N_693,N_2382);
and U4583 (N_4583,N_2279,N_2459);
and U4584 (N_4584,N_1205,N_1786);
and U4585 (N_4585,N_2317,N_1026);
or U4586 (N_4586,N_756,N_288);
and U4587 (N_4587,N_1728,N_280);
nand U4588 (N_4588,N_1323,N_469);
nor U4589 (N_4589,N_410,N_490);
nand U4590 (N_4590,N_1842,N_975);
or U4591 (N_4591,N_2294,N_1337);
or U4592 (N_4592,N_492,N_1080);
and U4593 (N_4593,N_90,N_199);
and U4594 (N_4594,N_971,N_2213);
and U4595 (N_4595,N_1909,N_1411);
nor U4596 (N_4596,N_557,N_2354);
nand U4597 (N_4597,N_1657,N_1755);
nand U4598 (N_4598,N_459,N_953);
nor U4599 (N_4599,N_2132,N_1393);
nand U4600 (N_4600,N_452,N_1552);
nor U4601 (N_4601,N_1972,N_201);
nor U4602 (N_4602,N_218,N_1975);
and U4603 (N_4603,N_378,N_648);
and U4604 (N_4604,N_2435,N_1308);
nand U4605 (N_4605,N_41,N_1967);
nand U4606 (N_4606,N_42,N_2270);
nor U4607 (N_4607,N_715,N_1198);
xor U4608 (N_4608,N_2270,N_1092);
and U4609 (N_4609,N_2030,N_1162);
nor U4610 (N_4610,N_1720,N_861);
nand U4611 (N_4611,N_219,N_499);
xnor U4612 (N_4612,N_1539,N_1993);
nand U4613 (N_4613,N_1734,N_1965);
or U4614 (N_4614,N_747,N_1920);
and U4615 (N_4615,N_510,N_696);
nor U4616 (N_4616,N_301,N_2013);
or U4617 (N_4617,N_2069,N_1121);
nand U4618 (N_4618,N_1320,N_614);
or U4619 (N_4619,N_703,N_787);
nor U4620 (N_4620,N_2491,N_2022);
nand U4621 (N_4621,N_609,N_1984);
nor U4622 (N_4622,N_1432,N_2374);
nor U4623 (N_4623,N_839,N_1299);
nor U4624 (N_4624,N_2158,N_1027);
or U4625 (N_4625,N_48,N_1053);
nor U4626 (N_4626,N_915,N_1914);
or U4627 (N_4627,N_2225,N_1097);
nand U4628 (N_4628,N_404,N_2195);
nor U4629 (N_4629,N_1121,N_1655);
nor U4630 (N_4630,N_1573,N_2353);
or U4631 (N_4631,N_314,N_471);
and U4632 (N_4632,N_357,N_1128);
and U4633 (N_4633,N_693,N_2021);
nand U4634 (N_4634,N_1801,N_2289);
nand U4635 (N_4635,N_1596,N_444);
nand U4636 (N_4636,N_872,N_1656);
and U4637 (N_4637,N_645,N_896);
nor U4638 (N_4638,N_20,N_516);
nor U4639 (N_4639,N_1384,N_864);
or U4640 (N_4640,N_2296,N_292);
nor U4641 (N_4641,N_438,N_1940);
nor U4642 (N_4642,N_29,N_691);
nand U4643 (N_4643,N_2342,N_922);
or U4644 (N_4644,N_1503,N_1163);
or U4645 (N_4645,N_1749,N_1836);
or U4646 (N_4646,N_122,N_225);
nand U4647 (N_4647,N_1544,N_411);
nor U4648 (N_4648,N_944,N_414);
and U4649 (N_4649,N_548,N_608);
nor U4650 (N_4650,N_2091,N_1327);
and U4651 (N_4651,N_1055,N_209);
nor U4652 (N_4652,N_2062,N_2312);
nor U4653 (N_4653,N_452,N_1440);
and U4654 (N_4654,N_1610,N_1261);
and U4655 (N_4655,N_1010,N_1026);
and U4656 (N_4656,N_1419,N_42);
nand U4657 (N_4657,N_2207,N_688);
or U4658 (N_4658,N_751,N_1072);
and U4659 (N_4659,N_1135,N_85);
nor U4660 (N_4660,N_1979,N_1334);
or U4661 (N_4661,N_90,N_1798);
nor U4662 (N_4662,N_1945,N_30);
or U4663 (N_4663,N_1463,N_1657);
nand U4664 (N_4664,N_247,N_1720);
or U4665 (N_4665,N_756,N_876);
nor U4666 (N_4666,N_123,N_2138);
and U4667 (N_4667,N_123,N_2163);
nor U4668 (N_4668,N_1560,N_1040);
nand U4669 (N_4669,N_1902,N_103);
or U4670 (N_4670,N_2408,N_817);
nor U4671 (N_4671,N_657,N_2336);
nor U4672 (N_4672,N_787,N_1064);
nor U4673 (N_4673,N_2176,N_2341);
nand U4674 (N_4674,N_271,N_1267);
and U4675 (N_4675,N_1582,N_1083);
nor U4676 (N_4676,N_2402,N_1900);
nand U4677 (N_4677,N_655,N_141);
or U4678 (N_4678,N_1856,N_1105);
or U4679 (N_4679,N_271,N_1221);
and U4680 (N_4680,N_804,N_89);
nand U4681 (N_4681,N_2362,N_1080);
nand U4682 (N_4682,N_447,N_833);
and U4683 (N_4683,N_1250,N_1824);
nor U4684 (N_4684,N_1470,N_2217);
nor U4685 (N_4685,N_2322,N_2173);
or U4686 (N_4686,N_1444,N_475);
nor U4687 (N_4687,N_887,N_737);
and U4688 (N_4688,N_1011,N_1647);
or U4689 (N_4689,N_1175,N_1622);
nor U4690 (N_4690,N_215,N_2082);
nand U4691 (N_4691,N_1737,N_1748);
and U4692 (N_4692,N_443,N_1344);
nor U4693 (N_4693,N_12,N_654);
nor U4694 (N_4694,N_2006,N_1732);
or U4695 (N_4695,N_1413,N_1154);
nand U4696 (N_4696,N_1441,N_243);
and U4697 (N_4697,N_1142,N_946);
nand U4698 (N_4698,N_1390,N_530);
nand U4699 (N_4699,N_1894,N_2497);
nor U4700 (N_4700,N_2119,N_1753);
or U4701 (N_4701,N_2017,N_1327);
and U4702 (N_4702,N_1178,N_2031);
and U4703 (N_4703,N_350,N_89);
and U4704 (N_4704,N_1235,N_317);
nor U4705 (N_4705,N_144,N_294);
nor U4706 (N_4706,N_2223,N_2089);
or U4707 (N_4707,N_1452,N_1284);
nand U4708 (N_4708,N_1353,N_173);
nand U4709 (N_4709,N_1109,N_244);
or U4710 (N_4710,N_54,N_561);
nand U4711 (N_4711,N_1053,N_1773);
nand U4712 (N_4712,N_2152,N_1985);
nor U4713 (N_4713,N_1376,N_612);
or U4714 (N_4714,N_1227,N_1529);
nor U4715 (N_4715,N_1621,N_1375);
or U4716 (N_4716,N_2312,N_773);
nor U4717 (N_4717,N_501,N_2170);
nand U4718 (N_4718,N_302,N_1386);
nor U4719 (N_4719,N_614,N_477);
nand U4720 (N_4720,N_382,N_1954);
and U4721 (N_4721,N_715,N_2488);
nand U4722 (N_4722,N_1087,N_1746);
nor U4723 (N_4723,N_457,N_1148);
or U4724 (N_4724,N_327,N_2269);
nor U4725 (N_4725,N_2098,N_1659);
and U4726 (N_4726,N_2006,N_181);
nor U4727 (N_4727,N_1588,N_2253);
nor U4728 (N_4728,N_1107,N_591);
or U4729 (N_4729,N_1603,N_163);
nor U4730 (N_4730,N_22,N_278);
nor U4731 (N_4731,N_2117,N_597);
and U4732 (N_4732,N_2191,N_1230);
or U4733 (N_4733,N_2221,N_995);
nor U4734 (N_4734,N_639,N_1291);
nand U4735 (N_4735,N_1805,N_1872);
and U4736 (N_4736,N_1688,N_239);
or U4737 (N_4737,N_2049,N_1838);
nor U4738 (N_4738,N_13,N_1229);
nor U4739 (N_4739,N_343,N_2266);
nand U4740 (N_4740,N_1339,N_2111);
nand U4741 (N_4741,N_188,N_1711);
or U4742 (N_4742,N_1360,N_580);
nor U4743 (N_4743,N_661,N_693);
or U4744 (N_4744,N_1416,N_1533);
nand U4745 (N_4745,N_836,N_1350);
or U4746 (N_4746,N_1138,N_1925);
nor U4747 (N_4747,N_2080,N_1438);
or U4748 (N_4748,N_462,N_182);
nor U4749 (N_4749,N_803,N_2397);
nand U4750 (N_4750,N_189,N_1019);
or U4751 (N_4751,N_2496,N_2340);
and U4752 (N_4752,N_374,N_1372);
nor U4753 (N_4753,N_2424,N_103);
nand U4754 (N_4754,N_1072,N_1121);
and U4755 (N_4755,N_368,N_585);
nor U4756 (N_4756,N_746,N_821);
and U4757 (N_4757,N_491,N_1851);
or U4758 (N_4758,N_955,N_774);
nor U4759 (N_4759,N_561,N_1097);
nand U4760 (N_4760,N_552,N_1046);
or U4761 (N_4761,N_1308,N_2240);
or U4762 (N_4762,N_2493,N_1685);
and U4763 (N_4763,N_300,N_2393);
or U4764 (N_4764,N_2221,N_1208);
nor U4765 (N_4765,N_2410,N_1182);
or U4766 (N_4766,N_826,N_854);
or U4767 (N_4767,N_163,N_671);
nor U4768 (N_4768,N_1070,N_1757);
nand U4769 (N_4769,N_1383,N_1793);
and U4770 (N_4770,N_1736,N_346);
or U4771 (N_4771,N_1807,N_71);
and U4772 (N_4772,N_1985,N_2428);
nand U4773 (N_4773,N_1768,N_151);
nor U4774 (N_4774,N_1634,N_2108);
nor U4775 (N_4775,N_1284,N_1652);
nand U4776 (N_4776,N_41,N_2226);
and U4777 (N_4777,N_896,N_842);
or U4778 (N_4778,N_504,N_1355);
nand U4779 (N_4779,N_330,N_167);
nand U4780 (N_4780,N_1444,N_2327);
and U4781 (N_4781,N_529,N_2247);
nand U4782 (N_4782,N_695,N_403);
nand U4783 (N_4783,N_934,N_679);
nor U4784 (N_4784,N_412,N_1369);
xor U4785 (N_4785,N_291,N_109);
and U4786 (N_4786,N_933,N_1232);
nor U4787 (N_4787,N_144,N_2473);
or U4788 (N_4788,N_700,N_890);
or U4789 (N_4789,N_293,N_1608);
and U4790 (N_4790,N_218,N_708);
and U4791 (N_4791,N_773,N_534);
nand U4792 (N_4792,N_1254,N_830);
and U4793 (N_4793,N_273,N_661);
nor U4794 (N_4794,N_2286,N_138);
or U4795 (N_4795,N_2446,N_628);
or U4796 (N_4796,N_657,N_1164);
or U4797 (N_4797,N_1287,N_2093);
nand U4798 (N_4798,N_918,N_686);
or U4799 (N_4799,N_2432,N_1174);
and U4800 (N_4800,N_186,N_1120);
nand U4801 (N_4801,N_1415,N_1059);
nand U4802 (N_4802,N_348,N_1696);
and U4803 (N_4803,N_255,N_670);
or U4804 (N_4804,N_392,N_1164);
and U4805 (N_4805,N_552,N_2289);
and U4806 (N_4806,N_1543,N_405);
and U4807 (N_4807,N_162,N_619);
and U4808 (N_4808,N_325,N_1103);
and U4809 (N_4809,N_128,N_148);
nand U4810 (N_4810,N_2446,N_2291);
and U4811 (N_4811,N_1878,N_200);
and U4812 (N_4812,N_1408,N_2405);
or U4813 (N_4813,N_906,N_466);
nor U4814 (N_4814,N_1287,N_225);
and U4815 (N_4815,N_103,N_2133);
nor U4816 (N_4816,N_55,N_1668);
or U4817 (N_4817,N_2108,N_1072);
or U4818 (N_4818,N_728,N_2185);
or U4819 (N_4819,N_722,N_1016);
and U4820 (N_4820,N_1683,N_2226);
or U4821 (N_4821,N_2386,N_125);
nor U4822 (N_4822,N_283,N_1088);
nand U4823 (N_4823,N_112,N_1369);
nor U4824 (N_4824,N_174,N_407);
nor U4825 (N_4825,N_1126,N_1361);
and U4826 (N_4826,N_133,N_1418);
and U4827 (N_4827,N_261,N_2368);
and U4828 (N_4828,N_2187,N_1116);
and U4829 (N_4829,N_1897,N_314);
nand U4830 (N_4830,N_1558,N_1062);
and U4831 (N_4831,N_922,N_740);
or U4832 (N_4832,N_1736,N_190);
or U4833 (N_4833,N_785,N_2293);
or U4834 (N_4834,N_521,N_1053);
nand U4835 (N_4835,N_1683,N_754);
nor U4836 (N_4836,N_557,N_154);
nor U4837 (N_4837,N_1501,N_445);
or U4838 (N_4838,N_1458,N_1876);
and U4839 (N_4839,N_1336,N_2398);
or U4840 (N_4840,N_165,N_1941);
nand U4841 (N_4841,N_692,N_1923);
and U4842 (N_4842,N_1069,N_1258);
or U4843 (N_4843,N_635,N_234);
or U4844 (N_4844,N_326,N_2214);
or U4845 (N_4845,N_1044,N_2111);
nor U4846 (N_4846,N_1898,N_2428);
nor U4847 (N_4847,N_1364,N_227);
or U4848 (N_4848,N_1238,N_1401);
or U4849 (N_4849,N_2011,N_2466);
or U4850 (N_4850,N_1877,N_577);
nor U4851 (N_4851,N_1930,N_1977);
nor U4852 (N_4852,N_609,N_253);
nor U4853 (N_4853,N_1091,N_2346);
nor U4854 (N_4854,N_443,N_1078);
nor U4855 (N_4855,N_331,N_1703);
nor U4856 (N_4856,N_434,N_2414);
nor U4857 (N_4857,N_567,N_1168);
or U4858 (N_4858,N_498,N_1778);
and U4859 (N_4859,N_1830,N_862);
and U4860 (N_4860,N_538,N_303);
nand U4861 (N_4861,N_991,N_1791);
or U4862 (N_4862,N_1246,N_1306);
and U4863 (N_4863,N_1466,N_2019);
or U4864 (N_4864,N_1860,N_1868);
and U4865 (N_4865,N_2321,N_865);
and U4866 (N_4866,N_635,N_2340);
or U4867 (N_4867,N_1132,N_2450);
or U4868 (N_4868,N_1517,N_1323);
nor U4869 (N_4869,N_206,N_847);
nand U4870 (N_4870,N_486,N_689);
nor U4871 (N_4871,N_1180,N_1001);
nor U4872 (N_4872,N_334,N_132);
and U4873 (N_4873,N_2125,N_1764);
or U4874 (N_4874,N_365,N_610);
nand U4875 (N_4875,N_2336,N_1886);
or U4876 (N_4876,N_798,N_2007);
nand U4877 (N_4877,N_2367,N_343);
or U4878 (N_4878,N_1483,N_617);
or U4879 (N_4879,N_1534,N_928);
and U4880 (N_4880,N_640,N_1378);
nand U4881 (N_4881,N_808,N_1692);
and U4882 (N_4882,N_1334,N_1845);
or U4883 (N_4883,N_824,N_1280);
nor U4884 (N_4884,N_1789,N_447);
or U4885 (N_4885,N_2237,N_2232);
and U4886 (N_4886,N_2183,N_506);
nor U4887 (N_4887,N_1908,N_2050);
nand U4888 (N_4888,N_1002,N_1554);
or U4889 (N_4889,N_1454,N_1109);
nand U4890 (N_4890,N_2223,N_315);
or U4891 (N_4891,N_857,N_1977);
nor U4892 (N_4892,N_471,N_208);
nor U4893 (N_4893,N_2206,N_1176);
nor U4894 (N_4894,N_1715,N_2498);
nor U4895 (N_4895,N_1405,N_2100);
and U4896 (N_4896,N_357,N_46);
and U4897 (N_4897,N_2409,N_1210);
or U4898 (N_4898,N_1073,N_2314);
or U4899 (N_4899,N_237,N_1958);
nand U4900 (N_4900,N_398,N_1014);
or U4901 (N_4901,N_122,N_1901);
nor U4902 (N_4902,N_1410,N_864);
and U4903 (N_4903,N_2120,N_577);
or U4904 (N_4904,N_226,N_2010);
xnor U4905 (N_4905,N_2,N_272);
or U4906 (N_4906,N_2479,N_2283);
nand U4907 (N_4907,N_1444,N_1472);
or U4908 (N_4908,N_2297,N_1509);
nand U4909 (N_4909,N_1396,N_2462);
or U4910 (N_4910,N_403,N_12);
or U4911 (N_4911,N_855,N_580);
and U4912 (N_4912,N_2054,N_23);
nor U4913 (N_4913,N_410,N_1635);
nor U4914 (N_4914,N_402,N_646);
or U4915 (N_4915,N_672,N_1033);
nand U4916 (N_4916,N_1440,N_153);
nor U4917 (N_4917,N_2491,N_348);
or U4918 (N_4918,N_31,N_2389);
or U4919 (N_4919,N_1020,N_238);
and U4920 (N_4920,N_1572,N_2128);
nand U4921 (N_4921,N_2415,N_177);
xnor U4922 (N_4922,N_105,N_180);
nor U4923 (N_4923,N_616,N_1248);
or U4924 (N_4924,N_1249,N_2168);
nor U4925 (N_4925,N_385,N_274);
nand U4926 (N_4926,N_1970,N_267);
nor U4927 (N_4927,N_799,N_1179);
and U4928 (N_4928,N_2350,N_374);
or U4929 (N_4929,N_2323,N_1170);
or U4930 (N_4930,N_2491,N_213);
nand U4931 (N_4931,N_1338,N_666);
or U4932 (N_4932,N_614,N_10);
nand U4933 (N_4933,N_1228,N_1670);
nand U4934 (N_4934,N_1087,N_989);
nand U4935 (N_4935,N_966,N_1330);
and U4936 (N_4936,N_944,N_536);
or U4937 (N_4937,N_1492,N_127);
and U4938 (N_4938,N_317,N_498);
and U4939 (N_4939,N_368,N_1982);
nor U4940 (N_4940,N_1076,N_2398);
or U4941 (N_4941,N_2222,N_1011);
and U4942 (N_4942,N_1409,N_1150);
or U4943 (N_4943,N_1258,N_283);
and U4944 (N_4944,N_2152,N_968);
nor U4945 (N_4945,N_90,N_62);
or U4946 (N_4946,N_2168,N_194);
nand U4947 (N_4947,N_1712,N_2321);
nand U4948 (N_4948,N_1466,N_544);
nor U4949 (N_4949,N_6,N_1988);
and U4950 (N_4950,N_460,N_1655);
nor U4951 (N_4951,N_1861,N_489);
or U4952 (N_4952,N_924,N_517);
nor U4953 (N_4953,N_1997,N_463);
nand U4954 (N_4954,N_2129,N_1019);
nor U4955 (N_4955,N_137,N_1901);
nand U4956 (N_4956,N_2111,N_2461);
and U4957 (N_4957,N_1257,N_152);
nor U4958 (N_4958,N_1879,N_1475);
nor U4959 (N_4959,N_707,N_1744);
or U4960 (N_4960,N_1887,N_2066);
nor U4961 (N_4961,N_1257,N_84);
or U4962 (N_4962,N_682,N_2412);
and U4963 (N_4963,N_119,N_1898);
or U4964 (N_4964,N_1850,N_349);
nor U4965 (N_4965,N_957,N_1438);
or U4966 (N_4966,N_295,N_1212);
or U4967 (N_4967,N_123,N_989);
nand U4968 (N_4968,N_1266,N_736);
nor U4969 (N_4969,N_1781,N_454);
nand U4970 (N_4970,N_668,N_73);
nor U4971 (N_4971,N_2380,N_527);
nand U4972 (N_4972,N_1110,N_2094);
nand U4973 (N_4973,N_695,N_719);
nor U4974 (N_4974,N_123,N_1634);
nand U4975 (N_4975,N_2175,N_1338);
and U4976 (N_4976,N_1465,N_2202);
nor U4977 (N_4977,N_2249,N_2027);
nor U4978 (N_4978,N_1251,N_475);
nand U4979 (N_4979,N_2295,N_288);
and U4980 (N_4980,N_1973,N_227);
or U4981 (N_4981,N_1121,N_390);
nand U4982 (N_4982,N_647,N_285);
and U4983 (N_4983,N_1906,N_1606);
or U4984 (N_4984,N_240,N_2107);
or U4985 (N_4985,N_1596,N_1344);
or U4986 (N_4986,N_1174,N_617);
or U4987 (N_4987,N_784,N_505);
nor U4988 (N_4988,N_1778,N_752);
nand U4989 (N_4989,N_1468,N_594);
and U4990 (N_4990,N_116,N_1848);
nor U4991 (N_4991,N_2000,N_854);
nor U4992 (N_4992,N_820,N_1167);
nor U4993 (N_4993,N_809,N_1690);
and U4994 (N_4994,N_1958,N_2066);
xor U4995 (N_4995,N_796,N_104);
and U4996 (N_4996,N_1256,N_315);
and U4997 (N_4997,N_78,N_476);
nor U4998 (N_4998,N_1086,N_252);
nand U4999 (N_4999,N_2235,N_1523);
and UO_0 (O_0,N_3464,N_4496);
nor UO_1 (O_1,N_4401,N_2604);
or UO_2 (O_2,N_4709,N_2767);
nand UO_3 (O_3,N_4142,N_4180);
or UO_4 (O_4,N_3305,N_3971);
or UO_5 (O_5,N_3928,N_3183);
or UO_6 (O_6,N_2684,N_4711);
nor UO_7 (O_7,N_4908,N_2859);
and UO_8 (O_8,N_4697,N_4375);
and UO_9 (O_9,N_4968,N_4706);
nor UO_10 (O_10,N_3722,N_2550);
or UO_11 (O_11,N_4211,N_4845);
and UO_12 (O_12,N_3534,N_2880);
nand UO_13 (O_13,N_2890,N_4194);
and UO_14 (O_14,N_2811,N_4482);
and UO_15 (O_15,N_3871,N_3606);
or UO_16 (O_16,N_4109,N_4485);
nor UO_17 (O_17,N_4251,N_4840);
or UO_18 (O_18,N_4701,N_3345);
nand UO_19 (O_19,N_2957,N_2678);
nand UO_20 (O_20,N_4616,N_3785);
and UO_21 (O_21,N_4869,N_4515);
nor UO_22 (O_22,N_3787,N_4549);
nand UO_23 (O_23,N_3241,N_2938);
and UO_24 (O_24,N_3297,N_3501);
nand UO_25 (O_25,N_2770,N_3993);
and UO_26 (O_26,N_4266,N_4831);
nand UO_27 (O_27,N_4511,N_2706);
nand UO_28 (O_28,N_4034,N_3095);
nor UO_29 (O_29,N_4483,N_3451);
and UO_30 (O_30,N_4976,N_4910);
and UO_31 (O_31,N_3438,N_3261);
nand UO_32 (O_32,N_4795,N_4522);
and UO_33 (O_33,N_3818,N_3576);
nand UO_34 (O_34,N_4823,N_4911);
nand UO_35 (O_35,N_3492,N_4956);
or UO_36 (O_36,N_3022,N_4882);
nor UO_37 (O_37,N_3967,N_4309);
and UO_38 (O_38,N_4407,N_3380);
or UO_39 (O_39,N_3815,N_2705);
nand UO_40 (O_40,N_3639,N_3503);
or UO_41 (O_41,N_3847,N_2873);
nor UO_42 (O_42,N_4978,N_2590);
or UO_43 (O_43,N_4741,N_2662);
nand UO_44 (O_44,N_3891,N_3770);
nand UO_45 (O_45,N_2820,N_4336);
or UO_46 (O_46,N_4565,N_3864);
and UO_47 (O_47,N_4044,N_3560);
and UO_48 (O_48,N_4261,N_4388);
and UO_49 (O_49,N_4271,N_2696);
nand UO_50 (O_50,N_3594,N_3861);
nand UO_51 (O_51,N_4042,N_4045);
or UO_52 (O_52,N_3513,N_4007);
and UO_53 (O_53,N_4439,N_3361);
and UO_54 (O_54,N_4158,N_4775);
nor UO_55 (O_55,N_3514,N_3913);
nand UO_56 (O_56,N_3491,N_3402);
nand UO_57 (O_57,N_4912,N_4416);
nor UO_58 (O_58,N_3349,N_3777);
or UO_59 (O_59,N_4464,N_4051);
or UO_60 (O_60,N_3055,N_4270);
nor UO_61 (O_61,N_3213,N_2986);
and UO_62 (O_62,N_2583,N_3024);
or UO_63 (O_63,N_4433,N_2872);
and UO_64 (O_64,N_4322,N_4521);
and UO_65 (O_65,N_3130,N_2911);
nand UO_66 (O_66,N_3086,N_4133);
and UO_67 (O_67,N_2596,N_3677);
and UO_68 (O_68,N_4806,N_4820);
or UO_69 (O_69,N_4932,N_3121);
nand UO_70 (O_70,N_2742,N_4573);
and UO_71 (O_71,N_4263,N_3564);
and UO_72 (O_72,N_4647,N_4118);
or UO_73 (O_73,N_3131,N_3911);
nor UO_74 (O_74,N_3873,N_4901);
nor UO_75 (O_75,N_4740,N_4591);
and UO_76 (O_76,N_2670,N_4724);
and UO_77 (O_77,N_2850,N_4649);
or UO_78 (O_78,N_3504,N_3552);
nor UO_79 (O_79,N_4644,N_4878);
and UO_80 (O_80,N_4124,N_4112);
and UO_81 (O_81,N_4026,N_2855);
nor UO_82 (O_82,N_4821,N_4449);
and UO_83 (O_83,N_4296,N_3903);
nand UO_84 (O_84,N_2537,N_4989);
nand UO_85 (O_85,N_4499,N_3017);
and UO_86 (O_86,N_4488,N_3869);
and UO_87 (O_87,N_2581,N_2856);
or UO_88 (O_88,N_4577,N_3962);
nand UO_89 (O_89,N_2649,N_4238);
nor UO_90 (O_90,N_2566,N_4964);
and UO_91 (O_91,N_3506,N_3879);
nand UO_92 (O_92,N_2614,N_3217);
and UO_93 (O_93,N_4281,N_2565);
nor UO_94 (O_94,N_4818,N_3343);
nor UO_95 (O_95,N_4279,N_4893);
nand UO_96 (O_96,N_3867,N_2740);
and UO_97 (O_97,N_4224,N_2992);
nand UO_98 (O_98,N_2782,N_4805);
nand UO_99 (O_99,N_4655,N_4606);
and UO_100 (O_100,N_4735,N_3308);
or UO_101 (O_101,N_4484,N_3381);
and UO_102 (O_102,N_4918,N_4313);
nand UO_103 (O_103,N_4207,N_3479);
or UO_104 (O_104,N_3240,N_4021);
and UO_105 (O_105,N_4759,N_4040);
or UO_106 (O_106,N_4345,N_3689);
nor UO_107 (O_107,N_3268,N_2758);
and UO_108 (O_108,N_3748,N_2579);
and UO_109 (O_109,N_2916,N_3754);
nor UO_110 (O_110,N_2936,N_4703);
and UO_111 (O_111,N_4425,N_4877);
or UO_112 (O_112,N_3016,N_3947);
xnor UO_113 (O_113,N_2682,N_2981);
or UO_114 (O_114,N_4039,N_4497);
nor UO_115 (O_115,N_2882,N_4841);
xnor UO_116 (O_116,N_4919,N_3649);
and UO_117 (O_117,N_4272,N_3979);
or UO_118 (O_118,N_2768,N_4122);
and UO_119 (O_119,N_4165,N_2697);
and UO_120 (O_120,N_4786,N_4492);
or UO_121 (O_121,N_3083,N_4922);
nand UO_122 (O_122,N_2704,N_4757);
and UO_123 (O_123,N_4125,N_4405);
or UO_124 (O_124,N_3037,N_4225);
nand UO_125 (O_125,N_4957,N_4063);
or UO_126 (O_126,N_4639,N_4412);
and UO_127 (O_127,N_2954,N_4060);
nand UO_128 (O_128,N_3001,N_3428);
and UO_129 (O_129,N_4787,N_4088);
or UO_130 (O_130,N_4603,N_3811);
nand UO_131 (O_131,N_4372,N_4779);
nor UO_132 (O_132,N_4175,N_2517);
or UO_133 (O_133,N_2750,N_4167);
nand UO_134 (O_134,N_2724,N_4363);
nand UO_135 (O_135,N_4601,N_2774);
nand UO_136 (O_136,N_3535,N_2643);
nand UO_137 (O_137,N_2666,N_3500);
and UO_138 (O_138,N_3419,N_4293);
nor UO_139 (O_139,N_4698,N_2533);
nand UO_140 (O_140,N_2642,N_4092);
nor UO_141 (O_141,N_3398,N_3696);
nand UO_142 (O_142,N_4370,N_4690);
nand UO_143 (O_143,N_3225,N_4410);
nor UO_144 (O_144,N_4982,N_2887);
and UO_145 (O_145,N_4904,N_2645);
nor UO_146 (O_146,N_4460,N_4585);
nor UO_147 (O_147,N_3161,N_4810);
nand UO_148 (O_148,N_4650,N_2549);
or UO_149 (O_149,N_3165,N_3334);
nor UO_150 (O_150,N_3020,N_4065);
or UO_151 (O_151,N_4053,N_2828);
nand UO_152 (O_152,N_3477,N_4012);
and UO_153 (O_153,N_4292,N_4003);
nand UO_154 (O_154,N_4862,N_3846);
nor UO_155 (O_155,N_3294,N_4215);
and UO_156 (O_156,N_4329,N_4500);
nor UO_157 (O_157,N_3484,N_4883);
nand UO_158 (O_158,N_3365,N_3544);
nand UO_159 (O_159,N_3453,N_3030);
nand UO_160 (O_160,N_4835,N_2814);
or UO_161 (O_161,N_3309,N_4994);
and UO_162 (O_162,N_2817,N_3210);
or UO_163 (O_163,N_3283,N_3561);
nor UO_164 (O_164,N_2807,N_4120);
nor UO_165 (O_165,N_2575,N_4283);
nor UO_166 (O_166,N_3949,N_4377);
and UO_167 (O_167,N_4437,N_2840);
and UO_168 (O_168,N_3641,N_4190);
nand UO_169 (O_169,N_3688,N_3863);
and UO_170 (O_170,N_2518,N_3434);
or UO_171 (O_171,N_2679,N_2578);
nor UO_172 (O_172,N_3937,N_3452);
or UO_173 (O_173,N_4632,N_4001);
nand UO_174 (O_174,N_4774,N_2803);
and UO_175 (O_175,N_4229,N_3202);
or UO_176 (O_176,N_4302,N_4260);
and UO_177 (O_177,N_4384,N_3566);
nand UO_178 (O_178,N_4895,N_4733);
and UO_179 (O_179,N_3736,N_2542);
nand UO_180 (O_180,N_4710,N_4570);
and UO_181 (O_181,N_3106,N_3096);
nor UO_182 (O_182,N_4725,N_3609);
and UO_183 (O_183,N_3812,N_4554);
or UO_184 (O_184,N_2528,N_4213);
xnor UO_185 (O_185,N_4974,N_3158);
and UO_186 (O_186,N_4659,N_4239);
and UO_187 (O_187,N_3247,N_3651);
and UO_188 (O_188,N_3836,N_3573);
xnor UO_189 (O_189,N_3321,N_2920);
or UO_190 (O_190,N_4430,N_3973);
or UO_191 (O_191,N_4324,N_3975);
or UO_192 (O_192,N_3068,N_4648);
nand UO_193 (O_193,N_3296,N_4576);
nand UO_194 (O_194,N_4767,N_3344);
and UO_195 (O_195,N_3896,N_4163);
and UO_196 (O_196,N_4590,N_3178);
nor UO_197 (O_197,N_4099,N_2551);
or UO_198 (O_198,N_2931,N_4343);
or UO_199 (O_199,N_4208,N_2910);
and UO_200 (O_200,N_3388,N_4214);
nor UO_201 (O_201,N_2744,N_3528);
nor UO_202 (O_202,N_3264,N_4742);
nor UO_203 (O_203,N_3656,N_4923);
and UO_204 (O_204,N_3745,N_3521);
nand UO_205 (O_205,N_2941,N_4396);
nand UO_206 (O_206,N_4945,N_3642);
nand UO_207 (O_207,N_2854,N_4962);
nor UO_208 (O_208,N_3843,N_4924);
nor UO_209 (O_209,N_3008,N_4609);
nand UO_210 (O_210,N_3422,N_3775);
nor UO_211 (O_211,N_4555,N_3222);
and UO_212 (O_212,N_4427,N_4376);
nor UO_213 (O_213,N_3051,N_4614);
nor UO_214 (O_214,N_2664,N_4716);
nand UO_215 (O_215,N_2563,N_4551);
and UO_216 (O_216,N_4715,N_2624);
nor UO_217 (O_217,N_3821,N_4930);
or UO_218 (O_218,N_4824,N_4816);
nand UO_219 (O_219,N_3760,N_4438);
and UO_220 (O_220,N_4074,N_3723);
and UO_221 (O_221,N_3957,N_4947);
nand UO_222 (O_222,N_4743,N_4838);
nand UO_223 (O_223,N_4385,N_3469);
or UO_224 (O_224,N_3553,N_3667);
or UO_225 (O_225,N_2825,N_2522);
or UO_226 (O_226,N_2857,N_4314);
nand UO_227 (O_227,N_3045,N_3331);
nor UO_228 (O_228,N_4046,N_2504);
and UO_229 (O_229,N_4006,N_2539);
and UO_230 (O_230,N_4894,N_2525);
or UO_231 (O_231,N_3442,N_4332);
and UO_232 (O_232,N_3819,N_4983);
or UO_233 (O_233,N_3483,N_2668);
nor UO_234 (O_234,N_3925,N_3671);
nor UO_235 (O_235,N_4140,N_4135);
nor UO_236 (O_236,N_4749,N_4888);
and UO_237 (O_237,N_3915,N_4847);
nor UO_238 (O_238,N_2714,N_4848);
and UO_239 (O_239,N_4812,N_4571);
and UO_240 (O_240,N_4705,N_3340);
or UO_241 (O_241,N_2646,N_4453);
nand UO_242 (O_242,N_4891,N_3265);
or UO_243 (O_243,N_4282,N_4037);
and UO_244 (O_244,N_4561,N_3946);
or UO_245 (O_245,N_4382,N_3263);
nand UO_246 (O_246,N_4575,N_3885);
nor UO_247 (O_247,N_4646,N_3177);
nand UO_248 (O_248,N_3236,N_3959);
nand UO_249 (O_249,N_3197,N_2901);
nor UO_250 (O_250,N_4326,N_4480);
xnor UO_251 (O_251,N_2636,N_2623);
and UO_252 (O_252,N_4604,N_4665);
nand UO_253 (O_253,N_3341,N_2798);
nand UO_254 (O_254,N_2665,N_3598);
nand UO_255 (O_255,N_3537,N_2589);
nor UO_256 (O_256,N_3989,N_2952);
nand UO_257 (O_257,N_3987,N_3984);
and UO_258 (O_258,N_4274,N_3953);
nor UO_259 (O_259,N_3726,N_3874);
nand UO_260 (O_260,N_4126,N_4955);
nand UO_261 (O_261,N_4052,N_4043);
or UO_262 (O_262,N_4783,N_4720);
nand UO_263 (O_263,N_2996,N_3169);
and UO_264 (O_264,N_3703,N_4971);
and UO_265 (O_265,N_2963,N_3735);
and UO_266 (O_266,N_3599,N_3362);
nor UO_267 (O_267,N_3659,N_4254);
nor UO_268 (O_268,N_4132,N_4247);
nand UO_269 (O_269,N_3548,N_3648);
nor UO_270 (O_270,N_2606,N_4212);
or UO_271 (O_271,N_4714,N_4670);
or UO_272 (O_272,N_3739,N_2779);
and UO_273 (O_273,N_3287,N_4033);
or UO_274 (O_274,N_4512,N_2567);
and UO_275 (O_275,N_4068,N_3123);
or UO_276 (O_276,N_4517,N_4243);
nand UO_277 (O_277,N_4794,N_4938);
nand UO_278 (O_278,N_4630,N_4594);
nand UO_279 (O_279,N_4798,N_3033);
nor UO_280 (O_280,N_3848,N_3729);
or UO_281 (O_281,N_3673,N_2893);
and UO_282 (O_282,N_3112,N_3732);
nor UO_283 (O_283,N_3413,N_2709);
nand UO_284 (O_284,N_4094,N_2757);
nor UO_285 (O_285,N_3851,N_2621);
nand UO_286 (O_286,N_2842,N_4420);
nand UO_287 (O_287,N_3793,N_3881);
and UO_288 (O_288,N_3716,N_4872);
or UO_289 (O_289,N_4490,N_3371);
or UO_290 (O_290,N_2783,N_2659);
nand UO_291 (O_291,N_2634,N_4032);
or UO_292 (O_292,N_2594,N_2677);
nand UO_293 (O_293,N_3808,N_3529);
and UO_294 (O_294,N_2833,N_2672);
or UO_295 (O_295,N_2964,N_3164);
or UO_296 (O_296,N_4530,N_3315);
nand UO_297 (O_297,N_2977,N_4297);
and UO_298 (O_298,N_4807,N_4860);
and UO_299 (O_299,N_2917,N_3618);
nand UO_300 (O_300,N_4117,N_3481);
nor UO_301 (O_301,N_3352,N_3107);
nand UO_302 (O_302,N_3917,N_2797);
nand UO_303 (O_303,N_4258,N_3249);
and UO_304 (O_304,N_3027,N_2681);
or UO_305 (O_305,N_2751,N_4441);
or UO_306 (O_306,N_3212,N_4036);
or UO_307 (O_307,N_4476,N_2710);
and UO_308 (O_308,N_4771,N_3619);
nand UO_309 (O_309,N_4310,N_4389);
nand UO_310 (O_310,N_3424,N_4839);
or UO_311 (O_311,N_4458,N_4093);
and UO_312 (O_312,N_4748,N_4651);
nand UO_313 (O_313,N_3623,N_4149);
nor UO_314 (O_314,N_3224,N_3436);
nor UO_315 (O_315,N_3172,N_3260);
nor UO_316 (O_316,N_2725,N_3731);
nand UO_317 (O_317,N_4641,N_4182);
or UO_318 (O_318,N_4766,N_2719);
or UO_319 (O_319,N_2573,N_3059);
or UO_320 (O_320,N_4726,N_4114);
or UO_321 (O_321,N_3638,N_2552);
nor UO_322 (O_322,N_4965,N_3404);
nor UO_323 (O_323,N_3556,N_3757);
or UO_324 (O_324,N_4568,N_2637);
and UO_325 (O_325,N_2948,N_4455);
or UO_326 (O_326,N_3567,N_3207);
or UO_327 (O_327,N_2547,N_3972);
nand UO_328 (O_328,N_3062,N_4809);
nor UO_329 (O_329,N_4588,N_4546);
and UO_330 (O_330,N_3936,N_3206);
or UO_331 (O_331,N_4231,N_4390);
and UO_332 (O_332,N_4984,N_3718);
and UO_333 (O_333,N_3870,N_3021);
nor UO_334 (O_334,N_4383,N_2657);
and UO_335 (O_335,N_4691,N_3075);
and UO_336 (O_336,N_3565,N_4491);
nand UO_337 (O_337,N_2958,N_4791);
nand UO_338 (O_338,N_2892,N_2946);
and UO_339 (O_339,N_4526,N_3531);
or UO_340 (O_340,N_3216,N_4369);
and UO_341 (O_341,N_4527,N_2739);
and UO_342 (O_342,N_4472,N_4428);
or UO_343 (O_343,N_2876,N_3658);
or UO_344 (O_344,N_4252,N_4284);
nor UO_345 (O_345,N_3295,N_3596);
or UO_346 (O_346,N_4054,N_3052);
nand UO_347 (O_347,N_3546,N_4746);
nor UO_348 (O_348,N_3910,N_4739);
nand UO_349 (O_349,N_3899,N_3789);
nor UO_350 (O_350,N_3683,N_4071);
nand UO_351 (O_351,N_4764,N_4137);
and UO_352 (O_352,N_4150,N_3111);
nor UO_353 (O_353,N_3144,N_4374);
xnor UO_354 (O_354,N_2960,N_3580);
and UO_355 (O_355,N_2804,N_3826);
nor UO_356 (O_356,N_4628,N_2538);
and UO_357 (O_357,N_4223,N_2994);
nand UO_358 (O_358,N_2717,N_2795);
or UO_359 (O_359,N_4334,N_4981);
or UO_360 (O_360,N_3809,N_4990);
nand UO_361 (O_361,N_4347,N_4881);
or UO_362 (O_362,N_3496,N_4879);
nor UO_363 (O_363,N_4654,N_4718);
nor UO_364 (O_364,N_3516,N_3113);
or UO_365 (O_365,N_3640,N_4176);
and UO_366 (O_366,N_3187,N_2592);
or UO_367 (O_367,N_4159,N_4929);
nor UO_368 (O_368,N_4531,N_4304);
nand UO_369 (O_369,N_3983,N_3174);
nand UO_370 (O_370,N_4803,N_3298);
nand UO_371 (O_371,N_3900,N_2712);
and UO_372 (O_372,N_4010,N_4085);
or UO_373 (O_373,N_2867,N_4459);
nand UO_374 (O_374,N_3682,N_2534);
and UO_375 (O_375,N_4379,N_2969);
nor UO_376 (O_376,N_2500,N_3978);
nor UO_377 (O_377,N_4529,N_3833);
nand UO_378 (O_378,N_3200,N_3148);
xor UO_379 (O_379,N_4998,N_2970);
or UO_380 (O_380,N_2937,N_4059);
nand UO_381 (O_381,N_2950,N_2633);
and UO_382 (O_382,N_4465,N_3592);
and UO_383 (O_383,N_4960,N_4935);
and UO_384 (O_384,N_2588,N_3134);
nand UO_385 (O_385,N_3149,N_4269);
nand UO_386 (O_386,N_4095,N_3214);
or UO_387 (O_387,N_4096,N_3319);
nand UO_388 (O_388,N_2685,N_4753);
and UO_389 (O_389,N_4166,N_4867);
nand UO_390 (O_390,N_3525,N_4770);
nand UO_391 (O_391,N_3590,N_2830);
or UO_392 (O_392,N_4975,N_2555);
and UO_393 (O_393,N_3768,N_4752);
or UO_394 (O_394,N_2663,N_4111);
or UO_395 (O_395,N_3088,N_3327);
nor UO_396 (O_396,N_3255,N_4129);
nor UO_397 (O_397,N_4602,N_3125);
or UO_398 (O_398,N_3907,N_2962);
nor UO_399 (O_399,N_3003,N_3154);
nor UO_400 (O_400,N_3737,N_3834);
and UO_401 (O_401,N_2955,N_4466);
or UO_402 (O_402,N_2928,N_3661);
nand UO_403 (O_403,N_4730,N_4552);
or UO_404 (O_404,N_2915,N_3990);
and UO_405 (O_405,N_3796,N_4519);
nand UO_406 (O_406,N_2809,N_2999);
or UO_407 (O_407,N_3932,N_2612);
nor UO_408 (O_408,N_2722,N_3663);
nor UO_409 (O_409,N_4550,N_3244);
or UO_410 (O_410,N_3447,N_4119);
nand UO_411 (O_411,N_4024,N_4198);
nor UO_412 (O_412,N_4950,N_4253);
or UO_413 (O_413,N_4836,N_4676);
nand UO_414 (O_414,N_4744,N_3435);
or UO_415 (O_415,N_4049,N_3390);
and UO_416 (O_416,N_4317,N_3559);
nor UO_417 (O_417,N_4843,N_4168);
nor UO_418 (O_418,N_3524,N_4355);
nor UO_419 (O_419,N_3046,N_3547);
and UO_420 (O_420,N_4429,N_4091);
and UO_421 (O_421,N_3761,N_4327);
nor UO_422 (O_422,N_3935,N_2597);
nand UO_423 (O_423,N_2667,N_3769);
nand UO_424 (O_424,N_3188,N_3968);
nor UO_425 (O_425,N_3281,N_2802);
or UO_426 (O_426,N_2731,N_4184);
nor UO_427 (O_427,N_2847,N_2713);
nor UO_428 (O_428,N_4226,N_4436);
and UO_429 (O_429,N_3539,N_3883);
nor UO_430 (O_430,N_2790,N_3961);
and UO_431 (O_431,N_4341,N_4451);
and UO_432 (O_432,N_4897,N_2919);
and UO_433 (O_433,N_2718,N_4196);
nand UO_434 (O_434,N_4693,N_2998);
nor UO_435 (O_435,N_4855,N_4217);
and UO_436 (O_436,N_4325,N_3880);
nor UO_437 (O_437,N_2843,N_4435);
or UO_438 (O_438,N_4944,N_4335);
nand UO_439 (O_439,N_4344,N_3964);
or UO_440 (O_440,N_4699,N_3747);
and UO_441 (O_441,N_3430,N_2698);
or UO_442 (O_442,N_2647,N_4916);
nor UO_443 (O_443,N_4863,N_2769);
nand UO_444 (O_444,N_2953,N_3952);
nand UO_445 (O_445,N_4853,N_4925);
and UO_446 (O_446,N_3720,N_2985);
or UO_447 (O_447,N_4642,N_4827);
nor UO_448 (O_448,N_4582,N_4751);
or UO_449 (O_449,N_3143,N_2808);
nand UO_450 (O_450,N_3043,N_2516);
nor UO_451 (O_451,N_4536,N_4173);
nand UO_452 (O_452,N_4183,N_3938);
and UO_453 (O_453,N_3969,N_4967);
nand UO_454 (O_454,N_3629,N_2826);
and UO_455 (O_455,N_2568,N_3314);
nor UO_456 (O_456,N_4949,N_4666);
and UO_457 (O_457,N_3470,N_3129);
nor UO_458 (O_458,N_3627,N_4569);
and UO_459 (O_459,N_4444,N_4909);
and UO_460 (O_460,N_4424,N_3098);
or UO_461 (O_461,N_2754,N_3707);
nand UO_462 (O_462,N_4315,N_4834);
nand UO_463 (O_463,N_4220,N_4478);
nor UO_464 (O_464,N_4899,N_4102);
nor UO_465 (O_465,N_3063,N_3660);
or UO_466 (O_466,N_3416,N_2894);
nand UO_467 (O_467,N_4084,N_3117);
or UO_468 (O_468,N_2676,N_4789);
nand UO_469 (O_469,N_2607,N_3414);
or UO_470 (O_470,N_4108,N_4278);
or UO_471 (O_471,N_3744,N_4702);
nor UO_472 (O_472,N_3898,N_4747);
nand UO_473 (O_473,N_2875,N_4505);
and UO_474 (O_474,N_3026,N_4494);
and UO_475 (O_475,N_3060,N_4640);
nand UO_476 (O_476,N_2973,N_3854);
nand UO_477 (O_477,N_4161,N_3005);
xor UO_478 (O_478,N_3693,N_3480);
or UO_479 (O_479,N_4409,N_4760);
and UO_480 (O_480,N_3887,N_3914);
nor UO_481 (O_481,N_3208,N_4399);
xor UO_482 (O_482,N_3613,N_4889);
and UO_483 (O_483,N_2562,N_4584);
nand UO_484 (O_484,N_3692,N_4493);
or UO_485 (O_485,N_3625,N_3509);
and UO_486 (O_486,N_2896,N_4819);
nand UO_487 (O_487,N_4262,N_3056);
nor UO_488 (O_488,N_2693,N_4660);
nor UO_489 (O_489,N_2519,N_3691);
nor UO_490 (O_490,N_3790,N_4768);
nor UO_491 (O_491,N_3690,N_2511);
and UO_492 (O_492,N_3409,N_4447);
or UO_493 (O_493,N_4115,N_2793);
or UO_494 (O_494,N_2741,N_4222);
nand UO_495 (O_495,N_4294,N_4062);
or UO_496 (O_496,N_4020,N_4018);
nor UO_497 (O_497,N_4152,N_2865);
nor UO_498 (O_498,N_2918,N_4580);
nand UO_499 (O_499,N_2675,N_4917);
and UO_500 (O_500,N_3151,N_4928);
or UO_501 (O_501,N_4535,N_4242);
and UO_502 (O_502,N_3905,N_3205);
and UO_503 (O_503,N_2587,N_4027);
nand UO_504 (O_504,N_4470,N_3377);
nand UO_505 (O_505,N_2961,N_2836);
nor UO_506 (O_506,N_3289,N_3122);
nor UO_507 (O_507,N_3162,N_3374);
and UO_508 (O_508,N_3802,N_3185);
nor UO_509 (O_509,N_3817,N_4187);
nor UO_510 (O_510,N_4722,N_4524);
and UO_511 (O_511,N_4219,N_4351);
nand UO_512 (O_512,N_2619,N_3238);
or UO_513 (O_513,N_3612,N_4874);
xnor UO_514 (O_514,N_4564,N_3595);
and UO_515 (O_515,N_4547,N_3742);
nor UO_516 (O_516,N_2778,N_3921);
or UO_517 (O_517,N_3459,N_2557);
and UO_518 (O_518,N_3042,N_3448);
nand UO_519 (O_519,N_3792,N_3044);
and UO_520 (O_520,N_3773,N_4792);
nor UO_521 (O_521,N_4643,N_3814);
nand UO_522 (O_522,N_2766,N_4685);
nand UO_523 (O_523,N_4946,N_3300);
or UO_524 (O_524,N_4307,N_3090);
nand UO_525 (O_525,N_3057,N_4110);
nand UO_526 (O_526,N_4157,N_2586);
nor UO_527 (O_527,N_3230,N_3600);
nor UO_528 (O_528,N_3399,N_4474);
or UO_529 (O_529,N_2846,N_4360);
nand UO_530 (O_530,N_3784,N_4599);
nor UO_531 (O_531,N_4127,N_3530);
or UO_532 (O_532,N_4200,N_3002);
or UO_533 (O_533,N_4558,N_4128);
nand UO_534 (O_534,N_4011,N_3010);
and UO_535 (O_535,N_3137,N_4134);
or UO_536 (O_536,N_2810,N_3709);
nand UO_537 (O_537,N_3634,N_3382);
nand UO_538 (O_538,N_4395,N_3498);
nor UO_539 (O_539,N_3680,N_2787);
or UO_540 (O_540,N_4319,N_3527);
or UO_541 (O_541,N_4413,N_4082);
nor UO_542 (O_542,N_4510,N_3633);
nand UO_543 (O_543,N_3115,N_3223);
nor UO_544 (O_544,N_3065,N_4454);
or UO_545 (O_545,N_2702,N_2593);
nor UO_546 (O_546,N_4331,N_3909);
and UO_547 (O_547,N_3246,N_4559);
nand UO_548 (O_548,N_4009,N_4321);
or UO_549 (O_549,N_2510,N_3934);
nand UO_550 (O_550,N_4081,N_3471);
nor UO_551 (O_551,N_3857,N_3048);
nor UO_552 (O_552,N_4452,N_4811);
nand UO_553 (O_553,N_4754,N_2776);
or UO_554 (O_554,N_3568,N_3320);
or UO_555 (O_555,N_2818,N_3505);
and UO_556 (O_556,N_3713,N_2883);
nor UO_557 (O_557,N_3458,N_4896);
nor UO_558 (O_558,N_4386,N_2860);
or UO_559 (O_559,N_2669,N_4473);
and UO_560 (O_560,N_3269,N_4057);
nor UO_561 (O_561,N_3810,N_3621);
nand UO_562 (O_562,N_3194,N_3771);
or UO_563 (O_563,N_3000,N_4857);
and UO_564 (O_564,N_2939,N_4680);
or UO_565 (O_565,N_4445,N_4291);
nor UO_566 (O_566,N_3868,N_3228);
or UO_567 (O_567,N_4988,N_2755);
or UO_568 (O_568,N_4008,N_4397);
and UO_569 (O_569,N_4856,N_3943);
or UO_570 (O_570,N_3473,N_3695);
or UO_571 (O_571,N_3325,N_4723);
nand UO_572 (O_572,N_2945,N_3091);
nor UO_573 (O_573,N_4629,N_2515);
nor UO_574 (O_574,N_4696,N_4089);
and UO_575 (O_575,N_3799,N_2653);
or UO_576 (O_576,N_4402,N_4832);
nand UO_577 (O_577,N_3421,N_2753);
or UO_578 (O_578,N_4457,N_2532);
or UO_579 (O_579,N_3607,N_2618);
nor UO_580 (O_580,N_4221,N_4563);
or UO_581 (O_581,N_2691,N_2580);
nand UO_582 (O_582,N_3211,N_4804);
and UO_583 (O_583,N_4892,N_3545);
nand UO_584 (O_584,N_3991,N_2801);
or UO_585 (O_585,N_3348,N_4669);
nand UO_586 (O_586,N_3085,N_2904);
and UO_587 (O_587,N_3630,N_3047);
nand UO_588 (O_588,N_2800,N_3681);
and UO_589 (O_589,N_3175,N_3614);
or UO_590 (O_590,N_3375,N_3822);
nor UO_591 (O_591,N_2570,N_4544);
nand UO_592 (O_592,N_3646,N_4342);
and UO_593 (O_593,N_2848,N_4016);
and UO_594 (O_594,N_3965,N_2824);
or UO_595 (O_595,N_4963,N_4712);
and UO_596 (O_596,N_4610,N_4041);
nor UO_597 (O_597,N_3862,N_3476);
and UO_598 (O_598,N_3078,N_3092);
nand UO_599 (O_599,N_3697,N_2674);
or UO_600 (O_600,N_3931,N_2902);
nand UO_601 (O_601,N_4479,N_3800);
nor UO_602 (O_602,N_4566,N_3356);
nor UO_603 (O_603,N_4777,N_3040);
nand UO_604 (O_604,N_2687,N_4267);
and UO_605 (O_605,N_3866,N_3251);
or UO_606 (O_606,N_4339,N_4619);
nand UO_607 (O_607,N_3120,N_3376);
and UO_608 (O_608,N_3778,N_3587);
and UO_609 (O_609,N_2660,N_2815);
xor UO_610 (O_610,N_4244,N_2526);
or UO_611 (O_611,N_2777,N_4788);
nand UO_612 (O_612,N_3486,N_3615);
nand UO_613 (O_613,N_3926,N_3258);
or UO_614 (O_614,N_2987,N_2514);
and UO_615 (O_615,N_4340,N_3855);
and UO_616 (O_616,N_3945,N_2523);
nand UO_617 (O_617,N_3555,N_2879);
nand UO_618 (O_618,N_3373,N_3977);
and UO_619 (O_619,N_3155,N_2967);
nor UO_620 (O_620,N_3838,N_2791);
and UO_621 (O_621,N_2582,N_4953);
nand UO_622 (O_622,N_2701,N_3357);
nor UO_623 (O_623,N_3582,N_2849);
or UO_624 (O_624,N_3620,N_2834);
nand UO_625 (O_625,N_4612,N_3190);
nand UO_626 (O_626,N_3895,N_3084);
or UO_627 (O_627,N_2535,N_4406);
nand UO_628 (O_628,N_3759,N_3393);
and UO_629 (O_629,N_2527,N_3280);
or UO_630 (O_630,N_4498,N_2838);
nor UO_631 (O_631,N_4154,N_2655);
nor UO_632 (O_632,N_3765,N_3329);
and UO_633 (O_633,N_4308,N_2979);
and UO_634 (O_634,N_3665,N_3578);
and UO_635 (O_635,N_4298,N_3215);
or UO_636 (O_636,N_2652,N_2771);
nand UO_637 (O_637,N_4790,N_3468);
nand UO_638 (O_638,N_4188,N_4675);
or UO_639 (O_639,N_4233,N_4635);
or UO_640 (O_640,N_2821,N_4461);
nand UO_641 (O_641,N_2900,N_3849);
and UO_642 (O_642,N_3039,N_3837);
nor UO_643 (O_643,N_2898,N_3363);
nand UO_644 (O_644,N_3250,N_4240);
or UO_645 (O_645,N_4533,N_4545);
nor UO_646 (O_646,N_2749,N_4357);
or UO_647 (O_647,N_3551,N_2829);
nand UO_648 (O_648,N_4980,N_3694);
nor UO_649 (O_649,N_4440,N_4905);
and UO_650 (O_650,N_2703,N_4268);
nor UO_651 (O_651,N_4781,N_3082);
and UO_652 (O_652,N_4023,N_4509);
nor UO_653 (O_653,N_4029,N_2827);
and UO_654 (O_654,N_2819,N_4264);
xor UO_655 (O_655,N_3974,N_4209);
or UO_656 (O_656,N_3929,N_4667);
nor UO_657 (O_657,N_2881,N_3804);
nor UO_658 (O_658,N_3467,N_4875);
and UO_659 (O_659,N_4653,N_3499);
nand UO_660 (O_660,N_3278,N_4915);
nand UO_661 (O_661,N_4323,N_2585);
nand UO_662 (O_662,N_2913,N_3781);
or UO_663 (O_663,N_3571,N_3272);
nand UO_664 (O_664,N_3050,N_3727);
and UO_665 (O_665,N_4362,N_4387);
nand UO_666 (O_666,N_3858,N_3077);
and UO_667 (O_667,N_4815,N_3307);
nor UO_668 (O_668,N_3142,N_2512);
and UO_669 (O_669,N_3860,N_3454);
nor UO_670 (O_670,N_2839,N_2812);
nor UO_671 (O_671,N_4080,N_4528);
nand UO_672 (O_672,N_4328,N_2775);
and UO_673 (O_673,N_4939,N_3825);
and UO_674 (O_674,N_4539,N_3192);
nand UO_675 (O_675,N_4178,N_3508);
nor UO_676 (O_676,N_4822,N_2506);
nand UO_677 (O_677,N_2844,N_3751);
nor UO_678 (O_678,N_2715,N_4400);
nand UO_679 (O_679,N_3036,N_4486);
and UO_680 (O_680,N_2784,N_3266);
nand UO_681 (O_681,N_4255,N_4828);
or UO_682 (O_682,N_3463,N_3139);
and UO_683 (O_683,N_2899,N_2609);
nor UO_684 (O_684,N_3622,N_3664);
or UO_685 (O_685,N_4391,N_4578);
or UO_686 (O_686,N_4002,N_3339);
nor UO_687 (O_687,N_3644,N_3522);
and UO_688 (O_688,N_4311,N_3355);
nand UO_689 (O_689,N_3996,N_2628);
and UO_690 (O_690,N_3859,N_2591);
or UO_691 (O_691,N_3684,N_2978);
nand UO_692 (O_692,N_3741,N_3193);
and UO_693 (O_693,N_2907,N_4287);
nor UO_694 (O_694,N_4678,N_4191);
and UO_695 (O_695,N_2509,N_4557);
xnor UO_696 (O_696,N_3888,N_3105);
nor UO_697 (O_697,N_3418,N_4356);
nor UO_698 (O_698,N_2651,N_4469);
or UO_699 (O_699,N_3306,N_4797);
nor UO_700 (O_700,N_2940,N_3176);
or UO_701 (O_701,N_3071,N_4574);
and UO_702 (O_702,N_3712,N_3706);
and UO_703 (O_703,N_4941,N_3455);
nor UO_704 (O_704,N_3061,N_3293);
and UO_705 (O_705,N_2641,N_4179);
nor UO_706 (O_706,N_4019,N_3890);
nand UO_707 (O_707,N_4589,N_3366);
nor UO_708 (O_708,N_3893,N_4898);
nand UO_709 (O_709,N_4055,N_3332);
nor UO_710 (O_710,N_3705,N_4677);
xor UO_711 (O_711,N_3816,N_2761);
nand UO_712 (O_712,N_3097,N_3322);
nand UO_713 (O_713,N_2871,N_3820);
and UO_714 (O_714,N_3515,N_2572);
nand UO_715 (O_715,N_4885,N_3719);
nand UO_716 (O_716,N_4160,N_4761);
and UO_717 (O_717,N_3444,N_2789);
nand UO_718 (O_718,N_3733,N_3310);
and UO_719 (O_719,N_2733,N_4503);
nor UO_720 (O_720,N_3940,N_4679);
or UO_721 (O_721,N_2870,N_2541);
or UO_722 (O_722,N_2760,N_3412);
nor UO_723 (O_723,N_2942,N_4596);
and UO_724 (O_724,N_4123,N_4234);
and UO_725 (O_725,N_4849,N_2520);
nand UO_726 (O_726,N_3317,N_3274);
nand UO_727 (O_727,N_4130,N_3668);
nand UO_728 (O_728,N_3132,N_3563);
nand UO_729 (O_729,N_4700,N_2536);
and UO_730 (O_730,N_3389,N_2930);
or UO_731 (O_731,N_3562,N_4906);
or UO_732 (O_732,N_3852,N_4404);
nor UO_733 (O_733,N_4017,N_4237);
or UO_734 (O_734,N_4662,N_3842);
nand UO_735 (O_735,N_3081,N_3532);
and UO_736 (O_736,N_3290,N_2507);
nor UO_737 (O_737,N_3806,N_3714);
or UO_738 (O_738,N_3432,N_4870);
nand UO_739 (O_739,N_3725,N_2956);
nor UO_740 (O_740,N_3227,N_4638);
nand UO_741 (O_741,N_3805,N_3461);
or UO_742 (O_742,N_2897,N_3196);
nor UO_743 (O_743,N_3602,N_3558);
or UO_744 (O_744,N_2635,N_3303);
and UO_745 (O_745,N_3338,N_4631);
and UO_746 (O_746,N_4131,N_3066);
or UO_747 (O_747,N_4784,N_3878);
or UO_748 (O_748,N_4350,N_3839);
or UO_749 (O_749,N_3403,N_3153);
or UO_750 (O_750,N_4607,N_4852);
nand UO_751 (O_751,N_4618,N_4713);
and UO_752 (O_752,N_4169,N_4961);
nand UO_753 (O_753,N_4289,N_4256);
nand UO_754 (O_754,N_3465,N_4997);
and UO_755 (O_755,N_2630,N_2508);
nor UO_756 (O_756,N_2743,N_4448);
and UO_757 (O_757,N_3256,N_3856);
or UO_758 (O_758,N_4958,N_4728);
nor UO_759 (O_759,N_4513,N_3201);
and UO_760 (O_760,N_3986,N_2721);
or UO_761 (O_761,N_3894,N_4966);
nand UO_762 (O_762,N_2626,N_4868);
and UO_763 (O_763,N_3014,N_2617);
nand UO_764 (O_764,N_3743,N_3884);
nor UO_765 (O_765,N_3286,N_2764);
and UO_766 (O_766,N_3203,N_4079);
and UO_767 (O_767,N_3579,N_4259);
or UO_768 (O_768,N_2935,N_3877);
and UO_769 (O_769,N_3942,N_4846);
nor UO_770 (O_770,N_2748,N_4796);
nor UO_771 (O_771,N_4228,N_2735);
nor UO_772 (O_772,N_2991,N_4050);
and UO_773 (O_773,N_2648,N_2982);
nand UO_774 (O_774,N_3074,N_2658);
or UO_775 (O_775,N_4762,N_4534);
nor UO_776 (O_776,N_2959,N_4197);
and UO_777 (O_777,N_4734,N_4717);
and UO_778 (O_778,N_3433,N_4542);
and UO_779 (O_779,N_4116,N_3672);
and UO_780 (O_780,N_2874,N_3850);
nor UO_781 (O_781,N_3446,N_2785);
nor UO_782 (O_782,N_2944,N_3426);
nand UO_783 (O_783,N_4038,N_3259);
nand UO_784 (O_784,N_3335,N_4463);
nand UO_785 (O_785,N_3346,N_3876);
nand UO_786 (O_786,N_3234,N_3439);
or UO_787 (O_787,N_2692,N_4814);
nor UO_788 (O_788,N_4245,N_2524);
nor UO_789 (O_789,N_4972,N_3411);
and UO_790 (O_790,N_2690,N_4411);
or UO_791 (O_791,N_3449,N_4305);
or UO_792 (O_792,N_2529,N_4393);
nor UO_793 (O_793,N_3950,N_2831);
nor UO_794 (O_794,N_3763,N_3941);
nor UO_795 (O_795,N_3581,N_3282);
or UO_796 (O_796,N_3526,N_3507);
nand UO_797 (O_797,N_4987,N_3012);
nor UO_798 (O_798,N_2558,N_2673);
or UO_799 (O_799,N_3220,N_2661);
and UO_800 (O_800,N_4073,N_4232);
nand UO_801 (O_801,N_4218,N_4951);
nor UO_802 (O_802,N_2720,N_4136);
and UO_803 (O_803,N_3072,N_2869);
nor UO_804 (O_804,N_3540,N_2559);
or UO_805 (O_805,N_4622,N_2695);
nand UO_806 (O_806,N_4306,N_3013);
nand UO_807 (O_807,N_4907,N_4138);
or UO_808 (O_808,N_3488,N_3813);
and UO_809 (O_809,N_2947,N_2759);
and UO_810 (O_810,N_2921,N_4652);
and UO_811 (O_811,N_4067,N_3301);
nand UO_812 (O_812,N_3383,N_3429);
and UO_813 (O_813,N_4581,N_3536);
nand UO_814 (O_814,N_4076,N_4475);
and UO_815 (O_815,N_3538,N_4993);
and UO_816 (O_816,N_3311,N_4850);
nor UO_817 (O_817,N_4432,N_3632);
or UO_818 (O_818,N_4973,N_4337);
or UO_819 (O_819,N_3038,N_3391);
and UO_820 (O_820,N_3549,N_4608);
and UO_821 (O_821,N_3650,N_4069);
and UO_822 (O_822,N_4113,N_3254);
nand UO_823 (O_823,N_2640,N_3933);
nor UO_824 (O_824,N_4210,N_3992);
nand UO_825 (O_825,N_2763,N_4467);
nor UO_826 (O_826,N_4913,N_4415);
nand UO_827 (O_827,N_4022,N_2781);
nor UO_828 (O_828,N_2806,N_3466);
nand UO_829 (O_829,N_4368,N_3495);
nand UO_830 (O_830,N_4265,N_4694);
nor UO_831 (O_831,N_4004,N_3009);
nor UO_832 (O_832,N_4829,N_3396);
or UO_833 (O_833,N_4600,N_4933);
nor UO_834 (O_834,N_3474,N_2990);
or UO_835 (O_835,N_3715,N_4854);
nand UO_836 (O_836,N_4030,N_4661);
or UO_837 (O_837,N_4674,N_3772);
nor UO_838 (O_838,N_2707,N_3724);
nand UO_839 (O_839,N_3157,N_4934);
xor UO_840 (O_840,N_4686,N_4992);
nor UO_841 (O_841,N_4139,N_3094);
and UO_842 (O_842,N_3209,N_4884);
and UO_843 (O_843,N_4403,N_4174);
nor UO_844 (O_844,N_3670,N_3603);
nor UO_845 (O_845,N_3631,N_3271);
or UO_846 (O_846,N_3035,N_4773);
and UO_847 (O_847,N_3179,N_4367);
xor UO_848 (O_848,N_3520,N_2595);
and UO_849 (O_849,N_3248,N_2688);
nor UO_850 (O_850,N_3350,N_2983);
and UO_851 (O_851,N_4450,N_4170);
and UO_852 (O_852,N_3675,N_3019);
nand UO_853 (O_853,N_3628,N_3031);
and UO_854 (O_854,N_3494,N_4873);
nand UO_855 (O_855,N_4621,N_3114);
nand UO_856 (O_856,N_3756,N_4532);
nand UO_857 (O_857,N_3360,N_4756);
nand UO_858 (O_858,N_3611,N_4683);
or UO_859 (O_859,N_3517,N_2912);
nand UO_860 (O_860,N_4199,N_4763);
nor UO_861 (O_861,N_3239,N_4538);
and UO_862 (O_862,N_4844,N_3542);
nor UO_863 (O_863,N_3653,N_3368);
nand UO_864 (O_864,N_4959,N_2600);
or UO_865 (O_865,N_4750,N_3276);
and UO_866 (O_866,N_2995,N_3605);
or UO_867 (O_867,N_4014,N_2708);
or UO_868 (O_868,N_4689,N_3982);
and UO_869 (O_869,N_2711,N_2584);
or UO_870 (O_870,N_3342,N_4358);
and UO_871 (O_871,N_3586,N_4780);
nor UO_872 (O_872,N_3919,N_2989);
nand UO_873 (O_873,N_4926,N_3601);
nand UO_874 (O_874,N_2622,N_3669);
nand UO_875 (O_875,N_4078,N_2625);
xor UO_876 (O_876,N_3167,N_3326);
or UO_877 (O_877,N_3277,N_4204);
nand UO_878 (O_878,N_4100,N_4937);
nor UO_879 (O_879,N_4246,N_3087);
nor UO_880 (O_880,N_4481,N_3103);
nand UO_881 (O_881,N_2788,N_3626);
nand UO_882 (O_882,N_2599,N_4842);
or UO_883 (O_883,N_3457,N_4431);
and UO_884 (O_884,N_3288,N_3762);
or UO_885 (O_885,N_4625,N_2841);
nand UO_886 (O_886,N_2556,N_4107);
nor UO_887 (O_887,N_4177,N_3604);
or UO_888 (O_888,N_3550,N_4732);
or UO_889 (O_889,N_3511,N_2730);
nand UO_890 (O_890,N_3386,N_2571);
nand UO_891 (O_891,N_2837,N_4276);
and UO_892 (O_892,N_4361,N_4275);
nor UO_893 (O_893,N_4903,N_2858);
nand UO_894 (O_894,N_2943,N_2644);
nor UO_895 (O_895,N_4285,N_4185);
and UO_896 (O_896,N_3510,N_2905);
or UO_897 (O_897,N_2561,N_3336);
or UO_898 (O_898,N_2780,N_2813);
nor UO_899 (O_899,N_3291,N_3128);
nor UO_900 (O_900,N_2773,N_4206);
nand UO_901 (O_901,N_2699,N_4141);
nor UO_902 (O_902,N_4560,N_3750);
xor UO_903 (O_903,N_3902,N_4736);
nand UO_904 (O_904,N_4392,N_3999);
and UO_905 (O_905,N_2993,N_4417);
nand UO_906 (O_906,N_3676,N_4248);
nor UO_907 (O_907,N_4979,N_4634);
and UO_908 (O_908,N_2765,N_2974);
nor UO_909 (O_909,N_4927,N_3273);
or UO_910 (O_910,N_4365,N_3369);
xor UO_911 (O_911,N_4540,N_3118);
nor UO_912 (O_912,N_2823,N_3845);
nand UO_913 (O_913,N_2530,N_2716);
or UO_914 (O_914,N_2543,N_2620);
nand UO_915 (O_915,N_4583,N_4145);
nor UO_916 (O_916,N_4338,N_2548);
nor UO_917 (O_917,N_4202,N_4518);
nor UO_918 (O_918,N_3119,N_3637);
nor UO_919 (O_919,N_2884,N_4826);
nor UO_920 (O_920,N_3801,N_2627);
nor UO_921 (O_921,N_4620,N_3367);
nor UO_922 (O_922,N_3647,N_2615);
nand UO_923 (O_923,N_4181,N_3823);
nand UO_924 (O_924,N_4000,N_4942);
nor UO_925 (O_925,N_3299,N_3163);
nand UO_926 (O_926,N_3865,N_4708);
or UO_927 (O_927,N_4423,N_3219);
nand UO_928 (O_928,N_4587,N_2564);
nand UO_929 (O_929,N_3569,N_3717);
nor UO_930 (O_930,N_3927,N_4721);
nand UO_931 (O_931,N_2576,N_4155);
or UO_932 (O_932,N_4658,N_2925);
nor UO_933 (O_933,N_4147,N_4785);
nand UO_934 (O_934,N_3313,N_4866);
and UO_935 (O_935,N_3195,N_4462);
nor UO_936 (O_936,N_4290,N_3958);
and UO_937 (O_937,N_4886,N_3577);
nor UO_938 (O_938,N_4541,N_3584);
nor UO_939 (O_939,N_2914,N_3575);
nor UO_940 (O_940,N_2908,N_3337);
nor UO_941 (O_941,N_3099,N_4977);
or UO_942 (O_942,N_4047,N_2531);
xnor UO_943 (O_943,N_4830,N_4303);
nand UO_944 (O_944,N_4861,N_2868);
nand UO_945 (O_945,N_4364,N_2949);
or UO_946 (O_946,N_4986,N_4772);
nor UO_947 (O_947,N_2933,N_3708);
nand UO_948 (O_948,N_2603,N_3124);
nor UO_949 (O_949,N_4567,N_2700);
or UO_950 (O_950,N_4504,N_3478);
and UO_951 (O_951,N_4837,N_3100);
and UO_952 (O_952,N_3841,N_2888);
and UO_953 (O_953,N_3679,N_4468);
or UO_954 (O_954,N_2608,N_4825);
and UO_955 (O_955,N_2680,N_2951);
and UO_956 (O_956,N_3226,N_4681);
nand UO_957 (O_957,N_2889,N_3779);
nand UO_958 (O_958,N_3353,N_4381);
nand UO_959 (O_959,N_4624,N_3101);
nor UO_960 (O_960,N_3798,N_4015);
or UO_961 (O_961,N_4999,N_2862);
nand UO_962 (O_962,N_3032,N_4664);
or UO_963 (O_963,N_4348,N_2610);
and UO_964 (O_964,N_3126,N_3951);
and UO_965 (O_965,N_4598,N_3487);
and UO_966 (O_966,N_3746,N_3828);
and UO_967 (O_967,N_3889,N_2909);
nor UO_968 (O_968,N_3966,N_3410);
or UO_969 (O_969,N_4487,N_4523);
nor UO_970 (O_970,N_3704,N_3407);
and UO_971 (O_971,N_3450,N_3782);
or UO_972 (O_972,N_3512,N_2521);
nor UO_973 (O_973,N_2747,N_4793);
or UO_974 (O_974,N_4778,N_4330);
or UO_975 (O_975,N_3218,N_4143);
or UO_976 (O_976,N_2980,N_2732);
or UO_977 (O_977,N_3830,N_3443);
nand UO_978 (O_978,N_4373,N_3152);
nand UO_979 (O_979,N_4312,N_3440);
nand UO_980 (O_980,N_2605,N_4623);
and UO_981 (O_981,N_3774,N_4098);
nand UO_982 (O_982,N_4164,N_4235);
nor UO_983 (O_983,N_3976,N_3159);
nand UO_984 (O_984,N_2805,N_4695);
and UO_985 (O_985,N_4707,N_4230);
nor UO_986 (O_986,N_4758,N_4613);
or UO_987 (O_987,N_4398,N_3312);
nand UO_988 (O_988,N_4525,N_3460);
nor UO_989 (O_989,N_4672,N_4996);
nor UO_990 (O_990,N_4586,N_2734);
and UO_991 (O_991,N_4688,N_4902);
nand UO_992 (O_992,N_3583,N_3832);
nor UO_993 (O_993,N_4394,N_4687);
or UO_994 (O_994,N_3904,N_3541);
nand UO_995 (O_995,N_4426,N_3182);
and UO_996 (O_996,N_4887,N_4153);
nand UO_997 (O_997,N_3420,N_3267);
nor UO_998 (O_998,N_3930,N_2503);
and UO_999 (O_999,N_4072,N_3918);
endmodule