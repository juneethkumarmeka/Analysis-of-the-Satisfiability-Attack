module basic_500_3000_500_40_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_295,In_287);
and U1 (N_1,In_312,In_294);
nand U2 (N_2,In_37,In_259);
nor U3 (N_3,In_416,In_176);
and U4 (N_4,In_471,In_379);
or U5 (N_5,In_173,In_372);
or U6 (N_6,In_154,In_207);
nand U7 (N_7,In_419,In_165);
nor U8 (N_8,In_410,In_357);
and U9 (N_9,In_111,In_297);
nor U10 (N_10,In_202,In_393);
and U11 (N_11,In_182,In_333);
nand U12 (N_12,In_387,In_134);
nand U13 (N_13,In_274,In_57);
nand U14 (N_14,In_221,In_69);
or U15 (N_15,In_195,In_412);
and U16 (N_16,In_121,In_28);
or U17 (N_17,In_230,In_449);
xnor U18 (N_18,In_417,In_13);
nand U19 (N_19,In_81,In_286);
nand U20 (N_20,In_169,In_143);
nand U21 (N_21,In_115,In_124);
nor U22 (N_22,In_461,In_348);
or U23 (N_23,In_367,In_443);
and U24 (N_24,In_237,In_76);
and U25 (N_25,In_30,In_2);
and U26 (N_26,In_240,In_214);
or U27 (N_27,In_481,In_332);
xor U28 (N_28,In_229,In_170);
nand U29 (N_29,In_324,In_263);
nor U30 (N_30,In_23,In_252);
or U31 (N_31,In_268,In_160);
nand U32 (N_32,In_14,In_90);
nand U33 (N_33,In_460,In_109);
xnor U34 (N_34,In_466,In_371);
or U35 (N_35,In_474,In_453);
or U36 (N_36,In_288,In_95);
or U37 (N_37,In_212,In_465);
or U38 (N_38,In_411,In_210);
and U39 (N_39,In_125,In_38);
nand U40 (N_40,In_52,In_83);
and U41 (N_41,In_456,In_484);
and U42 (N_42,In_437,In_187);
and U43 (N_43,In_175,In_459);
and U44 (N_44,In_440,In_236);
or U45 (N_45,In_36,In_382);
nand U46 (N_46,In_6,In_421);
and U47 (N_47,In_424,In_255);
nand U48 (N_48,In_241,In_475);
or U49 (N_49,In_362,In_491);
nor U50 (N_50,In_395,In_157);
nand U51 (N_51,In_46,In_188);
or U52 (N_52,In_281,In_155);
or U53 (N_53,In_470,In_423);
nand U54 (N_54,In_266,In_29);
nand U55 (N_55,In_129,In_303);
xor U56 (N_56,In_84,In_360);
and U57 (N_57,In_467,In_445);
nor U58 (N_58,In_388,In_359);
nor U59 (N_59,In_334,In_189);
nor U60 (N_60,In_211,In_427);
nand U61 (N_61,In_326,In_4);
or U62 (N_62,In_67,In_140);
or U63 (N_63,In_486,In_374);
or U64 (N_64,In_101,In_163);
or U65 (N_65,In_253,In_448);
nand U66 (N_66,In_112,In_350);
nand U67 (N_67,In_289,In_321);
xor U68 (N_68,In_161,In_493);
and U69 (N_69,In_331,In_78);
nand U70 (N_70,In_123,In_432);
or U71 (N_71,In_58,In_298);
or U72 (N_72,In_43,In_64);
and U73 (N_73,In_264,In_299);
nor U74 (N_74,In_70,In_269);
or U75 (N_75,In_267,In_63);
nor U76 (N_76,In_490,In_329);
nand U77 (N_77,In_290,In_420);
nand U78 (N_78,In_180,N_33);
and U79 (N_79,In_479,N_29);
and U80 (N_80,In_291,In_194);
nand U81 (N_81,In_311,In_378);
or U82 (N_82,In_409,In_216);
or U83 (N_83,In_150,In_179);
and U84 (N_84,In_5,In_248);
nand U85 (N_85,In_80,In_270);
or U86 (N_86,In_239,In_60);
or U87 (N_87,In_283,In_201);
nand U88 (N_88,In_363,In_122);
nand U89 (N_89,In_137,In_231);
xnor U90 (N_90,N_68,N_71);
and U91 (N_91,In_234,In_462);
nand U92 (N_92,In_177,In_10);
xnor U93 (N_93,In_65,In_158);
nor U94 (N_94,N_35,In_454);
and U95 (N_95,N_57,In_463);
nand U96 (N_96,In_31,N_10);
nor U97 (N_97,In_394,N_74);
nor U98 (N_98,In_322,In_349);
and U99 (N_99,In_213,In_108);
nor U100 (N_100,In_261,In_296);
and U101 (N_101,In_429,In_314);
or U102 (N_102,In_309,In_389);
nor U103 (N_103,N_39,In_1);
and U104 (N_104,In_426,In_205);
and U105 (N_105,In_337,In_209);
nand U106 (N_106,In_247,N_30);
nand U107 (N_107,In_144,In_439);
nand U108 (N_108,In_342,In_345);
or U109 (N_109,In_330,N_12);
or U110 (N_110,In_398,In_167);
nor U111 (N_111,In_232,In_319);
nor U112 (N_112,In_141,In_116);
or U113 (N_113,In_190,In_438);
nor U114 (N_114,In_271,N_47);
or U115 (N_115,N_53,In_442);
nor U116 (N_116,In_383,In_22);
nand U117 (N_117,In_185,In_219);
nand U118 (N_118,N_32,In_495);
nand U119 (N_119,In_223,N_7);
or U120 (N_120,N_21,In_128);
or U121 (N_121,N_14,In_56);
nand U122 (N_122,In_73,In_482);
nor U123 (N_123,N_24,In_301);
or U124 (N_124,In_92,In_145);
nand U125 (N_125,In_27,In_18);
nor U126 (N_126,In_477,In_338);
nand U127 (N_127,In_184,In_104);
or U128 (N_128,In_405,N_27);
nor U129 (N_129,In_20,In_469);
xor U130 (N_130,In_156,In_9);
nand U131 (N_131,In_352,N_61);
or U132 (N_132,In_181,In_215);
nor U133 (N_133,In_135,In_132);
nand U134 (N_134,N_52,N_5);
nand U135 (N_135,In_71,N_58);
and U136 (N_136,In_318,In_226);
nor U137 (N_137,In_48,N_73);
nand U138 (N_138,In_39,In_256);
or U139 (N_139,In_340,In_91);
and U140 (N_140,In_12,In_483);
and U141 (N_141,In_55,In_280);
xor U142 (N_142,In_66,N_1);
or U143 (N_143,In_341,In_87);
and U144 (N_144,In_159,In_40);
nor U145 (N_145,In_191,In_59);
nand U146 (N_146,In_168,In_316);
nor U147 (N_147,In_17,In_183);
or U148 (N_148,In_244,N_55);
nor U149 (N_149,In_285,In_323);
or U150 (N_150,In_220,N_23);
nor U151 (N_151,In_361,In_164);
or U152 (N_152,In_254,In_381);
nand U153 (N_153,N_99,In_431);
nor U154 (N_154,N_128,N_104);
nand U155 (N_155,In_130,N_63);
and U156 (N_156,N_31,In_196);
nor U157 (N_157,N_40,In_139);
or U158 (N_158,N_4,N_93);
nor U159 (N_159,N_94,In_276);
nor U160 (N_160,N_34,N_116);
or U161 (N_161,N_50,In_284);
nand U162 (N_162,In_396,N_42);
xnor U163 (N_163,In_488,In_89);
or U164 (N_164,In_310,N_119);
nand U165 (N_165,In_217,N_108);
nor U166 (N_166,In_273,In_119);
or U167 (N_167,N_111,In_250);
xor U168 (N_168,N_28,N_103);
and U169 (N_169,N_101,In_433);
nand U170 (N_170,In_278,In_305);
nor U171 (N_171,In_428,In_402);
nor U172 (N_172,N_113,In_408);
nor U173 (N_173,N_66,N_90);
nand U174 (N_174,In_246,N_8);
nor U175 (N_175,N_132,In_0);
and U176 (N_176,In_45,In_390);
and U177 (N_177,In_114,In_368);
nor U178 (N_178,N_88,N_114);
and U179 (N_179,In_293,In_222);
nor U180 (N_180,In_110,In_472);
and U181 (N_181,In_494,In_85);
nor U182 (N_182,In_47,N_60);
nor U183 (N_183,N_124,In_399);
and U184 (N_184,In_464,N_125);
nor U185 (N_185,N_91,N_146);
nor U186 (N_186,N_107,In_489);
or U187 (N_187,In_384,In_444);
nand U188 (N_188,In_162,In_243);
nor U189 (N_189,In_172,In_192);
and U190 (N_190,In_304,In_203);
and U191 (N_191,N_56,In_492);
xnor U192 (N_192,N_105,In_136);
nand U193 (N_193,In_3,N_3);
and U194 (N_194,In_458,In_335);
nor U195 (N_195,In_391,N_83);
nand U196 (N_196,In_88,N_77);
nor U197 (N_197,In_369,In_166);
nand U198 (N_198,In_468,In_44);
nand U199 (N_199,In_320,N_129);
or U200 (N_200,In_497,In_118);
or U201 (N_201,N_38,In_74);
nor U202 (N_202,N_45,In_450);
nand U203 (N_203,N_95,N_82);
or U204 (N_204,In_249,In_282);
or U205 (N_205,N_51,In_251);
and U206 (N_206,N_96,N_138);
nand U207 (N_207,In_265,In_366);
and U208 (N_208,N_70,N_123);
or U209 (N_209,In_356,N_121);
nand U210 (N_210,In_86,In_328);
nand U211 (N_211,N_41,In_49);
nand U212 (N_212,In_430,N_134);
nor U213 (N_213,N_122,N_118);
or U214 (N_214,In_364,In_93);
and U215 (N_215,N_43,In_127);
and U216 (N_216,In_106,In_392);
and U217 (N_217,In_292,In_53);
nor U218 (N_218,In_422,In_401);
nor U219 (N_219,In_197,In_242);
and U220 (N_220,In_50,N_17);
xnor U221 (N_221,N_0,In_302);
or U222 (N_222,In_94,N_75);
nand U223 (N_223,In_376,In_26);
and U224 (N_224,N_25,N_11);
nand U225 (N_225,In_151,In_346);
nor U226 (N_226,N_19,In_407);
nand U227 (N_227,N_136,In_414);
nand U228 (N_228,N_157,N_141);
nor U229 (N_229,In_224,In_72);
nor U230 (N_230,N_191,In_377);
xnor U231 (N_231,N_178,N_176);
and U232 (N_232,N_184,In_206);
nor U233 (N_233,In_275,In_133);
nand U234 (N_234,In_355,In_33);
nand U235 (N_235,N_115,In_262);
and U236 (N_236,N_120,N_211);
and U237 (N_237,N_203,In_307);
or U238 (N_238,In_434,N_148);
nand U239 (N_239,N_160,In_7);
nor U240 (N_240,In_96,In_446);
nor U241 (N_241,In_113,In_476);
nand U242 (N_242,In_228,N_2);
nand U243 (N_243,N_150,In_403);
nand U244 (N_244,N_181,In_308);
nand U245 (N_245,N_85,N_216);
or U246 (N_246,N_201,N_152);
nor U247 (N_247,N_164,In_98);
nor U248 (N_248,N_18,N_190);
and U249 (N_249,In_198,In_441);
or U250 (N_250,In_339,N_109);
nor U251 (N_251,N_54,In_385);
nor U252 (N_252,N_218,In_277);
nor U253 (N_253,N_126,In_99);
and U254 (N_254,In_358,In_257);
nand U255 (N_255,In_32,N_210);
and U256 (N_256,In_400,In_62);
and U257 (N_257,In_258,In_436);
nand U258 (N_258,N_221,In_153);
or U259 (N_259,N_194,In_24);
or U260 (N_260,In_418,In_452);
nor U261 (N_261,N_199,N_102);
nand U262 (N_262,N_222,N_220);
nand U263 (N_263,In_34,N_166);
or U264 (N_264,N_198,N_168);
nor U265 (N_265,N_97,In_82);
nand U266 (N_266,In_131,N_172);
nand U267 (N_267,N_207,In_487);
nand U268 (N_268,In_315,N_202);
nor U269 (N_269,In_300,N_145);
and U270 (N_270,N_155,In_375);
and U271 (N_271,N_209,N_147);
or U272 (N_272,N_140,N_100);
or U273 (N_273,In_42,In_54);
xnor U274 (N_274,In_107,In_415);
and U275 (N_275,N_44,N_144);
or U276 (N_276,N_185,N_162);
and U277 (N_277,In_404,In_306);
or U278 (N_278,In_138,N_133);
and U279 (N_279,In_41,N_177);
or U280 (N_280,N_112,N_98);
nor U281 (N_281,In_142,In_455);
or U282 (N_282,N_86,N_213);
or U283 (N_283,In_435,In_327);
and U284 (N_284,In_100,In_105);
nand U285 (N_285,N_180,N_174);
and U286 (N_286,N_153,In_457);
nand U287 (N_287,In_146,N_79);
nor U288 (N_288,N_81,N_224);
and U289 (N_289,In_480,In_238);
and U290 (N_290,N_76,In_227);
nand U291 (N_291,N_219,In_152);
nand U292 (N_292,In_102,N_131);
and U293 (N_293,N_13,In_171);
or U294 (N_294,N_158,In_21);
or U295 (N_295,N_204,In_225);
and U296 (N_296,N_188,N_106);
nor U297 (N_297,N_197,In_25);
or U298 (N_298,N_16,N_9);
nor U299 (N_299,N_59,N_159);
xor U300 (N_300,N_156,N_231);
nor U301 (N_301,In_499,N_187);
nor U302 (N_302,N_244,In_336);
nand U303 (N_303,N_291,N_151);
nand U304 (N_304,N_215,N_277);
or U305 (N_305,N_279,N_135);
nor U306 (N_306,N_171,In_148);
or U307 (N_307,N_232,N_253);
or U308 (N_308,In_260,In_11);
or U309 (N_309,N_127,N_92);
nor U310 (N_310,N_286,N_293);
nand U311 (N_311,N_230,N_284);
nor U312 (N_312,N_87,In_77);
and U313 (N_313,In_235,N_26);
nor U314 (N_314,N_46,In_478);
and U315 (N_315,N_254,N_161);
or U316 (N_316,N_243,N_72);
nor U317 (N_317,N_281,In_199);
nand U318 (N_318,N_233,N_239);
nand U319 (N_319,In_373,N_283);
or U320 (N_320,N_261,In_473);
or U321 (N_321,In_354,N_130);
nor U322 (N_322,N_214,N_186);
and U323 (N_323,In_380,N_274);
nand U324 (N_324,In_406,N_6);
or U325 (N_325,In_204,N_217);
nor U326 (N_326,N_289,In_233);
or U327 (N_327,In_68,N_205);
nor U328 (N_328,N_250,N_49);
nor U329 (N_329,N_169,N_117);
nor U330 (N_330,N_295,In_313);
and U331 (N_331,In_353,In_126);
or U332 (N_332,In_317,In_193);
and U333 (N_333,N_228,N_266);
nor U334 (N_334,N_139,In_103);
nor U335 (N_335,N_287,N_69);
nand U336 (N_336,In_149,N_292);
nor U337 (N_337,N_267,N_206);
nor U338 (N_338,N_299,N_225);
and U339 (N_339,In_498,N_285);
nor U340 (N_340,In_75,N_154);
nor U341 (N_341,N_275,N_62);
or U342 (N_342,N_110,N_170);
nor U343 (N_343,N_276,In_120);
or U344 (N_344,In_325,N_20);
or U345 (N_345,N_238,In_343);
nor U346 (N_346,N_227,N_260);
and U347 (N_347,N_258,N_280);
nand U348 (N_348,N_269,In_15);
nor U349 (N_349,N_234,In_178);
or U350 (N_350,N_296,N_149);
nand U351 (N_351,In_200,In_35);
or U352 (N_352,N_80,In_344);
nor U353 (N_353,N_268,N_65);
nor U354 (N_354,N_189,N_240);
or U355 (N_355,N_226,In_272);
nor U356 (N_356,N_137,In_16);
or U357 (N_357,N_278,N_183);
and U358 (N_358,N_248,In_218);
nand U359 (N_359,N_223,N_173);
nor U360 (N_360,N_245,N_237);
nor U361 (N_361,N_142,N_273);
nor U362 (N_362,N_256,In_485);
or U363 (N_363,N_282,N_271);
or U364 (N_364,N_78,In_496);
and U365 (N_365,N_288,In_351);
nand U366 (N_366,N_64,N_67);
and U367 (N_367,In_147,N_182);
and U368 (N_368,N_163,N_249);
or U369 (N_369,N_264,In_425);
nand U370 (N_370,In_451,N_48);
nand U371 (N_371,N_270,N_175);
nand U372 (N_372,N_242,N_265);
nand U373 (N_373,N_252,N_37);
or U374 (N_374,N_22,In_413);
or U375 (N_375,N_312,N_336);
nor U376 (N_376,N_355,N_322);
nand U377 (N_377,N_262,N_309);
or U378 (N_378,In_117,N_324);
or U379 (N_379,N_360,N_308);
or U380 (N_380,N_251,N_300);
nand U381 (N_381,N_357,N_236);
or U382 (N_382,In_365,N_167);
and U383 (N_383,N_347,N_359);
or U384 (N_384,N_349,In_447);
or U385 (N_385,In_208,N_319);
nand U386 (N_386,N_212,N_374);
or U387 (N_387,In_370,N_15);
nand U388 (N_388,N_193,In_397);
and U389 (N_389,N_330,N_165);
or U390 (N_390,N_290,N_338);
or U391 (N_391,N_302,In_386);
and U392 (N_392,N_326,N_297);
and U393 (N_393,N_361,N_365);
nor U394 (N_394,N_329,N_341);
nor U395 (N_395,N_257,N_255);
or U396 (N_396,In_347,In_245);
nand U397 (N_397,N_318,N_366);
nand U398 (N_398,N_334,N_323);
nor U399 (N_399,N_303,N_315);
and U400 (N_400,N_235,N_320);
nand U401 (N_401,N_246,N_84);
and U402 (N_402,N_304,N_310);
nand U403 (N_403,N_372,In_8);
and U404 (N_404,N_305,N_200);
nor U405 (N_405,N_208,N_332);
or U406 (N_406,N_307,N_298);
or U407 (N_407,N_354,N_351);
nand U408 (N_408,N_143,In_97);
or U409 (N_409,N_346,N_317);
nand U410 (N_410,N_350,In_51);
and U411 (N_411,N_352,N_314);
nor U412 (N_412,N_339,In_79);
nand U413 (N_413,N_321,N_333);
nor U414 (N_414,N_356,In_19);
or U415 (N_415,N_345,N_313);
or U416 (N_416,N_353,N_358);
xnor U417 (N_417,N_367,N_363);
or U418 (N_418,N_259,N_311);
or U419 (N_419,N_368,In_61);
nand U420 (N_420,In_186,N_371);
nor U421 (N_421,N_196,N_331);
nand U422 (N_422,N_369,In_174);
or U423 (N_423,N_335,N_272);
nor U424 (N_424,N_192,N_179);
nand U425 (N_425,N_343,N_89);
nand U426 (N_426,N_337,N_327);
nor U427 (N_427,N_247,N_229);
nor U428 (N_428,N_325,N_348);
and U429 (N_429,N_195,N_306);
and U430 (N_430,N_373,N_316);
nand U431 (N_431,N_241,N_294);
nand U432 (N_432,N_344,N_263);
xnor U433 (N_433,N_342,N_340);
nand U434 (N_434,N_328,N_364);
nor U435 (N_435,N_36,N_301);
nand U436 (N_436,In_279,N_370);
nand U437 (N_437,N_362,N_310);
nor U438 (N_438,N_297,N_307);
nor U439 (N_439,N_328,N_340);
nand U440 (N_440,N_318,N_247);
and U441 (N_441,N_322,N_304);
or U442 (N_442,In_97,In_347);
nand U443 (N_443,N_337,N_314);
and U444 (N_444,N_36,In_370);
nor U445 (N_445,In_61,N_364);
xor U446 (N_446,In_365,N_372);
nor U447 (N_447,N_200,N_368);
or U448 (N_448,In_347,N_336);
or U449 (N_449,N_196,N_315);
or U450 (N_450,N_410,N_415);
xnor U451 (N_451,N_411,N_413);
and U452 (N_452,N_377,N_408);
nor U453 (N_453,N_414,N_425);
nor U454 (N_454,N_435,N_383);
or U455 (N_455,N_449,N_402);
or U456 (N_456,N_444,N_380);
nand U457 (N_457,N_416,N_427);
nor U458 (N_458,N_433,N_422);
and U459 (N_459,N_421,N_379);
and U460 (N_460,N_385,N_438);
nor U461 (N_461,N_403,N_404);
xnor U462 (N_462,N_389,N_406);
nand U463 (N_463,N_442,N_405);
or U464 (N_464,N_401,N_390);
and U465 (N_465,N_446,N_376);
or U466 (N_466,N_439,N_440);
or U467 (N_467,N_429,N_428);
nor U468 (N_468,N_418,N_382);
or U469 (N_469,N_447,N_436);
nand U470 (N_470,N_419,N_395);
and U471 (N_471,N_420,N_394);
and U472 (N_472,N_384,N_397);
or U473 (N_473,N_443,N_375);
or U474 (N_474,N_426,N_391);
or U475 (N_475,N_398,N_392);
nor U476 (N_476,N_431,N_399);
nand U477 (N_477,N_412,N_430);
nor U478 (N_478,N_445,N_407);
and U479 (N_479,N_396,N_434);
nand U480 (N_480,N_378,N_400);
nand U481 (N_481,N_437,N_387);
nand U482 (N_482,N_441,N_424);
xnor U483 (N_483,N_423,N_448);
and U484 (N_484,N_417,N_432);
nand U485 (N_485,N_386,N_381);
and U486 (N_486,N_388,N_409);
nand U487 (N_487,N_393,N_386);
nand U488 (N_488,N_413,N_401);
or U489 (N_489,N_443,N_382);
nand U490 (N_490,N_418,N_429);
nand U491 (N_491,N_432,N_399);
or U492 (N_492,N_433,N_447);
nand U493 (N_493,N_413,N_435);
or U494 (N_494,N_396,N_403);
and U495 (N_495,N_412,N_380);
or U496 (N_496,N_439,N_412);
nand U497 (N_497,N_397,N_417);
nand U498 (N_498,N_409,N_439);
or U499 (N_499,N_431,N_388);
and U500 (N_500,N_379,N_436);
or U501 (N_501,N_440,N_407);
nor U502 (N_502,N_448,N_407);
or U503 (N_503,N_440,N_385);
or U504 (N_504,N_430,N_415);
nor U505 (N_505,N_399,N_430);
xor U506 (N_506,N_425,N_447);
xnor U507 (N_507,N_382,N_427);
nand U508 (N_508,N_381,N_407);
and U509 (N_509,N_429,N_401);
nand U510 (N_510,N_410,N_407);
xor U511 (N_511,N_401,N_381);
nand U512 (N_512,N_428,N_389);
or U513 (N_513,N_445,N_406);
nand U514 (N_514,N_423,N_443);
nor U515 (N_515,N_424,N_429);
nand U516 (N_516,N_384,N_399);
nor U517 (N_517,N_442,N_416);
or U518 (N_518,N_403,N_375);
nand U519 (N_519,N_383,N_444);
and U520 (N_520,N_375,N_412);
nor U521 (N_521,N_426,N_433);
nor U522 (N_522,N_432,N_430);
nand U523 (N_523,N_387,N_426);
nand U524 (N_524,N_375,N_389);
and U525 (N_525,N_488,N_493);
and U526 (N_526,N_455,N_498);
nand U527 (N_527,N_505,N_462);
nor U528 (N_528,N_466,N_510);
or U529 (N_529,N_506,N_456);
and U530 (N_530,N_523,N_521);
or U531 (N_531,N_509,N_503);
or U532 (N_532,N_458,N_501);
and U533 (N_533,N_467,N_491);
nor U534 (N_534,N_481,N_522);
nand U535 (N_535,N_460,N_475);
nand U536 (N_536,N_504,N_469);
and U537 (N_537,N_495,N_459);
nand U538 (N_538,N_507,N_518);
nor U539 (N_539,N_517,N_490);
nand U540 (N_540,N_451,N_489);
nand U541 (N_541,N_453,N_486);
or U542 (N_542,N_482,N_480);
nand U543 (N_543,N_472,N_502);
and U544 (N_544,N_476,N_524);
or U545 (N_545,N_464,N_471);
nor U546 (N_546,N_511,N_477);
and U547 (N_547,N_492,N_499);
nor U548 (N_548,N_483,N_463);
and U549 (N_549,N_500,N_494);
or U550 (N_550,N_457,N_461);
or U551 (N_551,N_470,N_452);
nor U552 (N_552,N_468,N_478);
or U553 (N_553,N_520,N_514);
nand U554 (N_554,N_513,N_512);
xor U555 (N_555,N_465,N_496);
and U556 (N_556,N_508,N_473);
and U557 (N_557,N_485,N_484);
nand U558 (N_558,N_450,N_479);
nor U559 (N_559,N_515,N_474);
and U560 (N_560,N_516,N_487);
or U561 (N_561,N_519,N_454);
or U562 (N_562,N_497,N_478);
or U563 (N_563,N_492,N_474);
nand U564 (N_564,N_450,N_460);
and U565 (N_565,N_459,N_481);
and U566 (N_566,N_491,N_501);
nor U567 (N_567,N_454,N_474);
nor U568 (N_568,N_486,N_491);
or U569 (N_569,N_513,N_463);
xnor U570 (N_570,N_473,N_459);
nand U571 (N_571,N_457,N_489);
or U572 (N_572,N_496,N_524);
and U573 (N_573,N_474,N_499);
or U574 (N_574,N_461,N_501);
nand U575 (N_575,N_484,N_461);
nor U576 (N_576,N_505,N_484);
and U577 (N_577,N_450,N_469);
and U578 (N_578,N_476,N_458);
nand U579 (N_579,N_502,N_487);
xor U580 (N_580,N_495,N_468);
or U581 (N_581,N_493,N_501);
nand U582 (N_582,N_479,N_497);
nor U583 (N_583,N_496,N_485);
and U584 (N_584,N_461,N_465);
or U585 (N_585,N_498,N_481);
or U586 (N_586,N_483,N_482);
nand U587 (N_587,N_505,N_501);
nand U588 (N_588,N_500,N_471);
or U589 (N_589,N_501,N_468);
nand U590 (N_590,N_461,N_488);
nand U591 (N_591,N_463,N_494);
or U592 (N_592,N_502,N_457);
nand U593 (N_593,N_490,N_483);
nand U594 (N_594,N_472,N_509);
or U595 (N_595,N_486,N_520);
nor U596 (N_596,N_472,N_505);
or U597 (N_597,N_507,N_500);
nand U598 (N_598,N_470,N_477);
or U599 (N_599,N_506,N_477);
or U600 (N_600,N_587,N_563);
nor U601 (N_601,N_577,N_539);
xor U602 (N_602,N_544,N_529);
nand U603 (N_603,N_556,N_575);
nand U604 (N_604,N_551,N_595);
or U605 (N_605,N_565,N_537);
nor U606 (N_606,N_567,N_553);
or U607 (N_607,N_591,N_588);
nand U608 (N_608,N_571,N_592);
nor U609 (N_609,N_530,N_576);
nand U610 (N_610,N_543,N_582);
and U611 (N_611,N_550,N_573);
nor U612 (N_612,N_578,N_585);
and U613 (N_613,N_542,N_546);
nand U614 (N_614,N_527,N_540);
nand U615 (N_615,N_581,N_526);
and U616 (N_616,N_594,N_549);
nand U617 (N_617,N_552,N_593);
nor U618 (N_618,N_548,N_538);
nor U619 (N_619,N_584,N_547);
nand U620 (N_620,N_590,N_545);
xor U621 (N_621,N_589,N_560);
or U622 (N_622,N_558,N_536);
nand U623 (N_623,N_554,N_533);
nand U624 (N_624,N_568,N_535);
or U625 (N_625,N_574,N_599);
nor U626 (N_626,N_531,N_597);
and U627 (N_627,N_541,N_569);
nand U628 (N_628,N_534,N_598);
and U629 (N_629,N_562,N_532);
or U630 (N_630,N_528,N_559);
and U631 (N_631,N_570,N_561);
nand U632 (N_632,N_566,N_572);
xor U633 (N_633,N_555,N_557);
nand U634 (N_634,N_583,N_564);
nand U635 (N_635,N_596,N_579);
nand U636 (N_636,N_586,N_580);
nor U637 (N_637,N_525,N_588);
nand U638 (N_638,N_534,N_593);
nand U639 (N_639,N_537,N_541);
or U640 (N_640,N_557,N_587);
nor U641 (N_641,N_570,N_528);
nand U642 (N_642,N_569,N_563);
and U643 (N_643,N_593,N_543);
and U644 (N_644,N_566,N_569);
nor U645 (N_645,N_528,N_599);
and U646 (N_646,N_576,N_525);
and U647 (N_647,N_531,N_569);
or U648 (N_648,N_566,N_585);
nor U649 (N_649,N_565,N_550);
nand U650 (N_650,N_586,N_560);
or U651 (N_651,N_573,N_535);
and U652 (N_652,N_582,N_564);
or U653 (N_653,N_568,N_596);
nor U654 (N_654,N_578,N_543);
nor U655 (N_655,N_571,N_542);
nor U656 (N_656,N_568,N_575);
nand U657 (N_657,N_530,N_546);
nand U658 (N_658,N_545,N_599);
nand U659 (N_659,N_586,N_554);
nand U660 (N_660,N_534,N_527);
or U661 (N_661,N_577,N_537);
nor U662 (N_662,N_531,N_549);
or U663 (N_663,N_536,N_544);
or U664 (N_664,N_599,N_596);
and U665 (N_665,N_590,N_555);
or U666 (N_666,N_525,N_578);
and U667 (N_667,N_563,N_527);
and U668 (N_668,N_582,N_578);
or U669 (N_669,N_583,N_532);
or U670 (N_670,N_533,N_562);
nor U671 (N_671,N_539,N_569);
and U672 (N_672,N_588,N_526);
nor U673 (N_673,N_530,N_560);
nand U674 (N_674,N_538,N_592);
nor U675 (N_675,N_617,N_636);
nor U676 (N_676,N_632,N_660);
or U677 (N_677,N_645,N_608);
or U678 (N_678,N_664,N_606);
nor U679 (N_679,N_613,N_641);
and U680 (N_680,N_662,N_647);
or U681 (N_681,N_670,N_671);
nand U682 (N_682,N_656,N_667);
nand U683 (N_683,N_614,N_669);
or U684 (N_684,N_639,N_674);
nand U685 (N_685,N_643,N_607);
nor U686 (N_686,N_666,N_651);
nor U687 (N_687,N_620,N_626);
nor U688 (N_688,N_630,N_629);
nand U689 (N_689,N_631,N_658);
nor U690 (N_690,N_638,N_673);
nand U691 (N_691,N_657,N_648);
or U692 (N_692,N_603,N_655);
nand U693 (N_693,N_640,N_637);
and U694 (N_694,N_646,N_622);
and U695 (N_695,N_623,N_625);
or U696 (N_696,N_659,N_612);
nor U697 (N_697,N_628,N_609);
and U698 (N_698,N_634,N_615);
nand U699 (N_699,N_672,N_668);
nor U700 (N_700,N_600,N_616);
and U701 (N_701,N_663,N_635);
or U702 (N_702,N_633,N_644);
nand U703 (N_703,N_619,N_654);
nand U704 (N_704,N_642,N_661);
nor U705 (N_705,N_653,N_605);
and U706 (N_706,N_602,N_610);
xnor U707 (N_707,N_611,N_650);
or U708 (N_708,N_618,N_624);
or U709 (N_709,N_652,N_649);
nand U710 (N_710,N_621,N_627);
and U711 (N_711,N_665,N_601);
nor U712 (N_712,N_604,N_638);
and U713 (N_713,N_625,N_609);
xnor U714 (N_714,N_605,N_622);
and U715 (N_715,N_668,N_618);
nand U716 (N_716,N_674,N_621);
or U717 (N_717,N_654,N_635);
nand U718 (N_718,N_619,N_660);
and U719 (N_719,N_656,N_663);
or U720 (N_720,N_617,N_646);
nor U721 (N_721,N_656,N_657);
xnor U722 (N_722,N_629,N_647);
nor U723 (N_723,N_660,N_641);
and U724 (N_724,N_670,N_609);
or U725 (N_725,N_608,N_662);
and U726 (N_726,N_627,N_659);
or U727 (N_727,N_667,N_605);
nor U728 (N_728,N_663,N_671);
or U729 (N_729,N_616,N_632);
nand U730 (N_730,N_634,N_613);
nand U731 (N_731,N_612,N_625);
or U732 (N_732,N_674,N_640);
nand U733 (N_733,N_651,N_624);
or U734 (N_734,N_613,N_600);
and U735 (N_735,N_664,N_624);
nand U736 (N_736,N_657,N_605);
nor U737 (N_737,N_641,N_621);
or U738 (N_738,N_607,N_604);
nand U739 (N_739,N_629,N_610);
nor U740 (N_740,N_668,N_669);
nor U741 (N_741,N_627,N_644);
nor U742 (N_742,N_652,N_634);
and U743 (N_743,N_624,N_655);
or U744 (N_744,N_607,N_628);
nor U745 (N_745,N_618,N_663);
nand U746 (N_746,N_663,N_674);
and U747 (N_747,N_659,N_625);
and U748 (N_748,N_647,N_656);
or U749 (N_749,N_612,N_636);
nor U750 (N_750,N_714,N_723);
nand U751 (N_751,N_737,N_748);
and U752 (N_752,N_729,N_733);
nor U753 (N_753,N_706,N_704);
nand U754 (N_754,N_745,N_701);
or U755 (N_755,N_718,N_710);
nand U756 (N_756,N_722,N_719);
nand U757 (N_757,N_711,N_739);
and U758 (N_758,N_698,N_728);
and U759 (N_759,N_712,N_708);
and U760 (N_760,N_736,N_717);
nor U761 (N_761,N_691,N_676);
nor U762 (N_762,N_743,N_678);
and U763 (N_763,N_705,N_740);
nor U764 (N_764,N_734,N_699);
nor U765 (N_765,N_731,N_697);
or U766 (N_766,N_707,N_689);
or U767 (N_767,N_680,N_686);
or U768 (N_768,N_742,N_735);
nor U769 (N_769,N_713,N_747);
or U770 (N_770,N_725,N_693);
nand U771 (N_771,N_692,N_715);
nor U772 (N_772,N_685,N_681);
nand U773 (N_773,N_675,N_696);
and U774 (N_774,N_732,N_684);
nor U775 (N_775,N_703,N_716);
nand U776 (N_776,N_702,N_727);
nand U777 (N_777,N_721,N_688);
and U778 (N_778,N_730,N_694);
or U779 (N_779,N_683,N_687);
nand U780 (N_780,N_700,N_746);
and U781 (N_781,N_677,N_679);
or U782 (N_782,N_682,N_738);
or U783 (N_783,N_726,N_749);
nor U784 (N_784,N_709,N_744);
and U785 (N_785,N_741,N_695);
or U786 (N_786,N_690,N_724);
nor U787 (N_787,N_720,N_749);
nor U788 (N_788,N_694,N_698);
nor U789 (N_789,N_675,N_727);
or U790 (N_790,N_686,N_717);
and U791 (N_791,N_749,N_692);
or U792 (N_792,N_686,N_745);
and U793 (N_793,N_712,N_699);
nand U794 (N_794,N_718,N_713);
or U795 (N_795,N_679,N_706);
xor U796 (N_796,N_744,N_716);
and U797 (N_797,N_694,N_696);
nand U798 (N_798,N_704,N_689);
and U799 (N_799,N_738,N_681);
and U800 (N_800,N_717,N_730);
xnor U801 (N_801,N_746,N_748);
nor U802 (N_802,N_749,N_736);
and U803 (N_803,N_705,N_707);
and U804 (N_804,N_714,N_677);
nor U805 (N_805,N_691,N_717);
nor U806 (N_806,N_742,N_699);
or U807 (N_807,N_726,N_738);
or U808 (N_808,N_700,N_686);
nand U809 (N_809,N_688,N_701);
nand U810 (N_810,N_694,N_739);
nor U811 (N_811,N_737,N_718);
or U812 (N_812,N_725,N_681);
or U813 (N_813,N_711,N_696);
nand U814 (N_814,N_727,N_701);
nand U815 (N_815,N_695,N_711);
and U816 (N_816,N_681,N_732);
xor U817 (N_817,N_747,N_742);
or U818 (N_818,N_727,N_706);
nand U819 (N_819,N_698,N_696);
or U820 (N_820,N_680,N_739);
nor U821 (N_821,N_681,N_704);
and U822 (N_822,N_704,N_680);
or U823 (N_823,N_689,N_725);
nand U824 (N_824,N_728,N_713);
nand U825 (N_825,N_761,N_811);
and U826 (N_826,N_784,N_777);
or U827 (N_827,N_787,N_806);
nand U828 (N_828,N_756,N_819);
nor U829 (N_829,N_758,N_753);
nand U830 (N_830,N_780,N_762);
or U831 (N_831,N_786,N_814);
nand U832 (N_832,N_801,N_817);
or U833 (N_833,N_822,N_769);
and U834 (N_834,N_773,N_754);
nor U835 (N_835,N_775,N_752);
nor U836 (N_836,N_813,N_824);
or U837 (N_837,N_750,N_792);
and U838 (N_838,N_794,N_767);
and U839 (N_839,N_798,N_788);
nand U840 (N_840,N_793,N_797);
and U841 (N_841,N_763,N_796);
and U842 (N_842,N_765,N_810);
nor U843 (N_843,N_781,N_812);
and U844 (N_844,N_772,N_778);
and U845 (N_845,N_755,N_803);
nor U846 (N_846,N_776,N_809);
and U847 (N_847,N_808,N_759);
and U848 (N_848,N_764,N_823);
or U849 (N_849,N_779,N_783);
nand U850 (N_850,N_768,N_795);
and U851 (N_851,N_751,N_805);
xor U852 (N_852,N_790,N_820);
or U853 (N_853,N_804,N_807);
nand U854 (N_854,N_766,N_821);
nor U855 (N_855,N_799,N_770);
nand U856 (N_856,N_815,N_785);
nor U857 (N_857,N_800,N_774);
and U858 (N_858,N_757,N_816);
or U859 (N_859,N_789,N_802);
and U860 (N_860,N_771,N_818);
nand U861 (N_861,N_760,N_791);
nor U862 (N_862,N_782,N_822);
nor U863 (N_863,N_802,N_787);
nor U864 (N_864,N_763,N_791);
nand U865 (N_865,N_790,N_791);
nand U866 (N_866,N_821,N_787);
or U867 (N_867,N_771,N_820);
nand U868 (N_868,N_766,N_803);
or U869 (N_869,N_814,N_824);
nor U870 (N_870,N_782,N_802);
nor U871 (N_871,N_790,N_754);
nor U872 (N_872,N_770,N_764);
nor U873 (N_873,N_808,N_819);
nand U874 (N_874,N_754,N_770);
nand U875 (N_875,N_786,N_790);
and U876 (N_876,N_797,N_778);
nand U877 (N_877,N_813,N_820);
nand U878 (N_878,N_805,N_786);
or U879 (N_879,N_763,N_780);
or U880 (N_880,N_786,N_788);
nor U881 (N_881,N_793,N_779);
or U882 (N_882,N_793,N_788);
nand U883 (N_883,N_766,N_761);
or U884 (N_884,N_757,N_787);
nor U885 (N_885,N_788,N_796);
xor U886 (N_886,N_759,N_779);
nor U887 (N_887,N_774,N_786);
nor U888 (N_888,N_799,N_796);
nor U889 (N_889,N_788,N_813);
nand U890 (N_890,N_750,N_798);
nor U891 (N_891,N_789,N_824);
or U892 (N_892,N_791,N_821);
nand U893 (N_893,N_753,N_800);
nand U894 (N_894,N_795,N_762);
or U895 (N_895,N_767,N_780);
nor U896 (N_896,N_767,N_788);
and U897 (N_897,N_822,N_779);
and U898 (N_898,N_780,N_795);
nand U899 (N_899,N_774,N_803);
and U900 (N_900,N_864,N_867);
nor U901 (N_901,N_862,N_875);
nor U902 (N_902,N_831,N_891);
nor U903 (N_903,N_827,N_829);
and U904 (N_904,N_868,N_839);
and U905 (N_905,N_884,N_834);
nand U906 (N_906,N_832,N_855);
nor U907 (N_907,N_880,N_860);
nand U908 (N_908,N_887,N_836);
and U909 (N_909,N_879,N_876);
and U910 (N_910,N_894,N_872);
nor U911 (N_911,N_886,N_892);
and U912 (N_912,N_874,N_859);
nor U913 (N_913,N_853,N_895);
or U914 (N_914,N_888,N_845);
xnor U915 (N_915,N_835,N_897);
or U916 (N_916,N_838,N_896);
or U917 (N_917,N_847,N_883);
nand U918 (N_918,N_863,N_885);
nor U919 (N_919,N_846,N_851);
nand U920 (N_920,N_843,N_828);
nand U921 (N_921,N_850,N_890);
and U922 (N_922,N_837,N_854);
xnor U923 (N_923,N_830,N_871);
nor U924 (N_924,N_840,N_866);
or U925 (N_925,N_865,N_825);
nand U926 (N_926,N_898,N_878);
or U927 (N_927,N_852,N_833);
nor U928 (N_928,N_881,N_882);
and U929 (N_929,N_841,N_893);
and U930 (N_930,N_889,N_856);
nand U931 (N_931,N_869,N_848);
and U932 (N_932,N_826,N_844);
nor U933 (N_933,N_873,N_861);
and U934 (N_934,N_849,N_842);
nand U935 (N_935,N_877,N_858);
and U936 (N_936,N_857,N_899);
or U937 (N_937,N_870,N_845);
or U938 (N_938,N_867,N_869);
and U939 (N_939,N_863,N_890);
or U940 (N_940,N_832,N_882);
nand U941 (N_941,N_868,N_838);
or U942 (N_942,N_852,N_848);
and U943 (N_943,N_892,N_851);
nor U944 (N_944,N_845,N_892);
or U945 (N_945,N_839,N_878);
and U946 (N_946,N_851,N_860);
nor U947 (N_947,N_862,N_837);
nor U948 (N_948,N_896,N_849);
or U949 (N_949,N_896,N_825);
or U950 (N_950,N_881,N_876);
or U951 (N_951,N_837,N_899);
nand U952 (N_952,N_828,N_854);
nor U953 (N_953,N_862,N_849);
and U954 (N_954,N_864,N_876);
or U955 (N_955,N_863,N_861);
nand U956 (N_956,N_840,N_880);
nor U957 (N_957,N_833,N_884);
nor U958 (N_958,N_826,N_890);
or U959 (N_959,N_858,N_872);
nor U960 (N_960,N_876,N_861);
xnor U961 (N_961,N_825,N_826);
nand U962 (N_962,N_843,N_881);
and U963 (N_963,N_894,N_826);
nor U964 (N_964,N_884,N_847);
nor U965 (N_965,N_869,N_887);
nor U966 (N_966,N_872,N_862);
nor U967 (N_967,N_862,N_826);
and U968 (N_968,N_833,N_885);
nand U969 (N_969,N_895,N_828);
or U970 (N_970,N_873,N_892);
and U971 (N_971,N_845,N_829);
or U972 (N_972,N_855,N_867);
nor U973 (N_973,N_842,N_834);
and U974 (N_974,N_825,N_891);
nand U975 (N_975,N_970,N_957);
and U976 (N_976,N_947,N_919);
nand U977 (N_977,N_930,N_940);
or U978 (N_978,N_964,N_914);
nor U979 (N_979,N_922,N_963);
or U980 (N_980,N_945,N_959);
xor U981 (N_981,N_933,N_909);
xor U982 (N_982,N_906,N_960);
nand U983 (N_983,N_951,N_902);
and U984 (N_984,N_961,N_962);
nor U985 (N_985,N_915,N_937);
nor U986 (N_986,N_953,N_916);
nand U987 (N_987,N_969,N_912);
nand U988 (N_988,N_955,N_966);
and U989 (N_989,N_967,N_904);
and U990 (N_990,N_905,N_903);
and U991 (N_991,N_913,N_934);
nor U992 (N_992,N_941,N_927);
or U993 (N_993,N_974,N_932);
nand U994 (N_994,N_965,N_971);
nand U995 (N_995,N_925,N_952);
nor U996 (N_996,N_924,N_936);
nor U997 (N_997,N_918,N_901);
or U998 (N_998,N_910,N_931);
and U999 (N_999,N_929,N_943);
nor U1000 (N_1000,N_946,N_911);
and U1001 (N_1001,N_948,N_949);
nand U1002 (N_1002,N_921,N_907);
or U1003 (N_1003,N_917,N_908);
xnor U1004 (N_1004,N_950,N_920);
and U1005 (N_1005,N_923,N_968);
nor U1006 (N_1006,N_942,N_928);
or U1007 (N_1007,N_972,N_956);
xnor U1008 (N_1008,N_900,N_958);
and U1009 (N_1009,N_926,N_935);
or U1010 (N_1010,N_954,N_938);
nor U1011 (N_1011,N_973,N_944);
and U1012 (N_1012,N_939,N_926);
or U1013 (N_1013,N_965,N_943);
nand U1014 (N_1014,N_955,N_959);
nor U1015 (N_1015,N_956,N_911);
nor U1016 (N_1016,N_919,N_911);
nor U1017 (N_1017,N_926,N_916);
nand U1018 (N_1018,N_920,N_960);
nor U1019 (N_1019,N_926,N_930);
and U1020 (N_1020,N_931,N_940);
nand U1021 (N_1021,N_938,N_969);
or U1022 (N_1022,N_950,N_953);
nor U1023 (N_1023,N_948,N_964);
and U1024 (N_1024,N_933,N_924);
nor U1025 (N_1025,N_950,N_931);
or U1026 (N_1026,N_914,N_900);
nor U1027 (N_1027,N_922,N_947);
and U1028 (N_1028,N_969,N_974);
and U1029 (N_1029,N_941,N_935);
and U1030 (N_1030,N_919,N_961);
xnor U1031 (N_1031,N_948,N_918);
nand U1032 (N_1032,N_920,N_917);
and U1033 (N_1033,N_902,N_936);
nand U1034 (N_1034,N_934,N_955);
nand U1035 (N_1035,N_969,N_945);
nand U1036 (N_1036,N_956,N_918);
or U1037 (N_1037,N_940,N_966);
nor U1038 (N_1038,N_900,N_970);
nor U1039 (N_1039,N_933,N_915);
nand U1040 (N_1040,N_970,N_961);
or U1041 (N_1041,N_934,N_911);
or U1042 (N_1042,N_941,N_947);
and U1043 (N_1043,N_961,N_959);
nor U1044 (N_1044,N_915,N_935);
nor U1045 (N_1045,N_908,N_900);
nand U1046 (N_1046,N_937,N_911);
or U1047 (N_1047,N_941,N_923);
nand U1048 (N_1048,N_945,N_901);
and U1049 (N_1049,N_936,N_919);
nor U1050 (N_1050,N_1029,N_1046);
or U1051 (N_1051,N_1049,N_1011);
nand U1052 (N_1052,N_1004,N_988);
xor U1053 (N_1053,N_1028,N_1014);
and U1054 (N_1054,N_1015,N_1007);
or U1055 (N_1055,N_1017,N_1025);
nor U1056 (N_1056,N_1006,N_1020);
nor U1057 (N_1057,N_976,N_992);
xor U1058 (N_1058,N_989,N_1018);
nor U1059 (N_1059,N_1002,N_1047);
nor U1060 (N_1060,N_1034,N_981);
or U1061 (N_1061,N_1032,N_1023);
or U1062 (N_1062,N_1043,N_1042);
or U1063 (N_1063,N_1030,N_1039);
nor U1064 (N_1064,N_1048,N_993);
nor U1065 (N_1065,N_996,N_975);
and U1066 (N_1066,N_1009,N_1013);
xor U1067 (N_1067,N_1012,N_978);
nor U1068 (N_1068,N_995,N_1005);
and U1069 (N_1069,N_1019,N_1037);
nand U1070 (N_1070,N_1038,N_982);
or U1071 (N_1071,N_984,N_1001);
or U1072 (N_1072,N_990,N_1008);
or U1073 (N_1073,N_983,N_1036);
and U1074 (N_1074,N_1040,N_1027);
nand U1075 (N_1075,N_979,N_1035);
and U1076 (N_1076,N_998,N_1024);
or U1077 (N_1077,N_980,N_1003);
nand U1078 (N_1078,N_1033,N_997);
or U1079 (N_1079,N_986,N_1016);
xor U1080 (N_1080,N_1010,N_1021);
or U1081 (N_1081,N_1026,N_1044);
nor U1082 (N_1082,N_1000,N_1041);
and U1083 (N_1083,N_999,N_991);
or U1084 (N_1084,N_1031,N_994);
and U1085 (N_1085,N_985,N_1045);
nor U1086 (N_1086,N_1022,N_987);
or U1087 (N_1087,N_977,N_1037);
xnor U1088 (N_1088,N_1021,N_1046);
and U1089 (N_1089,N_995,N_997);
or U1090 (N_1090,N_1044,N_1024);
xor U1091 (N_1091,N_988,N_1005);
nor U1092 (N_1092,N_1002,N_1003);
or U1093 (N_1093,N_990,N_981);
nor U1094 (N_1094,N_1032,N_1041);
nor U1095 (N_1095,N_977,N_1014);
nand U1096 (N_1096,N_1031,N_975);
and U1097 (N_1097,N_1027,N_1002);
xnor U1098 (N_1098,N_983,N_1012);
or U1099 (N_1099,N_1042,N_1021);
or U1100 (N_1100,N_1040,N_980);
nand U1101 (N_1101,N_981,N_984);
nand U1102 (N_1102,N_1010,N_1014);
nand U1103 (N_1103,N_1014,N_1024);
nand U1104 (N_1104,N_1030,N_1003);
or U1105 (N_1105,N_1039,N_1044);
nand U1106 (N_1106,N_1014,N_995);
or U1107 (N_1107,N_1022,N_1041);
or U1108 (N_1108,N_978,N_1007);
nor U1109 (N_1109,N_1021,N_1018);
and U1110 (N_1110,N_1025,N_1044);
or U1111 (N_1111,N_1005,N_1014);
xnor U1112 (N_1112,N_992,N_1035);
nor U1113 (N_1113,N_1041,N_1024);
nor U1114 (N_1114,N_990,N_991);
or U1115 (N_1115,N_1026,N_1015);
xnor U1116 (N_1116,N_1003,N_1012);
and U1117 (N_1117,N_985,N_992);
nor U1118 (N_1118,N_998,N_1010);
or U1119 (N_1119,N_1043,N_998);
or U1120 (N_1120,N_1021,N_987);
and U1121 (N_1121,N_1002,N_1026);
and U1122 (N_1122,N_1044,N_1040);
nor U1123 (N_1123,N_979,N_1011);
or U1124 (N_1124,N_1032,N_1006);
nor U1125 (N_1125,N_1087,N_1108);
nand U1126 (N_1126,N_1066,N_1069);
or U1127 (N_1127,N_1089,N_1085);
and U1128 (N_1128,N_1075,N_1095);
nor U1129 (N_1129,N_1058,N_1064);
or U1130 (N_1130,N_1073,N_1118);
and U1131 (N_1131,N_1055,N_1067);
nor U1132 (N_1132,N_1114,N_1115);
nand U1133 (N_1133,N_1119,N_1077);
and U1134 (N_1134,N_1112,N_1051);
and U1135 (N_1135,N_1120,N_1083);
nor U1136 (N_1136,N_1123,N_1063);
nand U1137 (N_1137,N_1098,N_1052);
nand U1138 (N_1138,N_1097,N_1101);
nand U1139 (N_1139,N_1068,N_1104);
nand U1140 (N_1140,N_1050,N_1122);
and U1141 (N_1141,N_1099,N_1081);
and U1142 (N_1142,N_1111,N_1116);
and U1143 (N_1143,N_1088,N_1092);
and U1144 (N_1144,N_1090,N_1102);
and U1145 (N_1145,N_1076,N_1121);
or U1146 (N_1146,N_1072,N_1057);
nor U1147 (N_1147,N_1074,N_1059);
or U1148 (N_1148,N_1106,N_1086);
nor U1149 (N_1149,N_1105,N_1103);
nand U1150 (N_1150,N_1096,N_1113);
or U1151 (N_1151,N_1056,N_1110);
nor U1152 (N_1152,N_1093,N_1062);
nor U1153 (N_1153,N_1070,N_1094);
nand U1154 (N_1154,N_1078,N_1065);
or U1155 (N_1155,N_1079,N_1084);
and U1156 (N_1156,N_1100,N_1107);
and U1157 (N_1157,N_1053,N_1080);
or U1158 (N_1158,N_1091,N_1109);
nor U1159 (N_1159,N_1117,N_1060);
nand U1160 (N_1160,N_1082,N_1054);
nand U1161 (N_1161,N_1071,N_1061);
nand U1162 (N_1162,N_1124,N_1094);
nor U1163 (N_1163,N_1057,N_1087);
and U1164 (N_1164,N_1058,N_1123);
or U1165 (N_1165,N_1088,N_1073);
or U1166 (N_1166,N_1073,N_1087);
nand U1167 (N_1167,N_1092,N_1081);
or U1168 (N_1168,N_1059,N_1116);
nand U1169 (N_1169,N_1058,N_1051);
nand U1170 (N_1170,N_1088,N_1114);
or U1171 (N_1171,N_1093,N_1104);
nor U1172 (N_1172,N_1061,N_1103);
nand U1173 (N_1173,N_1061,N_1055);
and U1174 (N_1174,N_1057,N_1058);
and U1175 (N_1175,N_1123,N_1089);
nor U1176 (N_1176,N_1103,N_1114);
and U1177 (N_1177,N_1092,N_1058);
or U1178 (N_1178,N_1052,N_1103);
or U1179 (N_1179,N_1087,N_1094);
and U1180 (N_1180,N_1077,N_1115);
nand U1181 (N_1181,N_1113,N_1120);
and U1182 (N_1182,N_1056,N_1118);
or U1183 (N_1183,N_1074,N_1123);
and U1184 (N_1184,N_1071,N_1091);
or U1185 (N_1185,N_1116,N_1054);
nand U1186 (N_1186,N_1088,N_1122);
or U1187 (N_1187,N_1061,N_1064);
and U1188 (N_1188,N_1060,N_1070);
and U1189 (N_1189,N_1080,N_1091);
nand U1190 (N_1190,N_1110,N_1092);
nand U1191 (N_1191,N_1075,N_1112);
nand U1192 (N_1192,N_1059,N_1062);
nand U1193 (N_1193,N_1082,N_1115);
or U1194 (N_1194,N_1082,N_1065);
nor U1195 (N_1195,N_1114,N_1084);
nand U1196 (N_1196,N_1051,N_1113);
nor U1197 (N_1197,N_1073,N_1084);
nor U1198 (N_1198,N_1095,N_1115);
nand U1199 (N_1199,N_1062,N_1097);
and U1200 (N_1200,N_1159,N_1185);
nor U1201 (N_1201,N_1157,N_1143);
nand U1202 (N_1202,N_1171,N_1130);
nand U1203 (N_1203,N_1132,N_1139);
and U1204 (N_1204,N_1191,N_1178);
or U1205 (N_1205,N_1195,N_1198);
nor U1206 (N_1206,N_1166,N_1151);
nand U1207 (N_1207,N_1158,N_1127);
nand U1208 (N_1208,N_1125,N_1141);
or U1209 (N_1209,N_1172,N_1148);
or U1210 (N_1210,N_1164,N_1169);
or U1211 (N_1211,N_1135,N_1156);
nand U1212 (N_1212,N_1155,N_1197);
nand U1213 (N_1213,N_1182,N_1176);
nor U1214 (N_1214,N_1140,N_1150);
or U1215 (N_1215,N_1180,N_1190);
and U1216 (N_1216,N_1173,N_1136);
nor U1217 (N_1217,N_1179,N_1153);
and U1218 (N_1218,N_1162,N_1154);
and U1219 (N_1219,N_1152,N_1144);
nand U1220 (N_1220,N_1128,N_1187);
and U1221 (N_1221,N_1170,N_1192);
or U1222 (N_1222,N_1138,N_1160);
nor U1223 (N_1223,N_1134,N_1161);
nor U1224 (N_1224,N_1163,N_1194);
and U1225 (N_1225,N_1193,N_1149);
and U1226 (N_1226,N_1175,N_1145);
or U1227 (N_1227,N_1188,N_1189);
xor U1228 (N_1228,N_1131,N_1199);
and U1229 (N_1229,N_1186,N_1137);
nand U1230 (N_1230,N_1133,N_1147);
nand U1231 (N_1231,N_1181,N_1142);
nand U1232 (N_1232,N_1168,N_1126);
and U1233 (N_1233,N_1184,N_1167);
nor U1234 (N_1234,N_1146,N_1183);
nand U1235 (N_1235,N_1177,N_1165);
xor U1236 (N_1236,N_1196,N_1129);
nand U1237 (N_1237,N_1174,N_1134);
nor U1238 (N_1238,N_1128,N_1164);
xnor U1239 (N_1239,N_1146,N_1180);
nor U1240 (N_1240,N_1166,N_1129);
and U1241 (N_1241,N_1167,N_1128);
and U1242 (N_1242,N_1150,N_1136);
and U1243 (N_1243,N_1171,N_1188);
nor U1244 (N_1244,N_1174,N_1139);
or U1245 (N_1245,N_1154,N_1140);
or U1246 (N_1246,N_1187,N_1199);
nand U1247 (N_1247,N_1165,N_1161);
nand U1248 (N_1248,N_1158,N_1139);
and U1249 (N_1249,N_1141,N_1180);
nand U1250 (N_1250,N_1157,N_1153);
nor U1251 (N_1251,N_1144,N_1142);
nand U1252 (N_1252,N_1137,N_1199);
and U1253 (N_1253,N_1184,N_1190);
or U1254 (N_1254,N_1171,N_1195);
nor U1255 (N_1255,N_1179,N_1170);
nand U1256 (N_1256,N_1139,N_1154);
or U1257 (N_1257,N_1188,N_1179);
nor U1258 (N_1258,N_1172,N_1189);
and U1259 (N_1259,N_1174,N_1141);
or U1260 (N_1260,N_1129,N_1163);
nor U1261 (N_1261,N_1182,N_1150);
nand U1262 (N_1262,N_1166,N_1127);
nand U1263 (N_1263,N_1189,N_1171);
nor U1264 (N_1264,N_1182,N_1154);
or U1265 (N_1265,N_1150,N_1176);
nand U1266 (N_1266,N_1137,N_1195);
and U1267 (N_1267,N_1180,N_1139);
and U1268 (N_1268,N_1157,N_1179);
or U1269 (N_1269,N_1148,N_1126);
or U1270 (N_1270,N_1179,N_1149);
or U1271 (N_1271,N_1189,N_1141);
or U1272 (N_1272,N_1187,N_1164);
or U1273 (N_1273,N_1198,N_1174);
or U1274 (N_1274,N_1155,N_1190);
nor U1275 (N_1275,N_1225,N_1240);
xnor U1276 (N_1276,N_1268,N_1272);
nor U1277 (N_1277,N_1250,N_1200);
nor U1278 (N_1278,N_1245,N_1261);
and U1279 (N_1279,N_1216,N_1253);
nor U1280 (N_1280,N_1243,N_1238);
and U1281 (N_1281,N_1235,N_1227);
and U1282 (N_1282,N_1274,N_1260);
nand U1283 (N_1283,N_1271,N_1257);
nor U1284 (N_1284,N_1208,N_1244);
and U1285 (N_1285,N_1218,N_1246);
or U1286 (N_1286,N_1255,N_1234);
and U1287 (N_1287,N_1259,N_1210);
and U1288 (N_1288,N_1270,N_1202);
nor U1289 (N_1289,N_1206,N_1262);
and U1290 (N_1290,N_1229,N_1264);
or U1291 (N_1291,N_1267,N_1247);
and U1292 (N_1292,N_1242,N_1248);
and U1293 (N_1293,N_1205,N_1252);
and U1294 (N_1294,N_1221,N_1207);
nand U1295 (N_1295,N_1251,N_1211);
or U1296 (N_1296,N_1241,N_1231);
nor U1297 (N_1297,N_1217,N_1204);
or U1298 (N_1298,N_1273,N_1228);
nand U1299 (N_1299,N_1266,N_1203);
nor U1300 (N_1300,N_1212,N_1239);
nor U1301 (N_1301,N_1213,N_1222);
or U1302 (N_1302,N_1265,N_1219);
or U1303 (N_1303,N_1249,N_1258);
nor U1304 (N_1304,N_1220,N_1256);
and U1305 (N_1305,N_1236,N_1263);
and U1306 (N_1306,N_1224,N_1269);
nor U1307 (N_1307,N_1223,N_1237);
nor U1308 (N_1308,N_1215,N_1214);
or U1309 (N_1309,N_1254,N_1233);
and U1310 (N_1310,N_1209,N_1226);
nand U1311 (N_1311,N_1232,N_1230);
and U1312 (N_1312,N_1201,N_1237);
nor U1313 (N_1313,N_1201,N_1242);
nor U1314 (N_1314,N_1235,N_1236);
or U1315 (N_1315,N_1230,N_1266);
nor U1316 (N_1316,N_1266,N_1228);
nor U1317 (N_1317,N_1247,N_1254);
and U1318 (N_1318,N_1273,N_1222);
or U1319 (N_1319,N_1200,N_1221);
and U1320 (N_1320,N_1210,N_1262);
nand U1321 (N_1321,N_1215,N_1213);
nand U1322 (N_1322,N_1251,N_1202);
nor U1323 (N_1323,N_1264,N_1254);
and U1324 (N_1324,N_1251,N_1231);
and U1325 (N_1325,N_1212,N_1265);
nand U1326 (N_1326,N_1217,N_1215);
nor U1327 (N_1327,N_1254,N_1208);
nand U1328 (N_1328,N_1212,N_1232);
nor U1329 (N_1329,N_1247,N_1253);
or U1330 (N_1330,N_1207,N_1227);
and U1331 (N_1331,N_1262,N_1273);
and U1332 (N_1332,N_1253,N_1217);
or U1333 (N_1333,N_1247,N_1263);
and U1334 (N_1334,N_1261,N_1210);
and U1335 (N_1335,N_1243,N_1203);
xor U1336 (N_1336,N_1260,N_1219);
or U1337 (N_1337,N_1209,N_1265);
nand U1338 (N_1338,N_1247,N_1266);
and U1339 (N_1339,N_1209,N_1242);
nor U1340 (N_1340,N_1209,N_1267);
xnor U1341 (N_1341,N_1224,N_1241);
nor U1342 (N_1342,N_1261,N_1255);
and U1343 (N_1343,N_1269,N_1237);
or U1344 (N_1344,N_1238,N_1246);
nand U1345 (N_1345,N_1244,N_1254);
and U1346 (N_1346,N_1204,N_1211);
and U1347 (N_1347,N_1241,N_1232);
nand U1348 (N_1348,N_1229,N_1256);
nand U1349 (N_1349,N_1222,N_1229);
nand U1350 (N_1350,N_1305,N_1325);
nand U1351 (N_1351,N_1292,N_1300);
nand U1352 (N_1352,N_1348,N_1313);
or U1353 (N_1353,N_1320,N_1344);
and U1354 (N_1354,N_1327,N_1307);
nand U1355 (N_1355,N_1346,N_1330);
nor U1356 (N_1356,N_1303,N_1279);
or U1357 (N_1357,N_1339,N_1287);
nand U1358 (N_1358,N_1321,N_1311);
nor U1359 (N_1359,N_1317,N_1302);
xnor U1360 (N_1360,N_1324,N_1290);
xor U1361 (N_1361,N_1291,N_1341);
nand U1362 (N_1362,N_1280,N_1277);
nor U1363 (N_1363,N_1296,N_1336);
or U1364 (N_1364,N_1276,N_1282);
and U1365 (N_1365,N_1319,N_1316);
nor U1366 (N_1366,N_1308,N_1284);
nor U1367 (N_1367,N_1289,N_1306);
nand U1368 (N_1368,N_1275,N_1334);
or U1369 (N_1369,N_1295,N_1298);
and U1370 (N_1370,N_1345,N_1342);
or U1371 (N_1371,N_1318,N_1301);
and U1372 (N_1372,N_1312,N_1338);
nor U1373 (N_1373,N_1322,N_1304);
or U1374 (N_1374,N_1340,N_1294);
nand U1375 (N_1375,N_1337,N_1349);
and U1376 (N_1376,N_1343,N_1326);
or U1377 (N_1377,N_1328,N_1281);
or U1378 (N_1378,N_1323,N_1347);
nand U1379 (N_1379,N_1310,N_1335);
or U1380 (N_1380,N_1333,N_1309);
nor U1381 (N_1381,N_1278,N_1293);
and U1382 (N_1382,N_1283,N_1297);
nand U1383 (N_1383,N_1288,N_1285);
or U1384 (N_1384,N_1299,N_1329);
nor U1385 (N_1385,N_1314,N_1332);
or U1386 (N_1386,N_1331,N_1315);
or U1387 (N_1387,N_1286,N_1295);
or U1388 (N_1388,N_1303,N_1286);
or U1389 (N_1389,N_1284,N_1311);
nand U1390 (N_1390,N_1291,N_1323);
nor U1391 (N_1391,N_1284,N_1295);
and U1392 (N_1392,N_1327,N_1287);
nand U1393 (N_1393,N_1329,N_1284);
nor U1394 (N_1394,N_1322,N_1286);
and U1395 (N_1395,N_1298,N_1315);
and U1396 (N_1396,N_1311,N_1296);
nor U1397 (N_1397,N_1301,N_1297);
nor U1398 (N_1398,N_1318,N_1344);
nand U1399 (N_1399,N_1283,N_1298);
nand U1400 (N_1400,N_1284,N_1283);
nor U1401 (N_1401,N_1310,N_1313);
and U1402 (N_1402,N_1318,N_1290);
nand U1403 (N_1403,N_1306,N_1333);
nor U1404 (N_1404,N_1335,N_1275);
and U1405 (N_1405,N_1312,N_1348);
nand U1406 (N_1406,N_1294,N_1287);
nand U1407 (N_1407,N_1317,N_1319);
nand U1408 (N_1408,N_1308,N_1311);
nand U1409 (N_1409,N_1321,N_1317);
nand U1410 (N_1410,N_1319,N_1321);
nor U1411 (N_1411,N_1281,N_1337);
and U1412 (N_1412,N_1319,N_1346);
or U1413 (N_1413,N_1320,N_1314);
nor U1414 (N_1414,N_1275,N_1318);
nand U1415 (N_1415,N_1293,N_1344);
nor U1416 (N_1416,N_1341,N_1278);
nor U1417 (N_1417,N_1330,N_1293);
nor U1418 (N_1418,N_1282,N_1310);
nor U1419 (N_1419,N_1310,N_1297);
and U1420 (N_1420,N_1339,N_1331);
or U1421 (N_1421,N_1331,N_1309);
and U1422 (N_1422,N_1290,N_1283);
nand U1423 (N_1423,N_1328,N_1282);
and U1424 (N_1424,N_1340,N_1326);
and U1425 (N_1425,N_1385,N_1416);
nand U1426 (N_1426,N_1398,N_1373);
nor U1427 (N_1427,N_1413,N_1396);
nand U1428 (N_1428,N_1382,N_1400);
or U1429 (N_1429,N_1423,N_1408);
nand U1430 (N_1430,N_1378,N_1401);
and U1431 (N_1431,N_1383,N_1357);
nand U1432 (N_1432,N_1368,N_1351);
nand U1433 (N_1433,N_1403,N_1404);
nor U1434 (N_1434,N_1419,N_1406);
and U1435 (N_1435,N_1374,N_1372);
nor U1436 (N_1436,N_1397,N_1392);
nand U1437 (N_1437,N_1358,N_1361);
or U1438 (N_1438,N_1424,N_1412);
nor U1439 (N_1439,N_1415,N_1367);
xor U1440 (N_1440,N_1370,N_1354);
nor U1441 (N_1441,N_1384,N_1389);
or U1442 (N_1442,N_1363,N_1411);
nor U1443 (N_1443,N_1420,N_1376);
or U1444 (N_1444,N_1422,N_1409);
nor U1445 (N_1445,N_1366,N_1377);
or U1446 (N_1446,N_1388,N_1410);
nand U1447 (N_1447,N_1418,N_1356);
and U1448 (N_1448,N_1402,N_1387);
xnor U1449 (N_1449,N_1417,N_1399);
nor U1450 (N_1450,N_1371,N_1421);
nor U1451 (N_1451,N_1375,N_1379);
or U1452 (N_1452,N_1359,N_1407);
nand U1453 (N_1453,N_1393,N_1394);
nand U1454 (N_1454,N_1395,N_1365);
or U1455 (N_1455,N_1360,N_1390);
or U1456 (N_1456,N_1380,N_1391);
or U1457 (N_1457,N_1369,N_1364);
nand U1458 (N_1458,N_1381,N_1353);
or U1459 (N_1459,N_1414,N_1386);
and U1460 (N_1460,N_1350,N_1352);
and U1461 (N_1461,N_1355,N_1405);
and U1462 (N_1462,N_1362,N_1389);
nor U1463 (N_1463,N_1370,N_1413);
and U1464 (N_1464,N_1387,N_1407);
nor U1465 (N_1465,N_1412,N_1419);
nor U1466 (N_1466,N_1378,N_1381);
or U1467 (N_1467,N_1367,N_1353);
and U1468 (N_1468,N_1390,N_1419);
and U1469 (N_1469,N_1390,N_1374);
nand U1470 (N_1470,N_1419,N_1365);
nor U1471 (N_1471,N_1351,N_1389);
or U1472 (N_1472,N_1408,N_1414);
nor U1473 (N_1473,N_1419,N_1351);
nor U1474 (N_1474,N_1422,N_1421);
or U1475 (N_1475,N_1366,N_1414);
or U1476 (N_1476,N_1384,N_1370);
and U1477 (N_1477,N_1409,N_1418);
nor U1478 (N_1478,N_1410,N_1359);
nor U1479 (N_1479,N_1378,N_1409);
nor U1480 (N_1480,N_1381,N_1351);
or U1481 (N_1481,N_1362,N_1352);
or U1482 (N_1482,N_1361,N_1367);
nand U1483 (N_1483,N_1393,N_1423);
or U1484 (N_1484,N_1358,N_1373);
nand U1485 (N_1485,N_1424,N_1409);
or U1486 (N_1486,N_1395,N_1410);
and U1487 (N_1487,N_1354,N_1416);
and U1488 (N_1488,N_1399,N_1386);
and U1489 (N_1489,N_1409,N_1373);
and U1490 (N_1490,N_1364,N_1415);
nand U1491 (N_1491,N_1363,N_1414);
and U1492 (N_1492,N_1356,N_1351);
nor U1493 (N_1493,N_1360,N_1404);
or U1494 (N_1494,N_1365,N_1408);
nor U1495 (N_1495,N_1352,N_1382);
nand U1496 (N_1496,N_1406,N_1386);
nor U1497 (N_1497,N_1384,N_1367);
nor U1498 (N_1498,N_1366,N_1396);
or U1499 (N_1499,N_1371,N_1390);
nand U1500 (N_1500,N_1426,N_1496);
nor U1501 (N_1501,N_1492,N_1462);
or U1502 (N_1502,N_1493,N_1434);
and U1503 (N_1503,N_1475,N_1445);
nand U1504 (N_1504,N_1464,N_1483);
or U1505 (N_1505,N_1490,N_1468);
or U1506 (N_1506,N_1436,N_1440);
nor U1507 (N_1507,N_1478,N_1441);
and U1508 (N_1508,N_1487,N_1469);
nor U1509 (N_1509,N_1453,N_1474);
or U1510 (N_1510,N_1473,N_1437);
and U1511 (N_1511,N_1489,N_1444);
nand U1512 (N_1512,N_1481,N_1472);
nor U1513 (N_1513,N_1463,N_1433);
nor U1514 (N_1514,N_1470,N_1448);
and U1515 (N_1515,N_1457,N_1425);
nand U1516 (N_1516,N_1480,N_1494);
nand U1517 (N_1517,N_1446,N_1455);
or U1518 (N_1518,N_1430,N_1467);
and U1519 (N_1519,N_1498,N_1465);
nand U1520 (N_1520,N_1497,N_1499);
or U1521 (N_1521,N_1442,N_1431);
or U1522 (N_1522,N_1439,N_1485);
nand U1523 (N_1523,N_1459,N_1447);
nand U1524 (N_1524,N_1458,N_1466);
and U1525 (N_1525,N_1488,N_1479);
and U1526 (N_1526,N_1476,N_1491);
and U1527 (N_1527,N_1495,N_1449);
and U1528 (N_1528,N_1451,N_1461);
and U1529 (N_1529,N_1450,N_1438);
or U1530 (N_1530,N_1471,N_1435);
nor U1531 (N_1531,N_1428,N_1454);
nor U1532 (N_1532,N_1432,N_1429);
or U1533 (N_1533,N_1427,N_1456);
and U1534 (N_1534,N_1486,N_1460);
nor U1535 (N_1535,N_1443,N_1484);
and U1536 (N_1536,N_1482,N_1477);
nor U1537 (N_1537,N_1452,N_1446);
nor U1538 (N_1538,N_1459,N_1442);
or U1539 (N_1539,N_1431,N_1434);
and U1540 (N_1540,N_1487,N_1496);
and U1541 (N_1541,N_1486,N_1438);
or U1542 (N_1542,N_1433,N_1476);
and U1543 (N_1543,N_1476,N_1442);
nor U1544 (N_1544,N_1458,N_1433);
and U1545 (N_1545,N_1447,N_1488);
and U1546 (N_1546,N_1428,N_1445);
nor U1547 (N_1547,N_1461,N_1486);
and U1548 (N_1548,N_1480,N_1431);
nor U1549 (N_1549,N_1440,N_1431);
nor U1550 (N_1550,N_1472,N_1492);
and U1551 (N_1551,N_1476,N_1445);
nor U1552 (N_1552,N_1433,N_1449);
nand U1553 (N_1553,N_1475,N_1426);
nor U1554 (N_1554,N_1482,N_1497);
or U1555 (N_1555,N_1431,N_1474);
xor U1556 (N_1556,N_1451,N_1490);
nor U1557 (N_1557,N_1480,N_1455);
and U1558 (N_1558,N_1454,N_1498);
or U1559 (N_1559,N_1426,N_1491);
or U1560 (N_1560,N_1476,N_1496);
and U1561 (N_1561,N_1498,N_1485);
and U1562 (N_1562,N_1467,N_1484);
and U1563 (N_1563,N_1470,N_1482);
nor U1564 (N_1564,N_1476,N_1470);
and U1565 (N_1565,N_1476,N_1426);
and U1566 (N_1566,N_1463,N_1444);
or U1567 (N_1567,N_1434,N_1439);
or U1568 (N_1568,N_1439,N_1481);
or U1569 (N_1569,N_1451,N_1430);
or U1570 (N_1570,N_1484,N_1486);
or U1571 (N_1571,N_1471,N_1494);
or U1572 (N_1572,N_1466,N_1474);
or U1573 (N_1573,N_1429,N_1486);
nand U1574 (N_1574,N_1478,N_1450);
nor U1575 (N_1575,N_1539,N_1551);
nor U1576 (N_1576,N_1520,N_1555);
and U1577 (N_1577,N_1535,N_1568);
and U1578 (N_1578,N_1558,N_1559);
and U1579 (N_1579,N_1511,N_1543);
nor U1580 (N_1580,N_1506,N_1532);
and U1581 (N_1581,N_1552,N_1529);
nand U1582 (N_1582,N_1534,N_1567);
or U1583 (N_1583,N_1565,N_1556);
nand U1584 (N_1584,N_1564,N_1547);
or U1585 (N_1585,N_1508,N_1530);
nand U1586 (N_1586,N_1516,N_1544);
nand U1587 (N_1587,N_1554,N_1522);
or U1588 (N_1588,N_1570,N_1509);
nor U1589 (N_1589,N_1546,N_1507);
and U1590 (N_1590,N_1571,N_1501);
and U1591 (N_1591,N_1525,N_1521);
or U1592 (N_1592,N_1536,N_1569);
and U1593 (N_1593,N_1526,N_1514);
xnor U1594 (N_1594,N_1553,N_1573);
and U1595 (N_1595,N_1561,N_1538);
nor U1596 (N_1596,N_1505,N_1510);
and U1597 (N_1597,N_1519,N_1515);
nand U1598 (N_1598,N_1566,N_1549);
xnor U1599 (N_1599,N_1537,N_1517);
or U1600 (N_1600,N_1500,N_1531);
or U1601 (N_1601,N_1563,N_1548);
or U1602 (N_1602,N_1512,N_1557);
nand U1603 (N_1603,N_1528,N_1542);
nand U1604 (N_1604,N_1518,N_1502);
and U1605 (N_1605,N_1540,N_1503);
xnor U1606 (N_1606,N_1504,N_1574);
nand U1607 (N_1607,N_1545,N_1562);
nor U1608 (N_1608,N_1541,N_1533);
nand U1609 (N_1609,N_1524,N_1550);
nor U1610 (N_1610,N_1527,N_1572);
nand U1611 (N_1611,N_1513,N_1560);
and U1612 (N_1612,N_1523,N_1548);
nand U1613 (N_1613,N_1551,N_1574);
and U1614 (N_1614,N_1536,N_1554);
nor U1615 (N_1615,N_1507,N_1554);
nand U1616 (N_1616,N_1530,N_1555);
nor U1617 (N_1617,N_1525,N_1541);
or U1618 (N_1618,N_1535,N_1563);
nor U1619 (N_1619,N_1505,N_1574);
or U1620 (N_1620,N_1523,N_1561);
or U1621 (N_1621,N_1503,N_1528);
nand U1622 (N_1622,N_1546,N_1556);
and U1623 (N_1623,N_1538,N_1562);
nand U1624 (N_1624,N_1516,N_1537);
and U1625 (N_1625,N_1515,N_1549);
or U1626 (N_1626,N_1524,N_1564);
xor U1627 (N_1627,N_1503,N_1515);
or U1628 (N_1628,N_1512,N_1532);
nor U1629 (N_1629,N_1506,N_1547);
or U1630 (N_1630,N_1552,N_1536);
or U1631 (N_1631,N_1567,N_1572);
nand U1632 (N_1632,N_1565,N_1526);
nand U1633 (N_1633,N_1562,N_1515);
nor U1634 (N_1634,N_1519,N_1568);
nor U1635 (N_1635,N_1536,N_1505);
or U1636 (N_1636,N_1568,N_1533);
and U1637 (N_1637,N_1524,N_1541);
nor U1638 (N_1638,N_1536,N_1564);
xor U1639 (N_1639,N_1508,N_1547);
nand U1640 (N_1640,N_1500,N_1574);
or U1641 (N_1641,N_1513,N_1501);
or U1642 (N_1642,N_1507,N_1509);
nor U1643 (N_1643,N_1542,N_1535);
and U1644 (N_1644,N_1551,N_1514);
nand U1645 (N_1645,N_1519,N_1523);
or U1646 (N_1646,N_1546,N_1555);
nor U1647 (N_1647,N_1528,N_1572);
or U1648 (N_1648,N_1502,N_1566);
nand U1649 (N_1649,N_1567,N_1508);
and U1650 (N_1650,N_1583,N_1599);
or U1651 (N_1651,N_1633,N_1619);
nand U1652 (N_1652,N_1594,N_1644);
and U1653 (N_1653,N_1609,N_1641);
or U1654 (N_1654,N_1611,N_1635);
or U1655 (N_1655,N_1595,N_1616);
nand U1656 (N_1656,N_1585,N_1590);
nor U1657 (N_1657,N_1601,N_1618);
and U1658 (N_1658,N_1578,N_1642);
nand U1659 (N_1659,N_1626,N_1605);
nor U1660 (N_1660,N_1587,N_1596);
nand U1661 (N_1661,N_1636,N_1612);
nand U1662 (N_1662,N_1593,N_1584);
xnor U1663 (N_1663,N_1648,N_1588);
nor U1664 (N_1664,N_1625,N_1598);
or U1665 (N_1665,N_1643,N_1576);
or U1666 (N_1666,N_1606,N_1575);
or U1667 (N_1667,N_1604,N_1645);
and U1668 (N_1668,N_1637,N_1586);
nor U1669 (N_1669,N_1589,N_1603);
and U1670 (N_1670,N_1621,N_1582);
nor U1671 (N_1671,N_1577,N_1613);
and U1672 (N_1672,N_1602,N_1580);
nor U1673 (N_1673,N_1617,N_1591);
or U1674 (N_1674,N_1630,N_1622);
nor U1675 (N_1675,N_1592,N_1607);
and U1676 (N_1676,N_1597,N_1629);
and U1677 (N_1677,N_1649,N_1600);
nor U1678 (N_1678,N_1615,N_1624);
or U1679 (N_1679,N_1628,N_1638);
nor U1680 (N_1680,N_1610,N_1608);
or U1681 (N_1681,N_1632,N_1623);
or U1682 (N_1682,N_1627,N_1646);
nand U1683 (N_1683,N_1634,N_1620);
nor U1684 (N_1684,N_1579,N_1639);
nand U1685 (N_1685,N_1631,N_1614);
nor U1686 (N_1686,N_1647,N_1581);
and U1687 (N_1687,N_1640,N_1607);
and U1688 (N_1688,N_1635,N_1614);
nor U1689 (N_1689,N_1583,N_1629);
nand U1690 (N_1690,N_1634,N_1583);
nor U1691 (N_1691,N_1635,N_1640);
or U1692 (N_1692,N_1584,N_1592);
nor U1693 (N_1693,N_1595,N_1604);
or U1694 (N_1694,N_1579,N_1601);
nand U1695 (N_1695,N_1625,N_1635);
nor U1696 (N_1696,N_1578,N_1580);
nor U1697 (N_1697,N_1630,N_1586);
nand U1698 (N_1698,N_1640,N_1636);
or U1699 (N_1699,N_1607,N_1600);
or U1700 (N_1700,N_1598,N_1622);
and U1701 (N_1701,N_1649,N_1582);
nor U1702 (N_1702,N_1598,N_1648);
or U1703 (N_1703,N_1598,N_1606);
xor U1704 (N_1704,N_1621,N_1635);
nand U1705 (N_1705,N_1590,N_1603);
or U1706 (N_1706,N_1579,N_1628);
and U1707 (N_1707,N_1614,N_1643);
nand U1708 (N_1708,N_1599,N_1640);
and U1709 (N_1709,N_1575,N_1631);
or U1710 (N_1710,N_1601,N_1603);
and U1711 (N_1711,N_1577,N_1624);
nor U1712 (N_1712,N_1596,N_1619);
nor U1713 (N_1713,N_1624,N_1583);
nand U1714 (N_1714,N_1622,N_1594);
nor U1715 (N_1715,N_1575,N_1580);
nand U1716 (N_1716,N_1594,N_1576);
and U1717 (N_1717,N_1632,N_1625);
nand U1718 (N_1718,N_1578,N_1628);
or U1719 (N_1719,N_1604,N_1647);
and U1720 (N_1720,N_1612,N_1622);
and U1721 (N_1721,N_1636,N_1632);
nor U1722 (N_1722,N_1618,N_1597);
nor U1723 (N_1723,N_1600,N_1614);
nand U1724 (N_1724,N_1646,N_1620);
and U1725 (N_1725,N_1709,N_1667);
or U1726 (N_1726,N_1722,N_1660);
nor U1727 (N_1727,N_1657,N_1673);
and U1728 (N_1728,N_1708,N_1712);
or U1729 (N_1729,N_1706,N_1698);
or U1730 (N_1730,N_1688,N_1680);
nand U1731 (N_1731,N_1677,N_1717);
nand U1732 (N_1732,N_1691,N_1699);
or U1733 (N_1733,N_1696,N_1681);
nor U1734 (N_1734,N_1675,N_1676);
nand U1735 (N_1735,N_1694,N_1672);
or U1736 (N_1736,N_1656,N_1690);
and U1737 (N_1737,N_1707,N_1679);
and U1738 (N_1738,N_1713,N_1669);
or U1739 (N_1739,N_1674,N_1670);
and U1740 (N_1740,N_1697,N_1711);
nand U1741 (N_1741,N_1651,N_1684);
or U1742 (N_1742,N_1650,N_1723);
and U1743 (N_1743,N_1720,N_1714);
or U1744 (N_1744,N_1715,N_1701);
nand U1745 (N_1745,N_1653,N_1658);
or U1746 (N_1746,N_1710,N_1683);
and U1747 (N_1747,N_1687,N_1659);
nor U1748 (N_1748,N_1721,N_1703);
or U1749 (N_1749,N_1671,N_1695);
or U1750 (N_1750,N_1700,N_1682);
or U1751 (N_1751,N_1655,N_1702);
or U1752 (N_1752,N_1719,N_1663);
nor U1753 (N_1753,N_1652,N_1662);
and U1754 (N_1754,N_1724,N_1718);
and U1755 (N_1755,N_1704,N_1666);
or U1756 (N_1756,N_1716,N_1705);
nor U1757 (N_1757,N_1686,N_1661);
nand U1758 (N_1758,N_1689,N_1668);
nand U1759 (N_1759,N_1693,N_1678);
and U1760 (N_1760,N_1664,N_1685);
nand U1761 (N_1761,N_1654,N_1665);
nor U1762 (N_1762,N_1692,N_1654);
nand U1763 (N_1763,N_1683,N_1698);
or U1764 (N_1764,N_1665,N_1651);
and U1765 (N_1765,N_1656,N_1682);
nor U1766 (N_1766,N_1705,N_1675);
nor U1767 (N_1767,N_1682,N_1674);
nor U1768 (N_1768,N_1696,N_1708);
nor U1769 (N_1769,N_1711,N_1694);
or U1770 (N_1770,N_1660,N_1720);
nor U1771 (N_1771,N_1669,N_1660);
and U1772 (N_1772,N_1708,N_1682);
nor U1773 (N_1773,N_1722,N_1683);
nand U1774 (N_1774,N_1678,N_1686);
or U1775 (N_1775,N_1711,N_1658);
nand U1776 (N_1776,N_1697,N_1677);
or U1777 (N_1777,N_1653,N_1707);
or U1778 (N_1778,N_1687,N_1720);
nand U1779 (N_1779,N_1691,N_1658);
and U1780 (N_1780,N_1656,N_1661);
or U1781 (N_1781,N_1688,N_1698);
and U1782 (N_1782,N_1675,N_1686);
nor U1783 (N_1783,N_1703,N_1719);
or U1784 (N_1784,N_1697,N_1655);
or U1785 (N_1785,N_1670,N_1660);
and U1786 (N_1786,N_1699,N_1698);
nor U1787 (N_1787,N_1684,N_1721);
and U1788 (N_1788,N_1685,N_1667);
or U1789 (N_1789,N_1708,N_1680);
and U1790 (N_1790,N_1658,N_1713);
and U1791 (N_1791,N_1705,N_1681);
nor U1792 (N_1792,N_1710,N_1656);
and U1793 (N_1793,N_1706,N_1669);
nand U1794 (N_1794,N_1695,N_1720);
nand U1795 (N_1795,N_1666,N_1670);
or U1796 (N_1796,N_1663,N_1720);
or U1797 (N_1797,N_1696,N_1668);
nand U1798 (N_1798,N_1656,N_1694);
nor U1799 (N_1799,N_1697,N_1663);
nor U1800 (N_1800,N_1737,N_1781);
or U1801 (N_1801,N_1750,N_1747);
nand U1802 (N_1802,N_1783,N_1787);
nand U1803 (N_1803,N_1752,N_1780);
and U1804 (N_1804,N_1771,N_1775);
or U1805 (N_1805,N_1735,N_1782);
nor U1806 (N_1806,N_1785,N_1754);
nand U1807 (N_1807,N_1763,N_1796);
nand U1808 (N_1808,N_1769,N_1766);
nor U1809 (N_1809,N_1776,N_1764);
or U1810 (N_1810,N_1795,N_1773);
or U1811 (N_1811,N_1740,N_1728);
or U1812 (N_1812,N_1765,N_1727);
nor U1813 (N_1813,N_1733,N_1784);
nand U1814 (N_1814,N_1738,N_1788);
nor U1815 (N_1815,N_1748,N_1791);
and U1816 (N_1816,N_1793,N_1742);
nand U1817 (N_1817,N_1760,N_1761);
or U1818 (N_1818,N_1757,N_1753);
and U1819 (N_1819,N_1768,N_1797);
nand U1820 (N_1820,N_1734,N_1725);
and U1821 (N_1821,N_1751,N_1799);
nor U1822 (N_1822,N_1794,N_1762);
nor U1823 (N_1823,N_1786,N_1729);
nor U1824 (N_1824,N_1767,N_1758);
or U1825 (N_1825,N_1744,N_1730);
nor U1826 (N_1826,N_1759,N_1726);
or U1827 (N_1827,N_1743,N_1770);
and U1828 (N_1828,N_1792,N_1790);
nand U1829 (N_1829,N_1777,N_1779);
and U1830 (N_1830,N_1741,N_1732);
or U1831 (N_1831,N_1798,N_1745);
nand U1832 (N_1832,N_1739,N_1731);
or U1833 (N_1833,N_1749,N_1756);
nand U1834 (N_1834,N_1774,N_1772);
nor U1835 (N_1835,N_1755,N_1736);
or U1836 (N_1836,N_1778,N_1746);
nor U1837 (N_1837,N_1789,N_1799);
or U1838 (N_1838,N_1757,N_1782);
and U1839 (N_1839,N_1756,N_1797);
or U1840 (N_1840,N_1728,N_1753);
nor U1841 (N_1841,N_1792,N_1745);
nor U1842 (N_1842,N_1754,N_1760);
nand U1843 (N_1843,N_1751,N_1788);
nand U1844 (N_1844,N_1736,N_1729);
nand U1845 (N_1845,N_1764,N_1781);
nor U1846 (N_1846,N_1749,N_1790);
or U1847 (N_1847,N_1792,N_1782);
nor U1848 (N_1848,N_1763,N_1742);
nor U1849 (N_1849,N_1785,N_1783);
or U1850 (N_1850,N_1726,N_1754);
nor U1851 (N_1851,N_1735,N_1769);
or U1852 (N_1852,N_1796,N_1746);
and U1853 (N_1853,N_1762,N_1755);
nand U1854 (N_1854,N_1773,N_1736);
or U1855 (N_1855,N_1766,N_1778);
nor U1856 (N_1856,N_1760,N_1782);
or U1857 (N_1857,N_1796,N_1783);
nand U1858 (N_1858,N_1777,N_1763);
nor U1859 (N_1859,N_1733,N_1786);
or U1860 (N_1860,N_1726,N_1788);
nor U1861 (N_1861,N_1757,N_1767);
or U1862 (N_1862,N_1763,N_1791);
or U1863 (N_1863,N_1782,N_1767);
nor U1864 (N_1864,N_1771,N_1785);
nand U1865 (N_1865,N_1748,N_1764);
or U1866 (N_1866,N_1769,N_1788);
and U1867 (N_1867,N_1790,N_1778);
or U1868 (N_1868,N_1797,N_1729);
or U1869 (N_1869,N_1737,N_1726);
and U1870 (N_1870,N_1763,N_1790);
nor U1871 (N_1871,N_1782,N_1725);
nand U1872 (N_1872,N_1759,N_1736);
nand U1873 (N_1873,N_1725,N_1799);
or U1874 (N_1874,N_1776,N_1752);
and U1875 (N_1875,N_1848,N_1851);
nor U1876 (N_1876,N_1850,N_1838);
and U1877 (N_1877,N_1818,N_1814);
nor U1878 (N_1878,N_1820,N_1816);
or U1879 (N_1879,N_1866,N_1823);
and U1880 (N_1880,N_1874,N_1858);
or U1881 (N_1881,N_1811,N_1841);
nor U1882 (N_1882,N_1821,N_1804);
and U1883 (N_1883,N_1831,N_1809);
or U1884 (N_1884,N_1819,N_1855);
xnor U1885 (N_1885,N_1810,N_1863);
nor U1886 (N_1886,N_1857,N_1853);
nand U1887 (N_1887,N_1812,N_1844);
nand U1888 (N_1888,N_1807,N_1822);
and U1889 (N_1889,N_1861,N_1830);
or U1890 (N_1890,N_1872,N_1828);
or U1891 (N_1891,N_1832,N_1849);
nor U1892 (N_1892,N_1871,N_1840);
or U1893 (N_1893,N_1865,N_1827);
nor U1894 (N_1894,N_1808,N_1847);
or U1895 (N_1895,N_1825,N_1860);
or U1896 (N_1896,N_1829,N_1864);
nor U1897 (N_1897,N_1852,N_1873);
and U1898 (N_1898,N_1805,N_1801);
nor U1899 (N_1899,N_1826,N_1800);
or U1900 (N_1900,N_1813,N_1839);
or U1901 (N_1901,N_1836,N_1806);
and U1902 (N_1902,N_1824,N_1837);
nand U1903 (N_1903,N_1870,N_1835);
nor U1904 (N_1904,N_1869,N_1859);
nor U1905 (N_1905,N_1834,N_1854);
nor U1906 (N_1906,N_1833,N_1802);
and U1907 (N_1907,N_1842,N_1846);
or U1908 (N_1908,N_1867,N_1843);
or U1909 (N_1909,N_1862,N_1803);
nand U1910 (N_1910,N_1868,N_1815);
nand U1911 (N_1911,N_1845,N_1856);
or U1912 (N_1912,N_1817,N_1862);
and U1913 (N_1913,N_1837,N_1861);
nor U1914 (N_1914,N_1828,N_1873);
and U1915 (N_1915,N_1826,N_1823);
and U1916 (N_1916,N_1828,N_1807);
nor U1917 (N_1917,N_1843,N_1847);
or U1918 (N_1918,N_1851,N_1861);
nor U1919 (N_1919,N_1803,N_1850);
and U1920 (N_1920,N_1816,N_1805);
nor U1921 (N_1921,N_1817,N_1870);
and U1922 (N_1922,N_1868,N_1802);
nand U1923 (N_1923,N_1813,N_1871);
nor U1924 (N_1924,N_1836,N_1847);
nor U1925 (N_1925,N_1827,N_1800);
or U1926 (N_1926,N_1836,N_1802);
and U1927 (N_1927,N_1861,N_1868);
nand U1928 (N_1928,N_1828,N_1806);
nor U1929 (N_1929,N_1824,N_1839);
and U1930 (N_1930,N_1860,N_1837);
nand U1931 (N_1931,N_1810,N_1860);
or U1932 (N_1932,N_1815,N_1801);
or U1933 (N_1933,N_1823,N_1867);
or U1934 (N_1934,N_1865,N_1830);
nand U1935 (N_1935,N_1802,N_1858);
nand U1936 (N_1936,N_1856,N_1865);
nand U1937 (N_1937,N_1811,N_1822);
and U1938 (N_1938,N_1845,N_1862);
or U1939 (N_1939,N_1859,N_1835);
xnor U1940 (N_1940,N_1812,N_1800);
or U1941 (N_1941,N_1803,N_1812);
nand U1942 (N_1942,N_1872,N_1858);
or U1943 (N_1943,N_1844,N_1822);
nor U1944 (N_1944,N_1849,N_1871);
nand U1945 (N_1945,N_1868,N_1826);
xor U1946 (N_1946,N_1807,N_1874);
nand U1947 (N_1947,N_1851,N_1866);
and U1948 (N_1948,N_1816,N_1851);
nor U1949 (N_1949,N_1834,N_1861);
nor U1950 (N_1950,N_1875,N_1902);
or U1951 (N_1951,N_1932,N_1887);
or U1952 (N_1952,N_1886,N_1941);
nand U1953 (N_1953,N_1912,N_1925);
and U1954 (N_1954,N_1882,N_1944);
xnor U1955 (N_1955,N_1933,N_1949);
or U1956 (N_1956,N_1896,N_1888);
nor U1957 (N_1957,N_1945,N_1880);
nand U1958 (N_1958,N_1895,N_1921);
xor U1959 (N_1959,N_1917,N_1915);
nor U1960 (N_1960,N_1891,N_1938);
and U1961 (N_1961,N_1922,N_1930);
and U1962 (N_1962,N_1934,N_1911);
nand U1963 (N_1963,N_1884,N_1924);
nand U1964 (N_1964,N_1878,N_1910);
and U1965 (N_1965,N_1889,N_1928);
or U1966 (N_1966,N_1920,N_1879);
or U1967 (N_1967,N_1883,N_1901);
or U1968 (N_1968,N_1897,N_1926);
or U1969 (N_1969,N_1892,N_1877);
nand U1970 (N_1970,N_1885,N_1929);
xor U1971 (N_1971,N_1909,N_1907);
nor U1972 (N_1972,N_1900,N_1890);
nor U1973 (N_1973,N_1904,N_1899);
nand U1974 (N_1974,N_1903,N_1935);
and U1975 (N_1975,N_1918,N_1894);
and U1976 (N_1976,N_1881,N_1942);
nor U1977 (N_1977,N_1913,N_1940);
xnor U1978 (N_1978,N_1906,N_1919);
nor U1979 (N_1979,N_1923,N_1927);
and U1980 (N_1980,N_1916,N_1946);
nor U1981 (N_1981,N_1908,N_1914);
nand U1982 (N_1982,N_1947,N_1937);
nor U1983 (N_1983,N_1876,N_1893);
nand U1984 (N_1984,N_1948,N_1943);
nand U1985 (N_1985,N_1931,N_1898);
nor U1986 (N_1986,N_1939,N_1905);
or U1987 (N_1987,N_1936,N_1909);
or U1988 (N_1988,N_1878,N_1897);
or U1989 (N_1989,N_1911,N_1877);
and U1990 (N_1990,N_1946,N_1930);
nand U1991 (N_1991,N_1901,N_1905);
nor U1992 (N_1992,N_1879,N_1918);
and U1993 (N_1993,N_1888,N_1948);
nor U1994 (N_1994,N_1931,N_1944);
or U1995 (N_1995,N_1901,N_1922);
xor U1996 (N_1996,N_1922,N_1887);
nor U1997 (N_1997,N_1911,N_1924);
and U1998 (N_1998,N_1928,N_1891);
xor U1999 (N_1999,N_1887,N_1931);
and U2000 (N_2000,N_1935,N_1948);
and U2001 (N_2001,N_1917,N_1939);
and U2002 (N_2002,N_1904,N_1930);
and U2003 (N_2003,N_1928,N_1937);
or U2004 (N_2004,N_1923,N_1948);
xnor U2005 (N_2005,N_1917,N_1876);
and U2006 (N_2006,N_1903,N_1901);
or U2007 (N_2007,N_1879,N_1937);
or U2008 (N_2008,N_1931,N_1895);
xnor U2009 (N_2009,N_1897,N_1895);
or U2010 (N_2010,N_1907,N_1888);
nand U2011 (N_2011,N_1916,N_1932);
and U2012 (N_2012,N_1903,N_1909);
nor U2013 (N_2013,N_1880,N_1905);
nand U2014 (N_2014,N_1946,N_1906);
or U2015 (N_2015,N_1906,N_1901);
and U2016 (N_2016,N_1932,N_1908);
nand U2017 (N_2017,N_1893,N_1934);
and U2018 (N_2018,N_1931,N_1924);
or U2019 (N_2019,N_1924,N_1918);
nor U2020 (N_2020,N_1948,N_1879);
nand U2021 (N_2021,N_1941,N_1924);
and U2022 (N_2022,N_1905,N_1920);
nor U2023 (N_2023,N_1935,N_1933);
or U2024 (N_2024,N_1888,N_1942);
or U2025 (N_2025,N_2011,N_2020);
nor U2026 (N_2026,N_1968,N_1984);
nor U2027 (N_2027,N_1987,N_1972);
nand U2028 (N_2028,N_1970,N_1982);
nor U2029 (N_2029,N_1954,N_1957);
and U2030 (N_2030,N_1994,N_1963);
and U2031 (N_2031,N_1992,N_1976);
or U2032 (N_2032,N_2008,N_2007);
or U2033 (N_2033,N_1952,N_1995);
xor U2034 (N_2034,N_2024,N_1958);
nand U2035 (N_2035,N_1997,N_1950);
nand U2036 (N_2036,N_2023,N_1960);
and U2037 (N_2037,N_1986,N_1974);
or U2038 (N_2038,N_1990,N_2013);
and U2039 (N_2039,N_1953,N_2019);
nand U2040 (N_2040,N_1985,N_2017);
nor U2041 (N_2041,N_2015,N_2018);
nor U2042 (N_2042,N_1993,N_2021);
nand U2043 (N_2043,N_1979,N_2006);
nand U2044 (N_2044,N_1966,N_1977);
nand U2045 (N_2045,N_1975,N_1998);
nand U2046 (N_2046,N_1962,N_1981);
or U2047 (N_2047,N_2004,N_2016);
nand U2048 (N_2048,N_2022,N_1989);
and U2049 (N_2049,N_1964,N_2001);
nor U2050 (N_2050,N_1969,N_1978);
and U2051 (N_2051,N_2000,N_1996);
nand U2052 (N_2052,N_2010,N_2003);
nor U2053 (N_2053,N_1980,N_1956);
nor U2054 (N_2054,N_1971,N_2009);
nor U2055 (N_2055,N_1991,N_1961);
nor U2056 (N_2056,N_1951,N_2014);
xor U2057 (N_2057,N_1965,N_1959);
nand U2058 (N_2058,N_1955,N_2002);
nor U2059 (N_2059,N_1999,N_2012);
xor U2060 (N_2060,N_1983,N_1967);
nor U2061 (N_2061,N_1988,N_1973);
nand U2062 (N_2062,N_2005,N_1999);
nor U2063 (N_2063,N_2024,N_1963);
or U2064 (N_2064,N_2017,N_2005);
and U2065 (N_2065,N_2015,N_2024);
nor U2066 (N_2066,N_1993,N_1969);
and U2067 (N_2067,N_1986,N_2000);
and U2068 (N_2068,N_1983,N_1965);
or U2069 (N_2069,N_1954,N_1979);
nand U2070 (N_2070,N_1995,N_2002);
or U2071 (N_2071,N_1970,N_1992);
nor U2072 (N_2072,N_1965,N_1957);
nand U2073 (N_2073,N_1994,N_1999);
nor U2074 (N_2074,N_2020,N_1967);
or U2075 (N_2075,N_1963,N_1992);
nor U2076 (N_2076,N_1963,N_2021);
or U2077 (N_2077,N_1977,N_2002);
nor U2078 (N_2078,N_1972,N_1984);
and U2079 (N_2079,N_2008,N_1957);
nand U2080 (N_2080,N_2009,N_1999);
and U2081 (N_2081,N_2020,N_1959);
nand U2082 (N_2082,N_1956,N_2004);
or U2083 (N_2083,N_2005,N_2015);
nand U2084 (N_2084,N_2022,N_1991);
nand U2085 (N_2085,N_2022,N_1951);
and U2086 (N_2086,N_1956,N_1952);
or U2087 (N_2087,N_1956,N_2018);
or U2088 (N_2088,N_1973,N_2006);
and U2089 (N_2089,N_1986,N_1968);
nor U2090 (N_2090,N_1998,N_2007);
or U2091 (N_2091,N_1968,N_1956);
and U2092 (N_2092,N_1955,N_1962);
nor U2093 (N_2093,N_2010,N_1950);
nor U2094 (N_2094,N_1975,N_1966);
or U2095 (N_2095,N_1957,N_1975);
xor U2096 (N_2096,N_1985,N_2005);
nor U2097 (N_2097,N_1982,N_1951);
or U2098 (N_2098,N_2001,N_1979);
nor U2099 (N_2099,N_1995,N_2019);
or U2100 (N_2100,N_2044,N_2040);
or U2101 (N_2101,N_2027,N_2097);
nand U2102 (N_2102,N_2026,N_2060);
and U2103 (N_2103,N_2080,N_2069);
nand U2104 (N_2104,N_2085,N_2043);
xnor U2105 (N_2105,N_2054,N_2071);
nand U2106 (N_2106,N_2066,N_2050);
nor U2107 (N_2107,N_2061,N_2079);
and U2108 (N_2108,N_2049,N_2032);
nor U2109 (N_2109,N_2095,N_2041);
nor U2110 (N_2110,N_2099,N_2093);
xnor U2111 (N_2111,N_2056,N_2064);
or U2112 (N_2112,N_2098,N_2075);
or U2113 (N_2113,N_2030,N_2055);
nand U2114 (N_2114,N_2067,N_2028);
and U2115 (N_2115,N_2051,N_2089);
and U2116 (N_2116,N_2076,N_2081);
and U2117 (N_2117,N_2045,N_2094);
or U2118 (N_2118,N_2052,N_2031);
or U2119 (N_2119,N_2087,N_2086);
nand U2120 (N_2120,N_2062,N_2083);
nor U2121 (N_2121,N_2092,N_2074);
nand U2122 (N_2122,N_2036,N_2053);
nor U2123 (N_2123,N_2088,N_2084);
nand U2124 (N_2124,N_2029,N_2033);
nand U2125 (N_2125,N_2025,N_2042);
and U2126 (N_2126,N_2096,N_2065);
and U2127 (N_2127,N_2063,N_2077);
and U2128 (N_2128,N_2038,N_2035);
or U2129 (N_2129,N_2047,N_2073);
or U2130 (N_2130,N_2068,N_2072);
nand U2131 (N_2131,N_2034,N_2090);
and U2132 (N_2132,N_2058,N_2091);
and U2133 (N_2133,N_2046,N_2057);
or U2134 (N_2134,N_2039,N_2078);
nor U2135 (N_2135,N_2082,N_2070);
or U2136 (N_2136,N_2059,N_2037);
nand U2137 (N_2137,N_2048,N_2071);
nand U2138 (N_2138,N_2034,N_2083);
and U2139 (N_2139,N_2087,N_2096);
xor U2140 (N_2140,N_2061,N_2064);
or U2141 (N_2141,N_2079,N_2055);
or U2142 (N_2142,N_2066,N_2063);
or U2143 (N_2143,N_2090,N_2056);
nor U2144 (N_2144,N_2043,N_2051);
and U2145 (N_2145,N_2055,N_2044);
or U2146 (N_2146,N_2083,N_2080);
nand U2147 (N_2147,N_2093,N_2088);
nor U2148 (N_2148,N_2035,N_2055);
xor U2149 (N_2149,N_2088,N_2095);
and U2150 (N_2150,N_2030,N_2067);
and U2151 (N_2151,N_2092,N_2042);
nand U2152 (N_2152,N_2043,N_2098);
and U2153 (N_2153,N_2067,N_2078);
nor U2154 (N_2154,N_2058,N_2035);
nand U2155 (N_2155,N_2055,N_2053);
or U2156 (N_2156,N_2092,N_2083);
or U2157 (N_2157,N_2091,N_2044);
and U2158 (N_2158,N_2070,N_2058);
xnor U2159 (N_2159,N_2057,N_2075);
xor U2160 (N_2160,N_2085,N_2077);
and U2161 (N_2161,N_2041,N_2078);
and U2162 (N_2162,N_2048,N_2065);
or U2163 (N_2163,N_2060,N_2063);
and U2164 (N_2164,N_2027,N_2046);
nand U2165 (N_2165,N_2044,N_2070);
and U2166 (N_2166,N_2073,N_2096);
and U2167 (N_2167,N_2088,N_2026);
nand U2168 (N_2168,N_2096,N_2037);
or U2169 (N_2169,N_2062,N_2049);
nand U2170 (N_2170,N_2082,N_2049);
or U2171 (N_2171,N_2056,N_2050);
nand U2172 (N_2172,N_2026,N_2098);
nand U2173 (N_2173,N_2053,N_2099);
nor U2174 (N_2174,N_2057,N_2074);
and U2175 (N_2175,N_2101,N_2102);
xor U2176 (N_2176,N_2127,N_2148);
nand U2177 (N_2177,N_2111,N_2112);
nor U2178 (N_2178,N_2159,N_2110);
nor U2179 (N_2179,N_2122,N_2119);
or U2180 (N_2180,N_2174,N_2107);
nor U2181 (N_2181,N_2108,N_2168);
nand U2182 (N_2182,N_2155,N_2170);
nor U2183 (N_2183,N_2104,N_2134);
and U2184 (N_2184,N_2121,N_2128);
nand U2185 (N_2185,N_2139,N_2131);
nor U2186 (N_2186,N_2136,N_2106);
or U2187 (N_2187,N_2167,N_2163);
or U2188 (N_2188,N_2124,N_2162);
nand U2189 (N_2189,N_2116,N_2133);
and U2190 (N_2190,N_2156,N_2150);
nor U2191 (N_2191,N_2153,N_2160);
nor U2192 (N_2192,N_2138,N_2171);
nand U2193 (N_2193,N_2135,N_2164);
or U2194 (N_2194,N_2132,N_2109);
xnor U2195 (N_2195,N_2105,N_2166);
or U2196 (N_2196,N_2118,N_2114);
nand U2197 (N_2197,N_2161,N_2157);
or U2198 (N_2198,N_2143,N_2172);
nor U2199 (N_2199,N_2137,N_2130);
nor U2200 (N_2200,N_2117,N_2120);
nand U2201 (N_2201,N_2145,N_2158);
or U2202 (N_2202,N_2113,N_2140);
nor U2203 (N_2203,N_2149,N_2100);
nand U2204 (N_2204,N_2169,N_2129);
or U2205 (N_2205,N_2103,N_2126);
nor U2206 (N_2206,N_2144,N_2152);
or U2207 (N_2207,N_2142,N_2173);
and U2208 (N_2208,N_2165,N_2154);
nor U2209 (N_2209,N_2141,N_2151);
or U2210 (N_2210,N_2123,N_2115);
nor U2211 (N_2211,N_2125,N_2147);
or U2212 (N_2212,N_2146,N_2155);
nor U2213 (N_2213,N_2116,N_2144);
nand U2214 (N_2214,N_2163,N_2143);
and U2215 (N_2215,N_2143,N_2165);
or U2216 (N_2216,N_2115,N_2111);
and U2217 (N_2217,N_2145,N_2134);
or U2218 (N_2218,N_2161,N_2120);
nor U2219 (N_2219,N_2139,N_2161);
or U2220 (N_2220,N_2109,N_2125);
nor U2221 (N_2221,N_2105,N_2167);
or U2222 (N_2222,N_2122,N_2173);
nand U2223 (N_2223,N_2160,N_2109);
or U2224 (N_2224,N_2113,N_2138);
nand U2225 (N_2225,N_2150,N_2118);
nor U2226 (N_2226,N_2119,N_2162);
and U2227 (N_2227,N_2132,N_2173);
and U2228 (N_2228,N_2166,N_2136);
nand U2229 (N_2229,N_2130,N_2149);
nand U2230 (N_2230,N_2112,N_2154);
and U2231 (N_2231,N_2130,N_2100);
and U2232 (N_2232,N_2167,N_2125);
or U2233 (N_2233,N_2100,N_2123);
xor U2234 (N_2234,N_2149,N_2152);
or U2235 (N_2235,N_2133,N_2155);
and U2236 (N_2236,N_2155,N_2159);
or U2237 (N_2237,N_2172,N_2169);
or U2238 (N_2238,N_2150,N_2170);
or U2239 (N_2239,N_2169,N_2133);
nand U2240 (N_2240,N_2152,N_2132);
and U2241 (N_2241,N_2153,N_2149);
nand U2242 (N_2242,N_2163,N_2115);
nor U2243 (N_2243,N_2168,N_2161);
or U2244 (N_2244,N_2103,N_2144);
nand U2245 (N_2245,N_2129,N_2140);
and U2246 (N_2246,N_2171,N_2129);
nand U2247 (N_2247,N_2142,N_2147);
nand U2248 (N_2248,N_2149,N_2113);
or U2249 (N_2249,N_2111,N_2132);
nand U2250 (N_2250,N_2227,N_2182);
nor U2251 (N_2251,N_2226,N_2192);
and U2252 (N_2252,N_2215,N_2210);
nor U2253 (N_2253,N_2208,N_2243);
and U2254 (N_2254,N_2216,N_2184);
nor U2255 (N_2255,N_2235,N_2202);
or U2256 (N_2256,N_2189,N_2178);
nor U2257 (N_2257,N_2218,N_2193);
nor U2258 (N_2258,N_2214,N_2187);
and U2259 (N_2259,N_2236,N_2200);
nand U2260 (N_2260,N_2203,N_2185);
nor U2261 (N_2261,N_2247,N_2217);
or U2262 (N_2262,N_2199,N_2188);
nor U2263 (N_2263,N_2225,N_2237);
nand U2264 (N_2264,N_2205,N_2244);
nor U2265 (N_2265,N_2198,N_2239);
or U2266 (N_2266,N_2246,N_2219);
nor U2267 (N_2267,N_2221,N_2248);
and U2268 (N_2268,N_2233,N_2213);
or U2269 (N_2269,N_2211,N_2249);
nor U2270 (N_2270,N_2234,N_2231);
nor U2271 (N_2271,N_2197,N_2228);
nor U2272 (N_2272,N_2242,N_2201);
and U2273 (N_2273,N_2222,N_2212);
and U2274 (N_2274,N_2190,N_2245);
nand U2275 (N_2275,N_2206,N_2183);
nor U2276 (N_2276,N_2196,N_2180);
nor U2277 (N_2277,N_2195,N_2176);
nand U2278 (N_2278,N_2229,N_2181);
nand U2279 (N_2279,N_2207,N_2240);
nor U2280 (N_2280,N_2241,N_2204);
or U2281 (N_2281,N_2238,N_2230);
and U2282 (N_2282,N_2209,N_2177);
and U2283 (N_2283,N_2191,N_2220);
and U2284 (N_2284,N_2232,N_2179);
or U2285 (N_2285,N_2194,N_2175);
nand U2286 (N_2286,N_2186,N_2223);
and U2287 (N_2287,N_2224,N_2202);
nor U2288 (N_2288,N_2245,N_2243);
nand U2289 (N_2289,N_2199,N_2186);
nand U2290 (N_2290,N_2224,N_2223);
nor U2291 (N_2291,N_2180,N_2198);
and U2292 (N_2292,N_2194,N_2242);
or U2293 (N_2293,N_2213,N_2201);
and U2294 (N_2294,N_2231,N_2240);
and U2295 (N_2295,N_2220,N_2214);
nor U2296 (N_2296,N_2188,N_2228);
and U2297 (N_2297,N_2182,N_2234);
or U2298 (N_2298,N_2210,N_2190);
and U2299 (N_2299,N_2188,N_2244);
xnor U2300 (N_2300,N_2199,N_2179);
nand U2301 (N_2301,N_2241,N_2195);
or U2302 (N_2302,N_2245,N_2197);
and U2303 (N_2303,N_2179,N_2204);
or U2304 (N_2304,N_2192,N_2232);
nor U2305 (N_2305,N_2192,N_2183);
and U2306 (N_2306,N_2248,N_2230);
nand U2307 (N_2307,N_2202,N_2223);
nor U2308 (N_2308,N_2199,N_2234);
or U2309 (N_2309,N_2222,N_2187);
nor U2310 (N_2310,N_2204,N_2184);
or U2311 (N_2311,N_2202,N_2186);
nand U2312 (N_2312,N_2203,N_2177);
nor U2313 (N_2313,N_2193,N_2195);
and U2314 (N_2314,N_2190,N_2233);
nor U2315 (N_2315,N_2220,N_2176);
nand U2316 (N_2316,N_2229,N_2222);
nor U2317 (N_2317,N_2238,N_2234);
or U2318 (N_2318,N_2247,N_2187);
or U2319 (N_2319,N_2238,N_2219);
or U2320 (N_2320,N_2211,N_2188);
nand U2321 (N_2321,N_2232,N_2221);
or U2322 (N_2322,N_2220,N_2246);
and U2323 (N_2323,N_2230,N_2235);
nor U2324 (N_2324,N_2201,N_2221);
or U2325 (N_2325,N_2308,N_2323);
nor U2326 (N_2326,N_2306,N_2250);
nor U2327 (N_2327,N_2268,N_2321);
nor U2328 (N_2328,N_2275,N_2271);
nor U2329 (N_2329,N_2266,N_2298);
nand U2330 (N_2330,N_2292,N_2304);
or U2331 (N_2331,N_2274,N_2282);
nor U2332 (N_2332,N_2261,N_2289);
and U2333 (N_2333,N_2252,N_2318);
and U2334 (N_2334,N_2270,N_2285);
and U2335 (N_2335,N_2302,N_2257);
or U2336 (N_2336,N_2303,N_2295);
nand U2337 (N_2337,N_2259,N_2272);
and U2338 (N_2338,N_2314,N_2301);
nand U2339 (N_2339,N_2284,N_2280);
nor U2340 (N_2340,N_2273,N_2286);
xor U2341 (N_2341,N_2269,N_2283);
and U2342 (N_2342,N_2312,N_2253);
nor U2343 (N_2343,N_2294,N_2305);
or U2344 (N_2344,N_2260,N_2299);
nor U2345 (N_2345,N_2293,N_2307);
and U2346 (N_2346,N_2262,N_2324);
and U2347 (N_2347,N_2309,N_2281);
and U2348 (N_2348,N_2256,N_2290);
and U2349 (N_2349,N_2319,N_2254);
or U2350 (N_2350,N_2291,N_2300);
xnor U2351 (N_2351,N_2277,N_2276);
nand U2352 (N_2352,N_2279,N_2263);
and U2353 (N_2353,N_2317,N_2288);
and U2354 (N_2354,N_2278,N_2287);
or U2355 (N_2355,N_2265,N_2267);
nor U2356 (N_2356,N_2264,N_2322);
and U2357 (N_2357,N_2310,N_2296);
or U2358 (N_2358,N_2311,N_2258);
and U2359 (N_2359,N_2316,N_2313);
or U2360 (N_2360,N_2255,N_2320);
nor U2361 (N_2361,N_2251,N_2297);
or U2362 (N_2362,N_2315,N_2324);
or U2363 (N_2363,N_2315,N_2310);
and U2364 (N_2364,N_2300,N_2299);
nor U2365 (N_2365,N_2271,N_2258);
or U2366 (N_2366,N_2310,N_2286);
xnor U2367 (N_2367,N_2321,N_2307);
and U2368 (N_2368,N_2274,N_2322);
or U2369 (N_2369,N_2294,N_2254);
xor U2370 (N_2370,N_2268,N_2295);
and U2371 (N_2371,N_2263,N_2260);
or U2372 (N_2372,N_2258,N_2266);
nand U2373 (N_2373,N_2299,N_2264);
and U2374 (N_2374,N_2280,N_2281);
and U2375 (N_2375,N_2269,N_2263);
and U2376 (N_2376,N_2313,N_2299);
or U2377 (N_2377,N_2321,N_2279);
nor U2378 (N_2378,N_2268,N_2273);
or U2379 (N_2379,N_2282,N_2302);
or U2380 (N_2380,N_2322,N_2270);
nand U2381 (N_2381,N_2283,N_2292);
nor U2382 (N_2382,N_2288,N_2251);
and U2383 (N_2383,N_2304,N_2299);
nor U2384 (N_2384,N_2253,N_2285);
xnor U2385 (N_2385,N_2314,N_2269);
nor U2386 (N_2386,N_2292,N_2253);
and U2387 (N_2387,N_2286,N_2282);
nand U2388 (N_2388,N_2293,N_2273);
nor U2389 (N_2389,N_2306,N_2323);
or U2390 (N_2390,N_2274,N_2259);
or U2391 (N_2391,N_2294,N_2299);
nand U2392 (N_2392,N_2307,N_2309);
or U2393 (N_2393,N_2255,N_2310);
nor U2394 (N_2394,N_2296,N_2300);
nor U2395 (N_2395,N_2316,N_2257);
nand U2396 (N_2396,N_2292,N_2261);
nor U2397 (N_2397,N_2308,N_2300);
nor U2398 (N_2398,N_2286,N_2259);
nand U2399 (N_2399,N_2318,N_2277);
nor U2400 (N_2400,N_2360,N_2327);
xor U2401 (N_2401,N_2383,N_2381);
nor U2402 (N_2402,N_2391,N_2330);
nand U2403 (N_2403,N_2364,N_2348);
and U2404 (N_2404,N_2347,N_2349);
or U2405 (N_2405,N_2357,N_2336);
and U2406 (N_2406,N_2395,N_2331);
and U2407 (N_2407,N_2388,N_2394);
or U2408 (N_2408,N_2371,N_2359);
and U2409 (N_2409,N_2363,N_2328);
or U2410 (N_2410,N_2326,N_2374);
xor U2411 (N_2411,N_2385,N_2333);
nor U2412 (N_2412,N_2335,N_2355);
and U2413 (N_2413,N_2353,N_2378);
or U2414 (N_2414,N_2325,N_2373);
and U2415 (N_2415,N_2346,N_2389);
or U2416 (N_2416,N_2338,N_2356);
and U2417 (N_2417,N_2386,N_2375);
and U2418 (N_2418,N_2387,N_2368);
and U2419 (N_2419,N_2334,N_2361);
nand U2420 (N_2420,N_2365,N_2350);
or U2421 (N_2421,N_2396,N_2342);
or U2422 (N_2422,N_2392,N_2352);
nor U2423 (N_2423,N_2376,N_2398);
nand U2424 (N_2424,N_2345,N_2384);
and U2425 (N_2425,N_2351,N_2390);
nand U2426 (N_2426,N_2379,N_2332);
and U2427 (N_2427,N_2377,N_2354);
or U2428 (N_2428,N_2380,N_2369);
nor U2429 (N_2429,N_2337,N_2370);
nor U2430 (N_2430,N_2399,N_2343);
nand U2431 (N_2431,N_2382,N_2358);
nor U2432 (N_2432,N_2339,N_2341);
or U2433 (N_2433,N_2340,N_2372);
or U2434 (N_2434,N_2344,N_2366);
and U2435 (N_2435,N_2329,N_2393);
nor U2436 (N_2436,N_2362,N_2397);
or U2437 (N_2437,N_2367,N_2372);
or U2438 (N_2438,N_2391,N_2355);
and U2439 (N_2439,N_2337,N_2392);
nand U2440 (N_2440,N_2329,N_2395);
nor U2441 (N_2441,N_2371,N_2327);
or U2442 (N_2442,N_2372,N_2362);
or U2443 (N_2443,N_2342,N_2355);
or U2444 (N_2444,N_2325,N_2333);
nand U2445 (N_2445,N_2345,N_2330);
nor U2446 (N_2446,N_2368,N_2396);
nand U2447 (N_2447,N_2364,N_2386);
nor U2448 (N_2448,N_2328,N_2350);
and U2449 (N_2449,N_2384,N_2376);
and U2450 (N_2450,N_2331,N_2374);
or U2451 (N_2451,N_2394,N_2396);
or U2452 (N_2452,N_2353,N_2381);
nand U2453 (N_2453,N_2399,N_2328);
nor U2454 (N_2454,N_2361,N_2371);
nand U2455 (N_2455,N_2378,N_2350);
or U2456 (N_2456,N_2357,N_2390);
or U2457 (N_2457,N_2378,N_2392);
and U2458 (N_2458,N_2347,N_2390);
and U2459 (N_2459,N_2383,N_2361);
xor U2460 (N_2460,N_2367,N_2374);
nor U2461 (N_2461,N_2343,N_2376);
or U2462 (N_2462,N_2338,N_2357);
nand U2463 (N_2463,N_2339,N_2371);
and U2464 (N_2464,N_2329,N_2328);
or U2465 (N_2465,N_2335,N_2390);
or U2466 (N_2466,N_2345,N_2362);
nor U2467 (N_2467,N_2332,N_2361);
xnor U2468 (N_2468,N_2367,N_2351);
and U2469 (N_2469,N_2339,N_2387);
nor U2470 (N_2470,N_2376,N_2395);
nand U2471 (N_2471,N_2394,N_2352);
and U2472 (N_2472,N_2338,N_2375);
and U2473 (N_2473,N_2388,N_2367);
nor U2474 (N_2474,N_2339,N_2393);
nor U2475 (N_2475,N_2432,N_2418);
nand U2476 (N_2476,N_2433,N_2411);
or U2477 (N_2477,N_2400,N_2435);
xor U2478 (N_2478,N_2417,N_2463);
and U2479 (N_2479,N_2462,N_2472);
and U2480 (N_2480,N_2402,N_2446);
nand U2481 (N_2481,N_2447,N_2403);
nand U2482 (N_2482,N_2427,N_2467);
nor U2483 (N_2483,N_2459,N_2468);
and U2484 (N_2484,N_2466,N_2470);
nand U2485 (N_2485,N_2428,N_2449);
nand U2486 (N_2486,N_2423,N_2457);
nor U2487 (N_2487,N_2421,N_2408);
nor U2488 (N_2488,N_2420,N_2437);
nand U2489 (N_2489,N_2406,N_2419);
and U2490 (N_2490,N_2453,N_2443);
nand U2491 (N_2491,N_2473,N_2426);
nor U2492 (N_2492,N_2405,N_2458);
and U2493 (N_2493,N_2456,N_2461);
or U2494 (N_2494,N_2425,N_2431);
and U2495 (N_2495,N_2407,N_2450);
nor U2496 (N_2496,N_2430,N_2444);
nand U2497 (N_2497,N_2404,N_2464);
or U2498 (N_2498,N_2416,N_2414);
nor U2499 (N_2499,N_2441,N_2410);
and U2500 (N_2500,N_2474,N_2412);
or U2501 (N_2501,N_2413,N_2429);
and U2502 (N_2502,N_2454,N_2451);
and U2503 (N_2503,N_2448,N_2445);
nand U2504 (N_2504,N_2424,N_2439);
and U2505 (N_2505,N_2409,N_2442);
nand U2506 (N_2506,N_2455,N_2401);
nand U2507 (N_2507,N_2438,N_2440);
and U2508 (N_2508,N_2434,N_2415);
nor U2509 (N_2509,N_2469,N_2436);
nor U2510 (N_2510,N_2471,N_2422);
nand U2511 (N_2511,N_2460,N_2465);
nor U2512 (N_2512,N_2452,N_2441);
nor U2513 (N_2513,N_2411,N_2473);
or U2514 (N_2514,N_2462,N_2415);
or U2515 (N_2515,N_2412,N_2432);
or U2516 (N_2516,N_2428,N_2452);
or U2517 (N_2517,N_2404,N_2405);
or U2518 (N_2518,N_2432,N_2427);
or U2519 (N_2519,N_2452,N_2422);
nor U2520 (N_2520,N_2467,N_2408);
nor U2521 (N_2521,N_2424,N_2419);
xor U2522 (N_2522,N_2404,N_2455);
or U2523 (N_2523,N_2464,N_2456);
nand U2524 (N_2524,N_2468,N_2460);
nand U2525 (N_2525,N_2431,N_2455);
or U2526 (N_2526,N_2459,N_2408);
and U2527 (N_2527,N_2414,N_2447);
nand U2528 (N_2528,N_2417,N_2410);
or U2529 (N_2529,N_2427,N_2457);
nor U2530 (N_2530,N_2445,N_2463);
nand U2531 (N_2531,N_2441,N_2466);
xnor U2532 (N_2532,N_2474,N_2415);
and U2533 (N_2533,N_2407,N_2472);
and U2534 (N_2534,N_2451,N_2431);
and U2535 (N_2535,N_2406,N_2450);
nand U2536 (N_2536,N_2418,N_2408);
nand U2537 (N_2537,N_2410,N_2464);
or U2538 (N_2538,N_2441,N_2414);
or U2539 (N_2539,N_2437,N_2459);
and U2540 (N_2540,N_2425,N_2454);
nand U2541 (N_2541,N_2402,N_2412);
nand U2542 (N_2542,N_2431,N_2405);
nand U2543 (N_2543,N_2409,N_2403);
nor U2544 (N_2544,N_2424,N_2415);
nand U2545 (N_2545,N_2413,N_2453);
and U2546 (N_2546,N_2446,N_2428);
xor U2547 (N_2547,N_2410,N_2467);
or U2548 (N_2548,N_2419,N_2463);
nor U2549 (N_2549,N_2444,N_2470);
nand U2550 (N_2550,N_2477,N_2503);
xor U2551 (N_2551,N_2506,N_2479);
or U2552 (N_2552,N_2507,N_2548);
nor U2553 (N_2553,N_2516,N_2523);
or U2554 (N_2554,N_2549,N_2476);
nor U2555 (N_2555,N_2545,N_2484);
and U2556 (N_2556,N_2527,N_2495);
or U2557 (N_2557,N_2522,N_2520);
nor U2558 (N_2558,N_2499,N_2490);
and U2559 (N_2559,N_2518,N_2525);
or U2560 (N_2560,N_2493,N_2538);
or U2561 (N_2561,N_2486,N_2514);
and U2562 (N_2562,N_2504,N_2539);
or U2563 (N_2563,N_2531,N_2512);
or U2564 (N_2564,N_2480,N_2536);
nor U2565 (N_2565,N_2491,N_2540);
nand U2566 (N_2566,N_2488,N_2482);
or U2567 (N_2567,N_2481,N_2485);
nand U2568 (N_2568,N_2489,N_2509);
or U2569 (N_2569,N_2494,N_2534);
nand U2570 (N_2570,N_2524,N_2501);
or U2571 (N_2571,N_2502,N_2505);
xor U2572 (N_2572,N_2483,N_2535);
or U2573 (N_2573,N_2475,N_2498);
or U2574 (N_2574,N_2541,N_2546);
or U2575 (N_2575,N_2497,N_2526);
or U2576 (N_2576,N_2515,N_2492);
and U2577 (N_2577,N_2487,N_2533);
or U2578 (N_2578,N_2544,N_2542);
and U2579 (N_2579,N_2521,N_2478);
nor U2580 (N_2580,N_2517,N_2530);
and U2581 (N_2581,N_2510,N_2532);
or U2582 (N_2582,N_2519,N_2537);
or U2583 (N_2583,N_2496,N_2508);
or U2584 (N_2584,N_2500,N_2547);
and U2585 (N_2585,N_2529,N_2511);
nand U2586 (N_2586,N_2528,N_2543);
nor U2587 (N_2587,N_2513,N_2514);
nand U2588 (N_2588,N_2537,N_2544);
nor U2589 (N_2589,N_2544,N_2539);
nand U2590 (N_2590,N_2541,N_2549);
nand U2591 (N_2591,N_2516,N_2548);
nand U2592 (N_2592,N_2514,N_2485);
nand U2593 (N_2593,N_2542,N_2545);
or U2594 (N_2594,N_2519,N_2548);
xor U2595 (N_2595,N_2486,N_2484);
nor U2596 (N_2596,N_2538,N_2479);
nand U2597 (N_2597,N_2538,N_2502);
nand U2598 (N_2598,N_2521,N_2515);
nand U2599 (N_2599,N_2504,N_2513);
nand U2600 (N_2600,N_2495,N_2512);
nand U2601 (N_2601,N_2499,N_2486);
xor U2602 (N_2602,N_2548,N_2538);
nand U2603 (N_2603,N_2518,N_2513);
or U2604 (N_2604,N_2537,N_2491);
nand U2605 (N_2605,N_2503,N_2495);
or U2606 (N_2606,N_2481,N_2515);
nand U2607 (N_2607,N_2498,N_2503);
or U2608 (N_2608,N_2543,N_2539);
and U2609 (N_2609,N_2489,N_2495);
or U2610 (N_2610,N_2487,N_2505);
nand U2611 (N_2611,N_2491,N_2489);
xor U2612 (N_2612,N_2546,N_2527);
nor U2613 (N_2613,N_2492,N_2523);
or U2614 (N_2614,N_2546,N_2523);
nand U2615 (N_2615,N_2505,N_2535);
nand U2616 (N_2616,N_2499,N_2514);
and U2617 (N_2617,N_2479,N_2533);
nand U2618 (N_2618,N_2523,N_2482);
and U2619 (N_2619,N_2490,N_2511);
or U2620 (N_2620,N_2526,N_2505);
nor U2621 (N_2621,N_2523,N_2529);
nand U2622 (N_2622,N_2539,N_2546);
nor U2623 (N_2623,N_2535,N_2518);
or U2624 (N_2624,N_2515,N_2544);
nor U2625 (N_2625,N_2610,N_2565);
nor U2626 (N_2626,N_2614,N_2580);
nor U2627 (N_2627,N_2597,N_2620);
nand U2628 (N_2628,N_2588,N_2550);
and U2629 (N_2629,N_2582,N_2605);
nand U2630 (N_2630,N_2572,N_2585);
and U2631 (N_2631,N_2554,N_2556);
nand U2632 (N_2632,N_2553,N_2579);
nand U2633 (N_2633,N_2559,N_2573);
nor U2634 (N_2634,N_2608,N_2566);
nand U2635 (N_2635,N_2593,N_2619);
nor U2636 (N_2636,N_2618,N_2551);
nand U2637 (N_2637,N_2595,N_2599);
nand U2638 (N_2638,N_2584,N_2570);
nand U2639 (N_2639,N_2586,N_2623);
nor U2640 (N_2640,N_2594,N_2576);
or U2641 (N_2641,N_2613,N_2592);
nor U2642 (N_2642,N_2589,N_2606);
or U2643 (N_2643,N_2555,N_2596);
and U2644 (N_2644,N_2564,N_2604);
nor U2645 (N_2645,N_2601,N_2558);
or U2646 (N_2646,N_2607,N_2574);
or U2647 (N_2647,N_2581,N_2571);
or U2648 (N_2648,N_2609,N_2563);
nor U2649 (N_2649,N_2568,N_2611);
nor U2650 (N_2650,N_2612,N_2615);
nor U2651 (N_2651,N_2587,N_2600);
or U2652 (N_2652,N_2598,N_2603);
and U2653 (N_2653,N_2561,N_2569);
nand U2654 (N_2654,N_2621,N_2575);
nor U2655 (N_2655,N_2616,N_2617);
nand U2656 (N_2656,N_2552,N_2560);
nand U2657 (N_2657,N_2622,N_2562);
and U2658 (N_2658,N_2602,N_2591);
or U2659 (N_2659,N_2578,N_2567);
nor U2660 (N_2660,N_2577,N_2583);
nor U2661 (N_2661,N_2624,N_2557);
or U2662 (N_2662,N_2590,N_2565);
nand U2663 (N_2663,N_2603,N_2612);
or U2664 (N_2664,N_2562,N_2587);
or U2665 (N_2665,N_2592,N_2599);
nand U2666 (N_2666,N_2563,N_2603);
or U2667 (N_2667,N_2562,N_2601);
or U2668 (N_2668,N_2620,N_2568);
or U2669 (N_2669,N_2556,N_2578);
nand U2670 (N_2670,N_2585,N_2607);
nand U2671 (N_2671,N_2595,N_2590);
nor U2672 (N_2672,N_2573,N_2564);
and U2673 (N_2673,N_2589,N_2579);
and U2674 (N_2674,N_2596,N_2567);
nor U2675 (N_2675,N_2556,N_2621);
nor U2676 (N_2676,N_2623,N_2621);
and U2677 (N_2677,N_2619,N_2570);
or U2678 (N_2678,N_2592,N_2572);
or U2679 (N_2679,N_2560,N_2585);
nor U2680 (N_2680,N_2580,N_2605);
and U2681 (N_2681,N_2603,N_2579);
or U2682 (N_2682,N_2586,N_2577);
nand U2683 (N_2683,N_2550,N_2590);
and U2684 (N_2684,N_2604,N_2594);
nor U2685 (N_2685,N_2573,N_2616);
nor U2686 (N_2686,N_2584,N_2596);
or U2687 (N_2687,N_2608,N_2612);
or U2688 (N_2688,N_2553,N_2596);
nand U2689 (N_2689,N_2593,N_2618);
nor U2690 (N_2690,N_2618,N_2579);
and U2691 (N_2691,N_2552,N_2563);
or U2692 (N_2692,N_2582,N_2559);
or U2693 (N_2693,N_2590,N_2618);
nor U2694 (N_2694,N_2609,N_2564);
or U2695 (N_2695,N_2575,N_2572);
or U2696 (N_2696,N_2616,N_2552);
and U2697 (N_2697,N_2576,N_2613);
nand U2698 (N_2698,N_2556,N_2602);
nor U2699 (N_2699,N_2607,N_2603);
or U2700 (N_2700,N_2695,N_2639);
xnor U2701 (N_2701,N_2657,N_2684);
nor U2702 (N_2702,N_2685,N_2689);
nor U2703 (N_2703,N_2654,N_2682);
nand U2704 (N_2704,N_2688,N_2660);
and U2705 (N_2705,N_2636,N_2647);
nor U2706 (N_2706,N_2696,N_2662);
or U2707 (N_2707,N_2648,N_2632);
nor U2708 (N_2708,N_2659,N_2631);
nand U2709 (N_2709,N_2675,N_2645);
or U2710 (N_2710,N_2633,N_2690);
nor U2711 (N_2711,N_2669,N_2678);
nor U2712 (N_2712,N_2634,N_2693);
nor U2713 (N_2713,N_2638,N_2651);
or U2714 (N_2714,N_2666,N_2627);
nand U2715 (N_2715,N_2642,N_2650);
and U2716 (N_2716,N_2630,N_2667);
nor U2717 (N_2717,N_2644,N_2683);
nand U2718 (N_2718,N_2656,N_2671);
and U2719 (N_2719,N_2672,N_2635);
and U2720 (N_2720,N_2692,N_2646);
and U2721 (N_2721,N_2643,N_2680);
and U2722 (N_2722,N_2641,N_2629);
or U2723 (N_2723,N_2686,N_2670);
nand U2724 (N_2724,N_2698,N_2677);
nand U2725 (N_2725,N_2679,N_2668);
and U2726 (N_2726,N_2661,N_2653);
xor U2727 (N_2727,N_2681,N_2625);
or U2728 (N_2728,N_2655,N_2626);
and U2729 (N_2729,N_2699,N_2676);
or U2730 (N_2730,N_2637,N_2652);
and U2731 (N_2731,N_2628,N_2665);
and U2732 (N_2732,N_2658,N_2640);
or U2733 (N_2733,N_2694,N_2674);
and U2734 (N_2734,N_2663,N_2673);
and U2735 (N_2735,N_2687,N_2664);
nor U2736 (N_2736,N_2697,N_2649);
nor U2737 (N_2737,N_2691,N_2657);
and U2738 (N_2738,N_2686,N_2669);
nor U2739 (N_2739,N_2673,N_2626);
nand U2740 (N_2740,N_2654,N_2643);
or U2741 (N_2741,N_2648,N_2638);
nand U2742 (N_2742,N_2683,N_2632);
and U2743 (N_2743,N_2660,N_2636);
nand U2744 (N_2744,N_2692,N_2639);
nand U2745 (N_2745,N_2684,N_2627);
nand U2746 (N_2746,N_2695,N_2652);
and U2747 (N_2747,N_2637,N_2628);
nand U2748 (N_2748,N_2686,N_2641);
nand U2749 (N_2749,N_2672,N_2657);
and U2750 (N_2750,N_2666,N_2658);
or U2751 (N_2751,N_2642,N_2648);
nor U2752 (N_2752,N_2656,N_2657);
nand U2753 (N_2753,N_2699,N_2656);
or U2754 (N_2754,N_2669,N_2653);
nand U2755 (N_2755,N_2688,N_2689);
and U2756 (N_2756,N_2661,N_2696);
and U2757 (N_2757,N_2682,N_2689);
nand U2758 (N_2758,N_2666,N_2667);
nor U2759 (N_2759,N_2675,N_2643);
nor U2760 (N_2760,N_2662,N_2680);
or U2761 (N_2761,N_2666,N_2635);
and U2762 (N_2762,N_2653,N_2658);
nand U2763 (N_2763,N_2691,N_2675);
nand U2764 (N_2764,N_2625,N_2637);
nand U2765 (N_2765,N_2653,N_2680);
nand U2766 (N_2766,N_2687,N_2684);
and U2767 (N_2767,N_2697,N_2694);
nand U2768 (N_2768,N_2672,N_2692);
nand U2769 (N_2769,N_2656,N_2665);
and U2770 (N_2770,N_2666,N_2638);
nand U2771 (N_2771,N_2629,N_2697);
and U2772 (N_2772,N_2679,N_2662);
or U2773 (N_2773,N_2630,N_2660);
and U2774 (N_2774,N_2627,N_2642);
nor U2775 (N_2775,N_2729,N_2764);
nor U2776 (N_2776,N_2744,N_2716);
or U2777 (N_2777,N_2703,N_2736);
and U2778 (N_2778,N_2771,N_2733);
nand U2779 (N_2779,N_2741,N_2728);
and U2780 (N_2780,N_2760,N_2700);
or U2781 (N_2781,N_2737,N_2718);
nand U2782 (N_2782,N_2767,N_2758);
or U2783 (N_2783,N_2756,N_2732);
nor U2784 (N_2784,N_2754,N_2711);
or U2785 (N_2785,N_2724,N_2740);
and U2786 (N_2786,N_2735,N_2713);
or U2787 (N_2787,N_2725,N_2739);
and U2788 (N_2788,N_2723,N_2706);
and U2789 (N_2789,N_2730,N_2768);
nand U2790 (N_2790,N_2747,N_2721);
or U2791 (N_2791,N_2770,N_2773);
nand U2792 (N_2792,N_2742,N_2757);
nand U2793 (N_2793,N_2769,N_2748);
nor U2794 (N_2794,N_2704,N_2714);
nand U2795 (N_2795,N_2749,N_2755);
nand U2796 (N_2796,N_2772,N_2745);
and U2797 (N_2797,N_2762,N_2726);
or U2798 (N_2798,N_2710,N_2722);
nor U2799 (N_2799,N_2705,N_2750);
or U2800 (N_2800,N_2746,N_2719);
nor U2801 (N_2801,N_2774,N_2727);
nor U2802 (N_2802,N_2765,N_2752);
or U2803 (N_2803,N_2717,N_2734);
nor U2804 (N_2804,N_2761,N_2701);
and U2805 (N_2805,N_2759,N_2738);
and U2806 (N_2806,N_2709,N_2743);
or U2807 (N_2807,N_2751,N_2731);
nand U2808 (N_2808,N_2707,N_2766);
or U2809 (N_2809,N_2712,N_2702);
nand U2810 (N_2810,N_2720,N_2763);
nor U2811 (N_2811,N_2753,N_2715);
and U2812 (N_2812,N_2708,N_2719);
nand U2813 (N_2813,N_2769,N_2738);
nor U2814 (N_2814,N_2768,N_2717);
nand U2815 (N_2815,N_2747,N_2751);
and U2816 (N_2816,N_2714,N_2764);
nor U2817 (N_2817,N_2753,N_2734);
nor U2818 (N_2818,N_2703,N_2774);
nor U2819 (N_2819,N_2736,N_2705);
and U2820 (N_2820,N_2720,N_2765);
nand U2821 (N_2821,N_2754,N_2744);
or U2822 (N_2822,N_2757,N_2700);
or U2823 (N_2823,N_2753,N_2774);
nor U2824 (N_2824,N_2761,N_2770);
and U2825 (N_2825,N_2732,N_2738);
nor U2826 (N_2826,N_2715,N_2772);
or U2827 (N_2827,N_2757,N_2721);
and U2828 (N_2828,N_2757,N_2735);
and U2829 (N_2829,N_2729,N_2772);
nor U2830 (N_2830,N_2722,N_2711);
and U2831 (N_2831,N_2721,N_2711);
nor U2832 (N_2832,N_2760,N_2732);
nor U2833 (N_2833,N_2716,N_2714);
nor U2834 (N_2834,N_2757,N_2726);
or U2835 (N_2835,N_2733,N_2752);
nand U2836 (N_2836,N_2728,N_2738);
nor U2837 (N_2837,N_2759,N_2760);
or U2838 (N_2838,N_2732,N_2703);
nand U2839 (N_2839,N_2774,N_2754);
nor U2840 (N_2840,N_2751,N_2773);
nand U2841 (N_2841,N_2702,N_2746);
and U2842 (N_2842,N_2752,N_2762);
nand U2843 (N_2843,N_2726,N_2760);
nand U2844 (N_2844,N_2753,N_2704);
nand U2845 (N_2845,N_2716,N_2772);
nand U2846 (N_2846,N_2700,N_2734);
and U2847 (N_2847,N_2756,N_2724);
and U2848 (N_2848,N_2743,N_2732);
or U2849 (N_2849,N_2760,N_2749);
nor U2850 (N_2850,N_2842,N_2844);
nor U2851 (N_2851,N_2783,N_2817);
nor U2852 (N_2852,N_2799,N_2775);
and U2853 (N_2853,N_2818,N_2848);
nand U2854 (N_2854,N_2789,N_2802);
nand U2855 (N_2855,N_2795,N_2806);
nor U2856 (N_2856,N_2837,N_2815);
and U2857 (N_2857,N_2822,N_2788);
and U2858 (N_2858,N_2781,N_2846);
xor U2859 (N_2859,N_2840,N_2841);
or U2860 (N_2860,N_2827,N_2787);
nor U2861 (N_2861,N_2819,N_2839);
and U2862 (N_2862,N_2830,N_2812);
nand U2863 (N_2863,N_2821,N_2790);
or U2864 (N_2864,N_2829,N_2780);
or U2865 (N_2865,N_2798,N_2800);
or U2866 (N_2866,N_2823,N_2814);
nand U2867 (N_2867,N_2847,N_2793);
nor U2868 (N_2868,N_2792,N_2838);
nand U2869 (N_2869,N_2796,N_2834);
nor U2870 (N_2870,N_2832,N_2797);
or U2871 (N_2871,N_2805,N_2843);
nand U2872 (N_2872,N_2777,N_2779);
or U2873 (N_2873,N_2824,N_2791);
and U2874 (N_2874,N_2826,N_2782);
nand U2875 (N_2875,N_2784,N_2825);
and U2876 (N_2876,N_2833,N_2801);
nand U2877 (N_2877,N_2820,N_2776);
or U2878 (N_2878,N_2849,N_2811);
and U2879 (N_2879,N_2803,N_2778);
nor U2880 (N_2880,N_2836,N_2809);
nor U2881 (N_2881,N_2831,N_2785);
and U2882 (N_2882,N_2813,N_2810);
and U2883 (N_2883,N_2845,N_2807);
nor U2884 (N_2884,N_2808,N_2804);
nor U2885 (N_2885,N_2786,N_2794);
or U2886 (N_2886,N_2816,N_2835);
or U2887 (N_2887,N_2828,N_2817);
nand U2888 (N_2888,N_2789,N_2812);
nor U2889 (N_2889,N_2819,N_2789);
or U2890 (N_2890,N_2836,N_2823);
or U2891 (N_2891,N_2810,N_2812);
xnor U2892 (N_2892,N_2780,N_2818);
or U2893 (N_2893,N_2849,N_2807);
and U2894 (N_2894,N_2804,N_2782);
or U2895 (N_2895,N_2832,N_2778);
nand U2896 (N_2896,N_2797,N_2802);
or U2897 (N_2897,N_2840,N_2809);
and U2898 (N_2898,N_2794,N_2833);
nor U2899 (N_2899,N_2832,N_2804);
or U2900 (N_2900,N_2813,N_2822);
or U2901 (N_2901,N_2839,N_2796);
nor U2902 (N_2902,N_2784,N_2785);
or U2903 (N_2903,N_2778,N_2825);
nor U2904 (N_2904,N_2845,N_2835);
and U2905 (N_2905,N_2780,N_2801);
nand U2906 (N_2906,N_2779,N_2788);
or U2907 (N_2907,N_2826,N_2811);
nor U2908 (N_2908,N_2800,N_2847);
and U2909 (N_2909,N_2845,N_2797);
nor U2910 (N_2910,N_2781,N_2811);
or U2911 (N_2911,N_2816,N_2784);
nand U2912 (N_2912,N_2840,N_2806);
nor U2913 (N_2913,N_2834,N_2781);
and U2914 (N_2914,N_2788,N_2833);
xnor U2915 (N_2915,N_2821,N_2824);
nor U2916 (N_2916,N_2835,N_2817);
and U2917 (N_2917,N_2794,N_2817);
and U2918 (N_2918,N_2838,N_2810);
or U2919 (N_2919,N_2833,N_2839);
nor U2920 (N_2920,N_2826,N_2787);
or U2921 (N_2921,N_2817,N_2844);
nor U2922 (N_2922,N_2786,N_2835);
xor U2923 (N_2923,N_2845,N_2832);
or U2924 (N_2924,N_2818,N_2788);
nand U2925 (N_2925,N_2905,N_2869);
and U2926 (N_2926,N_2858,N_2914);
and U2927 (N_2927,N_2879,N_2921);
and U2928 (N_2928,N_2865,N_2911);
nor U2929 (N_2929,N_2864,N_2877);
or U2930 (N_2930,N_2918,N_2886);
and U2931 (N_2931,N_2902,N_2907);
nor U2932 (N_2932,N_2900,N_2919);
nand U2933 (N_2933,N_2894,N_2880);
or U2934 (N_2934,N_2891,N_2870);
xor U2935 (N_2935,N_2873,N_2883);
and U2936 (N_2936,N_2857,N_2860);
nand U2937 (N_2937,N_2874,N_2917);
nor U2938 (N_2938,N_2901,N_2904);
nor U2939 (N_2939,N_2872,N_2884);
nand U2940 (N_2940,N_2915,N_2855);
or U2941 (N_2941,N_2892,N_2912);
and U2942 (N_2942,N_2896,N_2888);
nand U2943 (N_2943,N_2908,N_2887);
nand U2944 (N_2944,N_2889,N_2854);
nand U2945 (N_2945,N_2895,N_2890);
or U2946 (N_2946,N_2878,N_2871);
and U2947 (N_2947,N_2906,N_2923);
nor U2948 (N_2948,N_2851,N_2853);
nor U2949 (N_2949,N_2910,N_2867);
nand U2950 (N_2950,N_2861,N_2859);
or U2951 (N_2951,N_2898,N_2881);
xnor U2952 (N_2952,N_2899,N_2893);
or U2953 (N_2953,N_2862,N_2903);
nand U2954 (N_2954,N_2850,N_2885);
nand U2955 (N_2955,N_2882,N_2866);
or U2956 (N_2956,N_2922,N_2852);
and U2957 (N_2957,N_2920,N_2909);
or U2958 (N_2958,N_2863,N_2924);
and U2959 (N_2959,N_2856,N_2868);
nand U2960 (N_2960,N_2913,N_2897);
nor U2961 (N_2961,N_2875,N_2876);
nand U2962 (N_2962,N_2916,N_2919);
nor U2963 (N_2963,N_2917,N_2899);
or U2964 (N_2964,N_2891,N_2911);
nor U2965 (N_2965,N_2851,N_2889);
nor U2966 (N_2966,N_2885,N_2857);
nor U2967 (N_2967,N_2900,N_2865);
and U2968 (N_2968,N_2852,N_2853);
and U2969 (N_2969,N_2869,N_2913);
nand U2970 (N_2970,N_2870,N_2851);
nand U2971 (N_2971,N_2883,N_2908);
and U2972 (N_2972,N_2868,N_2881);
nand U2973 (N_2973,N_2859,N_2912);
nor U2974 (N_2974,N_2897,N_2900);
nor U2975 (N_2975,N_2915,N_2879);
xnor U2976 (N_2976,N_2919,N_2878);
or U2977 (N_2977,N_2856,N_2901);
nor U2978 (N_2978,N_2877,N_2862);
or U2979 (N_2979,N_2855,N_2913);
nand U2980 (N_2980,N_2867,N_2866);
nor U2981 (N_2981,N_2905,N_2912);
nand U2982 (N_2982,N_2874,N_2918);
nor U2983 (N_2983,N_2912,N_2852);
nand U2984 (N_2984,N_2853,N_2874);
or U2985 (N_2985,N_2913,N_2922);
nor U2986 (N_2986,N_2911,N_2875);
nand U2987 (N_2987,N_2852,N_2896);
nand U2988 (N_2988,N_2923,N_2920);
nor U2989 (N_2989,N_2882,N_2854);
nor U2990 (N_2990,N_2922,N_2910);
nand U2991 (N_2991,N_2858,N_2884);
or U2992 (N_2992,N_2886,N_2856);
or U2993 (N_2993,N_2914,N_2880);
nor U2994 (N_2994,N_2869,N_2862);
or U2995 (N_2995,N_2898,N_2872);
and U2996 (N_2996,N_2923,N_2903);
nand U2997 (N_2997,N_2904,N_2915);
nand U2998 (N_2998,N_2894,N_2923);
nor U2999 (N_2999,N_2867,N_2872);
xnor UO_0 (O_0,N_2953,N_2929);
nand UO_1 (O_1,N_2927,N_2984);
and UO_2 (O_2,N_2958,N_2976);
or UO_3 (O_3,N_2999,N_2972);
and UO_4 (O_4,N_2943,N_2963);
and UO_5 (O_5,N_2950,N_2995);
nor UO_6 (O_6,N_2945,N_2966);
or UO_7 (O_7,N_2987,N_2964);
nand UO_8 (O_8,N_2982,N_2959);
or UO_9 (O_9,N_2969,N_2944);
nand UO_10 (O_10,N_2938,N_2989);
and UO_11 (O_11,N_2983,N_2998);
and UO_12 (O_12,N_2956,N_2992);
and UO_13 (O_13,N_2947,N_2937);
and UO_14 (O_14,N_2961,N_2939);
nor UO_15 (O_15,N_2941,N_2936);
nand UO_16 (O_16,N_2968,N_2942);
nor UO_17 (O_17,N_2954,N_2971);
and UO_18 (O_18,N_2928,N_2948);
nand UO_19 (O_19,N_2974,N_2946);
or UO_20 (O_20,N_2970,N_2933);
or UO_21 (O_21,N_2997,N_2977);
or UO_22 (O_22,N_2962,N_2930);
nand UO_23 (O_23,N_2965,N_2981);
nand UO_24 (O_24,N_2949,N_2973);
and UO_25 (O_25,N_2957,N_2975);
and UO_26 (O_26,N_2985,N_2935);
or UO_27 (O_27,N_2990,N_2993);
nand UO_28 (O_28,N_2978,N_2952);
nand UO_29 (O_29,N_2996,N_2988);
or UO_30 (O_30,N_2994,N_2940);
nand UO_31 (O_31,N_2931,N_2925);
and UO_32 (O_32,N_2967,N_2979);
and UO_33 (O_33,N_2951,N_2980);
nand UO_34 (O_34,N_2991,N_2934);
nor UO_35 (O_35,N_2955,N_2926);
nand UO_36 (O_36,N_2986,N_2960);
and UO_37 (O_37,N_2932,N_2952);
or UO_38 (O_38,N_2997,N_2973);
nor UO_39 (O_39,N_2925,N_2934);
and UO_40 (O_40,N_2960,N_2991);
nor UO_41 (O_41,N_2975,N_2989);
nand UO_42 (O_42,N_2983,N_2929);
nor UO_43 (O_43,N_2958,N_2943);
and UO_44 (O_44,N_2953,N_2928);
and UO_45 (O_45,N_2965,N_2951);
nor UO_46 (O_46,N_2972,N_2993);
nand UO_47 (O_47,N_2927,N_2950);
or UO_48 (O_48,N_2926,N_2960);
nand UO_49 (O_49,N_2951,N_2933);
nor UO_50 (O_50,N_2933,N_2946);
and UO_51 (O_51,N_2931,N_2936);
nand UO_52 (O_52,N_2987,N_2946);
and UO_53 (O_53,N_2977,N_2933);
nor UO_54 (O_54,N_2948,N_2962);
and UO_55 (O_55,N_2930,N_2956);
or UO_56 (O_56,N_2960,N_2944);
or UO_57 (O_57,N_2998,N_2994);
and UO_58 (O_58,N_2949,N_2947);
or UO_59 (O_59,N_2993,N_2958);
nor UO_60 (O_60,N_2993,N_2970);
and UO_61 (O_61,N_2976,N_2959);
or UO_62 (O_62,N_2932,N_2931);
and UO_63 (O_63,N_2994,N_2985);
nor UO_64 (O_64,N_2974,N_2972);
nand UO_65 (O_65,N_2988,N_2941);
nor UO_66 (O_66,N_2929,N_2932);
nand UO_67 (O_67,N_2929,N_2967);
xnor UO_68 (O_68,N_2936,N_2986);
nor UO_69 (O_69,N_2974,N_2986);
and UO_70 (O_70,N_2992,N_2944);
or UO_71 (O_71,N_2993,N_2945);
nand UO_72 (O_72,N_2943,N_2933);
nand UO_73 (O_73,N_2962,N_2932);
nor UO_74 (O_74,N_2925,N_2969);
nor UO_75 (O_75,N_2952,N_2984);
or UO_76 (O_76,N_2958,N_2929);
nor UO_77 (O_77,N_2981,N_2986);
nand UO_78 (O_78,N_2928,N_2985);
and UO_79 (O_79,N_2941,N_2965);
nor UO_80 (O_80,N_2931,N_2959);
nand UO_81 (O_81,N_2940,N_2927);
or UO_82 (O_82,N_2991,N_2949);
and UO_83 (O_83,N_2963,N_2945);
or UO_84 (O_84,N_2942,N_2993);
and UO_85 (O_85,N_2972,N_2942);
or UO_86 (O_86,N_2944,N_2981);
nor UO_87 (O_87,N_2931,N_2994);
and UO_88 (O_88,N_2965,N_2979);
nor UO_89 (O_89,N_2989,N_2985);
and UO_90 (O_90,N_2990,N_2974);
or UO_91 (O_91,N_2970,N_2937);
and UO_92 (O_92,N_2951,N_2942);
or UO_93 (O_93,N_2981,N_2991);
and UO_94 (O_94,N_2944,N_2926);
or UO_95 (O_95,N_2957,N_2946);
and UO_96 (O_96,N_2947,N_2971);
or UO_97 (O_97,N_2986,N_2983);
nand UO_98 (O_98,N_2999,N_2969);
nor UO_99 (O_99,N_2927,N_2928);
and UO_100 (O_100,N_2993,N_2977);
nand UO_101 (O_101,N_2980,N_2927);
nor UO_102 (O_102,N_2925,N_2996);
and UO_103 (O_103,N_2950,N_2980);
nand UO_104 (O_104,N_2994,N_2949);
or UO_105 (O_105,N_2925,N_2994);
nand UO_106 (O_106,N_2987,N_2932);
or UO_107 (O_107,N_2993,N_2935);
or UO_108 (O_108,N_2925,N_2959);
and UO_109 (O_109,N_2982,N_2936);
nand UO_110 (O_110,N_2996,N_2964);
or UO_111 (O_111,N_2987,N_2951);
or UO_112 (O_112,N_2935,N_2943);
and UO_113 (O_113,N_2935,N_2930);
nor UO_114 (O_114,N_2932,N_2978);
nor UO_115 (O_115,N_2931,N_2960);
and UO_116 (O_116,N_2928,N_2960);
or UO_117 (O_117,N_2975,N_2985);
nand UO_118 (O_118,N_2954,N_2935);
and UO_119 (O_119,N_2959,N_2970);
xor UO_120 (O_120,N_2965,N_2994);
nand UO_121 (O_121,N_2986,N_2969);
nand UO_122 (O_122,N_2987,N_2939);
nand UO_123 (O_123,N_2960,N_2953);
nand UO_124 (O_124,N_2929,N_2972);
nand UO_125 (O_125,N_2935,N_2970);
or UO_126 (O_126,N_2997,N_2955);
and UO_127 (O_127,N_2963,N_2964);
nand UO_128 (O_128,N_2970,N_2952);
nand UO_129 (O_129,N_2961,N_2929);
or UO_130 (O_130,N_2930,N_2992);
nor UO_131 (O_131,N_2970,N_2941);
nand UO_132 (O_132,N_2932,N_2992);
nor UO_133 (O_133,N_2929,N_2947);
nor UO_134 (O_134,N_2975,N_2987);
nand UO_135 (O_135,N_2969,N_2982);
or UO_136 (O_136,N_2967,N_2946);
nor UO_137 (O_137,N_2988,N_2943);
and UO_138 (O_138,N_2926,N_2932);
and UO_139 (O_139,N_2979,N_2990);
nand UO_140 (O_140,N_2969,N_2991);
or UO_141 (O_141,N_2941,N_2942);
or UO_142 (O_142,N_2970,N_2929);
or UO_143 (O_143,N_2940,N_2955);
nor UO_144 (O_144,N_2988,N_2951);
nor UO_145 (O_145,N_2982,N_2940);
and UO_146 (O_146,N_2947,N_2973);
nor UO_147 (O_147,N_2940,N_2959);
nand UO_148 (O_148,N_2985,N_2984);
and UO_149 (O_149,N_2990,N_2932);
nor UO_150 (O_150,N_2936,N_2961);
or UO_151 (O_151,N_2930,N_2987);
nor UO_152 (O_152,N_2960,N_2967);
and UO_153 (O_153,N_2949,N_2959);
and UO_154 (O_154,N_2927,N_2968);
and UO_155 (O_155,N_2965,N_2974);
or UO_156 (O_156,N_2928,N_2979);
nand UO_157 (O_157,N_2947,N_2988);
and UO_158 (O_158,N_2930,N_2970);
nor UO_159 (O_159,N_2970,N_2954);
and UO_160 (O_160,N_2994,N_2941);
nor UO_161 (O_161,N_2980,N_2959);
nor UO_162 (O_162,N_2970,N_2951);
and UO_163 (O_163,N_2985,N_2953);
and UO_164 (O_164,N_2975,N_2935);
or UO_165 (O_165,N_2952,N_2957);
or UO_166 (O_166,N_2980,N_2945);
nor UO_167 (O_167,N_2937,N_2964);
nand UO_168 (O_168,N_2949,N_2985);
and UO_169 (O_169,N_2931,N_2927);
and UO_170 (O_170,N_2961,N_2960);
or UO_171 (O_171,N_2941,N_2939);
or UO_172 (O_172,N_2939,N_2975);
and UO_173 (O_173,N_2926,N_2987);
or UO_174 (O_174,N_2993,N_2980);
nor UO_175 (O_175,N_2984,N_2925);
nor UO_176 (O_176,N_2957,N_2992);
nor UO_177 (O_177,N_2990,N_2956);
and UO_178 (O_178,N_2946,N_2939);
nand UO_179 (O_179,N_2936,N_2942);
nand UO_180 (O_180,N_2977,N_2996);
and UO_181 (O_181,N_2952,N_2966);
and UO_182 (O_182,N_2955,N_2932);
and UO_183 (O_183,N_2977,N_2969);
nand UO_184 (O_184,N_2933,N_2953);
or UO_185 (O_185,N_2939,N_2943);
nor UO_186 (O_186,N_2955,N_2962);
nand UO_187 (O_187,N_2978,N_2979);
xnor UO_188 (O_188,N_2961,N_2977);
nand UO_189 (O_189,N_2947,N_2994);
nand UO_190 (O_190,N_2968,N_2928);
and UO_191 (O_191,N_2957,N_2991);
nand UO_192 (O_192,N_2990,N_2933);
and UO_193 (O_193,N_2957,N_2968);
and UO_194 (O_194,N_2995,N_2926);
nor UO_195 (O_195,N_2972,N_2990);
or UO_196 (O_196,N_2950,N_2944);
nor UO_197 (O_197,N_2995,N_2932);
xnor UO_198 (O_198,N_2943,N_2970);
and UO_199 (O_199,N_2927,N_2944);
and UO_200 (O_200,N_2997,N_2965);
nand UO_201 (O_201,N_2948,N_2957);
nor UO_202 (O_202,N_2943,N_2975);
or UO_203 (O_203,N_2969,N_2929);
nor UO_204 (O_204,N_2963,N_2956);
or UO_205 (O_205,N_2934,N_2977);
and UO_206 (O_206,N_2974,N_2932);
nand UO_207 (O_207,N_2927,N_2995);
nor UO_208 (O_208,N_2972,N_2943);
nor UO_209 (O_209,N_2950,N_2932);
and UO_210 (O_210,N_2976,N_2944);
nor UO_211 (O_211,N_2973,N_2994);
nor UO_212 (O_212,N_2933,N_2945);
nand UO_213 (O_213,N_2959,N_2941);
and UO_214 (O_214,N_2940,N_2999);
nand UO_215 (O_215,N_2988,N_2974);
nor UO_216 (O_216,N_2952,N_2941);
or UO_217 (O_217,N_2998,N_2948);
nor UO_218 (O_218,N_2998,N_2973);
nor UO_219 (O_219,N_2993,N_2986);
or UO_220 (O_220,N_2941,N_2962);
or UO_221 (O_221,N_2957,N_2940);
xnor UO_222 (O_222,N_2977,N_2950);
nand UO_223 (O_223,N_2972,N_2970);
nand UO_224 (O_224,N_2971,N_2974);
and UO_225 (O_225,N_2962,N_2935);
nor UO_226 (O_226,N_2941,N_2990);
or UO_227 (O_227,N_2946,N_2965);
or UO_228 (O_228,N_2928,N_2991);
nor UO_229 (O_229,N_2931,N_2944);
nand UO_230 (O_230,N_2965,N_2977);
and UO_231 (O_231,N_2958,N_2973);
or UO_232 (O_232,N_2999,N_2941);
nand UO_233 (O_233,N_2954,N_2937);
or UO_234 (O_234,N_2925,N_2929);
and UO_235 (O_235,N_2997,N_2938);
nor UO_236 (O_236,N_2948,N_2940);
and UO_237 (O_237,N_2987,N_2978);
or UO_238 (O_238,N_2959,N_2993);
and UO_239 (O_239,N_2992,N_2994);
nand UO_240 (O_240,N_2961,N_2958);
nor UO_241 (O_241,N_2948,N_2991);
and UO_242 (O_242,N_2996,N_2962);
xor UO_243 (O_243,N_2986,N_2994);
nand UO_244 (O_244,N_2967,N_2959);
nor UO_245 (O_245,N_2969,N_2959);
and UO_246 (O_246,N_2995,N_2966);
or UO_247 (O_247,N_2942,N_2982);
nor UO_248 (O_248,N_2989,N_2979);
nand UO_249 (O_249,N_2973,N_2995);
nand UO_250 (O_250,N_2937,N_2987);
xnor UO_251 (O_251,N_2988,N_2975);
and UO_252 (O_252,N_2931,N_2956);
xnor UO_253 (O_253,N_2933,N_2974);
nor UO_254 (O_254,N_2934,N_2960);
or UO_255 (O_255,N_2952,N_2986);
or UO_256 (O_256,N_2995,N_2935);
nor UO_257 (O_257,N_2976,N_2972);
nand UO_258 (O_258,N_2928,N_2984);
nor UO_259 (O_259,N_2936,N_2979);
and UO_260 (O_260,N_2928,N_2998);
nor UO_261 (O_261,N_2954,N_2930);
nor UO_262 (O_262,N_2926,N_2983);
nor UO_263 (O_263,N_2936,N_2930);
nand UO_264 (O_264,N_2933,N_2994);
nor UO_265 (O_265,N_2985,N_2967);
and UO_266 (O_266,N_2986,N_2979);
nor UO_267 (O_267,N_2959,N_2998);
xnor UO_268 (O_268,N_2986,N_2948);
or UO_269 (O_269,N_2996,N_2995);
or UO_270 (O_270,N_2925,N_2947);
and UO_271 (O_271,N_2980,N_2978);
nand UO_272 (O_272,N_2939,N_2937);
nor UO_273 (O_273,N_2948,N_2935);
nor UO_274 (O_274,N_2981,N_2964);
nor UO_275 (O_275,N_2941,N_2982);
or UO_276 (O_276,N_2945,N_2988);
and UO_277 (O_277,N_2961,N_2933);
nor UO_278 (O_278,N_2975,N_2958);
and UO_279 (O_279,N_2941,N_2928);
nor UO_280 (O_280,N_2979,N_2964);
xor UO_281 (O_281,N_2994,N_2978);
and UO_282 (O_282,N_2945,N_2983);
nor UO_283 (O_283,N_2946,N_2986);
xnor UO_284 (O_284,N_2936,N_2991);
or UO_285 (O_285,N_2972,N_2932);
nor UO_286 (O_286,N_2971,N_2999);
or UO_287 (O_287,N_2930,N_2993);
or UO_288 (O_288,N_2952,N_2983);
nor UO_289 (O_289,N_2999,N_2934);
and UO_290 (O_290,N_2993,N_2940);
or UO_291 (O_291,N_2975,N_2979);
or UO_292 (O_292,N_2970,N_2979);
or UO_293 (O_293,N_2962,N_2959);
nor UO_294 (O_294,N_2958,N_2942);
nand UO_295 (O_295,N_2956,N_2935);
nand UO_296 (O_296,N_2980,N_2983);
nand UO_297 (O_297,N_2993,N_2995);
nand UO_298 (O_298,N_2954,N_2939);
or UO_299 (O_299,N_2949,N_2960);
or UO_300 (O_300,N_2950,N_2963);
nor UO_301 (O_301,N_2954,N_2929);
nor UO_302 (O_302,N_2954,N_2963);
and UO_303 (O_303,N_2950,N_2955);
and UO_304 (O_304,N_2975,N_2982);
or UO_305 (O_305,N_2951,N_2994);
and UO_306 (O_306,N_2927,N_2960);
and UO_307 (O_307,N_2977,N_2930);
and UO_308 (O_308,N_2987,N_2935);
and UO_309 (O_309,N_2968,N_2966);
nand UO_310 (O_310,N_2986,N_2972);
or UO_311 (O_311,N_2979,N_2958);
and UO_312 (O_312,N_2975,N_2942);
or UO_313 (O_313,N_2947,N_2962);
nand UO_314 (O_314,N_2988,N_2960);
nor UO_315 (O_315,N_2984,N_2991);
nand UO_316 (O_316,N_2986,N_2957);
nand UO_317 (O_317,N_2997,N_2990);
nor UO_318 (O_318,N_2943,N_2974);
or UO_319 (O_319,N_2968,N_2976);
and UO_320 (O_320,N_2994,N_2961);
and UO_321 (O_321,N_2926,N_2966);
nor UO_322 (O_322,N_2962,N_2942);
nor UO_323 (O_323,N_2955,N_2930);
and UO_324 (O_324,N_2952,N_2995);
nor UO_325 (O_325,N_2931,N_2995);
nand UO_326 (O_326,N_2954,N_2945);
nor UO_327 (O_327,N_2937,N_2996);
and UO_328 (O_328,N_2975,N_2946);
nand UO_329 (O_329,N_2938,N_2934);
nand UO_330 (O_330,N_2926,N_2928);
nor UO_331 (O_331,N_2952,N_2976);
or UO_332 (O_332,N_2935,N_2997);
xor UO_333 (O_333,N_2993,N_2946);
and UO_334 (O_334,N_2996,N_2952);
or UO_335 (O_335,N_2933,N_2957);
nor UO_336 (O_336,N_2999,N_2962);
and UO_337 (O_337,N_2943,N_2985);
and UO_338 (O_338,N_2936,N_2999);
nand UO_339 (O_339,N_2987,N_2977);
and UO_340 (O_340,N_2955,N_2934);
and UO_341 (O_341,N_2960,N_2937);
and UO_342 (O_342,N_2964,N_2938);
xor UO_343 (O_343,N_2963,N_2990);
or UO_344 (O_344,N_2958,N_2990);
nand UO_345 (O_345,N_2951,N_2935);
or UO_346 (O_346,N_2943,N_2928);
nor UO_347 (O_347,N_2970,N_2950);
or UO_348 (O_348,N_2987,N_2992);
nor UO_349 (O_349,N_2992,N_2942);
and UO_350 (O_350,N_2985,N_2936);
nand UO_351 (O_351,N_2965,N_2983);
nor UO_352 (O_352,N_2954,N_2993);
or UO_353 (O_353,N_2930,N_2934);
nand UO_354 (O_354,N_2978,N_2996);
nor UO_355 (O_355,N_2982,N_2928);
and UO_356 (O_356,N_2926,N_2984);
and UO_357 (O_357,N_2995,N_2956);
nor UO_358 (O_358,N_2925,N_2972);
nor UO_359 (O_359,N_2950,N_2928);
or UO_360 (O_360,N_2969,N_2970);
nor UO_361 (O_361,N_2953,N_2937);
nand UO_362 (O_362,N_2997,N_2940);
or UO_363 (O_363,N_2984,N_2996);
and UO_364 (O_364,N_2961,N_2957);
or UO_365 (O_365,N_2995,N_2965);
or UO_366 (O_366,N_2974,N_2957);
or UO_367 (O_367,N_2949,N_2989);
or UO_368 (O_368,N_2971,N_2935);
nand UO_369 (O_369,N_2961,N_2971);
and UO_370 (O_370,N_2987,N_2976);
or UO_371 (O_371,N_2945,N_2965);
nand UO_372 (O_372,N_2948,N_2951);
or UO_373 (O_373,N_2974,N_2992);
and UO_374 (O_374,N_2997,N_2994);
and UO_375 (O_375,N_2953,N_2938);
and UO_376 (O_376,N_2994,N_2966);
or UO_377 (O_377,N_2944,N_2983);
nand UO_378 (O_378,N_2941,N_2946);
nor UO_379 (O_379,N_2996,N_2940);
nor UO_380 (O_380,N_2940,N_2972);
nor UO_381 (O_381,N_2933,N_2932);
nor UO_382 (O_382,N_2990,N_2946);
nor UO_383 (O_383,N_2952,N_2929);
or UO_384 (O_384,N_2999,N_2998);
or UO_385 (O_385,N_2990,N_2949);
or UO_386 (O_386,N_2931,N_2985);
and UO_387 (O_387,N_2946,N_2976);
nand UO_388 (O_388,N_2951,N_2982);
or UO_389 (O_389,N_2986,N_2964);
and UO_390 (O_390,N_2944,N_2935);
nor UO_391 (O_391,N_2937,N_2966);
nand UO_392 (O_392,N_2937,N_2993);
and UO_393 (O_393,N_2959,N_2946);
or UO_394 (O_394,N_2975,N_2945);
nor UO_395 (O_395,N_2969,N_2981);
or UO_396 (O_396,N_2959,N_2927);
nor UO_397 (O_397,N_2960,N_2968);
nor UO_398 (O_398,N_2954,N_2946);
nand UO_399 (O_399,N_2966,N_2991);
nand UO_400 (O_400,N_2937,N_2958);
and UO_401 (O_401,N_2926,N_2954);
nor UO_402 (O_402,N_2971,N_2977);
or UO_403 (O_403,N_2939,N_2964);
or UO_404 (O_404,N_2982,N_2984);
or UO_405 (O_405,N_2984,N_2953);
nor UO_406 (O_406,N_2961,N_2986);
or UO_407 (O_407,N_2948,N_2983);
and UO_408 (O_408,N_2946,N_2961);
or UO_409 (O_409,N_2968,N_2974);
nand UO_410 (O_410,N_2982,N_2966);
nand UO_411 (O_411,N_2973,N_2996);
nand UO_412 (O_412,N_2944,N_2986);
and UO_413 (O_413,N_2997,N_2943);
or UO_414 (O_414,N_2933,N_2958);
or UO_415 (O_415,N_2950,N_2954);
or UO_416 (O_416,N_2963,N_2958);
nand UO_417 (O_417,N_2992,N_2940);
or UO_418 (O_418,N_2970,N_2985);
nand UO_419 (O_419,N_2992,N_2984);
nand UO_420 (O_420,N_2998,N_2933);
or UO_421 (O_421,N_2987,N_2996);
nor UO_422 (O_422,N_2965,N_2928);
and UO_423 (O_423,N_2999,N_2937);
or UO_424 (O_424,N_2965,N_2996);
and UO_425 (O_425,N_2987,N_2958);
nand UO_426 (O_426,N_2998,N_2996);
or UO_427 (O_427,N_2945,N_2962);
nor UO_428 (O_428,N_2969,N_2935);
or UO_429 (O_429,N_2955,N_2976);
xor UO_430 (O_430,N_2991,N_2935);
and UO_431 (O_431,N_2953,N_2943);
nand UO_432 (O_432,N_2933,N_2938);
or UO_433 (O_433,N_2931,N_2940);
or UO_434 (O_434,N_2998,N_2974);
or UO_435 (O_435,N_2996,N_2963);
nor UO_436 (O_436,N_2972,N_2987);
nor UO_437 (O_437,N_2992,N_2926);
nor UO_438 (O_438,N_2960,N_2975);
nor UO_439 (O_439,N_2975,N_2976);
and UO_440 (O_440,N_2980,N_2931);
nand UO_441 (O_441,N_2947,N_2953);
xnor UO_442 (O_442,N_2997,N_2939);
or UO_443 (O_443,N_2965,N_2962);
nor UO_444 (O_444,N_2963,N_2937);
or UO_445 (O_445,N_2965,N_2964);
and UO_446 (O_446,N_2994,N_2984);
or UO_447 (O_447,N_2930,N_2984);
nor UO_448 (O_448,N_2931,N_2943);
nand UO_449 (O_449,N_2973,N_2929);
and UO_450 (O_450,N_2975,N_2929);
or UO_451 (O_451,N_2961,N_2927);
and UO_452 (O_452,N_2959,N_2994);
and UO_453 (O_453,N_2943,N_2982);
nand UO_454 (O_454,N_2945,N_2974);
nand UO_455 (O_455,N_2958,N_2932);
nand UO_456 (O_456,N_2931,N_2979);
nor UO_457 (O_457,N_2967,N_2977);
xor UO_458 (O_458,N_2992,N_2979);
nand UO_459 (O_459,N_2951,N_2972);
nand UO_460 (O_460,N_2945,N_2977);
and UO_461 (O_461,N_2957,N_2953);
nand UO_462 (O_462,N_2986,N_2985);
nor UO_463 (O_463,N_2993,N_2964);
nand UO_464 (O_464,N_2956,N_2928);
nand UO_465 (O_465,N_2948,N_2950);
and UO_466 (O_466,N_2957,N_2963);
nor UO_467 (O_467,N_2939,N_2938);
nor UO_468 (O_468,N_2942,N_2974);
or UO_469 (O_469,N_2998,N_2943);
or UO_470 (O_470,N_2976,N_2957);
and UO_471 (O_471,N_2980,N_2961);
nor UO_472 (O_472,N_2977,N_2976);
and UO_473 (O_473,N_2940,N_2981);
nor UO_474 (O_474,N_2949,N_2977);
xnor UO_475 (O_475,N_2965,N_2955);
or UO_476 (O_476,N_2952,N_2988);
or UO_477 (O_477,N_2967,N_2936);
and UO_478 (O_478,N_2934,N_2959);
or UO_479 (O_479,N_2960,N_2966);
nor UO_480 (O_480,N_2934,N_2989);
nor UO_481 (O_481,N_2974,N_2975);
nor UO_482 (O_482,N_2930,N_2952);
nor UO_483 (O_483,N_2934,N_2982);
nor UO_484 (O_484,N_2937,N_2968);
nor UO_485 (O_485,N_2956,N_2977);
nor UO_486 (O_486,N_2936,N_2974);
or UO_487 (O_487,N_2925,N_2949);
and UO_488 (O_488,N_2995,N_2967);
nand UO_489 (O_489,N_2996,N_2981);
nand UO_490 (O_490,N_2982,N_2965);
or UO_491 (O_491,N_2986,N_2976);
or UO_492 (O_492,N_2977,N_2959);
nand UO_493 (O_493,N_2967,N_2938);
nor UO_494 (O_494,N_2994,N_2977);
or UO_495 (O_495,N_2988,N_2957);
and UO_496 (O_496,N_2981,N_2999);
and UO_497 (O_497,N_2959,N_2974);
nor UO_498 (O_498,N_2998,N_2990);
nor UO_499 (O_499,N_2926,N_2999);
endmodule