module basic_5000_50000_5000_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_262,In_4747);
nor U1 (N_1,In_4217,In_3583);
nand U2 (N_2,In_65,In_895);
nand U3 (N_3,In_3356,In_4522);
and U4 (N_4,In_520,In_4991);
or U5 (N_5,In_4761,In_1295);
and U6 (N_6,In_4562,In_2104);
xnor U7 (N_7,In_3601,In_2961);
or U8 (N_8,In_2583,In_1671);
nand U9 (N_9,In_3213,In_64);
nand U10 (N_10,In_3972,In_2400);
xnor U11 (N_11,In_2378,In_1263);
nor U12 (N_12,In_2608,In_3649);
xnor U13 (N_13,In_2306,In_410);
nand U14 (N_14,In_2204,In_2933);
xnor U15 (N_15,In_664,In_967);
nand U16 (N_16,In_4682,In_1602);
nor U17 (N_17,In_18,In_354);
or U18 (N_18,In_3191,In_963);
or U19 (N_19,In_1825,In_2920);
xor U20 (N_20,In_2493,In_3065);
or U21 (N_21,In_4187,In_651);
nor U22 (N_22,In_188,In_2710);
and U23 (N_23,In_1929,In_468);
nand U24 (N_24,In_494,In_2633);
xnor U25 (N_25,In_3784,In_1636);
nor U26 (N_26,In_3690,In_3636);
xnor U27 (N_27,In_1326,In_275);
xnor U28 (N_28,In_662,In_3410);
or U29 (N_29,In_3225,In_4112);
nand U30 (N_30,In_3582,In_3140);
xnor U31 (N_31,In_297,In_564);
and U32 (N_32,In_1630,In_2977);
xor U33 (N_33,In_3192,In_3499);
nor U34 (N_34,In_4849,In_1612);
nor U35 (N_35,In_1845,In_1604);
or U36 (N_36,In_4156,In_1633);
or U37 (N_37,In_2112,In_2846);
or U38 (N_38,In_645,In_4732);
xor U39 (N_39,In_244,In_3640);
nor U40 (N_40,In_570,In_306);
nand U41 (N_41,In_1162,In_4139);
nand U42 (N_42,In_3044,In_3605);
xor U43 (N_43,In_754,In_3836);
xnor U44 (N_44,In_1288,In_4396);
nor U45 (N_45,In_3921,In_1559);
and U46 (N_46,In_3537,In_4371);
xor U47 (N_47,In_1331,In_3199);
and U48 (N_48,In_4153,In_3523);
and U49 (N_49,In_1672,In_2807);
and U50 (N_50,In_2757,In_4878);
or U51 (N_51,In_931,In_1275);
nand U52 (N_52,In_3984,In_4663);
or U53 (N_53,In_4226,In_4589);
xnor U54 (N_54,In_3956,In_4601);
xnor U55 (N_55,In_132,In_216);
xor U56 (N_56,In_1396,In_376);
or U57 (N_57,In_153,In_512);
and U58 (N_58,In_4475,In_948);
nor U59 (N_59,In_2407,In_3428);
or U60 (N_60,In_3378,In_471);
nor U61 (N_61,In_4310,In_1738);
xnor U62 (N_62,In_4972,In_4382);
nor U63 (N_63,In_1651,In_4800);
or U64 (N_64,In_688,In_2116);
nand U65 (N_65,In_3597,In_4468);
nand U66 (N_66,In_1567,In_2728);
and U67 (N_67,In_1476,In_4057);
or U68 (N_68,In_314,In_4042);
nand U69 (N_69,In_3619,In_4339);
xor U70 (N_70,In_4314,In_3206);
xnor U71 (N_71,In_122,In_3474);
nor U72 (N_72,In_4698,In_1367);
and U73 (N_73,In_2960,In_4242);
xnor U74 (N_74,In_2458,In_1104);
nor U75 (N_75,In_2232,In_1904);
or U76 (N_76,In_751,In_4911);
nand U77 (N_77,In_3067,In_247);
and U78 (N_78,In_941,In_3711);
nand U79 (N_79,In_1009,In_3749);
nand U80 (N_80,In_585,In_4889);
xnor U81 (N_81,In_355,In_4907);
nand U82 (N_82,In_2276,In_816);
xnor U83 (N_83,In_4062,In_2256);
nor U84 (N_84,In_3737,In_1042);
nand U85 (N_85,In_266,In_2936);
or U86 (N_86,In_545,In_2367);
nand U87 (N_87,In_1257,In_2878);
and U88 (N_88,In_556,In_415);
nand U89 (N_89,In_199,In_704);
and U90 (N_90,In_4517,In_804);
or U91 (N_91,In_272,In_3431);
xnor U92 (N_92,In_3674,In_2970);
nor U93 (N_93,In_2481,In_4600);
nand U94 (N_94,In_1281,In_4375);
and U95 (N_95,In_3261,In_2540);
nand U96 (N_96,In_3209,In_532);
or U97 (N_97,In_2001,In_1930);
or U98 (N_98,In_3832,In_3806);
nor U99 (N_99,In_2875,In_2840);
nor U100 (N_100,In_2981,In_91);
or U101 (N_101,In_1432,In_2330);
nand U102 (N_102,In_4291,In_4157);
or U103 (N_103,In_1858,In_3420);
and U104 (N_104,In_2855,In_1123);
nor U105 (N_105,In_4904,In_4304);
and U106 (N_106,In_1156,In_4367);
nor U107 (N_107,In_1780,In_752);
xnor U108 (N_108,In_261,In_4513);
nand U109 (N_109,In_2314,In_1193);
xnor U110 (N_110,In_3028,In_1054);
nor U111 (N_111,In_4587,In_3413);
and U112 (N_112,In_4539,In_489);
nor U113 (N_113,In_1371,In_345);
xnor U114 (N_114,In_4041,In_610);
xnor U115 (N_115,In_4084,In_3292);
nor U116 (N_116,In_4742,In_1942);
and U117 (N_117,In_2534,In_1032);
nor U118 (N_118,In_3501,In_825);
or U119 (N_119,In_2428,In_745);
and U120 (N_120,In_1495,In_1558);
xor U121 (N_121,In_4676,In_433);
nand U122 (N_122,In_2548,In_2226);
nor U123 (N_123,In_3091,In_829);
nand U124 (N_124,In_4701,In_3659);
nor U125 (N_125,In_235,In_2650);
nor U126 (N_126,In_1973,In_2081);
and U127 (N_127,In_1607,In_2909);
nor U128 (N_128,In_54,In_4709);
nand U129 (N_129,In_4995,In_2647);
nor U130 (N_130,In_3544,In_2562);
nor U131 (N_131,In_4903,In_1991);
or U132 (N_132,In_3119,In_4606);
and U133 (N_133,In_2423,In_2346);
xor U134 (N_134,In_403,In_4126);
and U135 (N_135,In_3020,In_4819);
nand U136 (N_136,In_1761,In_359);
xor U137 (N_137,In_1175,In_3023);
nor U138 (N_138,In_929,In_3114);
xor U139 (N_139,In_1664,In_909);
or U140 (N_140,In_3198,In_80);
and U141 (N_141,In_4428,In_971);
nand U142 (N_142,In_3155,In_102);
nand U143 (N_143,In_648,In_2582);
and U144 (N_144,In_4729,In_3968);
and U145 (N_145,In_1018,In_232);
nor U146 (N_146,In_4080,In_1874);
xor U147 (N_147,In_3258,In_2127);
nor U148 (N_148,In_1294,In_1817);
xor U149 (N_149,In_4093,In_2320);
or U150 (N_150,In_753,In_2337);
or U151 (N_151,In_4604,In_502);
or U152 (N_152,In_3918,In_707);
and U153 (N_153,In_4926,In_3170);
xor U154 (N_154,In_4221,In_861);
nand U155 (N_155,In_3411,In_500);
or U156 (N_156,In_224,In_4785);
and U157 (N_157,In_3855,In_3728);
nor U158 (N_158,In_2698,In_3657);
and U159 (N_159,In_2274,In_3087);
xor U160 (N_160,In_921,In_3571);
or U161 (N_161,In_1958,In_2721);
nor U162 (N_162,In_4982,In_414);
and U163 (N_163,In_4184,In_187);
xnor U164 (N_164,In_4104,In_3750);
nor U165 (N_165,In_3753,In_1730);
nand U166 (N_166,In_639,In_103);
or U167 (N_167,In_2445,In_332);
and U168 (N_168,In_2727,In_1434);
nand U169 (N_169,In_146,In_3117);
nor U170 (N_170,In_1499,In_2484);
nor U171 (N_171,In_3503,In_4832);
and U172 (N_172,In_2902,In_1028);
nor U173 (N_173,In_215,In_715);
nor U174 (N_174,In_624,In_3887);
nand U175 (N_175,In_1581,In_195);
nor U176 (N_176,In_789,In_172);
xor U177 (N_177,In_2305,In_3135);
or U178 (N_178,In_1964,In_2588);
and U179 (N_179,In_2043,In_4365);
and U180 (N_180,In_3600,In_1625);
nand U181 (N_181,In_2058,In_1024);
xor U182 (N_182,In_4658,In_2662);
nand U183 (N_183,In_66,In_2849);
and U184 (N_184,In_1226,In_1184);
or U185 (N_185,In_994,In_3061);
and U186 (N_186,In_2235,In_4256);
xnor U187 (N_187,In_4444,In_4462);
xor U188 (N_188,In_3025,In_2106);
nand U189 (N_189,In_3308,In_4614);
nor U190 (N_190,In_1595,In_4431);
or U191 (N_191,In_1613,In_577);
nor U192 (N_192,In_560,In_1401);
and U193 (N_193,In_3058,In_2790);
nand U194 (N_194,In_4870,In_2160);
or U195 (N_195,In_746,In_3365);
nor U196 (N_196,In_2244,In_3767);
and U197 (N_197,In_2778,In_2577);
xor U198 (N_198,In_543,In_2433);
and U199 (N_199,In_1348,In_1503);
and U200 (N_200,In_3884,In_12);
and U201 (N_201,In_2335,In_1884);
or U202 (N_202,In_4354,In_2336);
and U203 (N_203,In_818,In_2350);
and U204 (N_204,In_2990,In_2939);
and U205 (N_205,In_3970,In_2640);
or U206 (N_206,In_4790,In_154);
xnor U207 (N_207,In_4591,In_535);
or U208 (N_208,In_1366,In_4275);
nand U209 (N_209,In_661,In_4721);
xnor U210 (N_210,In_163,In_4131);
xor U211 (N_211,In_2464,In_69);
nor U212 (N_212,In_970,In_2556);
nor U213 (N_213,In_1161,In_1327);
or U214 (N_214,In_3374,In_2492);
nor U215 (N_215,In_2379,In_3184);
nor U216 (N_216,In_4830,In_3568);
nand U217 (N_217,In_17,In_358);
and U218 (N_218,In_3821,In_3684);
and U219 (N_219,In_4287,In_3775);
nor U220 (N_220,In_529,In_812);
and U221 (N_221,In_4605,In_4403);
or U222 (N_222,In_3340,In_125);
and U223 (N_223,In_311,In_522);
nor U224 (N_224,In_877,In_4755);
nor U225 (N_225,In_1287,In_2774);
nor U226 (N_226,In_469,In_2310);
nand U227 (N_227,In_4914,In_3536);
nand U228 (N_228,In_4681,In_3010);
xnor U229 (N_229,In_1227,In_3154);
xnor U230 (N_230,In_1598,In_1626);
xor U231 (N_231,In_1896,In_4265);
and U232 (N_232,In_350,In_2945);
or U233 (N_233,In_4316,In_4815);
xnor U234 (N_234,In_1159,In_3508);
xor U235 (N_235,In_2696,In_2820);
nor U236 (N_236,In_1648,In_811);
or U237 (N_237,In_2590,In_1860);
nor U238 (N_238,In_4295,In_3865);
nor U239 (N_239,In_760,In_4244);
xor U240 (N_240,In_2405,In_1336);
nor U241 (N_241,In_4413,In_807);
nor U242 (N_242,In_4264,In_583);
and U243 (N_243,In_1103,In_2730);
nand U244 (N_244,In_3997,In_4671);
or U245 (N_245,In_686,In_1324);
nor U246 (N_246,In_3335,In_2197);
or U247 (N_247,In_3532,In_4898);
or U248 (N_248,In_2821,In_4003);
or U249 (N_249,In_120,In_4398);
nand U250 (N_250,In_4888,In_4271);
xor U251 (N_251,In_1741,In_4777);
nand U252 (N_252,In_1554,In_2791);
or U253 (N_253,In_685,In_2927);
and U254 (N_254,In_3917,In_278);
nand U255 (N_255,In_4203,In_880);
or U256 (N_256,In_2083,In_3441);
nand U257 (N_257,In_3677,In_2580);
xor U258 (N_258,In_4844,In_4378);
or U259 (N_259,In_1208,In_3995);
xnor U260 (N_260,In_2731,In_3708);
and U261 (N_261,In_1143,In_4503);
nor U262 (N_262,In_340,In_2096);
and U263 (N_263,In_4306,In_3312);
xnor U264 (N_264,In_3455,In_2424);
xor U265 (N_265,In_620,In_4412);
nor U266 (N_266,In_1060,In_1519);
and U267 (N_267,In_1901,In_2039);
and U268 (N_268,In_2510,In_4569);
and U269 (N_269,In_4661,In_2829);
xor U270 (N_270,In_2622,In_2029);
nand U271 (N_271,In_2925,In_4665);
xor U272 (N_272,In_1497,In_3851);
and U273 (N_273,In_3320,In_4030);
xor U274 (N_274,In_4617,In_8);
nand U275 (N_275,In_2080,In_2281);
or U276 (N_276,In_2615,In_2668);
xor U277 (N_277,In_2308,In_3227);
nor U278 (N_278,In_365,In_1877);
and U279 (N_279,In_3498,In_3822);
nor U280 (N_280,In_1077,In_3400);
nor U281 (N_281,In_4703,In_2140);
xor U282 (N_282,In_1997,In_2701);
nand U283 (N_283,In_2653,In_428);
nand U284 (N_284,In_280,In_2142);
nor U285 (N_285,In_1518,In_178);
nand U286 (N_286,In_4654,In_3316);
nor U287 (N_287,In_1550,In_1752);
or U288 (N_288,In_955,In_4624);
nand U289 (N_289,In_3515,In_2296);
and U290 (N_290,In_2720,In_2794);
nand U291 (N_291,In_1763,In_4074);
nor U292 (N_292,In_94,In_4418);
xor U293 (N_293,In_2724,In_2661);
xnor U294 (N_294,In_2500,In_268);
nand U295 (N_295,In_1205,In_4842);
and U296 (N_296,In_4254,In_4100);
or U297 (N_297,In_2955,In_3004);
and U298 (N_298,In_2259,In_4115);
nand U299 (N_299,In_478,In_3736);
nand U300 (N_300,In_3768,In_3556);
xnor U301 (N_301,In_4469,In_4060);
and U302 (N_302,In_4890,In_606);
xnor U303 (N_303,In_3099,In_2738);
or U304 (N_304,In_900,In_554);
nor U305 (N_305,In_3969,In_1778);
xnor U306 (N_306,In_3481,In_1589);
nand U307 (N_307,In_4380,In_1873);
or U308 (N_308,In_3314,In_4646);
or U309 (N_309,In_1045,In_3440);
nor U310 (N_310,In_2365,In_3575);
xor U311 (N_311,In_1966,In_2028);
xor U312 (N_312,In_853,In_1674);
nor U313 (N_313,In_1306,In_4567);
and U314 (N_314,In_1806,In_2147);
or U315 (N_315,In_4399,In_61);
nor U316 (N_316,In_4236,In_4534);
nand U317 (N_317,In_2860,In_1109);
xor U318 (N_318,In_2587,In_2700);
or U319 (N_319,In_4099,In_4282);
xor U320 (N_320,In_1270,In_1391);
and U321 (N_321,In_352,In_4426);
xnor U322 (N_322,In_3263,In_708);
xor U323 (N_323,In_44,In_3304);
or U324 (N_324,In_2358,In_3562);
nor U325 (N_325,In_1443,In_2013);
nor U326 (N_326,In_4294,In_3414);
nand U327 (N_327,In_1023,In_3112);
or U328 (N_328,In_2623,In_3093);
or U329 (N_329,In_1900,In_3616);
and U330 (N_330,In_119,In_2628);
and U331 (N_331,In_4429,In_3422);
nor U332 (N_332,In_4633,In_2687);
and U333 (N_333,In_1491,In_164);
nand U334 (N_334,In_497,In_1774);
nand U335 (N_335,In_4554,In_1374);
or U336 (N_336,In_3942,In_456);
and U337 (N_337,In_3908,In_3927);
and U338 (N_338,In_1560,In_2268);
nor U339 (N_339,In_220,In_721);
or U340 (N_340,In_4067,In_798);
and U341 (N_341,In_2194,In_1838);
xor U342 (N_342,In_1526,In_765);
or U343 (N_343,In_4523,In_1556);
nor U344 (N_344,In_2191,In_1976);
and U345 (N_345,In_3149,In_1512);
xnor U346 (N_346,In_1398,In_3589);
nor U347 (N_347,In_3397,In_671);
xor U348 (N_348,In_697,In_4154);
nor U349 (N_349,In_231,In_2219);
or U350 (N_350,In_3476,In_1074);
nand U351 (N_351,In_4010,In_616);
or U352 (N_352,In_4861,In_2474);
nor U353 (N_353,In_4325,In_4002);
nor U354 (N_354,In_1236,In_3609);
and U355 (N_355,In_1911,In_2592);
nor U356 (N_356,In_677,In_3070);
nand U357 (N_357,In_4480,In_4223);
or U358 (N_358,In_2802,In_1949);
nor U359 (N_359,In_915,In_240);
and U360 (N_360,In_3847,In_3960);
nand U361 (N_361,In_3731,In_1245);
xor U362 (N_362,In_4374,In_1091);
nor U363 (N_363,In_2536,In_1540);
nor U364 (N_364,In_3788,In_3436);
nand U365 (N_365,In_1707,In_525);
xnor U366 (N_366,In_1988,In_2833);
nor U367 (N_367,In_482,In_1493);
xnor U368 (N_368,In_1421,In_3771);
and U369 (N_369,In_141,In_1785);
nor U370 (N_370,In_2678,In_4499);
xnor U371 (N_371,In_248,In_474);
nor U372 (N_372,In_4411,In_3951);
nand U373 (N_373,In_1676,In_2646);
xnor U374 (N_374,In_238,In_1428);
nor U375 (N_375,In_1320,In_1215);
nor U376 (N_376,In_883,In_1026);
nor U377 (N_377,In_2742,In_4088);
nor U378 (N_378,In_1583,In_969);
or U379 (N_379,In_3724,In_1268);
xor U380 (N_380,In_3306,In_4749);
and U381 (N_381,In_1642,In_3978);
nor U382 (N_382,In_1645,In_4805);
or U383 (N_383,In_3617,In_2971);
xnor U384 (N_384,In_479,In_2051);
or U385 (N_385,In_2439,In_3953);
nor U386 (N_386,In_4473,In_2324);
nor U387 (N_387,In_3376,In_3144);
nand U388 (N_388,In_1321,In_391);
nand U389 (N_389,In_168,In_3856);
and U390 (N_390,In_4147,In_4750);
nand U391 (N_391,In_2659,In_1766);
xor U392 (N_392,In_3699,In_2009);
nor U393 (N_393,In_553,In_1801);
xnor U394 (N_394,In_817,In_1235);
xor U395 (N_395,In_3870,In_680);
nor U396 (N_396,In_4497,In_4034);
nor U397 (N_397,In_1523,In_3224);
nor U398 (N_398,In_1001,In_2024);
xor U399 (N_399,In_2747,In_472);
nand U400 (N_400,In_2553,In_3014);
or U401 (N_401,In_4043,In_3277);
or U402 (N_402,In_334,In_1357);
nor U403 (N_403,In_1716,In_344);
nor U404 (N_404,In_2775,In_1809);
nand U405 (N_405,In_4559,In_3867);
nand U406 (N_406,In_892,In_4976);
or U407 (N_407,In_382,In_2811);
xor U408 (N_408,In_1600,In_4224);
nor U409 (N_409,In_3381,In_465);
nand U410 (N_410,In_4836,In_4470);
xnor U411 (N_411,In_3959,In_4450);
or U412 (N_412,In_4491,In_2621);
nand U413 (N_413,In_2542,In_1344);
xor U414 (N_414,In_1250,In_607);
or U415 (N_415,In_2409,In_922);
or U416 (N_416,In_1661,In_575);
nor U417 (N_417,In_1527,In_1836);
xor U418 (N_418,In_4183,In_4692);
and U419 (N_419,In_3437,In_4029);
nor U420 (N_420,In_2437,In_3835);
and U421 (N_421,In_4117,In_2507);
or U422 (N_422,In_3807,In_1865);
or U423 (N_423,In_3318,In_3449);
xor U424 (N_424,In_510,In_780);
or U425 (N_425,In_1262,In_4586);
nand U426 (N_426,In_4537,In_2416);
and U427 (N_427,In_1698,In_2515);
nor U428 (N_428,In_3818,In_4263);
and U429 (N_429,In_868,In_3006);
nand U430 (N_430,In_126,In_2550);
nand U431 (N_431,In_384,In_1889);
or U432 (N_432,In_4417,In_623);
and U433 (N_433,In_2918,In_329);
nor U434 (N_434,In_1631,In_702);
nand U435 (N_435,In_4745,In_1108);
and U436 (N_436,In_944,In_1217);
or U437 (N_437,In_3244,In_4969);
nand U438 (N_438,In_3220,In_3773);
and U439 (N_439,In_1974,In_108);
nor U440 (N_440,In_772,In_1906);
nor U441 (N_441,In_649,In_3379);
nand U442 (N_442,In_4728,In_4711);
nor U443 (N_443,In_3546,In_854);
xnor U444 (N_444,In_2125,In_399);
xor U445 (N_445,In_2393,In_3662);
and U446 (N_446,In_2797,In_3713);
nand U447 (N_447,In_914,In_2299);
nor U448 (N_448,In_339,In_2123);
nand U449 (N_449,In_4168,In_3247);
nor U450 (N_450,In_55,In_530);
and U451 (N_451,In_129,In_93);
xor U452 (N_452,In_4530,In_1282);
xor U453 (N_453,In_2697,In_4821);
and U454 (N_454,In_4174,In_2558);
or U455 (N_455,In_2394,In_4073);
or U456 (N_456,In_4794,In_86);
and U457 (N_457,In_1105,In_1767);
nand U458 (N_458,In_2810,In_2740);
xor U459 (N_459,In_3354,In_2755);
and U460 (N_460,In_612,In_3060);
nor U461 (N_461,In_206,In_3999);
and U462 (N_462,In_3069,In_875);
nor U463 (N_463,In_1811,In_4404);
and U464 (N_464,In_2218,In_3405);
or U465 (N_465,In_1992,In_4449);
or U466 (N_466,In_4405,In_3447);
nor U467 (N_467,In_790,In_3189);
nand U468 (N_468,In_1810,In_3257);
and U469 (N_469,In_3522,In_4039);
or U470 (N_470,In_3991,In_2386);
xnor U471 (N_471,In_4071,In_3913);
or U472 (N_472,In_2002,In_313);
and U473 (N_473,In_2538,In_4987);
nor U474 (N_474,In_3178,In_1004);
xnor U475 (N_475,In_4848,In_134);
and U476 (N_476,In_2010,In_4787);
nor U477 (N_477,In_1381,In_2207);
or U478 (N_478,In_518,In_3037);
and U479 (N_479,In_259,In_779);
and U480 (N_480,In_3327,In_4631);
nor U481 (N_481,In_2958,In_1885);
nand U482 (N_482,In_3309,In_3845);
nand U483 (N_483,In_390,In_2725);
nand U484 (N_484,In_4629,In_450);
nand U485 (N_485,In_1427,In_1043);
xor U486 (N_486,In_1148,In_4162);
and U487 (N_487,In_733,In_3939);
or U488 (N_488,In_748,In_1832);
nor U489 (N_489,In_3317,In_840);
xnor U490 (N_490,In_2520,In_1247);
nor U491 (N_491,In_2831,In_4940);
nor U492 (N_492,In_3620,In_11);
nor U493 (N_493,In_2351,In_1765);
xnor U494 (N_494,In_4760,In_726);
nor U495 (N_495,In_844,In_3602);
or U496 (N_496,In_145,In_1739);
and U497 (N_497,In_1177,In_888);
or U498 (N_498,In_3863,In_174);
and U499 (N_499,In_4596,In_3430);
or U500 (N_500,In_3324,In_605);
xor U501 (N_501,In_1228,In_2682);
xnor U502 (N_502,In_2457,In_4368);
and U503 (N_503,In_4735,In_4015);
or U504 (N_504,In_4258,In_750);
or U505 (N_505,In_2128,In_4445);
and U506 (N_506,In_1744,In_3697);
and U507 (N_507,In_4069,In_2851);
nand U508 (N_508,In_3359,In_3348);
nor U509 (N_509,In_1908,In_4044);
and U510 (N_510,In_1041,In_1561);
xor U511 (N_511,In_363,In_4619);
nor U512 (N_512,In_1463,In_1702);
nor U513 (N_513,In_855,In_3906);
nand U514 (N_514,In_3313,In_4137);
and U515 (N_515,In_2919,In_427);
and U516 (N_516,In_1999,In_4806);
xnor U517 (N_517,In_9,In_3796);
nor U518 (N_518,In_3294,In_3319);
and U519 (N_519,In_3056,In_1502);
or U520 (N_520,In_2799,In_3068);
xor U521 (N_521,In_2145,In_2169);
nand U522 (N_522,In_13,In_2767);
and U523 (N_523,In_1446,In_3326);
nand U524 (N_524,In_2282,In_1046);
xnor U525 (N_525,In_636,In_2077);
nand U526 (N_526,In_1229,In_1791);
and U527 (N_527,In_2297,In_3586);
nor U528 (N_528,In_2049,In_1037);
xor U529 (N_529,In_1160,In_3013);
nor U530 (N_530,In_3679,In_1875);
or U531 (N_531,In_2620,In_1426);
xor U532 (N_532,In_905,In_2143);
xor U533 (N_533,In_2756,In_643);
xor U534 (N_534,In_1418,In_3221);
and U535 (N_535,In_1242,In_1158);
or U536 (N_536,In_3071,In_630);
nor U537 (N_537,In_3564,In_2411);
or U538 (N_538,In_2449,In_4261);
or U539 (N_539,In_4362,In_3331);
xnor U540 (N_540,In_3607,In_4939);
or U541 (N_541,In_3459,In_2323);
and U542 (N_542,In_2450,In_3579);
xnor U543 (N_543,In_405,In_159);
nor U544 (N_544,In_185,In_1740);
xnor U545 (N_545,In_4989,In_4675);
nand U546 (N_546,In_3054,In_980);
nor U547 (N_547,In_58,In_4704);
nor U548 (N_548,In_4928,In_3641);
nand U549 (N_549,In_1945,In_3909);
nand U550 (N_550,In_4352,In_2788);
nand U551 (N_551,In_700,In_3098);
nand U552 (N_552,In_219,In_1380);
nand U553 (N_553,In_2941,In_4781);
and U554 (N_554,In_1311,In_2193);
nor U555 (N_555,In_4547,In_460);
and U556 (N_556,In_2005,In_204);
or U557 (N_557,In_3892,In_3686);
xnor U558 (N_558,In_258,In_1834);
and U559 (N_559,In_786,In_2059);
nor U560 (N_560,In_3525,In_2195);
xor U561 (N_561,In_1318,In_4259);
and U562 (N_562,In_4441,In_2518);
nor U563 (N_563,In_480,In_3841);
and U564 (N_564,In_3095,In_60);
nand U565 (N_565,In_1012,In_3236);
or U566 (N_566,In_1639,In_2825);
nand U567 (N_567,In_1545,In_4823);
nand U568 (N_568,In_4526,In_2604);
xor U569 (N_569,In_1587,In_2567);
nor U570 (N_570,In_590,In_1333);
nand U571 (N_571,In_3337,In_1453);
and U572 (N_572,In_444,In_3053);
nand U573 (N_573,In_2570,In_4772);
and U574 (N_574,In_2656,In_1793);
or U575 (N_575,In_3683,In_23);
or U576 (N_576,In_4479,In_1030);
nor U577 (N_577,In_2637,In_1853);
nand U578 (N_578,In_4007,In_4040);
xor U579 (N_579,In_4723,In_674);
nor U580 (N_580,In_3888,In_3262);
or U581 (N_581,In_2097,In_1307);
nand U582 (N_582,In_1925,In_4195);
xnor U583 (N_583,In_1285,In_2557);
nor U584 (N_584,In_1221,In_3299);
xor U585 (N_585,In_4072,In_4590);
or U586 (N_586,In_4260,In_4103);
xor U587 (N_587,In_3714,In_338);
or U588 (N_588,In_2236,In_4011);
xor U589 (N_589,In_2777,In_2261);
xor U590 (N_590,In_2470,In_4834);
and U591 (N_591,In_3592,In_372);
nand U592 (N_592,In_1951,In_189);
nor U593 (N_593,In_2911,In_1839);
nor U594 (N_594,In_1588,In_1922);
nand U595 (N_595,In_2907,In_1720);
nand U596 (N_596,In_2431,In_1376);
or U597 (N_597,In_1486,In_3982);
nor U598 (N_598,In_4102,In_3143);
and U599 (N_599,In_3175,In_2110);
and U600 (N_600,In_2359,In_641);
nand U601 (N_601,In_1691,In_631);
or U602 (N_602,In_995,In_1649);
nand U603 (N_603,In_2165,In_509);
nor U604 (N_604,In_3105,In_2965);
nand U605 (N_605,In_3783,In_3608);
xnor U606 (N_606,In_4063,In_273);
and U607 (N_607,In_3188,In_4886);
or U608 (N_608,In_1265,In_3465);
nor U609 (N_609,In_3086,In_4214);
nand U610 (N_610,In_1386,In_4638);
xnor U611 (N_611,In_1246,In_3829);
xnor U612 (N_612,In_4960,In_396);
or U613 (N_613,In_2111,In_296);
and U614 (N_614,In_2208,In_3384);
xnor U615 (N_615,In_2723,In_4563);
and U616 (N_616,In_4973,In_3748);
or U617 (N_617,In_4190,In_1356);
nor U618 (N_618,In_3889,In_2488);
xor U619 (N_619,In_2019,In_123);
nand U620 (N_620,In_533,In_4684);
nand U621 (N_621,In_2869,In_3047);
nor U622 (N_622,In_3973,In_3735);
or U623 (N_623,In_3936,In_4801);
and U624 (N_624,In_2769,In_4381);
and U625 (N_625,In_1851,In_2761);
and U626 (N_626,In_4970,In_254);
nor U627 (N_627,In_3089,In_3894);
or U628 (N_628,In_2000,In_4185);
nor U629 (N_629,In_3108,In_3007);
nand U630 (N_630,In_2609,In_4593);
nor U631 (N_631,In_1981,In_2912);
nand U632 (N_632,In_300,In_3229);
xor U633 (N_633,In_4509,In_588);
or U634 (N_634,In_766,In_2473);
xor U635 (N_635,In_4833,In_2192);
or U636 (N_636,In_4835,In_1803);
and U637 (N_637,In_3543,In_4076);
or U638 (N_638,In_100,In_3237);
xnor U639 (N_639,In_2313,In_2293);
nand U640 (N_640,In_3542,In_2749);
or U641 (N_641,In_516,In_3549);
xnor U642 (N_642,In_4127,In_1703);
nor U643 (N_643,In_511,In_1022);
nor U644 (N_644,In_4289,In_4786);
and U645 (N_645,In_1603,In_4822);
xnor U646 (N_646,In_466,In_589);
and U647 (N_647,In_4531,In_1125);
or U648 (N_648,In_39,In_1372);
nor U649 (N_649,In_2917,In_3922);
nand U650 (N_650,In_3201,In_871);
nor U651 (N_651,In_4387,In_3626);
and U652 (N_652,In_1243,In_3611);
xor U653 (N_653,In_2105,In_3353);
nand U654 (N_654,In_4472,In_3412);
xor U655 (N_655,In_2364,In_3520);
or U656 (N_656,In_594,In_441);
or U657 (N_657,In_214,In_2785);
and U658 (N_658,In_2499,In_4302);
and U659 (N_659,In_2490,In_3666);
nor U660 (N_660,In_852,In_1983);
xnor U661 (N_661,In_1111,In_521);
nand U662 (N_662,In_4485,In_4274);
or U663 (N_663,In_889,In_440);
nor U664 (N_664,In_1210,In_4390);
and U665 (N_665,In_2894,In_3780);
and U666 (N_666,In_3802,In_4333);
and U667 (N_667,In_3471,In_4828);
xnor U668 (N_668,In_2223,In_2036);
or U669 (N_669,In_2544,In_2442);
or U670 (N_670,In_1848,In_4452);
and U671 (N_671,In_3504,In_1820);
xor U672 (N_672,In_558,In_784);
nor U673 (N_673,In_252,In_3800);
and U674 (N_674,In_4825,In_162);
or U675 (N_675,In_2932,In_2676);
nand U676 (N_676,In_1341,In_3051);
nor U677 (N_677,In_4053,In_2453);
nand U678 (N_678,In_3925,In_4447);
or U679 (N_679,In_1541,In_2504);
and U680 (N_680,In_453,In_1025);
or U681 (N_681,In_437,In_4846);
and U682 (N_682,In_609,In_2861);
xnor U683 (N_683,In_2560,In_758);
nor U684 (N_684,In_2746,In_3179);
or U685 (N_685,In_3207,In_3588);
and U686 (N_686,In_2827,In_3529);
nor U687 (N_687,In_2418,In_1149);
or U688 (N_688,In_3814,In_3797);
nor U689 (N_689,In_2514,In_2549);
or U690 (N_690,In_2064,In_2602);
xor U691 (N_691,In_1117,In_1315);
nor U692 (N_692,In_2375,In_3985);
and U693 (N_693,In_1355,In_1776);
or U694 (N_694,In_4994,In_3637);
xnor U695 (N_695,In_3370,In_3387);
and U696 (N_696,In_4394,In_3103);
nand U697 (N_697,In_236,In_1469);
and U698 (N_698,In_4779,In_821);
nand U699 (N_699,In_847,In_3509);
nand U700 (N_700,In_1965,In_1358);
or U701 (N_701,In_169,In_3742);
and U702 (N_702,In_4016,In_336);
xor U703 (N_703,In_4005,In_2030);
xnor U704 (N_704,In_3919,In_4284);
or U705 (N_705,In_3940,In_2893);
or U706 (N_706,In_860,In_2652);
and U707 (N_707,In_1405,In_2501);
and U708 (N_708,In_327,In_928);
or U709 (N_709,In_863,In_2377);
xnor U710 (N_710,In_3618,In_2901);
xnor U711 (N_711,In_4237,In_3216);
nor U712 (N_712,In_1963,In_4199);
xnor U713 (N_713,In_3483,In_2750);
nor U714 (N_714,In_3603,In_2800);
or U715 (N_715,In_820,In_4668);
xnor U716 (N_716,In_898,In_1804);
nor U717 (N_717,In_3166,In_1340);
and U718 (N_718,In_2762,In_2946);
and U719 (N_719,In_109,In_2399);
nand U720 (N_720,In_1168,In_2130);
or U721 (N_721,In_3500,In_1750);
or U722 (N_722,In_2071,In_4720);
and U723 (N_723,In_4578,In_3701);
or U724 (N_724,In_1986,In_1058);
and U725 (N_725,In_3399,In_3297);
and U726 (N_726,In_4899,In_2613);
or U727 (N_727,In_418,In_1946);
nor U728 (N_728,In_2638,In_2717);
nor U729 (N_729,In_3810,In_2603);
nand U730 (N_730,In_1107,In_2951);
and U731 (N_731,In_3628,In_1048);
and U732 (N_732,In_2870,In_4094);
or U733 (N_733,In_3655,In_1189);
xnor U734 (N_734,In_1953,In_3896);
and U735 (N_735,In_4699,In_251);
xnor U736 (N_736,In_1116,In_2956);
nor U737 (N_737,In_3484,In_1085);
xor U738 (N_738,In_4118,In_3168);
or U739 (N_739,In_3475,In_4788);
or U740 (N_740,In_3260,In_452);
nand U741 (N_741,In_1521,In_582);
nor U742 (N_742,In_4607,In_4570);
nand U743 (N_743,In_4474,In_1186);
and U744 (N_744,In_3339,In_4196);
xnor U745 (N_745,In_1342,In_2171);
or U746 (N_746,In_4592,In_2781);
or U747 (N_747,In_1563,In_2612);
nor U748 (N_748,In_1579,In_2626);
nor U749 (N_749,In_2272,In_3516);
and U750 (N_750,In_4727,In_3816);
nor U751 (N_751,In_1578,In_3445);
and U752 (N_752,In_4383,In_703);
nand U753 (N_753,In_2984,In_4022);
or U754 (N_754,In_1950,In_1468);
nor U755 (N_755,In_4700,In_4487);
and U756 (N_756,In_2023,In_2595);
nor U757 (N_757,In_2610,In_972);
xnor U758 (N_758,In_1879,In_1566);
nand U759 (N_759,In_2391,In_2332);
nor U760 (N_760,In_1299,In_3083);
nor U761 (N_761,In_2325,In_849);
xnor U762 (N_762,In_3576,In_1802);
xor U763 (N_763,In_4033,In_4309);
and U764 (N_764,In_84,In_1547);
xor U765 (N_765,In_3528,In_2290);
nor U766 (N_766,In_4164,In_949);
nand U767 (N_767,In_679,In_429);
or U768 (N_768,In_4702,In_1297);
nor U769 (N_769,In_4824,In_654);
nand U770 (N_770,In_4863,In_3300);
nand U771 (N_771,In_19,In_1577);
xnor U772 (N_772,In_98,In_4296);
xor U773 (N_773,In_1683,In_487);
nor U774 (N_774,In_841,In_4783);
nor U775 (N_775,In_1417,In_4212);
or U776 (N_776,In_2456,In_3205);
nand U777 (N_777,In_3871,In_3720);
nand U778 (N_778,In_3223,In_4020);
and U779 (N_779,In_4955,In_2605);
and U780 (N_780,In_3805,In_4920);
nand U781 (N_781,In_2551,In_1938);
and U782 (N_782,In_1092,In_3785);
or U783 (N_783,In_4019,In_4440);
nand U784 (N_784,In_4054,In_4391);
or U785 (N_785,In_4211,In_136);
and U786 (N_786,In_2706,In_2994);
nand U787 (N_787,In_3124,In_2326);
or U788 (N_788,In_2180,In_2815);
and U789 (N_789,In_2976,In_2177);
xor U790 (N_790,In_4612,In_4155);
and U791 (N_791,In_2704,In_4966);
and U792 (N_792,In_2859,In_4205);
nand U793 (N_793,In_3506,In_256);
nand U794 (N_794,In_81,In_1689);
xor U795 (N_795,In_4142,In_2352);
nor U796 (N_796,In_2938,In_127);
nand U797 (N_797,In_2993,In_2921);
or U798 (N_798,In_2295,In_1047);
nand U799 (N_799,In_3254,In_3766);
xnor U800 (N_800,In_70,In_617);
nand U801 (N_801,In_422,In_4488);
or U802 (N_802,In_330,In_3204);
or U803 (N_803,In_1863,In_1667);
or U804 (N_804,In_2155,In_2497);
nand U805 (N_805,In_3203,In_1686);
or U806 (N_806,In_138,In_3338);
nand U807 (N_807,In_2373,In_1831);
nand U808 (N_808,In_4550,In_2889);
and U809 (N_809,In_4803,In_741);
nor U810 (N_810,In_4416,In_45);
or U811 (N_811,In_269,In_205);
or U812 (N_812,In_3837,In_302);
and U813 (N_813,In_2748,In_3897);
nor U814 (N_814,In_2220,In_3774);
nand U815 (N_815,In_4427,In_2086);
xnor U816 (N_816,In_1701,In_3126);
xor U817 (N_817,In_4331,In_357);
nand U818 (N_818,In_4,In_886);
or U819 (N_819,In_565,In_2506);
and U820 (N_820,In_1504,In_4881);
nor U821 (N_821,In_3893,In_4410);
and U822 (N_822,In_614,In_3330);
nand U823 (N_823,In_3752,In_3052);
and U824 (N_824,In_4300,In_2073);
and U825 (N_825,In_669,In_2436);
or U826 (N_826,In_353,In_3962);
nor U827 (N_827,In_3264,In_2702);
or U828 (N_828,In_3948,In_2923);
nand U829 (N_829,In_1605,In_2735);
nand U830 (N_830,In_3853,In_4009);
nand U831 (N_831,In_1029,In_1513);
and U832 (N_832,In_3090,In_201);
nand U833 (N_833,In_3315,In_2406);
or U834 (N_834,In_4350,In_3990);
xnor U835 (N_835,In_4198,In_308);
and U836 (N_836,In_4575,In_4999);
or U837 (N_837,In_3121,In_3820);
nand U838 (N_838,In_3351,In_4716);
nor U839 (N_839,In_3174,In_794);
and U840 (N_840,In_1987,In_1136);
xnor U841 (N_841,In_1346,In_78);
or U842 (N_842,In_1016,In_4630);
nand U843 (N_843,In_434,In_421);
nor U844 (N_844,In_4776,In_149);
xnor U845 (N_845,In_2528,In_714);
nor U846 (N_846,In_1480,In_245);
nand U847 (N_847,In_3687,In_3485);
and U848 (N_848,In_3293,In_4395);
xor U849 (N_849,In_4641,In_2202);
and U850 (N_850,In_4239,In_2928);
nand U851 (N_851,In_2692,In_3595);
and U852 (N_852,In_1697,In_4498);
and U853 (N_853,In_4909,In_1813);
and U854 (N_854,In_347,In_629);
xnor U855 (N_855,In_1027,In_2904);
nand U856 (N_856,In_874,In_2630);
or U857 (N_857,In_613,In_1439);
xor U858 (N_858,In_960,In_4222);
nor U859 (N_859,In_1926,In_3062);
nor U860 (N_860,In_602,In_891);
xnor U861 (N_861,In_1772,In_4770);
xnor U862 (N_862,In_3665,In_3514);
xor U863 (N_863,In_271,In_1485);
xnor U864 (N_864,In_1555,In_626);
nand U865 (N_865,In_4151,In_2316);
nand U866 (N_866,In_4406,In_1377);
xor U867 (N_867,In_4952,In_2806);
or U868 (N_868,In_2513,In_632);
or U869 (N_869,In_3798,In_1797);
xor U870 (N_870,In_1345,In_3267);
xnor U871 (N_871,In_2444,In_1002);
and U872 (N_872,In_1194,In_2175);
xor U873 (N_873,In_3015,In_1866);
or U874 (N_874,In_1814,In_4317);
or U875 (N_875,In_2693,In_4519);
and U876 (N_876,In_687,In_2524);
xnor U877 (N_877,In_1498,In_4255);
and U878 (N_878,In_3419,In_571);
and U879 (N_879,In_4111,In_756);
and U880 (N_880,In_2438,In_1783);
xor U881 (N_881,In_2784,In_1828);
xor U882 (N_882,In_467,In_242);
and U883 (N_883,In_1000,In_3904);
nand U884 (N_884,In_1790,In_3076);
xnor U885 (N_885,In_191,In_4762);
and U886 (N_886,In_1647,In_1655);
and U887 (N_887,In_2683,In_4713);
xnor U888 (N_888,In_1662,In_4081);
nor U889 (N_889,In_3804,In_3075);
and U890 (N_890,In_4566,In_1093);
nor U891 (N_891,In_2879,In_4876);
xor U892 (N_892,In_4867,In_1154);
or U893 (N_893,In_2287,In_4145);
nand U894 (N_894,In_3842,In_1735);
nand U895 (N_895,In_2312,In_4730);
xor U896 (N_896,In_906,In_1907);
nor U897 (N_897,In_4997,In_2119);
xnor U898 (N_898,In_1302,In_321);
or U899 (N_899,In_4268,In_1656);
nand U900 (N_900,In_3875,In_3958);
and U901 (N_901,In_2,In_569);
xnor U902 (N_902,In_4679,In_1267);
and U903 (N_903,In_4837,In_1844);
and U904 (N_904,In_2252,In_3470);
and U905 (N_905,In_4384,In_3578);
nor U906 (N_906,In_1462,In_4220);
xor U907 (N_907,In_423,In_2186);
nor U908 (N_908,In_3253,In_282);
xnor U909 (N_909,In_3610,In_918);
nand U910 (N_910,In_4574,In_1067);
nor U911 (N_911,In_1350,In_118);
nand U912 (N_912,In_800,In_4543);
nand U913 (N_913,In_1967,In_2913);
or U914 (N_914,In_723,In_1216);
and U915 (N_915,In_1233,In_360);
nand U916 (N_916,In_2291,In_3779);
nand U917 (N_917,In_3328,In_3332);
nand U918 (N_918,In_4913,In_1861);
and U919 (N_919,In_1237,In_1182);
nor U920 (N_920,In_4407,In_859);
nand U921 (N_921,In_1539,In_2521);
and U922 (N_922,In_1899,In_3497);
or U923 (N_923,In_2136,In_1139);
nor U924 (N_924,In_1757,In_1781);
nor U925 (N_925,In_1715,In_2527);
nor U926 (N_926,In_2196,In_1134);
nand U927 (N_927,In_749,In_3899);
nand U928 (N_928,In_2340,In_1163);
xor U929 (N_929,In_3190,In_3848);
or U930 (N_930,In_2052,In_3558);
or U931 (N_931,In_1035,In_2108);
or U932 (N_932,In_3963,In_792);
nor U933 (N_933,In_1126,In_2631);
nand U934 (N_934,In_4967,In_4098);
xnor U935 (N_935,In_684,In_2479);
nor U936 (N_936,In_393,In_4845);
nand U937 (N_937,In_1133,In_1223);
nor U938 (N_938,In_3427,In_1110);
nand U939 (N_939,In_4216,In_3833);
nor U940 (N_940,In_3496,In_633);
xnor U941 (N_941,In_3676,In_1102);
xor U942 (N_942,In_1565,In_361);
and U943 (N_943,In_4763,In_2174);
xor U944 (N_944,In_230,In_3077);
or U945 (N_945,In_1862,In_3467);
or U946 (N_946,In_4492,In_3347);
xnor U947 (N_947,In_1272,In_389);
nand U948 (N_948,In_1447,In_845);
or U949 (N_949,In_3290,In_4710);
nor U950 (N_950,In_1451,In_4545);
xnor U951 (N_951,In_4408,In_4925);
xor U952 (N_952,In_7,In_1152);
nor U953 (N_953,In_1179,In_499);
xnor U954 (N_954,In_666,In_3599);
or U955 (N_955,In_2547,In_737);
or U956 (N_956,In_2090,In_3839);
and U957 (N_957,In_2809,In_2262);
xor U958 (N_958,In_4588,In_559);
and U959 (N_959,In_3924,In_1699);
or U960 (N_960,In_4827,In_4860);
or U961 (N_961,In_3357,In_2288);
nand U962 (N_962,In_2823,In_1470);
nor U963 (N_963,In_4857,In_3702);
nor U964 (N_964,In_2099,In_1944);
or U965 (N_965,In_4726,In_343);
nor U966 (N_966,In_4854,In_2476);
nand U967 (N_967,In_2780,In_3593);
nand U968 (N_968,In_2619,In_1675);
nand U969 (N_969,In_4771,In_3177);
xor U970 (N_970,In_3046,In_2007);
nor U971 (N_971,In_4715,In_6);
or U972 (N_972,In_4233,In_317);
or U973 (N_973,In_3153,In_4923);
and U974 (N_974,In_2459,In_4957);
xor U975 (N_975,In_1248,In_4853);
nor U976 (N_976,In_1283,In_3828);
nand U977 (N_977,In_2853,In_1898);
or U978 (N_978,In_3992,In_292);
nor U979 (N_979,In_2532,In_4965);
nand U980 (N_980,In_2201,In_642);
and U981 (N_981,In_4089,In_1114);
nand U982 (N_982,In_4252,In_3587);
nand U983 (N_983,In_1773,In_4096);
nand U984 (N_984,In_3255,In_3048);
or U985 (N_985,In_1204,In_2472);
and U986 (N_986,In_3986,In_2465);
and U987 (N_987,In_3929,In_446);
xnor U988 (N_988,In_3946,In_194);
nand U989 (N_989,In_1916,In_3271);
and U990 (N_990,In_1852,In_2843);
and U991 (N_991,In_37,In_85);
xor U992 (N_992,In_924,In_2837);
and U993 (N_993,In_3429,In_1592);
xnor U994 (N_994,In_4228,In_416);
and U995 (N_995,In_923,In_1919);
xor U996 (N_996,In_1395,In_274);
nand U997 (N_997,In_4059,In_2995);
and U998 (N_998,In_1888,In_3761);
or U999 (N_999,In_2752,In_3944);
nor U1000 (N_1000,In_3627,In_2671);
nand U1001 (N_1001,In_143,In_3979);
nor U1002 (N_1002,In_1892,N_258);
xnor U1003 (N_1003,In_3418,In_3811);
nand U1004 (N_1004,In_1538,In_1404);
xnor U1005 (N_1005,In_3303,In_3038);
nand U1006 (N_1006,N_666,In_1349);
nor U1007 (N_1007,In_4028,In_773);
and U1008 (N_1008,In_79,In_1181);
nand U1009 (N_1009,N_286,N_273);
nor U1010 (N_1010,N_699,In_896);
and U1011 (N_1011,In_2440,In_99);
or U1012 (N_1012,In_1296,N_199);
nand U1013 (N_1013,In_3383,In_2224);
and U1014 (N_1014,In_3643,N_559);
nand U1015 (N_1015,N_647,N_762);
nor U1016 (N_1016,N_953,N_845);
and U1017 (N_1017,In_2283,In_1300);
nor U1018 (N_1018,In_1213,In_4576);
and U1019 (N_1019,In_3554,In_1982);
nand U1020 (N_1020,In_139,In_4092);
nor U1021 (N_1021,In_3466,In_2205);
nand U1022 (N_1022,N_648,In_1222);
nand U1023 (N_1023,In_4344,In_4924);
xor U1024 (N_1024,In_1531,In_4477);
or U1025 (N_1025,In_4434,In_3891);
nand U1026 (N_1026,In_2008,In_3561);
and U1027 (N_1027,In_2085,N_50);
nand U1028 (N_1028,In_557,In_2616);
or U1029 (N_1029,N_681,In_3248);
xor U1030 (N_1030,In_785,In_413);
nand U1031 (N_1031,N_89,In_2215);
nand U1032 (N_1032,In_4673,In_2354);
xnor U1033 (N_1033,In_4481,In_4049);
xnor U1034 (N_1034,In_771,In_83);
xor U1035 (N_1035,N_975,In_1280);
and U1036 (N_1036,N_491,In_165);
or U1037 (N_1037,In_1606,In_3646);
or U1038 (N_1038,In_1020,In_1872);
nor U1039 (N_1039,N_256,In_1472);
nor U1040 (N_1040,N_718,In_2344);
xor U1041 (N_1041,N_298,N_917);
xor U1042 (N_1042,In_4101,In_4150);
or U1043 (N_1043,In_0,In_3709);
xnor U1044 (N_1044,In_1220,In_524);
nor U1045 (N_1045,N_780,In_2880);
nand U1046 (N_1046,In_3989,In_2847);
nor U1047 (N_1047,In_755,N_138);
nor U1048 (N_1048,In_2818,In_2658);
nor U1049 (N_1049,N_69,In_4515);
xnor U1050 (N_1050,N_958,N_715);
or U1051 (N_1051,N_409,In_3234);
and U1052 (N_1052,In_2903,In_4858);
and U1053 (N_1053,In_1436,N_160);
nand U1054 (N_1054,In_4978,N_257);
xor U1055 (N_1055,In_1692,In_218);
or U1056 (N_1056,In_283,In_4163);
or U1057 (N_1057,In_1119,In_2079);
and U1058 (N_1058,In_1249,In_1170);
or U1059 (N_1059,In_2753,In_3782);
nor U1060 (N_1060,In_310,In_2867);
xor U1061 (N_1061,In_196,In_71);
and U1062 (N_1062,In_856,In_3212);
and U1063 (N_1063,In_4639,In_4359);
or U1064 (N_1064,N_36,In_1388);
or U1065 (N_1065,N_747,N_557);
xnor U1066 (N_1066,In_3488,In_2466);
nand U1067 (N_1067,In_4506,In_828);
and U1068 (N_1068,In_1303,In_2574);
and U1069 (N_1069,In_3751,N_175);
and U1070 (N_1070,In_2102,N_268);
and U1071 (N_1071,In_1039,In_3689);
xor U1072 (N_1072,In_1570,In_4880);
xor U1073 (N_1073,N_522,In_1277);
nor U1074 (N_1074,N_351,In_2461);
xnor U1075 (N_1075,In_1055,N_11);
nor U1076 (N_1076,In_2415,In_3398);
and U1077 (N_1077,In_4017,In_1960);
or U1078 (N_1078,In_676,In_4510);
xnor U1079 (N_1079,N_640,In_1553);
or U1080 (N_1080,In_3966,In_2152);
xor U1081 (N_1081,In_3521,In_2245);
nor U1082 (N_1082,In_3762,In_1279);
or U1083 (N_1083,In_3920,In_3270);
nand U1084 (N_1084,In_2699,In_951);
nand U1085 (N_1085,N_120,In_3739);
or U1086 (N_1086,In_1616,In_503);
nand U1087 (N_1087,In_842,In_1456);
nor U1088 (N_1088,In_318,N_963);
or U1089 (N_1089,N_914,In_1361);
nand U1090 (N_1090,In_289,In_930);
nand U1091 (N_1091,In_4608,In_43);
xor U1092 (N_1092,In_3692,In_2852);
or U1093 (N_1093,In_3868,In_3439);
and U1094 (N_1094,In_3305,In_640);
xor U1095 (N_1095,In_211,In_3606);
or U1096 (N_1096,In_3266,In_2511);
or U1097 (N_1097,In_1021,In_3131);
or U1098 (N_1098,N_506,In_2131);
nand U1099 (N_1099,N_961,N_669);
or U1100 (N_1100,In_4208,In_3573);
xnor U1101 (N_1101,In_377,In_1590);
xor U1102 (N_1102,N_21,In_1234);
and U1103 (N_1103,In_3541,N_827);
nor U1104 (N_1104,In_3663,In_4068);
nand U1105 (N_1105,In_3171,In_3834);
xor U1106 (N_1106,In_426,In_5);
xnor U1107 (N_1107,In_2997,In_4628);
xor U1108 (N_1108,In_4421,In_2834);
or U1109 (N_1109,N_578,N_763);
and U1110 (N_1110,N_508,In_4637);
nand U1111 (N_1111,N_438,In_3235);
nand U1112 (N_1112,N_363,In_3873);
nor U1113 (N_1113,In_2664,In_937);
nor U1114 (N_1114,N_526,In_4882);
or U1115 (N_1115,In_1073,In_1147);
or U1116 (N_1116,N_467,In_1815);
nand U1117 (N_1117,In_1542,In_3104);
or U1118 (N_1118,N_326,In_2645);
xnor U1119 (N_1119,N_493,In_1338);
nor U1120 (N_1120,In_2844,In_838);
nand U1121 (N_1121,In_4535,In_1745);
xor U1122 (N_1122,In_4106,In_1857);
and U1123 (N_1123,In_1634,In_1419);
xnor U1124 (N_1124,In_4789,In_3200);
or U1125 (N_1125,In_1910,In_77);
nor U1126 (N_1126,N_57,In_1088);
nand U1127 (N_1127,N_116,In_1659);
nor U1128 (N_1128,In_4290,In_2395);
nand U1129 (N_1129,In_1695,In_3673);
nor U1130 (N_1130,N_738,N_330);
or U1131 (N_1131,In_3790,In_1677);
or U1132 (N_1132,In_1694,N_193);
or U1133 (N_1133,In_3382,In_519);
and U1134 (N_1134,In_3685,In_1962);
nand U1135 (N_1135,N_472,In_3256);
nand U1136 (N_1136,In_22,In_890);
xor U1137 (N_1137,In_1609,In_3730);
nor U1138 (N_1138,In_2736,N_933);
xor U1139 (N_1139,In_601,N_187);
nand U1140 (N_1140,In_699,In_1343);
and U1141 (N_1141,N_774,In_4283);
and U1142 (N_1142,In_1723,In_3831);
and U1143 (N_1143,N_678,In_2522);
and U1144 (N_1144,In_4919,In_1360);
nand U1145 (N_1145,In_1688,In_4379);
xor U1146 (N_1146,N_152,In_4052);
or U1147 (N_1147,In_2292,N_205);
or U1148 (N_1148,In_3463,In_551);
nand U1149 (N_1149,N_730,In_3624);
and U1150 (N_1150,In_1954,In_4643);
xor U1151 (N_1151,N_532,In_1955);
or U1152 (N_1152,N_390,In_3653);
nor U1153 (N_1153,N_266,N_119);
or U1154 (N_1154,N_99,N_935);
and U1155 (N_1155,In_3268,In_2067);
and U1156 (N_1156,In_3194,In_728);
nor U1157 (N_1157,In_304,In_973);
or U1158 (N_1158,N_608,In_2065);
nand U1159 (N_1159,N_617,In_4324);
nand U1160 (N_1160,N_936,In_2813);
and U1161 (N_1161,In_299,N_909);
and U1162 (N_1162,In_505,In_3623);
and U1163 (N_1163,In_2531,N_476);
xnor U1164 (N_1164,N_551,In_226);
xor U1165 (N_1165,In_1407,N_389);
and U1166 (N_1166,In_3002,In_1173);
nor U1167 (N_1167,N_101,N_291);
and U1168 (N_1168,In_4696,In_3572);
nor U1169 (N_1169,In_473,In_3141);
nor U1170 (N_1170,In_1637,In_740);
or U1171 (N_1171,In_2040,In_2930);
and U1172 (N_1172,N_203,In_3669);
nor U1173 (N_1173,N_463,N_213);
and U1174 (N_1174,In_151,In_1643);
and U1175 (N_1175,In_3881,In_115);
xor U1176 (N_1176,In_4656,In_3622);
or U1177 (N_1177,In_4435,In_1444);
xor U1178 (N_1178,In_657,In_3957);
or U1179 (N_1179,In_1310,In_2137);
and U1180 (N_1180,In_1816,In_3022);
xor U1181 (N_1181,In_1008,In_2066);
or U1182 (N_1182,N_304,In_1883);
nand U1183 (N_1183,In_4433,N_745);
nand U1184 (N_1184,N_986,In_2822);
or U1185 (N_1185,N_80,In_3895);
and U1186 (N_1186,In_2271,In_1477);
nand U1187 (N_1187,In_1805,In_1571);
nand U1188 (N_1188,In_959,In_3453);
or U1189 (N_1189,In_2674,In_4875);
nor U1190 (N_1190,N_796,In_2625);
or U1191 (N_1191,In_2914,In_4466);
and U1192 (N_1192,In_1062,In_1251);
and U1193 (N_1193,In_2726,N_706);
nor U1194 (N_1194,In_2264,N_725);
xnor U1195 (N_1195,In_2078,N_834);
nand U1196 (N_1196,In_4238,N_893);
and U1197 (N_1197,In_1915,In_1933);
nand U1198 (N_1198,In_2675,N_265);
or U1199 (N_1199,In_316,In_4170);
and U1200 (N_1200,In_3151,N_582);
and U1201 (N_1201,In_124,N_993);
and U1202 (N_1202,In_2578,In_3981);
nor U1203 (N_1203,In_4599,In_1278);
or U1204 (N_1204,In_2016,In_2873);
nand U1205 (N_1205,In_3635,N_979);
or U1206 (N_1206,N_612,N_8);
or U1207 (N_1207,In_927,In_793);
and U1208 (N_1208,In_455,In_1274);
nand U1209 (N_1209,In_1069,N_433);
or U1210 (N_1210,In_3681,In_1492);
or U1211 (N_1211,In_386,In_2027);
or U1212 (N_1212,In_3134,In_727);
nand U1213 (N_1213,In_2303,In_1543);
and U1214 (N_1214,N_964,N_631);
nor U1215 (N_1215,In_1224,In_192);
nor U1216 (N_1216,In_1071,In_810);
and U1217 (N_1217,N_865,In_619);
nand U1218 (N_1218,In_943,In_4169);
or U1219 (N_1219,In_1365,In_3594);
xor U1220 (N_1220,In_2679,N_422);
or U1221 (N_1221,In_608,In_2842);
xor U1222 (N_1222,N_636,In_1238);
nor U1223 (N_1223,In_1770,In_203);
xnor U1224 (N_1224,N_705,In_3801);
xnor U1225 (N_1225,In_974,In_1078);
or U1226 (N_1226,In_4580,In_4896);
or U1227 (N_1227,N_573,In_1970);
or U1228 (N_1228,In_694,In_1089);
or U1229 (N_1229,In_2289,N_100);
nand U1230 (N_1230,In_1402,In_4516);
nor U1231 (N_1231,N_623,In_3150);
nand U1232 (N_1232,In_351,N_793);
nand U1233 (N_1233,In_14,N_923);
and U1234 (N_1234,In_1298,In_362);
nor U1235 (N_1235,In_1075,In_4232);
xor U1236 (N_1236,In_4341,In_527);
or U1237 (N_1237,In_4864,N_877);
nor U1238 (N_1238,In_1534,In_513);
xnor U1239 (N_1239,In_1199,In_2164);
nor U1240 (N_1240,In_3275,In_2886);
nor U1241 (N_1241,N_134,In_3001);
xor U1242 (N_1242,N_543,In_2897);
nand U1243 (N_1243,N_889,In_2101);
or U1244 (N_1244,In_3885,In_4484);
nand U1245 (N_1245,In_4975,In_1685);
nand U1246 (N_1246,In_2300,N_676);
or U1247 (N_1247,In_1557,In_4649);
nand U1248 (N_1248,In_4831,In_2053);
nand U1249 (N_1249,N_879,N_995);
and U1250 (N_1250,In_4160,In_2795);
and U1251 (N_1251,N_939,In_2413);
and U1252 (N_1252,N_468,In_3700);
and U1253 (N_1253,In_2494,In_4159);
and U1254 (N_1254,In_3050,In_2020);
and U1255 (N_1255,In_3901,In_3172);
nor U1256 (N_1256,In_2182,In_2685);
nor U1257 (N_1257,In_998,In_424);
or U1258 (N_1258,In_2883,In_3211);
and U1259 (N_1259,In_1269,In_3362);
or U1260 (N_1260,N_863,In_3923);
nor U1261 (N_1261,In_2250,In_976);
nor U1262 (N_1262,N_635,N_570);
or U1263 (N_1263,N_854,N_677);
or U1264 (N_1264,N_128,In_4581);
and U1265 (N_1265,In_1118,In_4865);
nand U1266 (N_1266,N_490,In_157);
and U1267 (N_1267,In_2839,In_4974);
xnor U1268 (N_1268,In_2681,In_4615);
or U1269 (N_1269,N_604,N_430);
xnor U1270 (N_1270,In_4471,In_1335);
xnor U1271 (N_1271,In_4766,In_2857);
nand U1272 (N_1272,In_4769,In_2267);
nand U1273 (N_1273,N_752,In_3218);
xor U1274 (N_1274,In_2667,In_2906);
nor U1275 (N_1275,In_3707,In_795);
xnor U1276 (N_1276,In_1941,In_4818);
and U1277 (N_1277,In_4708,In_3042);
xnor U1278 (N_1278,In_2184,N_216);
nand U1279 (N_1279,In_3819,In_932);
nor U1280 (N_1280,In_1057,In_4132);
xnor U1281 (N_1281,In_1100,In_3950);
nand U1282 (N_1282,In_3715,In_712);
or U1283 (N_1283,In_431,In_3843);
nor U1284 (N_1284,In_2978,In_4078);
nor U1285 (N_1285,In_4372,In_3705);
or U1286 (N_1286,N_700,N_118);
nand U1287 (N_1287,In_4386,In_3803);
and U1288 (N_1288,In_408,In_2238);
nor U1289 (N_1289,In_3334,In_4613);
xor U1290 (N_1290,N_484,In_3282);
nor U1291 (N_1291,In_463,In_1394);
nand U1292 (N_1292,In_4326,In_4482);
nor U1293 (N_1293,In_4495,In_2022);
and U1294 (N_1294,In_3791,In_2865);
or U1295 (N_1295,In_3096,In_2230);
xnor U1296 (N_1296,N_355,In_3367);
or U1297 (N_1297,N_161,In_3719);
and U1298 (N_1298,In_1886,N_575);
nor U1299 (N_1299,In_1798,In_3998);
nand U1300 (N_1300,N_296,In_1782);
or U1301 (N_1301,In_2943,In_3157);
xor U1302 (N_1302,In_3406,N_200);
nand U1303 (N_1303,N_924,N_810);
or U1304 (N_1304,In_2581,In_4954);
or U1305 (N_1305,In_3747,N_365);
or U1306 (N_1306,In_4023,In_4912);
nand U1307 (N_1307,In_2576,In_180);
nor U1308 (N_1308,In_2222,In_1696);
nand U1309 (N_1309,In_2934,N_43);
xor U1310 (N_1310,N_181,In_1614);
xor U1311 (N_1311,In_1652,In_3570);
and U1312 (N_1312,In_1094,N_883);
nor U1313 (N_1313,In_4585,In_1438);
nand U1314 (N_1314,In_3392,In_3815);
or U1315 (N_1315,N_798,In_2387);
xor U1316 (N_1316,N_220,N_142);
nor U1317 (N_1317,In_2385,In_4602);
nor U1318 (N_1318,N_284,In_288);
or U1319 (N_1319,In_1969,In_1464);
nand U1320 (N_1320,In_4273,N_54);
xnor U1321 (N_1321,In_1903,N_862);
xor U1322 (N_1322,In_3341,In_1188);
xor U1323 (N_1323,N_404,N_751);
and U1324 (N_1324,In_121,In_1905);
nand U1325 (N_1325,N_23,N_469);
nand U1326 (N_1326,In_439,In_3621);
nand U1327 (N_1327,In_1489,In_2905);
or U1328 (N_1328,In_1375,In_911);
nand U1329 (N_1329,In_2045,N_496);
xnor U1330 (N_1330,In_4353,N_135);
xnor U1331 (N_1331,In_3109,In_26);
xnor U1332 (N_1332,In_2012,In_2996);
xor U1333 (N_1333,In_4021,In_2338);
xor U1334 (N_1334,In_3682,In_2144);
or U1335 (N_1335,In_4808,In_3336);
and U1336 (N_1336,In_1090,In_788);
or U1337 (N_1337,In_4812,N_189);
nor U1338 (N_1338,In_1748,N_749);
nor U1339 (N_1339,In_4826,N_340);
and U1340 (N_1340,In_2596,In_1990);
and U1341 (N_1341,In_1325,In_4741);
nor U1342 (N_1342,N_238,In_3358);
and U1343 (N_1343,In_3003,In_4951);
and U1344 (N_1344,In_1146,In_2383);
xor U1345 (N_1345,In_3187,In_787);
xnor U1346 (N_1346,In_3438,In_961);
nand U1347 (N_1347,In_4409,In_2015);
or U1348 (N_1348,In_1622,In_263);
xnor U1349 (N_1349,In_3656,N_127);
and U1350 (N_1350,N_103,In_3580);
and U1351 (N_1351,N_501,In_1202);
and U1352 (N_1352,In_4871,In_1824);
nand U1353 (N_1353,In_1378,In_808);
and U1354 (N_1354,In_4500,In_2589);
and U1355 (N_1355,In_4561,N_28);
and U1356 (N_1356,In_4707,In_4678);
or U1357 (N_1357,N_269,In_656);
xor U1358 (N_1358,In_1363,N_156);
nand U1359 (N_1359,In_3360,In_1996);
nand U1360 (N_1360,In_4045,In_2021);
or U1361 (N_1361,N_223,N_447);
nand U1362 (N_1362,In_4303,In_1511);
or U1363 (N_1363,N_121,In_3952);
and U1364 (N_1364,In_1524,In_4149);
nor U1365 (N_1365,In_2452,In_2133);
nand U1366 (N_1366,In_1952,In_1731);
and U1367 (N_1367,N_139,N_987);
nand U1368 (N_1368,N_169,In_2963);
or U1369 (N_1369,N_425,N_0);
and U1370 (N_1370,In_46,In_233);
nand U1371 (N_1371,In_3493,In_4337);
and U1372 (N_1372,In_1635,N_253);
or U1373 (N_1373,In_2279,In_4250);
and U1374 (N_1374,In_3101,In_3059);
xor U1375 (N_1375,In_2356,In_1717);
xor U1376 (N_1376,N_144,In_1252);
or U1377 (N_1377,In_3817,In_4866);
nand U1378 (N_1378,In_778,In_2688);
or U1379 (N_1379,In_3574,N_451);
nand U1380 (N_1380,In_4820,In_902);
xor U1381 (N_1381,In_3019,N_47);
nand U1382 (N_1382,N_996,In_957);
xor U1383 (N_1383,In_1712,N_621);
or U1384 (N_1384,In_3138,N_474);
nor U1385 (N_1385,In_742,In_3878);
xor U1386 (N_1386,In_672,N_264);
xor U1387 (N_1387,In_572,In_374);
or U1388 (N_1388,N_949,N_664);
xor U1389 (N_1389,In_4527,In_4207);
and U1390 (N_1390,N_25,In_919);
nand U1391 (N_1391,N_420,N_354);
nor U1392 (N_1392,N_494,In_2286);
and U1393 (N_1393,In_32,N_734);
or U1394 (N_1394,In_3286,In_783);
xnor U1395 (N_1395,In_3364,In_381);
nor U1396 (N_1396,In_1721,In_2044);
or U1397 (N_1397,N_236,In_140);
nand U1398 (N_1398,In_1138,In_3106);
nand U1399 (N_1399,N_881,In_2561);
nor U1400 (N_1400,In_3394,N_530);
nand U1401 (N_1401,In_395,In_97);
nand U1402 (N_1402,In_2601,In_1063);
or U1403 (N_1403,In_1313,In_3063);
nor U1404 (N_1404,In_2991,In_3162);
nand U1405 (N_1405,In_2703,In_604);
nor U1406 (N_1406,In_1658,In_4636);
nor U1407 (N_1407,In_3208,In_1457);
xor U1408 (N_1408,In_2760,In_2796);
or U1409 (N_1409,In_3864,In_2670);
nor U1410 (N_1410,In_882,In_3217);
nor U1411 (N_1411,In_4129,N_591);
and U1412 (N_1412,In_2876,In_3704);
or U1413 (N_1413,N_267,In_894);
xnor U1414 (N_1414,In_4082,In_3722);
xor U1415 (N_1415,In_3830,In_3);
and U1416 (N_1416,In_370,In_3152);
nand U1417 (N_1417,N_9,In_4460);
and U1418 (N_1418,In_3540,In_1722);
or U1419 (N_1419,N_367,In_4938);
and U1420 (N_1420,In_4442,In_2783);
xor U1421 (N_1421,N_990,N_401);
nand U1422 (N_1422,N_411,N_182);
nand U1423 (N_1423,In_4349,In_1666);
nor U1424 (N_1424,N_146,In_3777);
xnor U1425 (N_1425,In_3487,In_4620);
nand U1426 (N_1426,In_2025,In_1203);
or U1427 (N_1427,In_4262,In_3242);
nand U1428 (N_1428,In_732,In_239);
or U1429 (N_1429,In_4584,In_904);
xnor U1430 (N_1430,N_464,In_1507);
nand U1431 (N_1431,N_724,In_62);
nor U1432 (N_1432,In_4840,In_1849);
xnor U1433 (N_1433,In_4097,In_2759);
nor U1434 (N_1434,N_978,In_2627);
and U1435 (N_1435,In_1789,N_811);
nand U1436 (N_1436,In_2334,In_3694);
or U1437 (N_1437,In_2564,In_4004);
nor U1438 (N_1438,In_4756,In_2517);
xor U1439 (N_1439,N_406,In_1796);
xor U1440 (N_1440,In_3511,In_3278);
and U1441 (N_1441,In_2862,In_4246);
and U1442 (N_1442,In_3703,In_2482);
and U1443 (N_1443,In_1719,In_3008);
xor U1444 (N_1444,N_277,In_835);
and U1445 (N_1445,In_2535,N_361);
and U1446 (N_1446,In_1180,In_4143);
and U1447 (N_1447,In_4347,In_701);
xor U1448 (N_1448,In_2069,In_2594);
or U1449 (N_1449,In_4553,In_2026);
xor U1450 (N_1450,In_1788,In_323);
xor U1451 (N_1451,In_1800,In_647);
and U1452 (N_1452,In_4616,N_599);
or U1453 (N_1453,In_850,N_86);
or U1454 (N_1454,N_306,N_315);
nor U1455 (N_1455,In_1747,In_4038);
nand U1456 (N_1456,N_515,In_1993);
nor U1457 (N_1457,In_981,N_310);
and U1458 (N_1458,In_4085,In_2212);
nand U1459 (N_1459,In_4141,In_2371);
xnor U1460 (N_1460,In_3478,In_3395);
or U1461 (N_1461,In_4598,In_2253);
nor U1462 (N_1462,N_246,N_67);
xor U1463 (N_1463,In_3226,In_942);
nor U1464 (N_1464,N_574,N_234);
xor U1465 (N_1465,In_4037,In_2384);
or U1466 (N_1466,In_3698,N_866);
nor U1467 (N_1467,In_2690,N_886);
nor U1468 (N_1468,In_1479,N_424);
and U1469 (N_1469,In_4075,In_3230);
nor U1470 (N_1470,In_4455,In_3111);
or U1471 (N_1471,In_3533,In_2629);
or U1472 (N_1472,In_2162,N_18);
and U1473 (N_1473,N_552,In_837);
or U1474 (N_1474,N_323,In_4272);
and U1475 (N_1475,N_345,In_3064);
nor U1476 (N_1476,In_3489,In_4292);
or U1477 (N_1477,In_486,In_1859);
nor U1478 (N_1478,N_819,In_2153);
and U1479 (N_1479,In_884,In_2114);
nand U1480 (N_1480,N_537,In_4321);
xor U1481 (N_1481,In_4622,In_2915);
and U1482 (N_1482,In_507,In_4947);
or U1483 (N_1483,In_3073,In_4956);
or U1484 (N_1484,In_735,In_1329);
or U1485 (N_1485,N_586,N_416);
nand U1486 (N_1486,In_2475,In_1641);
xor U1487 (N_1487,In_3080,In_2666);
nand U1488 (N_1488,In_1347,In_2575);
nand U1489 (N_1489,In_4135,N_479);
or U1490 (N_1490,In_2246,In_225);
nor U1491 (N_1491,N_370,In_3490);
nand U1492 (N_1492,In_3928,In_4743);
and U1493 (N_1493,In_4476,In_4892);
xor U1494 (N_1494,In_3473,In_447);
xor U1495 (N_1495,In_2999,In_1759);
and U1496 (N_1496,In_3799,In_2530);
nor U1497 (N_1497,In_2213,In_1549);
xor U1498 (N_1498,In_4422,N_96);
and U1499 (N_1499,In_250,In_2092);
or U1500 (N_1500,In_406,N_544);
nand U1501 (N_1501,N_153,N_357);
and U1502 (N_1502,N_316,In_4983);
or U1503 (N_1503,In_2311,N_450);
or U1504 (N_1504,N_655,In_4230);
nand U1505 (N_1505,In_4686,In_563);
and U1506 (N_1506,In_2091,In_3243);
nor U1507 (N_1507,In_3534,N_804);
or U1508 (N_1508,In_4791,In_4146);
and U1509 (N_1509,In_867,In_3133);
nand U1510 (N_1510,N_852,In_1190);
xnor U1511 (N_1511,In_621,In_41);
nor U1512 (N_1512,In_3712,In_2037);
or U1513 (N_1513,In_4971,In_4297);
or U1514 (N_1514,N_62,In_1516);
and U1515 (N_1515,In_2035,N_638);
nand U1516 (N_1516,In_1718,N_147);
and U1517 (N_1517,In_4859,In_4065);
nor U1518 (N_1518,N_722,N_856);
nor U1519 (N_1519,In_4961,In_4253);
nand U1520 (N_1520,In_4308,In_116);
or U1521 (N_1521,In_1036,N_59);
or U1522 (N_1522,N_502,In_4573);
xnor U1523 (N_1523,In_1155,N_667);
or U1524 (N_1524,In_2392,In_2887);
nand U1525 (N_1525,N_320,In_4241);
nor U1526 (N_1526,N_549,In_2353);
nand U1527 (N_1527,N_588,In_2333);
or U1528 (N_1528,In_4070,In_4180);
nand U1529 (N_1529,In_2054,In_4189);
and U1530 (N_1530,In_2972,In_4165);
xor U1531 (N_1531,N_697,N_5);
nand U1532 (N_1532,In_1003,In_2559);
or U1533 (N_1533,N_359,In_2979);
and U1534 (N_1534,In_209,In_182);
and U1535 (N_1535,N_194,N_817);
xor U1536 (N_1536,In_4752,In_2599);
and U1537 (N_1537,N_709,In_4953);
and U1538 (N_1538,N_982,In_3671);
nor U1539 (N_1539,In_665,In_4694);
nor U1540 (N_1540,In_4401,In_2109);
xor U1541 (N_1541,In_982,N_521);
or U1542 (N_1542,In_1033,In_658);
nor U1543 (N_1543,In_2248,N_743);
and U1544 (N_1544,In_2986,In_799);
xnor U1545 (N_1545,N_794,In_4436);
nor U1546 (N_1546,In_719,In_3850);
or U1547 (N_1547,In_2100,In_2665);
nand U1548 (N_1548,In_2804,In_1522);
nand U1549 (N_1549,In_3186,In_2266);
nor U1550 (N_1550,In_1878,In_4451);
and U1551 (N_1551,In_3945,N_460);
and U1552 (N_1552,In_747,In_1679);
or U1553 (N_1553,In_1403,In_1640);
and U1554 (N_1554,In_3911,In_1061);
xnor U1555 (N_1555,N_642,N_408);
nor U1556 (N_1556,In_3912,In_1753);
nor U1557 (N_1557,N_12,In_4551);
nand U1558 (N_1558,In_3757,In_2157);
nor U1559 (N_1559,In_1998,In_4504);
xnor U1560 (N_1560,In_4642,In_555);
nand U1561 (N_1561,In_2258,In_2427);
nor U1562 (N_1562,In_2095,N_379);
nand U1563 (N_1563,In_1975,In_3246);
xor U1564 (N_1564,In_3512,In_307);
or U1565 (N_1565,In_212,In_1309);
nand U1566 (N_1566,N_378,In_4276);
and U1567 (N_1567,In_3902,In_3808);
nor U1568 (N_1568,N_527,In_89);
and U1569 (N_1569,N_188,N_668);
and U1570 (N_1570,In_1317,In_4397);
xnor U1571 (N_1571,N_596,In_51);
or U1572 (N_1572,N_851,In_4122);
nor U1573 (N_1573,In_3738,In_2649);
and U1574 (N_1574,N_869,N_572);
or U1575 (N_1575,N_196,In_536);
or U1576 (N_1576,In_3880,In_2792);
and U1577 (N_1577,In_977,In_4234);
and U1578 (N_1578,In_1142,N_927);
and U1579 (N_1579,N_589,In_4990);
or U1580 (N_1580,N_329,In_4933);
nor U1581 (N_1581,In_2126,In_4736);
nor U1582 (N_1582,In_1176,In_644);
xor U1583 (N_1583,In_1440,N_412);
xnor U1584 (N_1584,In_4915,In_2068);
and U1585 (N_1585,In_1322,N_618);
xnor U1586 (N_1586,In_2401,In_4932);
and U1587 (N_1587,In_25,In_2451);
nor U1588 (N_1588,N_27,N_660);
and U1589 (N_1589,In_3569,N_457);
and U1590 (N_1590,In_74,In_3914);
nand U1591 (N_1591,In_2957,In_2877);
nor U1592 (N_1592,In_2686,In_27);
nor U1593 (N_1593,N_903,N_395);
nand U1594 (N_1594,In_646,In_3291);
xor U1595 (N_1595,In_3333,N_595);
or U1596 (N_1596,In_659,In_4248);
or U1597 (N_1597,In_4087,In_2614);
xor U1598 (N_1598,In_713,In_4315);
nand U1599 (N_1599,In_1769,In_4024);
nor U1600 (N_1600,In_2410,In_1708);
or U1601 (N_1601,In_4891,In_4757);
and U1602 (N_1602,In_4249,In_3502);
xnor U1603 (N_1603,In_1359,In_1214);
or U1604 (N_1604,In_285,In_3214);
nand U1605 (N_1605,In_4197,In_3249);
nor U1606 (N_1606,N_429,In_4392);
nor U1607 (N_1607,In_498,In_1638);
or U1608 (N_1608,In_3629,In_4158);
xnor U1609 (N_1609,In_3034,In_4176);
or U1610 (N_1610,In_144,In_1095);
nand U1611 (N_1611,In_3967,N_628);
or U1612 (N_1612,In_4984,In_2586);
or U1613 (N_1613,N_495,In_3018);
and U1614 (N_1614,In_1305,In_4179);
or U1615 (N_1615,In_3146,In_627);
xor U1616 (N_1616,N_533,In_3787);
nand U1617 (N_1617,In_2768,In_4121);
nand U1618 (N_1618,In_3994,N_629);
nor U1619 (N_1619,N_625,In_4439);
nor U1620 (N_1620,In_3740,In_470);
or U1621 (N_1621,In_4558,N_733);
xor U1622 (N_1622,In_4227,In_2552);
or U1623 (N_1623,In_3173,In_1490);
or U1624 (N_1624,In_768,In_595);
and U1625 (N_1625,In_2233,In_3307);
or U1626 (N_1626,N_83,In_202);
nand U1627 (N_1627,In_1856,N_971);
and U1628 (N_1628,In_4502,In_30);
nor U1629 (N_1629,In_3132,In_3343);
or U1630 (N_1630,In_2063,In_809);
or U1631 (N_1631,In_2672,In_3380);
and U1632 (N_1632,In_2047,N_920);
xor U1633 (N_1633,In_2734,In_1273);
or U1634 (N_1634,In_3219,In_3530);
nor U1635 (N_1635,N_613,N_801);
and U1636 (N_1636,In_3279,In_371);
or U1637 (N_1637,N_698,In_3813);
or U1638 (N_1638,In_4718,N_276);
or U1639 (N_1639,In_3861,In_35);
and U1640 (N_1640,In_4941,In_451);
nor U1641 (N_1641,N_252,In_4363);
nor U1642 (N_1642,N_290,In_1192);
nor U1643 (N_1643,In_3250,N_505);
nand U1644 (N_1644,In_1137,In_3197);
xor U1645 (N_1645,In_2600,In_1956);
xnor U1646 (N_1646,In_566,N_382);
and U1647 (N_1647,N_553,In_3183);
nor U1648 (N_1648,In_1328,In_4725);
nand U1649 (N_1649,In_4768,In_1693);
xor U1650 (N_1650,In_839,In_3045);
nand U1651 (N_1651,In_597,In_1411);
nand U1652 (N_1652,In_1034,In_3596);
or U1653 (N_1653,In_989,In_1596);
and U1654 (N_1654,In_4640,In_4373);
and U1655 (N_1655,N_968,In_2260);
xor U1656 (N_1656,In_4900,In_4235);
xor U1657 (N_1657,In_52,In_160);
xnor U1658 (N_1658,In_3849,In_4423);
nor U1659 (N_1659,N_170,In_2304);
and U1660 (N_1660,In_2983,In_2216);
and U1661 (N_1661,In_4921,N_720);
xor U1662 (N_1662,In_734,N_951);
nand U1663 (N_1663,In_3555,N_282);
xor U1664 (N_1664,N_755,In_2892);
and U1665 (N_1665,In_4764,In_1207);
nor U1666 (N_1666,In_885,In_567);
or U1667 (N_1667,In_1979,In_4454);
and U1668 (N_1668,In_3130,N_42);
and U1669 (N_1669,In_1316,In_4414);
nor U1670 (N_1670,In_1601,In_4862);
and U1671 (N_1671,In_3552,In_1728);
nor U1672 (N_1672,N_548,In_4648);
nand U1673 (N_1673,In_2835,In_1);
nor U1674 (N_1674,In_4611,N_859);
or U1675 (N_1675,N_91,N_358);
or U1676 (N_1676,In_260,In_2319);
and U1677 (N_1677,N_673,In_1211);
nor U1678 (N_1678,In_4278,In_4594);
nand U1679 (N_1679,In_179,N_414);
and U1680 (N_1680,In_2937,N_31);
xnor U1681 (N_1681,In_4508,In_2089);
nand U1682 (N_1682,In_4734,N_689);
or U1683 (N_1683,N_690,In_3716);
nand U1684 (N_1684,In_96,In_4489);
or U1685 (N_1685,In_3012,N_969);
nand U1686 (N_1686,In_4357,In_3547);
nand U1687 (N_1687,In_618,In_2502);
nand U1688 (N_1688,In_2814,In_380);
or U1689 (N_1689,In_1819,N_770);
and U1690 (N_1690,In_2368,In_2874);
and U1691 (N_1691,N_158,N_124);
nand U1692 (N_1692,In_246,In_375);
and U1693 (N_1693,In_724,In_2227);
and U1694 (N_1694,N_989,In_417);
nand U1695 (N_1695,In_4796,In_4852);
nor U1696 (N_1696,In_3823,In_1842);
and U1697 (N_1697,In_3507,In_3590);
or U1698 (N_1698,In_831,N_523);
xor U1699 (N_1699,In_2034,In_4651);
and U1700 (N_1700,In_1239,In_2151);
and U1701 (N_1701,In_1412,In_173);
and U1702 (N_1702,In_4632,N_108);
nand U1703 (N_1703,In_3729,In_1644);
xnor U1704 (N_1704,In_2178,N_908);
nor U1705 (N_1705,In_2254,N_897);
or U1706 (N_1706,In_161,In_4811);
xnor U1707 (N_1707,In_1422,N_580);
xor U1708 (N_1708,In_3789,In_1585);
or U1709 (N_1709,In_2989,In_2850);
and U1710 (N_1710,N_514,In_436);
nand U1711 (N_1711,In_1920,In_2198);
nor U1712 (N_1712,In_4124,In_1171);
or U1713 (N_1713,N_371,In_4342);
and U1714 (N_1714,N_214,In_2229);
or U1715 (N_1715,In_2751,N_754);
xor U1716 (N_1716,In_4346,In_1066);
or U1717 (N_1717,In_774,In_2848);
xnor U1718 (N_1718,N_861,In_1917);
nor U1719 (N_1719,In_2211,In_1597);
xor U1720 (N_1720,N_453,In_4784);
or U1721 (N_1721,In_858,In_2782);
nand U1722 (N_1722,In_4166,In_1732);
nor U1723 (N_1723,In_4929,In_4949);
and U1724 (N_1724,In_3491,In_1619);
nand U1725 (N_1725,In_2824,In_181);
xnor U1726 (N_1726,In_2190,In_1569);
or U1727 (N_1727,In_198,In_1460);
nor U1728 (N_1728,In_2134,In_379);
nor U1729 (N_1729,In_1011,In_1994);
xor U1730 (N_1730,In_4883,In_1657);
xor U1731 (N_1731,In_2498,In_4626);
and U1732 (N_1732,In_897,In_3123);
nand U1733 (N_1733,In_290,In_587);
and U1734 (N_1734,In_1937,N_531);
nor U1735 (N_1735,In_279,N_305);
or U1736 (N_1736,In_3613,In_3975);
nand U1737 (N_1737,In_1940,In_4181);
nand U1738 (N_1738,N_741,N_262);
nand U1739 (N_1739,In_2975,In_2255);
nor U1740 (N_1740,In_690,In_1663);
xor U1741 (N_1741,In_549,In_2360);
or U1742 (N_1742,In_869,N_212);
and U1743 (N_1743,In_2241,In_3916);
nand U1744 (N_1744,In_476,In_4753);
xor U1745 (N_1745,In_388,In_4318);
nand U1746 (N_1746,In_4048,In_4012);
nor U1747 (N_1747,N_289,N_884);
nor U1748 (N_1748,In_709,N_713);
nand U1749 (N_1749,N_946,In_2898);
or U1750 (N_1750,In_1912,In_4906);
xor U1751 (N_1751,In_490,In_4964);
and U1752 (N_1752,In_1891,In_2766);
or U1753 (N_1753,In_1435,In_445);
nand U1754 (N_1754,In_3165,In_1818);
xnor U1755 (N_1755,In_1308,In_4448);
or U1756 (N_1756,N_567,In_3156);
nor U1757 (N_1757,In_331,In_615);
nand U1758 (N_1758,In_879,In_1431);
or U1759 (N_1759,In_2737,N_564);
nor U1760 (N_1760,In_253,In_1209);
and U1761 (N_1761,In_2166,In_2712);
nor U1762 (N_1762,N_375,In_2495);
nand U1763 (N_1763,In_2343,In_3452);
nand U1764 (N_1764,In_4943,In_4916);
and U1765 (N_1765,In_1219,In_3457);
or U1766 (N_1766,In_2816,In_2129);
nand U1767 (N_1767,In_3425,N_413);
nand U1768 (N_1768,In_2776,In_3706);
nor U1769 (N_1769,In_1830,N_492);
or U1770 (N_1770,N_173,N_417);
nor U1771 (N_1771,In_1169,In_4319);
or U1772 (N_1772,In_4501,N_558);
xor U1773 (N_1773,N_761,N_183);
nor U1774 (N_1774,In_4731,In_4544);
nor U1775 (N_1775,N_757,In_3876);
nor U1776 (N_1776,In_1984,In_2181);
and U1777 (N_1777,In_3276,N_674);
xnor U1778 (N_1778,In_133,In_3718);
or U1779 (N_1779,N_313,N_34);
nor U1780 (N_1780,In_73,In_2885);
or U1781 (N_1781,In_1255,N_641);
or U1782 (N_1782,N_984,N_281);
xnor U1783 (N_1783,In_1843,In_1301);
nor U1784 (N_1784,In_710,N_10);
and U1785 (N_1785,In_3323,In_611);
nor U1786 (N_1786,In_2478,N_454);
and U1787 (N_1787,In_1611,N_767);
or U1788 (N_1788,In_1510,In_4931);
nand U1789 (N_1789,N_758,In_369);
or U1790 (N_1790,N_41,In_2046);
xor U1791 (N_1791,N_653,In_1031);
or U1792 (N_1792,N_858,In_2716);
xor U1793 (N_1793,In_2003,N_771);
nor U1794 (N_1794,In_2355,In_1864);
nand U1795 (N_1795,In_873,In_2715);
nor U1796 (N_1796,In_1151,In_3898);
nand U1797 (N_1797,In_1264,N_541);
or U1798 (N_1798,In_508,In_4557);
xnor U1799 (N_1799,In_2362,In_1441);
nor U1800 (N_1800,In_4754,In_1384);
xnor U1801 (N_1801,N_812,In_4669);
xor U1802 (N_1802,In_1196,N_872);
and U1803 (N_1803,In_4483,In_2033);
nor U1804 (N_1804,In_2744,N_955);
nand U1805 (N_1805,In_4175,N_68);
xor U1806 (N_1806,In_4719,In_4461);
nand U1807 (N_1807,In_4430,In_3385);
xor U1808 (N_1808,In_4267,In_2657);
and U1809 (N_1809,In_2968,In_2618);
nand U1810 (N_1810,In_1474,N_644);
xnor U1811 (N_1811,In_2695,In_1454);
or U1812 (N_1812,In_2845,In_3934);
or U1813 (N_1813,In_2209,N_434);
nor U1814 (N_1814,In_1924,N_911);
or U1815 (N_1815,In_3251,In_3825);
nor U1816 (N_1816,N_480,N_24);
xnor U1817 (N_1817,In_349,In_4047);
nor U1818 (N_1818,N_659,In_1430);
xor U1819 (N_1819,In_4552,In_4334);
or U1820 (N_1820,N_832,N_907);
or U1821 (N_1821,N_894,In_1044);
nand U1822 (N_1822,N_561,In_449);
and U1823 (N_1823,In_2635,In_2634);
nand U1824 (N_1824,In_1687,In_4627);
and U1825 (N_1825,N_318,In_673);
and U1826 (N_1826,In_2082,N_867);
and U1827 (N_1827,In_600,N_536);
xnor U1828 (N_1828,In_711,In_4992);
or U1829 (N_1829,In_155,In_4625);
and U1830 (N_1830,In_920,In_197);
xor U1831 (N_1831,In_716,In_2477);
or U1832 (N_1832,In_3877,N_20);
and U1833 (N_1833,In_4338,In_1700);
and U1834 (N_1834,In_901,In_1013);
nand U1835 (N_1835,In_1746,In_1520);
nor U1836 (N_1836,In_4644,N_516);
nor U1837 (N_1837,In_3563,In_1564);
or U1838 (N_1838,In_1373,In_3017);
xnor U1839 (N_1839,In_1936,In_2093);
xor U1840 (N_1840,In_454,N_113);
nor U1841 (N_1841,In_4335,N_723);
xor U1842 (N_1842,In_3854,In_2896);
nand U1843 (N_1843,In_3092,In_1968);
nor U1844 (N_1844,N_377,N_513);
or U1845 (N_1845,In_2496,In_1131);
and U1846 (N_1846,In_1876,In_346);
nor U1847 (N_1847,In_3393,In_1826);
nor U1848 (N_1848,In_1673,In_3302);
xnor U1849 (N_1849,N_540,In_3727);
and U1850 (N_1850,In_1533,N_292);
nand U1851 (N_1851,In_797,In_2402);
xnor U1852 (N_1852,In_462,In_1576);
nand U1853 (N_1853,In_400,N_649);
nand U1854 (N_1854,In_1122,In_4369);
xnor U1855 (N_1855,In_294,In_2651);
nand U1856 (N_1856,In_1854,N_19);
or U1857 (N_1857,In_493,In_1754);
nor U1858 (N_1858,In_1455,In_4895);
and U1859 (N_1859,In_893,In_2980);
and U1860 (N_1860,N_643,In_4298);
xor U1861 (N_1861,In_4597,In_4277);
or U1862 (N_1862,In_2505,In_2462);
and U1863 (N_1863,In_2593,N_249);
or U1864 (N_1864,In_1005,In_2161);
nand U1865 (N_1865,In_4458,In_4917);
nand U1866 (N_1866,In_4847,In_2636);
nor U1867 (N_1867,In_2446,In_496);
nor U1868 (N_1868,N_481,In_4281);
and U1869 (N_1869,In_4618,In_3415);
and U1870 (N_1870,In_4355,In_2048);
and U1871 (N_1871,In_293,In_2639);
xor U1872 (N_1872,N_339,In_95);
xor U1873 (N_1873,N_652,In_4345);
and U1874 (N_1874,In_2278,In_3368);
and U1875 (N_1875,N_308,In_3233);
nor U1876 (N_1876,In_3417,In_912);
xor U1877 (N_1877,In_983,In_3505);
and U1878 (N_1878,In_1191,In_1167);
nand U1879 (N_1879,In_2982,N_297);
nor U1880 (N_1880,In_284,In_4511);
nor U1881 (N_1881,N_321,N_885);
nand U1882 (N_1882,In_3295,In_1484);
xor U1883 (N_1883,In_528,N_563);
and U1884 (N_1884,In_2732,N_387);
or U1885 (N_1885,In_4443,In_4996);
xor U1886 (N_1886,N_443,In_348);
nor U1887 (N_1887,In_2309,N_598);
nor U1888 (N_1888,N_437,In_3746);
or U1889 (N_1889,In_4814,N_870);
xor U1890 (N_1890,In_4645,In_4018);
xor U1891 (N_1891,N_241,N_122);
or U1892 (N_1892,N_756,N_165);
and U1893 (N_1893,In_2321,In_2555);
xnor U1894 (N_1894,In_2654,N_294);
xor U1895 (N_1895,In_2327,In_938);
xor U1896 (N_1896,N_167,In_3409);
xnor U1897 (N_1897,N_683,N_686);
or U1898 (N_1898,In_2949,N_283);
and U1899 (N_1899,In_997,In_2284);
or U1900 (N_1900,In_3581,In_4872);
nand U1901 (N_1901,In_827,N_369);
xnor U1902 (N_1902,In_3287,In_1855);
nand U1903 (N_1903,In_2554,N_981);
nand U1904 (N_1904,In_1829,In_1017);
nor U1905 (N_1905,In_2969,In_1755);
xnor U1906 (N_1906,In_1140,In_1178);
xor U1907 (N_1907,In_4782,In_834);
or U1908 (N_1908,In_4910,In_3827);
or U1909 (N_1909,In_1076,N_6);
nand U1910 (N_1910,In_1985,In_2838);
and U1911 (N_1911,In_3639,In_1014);
and U1912 (N_1912,In_2339,In_291);
or U1913 (N_1913,N_415,N_560);
or U1914 (N_1914,In_739,In_2543);
nor U1915 (N_1915,In_736,In_539);
nor U1916 (N_1916,In_4520,N_455);
or U1917 (N_1917,In_1128,In_1758);
nand U1918 (N_1918,In_2179,In_2773);
or U1919 (N_1919,N_539,N_456);
or U1920 (N_1920,In_2243,In_1337);
or U1921 (N_1921,In_985,In_3389);
xnor U1922 (N_1922,In_325,N_159);
xnor U1923 (N_1923,N_823,In_4893);
and U1924 (N_1924,In_2199,N_913);
or U1925 (N_1925,In_2974,In_4659);
or U1926 (N_1926,In_2203,In_2388);
and U1927 (N_1927,N_278,In_4839);
nor U1928 (N_1928,In_2841,In_3033);
nor U1929 (N_1929,In_1624,In_4505);
and U1930 (N_1930,In_4329,In_3036);
nor U1931 (N_1931,In_2363,N_319);
xor U1932 (N_1932,In_171,In_3518);
nor U1933 (N_1933,In_50,In_3021);
and U1934 (N_1934,In_3585,In_3723);
nand U1935 (N_1935,In_4125,In_4817);
and U1936 (N_1936,In_3645,In_3651);
and U1937 (N_1937,N_130,N_499);
and U1938 (N_1938,In_1618,N_423);
or U1939 (N_1939,In_4565,In_1038);
nand U1940 (N_1940,In_4697,In_1286);
nor U1941 (N_1941,In_3404,In_301);
and U1942 (N_1942,In_4086,In_309);
and U1943 (N_1943,N_225,In_2441);
and U1944 (N_1944,N_88,In_3874);
and U1945 (N_1945,In_4993,In_200);
xor U1946 (N_1946,In_112,In_3661);
nor U1947 (N_1947,In_4621,In_4320);
or U1948 (N_1948,N_932,N_137);
nand U1949 (N_1949,In_1390,In_4689);
xnor U1950 (N_1950,N_2,In_1259);
xor U1951 (N_1951,In_3553,N_229);
or U1952 (N_1952,In_803,N_471);
and U1953 (N_1953,In_3285,In_2167);
nor U1954 (N_1954,In_4988,In_481);
nand U1955 (N_1955,In_4328,In_573);
or U1956 (N_1956,N_535,N_606);
xor U1957 (N_1957,In_2435,In_2966);
nand U1958 (N_1958,N_651,In_993);
nor U1959 (N_1959,N_775,In_3030);
nor U1960 (N_1960,N_875,In_4079);
or U1961 (N_1961,In_1174,N_17);
xor U1962 (N_1962,N_111,N_824);
and U1963 (N_1963,In_4229,In_668);
nor U1964 (N_1964,In_4288,In_4285);
and U1965 (N_1965,N_670,In_1379);
xor U1966 (N_1966,N_778,In_4690);
xor U1967 (N_1967,N_607,In_1293);
and U1968 (N_1968,N_991,N_594);
nand U1969 (N_1969,In_4792,In_1594);
nand U1970 (N_1970,N_942,In_3551);
xnor U1971 (N_1971,N_293,In_3078);
nand U1972 (N_1972,In_822,In_4740);
and U1973 (N_1973,N_611,In_2426);
nand U1974 (N_1974,In_2417,In_2566);
nor U1975 (N_1975,In_1751,N_219);
and U1976 (N_1976,In_3000,In_2916);
xnor U1977 (N_1977,In_1368,In_1452);
xnor U1978 (N_1978,In_4841,N_259);
and U1979 (N_1979,In_975,N_646);
nand U1980 (N_1980,In_4998,In_1339);
and U1981 (N_1981,In_2830,In_2503);
nand U1982 (N_1982,N_77,In_3612);
nand U1983 (N_1983,In_16,In_2454);
or U1984 (N_1984,In_999,In_1627);
or U1985 (N_1985,In_916,N_844);
nor U1986 (N_1986,In_156,In_1795);
nand U1987 (N_1987,N_898,In_2597);
nor U1988 (N_1988,N_123,In_4804);
or U1989 (N_1989,In_2798,In_1736);
and U1990 (N_1990,In_2863,In_763);
nor U1991 (N_1991,In_1668,In_3137);
nand U1992 (N_1992,In_3824,In_1141);
nor U1993 (N_1993,In_599,In_59);
and U1994 (N_1994,N_534,N_746);
and U1995 (N_1995,In_2519,In_4459);
nand U1996 (N_1996,In_364,In_2270);
or U1997 (N_1997,In_2122,N_3);
and U1998 (N_1998,In_1918,In_2819);
xnor U1999 (N_1999,In_925,In_3169);
xor U2000 (N_2000,N_488,In_4336);
xor U2001 (N_2001,In_3900,In_3444);
or U2002 (N_2002,In_3088,N_129);
nand U2003 (N_2003,In_443,N_226);
nor U2004 (N_2004,In_1425,In_1201);
nand U2005 (N_2005,N_828,N_1435);
and U2006 (N_2006,In_1711,In_4751);
or U2007 (N_2007,N_838,N_388);
xnor U2008 (N_2008,In_3648,N_1687);
and U2009 (N_2009,N_125,In_2812);
xnor U2010 (N_2010,In_2380,N_930);
nand U2011 (N_2011,N_1975,In_4032);
and U2012 (N_2012,N_1362,N_576);
nand U2013 (N_2013,N_905,In_3480);
xnor U2014 (N_2014,N_1407,In_3717);
or U2015 (N_2015,In_152,N_547);
nor U2016 (N_2016,In_4128,N_768);
xor U2017 (N_2017,N_1001,In_3915);
and U2018 (N_2018,N_1565,In_1473);
xnor U2019 (N_2019,N_1091,In_3781);
nor U2020 (N_2020,In_3344,N_904);
nor U2021 (N_2021,N_1296,In_3196);
nand U2022 (N_2022,In_4653,In_3288);
and U2023 (N_2023,In_4046,N_1962);
xnor U2024 (N_2024,N_1911,In_660);
nand U2025 (N_2025,In_2579,N_1358);
nor U2026 (N_2026,In_3139,In_4177);
and U2027 (N_2027,In_1706,N_1205);
nand U2028 (N_2028,N_1706,In_2432);
and U2029 (N_2029,In_1258,In_177);
nor U2030 (N_2030,In_3983,N_1639);
xnor U2031 (N_2031,N_1241,N_956);
or U2032 (N_2032,In_356,N_1018);
xor U2033 (N_2033,In_1458,In_3245);
and U2034 (N_2034,In_1690,N_222);
and U2035 (N_2035,In_775,N_1654);
nor U2036 (N_2036,N_92,N_890);
nor U2037 (N_2037,N_1336,In_2357);
nand U2038 (N_2038,N_769,N_1122);
nand U2039 (N_2039,In_2189,N_1031);
xor U2040 (N_2040,N_442,N_1934);
nand U2041 (N_2041,In_550,In_3464);
xor U2042 (N_2042,N_1788,In_3598);
or U2043 (N_2043,In_213,In_1351);
nand U2044 (N_2044,In_843,In_435);
nor U2045 (N_2045,In_1934,In_3346);
and U2046 (N_2046,N_1973,In_1115);
nor U2047 (N_2047,N_217,In_3210);
nand U2048 (N_2048,In_3980,In_3424);
nor U2049 (N_2049,In_147,In_4652);
nor U2050 (N_2050,N_38,N_1663);
and U2051 (N_2051,In_504,In_3468);
or U2052 (N_2052,In_580,In_67);
or U2053 (N_2053,N_1972,N_701);
nor U2054 (N_2054,In_4025,N_202);
nor U2055 (N_2055,In_2787,N_808);
or U2056 (N_2056,N_1938,In_2398);
or U2057 (N_2057,In_2508,In_2964);
or U2058 (N_2058,In_1195,N_802);
or U2059 (N_2059,In_4490,N_797);
nand U2060 (N_2060,N_1014,N_1851);
nand U2061 (N_2061,In_4134,In_3265);
xor U2062 (N_2062,N_172,N_1544);
xnor U2063 (N_2063,In_899,N_1789);
or U2064 (N_2064,In_2050,N_1088);
nor U2065 (N_2065,N_959,N_1381);
nor U2066 (N_2066,N_1287,N_1472);
xnor U2067 (N_2067,In_3658,In_3495);
xnor U2068 (N_2068,N_788,In_3883);
nand U2069 (N_2069,In_4979,In_1465);
nand U2070 (N_2070,In_4778,In_2280);
xor U2071 (N_2071,In_3869,N_1432);
nand U2072 (N_2072,N_696,In_4364);
nor U2073 (N_2073,In_4167,In_3758);
xnor U2074 (N_2074,In_1051,In_2247);
and U2075 (N_2075,N_1110,N_1019);
nand U2076 (N_2076,In_4457,N_764);
or U2077 (N_2077,N_126,In_1187);
nor U2078 (N_2078,In_1334,In_2307);
xnor U2079 (N_2079,N_337,N_1920);
nand U2080 (N_2080,N_1982,N_190);
nand U2081 (N_2081,In_2779,N_343);
and U2082 (N_2082,In_128,In_2150);
xor U2083 (N_2083,N_630,N_1971);
xor U2084 (N_2084,In_2899,In_3852);
nor U2085 (N_2085,In_1010,N_1061);
xnor U2086 (N_2086,In_4311,In_2509);
nor U2087 (N_2087,N_1299,N_1007);
nor U2088 (N_2088,N_1623,In_1049);
nor U2089 (N_2089,N_1216,N_1017);
xnor U2090 (N_2090,N_999,In_4688);
and U2091 (N_2091,N_1411,N_1426);
or U2092 (N_2092,In_4000,In_4874);
nand U2093 (N_2093,In_2632,N_601);
nor U2094 (N_2094,N_665,In_1475);
xnor U2095 (N_2095,In_4672,N_916);
nor U2096 (N_2096,N_1958,In_3548);
and U2097 (N_2097,In_4006,In_3432);
and U2098 (N_2098,N_892,In_3426);
or U2099 (N_2099,N_341,In_2159);
and U2100 (N_2100,N_1605,N_874);
nand U2101 (N_2101,In_1632,N_1087);
nand U2102 (N_2102,In_2032,N_154);
nand U2103 (N_2103,In_4802,In_1887);
nor U2104 (N_2104,In_4582,In_2075);
and U2105 (N_2105,In_966,N_65);
xor U2106 (N_2106,N_1234,N_1067);
and U2107 (N_2107,In_534,N_1829);
or U2108 (N_2108,In_1230,N_1064);
nor U2109 (N_2109,In_2141,In_913);
xnor U2110 (N_2110,In_3652,In_1551);
xor U2111 (N_2111,In_3907,N_1004);
nand U2112 (N_2112,In_1710,N_1609);
nand U2113 (N_2113,N_1330,N_1430);
and U2114 (N_2114,In_49,N_53);
or U2115 (N_2115,N_197,N_988);
nor U2116 (N_2116,In_4389,N_658);
and U2117 (N_2117,In_3477,In_1240);
or U2118 (N_2118,N_1508,N_1739);
and U2119 (N_2119,In_2882,N_1660);
or U2120 (N_2120,N_1461,N_421);
nand U2121 (N_2121,In_4647,N_1728);
nor U2122 (N_2122,In_538,In_4419);
nor U2123 (N_2123,N_1640,In_3433);
nor U2124 (N_2124,In_2713,In_4105);
and U2125 (N_2125,N_1046,N_603);
xor U2126 (N_2126,In_2349,In_4013);
xnor U2127 (N_2127,N_1986,In_1749);
and U2128 (N_2128,In_2836,N_1812);
xor U2129 (N_2129,N_45,In_1121);
and U2130 (N_2130,In_3615,In_3559);
or U2131 (N_2131,N_1587,N_143);
nor U2132 (N_2132,N_1783,N_1491);
and U2133 (N_2133,N_1438,N_1865);
xor U2134 (N_2134,N_1857,N_1755);
xor U2135 (N_2135,In_3638,N_1987);
nand U2136 (N_2136,In_683,In_2421);
and U2137 (N_2137,N_1132,N_826);
and U2138 (N_2138,In_281,In_3695);
nand U2139 (N_2139,In_593,In_3232);
xor U2140 (N_2140,N_528,In_1913);
and U2141 (N_2141,In_1332,N_1025);
xnor U2142 (N_2142,In_1200,In_113);
xor U2143 (N_2143,In_461,In_1387);
xnor U2144 (N_2144,In_3097,N_1860);
or U2145 (N_2145,In_4312,In_984);
nand U2146 (N_2146,N_1628,N_839);
and U2147 (N_2147,N_926,N_1968);
or U2148 (N_2148,In_3469,In_3390);
xor U2149 (N_2149,In_3377,In_1921);
nor U2150 (N_2150,N_1246,In_887);
or U2151 (N_2151,In_1762,N_162);
nor U2152 (N_2152,N_1331,In_717);
or U2153 (N_2153,N_302,N_1740);
and U2154 (N_2154,In_3460,N_1607);
xor U2155 (N_2155,In_3565,N_1191);
xor U2156 (N_2156,N_1166,N_1821);
or U2157 (N_2157,In_1959,N_1231);
or U2158 (N_2158,In_1734,N_1086);
xnor U2159 (N_2159,N_1634,N_772);
or U2160 (N_2160,N_682,In_3882);
nand U2161 (N_2161,N_1781,In_4935);
nand U2162 (N_2162,N_1147,N_1221);
and U2163 (N_2163,In_4855,N_410);
or U2164 (N_2164,N_1158,In_4963);
and U2165 (N_2165,N_1837,N_191);
nor U2166 (N_2166,N_891,In_3937);
and U2167 (N_2167,In_3281,N_498);
xnor U2168 (N_2168,N_1753,In_3786);
or U2169 (N_2169,In_542,N_1825);
nor U2170 (N_2170,In_2573,N_1344);
nand U2171 (N_2171,N_1917,In_4376);
nor U2172 (N_2172,N_1513,In_305);
xor U2173 (N_2173,In_3416,In_4635);
and U2174 (N_2174,In_4667,N_868);
nand U2175 (N_2175,In_2135,N_207);
xor U2176 (N_2176,In_3961,N_106);
xor U2177 (N_2177,N_1239,N_1408);
nand U2178 (N_2178,In_3016,In_3269);
nand U2179 (N_2179,In_2591,In_2729);
and U2180 (N_2180,In_2828,In_1684);
and U2181 (N_2181,N_1328,N_115);
xnor U2182 (N_2182,N_1916,N_748);
nor U2183 (N_2183,In_4327,N_242);
or U2184 (N_2184,In_3560,N_1270);
xor U2185 (N_2185,N_1473,N_740);
xnor U2186 (N_2186,In_2370,N_1350);
or U2187 (N_2187,In_4343,In_3932);
xor U2188 (N_2188,In_2103,In_1714);
nor U2189 (N_2189,In_598,N_1863);
and U2190 (N_2190,N_1049,In_2361);
nand U2191 (N_2191,N_1835,In_4120);
and U2192 (N_2192,N_1209,In_2660);
nand U2193 (N_2193,In_53,In_1084);
and U2194 (N_2194,N_328,In_3057);
or U2195 (N_2195,In_148,In_411);
nor U2196 (N_2196,N_1579,N_1774);
and U2197 (N_2197,N_1869,In_3329);
or U2198 (N_2198,In_1812,In_2006);
xnor U2199 (N_2199,In_2954,In_1323);
xor U2200 (N_2200,In_2864,In_4521);
or U2201 (N_2201,N_418,In_3239);
and U2202 (N_2202,N_56,In_2060);
nand U2203 (N_2203,In_4313,N_1349);
xor U2204 (N_2204,N_1923,N_1627);
or U2205 (N_2205,N_556,N_1596);
nand U2206 (N_2206,In_4541,In_477);
xnor U2207 (N_2207,In_183,In_4083);
and U2208 (N_2208,In_1978,In_4560);
xnor U2209 (N_2209,N_1608,N_274);
and U2210 (N_2210,In_2121,In_2120);
and U2211 (N_2211,In_217,In_2563);
nor U2212 (N_2212,In_2854,In_1212);
xnor U2213 (N_2213,In_4446,N_1632);
or U2214 (N_2214,N_965,In_432);
nor U2215 (N_2215,N_1372,In_1253);
or U2216 (N_2216,In_3094,In_2302);
nand U2217 (N_2217,N_1705,N_610);
or U2218 (N_2218,In_368,N_1416);
or U2219 (N_2219,N_1515,N_614);
nor U2220 (N_2220,N_1257,N_1141);
nor U2221 (N_2221,N_1090,In_412);
nor U2222 (N_2222,N_1227,N_1678);
nand U2223 (N_2223,N_307,N_1765);
xor U2224 (N_2224,In_1548,In_4192);
or U2225 (N_2225,N_504,N_1263);
nand U2226 (N_2226,In_4393,N_1855);
or U2227 (N_2227,In_667,N_692);
nor U2228 (N_2228,In_3310,In_3795);
and U2229 (N_2229,N_1383,In_1290);
or U2230 (N_2230,N_1887,In_249);
or U2231 (N_2231,N_1918,In_761);
or U2232 (N_2232,N_1359,N_1079);
and U2233 (N_2233,In_833,N_1945);
nor U2234 (N_2234,N_1386,N_1172);
nor U2235 (N_2235,N_1557,N_61);
xnor U2236 (N_2236,In_4014,In_1292);
and U2237 (N_2237,In_3462,N_1977);
nand U2238 (N_2238,In_1660,In_3128);
nand U2239 (N_2239,In_693,N_1572);
or U2240 (N_2240,In_2884,In_802);
nor U2241 (N_2241,N_950,In_1957);
or U2242 (N_2242,In_3872,N_1273);
nand U2243 (N_2243,N_841,In_1197);
or U2244 (N_2244,N_1827,In_3401);
nand U2245 (N_2245,N_311,In_3524);
nand U2246 (N_2246,N_1814,In_4107);
and U2247 (N_2247,In_2598,N_1114);
xor U2248 (N_2248,N_1462,In_110);
and U2249 (N_2249,N_1210,In_2973);
and U2250 (N_2250,In_1459,N_1709);
nand U2251 (N_2251,In_866,N_1307);
nand U2252 (N_2252,N_1524,In_3756);
nand U2253 (N_2253,In_15,In_341);
or U2254 (N_2254,N_1602,N_393);
and U2255 (N_2255,N_218,In_4685);
or U2256 (N_2256,In_3085,N_511);
or U2257 (N_2257,In_326,N_1115);
nand U2258 (N_2258,N_1698,N_568);
xor U2259 (N_2259,N_1242,In_3388);
nand U2260 (N_2260,In_1827,N_1040);
and U2261 (N_2261,N_459,In_2708);
and U2262 (N_2262,In_1525,N_63);
or U2263 (N_2263,N_633,N_1997);
xor U2264 (N_2264,N_1775,In_3110);
and U2265 (N_2265,In_4946,N_1525);
xor U2266 (N_2266,N_1492,In_652);
and U2267 (N_2267,In_675,N_1421);
and U2268 (N_2268,N_1779,In_3886);
nor U2269 (N_2269,N_1412,N_1801);
xnor U2270 (N_2270,N_394,N_76);
and U2271 (N_2271,N_1335,In_287);
and U2272 (N_2272,In_2234,In_3182);
or U2273 (N_2273,N_380,In_2770);
nor U2274 (N_2274,In_1183,N_49);
nor U2275 (N_2275,In_743,N_1218);
xnor U2276 (N_2276,N_1204,N_466);
nor U2277 (N_2277,N_254,N_279);
xor U2278 (N_2278,N_1020,In_3363);
nor U2279 (N_2279,N_1409,In_320);
xor U2280 (N_2280,N_1022,In_3158);
and U2281 (N_2281,N_848,N_737);
nand U2282 (N_2282,In_3167,In_4838);
or U2283 (N_2283,N_1294,In_2056);
and U2284 (N_2284,In_870,N_1308);
and U2285 (N_2285,N_110,N_1831);
and U2286 (N_2286,In_592,N_1228);
xnor U2287 (N_2287,N_791,N_1201);
and U2288 (N_2288,N_1763,N_1757);
nand U2289 (N_2289,N_1886,In_864);
and U2290 (N_2290,N_1889,N_1066);
xor U2291 (N_2291,In_1971,N_1690);
or U2292 (N_2292,N_1747,In_878);
xnor U2293 (N_2293,N_1562,N_1834);
nor U2294 (N_2294,N_366,In_1064);
xor U2295 (N_2295,N_895,In_1756);
or U2296 (N_2296,N_977,N_1219);
and U2297 (N_2297,In_2803,N_1392);
nand U2298 (N_2298,N_1870,In_448);
nor U2299 (N_2299,N_1071,N_1950);
nor U2300 (N_2300,N_1148,N_1039);
and U2301 (N_2301,N_1062,In_4868);
nand U2302 (N_2302,In_4036,In_1771);
nand U2303 (N_2303,N_1283,In_830);
nand U2304 (N_2304,In_2942,N_1567);
nor U2305 (N_2305,In_1500,N_792);
nor U2306 (N_2306,N_1028,In_3195);
and U2307 (N_2307,In_90,In_764);
xnor U2308 (N_2308,N_836,In_2808);
or U2309 (N_2309,In_1777,In_4388);
nand U2310 (N_2310,In_3259,In_3435);
or U2311 (N_2311,N_1326,In_4332);
and U2312 (N_2312,N_1838,N_1682);
and U2313 (N_2313,In_4774,N_1961);
and U2314 (N_2314,In_910,N_776);
and U2315 (N_2315,N_1005,In_2055);
nor U2316 (N_2316,N_928,In_3193);
nand U2317 (N_2317,In_552,N_1327);
nand U2318 (N_2318,N_1387,In_3082);
and U2319 (N_2319,In_4691,N_1966);
xor U2320 (N_2320,N_820,N_983);
and U2321 (N_2321,In_3350,N_1738);
or U2322 (N_2322,N_1406,N_7);
nor U2323 (N_2323,N_445,N_1182);
nand U2324 (N_2324,N_1999,In_4055);
nand U2325 (N_2325,N_271,In_952);
and U2326 (N_2326,In_813,In_4670);
nor U2327 (N_2327,N_402,In_653);
nand U2328 (N_2328,N_906,In_1573);
and U2329 (N_2329,N_1290,N_1688);
nand U2330 (N_2330,N_520,In_4968);
xor U2331 (N_2331,In_1530,N_1759);
nor U2332 (N_2332,N_1457,N_1969);
nand U2333 (N_2333,In_1787,In_2342);
xnor U2334 (N_2334,In_1129,In_4293);
xnor U2335 (N_2335,In_2537,In_1846);
and U2336 (N_2336,N_1536,N_232);
nor U2337 (N_2337,N_140,N_1670);
nand U2338 (N_2338,In_4894,In_2139);
xnor U2339 (N_2339,N_1681,N_1560);
and U2340 (N_2340,N_1828,N_1128);
or U2341 (N_2341,N_1211,N_1196);
nor U2342 (N_2342,N_900,In_1397);
or U2343 (N_2343,In_3760,N_1112);
xor U2344 (N_2344,N_224,N_1351);
nand U2345 (N_2345,In_1807,N_1144);
nand U2346 (N_2346,N_373,In_3726);
and U2347 (N_2347,N_1443,In_625);
or U2348 (N_2348,N_1098,N_1830);
nand U2349 (N_2349,N_1026,N_1174);
xnor U2350 (N_2350,N_671,In_4123);
and U2351 (N_2351,N_1037,N_1317);
nand U2352 (N_2352,N_1912,In_2469);
or U2353 (N_2353,In_2158,In_3100);
and U2354 (N_2354,In_4525,N_1667);
or U2355 (N_2355,In_4905,In_3974);
or U2356 (N_2356,N_148,In_1544);
nand U2357 (N_2357,N_1483,In_523);
and U2358 (N_2358,N_882,In_3043);
nand U2359 (N_2359,N_1901,In_4356);
nor U2360 (N_2360,N_929,N_1648);
nand U2361 (N_2361,N_1215,N_90);
or U2362 (N_2362,N_719,In_3721);
nand U2363 (N_2363,N_1319,N_1815);
xor U2364 (N_2364,N_1915,In_996);
xnor U2365 (N_2365,In_4370,In_1977);
or U2366 (N_2366,N_777,In_4879);
nor U2367 (N_2367,N_334,In_791);
xor U2368 (N_2368,In_1241,In_3976);
or U2369 (N_2369,In_3142,N_1162);
or U2370 (N_2370,N_1137,N_1506);
nor U2371 (N_2371,N_333,N_1168);
and U2372 (N_2372,N_1175,In_2763);
and U2373 (N_2373,N_1561,In_114);
nor U2374 (N_2374,In_2992,N_1744);
nor U2375 (N_2375,In_4486,N_853);
xor U2376 (N_2376,In_3492,N_1745);
nand U2377 (N_2377,N_1127,N_1729);
or U2378 (N_2378,In_1621,In_689);
xor U2379 (N_2379,In_3450,In_1725);
nand U2380 (N_2380,In_1353,In_1488);
xor U2381 (N_2381,In_1961,In_3539);
xnor U2382 (N_2382,N_1722,In_2366);
nand U2383 (N_2383,N_1503,In_1466);
nor U2384 (N_2384,N_1342,In_4693);
nand U2385 (N_2385,N_1282,N_198);
nand U2386 (N_2386,N_1391,In_29);
xnor U2387 (N_2387,In_2642,In_2546);
and U2388 (N_2388,N_1819,N_399);
or U2389 (N_2389,N_1160,N_1568);
and U2390 (N_2390,N_1708,N_40);
nand U2391 (N_2391,In_2866,N_1586);
xor U2392 (N_2392,In_3667,N_1873);
nand U2393 (N_2393,N_400,In_1737);
nand U2394 (N_2394,N_1456,In_221);
and U2395 (N_2395,N_1979,In_4051);
xor U2396 (N_2396,In_1650,In_3081);
nand U2397 (N_2397,In_4209,In_3113);
nor U2398 (N_2398,In_3040,N_703);
nand U2399 (N_2399,In_383,N_1006);
and U2400 (N_2400,N_1145,N_1723);
nand U2401 (N_2401,In_105,N_1555);
and U2402 (N_2402,N_766,In_3039);
nor U2403 (N_2403,N_938,N_1403);
nand U2404 (N_2404,N_1496,N_1277);
nand U2405 (N_2405,N_680,In_964);
xor U2406 (N_2406,N_1719,In_2317);
or U2407 (N_2407,In_2214,N_1305);
and U2408 (N_2408,N_1415,In_3032);
and U2409 (N_2409,N_1844,In_1995);
or U2410 (N_2410,In_1232,In_2176);
nor U2411 (N_2411,In_1902,In_3650);
or U2412 (N_2412,N_1849,N_943);
and U2413 (N_2413,N_79,N_1742);
nor U2414 (N_2414,N_1897,In_237);
nand U2415 (N_2415,In_3486,N_1832);
and U2416 (N_2416,In_4634,N_1377);
nand U2417 (N_2417,In_3472,N_97);
or U2418 (N_2418,N_1699,N_1113);
or U2419 (N_2419,N_1967,N_1905);
or U2420 (N_2420,In_2771,N_109);
nand U2421 (N_2421,N_1048,N_475);
or U2422 (N_2422,N_1038,In_1653);
xor U2423 (N_2423,In_4677,N_1970);
or U2424 (N_2424,N_1176,N_485);
or U2425 (N_2425,In_2786,N_1736);
xor U2426 (N_2426,N_1884,N_58);
nand U2427 (N_2427,In_3977,In_1369);
nor U2428 (N_2428,N_1974,In_4152);
xor U2429 (N_2429,In_1821,N_1631);
nand U2430 (N_2430,N_941,In_3550);
or U2431 (N_2431,In_1881,N_708);
xor U2432 (N_2432,N_645,In_4664);
nor U2433 (N_2433,N_1437,N_1139);
nand U2434 (N_2434,N_46,N_1766);
nand U2435 (N_2435,N_1206,N_1907);
or U2436 (N_2436,N_1208,N_627);
nand U2437 (N_2437,In_2429,In_1799);
nand U2438 (N_2438,N_1089,In_4305);
or U2439 (N_2439,N_239,In_2447);
nor U2440 (N_2440,N_372,N_1300);
nand U2441 (N_2441,In_2483,N_1778);
and U2442 (N_2442,N_555,N_1051);
or U2443 (N_2443,In_2041,In_2117);
nand U2444 (N_2444,N_1951,N_1414);
or U2445 (N_2445,In_475,In_3710);
or U2446 (N_2446,In_2718,In_2705);
nor U2447 (N_2447,N_728,N_1847);
or U2448 (N_2448,N_592,N_779);
xor U2449 (N_2449,N_1900,N_235);
or U2450 (N_2450,In_4655,N_1468);
and U2451 (N_2451,N_815,N_1425);
nand U2452 (N_2452,N_538,N_1680);
or U2453 (N_2453,In_1505,N_1780);
nor U2454 (N_2454,N_1750,In_3647);
xnor U2455 (N_2455,In_3301,N_1922);
or U2456 (N_2456,In_2739,N_517);
nand U2457 (N_2457,N_1297,In_2404);
xor U2458 (N_2458,In_20,N_830);
xor U2459 (N_2459,N_1546,In_3274);
nand U2460 (N_2460,In_3930,N_1612);
xnor U2461 (N_2461,N_1908,N_1802);
or U2462 (N_2462,In_826,In_2801);
nor U2463 (N_2463,N_1500,In_438);
or U2464 (N_2464,In_4400,In_337);
and U2465 (N_2465,N_1826,N_1685);
or U2466 (N_2466,In_4773,N_1029);
or U2467 (N_2467,In_2031,N_1240);
nand U2468 (N_2468,In_2257,N_571);
nand U2469 (N_2469,In_777,In_2924);
or U2470 (N_2470,In_1552,In_1871);
xnor U2471 (N_2471,N_919,N_1459);
or U2472 (N_2472,N_1380,N_1011);
and U2473 (N_2473,In_2707,In_1445);
or U2474 (N_2474,N_1479,In_4793);
nor U2475 (N_2475,N_436,N_1931);
or U2476 (N_2476,N_1932,In_186);
xor U2477 (N_2477,In_4738,In_2231);
and U2478 (N_2478,N_915,N_1485);
nor U2479 (N_2479,In_4494,N_1947);
xor U2480 (N_2480,In_670,N_1050);
nand U2481 (N_2481,N_1000,In_4843);
nor U2482 (N_2482,N_312,In_4243);
xnor U2483 (N_2483,In_2221,N_1985);
and U2484 (N_2484,N_1436,In_1448);
and U2485 (N_2485,N_250,In_4463);
or U2486 (N_2486,In_4438,In_3670);
or U2487 (N_2487,N_637,N_1746);
or U2488 (N_2488,N_1668,In_2758);
or U2489 (N_2489,In_402,N_1696);
xnor U2490 (N_2490,In_4225,N_177);
xnor U2491 (N_2491,N_1531,In_1098);
and U2492 (N_2492,In_4050,In_1724);
and U2493 (N_2493,N_910,N_1121);
nor U2494 (N_2494,N_1776,N_1057);
xor U2495 (N_2495,In_4536,N_1150);
nand U2496 (N_2496,N_1259,In_2585);
nor U2497 (N_2497,In_4299,In_3355);
xor U2498 (N_2498,N_384,In_4809);
xor U2499 (N_2499,N_1534,In_578);
xor U2500 (N_2500,N_1035,N_1078);
nand U2501 (N_2501,N_726,N_1702);
and U2502 (N_2502,In_1574,In_3147);
nor U2503 (N_2503,N_263,N_816);
and U2504 (N_2504,In_2491,N_435);
nand U2505 (N_2505,In_4415,N_684);
and U2506 (N_2506,In_409,In_947);
nand U2507 (N_2507,In_3298,In_2408);
and U2508 (N_2508,In_1478,N_1795);
nand U2509 (N_2509,N_1641,N_809);
or U2510 (N_2510,N_1771,N_1535);
or U2511 (N_2511,N_799,N_179);
and U2512 (N_2512,In_4807,In_2397);
xor U2513 (N_2513,N_1323,In_935);
nand U2514 (N_2514,In_3526,In_3933);
and U2515 (N_2515,In_4210,N_1677);
xor U2516 (N_2516,N_4,In_4201);
xor U2517 (N_2517,In_2952,N_1200);
nor U2518 (N_2518,N_1455,In_2185);
nor U2519 (N_2519,In_4465,N_325);
nand U2520 (N_2520,N_1023,N_1621);
nor U2521 (N_2521,In_3926,In_3272);
xor U2522 (N_2522,In_4514,N_887);
and U2523 (N_2523,N_1803,In_47);
xnor U2524 (N_2524,N_1820,In_2489);
xor U2525 (N_2525,N_546,In_222);
nor U2526 (N_2526,N_1340,N_1574);
or U2527 (N_2527,N_1116,N_233);
and U2528 (N_2528,In_986,In_2263);
xnor U2529 (N_2529,N_1163,In_3794);
or U2530 (N_2530,In_485,In_815);
nor U2531 (N_2531,In_1768,In_2940);
or U2532 (N_2532,N_1615,In_4231);
nor U2533 (N_2533,N_397,N_1314);
or U2534 (N_2534,In_4962,In_1890);
nor U2535 (N_2535,N_1402,In_2285);
xor U2536 (N_2536,In_33,In_4247);
nand U2537 (N_2537,In_442,In_3159);
and U2538 (N_2538,In_769,N_509);
or U2539 (N_2539,N_1734,N_221);
nand U2540 (N_2540,In_1096,In_2443);
nand U2541 (N_2541,N_1368,In_2425);
xor U2542 (N_2542,In_1072,In_4330);
nor U2543 (N_2543,N_1235,N_1254);
or U2544 (N_2544,In_2132,N_441);
and U2545 (N_2545,In_4850,N_1752);
nor U2546 (N_2546,N_529,In_579);
nor U2547 (N_2547,In_3386,N_270);
and U2548 (N_2548,In_1591,N_324);
nor U2549 (N_2549,In_1482,N_230);
nand U2550 (N_2550,N_192,N_1309);
xor U2551 (N_2551,In_1393,In_2680);
nor U2552 (N_2552,N_1142,N_1013);
and U2553 (N_2553,N_1100,N_1302);
xnor U2554 (N_2554,N_1543,In_3102);
or U2555 (N_2555,N_1054,N_1186);
nor U2556 (N_2556,N_1385,N_317);
nor U2557 (N_2557,In_1218,In_2606);
or U2558 (N_2558,In_1923,N_1528);
or U2559 (N_2559,N_1059,N_602);
or U2560 (N_2560,N_878,In_4556);
or U2561 (N_2561,In_1582,In_3296);
and U2562 (N_2562,In_464,N_1264);
xnor U2563 (N_2563,In_4108,N_1786);
and U2564 (N_2564,In_857,In_4936);
and U2565 (N_2565,N_1171,N_1509);
nand U2566 (N_2566,In_2390,In_1113);
or U2567 (N_2567,In_2985,In_1989);
nand U2568 (N_2568,N_1577,In_2617);
nand U2569 (N_2569,In_4958,N_184);
xnor U2570 (N_2570,N_831,N_1949);
nand U2571 (N_2571,N_1271,N_439);
and U2572 (N_2572,In_2584,N_1195);
xor U2573 (N_2573,In_2265,In_2188);
or U2574 (N_2574,N_35,In_836);
or U2575 (N_2575,In_2146,N_1626);
nand U2576 (N_2576,In_142,N_261);
and U2577 (N_2577,N_104,N_1484);
or U2578 (N_2578,N_695,N_1637);
nand U2579 (N_2579,In_1535,In_4136);
and U2580 (N_2580,In_720,N_1245);
nand U2581 (N_2581,N_1378,N_344);
nand U2582 (N_2582,In_3084,N_1032);
xor U2583 (N_2583,N_405,In_3252);
xnor U2584 (N_2584,N_1645,N_1512);
nor U2585 (N_2585,N_300,N_151);
nand U2586 (N_2586,N_1397,In_568);
and U2587 (N_2587,In_3734,In_2183);
and U2588 (N_2588,In_3026,N_1197);
xor U2589 (N_2589,N_1613,N_1604);
xnor U2590 (N_2590,In_517,In_4191);
xnor U2591 (N_2591,N_1143,In_4877);
nand U2592 (N_2592,In_1070,In_846);
nor U2593 (N_2593,N_837,In_2460);
xor U2594 (N_2594,In_286,N_1337);
nor U2595 (N_2595,N_1474,N_30);
or U2596 (N_2596,In_3631,In_3770);
nand U2597 (N_2597,In_1099,N_1096);
and U2598 (N_2598,In_1442,N_1043);
or U2599 (N_2599,In_1833,In_2228);
nor U2600 (N_2600,N_1646,N_1487);
nor U2601 (N_2601,In_4980,N_48);
and U2602 (N_2602,In_1629,In_979);
xor U2603 (N_2603,N_1903,In_4571);
or U2604 (N_2604,N_1181,N_1992);
nand U2605 (N_2605,N_1379,In_907);
or U2606 (N_2606,N_784,N_1823);
and U2607 (N_2607,In_3322,In_1794);
xnor U2608 (N_2608,In_107,N_654);
or U2609 (N_2609,In_958,In_3517);
nor U2610 (N_2610,N_634,In_650);
and U2611 (N_2611,N_1721,In_2655);
nand U2612 (N_2612,N_1471,In_4816);
xor U2613 (N_2613,N_1374,N_1291);
or U2614 (N_2614,In_1144,In_1471);
xnor U2615 (N_2615,N_702,In_696);
or U2616 (N_2616,N_1097,In_4095);
and U2617 (N_2617,N_155,In_3846);
xor U2618 (N_2618,N_448,In_1392);
nand U2619 (N_2619,N_1948,N_1643);
nor U2620 (N_2620,N_338,In_2754);
xor U2621 (N_2621,N_245,In_397);
xor U2622 (N_2622,N_1581,N_432);
and U2623 (N_2623,In_4810,In_1415);
nand U2624 (N_2624,N_1251,In_526);
nor U2625 (N_2625,In_398,N_39);
and U2626 (N_2626,In_111,In_1943);
and U2627 (N_2627,N_1151,N_1463);
xor U2628 (N_2628,N_1045,N_1784);
or U2629 (N_2629,N_1452,N_131);
and U2630 (N_2630,N_1935,In_137);
and U2631 (N_2631,N_1345,In_3122);
nand U2632 (N_2632,In_385,N_1260);
nand U2633 (N_2633,In_3996,N_1926);
xnor U2634 (N_2634,N_465,In_92);
and U2635 (N_2635,In_1670,In_1575);
xor U2636 (N_2636,N_694,In_3938);
or U2637 (N_2637,In_3510,In_1897);
or U2638 (N_2638,N_74,N_117);
and U2639 (N_2639,In_2689,In_3127);
or U2640 (N_2640,N_1275,N_1599);
or U2641 (N_2641,N_1848,In_2516);
or U2642 (N_2642,In_458,In_4493);
xor U2643 (N_2643,In_3680,In_4119);
nand U2644 (N_2644,N_1285,In_3859);
xor U2645 (N_2645,N_102,In_3862);
nor U2646 (N_2646,In_68,N_1178);
xor U2647 (N_2647,N_860,In_88);
xnor U2648 (N_2648,In_4922,N_1713);
and U2649 (N_2649,In_2922,In_1508);
nand U2650 (N_2650,N_1203,In_1882);
nor U2651 (N_2651,In_3228,In_4280);
nor U2652 (N_2652,N_347,In_2611);
nand U2653 (N_2653,N_998,In_3041);
xnor U2654 (N_2654,N_1707,N_1566);
or U2655 (N_2655,N_204,N_750);
xnor U2656 (N_2656,N_1140,N_1193);
nand U2657 (N_2657,In_2017,In_506);
nor U2658 (N_2658,In_407,In_4595);
nor U2659 (N_2659,In_4035,N_1867);
nand U2660 (N_2660,In_1868,In_175);
or U2661 (N_2661,In_1572,In_1779);
or U2662 (N_2662,In_2369,In_3634);
nor U2663 (N_2663,N_947,In_1410);
or U2664 (N_2664,N_1527,N_1434);
nand U2665 (N_2665,N_1548,N_176);
nor U2666 (N_2666,In_1260,In_1678);
and U2667 (N_2667,In_4885,N_174);
xor U2668 (N_2668,N_985,In_2908);
nand U2669 (N_2669,In_3107,In_2374);
and U2670 (N_2670,N_1504,N_1180);
nand U2671 (N_2671,In_1680,In_40);
nor U2672 (N_2672,N_1470,In_1389);
nand U2673 (N_2673,In_2168,In_298);
xnor U2674 (N_2674,N_1448,N_1904);
and U2675 (N_2675,In_4798,N_1694);
nand U2676 (N_2676,In_4351,N_1691);
and U2677 (N_2677,In_3321,N_157);
and U2678 (N_2678,N_1505,In_954);
or U2679 (N_2679,N_1617,N_843);
xnor U2680 (N_2680,N_1906,N_1980);
or U2681 (N_2681,N_1105,N_1895);
nand U2682 (N_2682,N_1518,In_3654);
nor U2683 (N_2683,In_4609,N_1395);
and U2684 (N_2684,N_1188,In_3812);
and U2685 (N_2685,In_1792,In_4897);
and U2686 (N_2686,In_2926,In_3633);
and U2687 (N_2687,N_1094,N_1659);
nor U2688 (N_2688,In_1423,N_60);
xnor U2689 (N_2689,In_2018,N_1214);
nor U2690 (N_2690,N_51,N_1711);
nor U2691 (N_2691,N_1808,N_1272);
or U2692 (N_2692,In_581,In_4286);
xor U2693 (N_2693,N_195,In_695);
nor U2694 (N_2694,N_1996,N_1450);
and U2695 (N_2695,In_3446,In_3283);
nand U2696 (N_2696,In_270,In_3352);
xnor U2697 (N_2697,In_934,In_1743);
or U2698 (N_2698,In_2871,In_257);
and U2699 (N_2699,In_514,N_744);
and U2700 (N_2700,In_4680,N_507);
xor U2701 (N_2701,In_515,In_3744);
nand U2702 (N_2702,In_4064,N_1055);
or U2703 (N_2703,N_597,In_2569);
nor U2704 (N_2704,In_1532,N_1511);
nand U2705 (N_2705,In_3844,In_953);
nor U2706 (N_2706,In_940,In_2070);
or U2707 (N_2707,In_3434,In_4538);
xnor U2708 (N_2708,N_1324,In_387);
or U2709 (N_2709,In_950,N_525);
or U2710 (N_2710,In_936,In_1608);
nor U2711 (N_2711,In_4829,N_1672);
xnor U2712 (N_2712,N_1710,N_322);
and U2713 (N_2713,N_288,N_1570);
or U2714 (N_2714,N_1124,N_1173);
and U2715 (N_2715,N_925,N_1356);
nor U2716 (N_2716,In_4568,In_1837);
nand U2717 (N_2717,N_33,N_1517);
and U2718 (N_2718,In_4266,N_1872);
nor U2719 (N_2719,N_569,In_3027);
nand U2720 (N_2720,N_1316,N_807);
or U2721 (N_2721,In_3765,N_1629);
nor U2722 (N_2722,In_1050,In_2929);
nor U2723 (N_2723,In_2962,N_107);
nand U2724 (N_2724,In_4188,In_1628);
nand U2725 (N_2725,In_241,In_988);
nand U2726 (N_2726,N_164,In_3280);
nand U2727 (N_2727,In_1312,In_1546);
nor U2728 (N_2728,N_1946,N_554);
nand U2729 (N_2729,In_2684,N_620);
nor U2730 (N_2730,In_3664,N_1068);
nor U2731 (N_2731,N_1021,In_4453);
or U2732 (N_2732,In_501,In_1681);
nand U2733 (N_2733,N_1928,N_1751);
and U2734 (N_2734,In_1847,In_2341);
xor U2735 (N_2735,In_2329,In_1537);
and U2736 (N_2736,In_170,In_2890);
nand U2737 (N_2737,In_806,In_404);
nand U2738 (N_2738,In_637,In_1599);
or U2739 (N_2739,In_3733,N_482);
xor U2740 (N_2740,N_71,N_1343);
and U2741 (N_2741,In_2745,In_1515);
xnor U2742 (N_2742,N_711,In_1665);
xor U2743 (N_2743,N_672,In_265);
and U2744 (N_2744,In_72,N_1422);
nor U2745 (N_2745,N_1117,In_2381);
nand U2746 (N_2746,In_3688,N_1401);
nand U2747 (N_2747,N_1594,In_2967);
xnor U2748 (N_2748,N_675,N_1217);
or U2749 (N_2749,N_966,In_3545);
or U2750 (N_2750,In_3461,N_82);
and U2751 (N_2751,N_1730,N_663);
and U2752 (N_2752,N_1366,N_1199);
or U2753 (N_2753,In_1481,N_1288);
xor U2754 (N_2754,N_710,In_4058);
xor U2755 (N_2755,In_3513,N_1119);
and U2756 (N_2756,N_1070,In_4138);
nand U2757 (N_2757,N_1318,In_1939);
xnor U2758 (N_2758,N_1253,In_3403);
or U2759 (N_2759,In_4366,N_512);
or U2760 (N_2760,In_718,In_2115);
xnor U2761 (N_2761,N_980,N_85);
or U2762 (N_2762,N_1754,In_2156);
and U2763 (N_2763,N_1301,In_131);
nor U2764 (N_2764,In_2541,N_1507);
nor U2765 (N_2765,N_1490,In_38);
xor U2766 (N_2766,N_1758,In_832);
nand U2767 (N_2767,In_4795,In_3454);
and U2768 (N_2768,In_324,N_1278);
xnor U2769 (N_2769,N_1770,N_1793);
xnor U2770 (N_2770,N_1060,In_488);
and U2771 (N_2771,N_1871,In_2485);
nand U2772 (N_2772,In_823,In_1870);
and U2773 (N_2773,In_1646,In_2448);
nand U2774 (N_2774,In_1164,In_628);
xor U2775 (N_2775,In_2118,In_3826);
or U2776 (N_2776,In_3778,N_562);
nand U2777 (N_2777,N_871,In_4737);
nand U2778 (N_2778,N_1249,In_824);
and U2779 (N_2779,N_1545,N_1082);
nand U2780 (N_2780,N_1878,In_4257);
nand U2781 (N_2781,N_1339,N_1125);
xor U2782 (N_2782,In_4683,In_2888);
xnor U2783 (N_2783,N_579,N_1811);
or U2784 (N_2784,In_3231,In_4478);
nand U2785 (N_2785,In_4765,In_1097);
xnor U2786 (N_2786,N_1303,In_4323);
nand U2787 (N_2787,In_2240,N_486);
nor U2788 (N_2788,In_3373,In_1775);
or U2789 (N_2789,N_1620,In_56);
nand U2790 (N_2790,In_1053,In_1362);
nand U2791 (N_2791,N_1306,In_223);
nor U2792 (N_2792,N_1675,In_3949);
nor U2793 (N_2793,N_735,N_64);
xor U2794 (N_2794,In_2947,N_1532);
nand U2795 (N_2795,In_229,In_3361);
and U2796 (N_2796,N_1890,N_1983);
and U2797 (N_2797,In_1330,In_3215);
nor U2798 (N_2798,N_1768,In_584);
nand U2799 (N_2799,In_1705,In_992);
and U2800 (N_2800,N_1441,N_1704);
or U2801 (N_2801,N_428,N_1649);
or U2802 (N_2802,In_1304,In_744);
nand U2803 (N_2803,In_1172,In_3366);
nor U2804 (N_2804,N_1537,N_1229);
or U2805 (N_2805,In_2376,In_2733);
nor U2806 (N_2806,N_912,N_1348);
and U2807 (N_2807,N_1787,N_1782);
nand U2808 (N_2808,In_3325,In_3009);
and U2809 (N_2809,N_55,In_2138);
and U2810 (N_2810,N_81,In_1880);
xnor U2811 (N_2811,N_1635,N_1822);
or U2812 (N_2812,N_1464,In_4001);
nand U2813 (N_2813,In_1733,N_1187);
xor U2814 (N_2814,N_1413,N_1274);
nand U2815 (N_2815,In_2345,N_13);
or U2816 (N_2816,N_622,In_2669);
and U2817 (N_2817,In_193,In_1580);
xor U2818 (N_2818,In_4218,In_4161);
or U2819 (N_2819,N_662,N_922);
nand U2820 (N_2820,In_2826,N_1625);
or U2821 (N_2821,N_1944,In_706);
and U2822 (N_2822,In_135,In_2998);
and U2823 (N_2823,In_234,In_3145);
nor U2824 (N_2824,In_4467,N_1072);
xor U2825 (N_2825,In_3840,N_1800);
or U2826 (N_2826,In_1166,N_1902);
or U2827 (N_2827,In_1786,In_4090);
xnor U2828 (N_2828,N_1213,N_141);
nand U2829 (N_2829,N_1875,In_1081);
or U2830 (N_2830,N_974,In_3118);
and U2831 (N_2831,In_2277,N_37);
nand U2832 (N_2832,In_483,In_3535);
or U2833 (N_2833,N_742,In_3567);
or U2834 (N_2834,In_1948,In_2107);
nand U2835 (N_2835,N_1295,In_2331);
and U2836 (N_2836,N_1666,N_1558);
xnor U2837 (N_2837,In_2294,In_3755);
or U2838 (N_2838,N_1899,N_1170);
and U2839 (N_2839,In_1383,N_1015);
nand U2840 (N_2840,N_1836,In_4130);
and U2841 (N_2841,N_243,N_1597);
or U2842 (N_2842,N_1236,In_4748);
or U2843 (N_2843,In_1408,N_1671);
nand U2844 (N_2844,N_149,In_1713);
nor U2845 (N_2845,In_1501,In_3442);
xor U2846 (N_2846,N_1353,N_542);
and U2847 (N_2847,N_1583,In_4610);
nand U2848 (N_2848,In_1276,N_1265);
or U2849 (N_2849,N_248,In_2910);
xnor U2850 (N_2850,N_1988,In_3240);
nor U2851 (N_2851,N_1322,N_1952);
nand U2852 (N_2852,In_3745,N_93);
nor U2853 (N_2853,N_1606,In_4918);
nor U2854 (N_2854,N_44,N_1683);
and U2855 (N_2855,N_1185,In_1850);
nor U2856 (N_2856,In_796,In_767);
or U2857 (N_2857,N_1909,N_1102);
or U2858 (N_2858,N_231,In_1509);
xor U2859 (N_2859,In_1726,In_1822);
nand U2860 (N_2860,N_1600,N_976);
or U2861 (N_2861,N_1898,N_1212);
and U2862 (N_2862,In_3759,In_1409);
xor U2863 (N_2863,In_881,In_2545);
or U2864 (N_2864,N_1638,N_1442);
and U2865 (N_2865,In_2088,In_3055);
xnor U2866 (N_2866,N_937,In_1382);
xor U2867 (N_2867,In_2529,N_1149);
nand U2868 (N_2868,N_303,N_331);
nand U2869 (N_2869,N_73,In_1593);
xnor U2870 (N_2870,In_638,N_524);
and U2871 (N_2871,In_75,In_3531);
or U2872 (N_2872,In_4733,N_1276);
or U2873 (N_2873,N_1933,In_2944);
or U2874 (N_2874,In_814,N_1611);
and U2875 (N_2875,In_4666,N_1310);
xnor U2876 (N_2876,In_1319,N_873);
xnor U2877 (N_2877,In_1068,In_322);
nor U2878 (N_2878,In_3372,In_4464);
and U2879 (N_2879,N_954,N_1154);
and U2880 (N_2880,N_1733,N_1269);
or U2881 (N_2881,In_2187,N_1376);
nor U2882 (N_2882,N_842,In_1314);
or U2883 (N_2883,In_1536,N_803);
or U2884 (N_2884,In_4533,N_1226);
and U2885 (N_2885,In_1909,N_185);
nor U2886 (N_2886,N_759,N_1762);
xor U2887 (N_2887,N_1647,N_896);
or U2888 (N_2888,N_1943,N_639);
nor U2889 (N_2889,In_4360,In_2014);
nor U2890 (N_2890,In_4674,N_519);
and U2891 (N_2891,N_16,In_4869);
nand U2892 (N_2892,N_95,In_546);
nor U2893 (N_2893,N_1410,N_1892);
or U2894 (N_2894,N_1879,In_3066);
or U2895 (N_2895,N_1080,N_1669);
or U2896 (N_2896,N_1603,In_805);
and U2897 (N_2897,In_210,In_4706);
and U2898 (N_2898,N_619,In_4705);
nand U2899 (N_2899,N_458,In_3238);
and U2900 (N_2900,N_503,N_1111);
xnor U2901 (N_2901,In_3443,N_829);
nand U2902 (N_2902,In_1086,In_3527);
or U2903 (N_2903,N_1530,In_1256);
and U2904 (N_2904,N_1773,In_1185);
nand U2905 (N_2905,In_2062,N_1230);
nor U2906 (N_2906,In_2648,In_1514);
xnor U2907 (N_2907,N_773,In_4518);
and U2908 (N_2908,N_753,N_208);
nand U2909 (N_2909,N_1093,In_1623);
nand U2910 (N_2910,N_427,In_596);
and U2911 (N_2911,In_1271,N_1136);
or U2912 (N_2912,N_227,N_1550);
xor U2913 (N_2913,In_2868,In_547);
nand U2914 (N_2914,N_1016,N_22);
or U2915 (N_2915,In_3222,In_76);
nor U2916 (N_2916,N_1279,N_577);
xnor U2917 (N_2917,In_2644,N_1104);
nor U2918 (N_2918,N_446,N_1888);
and U2919 (N_2919,In_3858,N_1589);
xnor U2920 (N_2920,In_2641,N_1418);
or U2921 (N_2921,N_1346,In_770);
xor U2922 (N_2922,In_3668,N_581);
nor U2923 (N_2923,N_864,In_926);
or U2924 (N_2924,N_1936,N_1585);
or U2925 (N_2925,In_4110,In_2249);
nand U2926 (N_2926,In_990,N_1417);
and U2927 (N_2927,N_973,N_1189);
and U2928 (N_2928,In_3890,In_2765);
nand U2929 (N_2929,In_2173,In_2872);
nor U2930 (N_2930,In_2348,In_2565);
xnor U2931 (N_2931,In_987,In_4148);
xor U2932 (N_2932,N_287,In_4528);
nor U2933 (N_2933,In_2891,In_1437);
nand U2934 (N_2934,In_82,In_4524);
nor U2935 (N_2935,N_822,N_1893);
nor U2936 (N_2936,N_1792,N_1304);
or U2937 (N_2937,N_1737,N_1542);
and U2938 (N_2938,N_1523,N_948);
and U2939 (N_2939,N_1268,In_4603);
xor U2940 (N_2940,In_2987,N_1538);
and U2941 (N_2941,N_1731,N_1693);
xor U2942 (N_2942,N_1856,N_1859);
nor U2943 (N_2943,In_2935,In_4623);
nand U2944 (N_2944,In_586,In_3809);
or U2945 (N_2945,N_687,N_1101);
nand U2946 (N_2946,In_1496,N_1458);
nand U2947 (N_2947,N_171,In_1914);
nand U2948 (N_2948,N_1717,N_1864);
xor U2949 (N_2949,N_376,N_1008);
or U2950 (N_2950,In_1266,In_3614);
xor U2951 (N_2951,N_1794,N_1202);
or U2952 (N_2952,N_260,In_562);
and U2953 (N_2953,N_352,N_739);
nor U2954 (N_2954,N_721,N_1616);
xnor U2955 (N_2955,N_518,N_1476);
and U2956 (N_2956,N_94,N_332);
nand U2957 (N_2957,In_4902,N_849);
or U2958 (N_2958,N_1580,In_2237);
xnor U2959 (N_2959,In_295,N_781);
nor U2960 (N_2960,In_4540,N_1598);
or U2961 (N_2961,N_1248,In_1764);
nand U2962 (N_2962,In_1433,N_1910);
nand U2963 (N_2963,In_2094,N_1553);
xor U2964 (N_2964,In_36,In_2172);
nand U2965 (N_2965,N_1394,N_1003);
nor U2966 (N_2966,In_1015,In_4031);
and U2967 (N_2967,N_962,N_426);
nor U2968 (N_2968,N_1718,N_1053);
xnor U2969 (N_2969,N_1161,In_4133);
nand U2970 (N_2970,N_1839,In_2038);
and U2971 (N_2971,In_603,N_716);
nand U2972 (N_2972,N_814,N_1965);
or U2973 (N_2973,N_1286,N_1311);
nand U2974 (N_2974,N_391,N_1400);
nor U2975 (N_2975,In_4767,In_2072);
and U2976 (N_2976,In_1231,N_1592);
nand U2977 (N_2977,In_2455,In_3910);
and U2978 (N_2978,N_1063,N_1595);
or U2979 (N_2979,N_1760,N_1460);
xnor U2980 (N_2980,In_4797,In_1927);
xor U2981 (N_2981,In_2691,In_3176);
and U2982 (N_2982,N_1076,N_1833);
xnor U2983 (N_2983,In_319,In_420);
and U2984 (N_2984,In_3180,N_857);
xor U2985 (N_2985,N_1516,In_1620);
nand U2986 (N_2986,N_1489,N_704);
nand U2987 (N_2987,N_736,In_4213);
nor U2988 (N_2988,N_1439,N_364);
and U2989 (N_2989,In_1487,In_2463);
nor U2990 (N_2990,In_1669,In_3160);
xor U2991 (N_2991,N_1398,N_1591);
xnor U2992 (N_2992,In_681,N_1074);
nand U2993 (N_2993,In_4496,In_277);
xor U2994 (N_2994,N_1636,In_903);
nor U2995 (N_2995,N_944,N_1103);
nand U2996 (N_2996,N_444,In_2931);
nand U2997 (N_2997,N_1083,In_430);
nor U2998 (N_2998,N_1370,In_3029);
or U2999 (N_2999,N_1360,In_373);
nor U3000 (N_3000,N_2481,In_3988);
xnor U3001 (N_3001,In_635,N_1712);
or U3002 (N_3002,N_2111,N_2020);
and U3003 (N_3003,N_2574,In_1840);
or U3004 (N_3004,N_2013,N_2681);
nor U3005 (N_3005,N_2402,N_2972);
xor U3006 (N_3006,N_1689,In_1019);
or U3007 (N_3007,N_960,N_2419);
nand U3008 (N_3008,N_626,N_2640);
or U3009 (N_3009,N_1767,N_2390);
and U3010 (N_3010,N_2517,N_1939);
nor U3011 (N_3011,N_2414,N_2473);
xnor U3012 (N_3012,N_1194,N_2825);
nand U3013 (N_3013,N_2172,N_360);
and U3014 (N_3014,In_1584,In_264);
nand U3015 (N_3015,N_1861,N_2137);
xnor U3016 (N_3016,N_1942,N_2675);
nor U3017 (N_3017,N_2154,In_3375);
or U3018 (N_3018,In_663,In_1400);
or U3019 (N_3019,In_1742,In_4714);
nor U3020 (N_3020,N_2794,N_2551);
nor U3021 (N_3021,In_968,N_2816);
and U3022 (N_3022,N_2082,In_3793);
or U3023 (N_3023,In_2568,In_4140);
nor U3024 (N_3024,N_1940,N_2889);
xnor U3025 (N_3025,N_1475,N_2294);
or U3026 (N_3026,N_1816,In_3273);
xnor U3027 (N_3027,N_2837,N_2429);
nand U3028 (N_3028,N_2593,N_2490);
or U3029 (N_3029,N_806,N_1081);
xnor U3030 (N_3030,N_787,N_2839);
xnor U3031 (N_3031,N_2325,N_2261);
or U3032 (N_3032,N_2477,In_4269);
xnor U3033 (N_3033,In_1615,In_104);
and U3034 (N_3034,N_2863,In_1416);
or U3035 (N_3035,N_1725,N_374);
and U3036 (N_3036,N_2973,N_105);
and U3037 (N_3037,N_2388,In_2895);
nor U3038 (N_3038,N_2712,N_1593);
and U3039 (N_3039,In_2624,N_2077);
and U3040 (N_3040,N_2401,In_3005);
nor U3041 (N_3041,N_2433,N_783);
or U3042 (N_3042,N_1357,N_1010);
and U3043 (N_3043,N_2416,In_738);
nand U3044 (N_3044,N_2190,In_150);
nor U3045 (N_3045,N_1817,N_2008);
or U3046 (N_3046,N_2443,N_2866);
nor U3047 (N_3047,N_1390,N_1030);
xor U3048 (N_3048,N_2649,N_2938);
nand U3049 (N_3049,In_956,N_244);
nand U3050 (N_3050,N_2377,N_2963);
nand U3051 (N_3051,In_4722,N_1652);
xnor U3052 (N_3052,N_1726,In_939);
or U3053 (N_3053,N_2102,N_2705);
nand U3054 (N_3054,N_2071,In_457);
xnor U3055 (N_3055,In_184,N_2186);
or U3056 (N_3056,N_2276,N_1192);
xor U3057 (N_3057,N_2731,N_2692);
and U3058 (N_3058,N_2363,N_2179);
nand U3059 (N_3059,N_2449,In_2817);
nand U3060 (N_3060,In_655,In_2743);
nand U3061 (N_3061,In_1972,In_1399);
or U3062 (N_3062,N_2515,N_1354);
xnor U3063 (N_3063,N_1735,In_3148);
and U3064 (N_3064,N_2607,N_2842);
and U3065 (N_3065,N_565,N_1913);
or U3066 (N_3066,N_2791,In_819);
or U3067 (N_3067,N_2903,N_1465);
and U3068 (N_3068,N_1042,N_1858);
xor U3069 (N_3069,N_2394,N_994);
and U3070 (N_3070,N_970,N_1255);
nand U3071 (N_3071,In_2953,N_2667);
and U3072 (N_3072,In_342,In_691);
nand U3073 (N_3073,N_407,In_1364);
nand U3074 (N_3074,N_2775,N_1454);
nand U3075 (N_3075,N_2312,N_2255);
nor U3076 (N_3076,N_1281,In_2420);
and U3077 (N_3077,N_1715,N_2764);
or U3078 (N_3078,In_2396,N_2003);
or U3079 (N_3079,N_2648,N_285);
nand U3080 (N_3080,N_2786,In_3408);
xnor U3081 (N_3081,N_1576,N_2941);
nand U3082 (N_3082,N_1420,In_2480);
xor U3083 (N_3083,N_2979,N_2254);
nor U3084 (N_3084,N_1041,N_1519);
and U3085 (N_3085,N_1184,N_2387);
xor U3086 (N_3086,N_2157,N_2208);
and U3087 (N_3087,In_4542,N_2766);
nand U3088 (N_3088,In_946,In_3857);
nand U3089 (N_3089,In_1056,In_3696);
xnor U3090 (N_3090,N_2026,N_2087);
xor U3091 (N_3091,N_2880,N_1854);
and U3092 (N_3092,N_1315,N_2730);
and U3093 (N_3093,N_2270,N_2760);
xor U3094 (N_3094,In_4402,N_2871);
xnor U3095 (N_3095,N_2501,N_1797);
xor U3096 (N_3096,N_2418,N_2537);
nand U3097 (N_3097,N_2439,N_1845);
and U3098 (N_3098,N_1547,N_1610);
and U3099 (N_3099,N_2400,In_3163);
nor U3100 (N_3100,In_3725,In_2148);
or U3101 (N_3101,N_2193,N_346);
xor U3102 (N_3102,N_2657,In_3371);
xor U3103 (N_3103,N_2030,N_2004);
nor U3104 (N_3104,N_2662,N_2788);
nor U3105 (N_3105,N_2006,N_1582);
or U3106 (N_3106,N_1881,N_2352);
and U3107 (N_3107,In_4425,N_2702);
or U3108 (N_3108,In_3678,N_2741);
nand U3109 (N_3109,N_1222,N_201);
or U3110 (N_3110,In_3955,In_2403);
or U3111 (N_3111,N_1325,N_2909);
nor U3112 (N_3112,N_2122,In_4200);
xnor U3113 (N_3113,N_2417,N_2398);
nand U3114 (N_3114,N_478,In_2057);
and U3115 (N_3115,N_1824,N_2344);
nor U3116 (N_3116,N_2762,N_2078);
or U3117 (N_3117,N_2868,N_1716);
or U3118 (N_3118,In_781,N_2001);
nand U3119 (N_3119,N_2559,N_1419);
nor U3120 (N_3120,In_312,In_3776);
nand U3121 (N_3121,N_2674,N_2497);
nand U3122 (N_3122,In_3241,N_1563);
xor U3123 (N_3123,N_2310,N_2425);
and U3124 (N_3124,N_1741,In_591);
or U3125 (N_3125,In_3011,N_2011);
nor U3126 (N_3126,N_1223,N_1978);
nand U3127 (N_3127,N_2059,In_392);
nor U3128 (N_3128,In_4577,N_2289);
xor U3129 (N_3129,In_3125,N_945);
nor U3130 (N_3130,In_1354,N_385);
xnor U3131 (N_3131,N_403,In_4959);
xor U3132 (N_3132,N_2703,N_2872);
nor U3133 (N_3133,N_2982,In_2677);
nor U3134 (N_3134,N_2132,In_4873);
nand U3135 (N_3135,N_2980,N_2733);
nor U3136 (N_3136,In_276,N_2295);
or U3137 (N_3137,In_3031,N_2984);
or U3138 (N_3138,N_2695,In_1007);
and U3139 (N_3139,N_2614,N_2052);
nand U3140 (N_3140,N_1469,In_1586);
nor U3141 (N_3141,In_1244,N_2850);
and U3142 (N_3142,N_2613,N_2396);
xor U3143 (N_3143,N_1772,N_2806);
and U3144 (N_3144,In_3120,N_813);
or U3145 (N_3145,N_1047,N_2765);
or U3146 (N_3146,N_2359,In_3772);
and U3147 (N_3147,In_4215,N_2879);
nor U3148 (N_3148,N_2736,In_4948);
or U3149 (N_3149,N_2829,N_1662);
and U3150 (N_3150,In_1080,N_2588);
nand U3151 (N_3151,N_934,In_3448);
or U3152 (N_3152,N_2911,N_921);
nor U3153 (N_3153,N_2891,N_2542);
nand U3154 (N_3154,N_2360,N_1369);
nand U3155 (N_3155,In_303,N_2426);
or U3156 (N_3156,N_386,N_1501);
nor U3157 (N_3157,N_1575,N_1877);
nor U3158 (N_3158,N_2287,N_940);
or U3159 (N_3159,N_593,In_2042);
xnor U3160 (N_3160,N_825,N_1075);
nor U3161 (N_3161,In_2098,In_725);
nand U3162 (N_3162,N_2203,In_4901);
nor U3163 (N_3163,N_2953,N_2841);
nor U3164 (N_3164,N_1642,N_2621);
nand U3165 (N_3165,N_2180,N_2992);
xnor U3166 (N_3166,N_1012,N_1289);
nor U3167 (N_3167,N_2809,N_2660);
nand U3168 (N_3168,In_492,N_1157);
xor U3169 (N_3169,N_1244,In_3342);
and U3170 (N_3170,N_2380,In_1823);
xnor U3171 (N_3171,N_2096,N_2063);
xor U3172 (N_3172,N_2256,N_2902);
xor U3173 (N_3173,In_3494,In_865);
xnor U3174 (N_3174,N_2466,N_2565);
xnor U3175 (N_3175,N_2707,In_2467);
nand U3176 (N_3176,N_2204,In_2251);
nor U3177 (N_3177,N_2442,N_2160);
nand U3178 (N_3178,N_1539,N_2822);
nor U3179 (N_3179,In_3421,N_550);
nand U3180 (N_3180,N_2091,N_2498);
and U3181 (N_3181,In_106,In_4662);
xnor U3182 (N_3182,N_2445,In_1052);
nor U3183 (N_3183,In_3479,N_1541);
nor U3184 (N_3184,N_992,In_3115);
and U3185 (N_3185,In_722,N_2409);
and U3186 (N_3186,N_800,N_1651);
xor U3187 (N_3187,N_383,N_2777);
xor U3188 (N_3188,N_2739,N_2321);
and U3189 (N_3189,In_2694,N_70);
nand U3190 (N_3190,N_1404,N_2696);
or U3191 (N_3191,In_2793,N_1256);
and U3192 (N_3192,N_2646,In_1450);
and U3193 (N_3193,In_2011,In_3931);
nor U3194 (N_3194,In_3423,In_540);
nand U3195 (N_3195,N_2309,N_790);
xor U3196 (N_3196,In_1006,N_2857);
nand U3197 (N_3197,N_1853,N_1165);
and U3198 (N_3198,N_2133,In_4027);
or U3199 (N_3199,N_2659,N_1655);
nor U3200 (N_3200,N_136,N_1488);
nand U3201 (N_3201,N_336,In_2422);
xnor U3202 (N_3202,N_1876,N_2487);
and U3203 (N_3203,N_2887,N_1874);
xnor U3204 (N_3204,N_2917,N_2427);
nor U3205 (N_3205,N_2751,N_2348);
nor U3206 (N_3206,N_2754,N_545);
nor U3207 (N_3207,N_431,N_2584);
or U3208 (N_3208,N_2688,In_228);
nor U3209 (N_3209,N_2625,N_247);
or U3210 (N_3210,N_1446,N_2556);
and U3211 (N_3211,N_2205,In_4358);
and U3212 (N_3212,N_2029,In_978);
or U3213 (N_3213,In_3947,N_2600);
nand U3214 (N_3214,N_2019,N_1665);
nor U3215 (N_3215,N_2906,N_2376);
nor U3216 (N_3216,In_1893,N_1953);
and U3217 (N_3217,In_3519,N_2301);
xor U3218 (N_3218,N_2399,N_2589);
nand U3219 (N_3219,In_419,In_3577);
and U3220 (N_3220,In_561,In_190);
xnor U3221 (N_3221,In_4546,N_1238);
nand U3222 (N_3222,N_2856,N_2238);
and U3223 (N_3223,N_2569,N_2511);
or U3224 (N_3224,N_2647,N_1449);
or U3225 (N_3225,N_2643,N_584);
xor U3226 (N_3226,N_2844,N_2934);
and U3227 (N_3227,N_2590,N_1258);
or U3228 (N_3228,N_2246,In_1261);
xnor U3229 (N_3229,In_4977,N_2357);
xnor U3230 (N_3230,N_2725,N_1850);
nand U3231 (N_3231,N_2127,N_1389);
nand U3232 (N_3232,N_2112,N_2074);
or U3233 (N_3233,N_1673,N_2368);
nor U3234 (N_3234,In_367,In_3456);
nand U3235 (N_3235,N_251,N_2025);
and U3236 (N_3236,In_3349,N_1564);
and U3237 (N_3237,N_2144,N_2790);
nor U3238 (N_3238,In_1157,N_2250);
nand U3239 (N_3239,N_72,N_2500);
nand U3240 (N_3240,N_1653,N_2770);
nor U3241 (N_3241,N_2056,N_1131);
nand U3242 (N_3242,N_419,N_163);
nor U3243 (N_3243,N_398,In_4219);
and U3244 (N_3244,N_1152,N_972);
or U3245 (N_3245,N_2252,N_2215);
nand U3246 (N_3246,N_1882,N_1084);
or U3247 (N_3247,In_3369,N_2420);
xnor U3248 (N_3248,N_2428,N_1919);
xnor U3249 (N_3249,N_2851,N_2039);
nor U3250 (N_3250,N_2704,N_2128);
xnor U3251 (N_3251,N_902,N_2499);
or U3252 (N_3252,In_3079,N_1365);
or U3253 (N_3253,N_2479,N_462);
xor U3254 (N_3254,In_2486,N_2612);
nor U3255 (N_3255,N_1695,N_1085);
nand U3256 (N_3256,N_2489,N_2966);
or U3257 (N_3257,N_2936,N_1614);
xor U3258 (N_3258,In_2200,N_87);
nor U3259 (N_3259,In_2571,In_3672);
nor U3260 (N_3260,N_210,N_2129);
nor U3261 (N_3261,N_1495,N_1777);
or U3262 (N_3262,N_166,N_1991);
xnor U3263 (N_3263,N_2905,In_2434);
xnor U3264 (N_3264,N_1077,N_2959);
nand U3265 (N_3265,In_872,N_2148);
and U3266 (N_3266,N_2230,N_2632);
nand U3267 (N_3267,N_2847,In_3035);
xor U3268 (N_3268,N_2010,N_2615);
nor U3269 (N_3269,In_1932,N_2768);
nor U3270 (N_3270,In_1083,In_4927);
and U3271 (N_3271,N_1533,In_2318);
xor U3272 (N_3272,N_2318,N_1493);
xnor U3273 (N_3273,N_2814,N_2969);
nand U3274 (N_3274,N_2828,N_2701);
nand U3275 (N_3275,In_3604,In_1132);
and U3276 (N_3276,N_2322,N_2159);
xor U3277 (N_3277,In_3181,N_1099);
nor U3278 (N_3278,In_1127,N_2535);
nand U3279 (N_3279,N_2073,In_1483);
nand U3280 (N_3280,In_1153,In_4799);
nor U3281 (N_3281,N_2840,N_2424);
and U3282 (N_3282,N_2478,N_1118);
xor U3283 (N_3283,N_1423,N_1262);
or U3284 (N_3284,N_2947,N_2916);
nand U3285 (N_3285,N_452,N_2224);
xnor U3286 (N_3286,In_1704,N_2991);
nor U3287 (N_3287,In_537,N_2221);
xnor U3288 (N_3288,N_1633,N_835);
and U3289 (N_3289,In_42,N_2308);
nor U3290 (N_3290,N_2366,In_1449);
nand U3291 (N_3291,N_2327,N_2534);
nand U3292 (N_3292,In_1040,N_1748);
and U3293 (N_3293,N_2738,In_759);
or U3294 (N_3294,In_698,N_1207);
xor U3295 (N_3295,N_2164,N_2552);
and U3296 (N_3296,In_1529,N_1549);
or U3297 (N_3297,In_3964,N_2470);
and U3298 (N_3298,N_2142,N_2198);
nand U3299 (N_3299,N_899,In_4981);
nor U3300 (N_3300,N_2329,N_876);
and U3301 (N_3301,N_2849,N_2624);
nand U3302 (N_3302,N_1521,In_2722);
or U3303 (N_3303,In_2419,In_227);
or U3304 (N_3304,In_1729,N_2838);
nor U3305 (N_3305,N_1280,N_2852);
xor U3306 (N_3306,N_2273,N_2507);
nor U3307 (N_3307,N_180,N_1578);
nor U3308 (N_3308,In_4660,N_2130);
nand U3309 (N_3309,N_2412,N_84);
and U3310 (N_3310,N_2407,In_2572);
nor U3311 (N_3311,N_327,N_2207);
or U3312 (N_3312,N_2661,N_2805);
or U3313 (N_3313,N_1292,N_2812);
nor U3314 (N_3314,N_850,N_1453);
nor U3315 (N_3315,N_2434,N_840);
nor U3316 (N_3316,N_2510,N_2286);
and U3317 (N_3317,In_1867,In_3993);
xnor U3318 (N_3318,In_1291,N_2283);
and U3319 (N_3319,N_2576,N_2898);
or U3320 (N_3320,N_2687,In_4056);
and U3321 (N_3321,N_2300,In_3284);
nand U3322 (N_3322,N_1433,N_2757);
or U3323 (N_3323,N_2910,N_2602);
or U3324 (N_3324,In_2988,N_2801);
nand U3325 (N_3325,N_2815,N_2663);
and U3326 (N_3326,N_1361,In_1784);
or U3327 (N_3327,N_2267,N_2275);
and U3328 (N_3328,N_1329,N_2521);
nand U3329 (N_3329,In_208,N_2105);
or U3330 (N_3330,N_2064,N_2494);
and U3331 (N_3331,N_2014,N_2608);
nor U3332 (N_3332,N_2367,N_2197);
nand U3333 (N_3333,N_2655,N_2901);
nand U3334 (N_3334,In_2741,In_4572);
nor U3335 (N_3335,N_2518,N_2457);
or U3336 (N_3336,N_2665,N_1526);
or U3337 (N_3337,In_3732,N_1451);
or U3338 (N_3338,In_4251,N_2579);
xnor U3339 (N_3339,N_2557,In_2347);
nor U3340 (N_3340,N_2861,N_1846);
nor U3341 (N_3341,N_2328,N_2233);
xnor U3342 (N_3342,N_2060,N_2672);
nor U3343 (N_3343,N_1120,N_2899);
and U3344 (N_3344,In_394,N_2818);
and U3345 (N_3345,N_2031,N_585);
and U3346 (N_3346,N_2932,In_3202);
xnor U3347 (N_3347,N_2247,N_2524);
nand U3348 (N_3348,In_682,N_1994);
and U3349 (N_3349,N_1866,In_1760);
and U3350 (N_3350,N_2664,In_4548);
and U3351 (N_3351,N_2878,N_2993);
xnor U3352 (N_3352,N_2285,N_2855);
or U3353 (N_3353,N_2732,In_2225);
xnor U3354 (N_3354,N_2054,N_2343);
nor U3355 (N_3355,N_2954,N_2034);
or U3356 (N_3356,N_2163,N_2351);
and U3357 (N_3357,N_2116,N_1601);
and U3358 (N_3358,N_2281,In_57);
nor U3359 (N_3359,N_2471,N_2015);
nand U3360 (N_3360,N_2787,N_2447);
or U3361 (N_3361,N_1156,N_2923);
and U3362 (N_3362,N_1743,N_66);
or U3363 (N_3363,N_2236,In_2526);
xor U3364 (N_3364,N_2436,In_1682);
nor U3365 (N_3365,In_130,In_2061);
or U3366 (N_3366,N_2249,N_2611);
or U3367 (N_3367,N_2622,In_4245);
nor U3368 (N_3368,In_2242,In_1145);
and U3369 (N_3369,N_2633,N_2166);
xnor U3370 (N_3370,N_2586,N_2362);
or U3371 (N_3371,N_2678,N_1679);
and U3372 (N_3372,N_2323,N_2131);
or U3373 (N_3373,In_484,N_661);
or U3374 (N_3374,N_2719,N_2846);
nand U3375 (N_3375,N_2884,N_2480);
nor U3376 (N_3376,N_1364,N_2104);
or U3377 (N_3377,N_2271,N_29);
nand U3378 (N_3378,N_2085,N_1427);
and U3379 (N_3379,In_4109,In_4908);
or U3380 (N_3380,N_2354,N_470);
nand U3381 (N_3381,N_2865,In_4171);
or U3382 (N_3382,N_2290,In_2643);
nor U3383 (N_3383,In_4950,N_657);
xor U3384 (N_3384,N_2571,In_3538);
or U3385 (N_3385,N_1,N_1805);
nand U3386 (N_3386,N_2922,N_2870);
or U3387 (N_3387,In_2709,N_2024);
nor U3388 (N_3388,N_489,In_1709);
or U3389 (N_3389,N_2773,In_634);
xor U3390 (N_3390,N_211,N_605);
nand U3391 (N_3391,In_167,N_1347);
nor U3392 (N_3392,In_678,N_2355);
or U3393 (N_3393,N_2737,In_1130);
nor U3394 (N_3394,N_2767,N_26);
or U3395 (N_3395,In_4361,In_4186);
and U3396 (N_3396,N_2342,N_1588);
or U3397 (N_3397,N_1981,N_2175);
nor U3398 (N_3398,N_2780,N_2968);
and U3399 (N_3399,N_2942,N_2642);
nand U3400 (N_3400,N_2432,N_2217);
nand U3401 (N_3401,In_4340,In_3769);
and U3402 (N_3402,N_2079,N_2605);
xor U3403 (N_3403,N_2926,N_1732);
nor U3404 (N_3404,N_2023,N_2279);
or U3405 (N_3405,N_1477,In_862);
and U3406 (N_3406,N_2562,N_2257);
xor U3407 (N_3407,N_2465,In_2084);
xnor U3408 (N_3408,In_851,In_2124);
and U3409 (N_3409,In_4114,N_888);
nand U3410 (N_3410,N_1159,N_2220);
xnor U3411 (N_3411,N_1954,N_2943);
nand U3412 (N_3412,N_1959,N_314);
or U3413 (N_3413,N_2057,N_2713);
nor U3414 (N_3414,N_2915,N_1445);
and U3415 (N_3415,N_2277,In_4813);
or U3416 (N_3416,In_255,N_2491);
nand U3417 (N_3417,In_1562,N_2151);
and U3418 (N_3418,In_4529,In_4240);
nor U3419 (N_3419,N_2201,In_1101);
nand U3420 (N_3420,N_1183,N_449);
xor U3421 (N_3421,N_2182,N_2046);
nor U3422 (N_3422,N_2748,N_1467);
or U3423 (N_3423,In_3630,N_2671);
nor U3424 (N_3424,N_1573,In_31);
and U3425 (N_3425,N_2729,N_1109);
nor U3426 (N_3426,In_2948,N_477);
xor U3427 (N_3427,N_2859,N_2550);
nand U3428 (N_3428,In_731,N_2033);
or U3429 (N_3429,N_309,N_2331);
nand U3430 (N_3430,In_4759,N_2796);
nor U3431 (N_3431,N_2330,N_2437);
nor U3432 (N_3432,N_2635,N_301);
xor U3433 (N_3433,N_78,N_2987);
xnor U3434 (N_3434,In_3660,In_4564);
nor U3435 (N_3435,N_2793,N_2913);
xnor U3436 (N_3436,In_2533,N_75);
nand U3437 (N_3437,N_2830,In_3943);
xor U3438 (N_3438,N_1697,In_495);
nand U3439 (N_3439,N_2320,In_1120);
nand U3440 (N_3440,N_2028,N_1701);
nand U3441 (N_3441,N_1169,N_1764);
nor U3442 (N_3442,N_1482,N_2545);
nor U3443 (N_3443,N_2100,N_2561);
xnor U3444 (N_3444,N_1724,In_3905);
or U3445 (N_3445,In_4348,N_2694);
and U3446 (N_3446,N_2858,N_2797);
or U3447 (N_3447,N_2684,N_2680);
and U3448 (N_3448,N_2546,N_2195);
xnor U3449 (N_3449,N_2188,In_2789);
or U3450 (N_3450,N_1569,In_3866);
nor U3451 (N_3451,N_2165,N_2848);
nor U3452 (N_3452,N_2774,N_1804);
nand U3453 (N_3453,N_2311,N_1440);
nand U3454 (N_3454,In_962,N_2231);
xor U3455 (N_3455,N_2874,N_1880);
or U3456 (N_3456,In_4549,N_186);
or U3457 (N_3457,N_1551,N_712);
nand U3458 (N_3458,In_2512,In_4270);
nor U3459 (N_3459,N_2800,N_299);
and U3460 (N_3460,N_1841,N_2293);
or U3461 (N_3461,N_2118,N_2749);
nand U3462 (N_3462,N_2629,N_2536);
nand U3463 (N_3463,N_2824,N_2564);
xnor U3464 (N_3464,N_901,N_1332);
and U3465 (N_3465,In_4746,In_2900);
or U3466 (N_3466,N_2080,In_3557);
or U3467 (N_3467,N_2623,In_1370);
nand U3468 (N_3468,N_2881,N_2404);
and U3469 (N_3469,In_4930,N_2075);
or U3470 (N_3470,N_1791,N_2715);
or U3471 (N_3471,N_1167,N_1293);
xnor U3472 (N_3472,N_2726,N_2650);
and U3473 (N_3473,In_4173,N_132);
nor U3474 (N_3474,In_4206,In_3164);
or U3475 (N_3475,N_2724,In_3741);
or U3476 (N_3476,N_2303,N_2027);
nor U3477 (N_3477,N_2582,N_2892);
or U3478 (N_3478,N_1027,N_2946);
nor U3479 (N_3479,N_2463,N_2742);
and U3480 (N_3480,N_2572,In_4579);
nor U3481 (N_3481,N_2088,N_2430);
or U3482 (N_3482,N_2389,N_2513);
or U3483 (N_3483,N_2985,N_2508);
xnor U3484 (N_3484,N_2723,In_1568);
xnor U3485 (N_3485,N_2689,In_4307);
and U3486 (N_3486,In_1413,N_2486);
or U3487 (N_3487,In_4091,In_3792);
xor U3488 (N_3488,In_3311,In_2301);
nor U3489 (N_3489,N_2802,N_2577);
and U3490 (N_3490,N_727,N_2598);
xnor U3491 (N_3491,N_2081,In_3971);
and U3492 (N_3492,N_2875,N_98);
or U3493 (N_3493,N_2107,N_32);
and U3494 (N_3494,N_2384,N_1650);
and U3495 (N_3495,N_2126,N_2539);
nor U3496 (N_3496,N_2720,N_1799);
xor U3497 (N_3497,In_10,In_101);
nor U3498 (N_3498,N_1727,N_1990);
nand U3499 (N_3499,N_2265,N_2072);
and U3500 (N_3500,In_2858,N_2406);
nand U3501 (N_3501,N_133,N_2976);
xor U3502 (N_3502,N_2361,N_1232);
xor U3503 (N_3503,N_2288,N_1756);
nor U3504 (N_3504,In_3743,N_2529);
xor U3505 (N_3505,In_2950,In_4116);
xor U3506 (N_3506,N_2299,N_1424);
nor U3507 (N_3507,N_2504,N_2967);
and U3508 (N_3508,N_2596,N_600);
nor U3509 (N_3509,N_632,N_2599);
or U3510 (N_3510,N_2683,N_2211);
or U3511 (N_3511,N_2940,N_2337);
and U3512 (N_3512,N_381,N_1494);
xnor U3513 (N_3513,N_2103,N_1298);
and U3514 (N_3514,In_4066,N_2804);
nor U3515 (N_3515,N_2807,N_1129);
nor U3516 (N_3516,N_14,N_2189);
nor U3517 (N_3517,N_2474,N_2956);
or U3518 (N_3518,In_1654,N_2717);
or U3519 (N_3519,N_114,N_1499);
or U3520 (N_3520,N_2155,N_2375);
or U3521 (N_3521,N_2540,N_1571);
or U3522 (N_3522,N_1481,In_2210);
nand U3523 (N_3523,N_2317,In_1112);
nor U3524 (N_3524,N_2234,N_52);
nor U3525 (N_3525,In_2275,N_1862);
and U3526 (N_3526,In_2412,In_1931);
or U3527 (N_3527,N_1657,N_342);
nand U3528 (N_3528,N_2668,In_2607);
or U3529 (N_3529,N_1956,N_2566);
nand U3530 (N_3530,N_2451,N_2709);
and U3531 (N_3531,N_2970,N_2483);
nor U3532 (N_3532,N_2378,N_2977);
nand U3533 (N_3533,N_2522,In_87);
or U3534 (N_3534,N_1590,N_1843);
or U3535 (N_3535,N_1714,In_1835);
nand U3536 (N_3536,In_34,In_729);
nor U3537 (N_3537,N_2627,N_1514);
nor U3538 (N_3538,In_2113,N_2974);
or U3539 (N_3539,N_2282,N_2769);
nor U3540 (N_3540,N_1052,N_2573);
or U3541 (N_3541,In_4194,N_2653);
nor U3542 (N_3542,N_2631,In_28);
nor U3543 (N_3543,In_3072,N_2185);
xor U3544 (N_3544,N_2527,In_1467);
nor U3545 (N_3545,N_1363,N_2042);
nor U3546 (N_3546,N_2505,N_1341);
nand U3547 (N_3547,N_1522,N_1622);
and U3548 (N_3548,N_2413,N_1790);
and U3549 (N_3549,N_2666,In_328);
and U3550 (N_3550,N_2746,N_2578);
nor U3551 (N_3551,In_4113,N_656);
or U3552 (N_3552,In_1506,N_2886);
nand U3553 (N_3553,N_2990,In_1617);
nand U3554 (N_3554,N_2435,N_2468);
or U3555 (N_3555,In_3407,N_2125);
xnor U3556 (N_3556,In_4739,In_4583);
or U3557 (N_3557,N_782,N_2333);
nand U3558 (N_3558,N_2475,N_2410);
or U3559 (N_3559,N_2949,N_957);
and U3560 (N_3560,N_1554,N_2656);
nor U3561 (N_3561,N_2392,N_2184);
xnor U3562 (N_3562,N_2708,N_2836);
xor U3563 (N_3563,N_2173,N_2782);
or U3564 (N_3564,N_2997,N_2372);
or U3565 (N_3565,In_1065,N_1447);
nor U3566 (N_3566,In_2149,In_207);
nor U3567 (N_3567,N_2677,N_2711);
nor U3568 (N_3568,N_1927,In_2087);
nand U3569 (N_3569,In_1895,N_2587);
or U3570 (N_3570,N_2338,In_3129);
xnor U3571 (N_3571,N_679,N_2520);
xnor U3572 (N_3572,N_1002,N_2066);
or U3573 (N_3573,N_2464,In_1980);
or U3574 (N_3574,N_2585,N_2146);
nand U3575 (N_3575,N_2798,N_2833);
or U3576 (N_3576,In_2154,N_2995);
xor U3577 (N_3577,N_2485,N_1644);
and U3578 (N_3578,In_1289,N_2191);
nor U3579 (N_3579,N_1399,In_2298);
and U3580 (N_3580,N_2482,N_1692);
or U3581 (N_3581,In_2269,In_63);
and U3582 (N_3582,N_2626,N_2113);
nand U3583 (N_3583,N_2168,N_483);
and U3584 (N_3584,N_2603,N_1153);
and U3585 (N_3585,N_272,N_2601);
or U3586 (N_3586,N_1486,N_1220);
xnor U3587 (N_3587,N_1984,In_48);
or U3588 (N_3588,N_209,N_2619);
nor U3589 (N_3589,In_267,N_2462);
and U3590 (N_3590,N_2722,N_2453);
nor U3591 (N_3591,N_2094,N_1761);
and U3592 (N_3592,N_2135,N_1266);
nand U3593 (N_3593,N_1937,N_1267);
xnor U3594 (N_3594,N_2706,In_1841);
or U3595 (N_3595,N_2506,In_4717);
nor U3596 (N_3596,N_2177,N_2349);
nor U3597 (N_3597,N_2339,In_459);
xnor U3598 (N_3598,In_4934,N_2553);
xor U3599 (N_3599,N_2636,N_2744);
or U3600 (N_3600,In_3965,N_2785);
and U3601 (N_3601,N_2693,N_2484);
xor U3602 (N_3602,N_2755,N_997);
xnor U3603 (N_3603,In_2163,N_2721);
or U3604 (N_3604,N_2883,N_2869);
or U3605 (N_3605,N_440,N_2176);
nor U3606 (N_3606,N_280,N_1429);
nor U3607 (N_3607,In_491,In_4061);
or U3608 (N_3608,N_1993,N_2761);
xor U3609 (N_3609,In_3691,N_2162);
nor U3610 (N_3610,N_2269,In_2468);
nand U3611 (N_3611,In_4942,N_1225);
xnor U3612 (N_3612,N_348,In_917);
nand U3613 (N_3613,N_1796,In_4986);
and U3614 (N_3614,N_349,N_2772);
xnor U3615 (N_3615,N_2036,N_2735);
xnor U3616 (N_3616,In_1135,N_2095);
nor U3617 (N_3617,In_908,N_2609);
nand U3618 (N_3618,In_4650,N_350);
xor U3619 (N_3619,N_2223,In_4945);
or U3620 (N_3620,N_2488,In_1254);
and U3621 (N_3621,In_2663,N_240);
nor U3622 (N_3622,N_15,N_1868);
nand U3623 (N_3623,N_2393,N_2108);
nand U3624 (N_3624,N_1798,N_2929);
nor U3625 (N_3625,N_1852,In_4695);
nand U3626 (N_3626,In_730,In_3482);
or U3627 (N_3627,N_2472,N_1396);
nand U3628 (N_3628,N_2700,In_3136);
nor U3629 (N_3629,N_616,In_2487);
nor U3630 (N_3630,N_1686,N_2876);
nand U3631 (N_3631,N_2356,N_2202);
and U3632 (N_3632,N_2897,In_1808);
or U3633 (N_3633,N_1885,In_2328);
xor U3634 (N_3634,N_2634,N_2759);
and U3635 (N_3635,N_2652,In_1461);
nor U3636 (N_3636,N_2931,N_2921);
nand U3637 (N_3637,N_2431,N_2047);
nand U3638 (N_3638,N_2843,In_1517);
or U3639 (N_3639,N_2810,N_1556);
or U3640 (N_3640,N_237,N_2262);
and U3641 (N_3641,N_2041,N_2181);
or U3642 (N_3642,N_2691,N_2213);
or U3643 (N_3643,N_1106,N_2939);
nand U3644 (N_3644,N_2495,N_2817);
xor U3645 (N_3645,N_2134,N_2408);
nor U3646 (N_3646,In_3591,N_2067);
nand U3647 (N_3647,N_2563,In_3289);
or U3648 (N_3648,N_2212,N_2583);
or U3649 (N_3649,N_1529,N_1552);
or U3650 (N_3650,N_1373,N_2304);
nand U3651 (N_3651,In_2382,N_2885);
and U3652 (N_3652,N_2170,In_3566);
nor U3653 (N_3653,N_2018,In_166);
and U3654 (N_3654,N_2525,N_2139);
and U3655 (N_3655,N_2448,In_1284);
and U3656 (N_3656,In_315,N_2385);
nor U3657 (N_3657,N_2560,In_3402);
nor U3658 (N_3658,N_2391,N_2654);
xnor U3659 (N_3659,N_2199,N_2548);
or U3660 (N_3660,N_2196,In_1947);
xor U3661 (N_3661,N_2192,In_4512);
and U3662 (N_3662,N_2458,N_2444);
nand U3663 (N_3663,N_2740,N_2957);
xnor U3664 (N_3664,In_335,N_1656);
and U3665 (N_3665,N_1243,N_2620);
xnor U3666 (N_3666,N_2306,N_2651);
and U3667 (N_3667,N_691,N_2187);
nor U3668 (N_3668,N_2335,In_1420);
nand U3669 (N_3669,In_3763,In_4780);
or U3670 (N_3670,N_1284,N_2747);
or U3671 (N_3671,N_2240,N_1431);
or U3672 (N_3672,In_4851,N_1092);
nor U3673 (N_3673,In_1198,N_2558);
nor U3674 (N_3674,N_1107,N_2789);
xor U3675 (N_3675,In_4193,N_2316);
nand U3676 (N_3676,N_2862,N_1960);
xnor U3677 (N_3677,N_2050,N_228);
xor U3678 (N_3678,N_952,N_1664);
nor U3679 (N_3679,N_1989,N_2114);
xor U3680 (N_3680,N_1842,In_848);
and U3681 (N_3681,N_2514,N_2888);
nor U3682 (N_3682,N_1126,N_2098);
and U3683 (N_3683,N_1674,N_1033);
nor U3684 (N_3684,N_2924,N_1252);
and U3685 (N_3685,N_2853,In_4532);
nor U3686 (N_3686,In_1894,In_4724);
nor U3687 (N_3687,N_2890,N_833);
nor U3688 (N_3688,N_1785,In_801);
or U3689 (N_3689,N_2919,N_2358);
or U3690 (N_3690,In_4432,N_178);
nand U3691 (N_3691,In_4424,N_2200);
nand U3692 (N_3692,N_473,N_2975);
xor U3693 (N_3693,In_176,N_2365);
nor U3694 (N_3694,N_2037,In_876);
xor U3695 (N_3695,N_1073,N_2637);
nor U3696 (N_3696,N_2783,N_2061);
xor U3697 (N_3697,N_2228,N_2978);
nor U3698 (N_3698,N_206,N_1338);
nor U3699 (N_3699,N_918,N_1130);
nand U3700 (N_3700,N_685,N_2771);
nand U3701 (N_3701,N_2278,N_2149);
nor U3702 (N_3702,N_2371,N_1371);
xnor U3703 (N_3703,N_396,N_2280);
xor U3704 (N_3704,N_1720,N_2106);
or U3705 (N_3705,N_461,N_1894);
nand U3706 (N_3706,N_2756,N_2998);
or U3707 (N_3707,N_2516,In_3860);
nand U3708 (N_3708,N_731,In_1869);
or U3709 (N_3709,N_2989,In_158);
nor U3710 (N_3710,N_1466,In_2719);
xor U3711 (N_3711,N_2592,N_2912);
nand U3712 (N_3712,In_2832,N_1095);
and U3713 (N_3713,N_2914,N_2835);
or U3714 (N_3714,N_2986,N_2594);
or U3715 (N_3715,N_2272,N_2541);
or U3716 (N_3716,In_4744,In_1150);
or U3717 (N_3717,In_2525,N_846);
nand U3718 (N_3718,N_1925,N_1177);
xor U3719 (N_3719,N_2049,N_2423);
nand U3720 (N_3720,In_3644,N_2364);
xnor U3721 (N_3721,N_2243,N_1480);
or U3722 (N_3722,In_4279,In_991);
or U3723 (N_3723,N_2699,N_2503);
or U3724 (N_3724,N_2567,N_2895);
or U3725 (N_3725,N_1618,N_1619);
xor U3726 (N_3726,In_574,N_1405);
nand U3727 (N_3727,N_2441,N_2381);
nor U3728 (N_3728,In_3632,N_2069);
xnor U3729 (N_3729,N_2948,N_2017);
nand U3730 (N_3730,In_2764,N_2930);
nor U3731 (N_3731,N_2658,N_255);
nand U3732 (N_3732,N_1498,N_1034);
nand U3733 (N_3733,N_2763,N_2750);
nor U3734 (N_3734,N_2955,N_2421);
nand U3735 (N_3735,N_2009,In_576);
or U3736 (N_3736,N_275,N_1658);
nor U3737 (N_3737,N_2044,N_1155);
nor U3738 (N_3738,N_2509,N_145);
or U3739 (N_3739,In_4657,N_1976);
and U3740 (N_3740,In_4385,N_1261);
nor U3741 (N_3741,N_2314,N_1233);
nor U3742 (N_3742,N_2641,N_2090);
or U3743 (N_3743,N_2682,N_2120);
nor U3744 (N_3744,N_2048,N_2141);
and U3745 (N_3745,N_2242,N_2092);
and U3746 (N_3746,In_2076,N_2673);
nand U3747 (N_3747,In_1225,N_2097);
nand U3748 (N_3748,In_3754,N_2455);
or U3749 (N_3749,N_2167,N_2803);
nand U3750 (N_3750,N_2676,N_2235);
and U3751 (N_3751,N_760,In_4144);
nand U3752 (N_3752,In_3396,N_1998);
and U3753 (N_3753,In_2315,In_4456);
and U3754 (N_3754,N_2904,N_2645);
xnor U3755 (N_3755,N_2259,N_2022);
or U3756 (N_3756,N_2826,N_2284);
xor U3757 (N_3757,N_650,In_4182);
xor U3758 (N_3758,N_2860,In_2239);
xnor U3759 (N_3759,N_2710,N_2918);
nor U3760 (N_3760,N_1957,N_2347);
xnor U3761 (N_3761,N_2965,N_818);
xnor U3762 (N_3762,N_2123,In_1087);
xnor U3763 (N_3763,N_2531,N_1247);
or U3764 (N_3764,N_2140,N_295);
and U3765 (N_3765,N_2893,In_2217);
nor U3766 (N_3766,In_243,In_2714);
nand U3767 (N_3767,N_2065,N_693);
nand U3768 (N_3768,N_2686,N_688);
xnor U3769 (N_3769,In_366,N_2628);
xnor U3770 (N_3770,N_2035,N_2827);
nor U3771 (N_3771,N_1352,In_2322);
and U3772 (N_3772,N_2227,N_1769);
nand U3773 (N_3773,In_3049,N_2983);
or U3774 (N_3774,N_2346,N_821);
nand U3775 (N_3775,N_707,In_2772);
and U3776 (N_3776,N_1502,N_2315);
xnor U3777 (N_3777,In_4775,N_2245);
and U3778 (N_3778,N_487,N_1382);
xor U3779 (N_3779,N_1883,N_2958);
nor U3780 (N_3780,N_2951,N_2000);
nand U3781 (N_3781,In_3458,N_2237);
and U3782 (N_3782,N_785,N_2937);
or U3783 (N_3783,In_2959,N_2222);
and U3784 (N_3784,N_2297,N_2147);
or U3785 (N_3785,N_2669,In_2539);
xnor U3786 (N_3786,N_795,N_2526);
nor U3787 (N_3787,In_1206,N_215);
nor U3788 (N_3788,In_425,N_2595);
nor U3789 (N_3789,In_2523,N_1510);
nor U3790 (N_3790,N_2178,N_2086);
xnor U3791 (N_3791,N_2174,N_2964);
nor U3792 (N_3792,N_2336,N_2543);
and U3793 (N_3793,N_1624,N_2411);
or U3794 (N_3794,N_2670,In_1124);
nand U3795 (N_3795,N_2002,N_2610);
and U3796 (N_3796,N_2145,In_4437);
xor U3797 (N_3797,N_2440,N_1024);
nand U3798 (N_3798,N_1809,N_2533);
xor U3799 (N_3799,In_3954,In_4687);
xnor U3800 (N_3800,N_2523,N_2604);
nand U3801 (N_3801,N_1964,N_2012);
nand U3802 (N_3802,N_2784,N_2823);
or U3803 (N_3803,N_2405,N_2734);
nor U3804 (N_3804,N_2927,In_782);
or U3805 (N_3805,N_2422,N_2994);
nor U3806 (N_3806,In_531,N_2618);
xor U3807 (N_3807,In_2430,N_1630);
or U3808 (N_3808,N_2055,In_2471);
or U3809 (N_3809,In_4712,In_2004);
or U3810 (N_3810,N_1367,In_4937);
nor U3811 (N_3811,N_1540,In_1352);
or U3812 (N_3812,N_2908,N_2727);
and U3813 (N_3813,N_2920,N_2461);
xnor U3814 (N_3814,N_2690,N_2032);
nor U3815 (N_3815,In_4377,N_2258);
nand U3816 (N_3816,N_2792,N_1108);
and U3817 (N_3817,N_1810,In_965);
and U3818 (N_3818,N_2038,N_2519);
and U3819 (N_3819,In_333,In_1727);
xor U3820 (N_3820,N_2274,In_3693);
and U3821 (N_3821,N_2831,N_1312);
and U3822 (N_3822,N_2446,N_786);
nor U3823 (N_3823,N_2143,N_2214);
or U3824 (N_3824,N_2950,In_2805);
nor U3825 (N_3825,N_510,In_1528);
nand U3826 (N_3826,In_4008,In_1429);
nor U3827 (N_3827,N_2379,N_2832);
xnor U3828 (N_3828,N_2819,In_3903);
nand U3829 (N_3829,In_757,N_2084);
nand U3830 (N_3830,N_2253,N_353);
and U3831 (N_3831,N_2110,N_1056);
and U3832 (N_3832,N_2450,N_2718);
or U3833 (N_3833,In_3584,N_1930);
nor U3834 (N_3834,N_2459,N_2169);
nand U3835 (N_3835,N_392,N_2900);
nor U3836 (N_3836,N_2156,In_4202);
nand U3837 (N_3837,N_2496,N_2894);
nor U3838 (N_3838,N_2369,N_2216);
and U3839 (N_3839,N_2291,In_2856);
xnor U3840 (N_3840,N_2225,N_1058);
nand U3841 (N_3841,N_2544,N_2743);
nor U3842 (N_3842,N_2326,N_2183);
xnor U3843 (N_3843,In_2414,N_2076);
and U3844 (N_3844,N_2403,N_2209);
and U3845 (N_3845,N_1478,In_4985);
or U3846 (N_3846,In_2711,N_2570);
xnor U3847 (N_3847,N_362,N_2753);
xor U3848 (N_3848,N_2040,N_1703);
or U3849 (N_3849,In_4555,N_880);
nor U3850 (N_3850,In_2389,N_1995);
xor U3851 (N_3851,In_1424,N_2062);
nor U3852 (N_3852,N_2241,In_2074);
xor U3853 (N_3853,N_1320,N_2580);
xor U3854 (N_3854,N_2644,N_2758);
or U3855 (N_3855,N_2845,N_1224);
xnor U3856 (N_3856,N_2319,N_1584);
or U3857 (N_3857,In_4322,N_2119);
and U3858 (N_3858,N_112,N_714);
nand U3859 (N_3859,N_1896,N_2996);
nand U3860 (N_3860,N_497,N_2210);
or U3861 (N_3861,N_2093,N_2053);
and U3862 (N_3862,In_4026,N_2395);
nor U3863 (N_3863,N_2538,N_2981);
nor U3864 (N_3864,N_1334,N_609);
xnor U3865 (N_3865,In_2170,N_2171);
or U3866 (N_3866,N_2251,In_541);
xnor U3867 (N_3867,N_2007,N_2971);
nor U3868 (N_3868,N_1840,In_24);
nand U3869 (N_3869,N_2016,N_566);
nand U3870 (N_3870,N_2298,N_1321);
or U3871 (N_3871,N_150,N_1444);
xnor U3872 (N_3872,N_2960,In_1494);
or U3873 (N_3873,N_1891,N_931);
or U3874 (N_3874,In_945,N_1036);
nand U3875 (N_3875,N_624,N_2383);
xor U3876 (N_3876,N_2933,N_729);
xor U3877 (N_3877,N_967,N_2554);
nor U3878 (N_3878,N_2268,N_2714);
nand U3879 (N_3879,N_2266,N_2685);
nand U3880 (N_3880,N_1355,N_500);
nor U3881 (N_3881,N_2776,N_2454);
nand U3882 (N_3882,N_2153,N_1428);
nand U3883 (N_3883,N_2350,N_2547);
nand U3884 (N_3884,N_2051,N_1520);
nand U3885 (N_3885,In_3935,N_2340);
nor U3886 (N_3886,N_2456,N_1684);
xor U3887 (N_3887,N_1941,N_1123);
xor U3888 (N_3888,N_1393,N_2101);
or U3889 (N_3889,N_789,In_3987);
nor U3890 (N_3890,N_1388,N_2679);
nor U3891 (N_3891,In_21,In_3879);
nand U3892 (N_3892,N_2962,N_1700);
nor U3893 (N_3893,N_1749,N_732);
nand U3894 (N_3894,N_1813,N_1179);
or U3895 (N_3895,In_2673,N_717);
and U3896 (N_3896,N_2502,N_1044);
nor U3897 (N_3897,N_2882,N_2697);
nand U3898 (N_3898,N_2795,N_2332);
or U3899 (N_3899,N_2935,In_1406);
nor U3900 (N_3900,N_2089,In_401);
xnor U3901 (N_3901,N_2307,In_2273);
nand U3902 (N_3902,N_2745,N_2296);
xor U3903 (N_3903,N_2334,In_1935);
and U3904 (N_3904,N_2043,In_3345);
nor U3905 (N_3905,N_2158,N_2530);
nor U3906 (N_3906,N_2374,N_1806);
and U3907 (N_3907,N_2469,N_2121);
nand U3908 (N_3908,N_2925,N_2616);
and U3909 (N_3909,In_3451,N_1924);
or U3910 (N_3910,N_1559,In_1385);
or U3911 (N_3911,N_1818,N_2549);
nor U3912 (N_3912,N_2161,N_1807);
and U3913 (N_3913,In_1079,N_2575);
nor U3914 (N_3914,N_2370,N_2808);
nor U3915 (N_3915,In_3024,N_1963);
or U3916 (N_3916,N_1250,N_1921);
nor U3917 (N_3917,N_2109,In_4507);
and U3918 (N_3918,N_2045,N_2988);
or U3919 (N_3919,N_2021,N_1955);
or U3920 (N_3920,N_335,N_2070);
xnor U3921 (N_3921,N_2928,N_855);
nand U3922 (N_3922,N_2896,In_1106);
nand U3923 (N_3923,N_2397,N_2811);
and U3924 (N_3924,In_4887,In_4758);
nor U3925 (N_3925,N_2952,In_3642);
or U3926 (N_3926,N_2728,N_2752);
nand U3927 (N_3927,In_548,N_2232);
or U3928 (N_3928,In_3625,N_2124);
nor U3929 (N_3929,N_2206,N_2492);
nor U3930 (N_3930,N_2373,N_2617);
nand U3931 (N_3931,In_4420,N_2778);
nand U3932 (N_3932,In_4172,N_2467);
nor U3933 (N_3933,N_1135,N_2821);
nand U3934 (N_3934,In_3764,N_2945);
or U3935 (N_3935,N_2799,In_2206);
nor U3936 (N_3936,N_2263,N_2219);
nand U3937 (N_3937,In_1082,N_1333);
or U3938 (N_3938,In_4178,In_3116);
and U3939 (N_3939,In_4856,N_2152);
or U3940 (N_3940,In_3185,N_1198);
or U3941 (N_3941,N_1133,N_2820);
and U3942 (N_3942,N_2591,N_2907);
nand U3943 (N_3943,N_2005,In_4884);
xnor U3944 (N_3944,N_1313,In_2881);
and U3945 (N_3945,N_2058,N_2083);
or U3946 (N_3946,N_356,N_2260);
or U3947 (N_3947,N_1497,In_3675);
nor U3948 (N_3948,In_1059,N_2864);
or U3949 (N_3949,N_1676,N_1914);
xor U3950 (N_3950,N_2305,In_378);
xor U3951 (N_3951,N_2630,N_2345);
xor U3952 (N_3952,In_117,N_2150);
nor U3953 (N_3953,N_2528,N_2218);
nor U3954 (N_3954,N_2493,N_1146);
and U3955 (N_3955,N_2353,N_2226);
nand U3956 (N_3956,N_2341,N_2194);
xnor U3957 (N_3957,N_1929,N_2244);
xor U3958 (N_3958,N_765,In_622);
nor U3959 (N_3959,N_2999,N_2834);
nor U3960 (N_3960,N_1237,N_2292);
nand U3961 (N_3961,In_1165,In_776);
and U3962 (N_3962,In_3391,In_1610);
and U3963 (N_3963,N_1190,N_2229);
or U3964 (N_3964,In_3941,N_2877);
and U3965 (N_3965,N_2606,N_2117);
nand U3966 (N_3966,In_762,N_1009);
xnor U3967 (N_3967,In_544,N_1065);
or U3968 (N_3968,In_4301,N_2532);
nand U3969 (N_3969,N_2438,N_2302);
nand U3970 (N_3970,N_1384,N_2698);
nand U3971 (N_3971,In_4944,N_2781);
xnor U3972 (N_3972,In_2372,N_2944);
nand U3973 (N_3973,N_2115,N_805);
xor U3974 (N_3974,N_590,N_2386);
nor U3975 (N_3975,In_933,N_615);
and U3976 (N_3976,N_1138,N_2415);
and U3977 (N_3977,N_2597,N_368);
nor U3978 (N_3978,N_2324,In_3838);
and U3979 (N_3979,In_692,N_2382);
nor U3980 (N_3980,N_2961,N_2264);
and U3981 (N_3981,N_847,N_2779);
and U3982 (N_3982,N_2867,N_1069);
and U3983 (N_3983,N_2452,N_2813);
nor U3984 (N_3984,N_2638,N_2854);
nor U3985 (N_3985,In_4077,N_1134);
nand U3986 (N_3986,N_1164,N_583);
or U3987 (N_3987,N_587,N_2239);
nor U3988 (N_3988,N_1661,In_1928);
nor U3989 (N_3989,N_2581,In_4204);
and U3990 (N_3990,N_168,N_2099);
or U3991 (N_3991,N_2568,N_2138);
or U3992 (N_3992,In_705,N_2476);
nor U3993 (N_3993,In_3161,N_2313);
nor U3994 (N_3994,N_2639,N_2555);
nor U3995 (N_3995,N_2873,N_2460);
nand U3996 (N_3996,In_3074,N_2248);
nand U3997 (N_3997,N_2512,N_2136);
and U3998 (N_3998,N_2068,In_1414);
or U3999 (N_3999,N_2716,N_1375);
or U4000 (N_4000,N_3144,N_3380);
or U4001 (N_4001,N_3430,N_3586);
nand U4002 (N_4002,N_3957,N_3459);
or U4003 (N_4003,N_3740,N_3089);
or U4004 (N_4004,N_3215,N_3719);
nor U4005 (N_4005,N_3945,N_3280);
and U4006 (N_4006,N_3796,N_3128);
and U4007 (N_4007,N_3631,N_3555);
nor U4008 (N_4008,N_3398,N_3568);
and U4009 (N_4009,N_3046,N_3387);
nor U4010 (N_4010,N_3899,N_3393);
and U4011 (N_4011,N_3080,N_3483);
xor U4012 (N_4012,N_3259,N_3882);
nor U4013 (N_4013,N_3635,N_3379);
nor U4014 (N_4014,N_3561,N_3867);
nor U4015 (N_4015,N_3407,N_3087);
or U4016 (N_4016,N_3200,N_3328);
and U4017 (N_4017,N_3012,N_3578);
xor U4018 (N_4018,N_3662,N_3120);
or U4019 (N_4019,N_3414,N_3893);
or U4020 (N_4020,N_3461,N_3843);
and U4021 (N_4021,N_3311,N_3180);
and U4022 (N_4022,N_3584,N_3032);
and U4023 (N_4023,N_3308,N_3876);
and U4024 (N_4024,N_3305,N_3658);
xnor U4025 (N_4025,N_3829,N_3906);
or U4026 (N_4026,N_3801,N_3902);
xnor U4027 (N_4027,N_3539,N_3491);
and U4028 (N_4028,N_3190,N_3695);
or U4029 (N_4029,N_3663,N_3714);
and U4030 (N_4030,N_3337,N_3637);
and U4031 (N_4031,N_3582,N_3581);
or U4032 (N_4032,N_3777,N_3276);
or U4033 (N_4033,N_3412,N_3840);
or U4034 (N_4034,N_3495,N_3834);
nand U4035 (N_4035,N_3440,N_3039);
nand U4036 (N_4036,N_3696,N_3002);
nand U4037 (N_4037,N_3604,N_3926);
or U4038 (N_4038,N_3060,N_3147);
or U4039 (N_4039,N_3929,N_3329);
xor U4040 (N_4040,N_3874,N_3293);
or U4041 (N_4041,N_3468,N_3507);
or U4042 (N_4042,N_3498,N_3527);
xor U4043 (N_4043,N_3226,N_3941);
or U4044 (N_4044,N_3709,N_3715);
nor U4045 (N_4045,N_3444,N_3804);
or U4046 (N_4046,N_3319,N_3047);
xor U4047 (N_4047,N_3477,N_3918);
xor U4048 (N_4048,N_3419,N_3710);
nor U4049 (N_4049,N_3471,N_3763);
nor U4050 (N_4050,N_3333,N_3399);
or U4051 (N_4051,N_3748,N_3923);
or U4052 (N_4052,N_3066,N_3655);
and U4053 (N_4053,N_3756,N_3921);
xor U4054 (N_4054,N_3282,N_3406);
and U4055 (N_4055,N_3102,N_3776);
nor U4056 (N_4056,N_3091,N_3048);
or U4057 (N_4057,N_3905,N_3737);
and U4058 (N_4058,N_3955,N_3974);
xnor U4059 (N_4059,N_3228,N_3352);
and U4060 (N_4060,N_3513,N_3605);
nor U4061 (N_4061,N_3775,N_3042);
or U4062 (N_4062,N_3236,N_3150);
xnor U4063 (N_4063,N_3057,N_3401);
nor U4064 (N_4064,N_3948,N_3919);
and U4065 (N_4065,N_3678,N_3169);
or U4066 (N_4066,N_3995,N_3699);
and U4067 (N_4067,N_3702,N_3628);
nand U4068 (N_4068,N_3205,N_3001);
and U4069 (N_4069,N_3608,N_3726);
nand U4070 (N_4070,N_3104,N_3881);
xor U4071 (N_4071,N_3667,N_3212);
nand U4072 (N_4072,N_3077,N_3184);
nand U4073 (N_4073,N_3518,N_3421);
xor U4074 (N_4074,N_3272,N_3589);
nor U4075 (N_4075,N_3460,N_3666);
or U4076 (N_4076,N_3478,N_3611);
nand U4077 (N_4077,N_3594,N_3908);
nand U4078 (N_4078,N_3836,N_3376);
xnor U4079 (N_4079,N_3670,N_3009);
nand U4080 (N_4080,N_3659,N_3729);
xor U4081 (N_4081,N_3723,N_3141);
nand U4082 (N_4082,N_3250,N_3958);
and U4083 (N_4083,N_3600,N_3053);
xnor U4084 (N_4084,N_3953,N_3500);
and U4085 (N_4085,N_3525,N_3837);
or U4086 (N_4086,N_3879,N_3064);
and U4087 (N_4087,N_3112,N_3105);
xnor U4088 (N_4088,N_3183,N_3315);
nor U4089 (N_4089,N_3520,N_3253);
xnor U4090 (N_4090,N_3361,N_3956);
nand U4091 (N_4091,N_3467,N_3014);
xor U4092 (N_4092,N_3573,N_3693);
nand U4093 (N_4093,N_3111,N_3725);
and U4094 (N_4094,N_3778,N_3254);
xnor U4095 (N_4095,N_3107,N_3360);
nand U4096 (N_4096,N_3307,N_3920);
and U4097 (N_4097,N_3760,N_3587);
and U4098 (N_4098,N_3552,N_3650);
or U4099 (N_4099,N_3660,N_3409);
nand U4100 (N_4100,N_3121,N_3773);
xnor U4101 (N_4101,N_3024,N_3618);
nand U4102 (N_4102,N_3367,N_3284);
or U4103 (N_4103,N_3869,N_3385);
or U4104 (N_4104,N_3971,N_3353);
or U4105 (N_4105,N_3952,N_3428);
xnor U4106 (N_4106,N_3781,N_3113);
or U4107 (N_4107,N_3934,N_3031);
xor U4108 (N_4108,N_3838,N_3167);
xor U4109 (N_4109,N_3951,N_3641);
nor U4110 (N_4110,N_3320,N_3157);
or U4111 (N_4111,N_3755,N_3232);
xor U4112 (N_4112,N_3441,N_3156);
or U4113 (N_4113,N_3526,N_3109);
nand U4114 (N_4114,N_3872,N_3427);
xor U4115 (N_4115,N_3632,N_3358);
nor U4116 (N_4116,N_3614,N_3241);
and U4117 (N_4117,N_3841,N_3375);
and U4118 (N_4118,N_3548,N_3607);
nand U4119 (N_4119,N_3770,N_3425);
and U4120 (N_4120,N_3197,N_3132);
nor U4121 (N_4121,N_3108,N_3529);
or U4122 (N_4122,N_3571,N_3900);
nand U4123 (N_4123,N_3005,N_3985);
nor U4124 (N_4124,N_3006,N_3751);
nand U4125 (N_4125,N_3317,N_3286);
nand U4126 (N_4126,N_3369,N_3251);
nand U4127 (N_4127,N_3731,N_3451);
xor U4128 (N_4128,N_3949,N_3870);
nor U4129 (N_4129,N_3033,N_3982);
xor U4130 (N_4130,N_3133,N_3558);
and U4131 (N_4131,N_3438,N_3472);
nand U4132 (N_4132,N_3544,N_3545);
nand U4133 (N_4133,N_3887,N_3198);
xor U4134 (N_4134,N_3886,N_3270);
xnor U4135 (N_4135,N_3512,N_3303);
nor U4136 (N_4136,N_3479,N_3283);
or U4137 (N_4137,N_3126,N_3813);
nand U4138 (N_4138,N_3590,N_3221);
or U4139 (N_4139,N_3803,N_3059);
or U4140 (N_4140,N_3866,N_3975);
and U4141 (N_4141,N_3455,N_3986);
and U4142 (N_4142,N_3531,N_3844);
xnor U4143 (N_4143,N_3807,N_3246);
nand U4144 (N_4144,N_3136,N_3967);
and U4145 (N_4145,N_3383,N_3160);
or U4146 (N_4146,N_3713,N_3166);
and U4147 (N_4147,N_3448,N_3368);
nand U4148 (N_4148,N_3370,N_3188);
nand U4149 (N_4149,N_3386,N_3862);
nor U4150 (N_4150,N_3155,N_3217);
nor U4151 (N_4151,N_3853,N_3707);
xor U4152 (N_4152,N_3027,N_3016);
and U4153 (N_4153,N_3187,N_3885);
nand U4154 (N_4154,N_3019,N_3179);
nand U4155 (N_4155,N_3532,N_3417);
or U4156 (N_4156,N_3818,N_3189);
and U4157 (N_4157,N_3884,N_3909);
nor U4158 (N_4158,N_3457,N_3429);
and U4159 (N_4159,N_3208,N_3435);
xnor U4160 (N_4160,N_3446,N_3331);
and U4161 (N_4161,N_3223,N_3359);
or U4162 (N_4162,N_3037,N_3922);
xor U4163 (N_4163,N_3405,N_3738);
or U4164 (N_4164,N_3613,N_3750);
xor U4165 (N_4165,N_3563,N_3903);
xor U4166 (N_4166,N_3959,N_3889);
xnor U4167 (N_4167,N_3809,N_3015);
nor U4168 (N_4168,N_3243,N_3944);
xnor U4169 (N_4169,N_3901,N_3939);
nor U4170 (N_4170,N_3300,N_3694);
nand U4171 (N_4171,N_3576,N_3351);
nand U4172 (N_4172,N_3222,N_3993);
or U4173 (N_4173,N_3690,N_3168);
nor U4174 (N_4174,N_3808,N_3514);
xnor U4175 (N_4175,N_3753,N_3186);
xor U4176 (N_4176,N_3612,N_3134);
or U4177 (N_4177,N_3240,N_3624);
and U4178 (N_4178,N_3022,N_3382);
nand U4179 (N_4179,N_3621,N_3335);
nor U4180 (N_4180,N_3049,N_3404);
xor U4181 (N_4181,N_3814,N_3633);
and U4182 (N_4182,N_3591,N_3860);
nand U4183 (N_4183,N_3038,N_3488);
nand U4184 (N_4184,N_3256,N_3546);
nand U4185 (N_4185,N_3969,N_3864);
and U4186 (N_4186,N_3443,N_3281);
nor U4187 (N_4187,N_3054,N_3026);
xnor U4188 (N_4188,N_3095,N_3799);
xnor U4189 (N_4189,N_3086,N_3090);
nor U4190 (N_4190,N_3721,N_3697);
nand U4191 (N_4191,N_3336,N_3063);
nor U4192 (N_4192,N_3625,N_3123);
and U4193 (N_4193,N_3787,N_3433);
xor U4194 (N_4194,N_3082,N_3069);
nor U4195 (N_4195,N_3285,N_3339);
nor U4196 (N_4196,N_3439,N_3313);
or U4197 (N_4197,N_3868,N_3823);
or U4198 (N_4198,N_3340,N_3671);
nor U4199 (N_4199,N_3540,N_3450);
nor U4200 (N_4200,N_3277,N_3692);
xor U4201 (N_4201,N_3541,N_3292);
xnor U4202 (N_4202,N_3538,N_3850);
nor U4203 (N_4203,N_3848,N_3263);
nand U4204 (N_4204,N_3274,N_3395);
or U4205 (N_4205,N_3269,N_3606);
and U4206 (N_4206,N_3220,N_3258);
xnor U4207 (N_4207,N_3654,N_3774);
nand U4208 (N_4208,N_3065,N_3790);
nor U4209 (N_4209,N_3023,N_3268);
nand U4210 (N_4210,N_3452,N_3865);
or U4211 (N_4211,N_3475,N_3330);
and U4212 (N_4212,N_3999,N_3646);
or U4213 (N_4213,N_3717,N_3354);
or U4214 (N_4214,N_3533,N_3378);
or U4215 (N_4215,N_3691,N_3542);
nand U4216 (N_4216,N_3266,N_3493);
xnor U4217 (N_4217,N_3932,N_3895);
nand U4218 (N_4218,N_3782,N_3580);
nand U4219 (N_4219,N_3296,N_3431);
nor U4220 (N_4220,N_3638,N_3636);
and U4221 (N_4221,N_3494,N_3422);
nor U4222 (N_4222,N_3474,N_3411);
nand U4223 (N_4223,N_3732,N_3977);
and U4224 (N_4224,N_3185,N_3597);
or U4225 (N_4225,N_3391,N_3365);
and U4226 (N_4226,N_3698,N_3152);
nor U4227 (N_4227,N_3505,N_3528);
and U4228 (N_4228,N_3201,N_3904);
nor U4229 (N_4229,N_3516,N_3757);
or U4230 (N_4230,N_3035,N_3878);
nand U4231 (N_4231,N_3793,N_3766);
and U4232 (N_4232,N_3079,N_3987);
nand U4233 (N_4233,N_3350,N_3828);
or U4234 (N_4234,N_3647,N_3000);
and U4235 (N_4235,N_3348,N_3029);
nor U4236 (N_4236,N_3453,N_3332);
xnor U4237 (N_4237,N_3768,N_3092);
and U4238 (N_4238,N_3791,N_3759);
xnor U4239 (N_4239,N_3289,N_3314);
and U4240 (N_4240,N_3554,N_3744);
or U4241 (N_4241,N_3464,N_3983);
or U4242 (N_4242,N_3159,N_3950);
nand U4243 (N_4243,N_3244,N_3075);
nor U4244 (N_4244,N_3989,N_3927);
xor U4245 (N_4245,N_3767,N_3789);
or U4246 (N_4246,N_3511,N_3871);
nor U4247 (N_4247,N_3783,N_3947);
and U4248 (N_4248,N_3960,N_3177);
and U4249 (N_4249,N_3372,N_3124);
xor U4250 (N_4250,N_3004,N_3550);
or U4251 (N_4251,N_3609,N_3273);
and U4252 (N_4252,N_3897,N_3734);
and U4253 (N_4253,N_3231,N_3786);
nand U4254 (N_4254,N_3362,N_3915);
nand U4255 (N_4255,N_3083,N_3835);
nand U4256 (N_4256,N_3465,N_3070);
and U4257 (N_4257,N_3418,N_3149);
xnor U4258 (N_4258,N_3521,N_3275);
nand U4259 (N_4259,N_3098,N_3326);
nor U4260 (N_4260,N_3400,N_3394);
nor U4261 (N_4261,N_3553,N_3668);
or U4262 (N_4262,N_3396,N_3785);
or U4263 (N_4263,N_3410,N_3980);
nor U4264 (N_4264,N_3937,N_3536);
nand U4265 (N_4265,N_3084,N_3374);
xnor U4266 (N_4266,N_3238,N_3517);
and U4267 (N_4267,N_3255,N_3924);
and U4268 (N_4268,N_3852,N_3306);
xnor U4269 (N_4269,N_3230,N_3547);
or U4270 (N_4270,N_3849,N_3278);
nand U4271 (N_4271,N_3562,N_3992);
nand U4272 (N_4272,N_3653,N_3925);
and U4273 (N_4273,N_3680,N_3146);
nand U4274 (N_4274,N_3788,N_3325);
nor U4275 (N_4275,N_3171,N_3316);
or U4276 (N_4276,N_3825,N_3954);
nand U4277 (N_4277,N_3816,N_3229);
nand U4278 (N_4278,N_3572,N_3499);
or U4279 (N_4279,N_3626,N_3469);
and U4280 (N_4280,N_3492,N_3742);
and U4281 (N_4281,N_3309,N_3570);
xnor U4282 (N_4282,N_3569,N_3020);
xnor U4283 (N_4283,N_3706,N_3261);
nor U4284 (N_4284,N_3481,N_3649);
nand U4285 (N_4285,N_3473,N_3762);
xor U4286 (N_4286,N_3323,N_3248);
or U4287 (N_4287,N_3703,N_3346);
nand U4288 (N_4288,N_3916,N_3687);
and U4289 (N_4289,N_3754,N_3008);
nor U4290 (N_4290,N_3935,N_3771);
xor U4291 (N_4291,N_3040,N_3142);
nor U4292 (N_4292,N_3883,N_3577);
nand U4293 (N_4293,N_3252,N_3802);
or U4294 (N_4294,N_3279,N_3482);
nor U4295 (N_4295,N_3007,N_3988);
xnor U4296 (N_4296,N_3454,N_3288);
xnor U4297 (N_4297,N_3898,N_3704);
and U4298 (N_4298,N_3815,N_3122);
nand U4299 (N_4299,N_3199,N_3373);
or U4300 (N_4300,N_3013,N_3010);
nor U4301 (N_4301,N_3392,N_3297);
or U4302 (N_4302,N_3349,N_3964);
xor U4303 (N_4303,N_3153,N_3745);
xor U4304 (N_4304,N_3101,N_3724);
and U4305 (N_4305,N_3312,N_3769);
nor U4306 (N_4306,N_3181,N_3722);
nand U4307 (N_4307,N_3991,N_3610);
nor U4308 (N_4308,N_3437,N_3863);
nand U4309 (N_4309,N_3055,N_3845);
and U4310 (N_4310,N_3746,N_3859);
nor U4311 (N_4311,N_3749,N_3017);
nand U4312 (N_4312,N_3826,N_3143);
xnor U4313 (N_4313,N_3490,N_3661);
nand U4314 (N_4314,N_3239,N_3942);
xor U4315 (N_4315,N_3970,N_3684);
xor U4316 (N_4316,N_3794,N_3242);
xor U4317 (N_4317,N_3968,N_3736);
xor U4318 (N_4318,N_3456,N_3851);
or U4319 (N_4319,N_3648,N_3644);
nand U4320 (N_4320,N_3797,N_3178);
xnor U4321 (N_4321,N_3928,N_3025);
and U4322 (N_4322,N_3096,N_3973);
nor U4323 (N_4323,N_3219,N_3543);
or U4324 (N_4324,N_3304,N_3629);
nand U4325 (N_4325,N_3994,N_3875);
or U4326 (N_4326,N_3366,N_3299);
xor U4327 (N_4327,N_3676,N_3485);
xor U4328 (N_4328,N_3135,N_3170);
and U4329 (N_4329,N_3739,N_3210);
or U4330 (N_4330,N_3415,N_3463);
or U4331 (N_4331,N_3287,N_3044);
xnor U4332 (N_4332,N_3524,N_3110);
nand U4333 (N_4333,N_3139,N_3912);
nor U4334 (N_4334,N_3592,N_3752);
and U4335 (N_4335,N_3896,N_3930);
or U4336 (N_4336,N_3209,N_3127);
and U4337 (N_4337,N_3138,N_3537);
xor U4338 (N_4338,N_3021,N_3462);
nand U4339 (N_4339,N_3164,N_3338);
nor U4340 (N_4340,N_3484,N_3593);
nor U4341 (N_4341,N_3619,N_3028);
and U4342 (N_4342,N_3355,N_3196);
and U4343 (N_4343,N_3798,N_3377);
nand U4344 (N_4344,N_3730,N_3817);
nor U4345 (N_4345,N_3997,N_3894);
or U4346 (N_4346,N_3117,N_3202);
nor U4347 (N_4347,N_3530,N_3195);
and U4348 (N_4348,N_3347,N_3535);
and U4349 (N_4349,N_3071,N_3093);
and U4350 (N_4350,N_3137,N_3129);
nand U4351 (N_4351,N_3257,N_3657);
nand U4352 (N_4352,N_3735,N_3161);
and U4353 (N_4353,N_3551,N_3779);
nand U4354 (N_4354,N_3733,N_3566);
and U4355 (N_4355,N_3203,N_3356);
and U4356 (N_4356,N_3996,N_3764);
nand U4357 (N_4357,N_3206,N_3842);
xor U4358 (N_4358,N_3642,N_3247);
or U4359 (N_4359,N_3810,N_3343);
nand U4360 (N_4360,N_3436,N_3389);
nand U4361 (N_4361,N_3615,N_3595);
and U4362 (N_4362,N_3708,N_3295);
nand U4363 (N_4363,N_3913,N_3442);
nor U4364 (N_4364,N_3131,N_3984);
nand U4365 (N_4365,N_3390,N_3681);
or U4366 (N_4366,N_3218,N_3043);
nand U4367 (N_4367,N_3602,N_3264);
nand U4368 (N_4368,N_3172,N_3408);
nand U4369 (N_4369,N_3596,N_3074);
nand U4370 (N_4370,N_3669,N_3832);
and U4371 (N_4371,N_3003,N_3728);
xor U4372 (N_4372,N_3034,N_3857);
or U4373 (N_4373,N_3085,N_3076);
or U4374 (N_4374,N_3966,N_3588);
or U4375 (N_4375,N_3599,N_3397);
nand U4376 (N_4376,N_3216,N_3716);
or U4377 (N_4377,N_3700,N_3858);
nor U4378 (N_4378,N_3780,N_3603);
nor U4379 (N_4379,N_3384,N_3194);
nor U4380 (N_4380,N_3234,N_3931);
or U4381 (N_4381,N_3727,N_3585);
nand U4382 (N_4382,N_3165,N_3846);
nor U4383 (N_4383,N_3891,N_3712);
xor U4384 (N_4384,N_3235,N_3861);
xnor U4385 (N_4385,N_3449,N_3933);
and U4386 (N_4386,N_3214,N_3741);
nand U4387 (N_4387,N_3173,N_3761);
or U4388 (N_4388,N_3298,N_3743);
nor U4389 (N_4389,N_3806,N_3998);
or U4390 (N_4390,N_3267,N_3036);
or U4391 (N_4391,N_3665,N_3503);
or U4392 (N_4392,N_3892,N_3420);
or U4393 (N_4393,N_3504,N_3097);
nand U4394 (N_4394,N_3342,N_3940);
or U4395 (N_4395,N_3174,N_3847);
xnor U4396 (N_4396,N_3322,N_3711);
nand U4397 (N_4397,N_3480,N_3962);
or U4398 (N_4398,N_3630,N_3683);
xor U4399 (N_4399,N_3062,N_3045);
nand U4400 (N_4400,N_3424,N_3664);
or U4401 (N_4401,N_3508,N_3327);
nor U4402 (N_4402,N_3510,N_3094);
and U4403 (N_4403,N_3880,N_3990);
xor U4404 (N_4404,N_3301,N_3938);
nor U4405 (N_4405,N_3118,N_3559);
xor U4406 (N_4406,N_3812,N_3402);
or U4407 (N_4407,N_3413,N_3622);
nand U4408 (N_4408,N_3403,N_3486);
nor U4409 (N_4409,N_3772,N_3119);
nand U4410 (N_4410,N_3620,N_3640);
nand U4411 (N_4411,N_3645,N_3078);
nand U4412 (N_4412,N_3100,N_3073);
and U4413 (N_4413,N_3682,N_3565);
and U4414 (N_4414,N_3050,N_3705);
and U4415 (N_4415,N_3639,N_3318);
nor U4416 (N_4416,N_3784,N_3081);
and U4417 (N_4417,N_3765,N_3673);
and U4418 (N_4418,N_3917,N_3911);
xnor U4419 (N_4419,N_3914,N_3509);
nor U4420 (N_4420,N_3225,N_3388);
and U4421 (N_4421,N_3502,N_3163);
nand U4422 (N_4422,N_3487,N_3344);
and U4423 (N_4423,N_3575,N_3564);
and U4424 (N_4424,N_3445,N_3341);
or U4425 (N_4425,N_3634,N_3758);
xor U4426 (N_4426,N_3627,N_3447);
xnor U4427 (N_4427,N_3067,N_3496);
or U4428 (N_4428,N_3207,N_3224);
and U4429 (N_4429,N_3371,N_3689);
nor U4430 (N_4430,N_3821,N_3811);
xor U4431 (N_4431,N_3291,N_3191);
nor U4432 (N_4432,N_3616,N_3675);
and U4433 (N_4433,N_3747,N_3961);
and U4434 (N_4434,N_3556,N_3416);
nand U4435 (N_4435,N_3839,N_3262);
or U4436 (N_4436,N_3116,N_3701);
and U4437 (N_4437,N_3458,N_3824);
xor U4438 (N_4438,N_3334,N_3260);
nand U4439 (N_4439,N_3497,N_3321);
or U4440 (N_4440,N_3506,N_3193);
nor U4441 (N_4441,N_3718,N_3833);
or U4442 (N_4442,N_3557,N_3058);
nor U4443 (N_4443,N_3534,N_3910);
xnor U4444 (N_4444,N_3489,N_3233);
nor U4445 (N_4445,N_3567,N_3115);
or U4446 (N_4446,N_3154,N_3158);
or U4447 (N_4447,N_3981,N_3476);
xnor U4448 (N_4448,N_3855,N_3583);
or U4449 (N_4449,N_3099,N_3979);
nor U4450 (N_4450,N_3432,N_3672);
or U4451 (N_4451,N_3651,N_3830);
and U4452 (N_4452,N_3265,N_3831);
or U4453 (N_4453,N_3051,N_3579);
xnor U4454 (N_4454,N_3720,N_3381);
or U4455 (N_4455,N_3972,N_3685);
nor U4456 (N_4456,N_3656,N_3245);
nand U4457 (N_4457,N_3800,N_3574);
xnor U4458 (N_4458,N_3677,N_3792);
and U4459 (N_4459,N_3237,N_3151);
nor U4460 (N_4460,N_3426,N_3854);
xor U4461 (N_4461,N_3674,N_3125);
xnor U4462 (N_4462,N_3175,N_3030);
nor U4463 (N_4463,N_3466,N_3145);
nor U4464 (N_4464,N_3088,N_3271);
nor U4465 (N_4465,N_3965,N_3114);
or U4466 (N_4466,N_3617,N_3827);
xor U4467 (N_4467,N_3522,N_3470);
nand U4468 (N_4468,N_3890,N_3148);
and U4469 (N_4469,N_3182,N_3888);
and U4470 (N_4470,N_3357,N_3061);
nand U4471 (N_4471,N_3907,N_3211);
nand U4472 (N_4472,N_3943,N_3805);
nor U4473 (N_4473,N_3213,N_3364);
nor U4474 (N_4474,N_3068,N_3363);
or U4475 (N_4475,N_3877,N_3601);
or U4476 (N_4476,N_3820,N_3688);
or U4477 (N_4477,N_3106,N_3936);
or U4478 (N_4478,N_3598,N_3822);
or U4479 (N_4479,N_3130,N_3249);
nor U4480 (N_4480,N_3623,N_3423);
nor U4481 (N_4481,N_3873,N_3192);
or U4482 (N_4482,N_3103,N_3549);
xor U4483 (N_4483,N_3345,N_3290);
nor U4484 (N_4484,N_3056,N_3679);
and U4485 (N_4485,N_3652,N_3162);
or U4486 (N_4486,N_3501,N_3523);
or U4487 (N_4487,N_3976,N_3294);
nand U4488 (N_4488,N_3515,N_3302);
nor U4489 (N_4489,N_3018,N_3978);
and U4490 (N_4490,N_3324,N_3052);
nand U4491 (N_4491,N_3856,N_3227);
and U4492 (N_4492,N_3140,N_3560);
xnor U4493 (N_4493,N_3643,N_3819);
xnor U4494 (N_4494,N_3176,N_3946);
xnor U4495 (N_4495,N_3204,N_3072);
and U4496 (N_4496,N_3310,N_3011);
or U4497 (N_4497,N_3686,N_3519);
or U4498 (N_4498,N_3434,N_3041);
nor U4499 (N_4499,N_3963,N_3795);
and U4500 (N_4500,N_3147,N_3870);
or U4501 (N_4501,N_3979,N_3577);
or U4502 (N_4502,N_3680,N_3559);
and U4503 (N_4503,N_3634,N_3276);
nor U4504 (N_4504,N_3672,N_3732);
and U4505 (N_4505,N_3694,N_3368);
or U4506 (N_4506,N_3360,N_3614);
and U4507 (N_4507,N_3126,N_3095);
or U4508 (N_4508,N_3420,N_3446);
or U4509 (N_4509,N_3422,N_3787);
nor U4510 (N_4510,N_3983,N_3232);
xnor U4511 (N_4511,N_3720,N_3484);
nor U4512 (N_4512,N_3292,N_3202);
and U4513 (N_4513,N_3401,N_3030);
and U4514 (N_4514,N_3761,N_3062);
nor U4515 (N_4515,N_3383,N_3047);
and U4516 (N_4516,N_3218,N_3037);
nand U4517 (N_4517,N_3276,N_3665);
or U4518 (N_4518,N_3357,N_3278);
xor U4519 (N_4519,N_3869,N_3800);
nor U4520 (N_4520,N_3610,N_3461);
nor U4521 (N_4521,N_3205,N_3384);
xor U4522 (N_4522,N_3203,N_3486);
nand U4523 (N_4523,N_3122,N_3036);
nand U4524 (N_4524,N_3016,N_3551);
xor U4525 (N_4525,N_3856,N_3447);
nand U4526 (N_4526,N_3519,N_3275);
and U4527 (N_4527,N_3666,N_3888);
nor U4528 (N_4528,N_3230,N_3502);
and U4529 (N_4529,N_3428,N_3804);
xnor U4530 (N_4530,N_3611,N_3470);
or U4531 (N_4531,N_3751,N_3361);
nor U4532 (N_4532,N_3774,N_3985);
nand U4533 (N_4533,N_3416,N_3320);
xor U4534 (N_4534,N_3232,N_3324);
nor U4535 (N_4535,N_3914,N_3165);
and U4536 (N_4536,N_3071,N_3464);
xnor U4537 (N_4537,N_3563,N_3042);
xnor U4538 (N_4538,N_3849,N_3436);
or U4539 (N_4539,N_3029,N_3556);
nand U4540 (N_4540,N_3829,N_3498);
xor U4541 (N_4541,N_3419,N_3628);
or U4542 (N_4542,N_3929,N_3257);
or U4543 (N_4543,N_3624,N_3730);
and U4544 (N_4544,N_3934,N_3508);
nand U4545 (N_4545,N_3046,N_3532);
xor U4546 (N_4546,N_3866,N_3701);
nor U4547 (N_4547,N_3054,N_3485);
nor U4548 (N_4548,N_3585,N_3805);
nand U4549 (N_4549,N_3919,N_3538);
and U4550 (N_4550,N_3895,N_3909);
xnor U4551 (N_4551,N_3836,N_3128);
xor U4552 (N_4552,N_3786,N_3217);
or U4553 (N_4553,N_3372,N_3325);
or U4554 (N_4554,N_3961,N_3824);
nand U4555 (N_4555,N_3101,N_3842);
nor U4556 (N_4556,N_3602,N_3708);
xnor U4557 (N_4557,N_3194,N_3728);
or U4558 (N_4558,N_3617,N_3781);
nor U4559 (N_4559,N_3744,N_3377);
nand U4560 (N_4560,N_3195,N_3341);
nand U4561 (N_4561,N_3023,N_3965);
xnor U4562 (N_4562,N_3368,N_3703);
and U4563 (N_4563,N_3089,N_3977);
xor U4564 (N_4564,N_3455,N_3348);
xnor U4565 (N_4565,N_3201,N_3411);
xnor U4566 (N_4566,N_3223,N_3624);
or U4567 (N_4567,N_3838,N_3783);
nor U4568 (N_4568,N_3077,N_3907);
and U4569 (N_4569,N_3129,N_3095);
or U4570 (N_4570,N_3126,N_3756);
nor U4571 (N_4571,N_3510,N_3934);
nand U4572 (N_4572,N_3306,N_3512);
nor U4573 (N_4573,N_3199,N_3522);
xor U4574 (N_4574,N_3217,N_3257);
nor U4575 (N_4575,N_3089,N_3909);
or U4576 (N_4576,N_3662,N_3815);
xor U4577 (N_4577,N_3429,N_3416);
nor U4578 (N_4578,N_3322,N_3791);
and U4579 (N_4579,N_3285,N_3749);
and U4580 (N_4580,N_3928,N_3075);
nor U4581 (N_4581,N_3657,N_3206);
or U4582 (N_4582,N_3676,N_3897);
nand U4583 (N_4583,N_3755,N_3639);
or U4584 (N_4584,N_3931,N_3841);
or U4585 (N_4585,N_3198,N_3967);
nand U4586 (N_4586,N_3580,N_3564);
nand U4587 (N_4587,N_3011,N_3263);
and U4588 (N_4588,N_3152,N_3875);
xnor U4589 (N_4589,N_3571,N_3234);
nor U4590 (N_4590,N_3462,N_3438);
nor U4591 (N_4591,N_3491,N_3337);
or U4592 (N_4592,N_3621,N_3566);
xor U4593 (N_4593,N_3482,N_3104);
nor U4594 (N_4594,N_3632,N_3926);
or U4595 (N_4595,N_3932,N_3400);
nor U4596 (N_4596,N_3595,N_3082);
or U4597 (N_4597,N_3861,N_3971);
or U4598 (N_4598,N_3274,N_3661);
and U4599 (N_4599,N_3855,N_3946);
or U4600 (N_4600,N_3925,N_3937);
or U4601 (N_4601,N_3908,N_3132);
nand U4602 (N_4602,N_3428,N_3557);
and U4603 (N_4603,N_3002,N_3856);
or U4604 (N_4604,N_3667,N_3792);
or U4605 (N_4605,N_3855,N_3313);
xnor U4606 (N_4606,N_3405,N_3562);
xor U4607 (N_4607,N_3270,N_3798);
nand U4608 (N_4608,N_3831,N_3171);
nor U4609 (N_4609,N_3525,N_3613);
nand U4610 (N_4610,N_3609,N_3525);
xor U4611 (N_4611,N_3896,N_3544);
xor U4612 (N_4612,N_3301,N_3809);
xnor U4613 (N_4613,N_3379,N_3930);
and U4614 (N_4614,N_3000,N_3230);
xor U4615 (N_4615,N_3643,N_3891);
and U4616 (N_4616,N_3033,N_3733);
xor U4617 (N_4617,N_3748,N_3459);
xnor U4618 (N_4618,N_3208,N_3008);
and U4619 (N_4619,N_3919,N_3916);
and U4620 (N_4620,N_3529,N_3147);
and U4621 (N_4621,N_3851,N_3735);
xor U4622 (N_4622,N_3296,N_3943);
xnor U4623 (N_4623,N_3910,N_3054);
nand U4624 (N_4624,N_3195,N_3722);
and U4625 (N_4625,N_3074,N_3020);
nand U4626 (N_4626,N_3129,N_3481);
or U4627 (N_4627,N_3325,N_3495);
xnor U4628 (N_4628,N_3738,N_3402);
nor U4629 (N_4629,N_3363,N_3076);
or U4630 (N_4630,N_3660,N_3195);
xnor U4631 (N_4631,N_3847,N_3250);
and U4632 (N_4632,N_3285,N_3669);
or U4633 (N_4633,N_3036,N_3178);
or U4634 (N_4634,N_3944,N_3155);
or U4635 (N_4635,N_3201,N_3175);
or U4636 (N_4636,N_3969,N_3991);
and U4637 (N_4637,N_3541,N_3016);
nor U4638 (N_4638,N_3963,N_3662);
or U4639 (N_4639,N_3098,N_3768);
nand U4640 (N_4640,N_3612,N_3007);
or U4641 (N_4641,N_3468,N_3605);
xnor U4642 (N_4642,N_3447,N_3395);
nand U4643 (N_4643,N_3950,N_3074);
nand U4644 (N_4644,N_3954,N_3284);
and U4645 (N_4645,N_3578,N_3475);
or U4646 (N_4646,N_3954,N_3629);
nor U4647 (N_4647,N_3580,N_3033);
or U4648 (N_4648,N_3416,N_3860);
or U4649 (N_4649,N_3278,N_3836);
or U4650 (N_4650,N_3217,N_3873);
and U4651 (N_4651,N_3683,N_3900);
xor U4652 (N_4652,N_3771,N_3781);
or U4653 (N_4653,N_3790,N_3326);
xnor U4654 (N_4654,N_3867,N_3193);
nor U4655 (N_4655,N_3675,N_3299);
nor U4656 (N_4656,N_3353,N_3806);
or U4657 (N_4657,N_3034,N_3258);
nor U4658 (N_4658,N_3238,N_3435);
xnor U4659 (N_4659,N_3594,N_3370);
or U4660 (N_4660,N_3135,N_3215);
or U4661 (N_4661,N_3578,N_3949);
and U4662 (N_4662,N_3131,N_3077);
nand U4663 (N_4663,N_3323,N_3132);
nand U4664 (N_4664,N_3089,N_3742);
xor U4665 (N_4665,N_3711,N_3292);
nor U4666 (N_4666,N_3849,N_3573);
nor U4667 (N_4667,N_3905,N_3481);
nor U4668 (N_4668,N_3766,N_3670);
xor U4669 (N_4669,N_3575,N_3338);
xor U4670 (N_4670,N_3914,N_3375);
nand U4671 (N_4671,N_3037,N_3480);
and U4672 (N_4672,N_3394,N_3087);
and U4673 (N_4673,N_3335,N_3472);
xnor U4674 (N_4674,N_3946,N_3288);
nor U4675 (N_4675,N_3468,N_3737);
nand U4676 (N_4676,N_3335,N_3365);
and U4677 (N_4677,N_3579,N_3820);
and U4678 (N_4678,N_3677,N_3784);
nand U4679 (N_4679,N_3883,N_3026);
or U4680 (N_4680,N_3310,N_3742);
and U4681 (N_4681,N_3038,N_3216);
nand U4682 (N_4682,N_3762,N_3787);
nor U4683 (N_4683,N_3517,N_3537);
nor U4684 (N_4684,N_3865,N_3567);
nor U4685 (N_4685,N_3676,N_3013);
xor U4686 (N_4686,N_3635,N_3644);
and U4687 (N_4687,N_3129,N_3475);
or U4688 (N_4688,N_3438,N_3269);
and U4689 (N_4689,N_3701,N_3427);
and U4690 (N_4690,N_3348,N_3779);
nor U4691 (N_4691,N_3830,N_3146);
nor U4692 (N_4692,N_3879,N_3055);
xnor U4693 (N_4693,N_3630,N_3949);
nand U4694 (N_4694,N_3688,N_3910);
xnor U4695 (N_4695,N_3422,N_3440);
and U4696 (N_4696,N_3610,N_3761);
xor U4697 (N_4697,N_3919,N_3021);
and U4698 (N_4698,N_3874,N_3182);
xnor U4699 (N_4699,N_3235,N_3754);
and U4700 (N_4700,N_3755,N_3990);
nor U4701 (N_4701,N_3239,N_3221);
nand U4702 (N_4702,N_3203,N_3194);
nand U4703 (N_4703,N_3921,N_3099);
nand U4704 (N_4704,N_3589,N_3477);
nor U4705 (N_4705,N_3917,N_3073);
or U4706 (N_4706,N_3480,N_3932);
xor U4707 (N_4707,N_3421,N_3753);
xor U4708 (N_4708,N_3615,N_3432);
nor U4709 (N_4709,N_3467,N_3369);
xnor U4710 (N_4710,N_3995,N_3402);
nand U4711 (N_4711,N_3852,N_3929);
or U4712 (N_4712,N_3810,N_3210);
xnor U4713 (N_4713,N_3555,N_3442);
or U4714 (N_4714,N_3974,N_3531);
nor U4715 (N_4715,N_3401,N_3156);
or U4716 (N_4716,N_3682,N_3891);
and U4717 (N_4717,N_3133,N_3860);
nand U4718 (N_4718,N_3548,N_3070);
nand U4719 (N_4719,N_3090,N_3142);
or U4720 (N_4720,N_3903,N_3304);
or U4721 (N_4721,N_3700,N_3043);
or U4722 (N_4722,N_3652,N_3842);
nand U4723 (N_4723,N_3006,N_3238);
xor U4724 (N_4724,N_3608,N_3214);
and U4725 (N_4725,N_3227,N_3332);
nand U4726 (N_4726,N_3694,N_3489);
and U4727 (N_4727,N_3883,N_3760);
nor U4728 (N_4728,N_3415,N_3071);
nand U4729 (N_4729,N_3931,N_3637);
and U4730 (N_4730,N_3009,N_3812);
and U4731 (N_4731,N_3299,N_3753);
or U4732 (N_4732,N_3939,N_3906);
nand U4733 (N_4733,N_3179,N_3273);
xor U4734 (N_4734,N_3116,N_3787);
xnor U4735 (N_4735,N_3591,N_3960);
and U4736 (N_4736,N_3836,N_3143);
or U4737 (N_4737,N_3635,N_3033);
and U4738 (N_4738,N_3360,N_3648);
or U4739 (N_4739,N_3464,N_3060);
nand U4740 (N_4740,N_3836,N_3749);
and U4741 (N_4741,N_3347,N_3575);
and U4742 (N_4742,N_3149,N_3415);
nand U4743 (N_4743,N_3106,N_3291);
nand U4744 (N_4744,N_3688,N_3126);
xor U4745 (N_4745,N_3913,N_3929);
nor U4746 (N_4746,N_3706,N_3649);
or U4747 (N_4747,N_3401,N_3523);
nand U4748 (N_4748,N_3383,N_3236);
xor U4749 (N_4749,N_3772,N_3579);
and U4750 (N_4750,N_3654,N_3960);
nand U4751 (N_4751,N_3445,N_3308);
or U4752 (N_4752,N_3924,N_3497);
nor U4753 (N_4753,N_3832,N_3193);
nand U4754 (N_4754,N_3908,N_3952);
nand U4755 (N_4755,N_3799,N_3299);
nor U4756 (N_4756,N_3991,N_3422);
nand U4757 (N_4757,N_3437,N_3812);
nand U4758 (N_4758,N_3091,N_3445);
nor U4759 (N_4759,N_3683,N_3160);
nor U4760 (N_4760,N_3935,N_3405);
nand U4761 (N_4761,N_3949,N_3575);
nor U4762 (N_4762,N_3654,N_3844);
and U4763 (N_4763,N_3578,N_3254);
or U4764 (N_4764,N_3513,N_3325);
nand U4765 (N_4765,N_3436,N_3161);
and U4766 (N_4766,N_3836,N_3085);
and U4767 (N_4767,N_3744,N_3555);
xor U4768 (N_4768,N_3083,N_3891);
or U4769 (N_4769,N_3378,N_3456);
nand U4770 (N_4770,N_3925,N_3493);
nand U4771 (N_4771,N_3118,N_3197);
nand U4772 (N_4772,N_3753,N_3121);
xor U4773 (N_4773,N_3598,N_3801);
nand U4774 (N_4774,N_3773,N_3223);
nor U4775 (N_4775,N_3732,N_3608);
or U4776 (N_4776,N_3558,N_3266);
or U4777 (N_4777,N_3853,N_3305);
or U4778 (N_4778,N_3044,N_3233);
and U4779 (N_4779,N_3347,N_3400);
and U4780 (N_4780,N_3746,N_3459);
or U4781 (N_4781,N_3301,N_3376);
and U4782 (N_4782,N_3827,N_3861);
nor U4783 (N_4783,N_3128,N_3333);
and U4784 (N_4784,N_3227,N_3277);
nor U4785 (N_4785,N_3172,N_3766);
or U4786 (N_4786,N_3101,N_3409);
or U4787 (N_4787,N_3488,N_3845);
xnor U4788 (N_4788,N_3543,N_3865);
and U4789 (N_4789,N_3319,N_3662);
nand U4790 (N_4790,N_3558,N_3283);
xor U4791 (N_4791,N_3189,N_3551);
nand U4792 (N_4792,N_3269,N_3248);
nor U4793 (N_4793,N_3534,N_3933);
or U4794 (N_4794,N_3942,N_3069);
nand U4795 (N_4795,N_3071,N_3916);
and U4796 (N_4796,N_3367,N_3214);
nor U4797 (N_4797,N_3496,N_3517);
xnor U4798 (N_4798,N_3396,N_3909);
and U4799 (N_4799,N_3711,N_3638);
nand U4800 (N_4800,N_3103,N_3744);
nor U4801 (N_4801,N_3719,N_3026);
nand U4802 (N_4802,N_3920,N_3451);
and U4803 (N_4803,N_3928,N_3040);
nand U4804 (N_4804,N_3440,N_3595);
or U4805 (N_4805,N_3964,N_3425);
xnor U4806 (N_4806,N_3988,N_3211);
xor U4807 (N_4807,N_3558,N_3980);
or U4808 (N_4808,N_3945,N_3145);
and U4809 (N_4809,N_3001,N_3600);
xor U4810 (N_4810,N_3652,N_3034);
or U4811 (N_4811,N_3665,N_3097);
or U4812 (N_4812,N_3675,N_3167);
xor U4813 (N_4813,N_3299,N_3877);
and U4814 (N_4814,N_3912,N_3512);
xnor U4815 (N_4815,N_3346,N_3685);
and U4816 (N_4816,N_3389,N_3491);
xor U4817 (N_4817,N_3838,N_3554);
or U4818 (N_4818,N_3858,N_3212);
nor U4819 (N_4819,N_3588,N_3753);
and U4820 (N_4820,N_3325,N_3059);
nor U4821 (N_4821,N_3552,N_3182);
nor U4822 (N_4822,N_3605,N_3232);
and U4823 (N_4823,N_3045,N_3184);
xor U4824 (N_4824,N_3181,N_3942);
nor U4825 (N_4825,N_3472,N_3586);
or U4826 (N_4826,N_3360,N_3044);
or U4827 (N_4827,N_3078,N_3238);
or U4828 (N_4828,N_3129,N_3176);
xnor U4829 (N_4829,N_3468,N_3104);
and U4830 (N_4830,N_3598,N_3896);
or U4831 (N_4831,N_3427,N_3466);
and U4832 (N_4832,N_3535,N_3276);
nor U4833 (N_4833,N_3895,N_3342);
xor U4834 (N_4834,N_3541,N_3916);
or U4835 (N_4835,N_3005,N_3848);
nor U4836 (N_4836,N_3832,N_3086);
and U4837 (N_4837,N_3749,N_3163);
xor U4838 (N_4838,N_3922,N_3801);
nor U4839 (N_4839,N_3021,N_3296);
and U4840 (N_4840,N_3566,N_3272);
xnor U4841 (N_4841,N_3158,N_3749);
xnor U4842 (N_4842,N_3327,N_3518);
or U4843 (N_4843,N_3443,N_3799);
and U4844 (N_4844,N_3211,N_3741);
or U4845 (N_4845,N_3856,N_3243);
and U4846 (N_4846,N_3007,N_3045);
nor U4847 (N_4847,N_3256,N_3807);
and U4848 (N_4848,N_3676,N_3575);
nor U4849 (N_4849,N_3169,N_3732);
xnor U4850 (N_4850,N_3159,N_3433);
or U4851 (N_4851,N_3952,N_3482);
and U4852 (N_4852,N_3407,N_3651);
or U4853 (N_4853,N_3529,N_3949);
xor U4854 (N_4854,N_3123,N_3619);
xor U4855 (N_4855,N_3037,N_3700);
xnor U4856 (N_4856,N_3647,N_3238);
nor U4857 (N_4857,N_3266,N_3708);
nand U4858 (N_4858,N_3998,N_3941);
nor U4859 (N_4859,N_3425,N_3643);
or U4860 (N_4860,N_3753,N_3201);
or U4861 (N_4861,N_3396,N_3452);
and U4862 (N_4862,N_3573,N_3349);
and U4863 (N_4863,N_3792,N_3832);
nor U4864 (N_4864,N_3804,N_3133);
or U4865 (N_4865,N_3112,N_3953);
xor U4866 (N_4866,N_3150,N_3771);
and U4867 (N_4867,N_3731,N_3815);
and U4868 (N_4868,N_3911,N_3036);
xor U4869 (N_4869,N_3357,N_3654);
nor U4870 (N_4870,N_3884,N_3808);
nor U4871 (N_4871,N_3124,N_3026);
or U4872 (N_4872,N_3246,N_3027);
nor U4873 (N_4873,N_3774,N_3243);
or U4874 (N_4874,N_3817,N_3166);
nand U4875 (N_4875,N_3180,N_3445);
and U4876 (N_4876,N_3963,N_3461);
nor U4877 (N_4877,N_3641,N_3739);
and U4878 (N_4878,N_3568,N_3145);
or U4879 (N_4879,N_3573,N_3815);
nor U4880 (N_4880,N_3401,N_3881);
nand U4881 (N_4881,N_3661,N_3959);
and U4882 (N_4882,N_3448,N_3171);
and U4883 (N_4883,N_3839,N_3498);
xor U4884 (N_4884,N_3787,N_3844);
or U4885 (N_4885,N_3342,N_3387);
and U4886 (N_4886,N_3501,N_3444);
nand U4887 (N_4887,N_3532,N_3535);
nor U4888 (N_4888,N_3242,N_3368);
nand U4889 (N_4889,N_3939,N_3367);
nand U4890 (N_4890,N_3965,N_3929);
or U4891 (N_4891,N_3948,N_3709);
nor U4892 (N_4892,N_3770,N_3564);
or U4893 (N_4893,N_3315,N_3732);
or U4894 (N_4894,N_3290,N_3976);
nand U4895 (N_4895,N_3062,N_3345);
and U4896 (N_4896,N_3783,N_3475);
xor U4897 (N_4897,N_3499,N_3590);
or U4898 (N_4898,N_3284,N_3040);
and U4899 (N_4899,N_3401,N_3754);
nand U4900 (N_4900,N_3734,N_3801);
or U4901 (N_4901,N_3247,N_3418);
nor U4902 (N_4902,N_3940,N_3629);
and U4903 (N_4903,N_3733,N_3542);
and U4904 (N_4904,N_3820,N_3517);
xnor U4905 (N_4905,N_3411,N_3328);
nor U4906 (N_4906,N_3532,N_3943);
and U4907 (N_4907,N_3334,N_3506);
and U4908 (N_4908,N_3973,N_3730);
nand U4909 (N_4909,N_3882,N_3301);
or U4910 (N_4910,N_3891,N_3146);
xor U4911 (N_4911,N_3310,N_3820);
and U4912 (N_4912,N_3893,N_3960);
nand U4913 (N_4913,N_3066,N_3172);
nand U4914 (N_4914,N_3695,N_3536);
or U4915 (N_4915,N_3317,N_3111);
nor U4916 (N_4916,N_3492,N_3923);
or U4917 (N_4917,N_3917,N_3112);
nand U4918 (N_4918,N_3721,N_3596);
and U4919 (N_4919,N_3952,N_3503);
nand U4920 (N_4920,N_3176,N_3682);
nor U4921 (N_4921,N_3053,N_3631);
xor U4922 (N_4922,N_3036,N_3425);
nor U4923 (N_4923,N_3700,N_3733);
and U4924 (N_4924,N_3081,N_3837);
or U4925 (N_4925,N_3270,N_3775);
nand U4926 (N_4926,N_3069,N_3328);
and U4927 (N_4927,N_3568,N_3099);
or U4928 (N_4928,N_3578,N_3411);
and U4929 (N_4929,N_3072,N_3108);
or U4930 (N_4930,N_3415,N_3663);
nor U4931 (N_4931,N_3300,N_3350);
nand U4932 (N_4932,N_3108,N_3726);
nor U4933 (N_4933,N_3729,N_3400);
or U4934 (N_4934,N_3996,N_3636);
xnor U4935 (N_4935,N_3627,N_3755);
or U4936 (N_4936,N_3625,N_3857);
xor U4937 (N_4937,N_3703,N_3942);
or U4938 (N_4938,N_3927,N_3178);
nor U4939 (N_4939,N_3824,N_3316);
and U4940 (N_4940,N_3766,N_3836);
or U4941 (N_4941,N_3145,N_3916);
nand U4942 (N_4942,N_3912,N_3740);
nor U4943 (N_4943,N_3229,N_3290);
nor U4944 (N_4944,N_3855,N_3005);
and U4945 (N_4945,N_3245,N_3101);
xnor U4946 (N_4946,N_3881,N_3107);
and U4947 (N_4947,N_3971,N_3057);
nand U4948 (N_4948,N_3585,N_3344);
or U4949 (N_4949,N_3767,N_3788);
nand U4950 (N_4950,N_3720,N_3733);
and U4951 (N_4951,N_3455,N_3378);
nor U4952 (N_4952,N_3328,N_3618);
or U4953 (N_4953,N_3912,N_3502);
nand U4954 (N_4954,N_3866,N_3404);
and U4955 (N_4955,N_3854,N_3726);
and U4956 (N_4956,N_3869,N_3085);
xnor U4957 (N_4957,N_3250,N_3056);
and U4958 (N_4958,N_3839,N_3349);
nand U4959 (N_4959,N_3416,N_3952);
and U4960 (N_4960,N_3883,N_3662);
nor U4961 (N_4961,N_3363,N_3438);
nor U4962 (N_4962,N_3800,N_3593);
or U4963 (N_4963,N_3155,N_3819);
nand U4964 (N_4964,N_3343,N_3008);
nand U4965 (N_4965,N_3852,N_3157);
nor U4966 (N_4966,N_3666,N_3571);
or U4967 (N_4967,N_3260,N_3463);
nor U4968 (N_4968,N_3534,N_3229);
or U4969 (N_4969,N_3245,N_3961);
nor U4970 (N_4970,N_3838,N_3713);
nor U4971 (N_4971,N_3429,N_3292);
nor U4972 (N_4972,N_3466,N_3653);
nor U4973 (N_4973,N_3959,N_3468);
nor U4974 (N_4974,N_3091,N_3018);
xnor U4975 (N_4975,N_3411,N_3779);
or U4976 (N_4976,N_3919,N_3263);
nor U4977 (N_4977,N_3503,N_3569);
nor U4978 (N_4978,N_3206,N_3466);
and U4979 (N_4979,N_3569,N_3554);
or U4980 (N_4980,N_3400,N_3144);
and U4981 (N_4981,N_3346,N_3568);
or U4982 (N_4982,N_3920,N_3614);
nand U4983 (N_4983,N_3487,N_3784);
and U4984 (N_4984,N_3480,N_3933);
nand U4985 (N_4985,N_3377,N_3045);
xnor U4986 (N_4986,N_3709,N_3345);
or U4987 (N_4987,N_3184,N_3933);
nand U4988 (N_4988,N_3777,N_3217);
and U4989 (N_4989,N_3969,N_3383);
and U4990 (N_4990,N_3056,N_3893);
and U4991 (N_4991,N_3636,N_3864);
and U4992 (N_4992,N_3951,N_3327);
nor U4993 (N_4993,N_3631,N_3651);
and U4994 (N_4994,N_3890,N_3507);
nand U4995 (N_4995,N_3233,N_3699);
and U4996 (N_4996,N_3304,N_3091);
and U4997 (N_4997,N_3030,N_3350);
nor U4998 (N_4998,N_3211,N_3968);
nor U4999 (N_4999,N_3593,N_3190);
xnor U5000 (N_5000,N_4954,N_4669);
or U5001 (N_5001,N_4958,N_4955);
nor U5002 (N_5002,N_4066,N_4260);
xor U5003 (N_5003,N_4381,N_4079);
and U5004 (N_5004,N_4091,N_4598);
xor U5005 (N_5005,N_4285,N_4440);
xnor U5006 (N_5006,N_4406,N_4607);
nor U5007 (N_5007,N_4127,N_4554);
or U5008 (N_5008,N_4973,N_4452);
nor U5009 (N_5009,N_4347,N_4370);
xor U5010 (N_5010,N_4070,N_4307);
and U5011 (N_5011,N_4912,N_4418);
nand U5012 (N_5012,N_4638,N_4969);
nor U5013 (N_5013,N_4610,N_4466);
xnor U5014 (N_5014,N_4795,N_4908);
and U5015 (N_5015,N_4504,N_4957);
xor U5016 (N_5016,N_4904,N_4422);
nand U5017 (N_5017,N_4575,N_4629);
or U5018 (N_5018,N_4801,N_4978);
nor U5019 (N_5019,N_4753,N_4552);
or U5020 (N_5020,N_4008,N_4930);
or U5021 (N_5021,N_4691,N_4674);
and U5022 (N_5022,N_4322,N_4605);
or U5023 (N_5023,N_4541,N_4965);
xor U5024 (N_5024,N_4297,N_4301);
or U5025 (N_5025,N_4027,N_4025);
xor U5026 (N_5026,N_4895,N_4609);
xor U5027 (N_5027,N_4337,N_4007);
nor U5028 (N_5028,N_4961,N_4011);
and U5029 (N_5029,N_4256,N_4359);
nand U5030 (N_5030,N_4253,N_4143);
xor U5031 (N_5031,N_4572,N_4619);
nand U5032 (N_5032,N_4524,N_4796);
or U5033 (N_5033,N_4195,N_4875);
nor U5034 (N_5034,N_4684,N_4162);
nand U5035 (N_5035,N_4456,N_4943);
nor U5036 (N_5036,N_4232,N_4647);
and U5037 (N_5037,N_4124,N_4457);
and U5038 (N_5038,N_4243,N_4509);
xnor U5039 (N_5039,N_4306,N_4389);
nor U5040 (N_5040,N_4172,N_4246);
xnor U5041 (N_5041,N_4938,N_4198);
and U5042 (N_5042,N_4502,N_4429);
nand U5043 (N_5043,N_4272,N_4491);
or U5044 (N_5044,N_4987,N_4262);
or U5045 (N_5045,N_4342,N_4014);
nor U5046 (N_5046,N_4850,N_4661);
and U5047 (N_5047,N_4768,N_4146);
and U5048 (N_5048,N_4785,N_4588);
and U5049 (N_5049,N_4950,N_4542);
nor U5050 (N_5050,N_4486,N_4846);
xor U5051 (N_5051,N_4992,N_4341);
nor U5052 (N_5052,N_4516,N_4681);
and U5053 (N_5053,N_4882,N_4731);
nor U5054 (N_5054,N_4196,N_4676);
xor U5055 (N_5055,N_4211,N_4490);
and U5056 (N_5056,N_4383,N_4784);
nor U5057 (N_5057,N_4547,N_4929);
nor U5058 (N_5058,N_4225,N_4927);
or U5059 (N_5059,N_4845,N_4385);
nor U5060 (N_5060,N_4841,N_4743);
nand U5061 (N_5061,N_4577,N_4374);
or U5062 (N_5062,N_4058,N_4673);
xor U5063 (N_5063,N_4224,N_4264);
or U5064 (N_5064,N_4686,N_4781);
nand U5065 (N_5065,N_4106,N_4703);
and U5066 (N_5066,N_4964,N_4290);
nand U5067 (N_5067,N_4094,N_4428);
or U5068 (N_5068,N_4453,N_4069);
xnor U5069 (N_5069,N_4960,N_4581);
xor U5070 (N_5070,N_4261,N_4117);
xor U5071 (N_5071,N_4037,N_4849);
and U5072 (N_5072,N_4537,N_4837);
nor U5073 (N_5073,N_4983,N_4847);
xnor U5074 (N_5074,N_4636,N_4273);
nor U5075 (N_5075,N_4741,N_4320);
or U5076 (N_5076,N_4518,N_4152);
and U5077 (N_5077,N_4072,N_4494);
and U5078 (N_5078,N_4183,N_4748);
xnor U5079 (N_5079,N_4650,N_4121);
xnor U5080 (N_5080,N_4632,N_4639);
or U5081 (N_5081,N_4171,N_4956);
xor U5082 (N_5082,N_4065,N_4874);
xor U5083 (N_5083,N_4915,N_4946);
or U5084 (N_5084,N_4551,N_4207);
xnor U5085 (N_5085,N_4334,N_4568);
or U5086 (N_5086,N_4254,N_4028);
nor U5087 (N_5087,N_4009,N_4852);
nor U5088 (N_5088,N_4061,N_4530);
and U5089 (N_5089,N_4570,N_4561);
xnor U5090 (N_5090,N_4996,N_4396);
and U5091 (N_5091,N_4214,N_4371);
nand U5092 (N_5092,N_4208,N_4591);
xnor U5093 (N_5093,N_4696,N_4595);
nand U5094 (N_5094,N_4085,N_4442);
nor U5095 (N_5095,N_4180,N_4154);
and U5096 (N_5096,N_4975,N_4810);
xor U5097 (N_5097,N_4168,N_4077);
nor U5098 (N_5098,N_4791,N_4543);
xnor U5099 (N_5099,N_4545,N_4910);
nor U5100 (N_5100,N_4454,N_4289);
or U5101 (N_5101,N_4574,N_4831);
or U5102 (N_5102,N_4790,N_4878);
and U5103 (N_5103,N_4798,N_4532);
and U5104 (N_5104,N_4515,N_4693);
nand U5105 (N_5105,N_4677,N_4824);
nor U5106 (N_5106,N_4259,N_4567);
xor U5107 (N_5107,N_4078,N_4525);
nand U5108 (N_5108,N_4176,N_4191);
nor U5109 (N_5109,N_4348,N_4046);
nand U5110 (N_5110,N_4872,N_4326);
and U5111 (N_5111,N_4864,N_4974);
or U5112 (N_5112,N_4779,N_4174);
xor U5113 (N_5113,N_4734,N_4199);
nor U5114 (N_5114,N_4404,N_4982);
nor U5115 (N_5115,N_4923,N_4675);
and U5116 (N_5116,N_4646,N_4944);
nor U5117 (N_5117,N_4902,N_4424);
nor U5118 (N_5118,N_4892,N_4001);
or U5119 (N_5119,N_4080,N_4692);
xnor U5120 (N_5120,N_4862,N_4933);
xnor U5121 (N_5121,N_4576,N_4680);
nor U5122 (N_5122,N_4776,N_4349);
nor U5123 (N_5123,N_4156,N_4287);
nor U5124 (N_5124,N_4514,N_4459);
and U5125 (N_5125,N_4830,N_4817);
nand U5126 (N_5126,N_4031,N_4412);
nand U5127 (N_5127,N_4986,N_4690);
xor U5128 (N_5128,N_4203,N_4278);
or U5129 (N_5129,N_4701,N_4060);
xnor U5130 (N_5130,N_4835,N_4787);
xnor U5131 (N_5131,N_4750,N_4251);
nand U5132 (N_5132,N_4186,N_4310);
nor U5133 (N_5133,N_4427,N_4193);
xnor U5134 (N_5134,N_4299,N_4110);
nand U5135 (N_5135,N_4388,N_4062);
or U5136 (N_5136,N_4737,N_4484);
and U5137 (N_5137,N_4560,N_4147);
nor U5138 (N_5138,N_4922,N_4599);
nor U5139 (N_5139,N_4997,N_4096);
and U5140 (N_5140,N_4901,N_4237);
nand U5141 (N_5141,N_4697,N_4479);
nand U5142 (N_5142,N_4399,N_4369);
xor U5143 (N_5143,N_4707,N_4338);
nor U5144 (N_5144,N_4336,N_4064);
and U5145 (N_5145,N_4135,N_4648);
nand U5146 (N_5146,N_4470,N_4282);
nor U5147 (N_5147,N_4662,N_4402);
nor U5148 (N_5148,N_4308,N_4688);
nor U5149 (N_5149,N_4103,N_4618);
or U5150 (N_5150,N_4582,N_4393);
nor U5151 (N_5151,N_4709,N_4055);
nor U5152 (N_5152,N_4573,N_4002);
and U5153 (N_5153,N_4372,N_4565);
and U5154 (N_5154,N_4050,N_4919);
nor U5155 (N_5155,N_4765,N_4119);
and U5156 (N_5156,N_4722,N_4640);
or U5157 (N_5157,N_4694,N_4770);
and U5158 (N_5158,N_4536,N_4434);
xor U5159 (N_5159,N_4894,N_4660);
nor U5160 (N_5160,N_4248,N_4441);
xnor U5161 (N_5161,N_4507,N_4728);
or U5162 (N_5162,N_4405,N_4600);
nor U5163 (N_5163,N_4948,N_4040);
nor U5164 (N_5164,N_4090,N_4579);
nor U5165 (N_5165,N_4578,N_4130);
nor U5166 (N_5166,N_4084,N_4799);
and U5167 (N_5167,N_4730,N_4448);
and U5168 (N_5168,N_4968,N_4473);
nor U5169 (N_5169,N_4111,N_4052);
nor U5170 (N_5170,N_4082,N_4458);
and U5171 (N_5171,N_4655,N_4021);
xor U5172 (N_5172,N_4433,N_4339);
nand U5173 (N_5173,N_4813,N_4221);
xnor U5174 (N_5174,N_4746,N_4379);
nand U5175 (N_5175,N_4989,N_4220);
nand U5176 (N_5176,N_4148,N_4833);
or U5177 (N_5177,N_4380,N_4634);
or U5178 (N_5178,N_4375,N_4866);
xnor U5179 (N_5179,N_4526,N_4410);
nand U5180 (N_5180,N_4329,N_4447);
nand U5181 (N_5181,N_4140,N_4777);
nor U5182 (N_5182,N_4268,N_4580);
or U5183 (N_5183,N_4086,N_4937);
or U5184 (N_5184,N_4421,N_4343);
xor U5185 (N_5185,N_4840,N_4335);
nor U5186 (N_5186,N_4877,N_4719);
nor U5187 (N_5187,N_4825,N_4718);
or U5188 (N_5188,N_4685,N_4498);
and U5189 (N_5189,N_4544,N_4962);
nor U5190 (N_5190,N_4108,N_4275);
nand U5191 (N_5191,N_4775,N_4330);
nor U5192 (N_5192,N_4012,N_4182);
and U5193 (N_5193,N_4144,N_4981);
nor U5194 (N_5194,N_4557,N_4250);
and U5195 (N_5195,N_4528,N_4185);
and U5196 (N_5196,N_4708,N_4621);
and U5197 (N_5197,N_4823,N_4668);
xor U5198 (N_5198,N_4226,N_4026);
or U5199 (N_5199,N_4449,N_4257);
or U5200 (N_5200,N_4157,N_4240);
nor U5201 (N_5201,N_4683,N_4294);
nand U5202 (N_5202,N_4415,N_4202);
nand U5203 (N_5203,N_4711,N_4303);
or U5204 (N_5204,N_4286,N_4888);
and U5205 (N_5205,N_4539,N_4317);
nor U5206 (N_5206,N_4714,N_4102);
nand U5207 (N_5207,N_4219,N_4553);
nor U5208 (N_5208,N_4505,N_4201);
nor U5209 (N_5209,N_4137,N_4819);
nand U5210 (N_5210,N_4903,N_4178);
and U5211 (N_5211,N_4047,N_4395);
and U5212 (N_5212,N_4721,N_4990);
nand U5213 (N_5213,N_4327,N_4735);
xnor U5214 (N_5214,N_4266,N_4726);
nand U5215 (N_5215,N_4107,N_4885);
nand U5216 (N_5216,N_4120,N_4985);
and U5217 (N_5217,N_4401,N_4928);
or U5218 (N_5218,N_4408,N_4942);
xor U5219 (N_5219,N_4503,N_4476);
or U5220 (N_5220,N_4175,N_4030);
nand U5221 (N_5221,N_4717,N_4361);
nand U5222 (N_5222,N_4896,N_4884);
and U5223 (N_5223,N_4481,N_4851);
nand U5224 (N_5224,N_4426,N_4994);
nand U5225 (N_5225,N_4350,N_4854);
or U5226 (N_5226,N_4043,N_4450);
and U5227 (N_5227,N_4419,N_4315);
xor U5228 (N_5228,N_4867,N_4756);
nand U5229 (N_5229,N_4533,N_4739);
or U5230 (N_5230,N_4075,N_4853);
nor U5231 (N_5231,N_4036,N_4856);
xnor U5232 (N_5232,N_4056,N_4133);
xnor U5233 (N_5233,N_4635,N_4935);
xnor U5234 (N_5234,N_4963,N_4794);
nor U5235 (N_5235,N_4751,N_4475);
xor U5236 (N_5236,N_4644,N_4270);
nand U5237 (N_5237,N_4625,N_4384);
or U5238 (N_5238,N_4988,N_4455);
nand U5239 (N_5239,N_4305,N_4059);
and U5240 (N_5240,N_4742,N_4815);
and U5241 (N_5241,N_4952,N_4754);
and U5242 (N_5242,N_4416,N_4637);
nor U5243 (N_5243,N_4497,N_4967);
and U5244 (N_5244,N_4564,N_4160);
or U5245 (N_5245,N_4816,N_4020);
nor U5246 (N_5246,N_4229,N_4436);
nor U5247 (N_5247,N_4772,N_4015);
or U5248 (N_5248,N_4870,N_4814);
and U5249 (N_5249,N_4925,N_4767);
nand U5250 (N_5250,N_4909,N_4489);
or U5251 (N_5251,N_4465,N_4809);
xor U5252 (N_5252,N_4071,N_4019);
nand U5253 (N_5253,N_4720,N_4354);
or U5254 (N_5254,N_4880,N_4757);
nor U5255 (N_5255,N_4774,N_4093);
nand U5256 (N_5256,N_4344,N_4227);
nor U5257 (N_5257,N_4116,N_4540);
nor U5258 (N_5258,N_4122,N_4432);
nand U5259 (N_5259,N_4420,N_4736);
or U5260 (N_5260,N_4241,N_4245);
nand U5261 (N_5261,N_4562,N_4889);
or U5262 (N_5262,N_4187,N_4067);
xnor U5263 (N_5263,N_4594,N_4871);
xor U5264 (N_5264,N_4920,N_4463);
nor U5265 (N_5265,N_4861,N_4620);
or U5266 (N_5266,N_4704,N_4488);
nand U5267 (N_5267,N_4869,N_4493);
nor U5268 (N_5268,N_4284,N_4971);
nor U5269 (N_5269,N_4670,N_4511);
nand U5270 (N_5270,N_4197,N_4807);
nor U5271 (N_5271,N_4702,N_4265);
nor U5272 (N_5272,N_4271,N_4048);
or U5273 (N_5273,N_4951,N_4480);
nand U5274 (N_5274,N_4045,N_4585);
xnor U5275 (N_5275,N_4423,N_4766);
nor U5276 (N_5276,N_4771,N_4368);
and U5277 (N_5277,N_4510,N_4729);
nand U5278 (N_5278,N_4656,N_4900);
and U5279 (N_5279,N_4394,N_4312);
nand U5280 (N_5280,N_4478,N_4659);
xnor U5281 (N_5281,N_4018,N_4141);
xor U5282 (N_5282,N_4941,N_4976);
or U5283 (N_5283,N_4612,N_4710);
nand U5284 (N_5284,N_4083,N_4804);
nand U5285 (N_5285,N_4319,N_4555);
nor U5286 (N_5286,N_4517,N_4727);
nand U5287 (N_5287,N_4977,N_4806);
nand U5288 (N_5288,N_4715,N_4838);
nand U5289 (N_5289,N_4550,N_4044);
nand U5290 (N_5290,N_4189,N_4166);
nor U5291 (N_5291,N_4364,N_4664);
or U5292 (N_5292,N_4616,N_4378);
or U5293 (N_5293,N_4430,N_4602);
or U5294 (N_5294,N_4842,N_4812);
nor U5295 (N_5295,N_4357,N_4355);
and U5296 (N_5296,N_4017,N_4939);
and U5297 (N_5297,N_4913,N_4628);
nand U5298 (N_5298,N_4365,N_4035);
nor U5299 (N_5299,N_4800,N_4700);
xnor U5300 (N_5300,N_4444,N_4288);
nor U5301 (N_5301,N_4844,N_4216);
and U5302 (N_5302,N_4006,N_4145);
xor U5303 (N_5303,N_4758,N_4387);
xnor U5304 (N_5304,N_4808,N_4414);
and U5305 (N_5305,N_4863,N_4991);
and U5306 (N_5306,N_4911,N_4471);
nor U5307 (N_5307,N_4522,N_4811);
nand U5308 (N_5308,N_4013,N_4860);
and U5309 (N_5309,N_4993,N_4949);
and U5310 (N_5310,N_4906,N_4435);
or U5311 (N_5311,N_4099,N_4249);
xnor U5312 (N_5312,N_4425,N_4645);
xor U5313 (N_5313,N_4611,N_4164);
xor U5314 (N_5314,N_4897,N_4010);
and U5315 (N_5315,N_4280,N_4445);
xor U5316 (N_5316,N_4192,N_4678);
or U5317 (N_5317,N_4382,N_4293);
nand U5318 (N_5318,N_4786,N_4366);
xnor U5319 (N_5319,N_4105,N_4403);
and U5320 (N_5320,N_4725,N_4699);
xnor U5321 (N_5321,N_4321,N_4205);
xor U5322 (N_5322,N_4608,N_4512);
nand U5323 (N_5323,N_4376,N_4821);
nor U5324 (N_5324,N_4829,N_4797);
or U5325 (N_5325,N_4613,N_4496);
xnor U5326 (N_5326,N_4109,N_4331);
nand U5327 (N_5327,N_4666,N_4360);
xor U5328 (N_5328,N_4995,N_4151);
nor U5329 (N_5329,N_4460,N_4390);
xnor U5330 (N_5330,N_4793,N_4206);
nand U5331 (N_5331,N_4857,N_4115);
nor U5332 (N_5332,N_4231,N_4098);
and U5333 (N_5333,N_4828,N_4104);
xnor U5334 (N_5334,N_4534,N_4859);
or U5335 (N_5335,N_4004,N_4467);
and U5336 (N_5336,N_4641,N_4789);
or U5337 (N_5337,N_4752,N_4559);
xnor U5338 (N_5338,N_4477,N_4153);
and U5339 (N_5339,N_4820,N_4302);
or U5340 (N_5340,N_4836,N_4333);
or U5341 (N_5341,N_4318,N_4931);
xor U5342 (N_5342,N_4234,N_4034);
nand U5343 (N_5343,N_4316,N_4215);
and U5344 (N_5344,N_4500,N_4966);
or U5345 (N_5345,N_4617,N_4917);
nor U5346 (N_5346,N_4188,N_4716);
or U5347 (N_5347,N_4563,N_4095);
nand U5348 (N_5348,N_4918,N_4643);
xor U5349 (N_5349,N_4170,N_4745);
and U5350 (N_5350,N_4980,N_4469);
nor U5351 (N_5351,N_4397,N_4546);
and U5352 (N_5352,N_4883,N_4267);
nor U5353 (N_5353,N_4413,N_4165);
and U5354 (N_5354,N_4592,N_4778);
xnor U5355 (N_5355,N_4114,N_4843);
and U5356 (N_5356,N_4129,N_4300);
nand U5357 (N_5357,N_4868,N_4506);
xor U5358 (N_5358,N_4088,N_4053);
nor U5359 (N_5359,N_4029,N_4295);
nand U5360 (N_5360,N_4163,N_4003);
nand U5361 (N_5361,N_4571,N_4914);
and U5362 (N_5362,N_4805,N_4332);
or U5363 (N_5363,N_4926,N_4092);
nor U5364 (N_5364,N_4657,N_4311);
nor U5365 (N_5365,N_4244,N_4905);
nand U5366 (N_5366,N_4247,N_4826);
nor U5367 (N_5367,N_4113,N_4566);
nor U5368 (N_5368,N_4626,N_4590);
nor U5369 (N_5369,N_4865,N_4642);
and U5370 (N_5370,N_4529,N_4438);
nor U5371 (N_5371,N_4346,N_4184);
or U5372 (N_5372,N_4016,N_4916);
or U5373 (N_5373,N_4472,N_4296);
nand U5374 (N_5374,N_4947,N_4839);
nor U5375 (N_5375,N_4169,N_4269);
xor U5376 (N_5376,N_4367,N_4936);
xnor U5377 (N_5377,N_4593,N_4309);
and U5378 (N_5378,N_4125,N_4858);
nor U5379 (N_5379,N_4682,N_4446);
nand U5380 (N_5380,N_4687,N_4932);
or U5381 (N_5381,N_4051,N_4398);
and U5382 (N_5382,N_4161,N_4213);
xnor U5383 (N_5383,N_4462,N_4788);
and U5384 (N_5384,N_4358,N_4508);
and U5385 (N_5385,N_4597,N_4194);
xor U5386 (N_5386,N_4706,N_4780);
nor U5387 (N_5387,N_4689,N_4042);
and U5388 (N_5388,N_4138,N_4304);
nor U5389 (N_5389,N_4970,N_4487);
or U5390 (N_5390,N_4671,N_4217);
nor U5391 (N_5391,N_4832,N_4654);
xnor U5392 (N_5392,N_4615,N_4179);
xnor U5393 (N_5393,N_4136,N_4118);
xor U5394 (N_5394,N_4238,N_4601);
or U5395 (N_5395,N_4520,N_4167);
and U5396 (N_5396,N_4313,N_4940);
and U5397 (N_5397,N_4899,N_4755);
nand U5398 (N_5398,N_4898,N_4822);
nand U5399 (N_5399,N_4150,N_4979);
nand U5400 (N_5400,N_4523,N_4101);
or U5401 (N_5401,N_4492,N_4235);
nand U5402 (N_5402,N_4891,N_4439);
nand U5403 (N_5403,N_4209,N_4112);
or U5404 (N_5404,N_4222,N_4377);
xor U5405 (N_5405,N_4998,N_4263);
nand U5406 (N_5406,N_4057,N_4584);
xnor U5407 (N_5407,N_4945,N_4392);
nand U5408 (N_5408,N_4291,N_4212);
or U5409 (N_5409,N_4074,N_4210);
nor U5410 (N_5410,N_4005,N_4100);
xnor U5411 (N_5411,N_4651,N_4759);
nand U5412 (N_5412,N_4614,N_4782);
or U5413 (N_5413,N_4959,N_4818);
or U5414 (N_5414,N_4658,N_4649);
nand U5415 (N_5415,N_4972,N_4190);
or U5416 (N_5416,N_4200,N_4893);
xor U5417 (N_5417,N_4173,N_4749);
xor U5418 (N_5418,N_4834,N_4352);
or U5419 (N_5419,N_4242,N_4277);
nand U5420 (N_5420,N_4876,N_4073);
nor U5421 (N_5421,N_4292,N_4740);
xnor U5422 (N_5422,N_4236,N_4783);
or U5423 (N_5423,N_4417,N_4233);
and U5424 (N_5424,N_4032,N_4076);
xor U5425 (N_5425,N_4633,N_4323);
or U5426 (N_5426,N_4953,N_4386);
or U5427 (N_5427,N_4848,N_4769);
and U5428 (N_5428,N_4063,N_4501);
nor U5429 (N_5429,N_4744,N_4999);
or U5430 (N_5430,N_4033,N_4142);
or U5431 (N_5431,N_4230,N_4698);
xor U5432 (N_5432,N_4606,N_4855);
and U5433 (N_5433,N_4732,N_4747);
xnor U5434 (N_5434,N_4556,N_4622);
xor U5435 (N_5435,N_4177,N_4762);
xor U5436 (N_5436,N_4362,N_4934);
or U5437 (N_5437,N_4391,N_4039);
and U5438 (N_5438,N_4924,N_4764);
and U5439 (N_5439,N_4713,N_4023);
and U5440 (N_5440,N_4483,N_4155);
or U5441 (N_5441,N_4218,N_4627);
xor U5442 (N_5442,N_4283,N_4586);
nand U5443 (N_5443,N_4667,N_4604);
nor U5444 (N_5444,N_4279,N_4723);
or U5445 (N_5445,N_4400,N_4631);
nand U5446 (N_5446,N_4761,N_4134);
xnor U5447 (N_5447,N_4873,N_4589);
xor U5448 (N_5448,N_4724,N_4624);
or U5449 (N_5449,N_4760,N_4679);
nor U5450 (N_5450,N_4773,N_4068);
and U5451 (N_5451,N_4128,N_4464);
or U5452 (N_5452,N_4695,N_4054);
or U5453 (N_5453,N_4325,N_4886);
or U5454 (N_5454,N_4274,N_4623);
nor U5455 (N_5455,N_4583,N_4519);
and U5456 (N_5456,N_4738,N_4131);
xnor U5457 (N_5457,N_4663,N_4373);
and U5458 (N_5458,N_4596,N_4569);
and U5459 (N_5459,N_4468,N_4827);
and U5460 (N_5460,N_4411,N_4351);
nand U5461 (N_5461,N_4356,N_4409);
nand U5462 (N_5462,N_4363,N_4081);
or U5463 (N_5463,N_4603,N_4665);
xnor U5464 (N_5464,N_4087,N_4437);
xor U5465 (N_5465,N_4474,N_4041);
and U5466 (N_5466,N_4792,N_4881);
and U5467 (N_5467,N_4239,N_4548);
xor U5468 (N_5468,N_4298,N_4049);
nand U5469 (N_5469,N_4803,N_4123);
xnor U5470 (N_5470,N_4921,N_4802);
nor U5471 (N_5471,N_4538,N_4984);
xnor U5472 (N_5472,N_4451,N_4204);
and U5473 (N_5473,N_4879,N_4672);
nand U5474 (N_5474,N_4705,N_4255);
and U5475 (N_5475,N_4258,N_4907);
xor U5476 (N_5476,N_4890,N_4630);
or U5477 (N_5477,N_4407,N_4558);
xor U5478 (N_5478,N_4887,N_4328);
xor U5479 (N_5479,N_4712,N_4314);
or U5480 (N_5480,N_4653,N_4527);
and U5481 (N_5481,N_4521,N_4097);
xnor U5482 (N_5482,N_4531,N_4038);
nor U5483 (N_5483,N_4461,N_4733);
nor U5484 (N_5484,N_4353,N_4340);
and U5485 (N_5485,N_4345,N_4495);
nor U5486 (N_5486,N_4000,N_4513);
xor U5487 (N_5487,N_4022,N_4139);
and U5488 (N_5488,N_4535,N_4276);
xnor U5489 (N_5489,N_4431,N_4482);
nand U5490 (N_5490,N_4126,N_4324);
nor U5491 (N_5491,N_4089,N_4485);
or U5492 (N_5492,N_4652,N_4024);
or U5493 (N_5493,N_4159,N_4228);
xor U5494 (N_5494,N_4549,N_4499);
or U5495 (N_5495,N_4223,N_4281);
and U5496 (N_5496,N_4587,N_4181);
and U5497 (N_5497,N_4252,N_4149);
xor U5498 (N_5498,N_4132,N_4443);
nor U5499 (N_5499,N_4158,N_4763);
xor U5500 (N_5500,N_4946,N_4560);
or U5501 (N_5501,N_4591,N_4206);
or U5502 (N_5502,N_4431,N_4904);
and U5503 (N_5503,N_4817,N_4266);
and U5504 (N_5504,N_4153,N_4585);
nor U5505 (N_5505,N_4225,N_4342);
or U5506 (N_5506,N_4654,N_4465);
xnor U5507 (N_5507,N_4133,N_4864);
and U5508 (N_5508,N_4337,N_4637);
or U5509 (N_5509,N_4451,N_4939);
or U5510 (N_5510,N_4923,N_4636);
nand U5511 (N_5511,N_4986,N_4594);
or U5512 (N_5512,N_4660,N_4962);
nor U5513 (N_5513,N_4123,N_4871);
nand U5514 (N_5514,N_4892,N_4466);
nor U5515 (N_5515,N_4775,N_4667);
nand U5516 (N_5516,N_4790,N_4349);
xnor U5517 (N_5517,N_4493,N_4741);
xor U5518 (N_5518,N_4129,N_4718);
and U5519 (N_5519,N_4162,N_4665);
or U5520 (N_5520,N_4307,N_4040);
xor U5521 (N_5521,N_4293,N_4726);
or U5522 (N_5522,N_4647,N_4943);
nor U5523 (N_5523,N_4390,N_4900);
nor U5524 (N_5524,N_4290,N_4168);
xor U5525 (N_5525,N_4349,N_4148);
nand U5526 (N_5526,N_4516,N_4267);
nor U5527 (N_5527,N_4411,N_4871);
xnor U5528 (N_5528,N_4200,N_4057);
or U5529 (N_5529,N_4129,N_4275);
xnor U5530 (N_5530,N_4400,N_4886);
nand U5531 (N_5531,N_4512,N_4533);
or U5532 (N_5532,N_4439,N_4909);
nor U5533 (N_5533,N_4072,N_4213);
nor U5534 (N_5534,N_4825,N_4962);
nor U5535 (N_5535,N_4005,N_4630);
or U5536 (N_5536,N_4754,N_4084);
and U5537 (N_5537,N_4570,N_4928);
nor U5538 (N_5538,N_4486,N_4786);
or U5539 (N_5539,N_4230,N_4692);
xor U5540 (N_5540,N_4202,N_4521);
and U5541 (N_5541,N_4910,N_4370);
and U5542 (N_5542,N_4079,N_4484);
nand U5543 (N_5543,N_4083,N_4392);
nand U5544 (N_5544,N_4895,N_4302);
or U5545 (N_5545,N_4546,N_4074);
nand U5546 (N_5546,N_4973,N_4014);
and U5547 (N_5547,N_4380,N_4038);
nor U5548 (N_5548,N_4887,N_4555);
or U5549 (N_5549,N_4571,N_4044);
or U5550 (N_5550,N_4623,N_4356);
and U5551 (N_5551,N_4811,N_4719);
xor U5552 (N_5552,N_4400,N_4855);
and U5553 (N_5553,N_4650,N_4874);
or U5554 (N_5554,N_4776,N_4388);
xor U5555 (N_5555,N_4738,N_4559);
xnor U5556 (N_5556,N_4027,N_4372);
nand U5557 (N_5557,N_4907,N_4868);
and U5558 (N_5558,N_4810,N_4267);
and U5559 (N_5559,N_4655,N_4062);
nor U5560 (N_5560,N_4735,N_4981);
xor U5561 (N_5561,N_4758,N_4081);
and U5562 (N_5562,N_4924,N_4125);
xnor U5563 (N_5563,N_4931,N_4104);
xnor U5564 (N_5564,N_4916,N_4517);
or U5565 (N_5565,N_4110,N_4468);
and U5566 (N_5566,N_4159,N_4560);
xor U5567 (N_5567,N_4774,N_4430);
nor U5568 (N_5568,N_4679,N_4205);
nor U5569 (N_5569,N_4252,N_4263);
nand U5570 (N_5570,N_4591,N_4520);
nand U5571 (N_5571,N_4577,N_4110);
nor U5572 (N_5572,N_4589,N_4881);
or U5573 (N_5573,N_4528,N_4647);
nand U5574 (N_5574,N_4540,N_4441);
nand U5575 (N_5575,N_4259,N_4985);
and U5576 (N_5576,N_4895,N_4062);
and U5577 (N_5577,N_4114,N_4794);
nor U5578 (N_5578,N_4104,N_4821);
xor U5579 (N_5579,N_4206,N_4466);
nand U5580 (N_5580,N_4956,N_4721);
or U5581 (N_5581,N_4968,N_4204);
xor U5582 (N_5582,N_4822,N_4602);
xor U5583 (N_5583,N_4932,N_4170);
and U5584 (N_5584,N_4801,N_4513);
nor U5585 (N_5585,N_4214,N_4335);
or U5586 (N_5586,N_4725,N_4536);
xor U5587 (N_5587,N_4832,N_4094);
or U5588 (N_5588,N_4961,N_4812);
xor U5589 (N_5589,N_4278,N_4126);
and U5590 (N_5590,N_4592,N_4168);
nor U5591 (N_5591,N_4985,N_4580);
and U5592 (N_5592,N_4620,N_4989);
and U5593 (N_5593,N_4765,N_4619);
nand U5594 (N_5594,N_4584,N_4685);
xnor U5595 (N_5595,N_4900,N_4522);
nor U5596 (N_5596,N_4609,N_4525);
or U5597 (N_5597,N_4578,N_4344);
and U5598 (N_5598,N_4973,N_4961);
nand U5599 (N_5599,N_4467,N_4633);
nor U5600 (N_5600,N_4722,N_4875);
xnor U5601 (N_5601,N_4542,N_4819);
or U5602 (N_5602,N_4194,N_4323);
or U5603 (N_5603,N_4560,N_4063);
xnor U5604 (N_5604,N_4870,N_4861);
xnor U5605 (N_5605,N_4729,N_4148);
and U5606 (N_5606,N_4199,N_4875);
or U5607 (N_5607,N_4459,N_4423);
nand U5608 (N_5608,N_4735,N_4526);
xor U5609 (N_5609,N_4946,N_4585);
xnor U5610 (N_5610,N_4439,N_4558);
and U5611 (N_5611,N_4057,N_4777);
nor U5612 (N_5612,N_4446,N_4560);
or U5613 (N_5613,N_4281,N_4959);
nor U5614 (N_5614,N_4888,N_4488);
and U5615 (N_5615,N_4358,N_4527);
and U5616 (N_5616,N_4275,N_4773);
nor U5617 (N_5617,N_4990,N_4598);
nor U5618 (N_5618,N_4632,N_4113);
or U5619 (N_5619,N_4297,N_4724);
nor U5620 (N_5620,N_4410,N_4578);
and U5621 (N_5621,N_4371,N_4578);
and U5622 (N_5622,N_4294,N_4016);
and U5623 (N_5623,N_4707,N_4139);
or U5624 (N_5624,N_4882,N_4110);
nor U5625 (N_5625,N_4705,N_4411);
and U5626 (N_5626,N_4714,N_4976);
and U5627 (N_5627,N_4116,N_4375);
nor U5628 (N_5628,N_4401,N_4167);
or U5629 (N_5629,N_4827,N_4125);
or U5630 (N_5630,N_4186,N_4596);
and U5631 (N_5631,N_4311,N_4855);
nor U5632 (N_5632,N_4840,N_4009);
and U5633 (N_5633,N_4713,N_4315);
nand U5634 (N_5634,N_4641,N_4181);
nand U5635 (N_5635,N_4547,N_4078);
xnor U5636 (N_5636,N_4442,N_4959);
xnor U5637 (N_5637,N_4550,N_4492);
xnor U5638 (N_5638,N_4726,N_4304);
and U5639 (N_5639,N_4783,N_4737);
and U5640 (N_5640,N_4509,N_4257);
and U5641 (N_5641,N_4650,N_4120);
xnor U5642 (N_5642,N_4114,N_4028);
nand U5643 (N_5643,N_4264,N_4019);
xor U5644 (N_5644,N_4233,N_4586);
and U5645 (N_5645,N_4465,N_4850);
and U5646 (N_5646,N_4644,N_4927);
nor U5647 (N_5647,N_4652,N_4422);
xor U5648 (N_5648,N_4688,N_4622);
nand U5649 (N_5649,N_4126,N_4628);
or U5650 (N_5650,N_4567,N_4171);
or U5651 (N_5651,N_4087,N_4239);
nor U5652 (N_5652,N_4675,N_4182);
and U5653 (N_5653,N_4269,N_4352);
nand U5654 (N_5654,N_4432,N_4799);
and U5655 (N_5655,N_4108,N_4594);
nand U5656 (N_5656,N_4782,N_4095);
nand U5657 (N_5657,N_4882,N_4071);
xnor U5658 (N_5658,N_4576,N_4950);
or U5659 (N_5659,N_4892,N_4705);
and U5660 (N_5660,N_4677,N_4007);
or U5661 (N_5661,N_4958,N_4806);
and U5662 (N_5662,N_4960,N_4715);
nor U5663 (N_5663,N_4553,N_4215);
xnor U5664 (N_5664,N_4746,N_4382);
nor U5665 (N_5665,N_4135,N_4138);
and U5666 (N_5666,N_4421,N_4698);
nor U5667 (N_5667,N_4584,N_4647);
xor U5668 (N_5668,N_4348,N_4488);
and U5669 (N_5669,N_4397,N_4663);
and U5670 (N_5670,N_4472,N_4212);
nand U5671 (N_5671,N_4222,N_4233);
nor U5672 (N_5672,N_4721,N_4191);
or U5673 (N_5673,N_4575,N_4318);
nand U5674 (N_5674,N_4342,N_4930);
or U5675 (N_5675,N_4139,N_4847);
nand U5676 (N_5676,N_4508,N_4138);
or U5677 (N_5677,N_4918,N_4110);
xnor U5678 (N_5678,N_4426,N_4012);
and U5679 (N_5679,N_4479,N_4110);
or U5680 (N_5680,N_4474,N_4779);
nand U5681 (N_5681,N_4282,N_4994);
and U5682 (N_5682,N_4737,N_4138);
nand U5683 (N_5683,N_4911,N_4150);
or U5684 (N_5684,N_4014,N_4089);
xor U5685 (N_5685,N_4930,N_4602);
or U5686 (N_5686,N_4813,N_4537);
or U5687 (N_5687,N_4447,N_4659);
nor U5688 (N_5688,N_4684,N_4641);
xnor U5689 (N_5689,N_4279,N_4036);
xor U5690 (N_5690,N_4666,N_4431);
nor U5691 (N_5691,N_4908,N_4602);
nand U5692 (N_5692,N_4587,N_4907);
or U5693 (N_5693,N_4930,N_4434);
nor U5694 (N_5694,N_4105,N_4899);
xor U5695 (N_5695,N_4935,N_4962);
nand U5696 (N_5696,N_4628,N_4021);
xnor U5697 (N_5697,N_4712,N_4723);
nand U5698 (N_5698,N_4355,N_4005);
nand U5699 (N_5699,N_4483,N_4610);
or U5700 (N_5700,N_4532,N_4912);
nor U5701 (N_5701,N_4953,N_4453);
nand U5702 (N_5702,N_4881,N_4049);
and U5703 (N_5703,N_4793,N_4183);
nor U5704 (N_5704,N_4610,N_4537);
xnor U5705 (N_5705,N_4137,N_4424);
and U5706 (N_5706,N_4625,N_4897);
or U5707 (N_5707,N_4830,N_4265);
nand U5708 (N_5708,N_4256,N_4814);
and U5709 (N_5709,N_4235,N_4274);
xor U5710 (N_5710,N_4489,N_4856);
nand U5711 (N_5711,N_4567,N_4468);
xnor U5712 (N_5712,N_4431,N_4441);
nand U5713 (N_5713,N_4906,N_4565);
and U5714 (N_5714,N_4402,N_4504);
nand U5715 (N_5715,N_4194,N_4873);
xor U5716 (N_5716,N_4461,N_4436);
nand U5717 (N_5717,N_4689,N_4069);
nand U5718 (N_5718,N_4985,N_4514);
xnor U5719 (N_5719,N_4936,N_4251);
or U5720 (N_5720,N_4715,N_4046);
and U5721 (N_5721,N_4674,N_4698);
xnor U5722 (N_5722,N_4742,N_4667);
nand U5723 (N_5723,N_4473,N_4276);
xor U5724 (N_5724,N_4619,N_4349);
nor U5725 (N_5725,N_4072,N_4562);
and U5726 (N_5726,N_4562,N_4761);
nand U5727 (N_5727,N_4193,N_4580);
nand U5728 (N_5728,N_4801,N_4453);
nand U5729 (N_5729,N_4937,N_4520);
nor U5730 (N_5730,N_4148,N_4806);
nand U5731 (N_5731,N_4168,N_4136);
nand U5732 (N_5732,N_4059,N_4418);
and U5733 (N_5733,N_4450,N_4078);
nor U5734 (N_5734,N_4783,N_4714);
and U5735 (N_5735,N_4629,N_4874);
or U5736 (N_5736,N_4219,N_4812);
nand U5737 (N_5737,N_4707,N_4370);
xnor U5738 (N_5738,N_4639,N_4495);
or U5739 (N_5739,N_4568,N_4566);
or U5740 (N_5740,N_4825,N_4370);
nand U5741 (N_5741,N_4386,N_4543);
nand U5742 (N_5742,N_4638,N_4053);
nor U5743 (N_5743,N_4324,N_4100);
nor U5744 (N_5744,N_4223,N_4725);
or U5745 (N_5745,N_4209,N_4509);
nand U5746 (N_5746,N_4184,N_4786);
xor U5747 (N_5747,N_4276,N_4476);
and U5748 (N_5748,N_4079,N_4865);
and U5749 (N_5749,N_4449,N_4987);
or U5750 (N_5750,N_4352,N_4714);
and U5751 (N_5751,N_4060,N_4391);
or U5752 (N_5752,N_4933,N_4391);
nor U5753 (N_5753,N_4702,N_4400);
nand U5754 (N_5754,N_4900,N_4959);
nand U5755 (N_5755,N_4618,N_4679);
nor U5756 (N_5756,N_4680,N_4203);
nand U5757 (N_5757,N_4665,N_4983);
or U5758 (N_5758,N_4165,N_4996);
and U5759 (N_5759,N_4766,N_4044);
or U5760 (N_5760,N_4524,N_4813);
nor U5761 (N_5761,N_4498,N_4952);
nor U5762 (N_5762,N_4124,N_4346);
nor U5763 (N_5763,N_4115,N_4240);
xnor U5764 (N_5764,N_4764,N_4685);
and U5765 (N_5765,N_4829,N_4537);
nor U5766 (N_5766,N_4234,N_4396);
and U5767 (N_5767,N_4038,N_4312);
or U5768 (N_5768,N_4779,N_4932);
nand U5769 (N_5769,N_4612,N_4540);
xnor U5770 (N_5770,N_4167,N_4902);
xnor U5771 (N_5771,N_4333,N_4923);
or U5772 (N_5772,N_4022,N_4707);
or U5773 (N_5773,N_4465,N_4497);
xnor U5774 (N_5774,N_4334,N_4531);
xnor U5775 (N_5775,N_4013,N_4739);
or U5776 (N_5776,N_4707,N_4646);
and U5777 (N_5777,N_4453,N_4960);
xnor U5778 (N_5778,N_4142,N_4607);
nand U5779 (N_5779,N_4880,N_4579);
nor U5780 (N_5780,N_4041,N_4731);
xnor U5781 (N_5781,N_4819,N_4421);
and U5782 (N_5782,N_4520,N_4483);
xor U5783 (N_5783,N_4493,N_4450);
xor U5784 (N_5784,N_4100,N_4126);
xnor U5785 (N_5785,N_4131,N_4810);
nor U5786 (N_5786,N_4050,N_4633);
xnor U5787 (N_5787,N_4443,N_4598);
and U5788 (N_5788,N_4255,N_4320);
nand U5789 (N_5789,N_4135,N_4064);
nor U5790 (N_5790,N_4481,N_4920);
and U5791 (N_5791,N_4113,N_4059);
xnor U5792 (N_5792,N_4885,N_4428);
or U5793 (N_5793,N_4277,N_4390);
xnor U5794 (N_5794,N_4333,N_4924);
or U5795 (N_5795,N_4490,N_4330);
nand U5796 (N_5796,N_4882,N_4682);
or U5797 (N_5797,N_4672,N_4905);
and U5798 (N_5798,N_4040,N_4364);
nor U5799 (N_5799,N_4529,N_4573);
xor U5800 (N_5800,N_4379,N_4248);
xnor U5801 (N_5801,N_4026,N_4520);
nand U5802 (N_5802,N_4484,N_4496);
or U5803 (N_5803,N_4158,N_4363);
nand U5804 (N_5804,N_4269,N_4383);
or U5805 (N_5805,N_4790,N_4893);
xor U5806 (N_5806,N_4862,N_4700);
nand U5807 (N_5807,N_4816,N_4717);
nand U5808 (N_5808,N_4082,N_4479);
nand U5809 (N_5809,N_4780,N_4016);
nand U5810 (N_5810,N_4141,N_4690);
nor U5811 (N_5811,N_4368,N_4568);
nor U5812 (N_5812,N_4086,N_4203);
xor U5813 (N_5813,N_4864,N_4284);
nand U5814 (N_5814,N_4234,N_4606);
or U5815 (N_5815,N_4605,N_4304);
and U5816 (N_5816,N_4160,N_4132);
nor U5817 (N_5817,N_4985,N_4835);
nor U5818 (N_5818,N_4666,N_4245);
xor U5819 (N_5819,N_4579,N_4662);
and U5820 (N_5820,N_4507,N_4627);
or U5821 (N_5821,N_4780,N_4286);
nor U5822 (N_5822,N_4564,N_4262);
and U5823 (N_5823,N_4537,N_4517);
nor U5824 (N_5824,N_4827,N_4766);
and U5825 (N_5825,N_4833,N_4272);
or U5826 (N_5826,N_4390,N_4684);
or U5827 (N_5827,N_4279,N_4395);
or U5828 (N_5828,N_4625,N_4965);
or U5829 (N_5829,N_4185,N_4634);
nand U5830 (N_5830,N_4124,N_4141);
xor U5831 (N_5831,N_4544,N_4082);
xnor U5832 (N_5832,N_4564,N_4279);
and U5833 (N_5833,N_4879,N_4705);
xnor U5834 (N_5834,N_4925,N_4074);
and U5835 (N_5835,N_4070,N_4478);
nor U5836 (N_5836,N_4054,N_4105);
nor U5837 (N_5837,N_4629,N_4142);
nand U5838 (N_5838,N_4427,N_4897);
or U5839 (N_5839,N_4396,N_4713);
or U5840 (N_5840,N_4020,N_4850);
nand U5841 (N_5841,N_4855,N_4426);
nor U5842 (N_5842,N_4412,N_4091);
nand U5843 (N_5843,N_4659,N_4945);
and U5844 (N_5844,N_4839,N_4306);
xor U5845 (N_5845,N_4435,N_4282);
xor U5846 (N_5846,N_4656,N_4863);
nand U5847 (N_5847,N_4081,N_4435);
or U5848 (N_5848,N_4193,N_4291);
xor U5849 (N_5849,N_4757,N_4948);
xnor U5850 (N_5850,N_4389,N_4349);
nor U5851 (N_5851,N_4211,N_4544);
xnor U5852 (N_5852,N_4893,N_4801);
xor U5853 (N_5853,N_4454,N_4387);
and U5854 (N_5854,N_4612,N_4140);
nand U5855 (N_5855,N_4703,N_4029);
nor U5856 (N_5856,N_4974,N_4500);
and U5857 (N_5857,N_4643,N_4189);
xnor U5858 (N_5858,N_4576,N_4617);
nor U5859 (N_5859,N_4038,N_4954);
xor U5860 (N_5860,N_4512,N_4477);
or U5861 (N_5861,N_4055,N_4338);
xor U5862 (N_5862,N_4071,N_4469);
xnor U5863 (N_5863,N_4842,N_4681);
or U5864 (N_5864,N_4995,N_4775);
or U5865 (N_5865,N_4728,N_4989);
nand U5866 (N_5866,N_4040,N_4581);
nor U5867 (N_5867,N_4002,N_4675);
xnor U5868 (N_5868,N_4808,N_4890);
xor U5869 (N_5869,N_4079,N_4796);
nand U5870 (N_5870,N_4063,N_4952);
or U5871 (N_5871,N_4103,N_4788);
nand U5872 (N_5872,N_4843,N_4099);
nor U5873 (N_5873,N_4415,N_4954);
nor U5874 (N_5874,N_4867,N_4002);
and U5875 (N_5875,N_4696,N_4917);
xor U5876 (N_5876,N_4595,N_4686);
nor U5877 (N_5877,N_4001,N_4951);
nor U5878 (N_5878,N_4115,N_4820);
nor U5879 (N_5879,N_4023,N_4069);
and U5880 (N_5880,N_4224,N_4183);
or U5881 (N_5881,N_4774,N_4079);
nor U5882 (N_5882,N_4954,N_4293);
nand U5883 (N_5883,N_4583,N_4513);
nor U5884 (N_5884,N_4654,N_4500);
nand U5885 (N_5885,N_4242,N_4056);
nand U5886 (N_5886,N_4011,N_4898);
or U5887 (N_5887,N_4784,N_4835);
or U5888 (N_5888,N_4580,N_4741);
nor U5889 (N_5889,N_4897,N_4803);
and U5890 (N_5890,N_4797,N_4359);
or U5891 (N_5891,N_4286,N_4787);
or U5892 (N_5892,N_4322,N_4348);
or U5893 (N_5893,N_4384,N_4163);
nor U5894 (N_5894,N_4271,N_4574);
nand U5895 (N_5895,N_4909,N_4110);
xor U5896 (N_5896,N_4551,N_4819);
xnor U5897 (N_5897,N_4338,N_4360);
or U5898 (N_5898,N_4187,N_4766);
nor U5899 (N_5899,N_4900,N_4993);
nand U5900 (N_5900,N_4608,N_4363);
or U5901 (N_5901,N_4917,N_4184);
xnor U5902 (N_5902,N_4141,N_4582);
xor U5903 (N_5903,N_4014,N_4117);
nand U5904 (N_5904,N_4765,N_4520);
xor U5905 (N_5905,N_4630,N_4813);
or U5906 (N_5906,N_4448,N_4766);
and U5907 (N_5907,N_4029,N_4607);
xnor U5908 (N_5908,N_4068,N_4567);
nor U5909 (N_5909,N_4497,N_4300);
or U5910 (N_5910,N_4909,N_4686);
or U5911 (N_5911,N_4754,N_4369);
nor U5912 (N_5912,N_4593,N_4048);
nand U5913 (N_5913,N_4568,N_4694);
nand U5914 (N_5914,N_4450,N_4753);
and U5915 (N_5915,N_4616,N_4566);
xnor U5916 (N_5916,N_4798,N_4996);
nand U5917 (N_5917,N_4269,N_4599);
nor U5918 (N_5918,N_4662,N_4514);
and U5919 (N_5919,N_4177,N_4737);
or U5920 (N_5920,N_4609,N_4159);
nand U5921 (N_5921,N_4869,N_4034);
xor U5922 (N_5922,N_4736,N_4718);
nand U5923 (N_5923,N_4001,N_4729);
nand U5924 (N_5924,N_4273,N_4153);
xor U5925 (N_5925,N_4923,N_4492);
nand U5926 (N_5926,N_4001,N_4314);
nand U5927 (N_5927,N_4926,N_4051);
nand U5928 (N_5928,N_4893,N_4826);
and U5929 (N_5929,N_4792,N_4660);
nor U5930 (N_5930,N_4060,N_4538);
and U5931 (N_5931,N_4924,N_4161);
xnor U5932 (N_5932,N_4370,N_4539);
nor U5933 (N_5933,N_4324,N_4960);
nand U5934 (N_5934,N_4097,N_4556);
and U5935 (N_5935,N_4839,N_4706);
nor U5936 (N_5936,N_4539,N_4399);
or U5937 (N_5937,N_4866,N_4471);
and U5938 (N_5938,N_4620,N_4586);
or U5939 (N_5939,N_4300,N_4422);
xnor U5940 (N_5940,N_4201,N_4067);
nor U5941 (N_5941,N_4023,N_4937);
nor U5942 (N_5942,N_4444,N_4419);
and U5943 (N_5943,N_4697,N_4986);
xnor U5944 (N_5944,N_4536,N_4274);
nor U5945 (N_5945,N_4861,N_4634);
xnor U5946 (N_5946,N_4409,N_4655);
xor U5947 (N_5947,N_4489,N_4564);
nor U5948 (N_5948,N_4574,N_4971);
and U5949 (N_5949,N_4584,N_4172);
and U5950 (N_5950,N_4842,N_4904);
or U5951 (N_5951,N_4541,N_4582);
nand U5952 (N_5952,N_4570,N_4815);
nor U5953 (N_5953,N_4662,N_4353);
and U5954 (N_5954,N_4781,N_4732);
nand U5955 (N_5955,N_4583,N_4601);
xor U5956 (N_5956,N_4771,N_4663);
nand U5957 (N_5957,N_4659,N_4390);
and U5958 (N_5958,N_4156,N_4888);
or U5959 (N_5959,N_4215,N_4783);
nand U5960 (N_5960,N_4136,N_4001);
xor U5961 (N_5961,N_4407,N_4822);
or U5962 (N_5962,N_4930,N_4297);
nor U5963 (N_5963,N_4167,N_4396);
nand U5964 (N_5964,N_4336,N_4956);
and U5965 (N_5965,N_4287,N_4281);
nor U5966 (N_5966,N_4225,N_4223);
or U5967 (N_5967,N_4719,N_4960);
nand U5968 (N_5968,N_4432,N_4444);
xor U5969 (N_5969,N_4778,N_4916);
or U5970 (N_5970,N_4942,N_4738);
and U5971 (N_5971,N_4563,N_4614);
xor U5972 (N_5972,N_4526,N_4930);
or U5973 (N_5973,N_4795,N_4381);
or U5974 (N_5974,N_4848,N_4187);
xnor U5975 (N_5975,N_4505,N_4623);
nand U5976 (N_5976,N_4158,N_4800);
and U5977 (N_5977,N_4478,N_4915);
xnor U5978 (N_5978,N_4150,N_4426);
xnor U5979 (N_5979,N_4700,N_4280);
nand U5980 (N_5980,N_4328,N_4578);
and U5981 (N_5981,N_4452,N_4617);
or U5982 (N_5982,N_4037,N_4805);
xor U5983 (N_5983,N_4221,N_4467);
nor U5984 (N_5984,N_4356,N_4876);
and U5985 (N_5985,N_4484,N_4728);
nand U5986 (N_5986,N_4486,N_4811);
and U5987 (N_5987,N_4422,N_4354);
xor U5988 (N_5988,N_4827,N_4200);
and U5989 (N_5989,N_4208,N_4249);
nand U5990 (N_5990,N_4536,N_4164);
xor U5991 (N_5991,N_4218,N_4083);
nor U5992 (N_5992,N_4069,N_4699);
and U5993 (N_5993,N_4023,N_4466);
or U5994 (N_5994,N_4967,N_4170);
or U5995 (N_5995,N_4069,N_4065);
nor U5996 (N_5996,N_4175,N_4121);
nor U5997 (N_5997,N_4966,N_4642);
nor U5998 (N_5998,N_4677,N_4586);
xor U5999 (N_5999,N_4628,N_4779);
nand U6000 (N_6000,N_5722,N_5848);
nor U6001 (N_6001,N_5914,N_5207);
nor U6002 (N_6002,N_5127,N_5922);
xnor U6003 (N_6003,N_5405,N_5155);
xnor U6004 (N_6004,N_5775,N_5825);
xnor U6005 (N_6005,N_5138,N_5813);
xnor U6006 (N_6006,N_5968,N_5894);
nand U6007 (N_6007,N_5644,N_5165);
nand U6008 (N_6008,N_5771,N_5421);
or U6009 (N_6009,N_5497,N_5224);
and U6010 (N_6010,N_5923,N_5759);
nand U6011 (N_6011,N_5426,N_5607);
nand U6012 (N_6012,N_5301,N_5599);
xnor U6013 (N_6013,N_5340,N_5755);
nor U6014 (N_6014,N_5799,N_5208);
or U6015 (N_6015,N_5663,N_5269);
or U6016 (N_6016,N_5436,N_5437);
or U6017 (N_6017,N_5697,N_5615);
or U6018 (N_6018,N_5820,N_5560);
and U6019 (N_6019,N_5788,N_5311);
and U6020 (N_6020,N_5559,N_5126);
xor U6021 (N_6021,N_5933,N_5478);
xor U6022 (N_6022,N_5756,N_5837);
xnor U6023 (N_6023,N_5416,N_5846);
or U6024 (N_6024,N_5080,N_5428);
and U6025 (N_6025,N_5708,N_5355);
nand U6026 (N_6026,N_5844,N_5243);
xor U6027 (N_6027,N_5612,N_5907);
xnor U6028 (N_6028,N_5040,N_5206);
or U6029 (N_6029,N_5971,N_5794);
xnor U6030 (N_6030,N_5537,N_5779);
xnor U6031 (N_6031,N_5806,N_5839);
xnor U6032 (N_6032,N_5459,N_5177);
nand U6033 (N_6033,N_5056,N_5001);
or U6034 (N_6034,N_5252,N_5186);
nand U6035 (N_6035,N_5577,N_5280);
xor U6036 (N_6036,N_5498,N_5992);
or U6037 (N_6037,N_5329,N_5656);
and U6038 (N_6038,N_5858,N_5276);
or U6039 (N_6039,N_5845,N_5620);
nor U6040 (N_6040,N_5944,N_5228);
and U6041 (N_6041,N_5400,N_5103);
nand U6042 (N_6042,N_5627,N_5489);
xnor U6043 (N_6043,N_5580,N_5823);
nand U6044 (N_6044,N_5624,N_5380);
xnor U6045 (N_6045,N_5928,N_5109);
nor U6046 (N_6046,N_5122,N_5991);
nand U6047 (N_6047,N_5125,N_5084);
xor U6048 (N_6048,N_5729,N_5955);
nor U6049 (N_6049,N_5027,N_5689);
or U6050 (N_6050,N_5540,N_5981);
or U6051 (N_6051,N_5524,N_5867);
and U6052 (N_6052,N_5891,N_5601);
nand U6053 (N_6053,N_5427,N_5157);
nor U6054 (N_6054,N_5574,N_5768);
and U6055 (N_6055,N_5895,N_5623);
nand U6056 (N_6056,N_5838,N_5645);
or U6057 (N_6057,N_5211,N_5541);
and U6058 (N_6058,N_5073,N_5116);
and U6059 (N_6059,N_5639,N_5287);
nand U6060 (N_6060,N_5758,N_5547);
xnor U6061 (N_6061,N_5055,N_5636);
xor U6062 (N_6062,N_5546,N_5835);
xnor U6063 (N_6063,N_5592,N_5007);
nand U6064 (N_6064,N_5019,N_5821);
and U6065 (N_6065,N_5316,N_5500);
nor U6066 (N_6066,N_5651,N_5936);
and U6067 (N_6067,N_5064,N_5807);
nand U6068 (N_6068,N_5602,N_5174);
and U6069 (N_6069,N_5849,N_5595);
and U6070 (N_6070,N_5888,N_5246);
nand U6071 (N_6071,N_5951,N_5370);
or U6072 (N_6072,N_5480,N_5088);
and U6073 (N_6073,N_5101,N_5544);
nor U6074 (N_6074,N_5764,N_5302);
and U6075 (N_6075,N_5474,N_5015);
nor U6076 (N_6076,N_5626,N_5596);
and U6077 (N_6077,N_5250,N_5876);
or U6078 (N_6078,N_5781,N_5131);
and U6079 (N_6079,N_5572,N_5665);
or U6080 (N_6080,N_5034,N_5536);
or U6081 (N_6081,N_5377,N_5969);
and U6082 (N_6082,N_5702,N_5908);
nor U6083 (N_6083,N_5790,N_5447);
or U6084 (N_6084,N_5096,N_5810);
nand U6085 (N_6085,N_5715,N_5909);
nand U6086 (N_6086,N_5318,N_5526);
or U6087 (N_6087,N_5430,N_5168);
xnor U6088 (N_6088,N_5898,N_5331);
xnor U6089 (N_6089,N_5660,N_5934);
nor U6090 (N_6090,N_5222,N_5255);
xor U6091 (N_6091,N_5952,N_5718);
xnor U6092 (N_6092,N_5957,N_5930);
nor U6093 (N_6093,N_5076,N_5905);
nand U6094 (N_6094,N_5324,N_5328);
nor U6095 (N_6095,N_5213,N_5522);
xor U6096 (N_6096,N_5904,N_5139);
nor U6097 (N_6097,N_5836,N_5210);
nor U6098 (N_6098,N_5110,N_5819);
and U6099 (N_6099,N_5528,N_5648);
nor U6100 (N_6100,N_5227,N_5391);
xnor U6101 (N_6101,N_5997,N_5966);
or U6102 (N_6102,N_5036,N_5225);
or U6103 (N_6103,N_5273,N_5798);
nor U6104 (N_6104,N_5583,N_5690);
nor U6105 (N_6105,N_5477,N_5071);
nand U6106 (N_6106,N_5214,N_5803);
xor U6107 (N_6107,N_5760,N_5284);
or U6108 (N_6108,N_5107,N_5467);
xnor U6109 (N_6109,N_5070,N_5632);
and U6110 (N_6110,N_5203,N_5286);
and U6111 (N_6111,N_5913,N_5613);
nand U6112 (N_6112,N_5319,N_5411);
nor U6113 (N_6113,N_5711,N_5024);
nand U6114 (N_6114,N_5156,N_5986);
xor U6115 (N_6115,N_5159,N_5667);
nand U6116 (N_6116,N_5066,N_5145);
xor U6117 (N_6117,N_5927,N_5698);
and U6118 (N_6118,N_5237,N_5153);
nor U6119 (N_6119,N_5098,N_5197);
or U6120 (N_6120,N_5988,N_5148);
or U6121 (N_6121,N_5093,N_5023);
or U6122 (N_6122,N_5360,N_5638);
or U6123 (N_6123,N_5121,N_5358);
and U6124 (N_6124,N_5916,N_5552);
or U6125 (N_6125,N_5832,N_5670);
nand U6126 (N_6126,N_5533,N_5095);
and U6127 (N_6127,N_5452,N_5005);
or U6128 (N_6128,N_5622,N_5531);
or U6129 (N_6129,N_5608,N_5162);
and U6130 (N_6130,N_5030,N_5339);
xnor U6131 (N_6131,N_5183,N_5661);
nand U6132 (N_6132,N_5432,N_5499);
nor U6133 (N_6133,N_5047,N_5990);
or U6134 (N_6134,N_5647,N_5422);
or U6135 (N_6135,N_5146,N_5899);
xnor U6136 (N_6136,N_5633,N_5052);
and U6137 (N_6137,N_5889,N_5600);
xnor U6138 (N_6138,N_5947,N_5641);
nor U6139 (N_6139,N_5397,N_5332);
and U6140 (N_6140,N_5965,N_5744);
nand U6141 (N_6141,N_5508,N_5884);
xor U6142 (N_6142,N_5124,N_5353);
nand U6143 (N_6143,N_5576,N_5494);
or U6144 (N_6144,N_5388,N_5506);
nor U6145 (N_6145,N_5719,N_5309);
nor U6146 (N_6146,N_5415,N_5188);
or U6147 (N_6147,N_5575,N_5772);
xor U6148 (N_6148,N_5535,N_5193);
nand U6149 (N_6149,N_5958,N_5363);
xnor U6150 (N_6150,N_5181,N_5960);
or U6151 (N_6151,N_5291,N_5014);
nor U6152 (N_6152,N_5762,N_5584);
and U6153 (N_6153,N_5439,N_5882);
nand U6154 (N_6154,N_5926,N_5650);
or U6155 (N_6155,N_5337,N_5588);
and U6156 (N_6156,N_5264,N_5619);
and U6157 (N_6157,N_5382,N_5598);
nand U6158 (N_6158,N_5298,N_5616);
nand U6159 (N_6159,N_5903,N_5266);
or U6160 (N_6160,N_5707,N_5470);
nor U6161 (N_6161,N_5860,N_5017);
xor U6162 (N_6162,N_5473,N_5814);
xnor U6163 (N_6163,N_5020,N_5362);
or U6164 (N_6164,N_5743,N_5730);
xnor U6165 (N_6165,N_5841,N_5677);
nor U6166 (N_6166,N_5581,N_5099);
nor U6167 (N_6167,N_5343,N_5379);
and U6168 (N_6168,N_5140,N_5396);
xnor U6169 (N_6169,N_5878,N_5414);
nand U6170 (N_6170,N_5950,N_5048);
nand U6171 (N_6171,N_5874,N_5075);
nor U6172 (N_6172,N_5578,N_5100);
xnor U6173 (N_6173,N_5006,N_5694);
xnor U6174 (N_6174,N_5802,N_5850);
nor U6175 (N_6175,N_5948,N_5369);
nand U6176 (N_6176,N_5142,N_5022);
and U6177 (N_6177,N_5275,N_5381);
nand U6178 (N_6178,N_5031,N_5129);
or U6179 (N_6179,N_5539,N_5325);
nor U6180 (N_6180,N_5853,N_5373);
and U6181 (N_6181,N_5978,N_5094);
and U6182 (N_6182,N_5683,N_5886);
nor U6183 (N_6183,N_5199,N_5606);
or U6184 (N_6184,N_5890,N_5834);
and U6185 (N_6185,N_5617,N_5726);
nand U6186 (N_6186,N_5424,N_5628);
nor U6187 (N_6187,N_5290,N_5939);
nor U6188 (N_6188,N_5793,N_5270);
and U6189 (N_6189,N_5238,N_5198);
xnor U6190 (N_6190,N_5441,N_5582);
and U6191 (N_6191,N_5163,N_5425);
xnor U6192 (N_6192,N_5488,N_5289);
nor U6193 (N_6193,N_5984,N_5236);
or U6194 (N_6194,N_5371,N_5631);
xor U6195 (N_6195,N_5881,N_5995);
nor U6196 (N_6196,N_5682,N_5517);
and U6197 (N_6197,N_5384,N_5032);
nand U6198 (N_6198,N_5215,N_5590);
or U6199 (N_6199,N_5941,N_5789);
or U6200 (N_6200,N_5242,N_5239);
and U6201 (N_6201,N_5471,N_5061);
xnor U6202 (N_6202,N_5999,N_5566);
nor U6203 (N_6203,N_5194,N_5390);
xor U6204 (N_6204,N_5209,N_5774);
xor U6205 (N_6205,N_5658,N_5151);
xnor U6206 (N_6206,N_5979,N_5953);
xor U6207 (N_6207,N_5681,N_5089);
nor U6208 (N_6208,N_5253,N_5120);
and U6209 (N_6209,N_5993,N_5462);
nor U6210 (N_6210,N_5410,N_5366);
nand U6211 (N_6211,N_5413,N_5136);
and U6212 (N_6212,N_5134,N_5357);
nor U6213 (N_6213,N_5254,N_5761);
or U6214 (N_6214,N_5178,N_5733);
or U6215 (N_6215,N_5684,N_5365);
nand U6216 (N_6216,N_5833,N_5545);
xnor U6217 (N_6217,N_5260,N_5490);
and U6218 (N_6218,N_5696,N_5161);
xor U6219 (N_6219,N_5423,N_5050);
or U6220 (N_6220,N_5664,N_5679);
xnor U6221 (N_6221,N_5495,N_5265);
or U6222 (N_6222,N_5593,N_5012);
nand U6223 (N_6223,N_5847,N_5586);
nor U6224 (N_6224,N_5464,N_5067);
nand U6225 (N_6225,N_5221,N_5879);
xor U6226 (N_6226,N_5330,N_5784);
and U6227 (N_6227,N_5857,N_5629);
nand U6228 (N_6228,N_5507,N_5297);
nand U6229 (N_6229,N_5486,N_5223);
xnor U6230 (N_6230,N_5515,N_5118);
xor U6231 (N_6231,N_5108,N_5081);
and U6232 (N_6232,N_5387,N_5457);
nor U6233 (N_6233,N_5282,N_5351);
xnor U6234 (N_6234,N_5935,N_5117);
or U6235 (N_6235,N_5097,N_5468);
or U6236 (N_6236,N_5205,N_5863);
or U6237 (N_6237,N_5640,N_5083);
or U6238 (N_6238,N_5505,N_5346);
or U6239 (N_6239,N_5637,N_5766);
or U6240 (N_6240,N_5322,N_5344);
and U6241 (N_6241,N_5465,N_5585);
and U6242 (N_6242,N_5668,N_5959);
nor U6243 (N_6243,N_5361,N_5705);
and U6244 (N_6244,N_5736,N_5402);
and U6245 (N_6245,N_5688,N_5554);
and U6246 (N_6246,N_5672,N_5292);
xor U6247 (N_6247,N_5232,N_5043);
xnor U6248 (N_6248,N_5175,N_5141);
or U6249 (N_6249,N_5069,N_5757);
nand U6250 (N_6250,N_5809,N_5695);
nand U6251 (N_6251,N_5469,N_5954);
nand U6252 (N_6252,N_5356,N_5856);
and U6253 (N_6253,N_5873,N_5158);
xor U6254 (N_6254,N_5634,N_5128);
nor U6255 (N_6255,N_5815,N_5202);
or U6256 (N_6256,N_5114,N_5160);
and U6257 (N_6257,N_5312,N_5182);
xor U6258 (N_6258,N_5249,N_5666);
nand U6259 (N_6259,N_5748,N_5618);
and U6260 (N_6260,N_5354,N_5399);
or U6261 (N_6261,N_5407,N_5776);
nand U6262 (N_6262,N_5314,N_5072);
nand U6263 (N_6263,N_5609,N_5087);
and U6264 (N_6264,N_5143,N_5485);
or U6265 (N_6265,N_5008,N_5782);
xnor U6266 (N_6266,N_5614,N_5750);
or U6267 (N_6267,N_5455,N_5333);
nand U6268 (N_6268,N_5173,N_5395);
and U6269 (N_6269,N_5044,N_5751);
xnor U6270 (N_6270,N_5149,N_5513);
nand U6271 (N_6271,N_5869,N_5970);
nand U6272 (N_6272,N_5822,N_5787);
or U6273 (N_6273,N_5179,N_5920);
or U6274 (N_6274,N_5394,N_5795);
nand U6275 (N_6275,N_5398,N_5530);
xor U6276 (N_6276,N_5058,N_5763);
xor U6277 (N_6277,N_5680,N_5918);
nor U6278 (N_6278,N_5435,N_5041);
or U6279 (N_6279,N_5229,N_5741);
nand U6280 (N_6280,N_5037,N_5724);
nor U6281 (N_6281,N_5453,N_5323);
nor U6282 (N_6282,N_5212,N_5851);
nor U6283 (N_6283,N_5937,N_5204);
nor U6284 (N_6284,N_5800,N_5998);
and U6285 (N_6285,N_5520,N_5137);
nor U6286 (N_6286,N_5277,N_5737);
nand U6287 (N_6287,N_5630,N_5230);
and U6288 (N_6288,N_5152,N_5233);
nand U6289 (N_6289,N_5987,N_5674);
or U6290 (N_6290,N_5932,N_5011);
nor U6291 (N_6291,N_5299,N_5321);
xor U6292 (N_6292,N_5712,N_5885);
nand U6293 (N_6293,N_5862,N_5678);
and U6294 (N_6294,N_5703,N_5259);
and U6295 (N_6295,N_5603,N_5549);
nand U6296 (N_6296,N_5409,N_5510);
or U6297 (N_6297,N_5456,N_5112);
nor U6298 (N_6298,N_5817,N_5150);
xnor U6299 (N_6299,N_5035,N_5113);
xor U6300 (N_6300,N_5967,N_5565);
nand U6301 (N_6301,N_5655,N_5383);
nand U6302 (N_6302,N_5818,N_5315);
xnor U6303 (N_6303,N_5563,N_5735);
nand U6304 (N_6304,N_5686,N_5523);
and U6305 (N_6305,N_5285,N_5912);
xor U6306 (N_6306,N_5555,N_5078);
nand U6307 (N_6307,N_5172,N_5676);
xor U6308 (N_6308,N_5514,N_5240);
and U6309 (N_6309,N_5982,N_5504);
xnor U6310 (N_6310,N_5942,N_5102);
and U6311 (N_6311,N_5349,N_5740);
nor U6312 (N_6312,N_5662,N_5304);
or U6313 (N_6313,N_5412,N_5293);
nor U6314 (N_6314,N_5170,N_5294);
or U6315 (N_6315,N_5693,N_5875);
xnor U6316 (N_6316,N_5446,N_5880);
xor U6317 (N_6317,N_5653,N_5063);
and U6318 (N_6318,N_5231,N_5192);
xor U6319 (N_6319,N_5773,N_5278);
nand U6320 (N_6320,N_5454,N_5444);
or U6321 (N_6321,N_5057,N_5701);
xnor U6322 (N_6322,N_5003,N_5753);
nand U6323 (N_6323,N_5115,N_5691);
and U6324 (N_6324,N_5654,N_5458);
nand U6325 (N_6325,N_5466,N_5189);
and U6326 (N_6326,N_5217,N_5538);
xor U6327 (N_6327,N_5961,N_5828);
or U6328 (N_6328,N_5267,N_5562);
nand U6329 (N_6329,N_5945,N_5419);
nand U6330 (N_6330,N_5765,N_5642);
nand U6331 (N_6331,N_5943,N_5408);
nand U6332 (N_6332,N_5000,N_5348);
xnor U6333 (N_6333,N_5604,N_5949);
nor U6334 (N_6334,N_5086,N_5461);
nor U6335 (N_6335,N_5625,N_5829);
nor U6336 (N_6336,N_5429,N_5451);
and U6337 (N_6337,N_5090,N_5046);
and U6338 (N_6338,N_5201,N_5579);
nor U6339 (N_6339,N_5487,N_5983);
nor U6340 (N_6340,N_5975,N_5434);
nor U6341 (N_6341,N_5016,N_5725);
xor U6342 (N_6342,N_5797,N_5235);
nand U6343 (N_6343,N_5974,N_5564);
xnor U6344 (N_6344,N_5010,N_5785);
xor U6345 (N_6345,N_5443,N_5714);
nor U6346 (N_6346,N_5347,N_5310);
xnor U6347 (N_6347,N_5296,N_5283);
or U6348 (N_6348,N_5169,N_5376);
or U6349 (N_6349,N_5897,N_5611);
nor U6350 (N_6350,N_5184,N_5901);
or U6351 (N_6351,N_5732,N_5144);
nand U6352 (N_6352,N_5327,N_5512);
nor U6353 (N_6353,N_5502,N_5338);
nand U6354 (N_6354,N_5720,N_5385);
or U6355 (N_6355,N_5483,N_5556);
nand U6356 (N_6356,N_5335,N_5418);
and U6357 (N_6357,N_5171,N_5597);
nor U6358 (N_6358,N_5994,N_5062);
nand U6359 (N_6359,N_5859,N_5657);
or U6360 (N_6360,N_5571,N_5386);
and U6361 (N_6361,N_5364,N_5792);
xor U6362 (N_6362,N_5717,N_5262);
nor U6363 (N_6363,N_5247,N_5866);
xor U6364 (N_6364,N_5706,N_5709);
or U6365 (N_6365,N_5111,N_5865);
nor U6366 (N_6366,N_5472,N_5187);
nand U6367 (N_6367,N_5996,N_5527);
nand U6368 (N_6368,N_5028,N_5045);
or U6369 (N_6369,N_5244,N_5728);
and U6370 (N_6370,N_5352,N_5021);
or U6371 (N_6371,N_5378,N_5742);
or U6372 (N_6372,N_5166,N_5033);
and U6373 (N_6373,N_5257,N_5830);
nor U6374 (N_6374,N_5985,N_5009);
nor U6375 (N_6375,N_5754,N_5059);
xnor U6376 (N_6376,N_5481,N_5479);
xor U6377 (N_6377,N_5068,N_5106);
xor U6378 (N_6378,N_5811,N_5827);
nor U6379 (N_6379,N_5924,N_5196);
xor U6380 (N_6380,N_5448,N_5569);
and U6381 (N_6381,N_5673,N_5389);
or U6382 (N_6382,N_5700,N_5445);
and U6383 (N_6383,N_5896,N_5219);
or U6384 (N_6384,N_5946,N_5216);
or U6385 (N_6385,N_5104,N_5018);
nand U6386 (N_6386,N_5973,N_5812);
nor U6387 (N_6387,N_5687,N_5659);
xnor U6388 (N_6388,N_5525,N_5917);
xnor U6389 (N_6389,N_5542,N_5704);
nor U6390 (N_6390,N_5092,N_5482);
nand U6391 (N_6391,N_5393,N_5404);
and U6392 (N_6392,N_5721,N_5870);
or U6393 (N_6393,N_5039,N_5902);
xnor U6394 (N_6394,N_5646,N_5440);
or U6395 (N_6395,N_5652,N_5516);
xnor U6396 (N_6396,N_5085,N_5940);
nand U6397 (N_6397,N_5558,N_5263);
nor U6398 (N_6398,N_5038,N_5727);
or U6399 (N_6399,N_5375,N_5861);
and U6400 (N_6400,N_5509,N_5307);
and U6401 (N_6401,N_5854,N_5872);
and U6402 (N_6402,N_5132,N_5496);
and U6403 (N_6403,N_5042,N_5518);
xor U6404 (N_6404,N_5906,N_5868);
xnor U6405 (N_6405,N_5900,N_5133);
and U6406 (N_6406,N_5801,N_5739);
nand U6407 (N_6407,N_5501,N_5268);
nand U6408 (N_6408,N_5077,N_5449);
or U6409 (N_6409,N_5791,N_5082);
nor U6410 (N_6410,N_5406,N_5271);
xor U6411 (N_6411,N_5519,N_5079);
nand U6412 (N_6412,N_5476,N_5783);
and U6413 (N_6413,N_5029,N_5147);
and U6414 (N_6414,N_5403,N_5723);
nor U6415 (N_6415,N_5374,N_5699);
nand U6416 (N_6416,N_5342,N_5503);
nor U6417 (N_6417,N_5915,N_5534);
or U6418 (N_6418,N_5484,N_5359);
or U6419 (N_6419,N_5635,N_5931);
and U6420 (N_6420,N_5326,N_5288);
xor U6421 (N_6421,N_5685,N_5220);
or U6422 (N_6422,N_5060,N_5752);
nor U6423 (N_6423,N_5747,N_5191);
xnor U6424 (N_6424,N_5303,N_5734);
nand U6425 (N_6425,N_5910,N_5731);
xnor U6426 (N_6426,N_5401,N_5855);
xor U6427 (N_6427,N_5218,N_5295);
nand U6428 (N_6428,N_5300,N_5074);
xnor U6429 (N_6429,N_5272,N_5568);
nand U6430 (N_6430,N_5883,N_5164);
xnor U6431 (N_6431,N_5180,N_5808);
or U6432 (N_6432,N_5274,N_5893);
nor U6433 (N_6433,N_5130,N_5929);
or U6434 (N_6434,N_5919,N_5119);
nor U6435 (N_6435,N_5543,N_5433);
xnor U6436 (N_6436,N_5521,N_5567);
and U6437 (N_6437,N_5013,N_5313);
nor U6438 (N_6438,N_5831,N_5258);
nor U6439 (N_6439,N_5345,N_5176);
and U6440 (N_6440,N_5805,N_5649);
or U6441 (N_6441,N_5643,N_5675);
nor U6442 (N_6442,N_5123,N_5532);
nand U6443 (N_6443,N_5621,N_5049);
and U6444 (N_6444,N_5840,N_5550);
xnor U6445 (N_6445,N_5956,N_5463);
xor U6446 (N_6446,N_5925,N_5442);
xnor U6447 (N_6447,N_5251,N_5892);
and U6448 (N_6448,N_5368,N_5460);
and U6449 (N_6449,N_5420,N_5417);
nand U6450 (N_6450,N_5025,N_5769);
or U6451 (N_6451,N_5551,N_5594);
nor U6452 (N_6452,N_5589,N_5852);
xnor U6453 (N_6453,N_5716,N_5051);
nor U6454 (N_6454,N_5713,N_5778);
xnor U6455 (N_6455,N_5305,N_5105);
or U6456 (N_6456,N_5054,N_5864);
xnor U6457 (N_6457,N_5306,N_5317);
nor U6458 (N_6458,N_5548,N_5241);
or U6459 (N_6459,N_5281,N_5135);
or U6460 (N_6460,N_5963,N_5770);
nor U6461 (N_6461,N_5976,N_5261);
and U6462 (N_6462,N_5749,N_5557);
xor U6463 (N_6463,N_5561,N_5392);
xnor U6464 (N_6464,N_5786,N_5279);
xnor U6465 (N_6465,N_5877,N_5671);
xor U6466 (N_6466,N_5320,N_5053);
or U6467 (N_6467,N_5843,N_5921);
or U6468 (N_6468,N_5185,N_5245);
nor U6469 (N_6469,N_5767,N_5553);
xor U6470 (N_6470,N_5710,N_5570);
nand U6471 (N_6471,N_5738,N_5796);
or U6472 (N_6472,N_5964,N_5573);
and U6473 (N_6473,N_5911,N_5511);
nand U6474 (N_6474,N_5154,N_5610);
and U6475 (N_6475,N_5587,N_5989);
xor U6476 (N_6476,N_5491,N_5334);
nor U6477 (N_6477,N_5367,N_5826);
xor U6478 (N_6478,N_5824,N_5004);
nor U6479 (N_6479,N_5002,N_5248);
nor U6480 (N_6480,N_5605,N_5529);
xor U6481 (N_6481,N_5887,N_5372);
and U6482 (N_6482,N_5256,N_5065);
or U6483 (N_6483,N_5200,N_5350);
xnor U6484 (N_6484,N_5842,N_5804);
or U6485 (N_6485,N_5190,N_5591);
nand U6486 (N_6486,N_5167,N_5438);
xnor U6487 (N_6487,N_5692,N_5980);
and U6488 (N_6488,N_5871,N_5816);
and U6489 (N_6489,N_5493,N_5195);
xor U6490 (N_6490,N_5234,N_5091);
or U6491 (N_6491,N_5492,N_5336);
xnor U6492 (N_6492,N_5938,N_5431);
and U6493 (N_6493,N_5026,N_5341);
nor U6494 (N_6494,N_5962,N_5977);
and U6495 (N_6495,N_5450,N_5475);
nand U6496 (N_6496,N_5777,N_5308);
nand U6497 (N_6497,N_5669,N_5745);
and U6498 (N_6498,N_5972,N_5226);
xnor U6499 (N_6499,N_5780,N_5746);
or U6500 (N_6500,N_5548,N_5796);
and U6501 (N_6501,N_5967,N_5316);
and U6502 (N_6502,N_5720,N_5895);
nor U6503 (N_6503,N_5738,N_5750);
or U6504 (N_6504,N_5522,N_5455);
xnor U6505 (N_6505,N_5903,N_5125);
nor U6506 (N_6506,N_5089,N_5050);
nand U6507 (N_6507,N_5637,N_5997);
nand U6508 (N_6508,N_5727,N_5544);
and U6509 (N_6509,N_5956,N_5434);
nor U6510 (N_6510,N_5327,N_5996);
nand U6511 (N_6511,N_5562,N_5531);
nor U6512 (N_6512,N_5109,N_5572);
nand U6513 (N_6513,N_5209,N_5267);
and U6514 (N_6514,N_5325,N_5677);
xor U6515 (N_6515,N_5057,N_5085);
and U6516 (N_6516,N_5640,N_5535);
or U6517 (N_6517,N_5656,N_5568);
nor U6518 (N_6518,N_5376,N_5613);
xnor U6519 (N_6519,N_5512,N_5202);
nand U6520 (N_6520,N_5072,N_5601);
xor U6521 (N_6521,N_5505,N_5385);
or U6522 (N_6522,N_5707,N_5050);
and U6523 (N_6523,N_5370,N_5111);
xnor U6524 (N_6524,N_5581,N_5997);
xnor U6525 (N_6525,N_5385,N_5253);
nor U6526 (N_6526,N_5708,N_5195);
nand U6527 (N_6527,N_5262,N_5070);
nor U6528 (N_6528,N_5400,N_5014);
xnor U6529 (N_6529,N_5326,N_5650);
nand U6530 (N_6530,N_5714,N_5133);
or U6531 (N_6531,N_5974,N_5627);
and U6532 (N_6532,N_5532,N_5131);
nand U6533 (N_6533,N_5778,N_5285);
and U6534 (N_6534,N_5081,N_5284);
nor U6535 (N_6535,N_5238,N_5639);
nor U6536 (N_6536,N_5307,N_5342);
or U6537 (N_6537,N_5168,N_5964);
nor U6538 (N_6538,N_5923,N_5177);
nand U6539 (N_6539,N_5003,N_5805);
xnor U6540 (N_6540,N_5153,N_5992);
xnor U6541 (N_6541,N_5789,N_5049);
nor U6542 (N_6542,N_5226,N_5675);
xnor U6543 (N_6543,N_5366,N_5963);
nand U6544 (N_6544,N_5713,N_5620);
and U6545 (N_6545,N_5893,N_5815);
and U6546 (N_6546,N_5442,N_5730);
nor U6547 (N_6547,N_5638,N_5406);
or U6548 (N_6548,N_5219,N_5357);
nor U6549 (N_6549,N_5503,N_5080);
nor U6550 (N_6550,N_5841,N_5691);
nand U6551 (N_6551,N_5557,N_5110);
or U6552 (N_6552,N_5503,N_5070);
and U6553 (N_6553,N_5344,N_5535);
or U6554 (N_6554,N_5625,N_5060);
and U6555 (N_6555,N_5089,N_5030);
or U6556 (N_6556,N_5485,N_5711);
and U6557 (N_6557,N_5707,N_5030);
xor U6558 (N_6558,N_5019,N_5483);
or U6559 (N_6559,N_5747,N_5468);
xnor U6560 (N_6560,N_5458,N_5456);
xnor U6561 (N_6561,N_5991,N_5587);
nand U6562 (N_6562,N_5723,N_5429);
xor U6563 (N_6563,N_5195,N_5449);
xor U6564 (N_6564,N_5612,N_5974);
and U6565 (N_6565,N_5697,N_5112);
nor U6566 (N_6566,N_5987,N_5582);
nand U6567 (N_6567,N_5652,N_5848);
nand U6568 (N_6568,N_5816,N_5686);
or U6569 (N_6569,N_5630,N_5993);
or U6570 (N_6570,N_5404,N_5667);
and U6571 (N_6571,N_5974,N_5639);
xor U6572 (N_6572,N_5828,N_5902);
nor U6573 (N_6573,N_5456,N_5765);
nand U6574 (N_6574,N_5688,N_5908);
and U6575 (N_6575,N_5637,N_5869);
and U6576 (N_6576,N_5278,N_5470);
nand U6577 (N_6577,N_5703,N_5163);
or U6578 (N_6578,N_5773,N_5706);
or U6579 (N_6579,N_5071,N_5957);
or U6580 (N_6580,N_5669,N_5302);
and U6581 (N_6581,N_5628,N_5820);
nand U6582 (N_6582,N_5128,N_5150);
xnor U6583 (N_6583,N_5382,N_5789);
or U6584 (N_6584,N_5561,N_5379);
or U6585 (N_6585,N_5685,N_5356);
nor U6586 (N_6586,N_5871,N_5334);
nor U6587 (N_6587,N_5797,N_5957);
or U6588 (N_6588,N_5084,N_5424);
nor U6589 (N_6589,N_5939,N_5687);
nand U6590 (N_6590,N_5144,N_5107);
or U6591 (N_6591,N_5327,N_5490);
nor U6592 (N_6592,N_5225,N_5243);
xnor U6593 (N_6593,N_5524,N_5597);
xnor U6594 (N_6594,N_5227,N_5696);
and U6595 (N_6595,N_5942,N_5933);
xor U6596 (N_6596,N_5150,N_5218);
nor U6597 (N_6597,N_5819,N_5474);
or U6598 (N_6598,N_5890,N_5325);
and U6599 (N_6599,N_5541,N_5218);
nand U6600 (N_6600,N_5298,N_5542);
nor U6601 (N_6601,N_5027,N_5343);
and U6602 (N_6602,N_5036,N_5527);
and U6603 (N_6603,N_5019,N_5947);
nor U6604 (N_6604,N_5670,N_5312);
nor U6605 (N_6605,N_5558,N_5642);
or U6606 (N_6606,N_5400,N_5888);
nand U6607 (N_6607,N_5942,N_5486);
xor U6608 (N_6608,N_5099,N_5775);
nor U6609 (N_6609,N_5235,N_5157);
nand U6610 (N_6610,N_5905,N_5661);
xnor U6611 (N_6611,N_5817,N_5321);
xor U6612 (N_6612,N_5674,N_5428);
xor U6613 (N_6613,N_5962,N_5052);
and U6614 (N_6614,N_5257,N_5487);
xor U6615 (N_6615,N_5177,N_5891);
nand U6616 (N_6616,N_5470,N_5703);
nor U6617 (N_6617,N_5331,N_5270);
xnor U6618 (N_6618,N_5414,N_5913);
or U6619 (N_6619,N_5345,N_5340);
or U6620 (N_6620,N_5658,N_5017);
nand U6621 (N_6621,N_5695,N_5394);
and U6622 (N_6622,N_5411,N_5799);
and U6623 (N_6623,N_5331,N_5035);
and U6624 (N_6624,N_5458,N_5550);
or U6625 (N_6625,N_5877,N_5095);
xnor U6626 (N_6626,N_5004,N_5230);
nor U6627 (N_6627,N_5785,N_5977);
xnor U6628 (N_6628,N_5566,N_5693);
nor U6629 (N_6629,N_5409,N_5149);
xnor U6630 (N_6630,N_5239,N_5197);
or U6631 (N_6631,N_5704,N_5628);
or U6632 (N_6632,N_5674,N_5222);
nor U6633 (N_6633,N_5128,N_5159);
xnor U6634 (N_6634,N_5927,N_5040);
or U6635 (N_6635,N_5284,N_5899);
or U6636 (N_6636,N_5845,N_5520);
or U6637 (N_6637,N_5472,N_5774);
and U6638 (N_6638,N_5822,N_5849);
or U6639 (N_6639,N_5602,N_5438);
nand U6640 (N_6640,N_5365,N_5375);
nor U6641 (N_6641,N_5094,N_5861);
xnor U6642 (N_6642,N_5316,N_5359);
xor U6643 (N_6643,N_5326,N_5195);
xnor U6644 (N_6644,N_5826,N_5829);
nand U6645 (N_6645,N_5329,N_5931);
and U6646 (N_6646,N_5640,N_5356);
or U6647 (N_6647,N_5659,N_5144);
nand U6648 (N_6648,N_5055,N_5831);
nor U6649 (N_6649,N_5042,N_5498);
xnor U6650 (N_6650,N_5350,N_5571);
xnor U6651 (N_6651,N_5550,N_5160);
nand U6652 (N_6652,N_5621,N_5042);
nand U6653 (N_6653,N_5256,N_5850);
and U6654 (N_6654,N_5181,N_5729);
nand U6655 (N_6655,N_5264,N_5924);
nor U6656 (N_6656,N_5589,N_5462);
or U6657 (N_6657,N_5252,N_5719);
and U6658 (N_6658,N_5676,N_5035);
nand U6659 (N_6659,N_5363,N_5075);
xor U6660 (N_6660,N_5687,N_5726);
xor U6661 (N_6661,N_5332,N_5743);
nand U6662 (N_6662,N_5372,N_5030);
nor U6663 (N_6663,N_5250,N_5804);
or U6664 (N_6664,N_5577,N_5766);
nand U6665 (N_6665,N_5593,N_5908);
xnor U6666 (N_6666,N_5970,N_5842);
nor U6667 (N_6667,N_5866,N_5181);
or U6668 (N_6668,N_5284,N_5419);
or U6669 (N_6669,N_5005,N_5711);
or U6670 (N_6670,N_5824,N_5780);
nor U6671 (N_6671,N_5085,N_5391);
nor U6672 (N_6672,N_5233,N_5160);
xnor U6673 (N_6673,N_5999,N_5251);
or U6674 (N_6674,N_5724,N_5983);
and U6675 (N_6675,N_5081,N_5598);
nor U6676 (N_6676,N_5305,N_5485);
xnor U6677 (N_6677,N_5425,N_5493);
nor U6678 (N_6678,N_5934,N_5312);
nor U6679 (N_6679,N_5203,N_5125);
nand U6680 (N_6680,N_5707,N_5849);
and U6681 (N_6681,N_5362,N_5927);
nor U6682 (N_6682,N_5954,N_5787);
nand U6683 (N_6683,N_5986,N_5407);
or U6684 (N_6684,N_5273,N_5754);
or U6685 (N_6685,N_5659,N_5566);
and U6686 (N_6686,N_5772,N_5621);
nand U6687 (N_6687,N_5752,N_5910);
and U6688 (N_6688,N_5206,N_5176);
xor U6689 (N_6689,N_5392,N_5274);
xor U6690 (N_6690,N_5431,N_5206);
xnor U6691 (N_6691,N_5458,N_5904);
nand U6692 (N_6692,N_5427,N_5501);
or U6693 (N_6693,N_5728,N_5036);
and U6694 (N_6694,N_5880,N_5304);
xor U6695 (N_6695,N_5157,N_5781);
nor U6696 (N_6696,N_5893,N_5054);
xnor U6697 (N_6697,N_5329,N_5977);
xor U6698 (N_6698,N_5768,N_5908);
nor U6699 (N_6699,N_5494,N_5248);
xnor U6700 (N_6700,N_5301,N_5154);
or U6701 (N_6701,N_5460,N_5345);
nand U6702 (N_6702,N_5915,N_5276);
or U6703 (N_6703,N_5331,N_5517);
or U6704 (N_6704,N_5516,N_5333);
nand U6705 (N_6705,N_5871,N_5596);
xor U6706 (N_6706,N_5240,N_5244);
nor U6707 (N_6707,N_5511,N_5524);
nand U6708 (N_6708,N_5201,N_5167);
nand U6709 (N_6709,N_5081,N_5347);
and U6710 (N_6710,N_5736,N_5181);
and U6711 (N_6711,N_5361,N_5401);
and U6712 (N_6712,N_5285,N_5152);
nor U6713 (N_6713,N_5691,N_5974);
or U6714 (N_6714,N_5154,N_5187);
and U6715 (N_6715,N_5332,N_5112);
or U6716 (N_6716,N_5754,N_5644);
nand U6717 (N_6717,N_5538,N_5750);
or U6718 (N_6718,N_5741,N_5107);
nor U6719 (N_6719,N_5948,N_5892);
nor U6720 (N_6720,N_5630,N_5090);
nand U6721 (N_6721,N_5763,N_5926);
and U6722 (N_6722,N_5578,N_5298);
nor U6723 (N_6723,N_5678,N_5864);
nand U6724 (N_6724,N_5916,N_5853);
or U6725 (N_6725,N_5227,N_5259);
xnor U6726 (N_6726,N_5226,N_5787);
nand U6727 (N_6727,N_5991,N_5117);
nor U6728 (N_6728,N_5259,N_5828);
nor U6729 (N_6729,N_5887,N_5463);
and U6730 (N_6730,N_5046,N_5887);
xnor U6731 (N_6731,N_5795,N_5495);
xnor U6732 (N_6732,N_5198,N_5152);
or U6733 (N_6733,N_5876,N_5999);
nand U6734 (N_6734,N_5948,N_5555);
or U6735 (N_6735,N_5123,N_5618);
xor U6736 (N_6736,N_5801,N_5142);
and U6737 (N_6737,N_5336,N_5298);
or U6738 (N_6738,N_5061,N_5221);
and U6739 (N_6739,N_5148,N_5138);
nor U6740 (N_6740,N_5361,N_5527);
nor U6741 (N_6741,N_5947,N_5228);
xnor U6742 (N_6742,N_5991,N_5777);
nand U6743 (N_6743,N_5333,N_5098);
xor U6744 (N_6744,N_5495,N_5990);
xor U6745 (N_6745,N_5565,N_5767);
nand U6746 (N_6746,N_5804,N_5019);
nor U6747 (N_6747,N_5455,N_5916);
nand U6748 (N_6748,N_5259,N_5283);
nand U6749 (N_6749,N_5998,N_5104);
nor U6750 (N_6750,N_5960,N_5802);
or U6751 (N_6751,N_5369,N_5556);
nor U6752 (N_6752,N_5752,N_5779);
xnor U6753 (N_6753,N_5486,N_5253);
or U6754 (N_6754,N_5117,N_5378);
xor U6755 (N_6755,N_5283,N_5919);
xnor U6756 (N_6756,N_5395,N_5330);
or U6757 (N_6757,N_5204,N_5479);
nand U6758 (N_6758,N_5087,N_5421);
xnor U6759 (N_6759,N_5163,N_5750);
or U6760 (N_6760,N_5020,N_5895);
and U6761 (N_6761,N_5671,N_5483);
nor U6762 (N_6762,N_5783,N_5750);
nand U6763 (N_6763,N_5695,N_5229);
nor U6764 (N_6764,N_5538,N_5617);
and U6765 (N_6765,N_5141,N_5417);
or U6766 (N_6766,N_5453,N_5040);
nor U6767 (N_6767,N_5029,N_5967);
nand U6768 (N_6768,N_5192,N_5560);
or U6769 (N_6769,N_5211,N_5151);
and U6770 (N_6770,N_5738,N_5252);
or U6771 (N_6771,N_5087,N_5173);
nor U6772 (N_6772,N_5879,N_5019);
nand U6773 (N_6773,N_5332,N_5886);
xor U6774 (N_6774,N_5905,N_5218);
nor U6775 (N_6775,N_5928,N_5356);
xnor U6776 (N_6776,N_5670,N_5039);
and U6777 (N_6777,N_5609,N_5450);
xor U6778 (N_6778,N_5807,N_5958);
xor U6779 (N_6779,N_5080,N_5722);
or U6780 (N_6780,N_5671,N_5770);
nand U6781 (N_6781,N_5259,N_5632);
or U6782 (N_6782,N_5029,N_5935);
or U6783 (N_6783,N_5023,N_5842);
xor U6784 (N_6784,N_5785,N_5604);
nor U6785 (N_6785,N_5981,N_5175);
and U6786 (N_6786,N_5579,N_5392);
nor U6787 (N_6787,N_5547,N_5609);
or U6788 (N_6788,N_5824,N_5751);
xnor U6789 (N_6789,N_5142,N_5466);
xor U6790 (N_6790,N_5020,N_5397);
nor U6791 (N_6791,N_5149,N_5046);
and U6792 (N_6792,N_5347,N_5970);
nor U6793 (N_6793,N_5250,N_5149);
nor U6794 (N_6794,N_5375,N_5592);
nand U6795 (N_6795,N_5108,N_5300);
and U6796 (N_6796,N_5262,N_5023);
xor U6797 (N_6797,N_5517,N_5084);
nand U6798 (N_6798,N_5717,N_5942);
nand U6799 (N_6799,N_5449,N_5792);
nor U6800 (N_6800,N_5324,N_5899);
or U6801 (N_6801,N_5179,N_5997);
xnor U6802 (N_6802,N_5707,N_5123);
or U6803 (N_6803,N_5969,N_5610);
xnor U6804 (N_6804,N_5104,N_5898);
nor U6805 (N_6805,N_5365,N_5322);
nand U6806 (N_6806,N_5874,N_5100);
nor U6807 (N_6807,N_5650,N_5444);
and U6808 (N_6808,N_5643,N_5738);
nand U6809 (N_6809,N_5181,N_5583);
or U6810 (N_6810,N_5911,N_5378);
and U6811 (N_6811,N_5885,N_5185);
xnor U6812 (N_6812,N_5268,N_5774);
and U6813 (N_6813,N_5004,N_5655);
nand U6814 (N_6814,N_5373,N_5671);
or U6815 (N_6815,N_5956,N_5654);
nor U6816 (N_6816,N_5005,N_5614);
nor U6817 (N_6817,N_5057,N_5453);
nor U6818 (N_6818,N_5399,N_5182);
nand U6819 (N_6819,N_5378,N_5819);
or U6820 (N_6820,N_5963,N_5506);
nand U6821 (N_6821,N_5346,N_5242);
and U6822 (N_6822,N_5323,N_5655);
and U6823 (N_6823,N_5246,N_5954);
xnor U6824 (N_6824,N_5478,N_5697);
nor U6825 (N_6825,N_5156,N_5852);
nand U6826 (N_6826,N_5301,N_5632);
or U6827 (N_6827,N_5633,N_5837);
nand U6828 (N_6828,N_5949,N_5413);
or U6829 (N_6829,N_5231,N_5492);
nor U6830 (N_6830,N_5748,N_5706);
and U6831 (N_6831,N_5173,N_5646);
nor U6832 (N_6832,N_5098,N_5040);
nor U6833 (N_6833,N_5414,N_5054);
nor U6834 (N_6834,N_5994,N_5880);
or U6835 (N_6835,N_5525,N_5933);
nand U6836 (N_6836,N_5722,N_5494);
and U6837 (N_6837,N_5480,N_5829);
or U6838 (N_6838,N_5016,N_5215);
xor U6839 (N_6839,N_5354,N_5705);
and U6840 (N_6840,N_5778,N_5506);
xor U6841 (N_6841,N_5802,N_5798);
nand U6842 (N_6842,N_5191,N_5402);
and U6843 (N_6843,N_5123,N_5142);
or U6844 (N_6844,N_5617,N_5404);
and U6845 (N_6845,N_5938,N_5342);
or U6846 (N_6846,N_5691,N_5527);
nor U6847 (N_6847,N_5933,N_5699);
and U6848 (N_6848,N_5879,N_5710);
nand U6849 (N_6849,N_5421,N_5135);
or U6850 (N_6850,N_5433,N_5835);
or U6851 (N_6851,N_5370,N_5441);
nor U6852 (N_6852,N_5749,N_5442);
xor U6853 (N_6853,N_5993,N_5112);
xnor U6854 (N_6854,N_5740,N_5818);
nor U6855 (N_6855,N_5296,N_5098);
and U6856 (N_6856,N_5869,N_5460);
and U6857 (N_6857,N_5607,N_5898);
or U6858 (N_6858,N_5097,N_5231);
nand U6859 (N_6859,N_5635,N_5623);
or U6860 (N_6860,N_5183,N_5997);
nand U6861 (N_6861,N_5874,N_5359);
nor U6862 (N_6862,N_5766,N_5476);
nand U6863 (N_6863,N_5826,N_5883);
xor U6864 (N_6864,N_5144,N_5400);
xor U6865 (N_6865,N_5970,N_5515);
nand U6866 (N_6866,N_5478,N_5435);
xor U6867 (N_6867,N_5487,N_5191);
nor U6868 (N_6868,N_5206,N_5367);
nand U6869 (N_6869,N_5822,N_5586);
nand U6870 (N_6870,N_5537,N_5190);
nand U6871 (N_6871,N_5302,N_5122);
xor U6872 (N_6872,N_5109,N_5885);
or U6873 (N_6873,N_5000,N_5055);
and U6874 (N_6874,N_5855,N_5085);
nor U6875 (N_6875,N_5711,N_5742);
or U6876 (N_6876,N_5500,N_5013);
xnor U6877 (N_6877,N_5816,N_5807);
nand U6878 (N_6878,N_5020,N_5548);
xor U6879 (N_6879,N_5780,N_5898);
and U6880 (N_6880,N_5038,N_5188);
nand U6881 (N_6881,N_5025,N_5164);
xor U6882 (N_6882,N_5410,N_5276);
and U6883 (N_6883,N_5421,N_5544);
xor U6884 (N_6884,N_5689,N_5224);
nor U6885 (N_6885,N_5875,N_5609);
nor U6886 (N_6886,N_5984,N_5814);
and U6887 (N_6887,N_5549,N_5936);
or U6888 (N_6888,N_5214,N_5776);
or U6889 (N_6889,N_5940,N_5111);
xor U6890 (N_6890,N_5477,N_5878);
or U6891 (N_6891,N_5700,N_5393);
xor U6892 (N_6892,N_5027,N_5464);
nand U6893 (N_6893,N_5683,N_5184);
and U6894 (N_6894,N_5826,N_5571);
nor U6895 (N_6895,N_5777,N_5114);
or U6896 (N_6896,N_5037,N_5277);
or U6897 (N_6897,N_5704,N_5792);
or U6898 (N_6898,N_5934,N_5991);
and U6899 (N_6899,N_5045,N_5621);
xor U6900 (N_6900,N_5926,N_5641);
nor U6901 (N_6901,N_5567,N_5997);
nor U6902 (N_6902,N_5224,N_5650);
or U6903 (N_6903,N_5586,N_5560);
xnor U6904 (N_6904,N_5066,N_5272);
nor U6905 (N_6905,N_5402,N_5888);
nor U6906 (N_6906,N_5177,N_5562);
nand U6907 (N_6907,N_5293,N_5208);
nor U6908 (N_6908,N_5210,N_5751);
xor U6909 (N_6909,N_5951,N_5948);
nor U6910 (N_6910,N_5105,N_5820);
nor U6911 (N_6911,N_5362,N_5538);
or U6912 (N_6912,N_5773,N_5665);
nor U6913 (N_6913,N_5297,N_5677);
and U6914 (N_6914,N_5190,N_5484);
nand U6915 (N_6915,N_5358,N_5021);
and U6916 (N_6916,N_5659,N_5028);
xor U6917 (N_6917,N_5140,N_5676);
nor U6918 (N_6918,N_5269,N_5571);
nor U6919 (N_6919,N_5978,N_5118);
and U6920 (N_6920,N_5408,N_5947);
or U6921 (N_6921,N_5890,N_5166);
or U6922 (N_6922,N_5710,N_5491);
or U6923 (N_6923,N_5282,N_5206);
nand U6924 (N_6924,N_5308,N_5340);
and U6925 (N_6925,N_5683,N_5066);
xor U6926 (N_6926,N_5032,N_5215);
or U6927 (N_6927,N_5208,N_5071);
or U6928 (N_6928,N_5049,N_5828);
nand U6929 (N_6929,N_5677,N_5077);
xnor U6930 (N_6930,N_5443,N_5033);
nor U6931 (N_6931,N_5096,N_5988);
nor U6932 (N_6932,N_5524,N_5386);
nor U6933 (N_6933,N_5017,N_5780);
or U6934 (N_6934,N_5002,N_5588);
or U6935 (N_6935,N_5599,N_5071);
nand U6936 (N_6936,N_5526,N_5097);
nand U6937 (N_6937,N_5106,N_5517);
nor U6938 (N_6938,N_5970,N_5657);
xnor U6939 (N_6939,N_5559,N_5046);
nor U6940 (N_6940,N_5856,N_5713);
nand U6941 (N_6941,N_5372,N_5195);
nor U6942 (N_6942,N_5673,N_5921);
and U6943 (N_6943,N_5607,N_5045);
xnor U6944 (N_6944,N_5097,N_5170);
nand U6945 (N_6945,N_5256,N_5848);
and U6946 (N_6946,N_5581,N_5235);
or U6947 (N_6947,N_5558,N_5559);
or U6948 (N_6948,N_5107,N_5000);
nor U6949 (N_6949,N_5137,N_5585);
or U6950 (N_6950,N_5498,N_5884);
xnor U6951 (N_6951,N_5642,N_5059);
nand U6952 (N_6952,N_5568,N_5054);
xnor U6953 (N_6953,N_5220,N_5471);
xnor U6954 (N_6954,N_5887,N_5326);
nor U6955 (N_6955,N_5653,N_5596);
xor U6956 (N_6956,N_5392,N_5440);
nor U6957 (N_6957,N_5781,N_5431);
nand U6958 (N_6958,N_5942,N_5144);
nand U6959 (N_6959,N_5922,N_5949);
or U6960 (N_6960,N_5973,N_5131);
xnor U6961 (N_6961,N_5419,N_5250);
nor U6962 (N_6962,N_5499,N_5513);
nand U6963 (N_6963,N_5377,N_5994);
nand U6964 (N_6964,N_5462,N_5846);
nor U6965 (N_6965,N_5410,N_5194);
and U6966 (N_6966,N_5598,N_5208);
xor U6967 (N_6967,N_5872,N_5702);
and U6968 (N_6968,N_5505,N_5943);
and U6969 (N_6969,N_5969,N_5835);
xor U6970 (N_6970,N_5844,N_5275);
nand U6971 (N_6971,N_5002,N_5761);
nand U6972 (N_6972,N_5626,N_5561);
nand U6973 (N_6973,N_5627,N_5593);
and U6974 (N_6974,N_5772,N_5499);
nand U6975 (N_6975,N_5773,N_5694);
or U6976 (N_6976,N_5935,N_5610);
and U6977 (N_6977,N_5505,N_5904);
nand U6978 (N_6978,N_5634,N_5305);
or U6979 (N_6979,N_5542,N_5478);
xor U6980 (N_6980,N_5253,N_5440);
xnor U6981 (N_6981,N_5171,N_5617);
nor U6982 (N_6982,N_5426,N_5553);
or U6983 (N_6983,N_5064,N_5748);
xor U6984 (N_6984,N_5630,N_5057);
xor U6985 (N_6985,N_5405,N_5566);
and U6986 (N_6986,N_5599,N_5159);
xor U6987 (N_6987,N_5657,N_5190);
xnor U6988 (N_6988,N_5004,N_5224);
nand U6989 (N_6989,N_5305,N_5223);
and U6990 (N_6990,N_5594,N_5236);
nor U6991 (N_6991,N_5746,N_5117);
or U6992 (N_6992,N_5761,N_5641);
xor U6993 (N_6993,N_5701,N_5980);
and U6994 (N_6994,N_5474,N_5051);
and U6995 (N_6995,N_5642,N_5053);
nor U6996 (N_6996,N_5433,N_5679);
and U6997 (N_6997,N_5330,N_5685);
and U6998 (N_6998,N_5734,N_5331);
and U6999 (N_6999,N_5897,N_5766);
nand U7000 (N_7000,N_6283,N_6698);
or U7001 (N_7001,N_6008,N_6503);
nand U7002 (N_7002,N_6384,N_6299);
and U7003 (N_7003,N_6089,N_6724);
and U7004 (N_7004,N_6173,N_6940);
or U7005 (N_7005,N_6301,N_6810);
nor U7006 (N_7006,N_6360,N_6543);
and U7007 (N_7007,N_6766,N_6273);
nor U7008 (N_7008,N_6793,N_6842);
nand U7009 (N_7009,N_6968,N_6800);
or U7010 (N_7010,N_6477,N_6460);
nand U7011 (N_7011,N_6179,N_6974);
and U7012 (N_7012,N_6499,N_6757);
nand U7013 (N_7013,N_6669,N_6535);
xor U7014 (N_7014,N_6635,N_6030);
and U7015 (N_7015,N_6654,N_6402);
and U7016 (N_7016,N_6216,N_6506);
xnor U7017 (N_7017,N_6466,N_6470);
or U7018 (N_7018,N_6518,N_6650);
nor U7019 (N_7019,N_6243,N_6648);
nor U7020 (N_7020,N_6309,N_6451);
xnor U7021 (N_7021,N_6849,N_6742);
or U7022 (N_7022,N_6364,N_6036);
nand U7023 (N_7023,N_6469,N_6715);
and U7024 (N_7024,N_6716,N_6314);
or U7025 (N_7025,N_6446,N_6576);
xnor U7026 (N_7026,N_6428,N_6124);
xor U7027 (N_7027,N_6943,N_6893);
xor U7028 (N_7028,N_6408,N_6702);
nor U7029 (N_7029,N_6726,N_6075);
xor U7030 (N_7030,N_6671,N_6989);
and U7031 (N_7031,N_6288,N_6510);
or U7032 (N_7032,N_6372,N_6330);
or U7033 (N_7033,N_6111,N_6542);
xor U7034 (N_7034,N_6573,N_6382);
xnor U7035 (N_7035,N_6020,N_6000);
nor U7036 (N_7036,N_6951,N_6675);
nand U7037 (N_7037,N_6125,N_6975);
or U7038 (N_7038,N_6254,N_6291);
nand U7039 (N_7039,N_6444,N_6528);
or U7040 (N_7040,N_6206,N_6571);
nor U7041 (N_7041,N_6185,N_6165);
nand U7042 (N_7042,N_6655,N_6353);
xor U7043 (N_7043,N_6971,N_6607);
nor U7044 (N_7044,N_6608,N_6763);
xor U7045 (N_7045,N_6365,N_6997);
xnor U7046 (N_7046,N_6802,N_6797);
nand U7047 (N_7047,N_6632,N_6356);
nand U7048 (N_7048,N_6526,N_6533);
and U7049 (N_7049,N_6773,N_6912);
nor U7050 (N_7050,N_6452,N_6539);
and U7051 (N_7051,N_6728,N_6256);
and U7052 (N_7052,N_6690,N_6500);
or U7053 (N_7053,N_6917,N_6099);
xor U7054 (N_7054,N_6227,N_6144);
xnor U7055 (N_7055,N_6117,N_6455);
and U7056 (N_7056,N_6722,N_6848);
or U7057 (N_7057,N_6721,N_6198);
nor U7058 (N_7058,N_6113,N_6937);
nor U7059 (N_7059,N_6588,N_6122);
or U7060 (N_7060,N_6942,N_6473);
xor U7061 (N_7061,N_6718,N_6415);
or U7062 (N_7062,N_6764,N_6979);
nor U7063 (N_7063,N_6609,N_6816);
nand U7064 (N_7064,N_6884,N_6121);
and U7065 (N_7065,N_6935,N_6390);
nor U7066 (N_7066,N_6171,N_6739);
or U7067 (N_7067,N_6569,N_6164);
nor U7068 (N_7068,N_6960,N_6732);
or U7069 (N_7069,N_6063,N_6479);
nor U7070 (N_7070,N_6183,N_6964);
or U7071 (N_7071,N_6277,N_6925);
and U7072 (N_7072,N_6594,N_6775);
nor U7073 (N_7073,N_6443,N_6754);
or U7074 (N_7074,N_6765,N_6620);
and U7075 (N_7075,N_6044,N_6991);
nor U7076 (N_7076,N_6661,N_6647);
and U7077 (N_7077,N_6846,N_6965);
nor U7078 (N_7078,N_6705,N_6134);
xor U7079 (N_7079,N_6791,N_6694);
and U7080 (N_7080,N_6795,N_6474);
and U7081 (N_7081,N_6596,N_6229);
nand U7082 (N_7082,N_6221,N_6251);
nor U7083 (N_7083,N_6613,N_6205);
nor U7084 (N_7084,N_6271,N_6417);
xor U7085 (N_7085,N_6794,N_6264);
or U7086 (N_7086,N_6636,N_6047);
and U7087 (N_7087,N_6286,N_6200);
nand U7088 (N_7088,N_6045,N_6430);
and U7089 (N_7089,N_6901,N_6519);
nand U7090 (N_7090,N_6798,N_6274);
or U7091 (N_7091,N_6805,N_6593);
nand U7092 (N_7092,N_6651,N_6380);
xnor U7093 (N_7093,N_6984,N_6310);
or U7094 (N_7094,N_6666,N_6037);
nor U7095 (N_7095,N_6701,N_6293);
and U7096 (N_7096,N_6860,N_6048);
xnor U7097 (N_7097,N_6550,N_6263);
xnor U7098 (N_7098,N_6879,N_6736);
nor U7099 (N_7099,N_6103,N_6714);
nand U7100 (N_7100,N_6313,N_6850);
and U7101 (N_7101,N_6300,N_6143);
xnor U7102 (N_7102,N_6231,N_6489);
xor U7103 (N_7103,N_6447,N_6628);
or U7104 (N_7104,N_6371,N_6189);
xnor U7105 (N_7105,N_6803,N_6320);
xnor U7106 (N_7106,N_6821,N_6999);
nor U7107 (N_7107,N_6919,N_6983);
nand U7108 (N_7108,N_6396,N_6012);
nor U7109 (N_7109,N_6748,N_6230);
and U7110 (N_7110,N_6804,N_6723);
nor U7111 (N_7111,N_6426,N_6953);
and U7112 (N_7112,N_6076,N_6475);
and U7113 (N_7113,N_6969,N_6498);
nor U7114 (N_7114,N_6239,N_6049);
nor U7115 (N_7115,N_6545,N_6297);
xnor U7116 (N_7116,N_6188,N_6400);
or U7117 (N_7117,N_6411,N_6740);
xor U7118 (N_7118,N_6308,N_6375);
xnor U7119 (N_7119,N_6412,N_6696);
or U7120 (N_7120,N_6349,N_6427);
xnor U7121 (N_7121,N_6461,N_6042);
xor U7122 (N_7122,N_6900,N_6232);
and U7123 (N_7123,N_6249,N_6830);
and U7124 (N_7124,N_6602,N_6825);
or U7125 (N_7125,N_6978,N_6952);
or U7126 (N_7126,N_6495,N_6130);
nor U7127 (N_7127,N_6255,N_6357);
nor U7128 (N_7128,N_6483,N_6785);
nand U7129 (N_7129,N_6990,N_6224);
xor U7130 (N_7130,N_6343,N_6208);
and U7131 (N_7131,N_6015,N_6911);
nor U7132 (N_7132,N_6649,N_6304);
or U7133 (N_7133,N_6374,N_6465);
nand U7134 (N_7134,N_6448,N_6234);
and U7135 (N_7135,N_6839,N_6361);
nand U7136 (N_7136,N_6369,N_6982);
nor U7137 (N_7137,N_6598,N_6284);
xnor U7138 (N_7138,N_6688,N_6138);
xnor U7139 (N_7139,N_6325,N_6141);
or U7140 (N_7140,N_6634,N_6359);
nor U7141 (N_7141,N_6157,N_6644);
nor U7142 (N_7142,N_6406,N_6782);
xnor U7143 (N_7143,N_6084,N_6626);
nand U7144 (N_7144,N_6486,N_6679);
xor U7145 (N_7145,N_6615,N_6378);
nand U7146 (N_7146,N_6756,N_6098);
nand U7147 (N_7147,N_6868,N_6567);
nand U7148 (N_7148,N_6302,N_6881);
xor U7149 (N_7149,N_6921,N_6737);
nand U7150 (N_7150,N_6140,N_6938);
nand U7151 (N_7151,N_6522,N_6267);
nor U7152 (N_7152,N_6998,N_6811);
or U7153 (N_7153,N_6462,N_6203);
nand U7154 (N_7154,N_6551,N_6882);
nor U7155 (N_7155,N_6172,N_6060);
nor U7156 (N_7156,N_6876,N_6502);
and U7157 (N_7157,N_6069,N_6210);
xnor U7158 (N_7158,N_6908,N_6970);
xnor U7159 (N_7159,N_6516,N_6834);
nand U7160 (N_7160,N_6066,N_6664);
xor U7161 (N_7161,N_6070,N_6222);
nand U7162 (N_7162,N_6591,N_6156);
or U7163 (N_7163,N_6959,N_6269);
nand U7164 (N_7164,N_6823,N_6924);
nand U7165 (N_7165,N_6874,N_6676);
and U7166 (N_7166,N_6241,N_6425);
nand U7167 (N_7167,N_6092,N_6105);
or U7168 (N_7168,N_6133,N_6315);
or U7169 (N_7169,N_6824,N_6601);
nor U7170 (N_7170,N_6776,N_6324);
xnor U7171 (N_7171,N_6484,N_6788);
and U7172 (N_7172,N_6480,N_6719);
xnor U7173 (N_7173,N_6292,N_6897);
nand U7174 (N_7174,N_6871,N_6026);
or U7175 (N_7175,N_6238,N_6061);
and U7176 (N_7176,N_6948,N_6945);
or U7177 (N_7177,N_6319,N_6294);
xor U7178 (N_7178,N_6096,N_6665);
nand U7179 (N_7179,N_6864,N_6856);
xor U7180 (N_7180,N_6918,N_6219);
nor U7181 (N_7181,N_6672,N_6316);
or U7182 (N_7182,N_6629,N_6307);
nor U7183 (N_7183,N_6295,N_6738);
nor U7184 (N_7184,N_6563,N_6812);
nor U7185 (N_7185,N_6577,N_6837);
or U7186 (N_7186,N_6225,N_6611);
and U7187 (N_7187,N_6789,N_6858);
nand U7188 (N_7188,N_6685,N_6150);
xor U7189 (N_7189,N_6253,N_6114);
or U7190 (N_7190,N_6914,N_6091);
and U7191 (N_7191,N_6029,N_6581);
nand U7192 (N_7192,N_6708,N_6866);
xnor U7193 (N_7193,N_6014,N_6552);
nor U7194 (N_7194,N_6456,N_6927);
nand U7195 (N_7195,N_6407,N_6196);
nand U7196 (N_7196,N_6836,N_6278);
and U7197 (N_7197,N_6889,N_6471);
or U7198 (N_7198,N_6599,N_6128);
or U7199 (N_7199,N_6487,N_6910);
nand U7200 (N_7200,N_6025,N_6041);
nand U7201 (N_7201,N_6660,N_6323);
nand U7202 (N_7202,N_6115,N_6187);
nand U7203 (N_7203,N_6265,N_6281);
and U7204 (N_7204,N_6658,N_6605);
or U7205 (N_7205,N_6306,N_6760);
nand U7206 (N_7206,N_6769,N_6614);
xnor U7207 (N_7207,N_6815,N_6833);
nor U7208 (N_7208,N_6541,N_6734);
or U7209 (N_7209,N_6488,N_6051);
nand U7210 (N_7210,N_6363,N_6376);
nor U7211 (N_7211,N_6478,N_6963);
and U7212 (N_7212,N_6832,N_6340);
and U7213 (N_7213,N_6167,N_6184);
nand U7214 (N_7214,N_6529,N_6246);
nand U7215 (N_7215,N_6418,N_6016);
or U7216 (N_7216,N_6600,N_6215);
nand U7217 (N_7217,N_6907,N_6348);
or U7218 (N_7218,N_6368,N_6090);
nor U7219 (N_7219,N_6645,N_6829);
xor U7220 (N_7220,N_6019,N_6986);
nor U7221 (N_7221,N_6245,N_6414);
or U7222 (N_7222,N_6059,N_6341);
xnor U7223 (N_7223,N_6028,N_6904);
and U7224 (N_7224,N_6413,N_6178);
nor U7225 (N_7225,N_6903,N_6181);
and U7226 (N_7226,N_6958,N_6784);
and U7227 (N_7227,N_6244,N_6770);
nor U7228 (N_7228,N_6298,N_6562);
and U7229 (N_7229,N_6336,N_6064);
or U7230 (N_7230,N_6139,N_6102);
nor U7231 (N_7231,N_6485,N_6335);
nor U7232 (N_7232,N_6922,N_6709);
xor U7233 (N_7233,N_6553,N_6158);
nor U7234 (N_7234,N_6840,N_6713);
or U7235 (N_7235,N_6886,N_6381);
and U7236 (N_7236,N_6725,N_6339);
nand U7237 (N_7237,N_6112,N_6322);
or U7238 (N_7238,N_6689,N_6513);
and U7239 (N_7239,N_6056,N_6578);
nor U7240 (N_7240,N_6010,N_6711);
nor U7241 (N_7241,N_6104,N_6226);
and U7242 (N_7242,N_6887,N_6779);
and U7243 (N_7243,N_6746,N_6625);
xor U7244 (N_7244,N_6079,N_6652);
and U7245 (N_7245,N_6585,N_6345);
xor U7246 (N_7246,N_6610,N_6204);
nor U7247 (N_7247,N_6275,N_6508);
or U7248 (N_7248,N_6137,N_6890);
nor U7249 (N_7249,N_6633,N_6437);
nand U7250 (N_7250,N_6279,N_6442);
xor U7251 (N_7251,N_6399,N_6643);
and U7252 (N_7252,N_6538,N_6640);
and U7253 (N_7253,N_6768,N_6561);
nand U7254 (N_7254,N_6853,N_6367);
and U7255 (N_7255,N_6129,N_6898);
nor U7256 (N_7256,N_6317,N_6035);
and U7257 (N_7257,N_6252,N_6962);
nand U7258 (N_7258,N_6397,N_6373);
nand U7259 (N_7259,N_6646,N_6262);
and U7260 (N_7260,N_6052,N_6186);
and U7261 (N_7261,N_6395,N_6386);
nand U7262 (N_7262,N_6023,N_6257);
nor U7263 (N_7263,N_6459,N_6088);
nand U7264 (N_7264,N_6995,N_6132);
or U7265 (N_7265,N_6175,N_6828);
and U7266 (N_7266,N_6002,N_6354);
and U7267 (N_7267,N_6154,N_6806);
and U7268 (N_7268,N_6831,N_6944);
nand U7269 (N_7269,N_6272,N_6575);
or U7270 (N_7270,N_6383,N_6046);
xnor U7271 (N_7271,N_6153,N_6851);
xor U7272 (N_7272,N_6394,N_6807);
nand U7273 (N_7273,N_6501,N_6949);
or U7274 (N_7274,N_6270,N_6586);
or U7275 (N_7275,N_6440,N_6347);
and U7276 (N_7276,N_6107,N_6928);
and U7277 (N_7277,N_6201,N_6835);
or U7278 (N_7278,N_6468,N_6136);
nand U7279 (N_7279,N_6190,N_6845);
nand U7280 (N_7280,N_6967,N_6813);
and U7281 (N_7281,N_6355,N_6142);
or U7282 (N_7282,N_6033,N_6532);
or U7283 (N_7283,N_6767,N_6973);
and U7284 (N_7284,N_6078,N_6276);
xnor U7285 (N_7285,N_6631,N_6878);
xnor U7286 (N_7286,N_6476,N_6280);
xor U7287 (N_7287,N_6667,N_6496);
nand U7288 (N_7288,N_6521,N_6771);
nand U7289 (N_7289,N_6638,N_6071);
xor U7290 (N_7290,N_6393,N_6534);
xnor U7291 (N_7291,N_6867,N_6662);
xnor U7292 (N_7292,N_6050,N_6398);
nand U7293 (N_7293,N_6106,N_6604);
or U7294 (N_7294,N_6684,N_6560);
and U7295 (N_7295,N_6419,N_6548);
nand U7296 (N_7296,N_6009,N_6870);
nor U7297 (N_7297,N_6570,N_6405);
xor U7298 (N_7298,N_6031,N_6155);
nand U7299 (N_7299,N_6926,N_6544);
xnor U7300 (N_7300,N_6618,N_6482);
nor U7301 (N_7301,N_6131,N_6799);
or U7302 (N_7302,N_6761,N_6857);
xor U7303 (N_7303,N_6682,N_6450);
xnor U7304 (N_7304,N_6388,N_6344);
nor U7305 (N_7305,N_6093,N_6843);
nand U7306 (N_7306,N_6555,N_6656);
nor U7307 (N_7307,N_6915,N_6220);
or U7308 (N_7308,N_6527,N_6458);
nand U7309 (N_7309,N_6939,N_6584);
or U7310 (N_7310,N_6193,N_6233);
or U7311 (N_7311,N_6996,N_6670);
nor U7312 (N_7312,N_6163,N_6362);
nor U7313 (N_7313,N_6120,N_6118);
xor U7314 (N_7314,N_6085,N_6556);
or U7315 (N_7315,N_6192,N_6086);
nor U7316 (N_7316,N_6013,N_6159);
xor U7317 (N_7317,N_6449,N_6759);
and U7318 (N_7318,N_6438,N_6424);
nand U7319 (N_7319,N_6018,N_6540);
nor U7320 (N_7320,N_6454,N_6977);
xnor U7321 (N_7321,N_6587,N_6595);
nor U7322 (N_7322,N_6217,N_6745);
or U7323 (N_7323,N_6727,N_6720);
and U7324 (N_7324,N_6083,N_6494);
or U7325 (N_7325,N_6385,N_6236);
or U7326 (N_7326,N_6902,N_6622);
nand U7327 (N_7327,N_6781,N_6250);
nor U7328 (N_7328,N_6100,N_6289);
nor U7329 (N_7329,N_6027,N_6366);
nor U7330 (N_7330,N_6017,N_6683);
xnor U7331 (N_7331,N_6572,N_6957);
xnor U7332 (N_7332,N_6936,N_6021);
xor U7333 (N_7333,N_6703,N_6976);
or U7334 (N_7334,N_6235,N_6170);
nand U7335 (N_7335,N_6565,N_6180);
nor U7336 (N_7336,N_6616,N_6077);
nor U7337 (N_7337,N_6992,N_6214);
nor U7338 (N_7338,N_6744,N_6195);
or U7339 (N_7339,N_6073,N_6067);
xnor U7340 (N_7340,N_6961,N_6772);
and U7341 (N_7341,N_6337,N_6820);
or U7342 (N_7342,N_6743,N_6296);
xor U7343 (N_7343,N_6906,N_6282);
xnor U7344 (N_7344,N_6659,N_6603);
nand U7345 (N_7345,N_6753,N_6814);
xor U7346 (N_7346,N_6074,N_6116);
xnor U7347 (N_7347,N_6197,N_6237);
or U7348 (N_7348,N_6891,N_6929);
or U7349 (N_7349,N_6087,N_6681);
and U7350 (N_7350,N_6094,N_6801);
nor U7351 (N_7351,N_6699,N_6966);
and U7352 (N_7352,N_6880,N_6436);
nand U7353 (N_7353,N_6692,N_6826);
xnor U7354 (N_7354,N_6861,N_6980);
xor U7355 (N_7355,N_6700,N_6895);
nand U7356 (N_7356,N_6285,N_6326);
xor U7357 (N_7357,N_6751,N_6146);
nand U7358 (N_7358,N_6956,N_6733);
nor U7359 (N_7359,N_6057,N_6930);
or U7360 (N_7360,N_6492,N_6248);
or U7361 (N_7361,N_6580,N_6433);
and U7362 (N_7362,N_6321,N_6827);
or U7363 (N_7363,N_6592,N_6762);
xor U7364 (N_7364,N_6081,N_6920);
and U7365 (N_7365,N_6401,N_6512);
and U7366 (N_7366,N_6885,N_6673);
or U7367 (N_7367,N_6260,N_6520);
xor U7368 (N_7368,N_6370,N_6597);
and U7369 (N_7369,N_6043,N_6695);
or U7370 (N_7370,N_6985,N_6932);
nand U7371 (N_7371,N_6119,N_6329);
or U7372 (N_7372,N_6623,N_6182);
and U7373 (N_7373,N_6511,N_6574);
and U7374 (N_7374,N_6097,N_6844);
or U7375 (N_7375,N_6358,N_6993);
and U7376 (N_7376,N_6729,N_6712);
nor U7377 (N_7377,N_6505,N_6377);
and U7378 (N_7378,N_6007,N_6988);
xor U7379 (N_7379,N_6515,N_6677);
and U7380 (N_7380,N_6859,N_6663);
nand U7381 (N_7381,N_6391,N_6954);
nand U7382 (N_7382,N_6892,N_6972);
nand U7383 (N_7383,N_6177,N_6749);
xnor U7384 (N_7384,N_6004,N_6202);
or U7385 (N_7385,N_6687,N_6582);
nor U7386 (N_7386,N_6717,N_6457);
and U7387 (N_7387,N_6389,N_6525);
nand U7388 (N_7388,N_6082,N_6822);
or U7389 (N_7389,N_6410,N_6579);
or U7390 (N_7390,N_6223,N_6792);
or U7391 (N_7391,N_6531,N_6735);
or U7392 (N_7392,N_6854,N_6404);
and U7393 (N_7393,N_6431,N_6068);
and U7394 (N_7394,N_6127,N_6873);
nor U7395 (N_7395,N_6174,N_6493);
or U7396 (N_7396,N_6392,N_6053);
and U7397 (N_7397,N_6863,N_6946);
nor U7398 (N_7398,N_6564,N_6032);
nor U7399 (N_7399,N_6707,N_6786);
or U7400 (N_7400,N_6750,N_6022);
xnor U7401 (N_7401,N_6467,N_6504);
and U7402 (N_7402,N_6875,N_6606);
or U7403 (N_7403,N_6491,N_6916);
xor U7404 (N_7404,N_6808,N_6218);
xor U7405 (N_7405,N_6148,N_6865);
and U7406 (N_7406,N_6642,N_6240);
xor U7407 (N_7407,N_6536,N_6619);
or U7408 (N_7408,N_6191,N_6387);
nor U7409 (N_7409,N_6062,N_6706);
and U7410 (N_7410,N_6617,N_6338);
nor U7411 (N_7411,N_6472,N_6637);
xnor U7412 (N_7412,N_6123,N_6796);
nor U7413 (N_7413,N_6627,N_6778);
xnor U7414 (N_7414,N_6126,N_6869);
and U7415 (N_7415,N_6258,N_6730);
or U7416 (N_7416,N_6169,N_6855);
nand U7417 (N_7417,N_6108,N_6755);
nand U7418 (N_7418,N_6266,N_6168);
xnor U7419 (N_7419,N_6758,N_6416);
nor U7420 (N_7420,N_6896,N_6199);
and U7421 (N_7421,N_6710,N_6209);
nor U7422 (N_7422,N_6481,N_6441);
and U7423 (N_7423,N_6693,N_6639);
nand U7424 (N_7424,N_6403,N_6318);
nor U7425 (N_7425,N_6490,N_6328);
nor U7426 (N_7426,N_6691,N_6261);
xnor U7427 (N_7427,N_6497,N_6883);
nor U7428 (N_7428,N_6894,N_6247);
or U7429 (N_7429,N_6838,N_6242);
and U7430 (N_7430,N_6847,N_6621);
or U7431 (N_7431,N_6819,N_6590);
xnor U7432 (N_7432,N_6589,N_6290);
and U7433 (N_7433,N_6039,N_6537);
xnor U7434 (N_7434,N_6342,N_6211);
nand U7435 (N_7435,N_6818,N_6787);
or U7436 (N_7436,N_6657,N_6862);
nand U7437 (N_7437,N_6624,N_6809);
xor U7438 (N_7438,N_6212,N_6334);
or U7439 (N_7439,N_6704,N_6003);
and U7440 (N_7440,N_6303,N_6054);
or U7441 (N_7441,N_6162,N_6101);
nor U7442 (N_7442,N_6072,N_6034);
or U7443 (N_7443,N_6987,N_6147);
or U7444 (N_7444,N_6841,N_6024);
or U7445 (N_7445,N_6777,N_6305);
or U7446 (N_7446,N_6557,N_6523);
nand U7447 (N_7447,N_6011,N_6332);
nor U7448 (N_7448,N_6549,N_6287);
or U7449 (N_7449,N_6423,N_6686);
xnor U7450 (N_7450,N_6259,N_6674);
or U7451 (N_7451,N_6955,N_6877);
nand U7452 (N_7452,N_6311,N_6422);
or U7453 (N_7453,N_6038,N_6434);
or U7454 (N_7454,N_6546,N_6559);
or U7455 (N_7455,N_6934,N_6530);
nand U7456 (N_7456,N_6080,N_6566);
xor U7457 (N_7457,N_6161,N_6554);
or U7458 (N_7458,N_6680,N_6909);
nand U7459 (N_7459,N_6001,N_6933);
and U7460 (N_7460,N_6464,N_6435);
xor U7461 (N_7461,N_6509,N_6931);
and U7462 (N_7462,N_6409,N_6194);
or U7463 (N_7463,N_6006,N_6095);
nand U7464 (N_7464,N_6207,N_6852);
or U7465 (N_7465,N_6941,N_6145);
nor U7466 (N_7466,N_6568,N_6421);
nor U7467 (N_7467,N_6327,N_6783);
and U7468 (N_7468,N_6331,N_6547);
nand U7469 (N_7469,N_6913,N_6160);
or U7470 (N_7470,N_6517,N_6899);
nor U7471 (N_7471,N_6558,N_6947);
or U7472 (N_7472,N_6312,N_6507);
xnor U7473 (N_7473,N_6731,N_6872);
nand U7474 (N_7474,N_6774,N_6994);
xnor U7475 (N_7475,N_6346,N_6420);
or U7476 (N_7476,N_6453,N_6065);
xor U7477 (N_7477,N_6653,N_6524);
and U7478 (N_7478,N_6432,N_6630);
and U7479 (N_7479,N_6350,N_6352);
xor U7480 (N_7480,N_6697,N_6228);
and U7481 (N_7481,N_6005,N_6152);
and U7482 (N_7482,N_6166,N_6151);
nand U7483 (N_7483,N_6741,N_6439);
nor U7484 (N_7484,N_6678,N_6923);
nor U7485 (N_7485,N_6109,N_6110);
nor U7486 (N_7486,N_6888,N_6514);
nor U7487 (N_7487,N_6950,N_6463);
or U7488 (N_7488,N_6379,N_6817);
nand U7489 (N_7489,N_6445,N_6176);
nand U7490 (N_7490,N_6905,N_6790);
or U7491 (N_7491,N_6981,N_6429);
and U7492 (N_7492,N_6149,N_6058);
xor U7493 (N_7493,N_6668,N_6055);
nand U7494 (N_7494,N_6040,N_6213);
xor U7495 (N_7495,N_6641,N_6135);
nor U7496 (N_7496,N_6333,N_6752);
nand U7497 (N_7497,N_6583,N_6747);
nand U7498 (N_7498,N_6268,N_6612);
xnor U7499 (N_7499,N_6351,N_6780);
and U7500 (N_7500,N_6639,N_6744);
and U7501 (N_7501,N_6532,N_6007);
and U7502 (N_7502,N_6692,N_6944);
xor U7503 (N_7503,N_6809,N_6486);
nor U7504 (N_7504,N_6806,N_6521);
xnor U7505 (N_7505,N_6779,N_6906);
and U7506 (N_7506,N_6933,N_6794);
and U7507 (N_7507,N_6028,N_6989);
nand U7508 (N_7508,N_6573,N_6869);
or U7509 (N_7509,N_6451,N_6357);
or U7510 (N_7510,N_6681,N_6717);
nor U7511 (N_7511,N_6440,N_6647);
or U7512 (N_7512,N_6798,N_6478);
and U7513 (N_7513,N_6284,N_6462);
nor U7514 (N_7514,N_6487,N_6766);
or U7515 (N_7515,N_6250,N_6343);
xor U7516 (N_7516,N_6796,N_6780);
nand U7517 (N_7517,N_6576,N_6372);
and U7518 (N_7518,N_6629,N_6298);
or U7519 (N_7519,N_6391,N_6769);
nand U7520 (N_7520,N_6903,N_6760);
xnor U7521 (N_7521,N_6964,N_6902);
nor U7522 (N_7522,N_6967,N_6057);
nand U7523 (N_7523,N_6312,N_6882);
and U7524 (N_7524,N_6048,N_6794);
nor U7525 (N_7525,N_6072,N_6619);
nor U7526 (N_7526,N_6143,N_6409);
and U7527 (N_7527,N_6557,N_6129);
nor U7528 (N_7528,N_6852,N_6880);
or U7529 (N_7529,N_6503,N_6370);
and U7530 (N_7530,N_6254,N_6866);
nand U7531 (N_7531,N_6498,N_6388);
and U7532 (N_7532,N_6109,N_6690);
nand U7533 (N_7533,N_6651,N_6754);
or U7534 (N_7534,N_6147,N_6421);
xnor U7535 (N_7535,N_6175,N_6859);
and U7536 (N_7536,N_6015,N_6026);
xor U7537 (N_7537,N_6240,N_6589);
nand U7538 (N_7538,N_6323,N_6954);
and U7539 (N_7539,N_6931,N_6831);
nand U7540 (N_7540,N_6866,N_6343);
or U7541 (N_7541,N_6786,N_6421);
nand U7542 (N_7542,N_6935,N_6992);
xnor U7543 (N_7543,N_6258,N_6300);
xor U7544 (N_7544,N_6755,N_6589);
and U7545 (N_7545,N_6745,N_6766);
nand U7546 (N_7546,N_6290,N_6336);
and U7547 (N_7547,N_6366,N_6918);
xnor U7548 (N_7548,N_6980,N_6925);
xor U7549 (N_7549,N_6190,N_6194);
and U7550 (N_7550,N_6188,N_6602);
and U7551 (N_7551,N_6426,N_6338);
xor U7552 (N_7552,N_6076,N_6287);
nor U7553 (N_7553,N_6467,N_6919);
nor U7554 (N_7554,N_6257,N_6957);
or U7555 (N_7555,N_6313,N_6587);
xor U7556 (N_7556,N_6507,N_6472);
nand U7557 (N_7557,N_6433,N_6474);
or U7558 (N_7558,N_6317,N_6729);
xnor U7559 (N_7559,N_6048,N_6632);
and U7560 (N_7560,N_6359,N_6961);
xnor U7561 (N_7561,N_6889,N_6864);
or U7562 (N_7562,N_6706,N_6878);
nand U7563 (N_7563,N_6620,N_6002);
xor U7564 (N_7564,N_6842,N_6153);
xnor U7565 (N_7565,N_6358,N_6526);
or U7566 (N_7566,N_6965,N_6933);
or U7567 (N_7567,N_6480,N_6358);
nor U7568 (N_7568,N_6278,N_6337);
nand U7569 (N_7569,N_6432,N_6943);
and U7570 (N_7570,N_6666,N_6430);
nor U7571 (N_7571,N_6953,N_6313);
nand U7572 (N_7572,N_6883,N_6159);
or U7573 (N_7573,N_6430,N_6064);
nand U7574 (N_7574,N_6124,N_6950);
and U7575 (N_7575,N_6622,N_6772);
xor U7576 (N_7576,N_6877,N_6273);
or U7577 (N_7577,N_6425,N_6817);
xnor U7578 (N_7578,N_6300,N_6155);
and U7579 (N_7579,N_6689,N_6796);
nand U7580 (N_7580,N_6960,N_6757);
nor U7581 (N_7581,N_6779,N_6438);
and U7582 (N_7582,N_6811,N_6814);
and U7583 (N_7583,N_6247,N_6119);
nand U7584 (N_7584,N_6753,N_6841);
nor U7585 (N_7585,N_6734,N_6736);
xor U7586 (N_7586,N_6206,N_6297);
nand U7587 (N_7587,N_6909,N_6803);
nand U7588 (N_7588,N_6262,N_6459);
nand U7589 (N_7589,N_6299,N_6032);
and U7590 (N_7590,N_6171,N_6836);
nand U7591 (N_7591,N_6691,N_6779);
nand U7592 (N_7592,N_6107,N_6545);
nor U7593 (N_7593,N_6990,N_6750);
nor U7594 (N_7594,N_6653,N_6907);
and U7595 (N_7595,N_6924,N_6727);
nand U7596 (N_7596,N_6007,N_6260);
or U7597 (N_7597,N_6021,N_6697);
nor U7598 (N_7598,N_6770,N_6889);
xor U7599 (N_7599,N_6383,N_6096);
or U7600 (N_7600,N_6566,N_6267);
or U7601 (N_7601,N_6735,N_6852);
xnor U7602 (N_7602,N_6337,N_6417);
nand U7603 (N_7603,N_6270,N_6723);
xor U7604 (N_7604,N_6833,N_6455);
and U7605 (N_7605,N_6798,N_6460);
nor U7606 (N_7606,N_6217,N_6836);
and U7607 (N_7607,N_6561,N_6506);
xnor U7608 (N_7608,N_6277,N_6806);
and U7609 (N_7609,N_6174,N_6594);
and U7610 (N_7610,N_6192,N_6364);
and U7611 (N_7611,N_6401,N_6504);
or U7612 (N_7612,N_6895,N_6794);
xor U7613 (N_7613,N_6318,N_6118);
nor U7614 (N_7614,N_6407,N_6552);
nor U7615 (N_7615,N_6836,N_6058);
and U7616 (N_7616,N_6769,N_6365);
or U7617 (N_7617,N_6053,N_6950);
nor U7618 (N_7618,N_6524,N_6867);
or U7619 (N_7619,N_6247,N_6858);
or U7620 (N_7620,N_6953,N_6168);
nand U7621 (N_7621,N_6464,N_6231);
xor U7622 (N_7622,N_6490,N_6502);
and U7623 (N_7623,N_6412,N_6770);
and U7624 (N_7624,N_6226,N_6467);
xor U7625 (N_7625,N_6757,N_6273);
xnor U7626 (N_7626,N_6898,N_6097);
or U7627 (N_7627,N_6754,N_6001);
and U7628 (N_7628,N_6975,N_6250);
and U7629 (N_7629,N_6673,N_6464);
nand U7630 (N_7630,N_6714,N_6560);
xnor U7631 (N_7631,N_6287,N_6471);
nand U7632 (N_7632,N_6429,N_6971);
or U7633 (N_7633,N_6743,N_6233);
xor U7634 (N_7634,N_6545,N_6021);
nand U7635 (N_7635,N_6609,N_6017);
or U7636 (N_7636,N_6229,N_6801);
xor U7637 (N_7637,N_6489,N_6855);
or U7638 (N_7638,N_6088,N_6272);
or U7639 (N_7639,N_6666,N_6018);
xnor U7640 (N_7640,N_6103,N_6923);
nor U7641 (N_7641,N_6343,N_6729);
and U7642 (N_7642,N_6448,N_6239);
nor U7643 (N_7643,N_6930,N_6505);
xor U7644 (N_7644,N_6273,N_6911);
xor U7645 (N_7645,N_6225,N_6311);
or U7646 (N_7646,N_6554,N_6846);
or U7647 (N_7647,N_6266,N_6000);
xnor U7648 (N_7648,N_6645,N_6468);
nand U7649 (N_7649,N_6556,N_6996);
nand U7650 (N_7650,N_6058,N_6344);
xnor U7651 (N_7651,N_6761,N_6823);
nand U7652 (N_7652,N_6621,N_6216);
and U7653 (N_7653,N_6179,N_6216);
or U7654 (N_7654,N_6486,N_6709);
nor U7655 (N_7655,N_6246,N_6485);
xnor U7656 (N_7656,N_6353,N_6052);
and U7657 (N_7657,N_6154,N_6324);
nor U7658 (N_7658,N_6040,N_6657);
and U7659 (N_7659,N_6786,N_6929);
and U7660 (N_7660,N_6775,N_6178);
or U7661 (N_7661,N_6729,N_6184);
or U7662 (N_7662,N_6173,N_6670);
nor U7663 (N_7663,N_6095,N_6435);
nand U7664 (N_7664,N_6573,N_6797);
or U7665 (N_7665,N_6058,N_6946);
xor U7666 (N_7666,N_6383,N_6154);
xor U7667 (N_7667,N_6513,N_6982);
nor U7668 (N_7668,N_6992,N_6963);
or U7669 (N_7669,N_6079,N_6056);
nor U7670 (N_7670,N_6327,N_6886);
nor U7671 (N_7671,N_6276,N_6847);
nor U7672 (N_7672,N_6482,N_6275);
xnor U7673 (N_7673,N_6460,N_6099);
xnor U7674 (N_7674,N_6606,N_6509);
or U7675 (N_7675,N_6883,N_6083);
nand U7676 (N_7676,N_6784,N_6482);
and U7677 (N_7677,N_6303,N_6522);
nand U7678 (N_7678,N_6825,N_6282);
nor U7679 (N_7679,N_6075,N_6111);
or U7680 (N_7680,N_6030,N_6978);
or U7681 (N_7681,N_6595,N_6542);
nand U7682 (N_7682,N_6147,N_6873);
nor U7683 (N_7683,N_6745,N_6492);
nor U7684 (N_7684,N_6641,N_6025);
xor U7685 (N_7685,N_6455,N_6879);
nor U7686 (N_7686,N_6930,N_6034);
and U7687 (N_7687,N_6605,N_6678);
nor U7688 (N_7688,N_6673,N_6880);
xnor U7689 (N_7689,N_6856,N_6760);
nor U7690 (N_7690,N_6084,N_6807);
nand U7691 (N_7691,N_6030,N_6308);
xnor U7692 (N_7692,N_6124,N_6161);
nor U7693 (N_7693,N_6258,N_6118);
and U7694 (N_7694,N_6930,N_6368);
or U7695 (N_7695,N_6489,N_6420);
nand U7696 (N_7696,N_6932,N_6516);
nor U7697 (N_7697,N_6895,N_6550);
or U7698 (N_7698,N_6739,N_6152);
nor U7699 (N_7699,N_6355,N_6090);
nand U7700 (N_7700,N_6185,N_6607);
or U7701 (N_7701,N_6440,N_6335);
nor U7702 (N_7702,N_6716,N_6410);
xnor U7703 (N_7703,N_6106,N_6336);
or U7704 (N_7704,N_6383,N_6104);
nor U7705 (N_7705,N_6515,N_6015);
or U7706 (N_7706,N_6208,N_6624);
nand U7707 (N_7707,N_6114,N_6646);
and U7708 (N_7708,N_6077,N_6589);
or U7709 (N_7709,N_6527,N_6198);
nand U7710 (N_7710,N_6496,N_6243);
and U7711 (N_7711,N_6056,N_6256);
nand U7712 (N_7712,N_6758,N_6993);
nor U7713 (N_7713,N_6985,N_6223);
xnor U7714 (N_7714,N_6385,N_6066);
nor U7715 (N_7715,N_6387,N_6636);
nor U7716 (N_7716,N_6267,N_6968);
and U7717 (N_7717,N_6273,N_6753);
xor U7718 (N_7718,N_6946,N_6250);
and U7719 (N_7719,N_6154,N_6139);
nor U7720 (N_7720,N_6575,N_6311);
nand U7721 (N_7721,N_6883,N_6923);
xor U7722 (N_7722,N_6609,N_6978);
or U7723 (N_7723,N_6655,N_6879);
or U7724 (N_7724,N_6793,N_6811);
and U7725 (N_7725,N_6119,N_6665);
or U7726 (N_7726,N_6716,N_6051);
or U7727 (N_7727,N_6475,N_6546);
nor U7728 (N_7728,N_6330,N_6134);
nand U7729 (N_7729,N_6859,N_6766);
nor U7730 (N_7730,N_6687,N_6281);
xnor U7731 (N_7731,N_6364,N_6834);
xnor U7732 (N_7732,N_6526,N_6541);
nor U7733 (N_7733,N_6239,N_6087);
nor U7734 (N_7734,N_6037,N_6687);
nor U7735 (N_7735,N_6216,N_6841);
nor U7736 (N_7736,N_6548,N_6802);
and U7737 (N_7737,N_6875,N_6369);
nand U7738 (N_7738,N_6984,N_6682);
xnor U7739 (N_7739,N_6745,N_6261);
nand U7740 (N_7740,N_6635,N_6867);
nor U7741 (N_7741,N_6147,N_6258);
or U7742 (N_7742,N_6299,N_6937);
nand U7743 (N_7743,N_6550,N_6329);
and U7744 (N_7744,N_6431,N_6472);
or U7745 (N_7745,N_6101,N_6699);
nor U7746 (N_7746,N_6725,N_6848);
nand U7747 (N_7747,N_6855,N_6521);
nand U7748 (N_7748,N_6289,N_6269);
nor U7749 (N_7749,N_6622,N_6346);
xnor U7750 (N_7750,N_6793,N_6278);
xnor U7751 (N_7751,N_6651,N_6104);
xnor U7752 (N_7752,N_6468,N_6029);
and U7753 (N_7753,N_6587,N_6170);
nor U7754 (N_7754,N_6714,N_6543);
nor U7755 (N_7755,N_6722,N_6452);
and U7756 (N_7756,N_6324,N_6797);
xnor U7757 (N_7757,N_6130,N_6187);
nand U7758 (N_7758,N_6998,N_6813);
and U7759 (N_7759,N_6041,N_6099);
and U7760 (N_7760,N_6092,N_6637);
or U7761 (N_7761,N_6190,N_6883);
nand U7762 (N_7762,N_6398,N_6855);
or U7763 (N_7763,N_6095,N_6283);
nand U7764 (N_7764,N_6393,N_6090);
nand U7765 (N_7765,N_6083,N_6646);
and U7766 (N_7766,N_6752,N_6392);
xor U7767 (N_7767,N_6449,N_6580);
nand U7768 (N_7768,N_6290,N_6987);
xor U7769 (N_7769,N_6071,N_6848);
xnor U7770 (N_7770,N_6968,N_6616);
nand U7771 (N_7771,N_6372,N_6184);
nand U7772 (N_7772,N_6167,N_6025);
nor U7773 (N_7773,N_6092,N_6782);
nand U7774 (N_7774,N_6892,N_6831);
nand U7775 (N_7775,N_6881,N_6051);
nand U7776 (N_7776,N_6304,N_6425);
and U7777 (N_7777,N_6454,N_6593);
nor U7778 (N_7778,N_6035,N_6979);
or U7779 (N_7779,N_6865,N_6676);
or U7780 (N_7780,N_6966,N_6131);
nor U7781 (N_7781,N_6974,N_6457);
nor U7782 (N_7782,N_6583,N_6745);
nor U7783 (N_7783,N_6677,N_6765);
nor U7784 (N_7784,N_6449,N_6324);
nand U7785 (N_7785,N_6816,N_6253);
and U7786 (N_7786,N_6613,N_6444);
nand U7787 (N_7787,N_6038,N_6032);
nand U7788 (N_7788,N_6046,N_6971);
and U7789 (N_7789,N_6687,N_6489);
nor U7790 (N_7790,N_6810,N_6237);
or U7791 (N_7791,N_6188,N_6898);
nand U7792 (N_7792,N_6899,N_6572);
and U7793 (N_7793,N_6031,N_6801);
or U7794 (N_7794,N_6641,N_6346);
nand U7795 (N_7795,N_6590,N_6664);
xnor U7796 (N_7796,N_6391,N_6665);
and U7797 (N_7797,N_6909,N_6717);
nor U7798 (N_7798,N_6795,N_6300);
nand U7799 (N_7799,N_6486,N_6947);
and U7800 (N_7800,N_6463,N_6050);
nand U7801 (N_7801,N_6312,N_6182);
nand U7802 (N_7802,N_6771,N_6945);
nand U7803 (N_7803,N_6077,N_6624);
nor U7804 (N_7804,N_6612,N_6050);
xnor U7805 (N_7805,N_6139,N_6170);
or U7806 (N_7806,N_6476,N_6918);
nor U7807 (N_7807,N_6635,N_6015);
nand U7808 (N_7808,N_6843,N_6469);
xnor U7809 (N_7809,N_6692,N_6408);
nor U7810 (N_7810,N_6685,N_6199);
nand U7811 (N_7811,N_6689,N_6897);
xor U7812 (N_7812,N_6403,N_6914);
or U7813 (N_7813,N_6500,N_6998);
nand U7814 (N_7814,N_6833,N_6338);
nand U7815 (N_7815,N_6767,N_6286);
nand U7816 (N_7816,N_6801,N_6516);
xnor U7817 (N_7817,N_6469,N_6451);
nor U7818 (N_7818,N_6688,N_6900);
nand U7819 (N_7819,N_6532,N_6110);
nand U7820 (N_7820,N_6050,N_6274);
xor U7821 (N_7821,N_6632,N_6446);
nand U7822 (N_7822,N_6930,N_6017);
xnor U7823 (N_7823,N_6221,N_6597);
nor U7824 (N_7824,N_6322,N_6195);
nor U7825 (N_7825,N_6049,N_6158);
or U7826 (N_7826,N_6136,N_6927);
or U7827 (N_7827,N_6516,N_6398);
and U7828 (N_7828,N_6211,N_6327);
or U7829 (N_7829,N_6467,N_6653);
nor U7830 (N_7830,N_6112,N_6954);
and U7831 (N_7831,N_6250,N_6407);
nand U7832 (N_7832,N_6012,N_6593);
xor U7833 (N_7833,N_6865,N_6740);
xor U7834 (N_7834,N_6198,N_6231);
and U7835 (N_7835,N_6138,N_6115);
nor U7836 (N_7836,N_6499,N_6332);
nand U7837 (N_7837,N_6778,N_6095);
xnor U7838 (N_7838,N_6371,N_6929);
or U7839 (N_7839,N_6946,N_6969);
nor U7840 (N_7840,N_6287,N_6694);
nor U7841 (N_7841,N_6305,N_6068);
nor U7842 (N_7842,N_6014,N_6428);
nand U7843 (N_7843,N_6293,N_6844);
nor U7844 (N_7844,N_6492,N_6475);
nand U7845 (N_7845,N_6908,N_6002);
xor U7846 (N_7846,N_6734,N_6338);
xnor U7847 (N_7847,N_6827,N_6974);
nor U7848 (N_7848,N_6113,N_6042);
nor U7849 (N_7849,N_6946,N_6878);
nand U7850 (N_7850,N_6050,N_6846);
nand U7851 (N_7851,N_6351,N_6843);
xnor U7852 (N_7852,N_6455,N_6368);
and U7853 (N_7853,N_6450,N_6022);
nand U7854 (N_7854,N_6403,N_6775);
and U7855 (N_7855,N_6314,N_6484);
and U7856 (N_7856,N_6748,N_6983);
and U7857 (N_7857,N_6544,N_6246);
and U7858 (N_7858,N_6991,N_6219);
nand U7859 (N_7859,N_6810,N_6427);
xnor U7860 (N_7860,N_6291,N_6322);
nor U7861 (N_7861,N_6249,N_6357);
nor U7862 (N_7862,N_6875,N_6954);
xor U7863 (N_7863,N_6577,N_6300);
xor U7864 (N_7864,N_6004,N_6788);
nand U7865 (N_7865,N_6722,N_6077);
or U7866 (N_7866,N_6018,N_6922);
or U7867 (N_7867,N_6114,N_6109);
and U7868 (N_7868,N_6991,N_6920);
nand U7869 (N_7869,N_6180,N_6280);
nand U7870 (N_7870,N_6325,N_6361);
nand U7871 (N_7871,N_6973,N_6403);
or U7872 (N_7872,N_6783,N_6254);
or U7873 (N_7873,N_6934,N_6722);
nand U7874 (N_7874,N_6819,N_6358);
nor U7875 (N_7875,N_6042,N_6871);
nand U7876 (N_7876,N_6682,N_6335);
or U7877 (N_7877,N_6188,N_6579);
or U7878 (N_7878,N_6587,N_6095);
nor U7879 (N_7879,N_6891,N_6254);
xnor U7880 (N_7880,N_6335,N_6861);
and U7881 (N_7881,N_6154,N_6250);
nor U7882 (N_7882,N_6397,N_6624);
xor U7883 (N_7883,N_6460,N_6461);
nand U7884 (N_7884,N_6996,N_6636);
and U7885 (N_7885,N_6524,N_6030);
xnor U7886 (N_7886,N_6801,N_6561);
or U7887 (N_7887,N_6714,N_6138);
nand U7888 (N_7888,N_6334,N_6522);
xnor U7889 (N_7889,N_6701,N_6606);
or U7890 (N_7890,N_6856,N_6254);
and U7891 (N_7891,N_6906,N_6072);
or U7892 (N_7892,N_6311,N_6367);
or U7893 (N_7893,N_6105,N_6559);
xor U7894 (N_7894,N_6931,N_6364);
and U7895 (N_7895,N_6682,N_6990);
nand U7896 (N_7896,N_6622,N_6623);
xor U7897 (N_7897,N_6053,N_6067);
nor U7898 (N_7898,N_6036,N_6873);
nor U7899 (N_7899,N_6680,N_6575);
or U7900 (N_7900,N_6076,N_6991);
xor U7901 (N_7901,N_6225,N_6665);
nor U7902 (N_7902,N_6662,N_6435);
nand U7903 (N_7903,N_6032,N_6678);
or U7904 (N_7904,N_6010,N_6108);
nor U7905 (N_7905,N_6308,N_6521);
nor U7906 (N_7906,N_6114,N_6575);
or U7907 (N_7907,N_6855,N_6185);
and U7908 (N_7908,N_6984,N_6897);
or U7909 (N_7909,N_6681,N_6827);
nand U7910 (N_7910,N_6979,N_6005);
and U7911 (N_7911,N_6642,N_6647);
and U7912 (N_7912,N_6821,N_6825);
xnor U7913 (N_7913,N_6445,N_6146);
nand U7914 (N_7914,N_6603,N_6089);
nor U7915 (N_7915,N_6401,N_6093);
nor U7916 (N_7916,N_6706,N_6837);
nor U7917 (N_7917,N_6619,N_6457);
or U7918 (N_7918,N_6681,N_6186);
nor U7919 (N_7919,N_6416,N_6055);
and U7920 (N_7920,N_6406,N_6601);
xnor U7921 (N_7921,N_6621,N_6743);
nand U7922 (N_7922,N_6757,N_6859);
or U7923 (N_7923,N_6896,N_6341);
or U7924 (N_7924,N_6108,N_6133);
or U7925 (N_7925,N_6063,N_6987);
or U7926 (N_7926,N_6077,N_6640);
nor U7927 (N_7927,N_6104,N_6652);
or U7928 (N_7928,N_6918,N_6070);
nand U7929 (N_7929,N_6110,N_6365);
or U7930 (N_7930,N_6299,N_6279);
nor U7931 (N_7931,N_6420,N_6766);
xnor U7932 (N_7932,N_6045,N_6989);
and U7933 (N_7933,N_6756,N_6839);
nand U7934 (N_7934,N_6860,N_6252);
and U7935 (N_7935,N_6128,N_6155);
or U7936 (N_7936,N_6005,N_6503);
and U7937 (N_7937,N_6271,N_6608);
and U7938 (N_7938,N_6105,N_6684);
nand U7939 (N_7939,N_6942,N_6717);
nand U7940 (N_7940,N_6583,N_6472);
and U7941 (N_7941,N_6211,N_6043);
nor U7942 (N_7942,N_6302,N_6866);
and U7943 (N_7943,N_6762,N_6345);
xnor U7944 (N_7944,N_6080,N_6567);
or U7945 (N_7945,N_6562,N_6825);
nand U7946 (N_7946,N_6708,N_6496);
or U7947 (N_7947,N_6898,N_6131);
xor U7948 (N_7948,N_6776,N_6088);
xor U7949 (N_7949,N_6793,N_6478);
nor U7950 (N_7950,N_6249,N_6800);
or U7951 (N_7951,N_6515,N_6212);
nor U7952 (N_7952,N_6188,N_6607);
nor U7953 (N_7953,N_6367,N_6606);
or U7954 (N_7954,N_6266,N_6013);
nor U7955 (N_7955,N_6730,N_6441);
nor U7956 (N_7956,N_6331,N_6034);
nand U7957 (N_7957,N_6413,N_6704);
or U7958 (N_7958,N_6119,N_6261);
nor U7959 (N_7959,N_6454,N_6922);
nor U7960 (N_7960,N_6891,N_6098);
and U7961 (N_7961,N_6628,N_6928);
nand U7962 (N_7962,N_6624,N_6267);
and U7963 (N_7963,N_6770,N_6762);
and U7964 (N_7964,N_6058,N_6320);
nor U7965 (N_7965,N_6910,N_6509);
or U7966 (N_7966,N_6308,N_6439);
nand U7967 (N_7967,N_6516,N_6973);
or U7968 (N_7968,N_6300,N_6089);
nand U7969 (N_7969,N_6580,N_6707);
and U7970 (N_7970,N_6561,N_6333);
and U7971 (N_7971,N_6996,N_6044);
xor U7972 (N_7972,N_6474,N_6806);
and U7973 (N_7973,N_6292,N_6573);
xnor U7974 (N_7974,N_6946,N_6926);
xnor U7975 (N_7975,N_6659,N_6255);
xor U7976 (N_7976,N_6009,N_6594);
nor U7977 (N_7977,N_6818,N_6949);
nand U7978 (N_7978,N_6821,N_6340);
and U7979 (N_7979,N_6279,N_6583);
or U7980 (N_7980,N_6912,N_6325);
and U7981 (N_7981,N_6281,N_6918);
nand U7982 (N_7982,N_6270,N_6065);
and U7983 (N_7983,N_6804,N_6163);
nand U7984 (N_7984,N_6082,N_6405);
nor U7985 (N_7985,N_6566,N_6417);
nand U7986 (N_7986,N_6142,N_6243);
xor U7987 (N_7987,N_6252,N_6302);
nor U7988 (N_7988,N_6947,N_6631);
and U7989 (N_7989,N_6805,N_6705);
and U7990 (N_7990,N_6112,N_6075);
or U7991 (N_7991,N_6136,N_6171);
nand U7992 (N_7992,N_6096,N_6413);
nand U7993 (N_7993,N_6551,N_6432);
and U7994 (N_7994,N_6625,N_6295);
nor U7995 (N_7995,N_6579,N_6516);
and U7996 (N_7996,N_6631,N_6425);
nand U7997 (N_7997,N_6291,N_6199);
or U7998 (N_7998,N_6539,N_6025);
and U7999 (N_7999,N_6679,N_6128);
xnor U8000 (N_8000,N_7116,N_7204);
and U8001 (N_8001,N_7548,N_7009);
and U8002 (N_8002,N_7392,N_7743);
nand U8003 (N_8003,N_7682,N_7039);
xnor U8004 (N_8004,N_7805,N_7187);
nand U8005 (N_8005,N_7539,N_7549);
and U8006 (N_8006,N_7339,N_7030);
or U8007 (N_8007,N_7178,N_7474);
nand U8008 (N_8008,N_7780,N_7818);
or U8009 (N_8009,N_7603,N_7936);
or U8010 (N_8010,N_7156,N_7438);
nor U8011 (N_8011,N_7348,N_7031);
nor U8012 (N_8012,N_7423,N_7913);
nand U8013 (N_8013,N_7279,N_7925);
and U8014 (N_8014,N_7674,N_7550);
xor U8015 (N_8015,N_7821,N_7620);
or U8016 (N_8016,N_7498,N_7753);
and U8017 (N_8017,N_7654,N_7459);
or U8018 (N_8018,N_7355,N_7115);
nand U8019 (N_8019,N_7749,N_7789);
or U8020 (N_8020,N_7737,N_7456);
nor U8021 (N_8021,N_7250,N_7242);
nor U8022 (N_8022,N_7867,N_7436);
nand U8023 (N_8023,N_7838,N_7827);
nor U8024 (N_8024,N_7061,N_7522);
nand U8025 (N_8025,N_7767,N_7702);
xor U8026 (N_8026,N_7732,N_7139);
or U8027 (N_8027,N_7980,N_7247);
nor U8028 (N_8028,N_7811,N_7306);
or U8029 (N_8029,N_7680,N_7644);
nand U8030 (N_8030,N_7834,N_7312);
nand U8031 (N_8031,N_7128,N_7055);
or U8032 (N_8032,N_7516,N_7470);
nand U8033 (N_8033,N_7349,N_7280);
xnor U8034 (N_8034,N_7712,N_7440);
or U8035 (N_8035,N_7119,N_7077);
or U8036 (N_8036,N_7759,N_7611);
nand U8037 (N_8037,N_7006,N_7054);
and U8038 (N_8038,N_7394,N_7016);
xor U8039 (N_8039,N_7940,N_7506);
nor U8040 (N_8040,N_7685,N_7018);
xor U8041 (N_8041,N_7511,N_7337);
nand U8042 (N_8042,N_7001,N_7199);
or U8043 (N_8043,N_7399,N_7807);
and U8044 (N_8044,N_7802,N_7798);
xnor U8045 (N_8045,N_7331,N_7970);
nand U8046 (N_8046,N_7426,N_7836);
nor U8047 (N_8047,N_7884,N_7776);
and U8048 (N_8048,N_7701,N_7037);
xnor U8049 (N_8049,N_7411,N_7959);
and U8050 (N_8050,N_7092,N_7461);
or U8051 (N_8051,N_7666,N_7915);
xor U8052 (N_8052,N_7024,N_7245);
and U8053 (N_8053,N_7237,N_7546);
xor U8054 (N_8054,N_7453,N_7131);
and U8055 (N_8055,N_7047,N_7332);
and U8056 (N_8056,N_7314,N_7471);
nand U8057 (N_8057,N_7317,N_7750);
or U8058 (N_8058,N_7891,N_7845);
nor U8059 (N_8059,N_7153,N_7171);
nor U8060 (N_8060,N_7130,N_7466);
and U8061 (N_8061,N_7142,N_7484);
and U8062 (N_8062,N_7883,N_7552);
xnor U8063 (N_8063,N_7997,N_7598);
nor U8064 (N_8064,N_7259,N_7034);
nor U8065 (N_8065,N_7212,N_7599);
xor U8066 (N_8066,N_7170,N_7447);
nand U8067 (N_8067,N_7448,N_7455);
or U8068 (N_8068,N_7725,N_7796);
nor U8069 (N_8069,N_7833,N_7602);
nand U8070 (N_8070,N_7158,N_7008);
nor U8071 (N_8071,N_7748,N_7076);
xnor U8072 (N_8072,N_7521,N_7637);
and U8073 (N_8073,N_7433,N_7782);
xor U8074 (N_8074,N_7799,N_7487);
nor U8075 (N_8075,N_7882,N_7129);
or U8076 (N_8076,N_7995,N_7230);
xnor U8077 (N_8077,N_7301,N_7169);
and U8078 (N_8078,N_7790,N_7005);
nor U8079 (N_8079,N_7416,N_7662);
nor U8080 (N_8080,N_7120,N_7901);
and U8081 (N_8081,N_7262,N_7996);
nor U8082 (N_8082,N_7870,N_7389);
nand U8083 (N_8083,N_7402,N_7098);
nor U8084 (N_8084,N_7072,N_7203);
xor U8085 (N_8085,N_7999,N_7698);
xnor U8086 (N_8086,N_7524,N_7612);
nor U8087 (N_8087,N_7189,N_7815);
nand U8088 (N_8088,N_7002,N_7106);
and U8089 (N_8089,N_7021,N_7617);
and U8090 (N_8090,N_7136,N_7198);
nand U8091 (N_8091,N_7963,N_7645);
or U8092 (N_8092,N_7810,N_7515);
and U8093 (N_8093,N_7500,N_7291);
xor U8094 (N_8094,N_7185,N_7669);
nor U8095 (N_8095,N_7509,N_7017);
or U8096 (N_8096,N_7874,N_7308);
xor U8097 (N_8097,N_7555,N_7226);
or U8098 (N_8098,N_7482,N_7731);
and U8099 (N_8099,N_7003,N_7921);
and U8100 (N_8100,N_7825,N_7544);
nor U8101 (N_8101,N_7571,N_7462);
nor U8102 (N_8102,N_7792,N_7880);
nor U8103 (N_8103,N_7764,N_7257);
and U8104 (N_8104,N_7860,N_7049);
nor U8105 (N_8105,N_7920,N_7930);
nor U8106 (N_8106,N_7892,N_7080);
nor U8107 (N_8107,N_7527,N_7956);
or U8108 (N_8108,N_7371,N_7241);
nor U8109 (N_8109,N_7268,N_7961);
nand U8110 (N_8110,N_7557,N_7797);
nand U8111 (N_8111,N_7889,N_7275);
xnor U8112 (N_8112,N_7027,N_7528);
xor U8113 (N_8113,N_7982,N_7504);
and U8114 (N_8114,N_7298,N_7852);
nor U8115 (N_8115,N_7859,N_7358);
nor U8116 (N_8116,N_7763,N_7962);
and U8117 (N_8117,N_7619,N_7992);
and U8118 (N_8118,N_7781,N_7007);
or U8119 (N_8119,N_7014,N_7439);
xnor U8120 (N_8120,N_7386,N_7861);
and U8121 (N_8121,N_7765,N_7795);
nor U8122 (N_8122,N_7512,N_7957);
or U8123 (N_8123,N_7812,N_7288);
or U8124 (N_8124,N_7026,N_7218);
and U8125 (N_8125,N_7430,N_7499);
nand U8126 (N_8126,N_7652,N_7217);
xor U8127 (N_8127,N_7019,N_7053);
and U8128 (N_8128,N_7363,N_7517);
xor U8129 (N_8129,N_7322,N_7877);
nor U8130 (N_8130,N_7850,N_7532);
or U8131 (N_8131,N_7473,N_7761);
nor U8132 (N_8132,N_7045,N_7633);
nor U8133 (N_8133,N_7066,N_7965);
and U8134 (N_8134,N_7887,N_7973);
or U8135 (N_8135,N_7117,N_7243);
nand U8136 (N_8136,N_7103,N_7932);
and U8137 (N_8137,N_7425,N_7908);
xor U8138 (N_8138,N_7719,N_7161);
nand U8139 (N_8139,N_7292,N_7104);
nand U8140 (N_8140,N_7122,N_7406);
nor U8141 (N_8141,N_7491,N_7286);
nor U8142 (N_8142,N_7109,N_7254);
and U8143 (N_8143,N_7351,N_7927);
nor U8144 (N_8144,N_7771,N_7862);
and U8145 (N_8145,N_7478,N_7563);
nor U8146 (N_8146,N_7900,N_7824);
nor U8147 (N_8147,N_7952,N_7646);
and U8148 (N_8148,N_7475,N_7046);
nand U8149 (N_8149,N_7739,N_7559);
xor U8150 (N_8150,N_7875,N_7543);
xor U8151 (N_8151,N_7533,N_7806);
or U8152 (N_8152,N_7266,N_7064);
nand U8153 (N_8153,N_7094,N_7486);
or U8154 (N_8154,N_7197,N_7586);
nor U8155 (N_8155,N_7377,N_7830);
nor U8156 (N_8156,N_7011,N_7935);
and U8157 (N_8157,N_7148,N_7040);
or U8158 (N_8158,N_7012,N_7396);
xor U8159 (N_8159,N_7225,N_7525);
or U8160 (N_8160,N_7388,N_7686);
nand U8161 (N_8161,N_7706,N_7446);
and U8162 (N_8162,N_7488,N_7597);
xor U8163 (N_8163,N_7144,N_7989);
nand U8164 (N_8164,N_7979,N_7950);
xor U8165 (N_8165,N_7490,N_7657);
nand U8166 (N_8166,N_7501,N_7541);
or U8167 (N_8167,N_7653,N_7369);
and U8168 (N_8168,N_7335,N_7100);
nor U8169 (N_8169,N_7760,N_7508);
xor U8170 (N_8170,N_7420,N_7934);
and U8171 (N_8171,N_7710,N_7492);
nor U8172 (N_8172,N_7945,N_7062);
and U8173 (N_8173,N_7215,N_7639);
xnor U8174 (N_8174,N_7274,N_7697);
or U8175 (N_8175,N_7804,N_7162);
and U8176 (N_8176,N_7881,N_7551);
or U8177 (N_8177,N_7495,N_7736);
nand U8178 (N_8178,N_7323,N_7670);
and U8179 (N_8179,N_7942,N_7744);
and U8180 (N_8180,N_7582,N_7253);
nand U8181 (N_8181,N_7756,N_7630);
xor U8182 (N_8182,N_7362,N_7088);
or U8183 (N_8183,N_7069,N_7147);
and U8184 (N_8184,N_7616,N_7407);
and U8185 (N_8185,N_7256,N_7890);
xor U8186 (N_8186,N_7841,N_7871);
nor U8187 (N_8187,N_7745,N_7886);
xor U8188 (N_8188,N_7099,N_7542);
nor U8189 (N_8189,N_7329,N_7676);
xnor U8190 (N_8190,N_7318,N_7667);
or U8191 (N_8191,N_7829,N_7477);
xnor U8192 (N_8192,N_7664,N_7071);
or U8193 (N_8193,N_7346,N_7740);
xor U8194 (N_8194,N_7758,N_7704);
nor U8195 (N_8195,N_7911,N_7735);
or U8196 (N_8196,N_7287,N_7726);
or U8197 (N_8197,N_7300,N_7648);
or U8198 (N_8198,N_7954,N_7537);
xor U8199 (N_8199,N_7151,N_7975);
nor U8200 (N_8200,N_7857,N_7757);
nor U8201 (N_8201,N_7787,N_7352);
or U8202 (N_8202,N_7568,N_7101);
nand U8203 (N_8203,N_7978,N_7336);
xor U8204 (N_8204,N_7953,N_7819);
xor U8205 (N_8205,N_7413,N_7342);
nand U8206 (N_8206,N_7554,N_7350);
and U8207 (N_8207,N_7727,N_7502);
and U8208 (N_8208,N_7232,N_7600);
and U8209 (N_8209,N_7949,N_7747);
and U8210 (N_8210,N_7847,N_7803);
and U8211 (N_8211,N_7343,N_7194);
or U8212 (N_8212,N_7910,N_7041);
and U8213 (N_8213,N_7746,N_7347);
xnor U8214 (N_8214,N_7025,N_7097);
nor U8215 (N_8215,N_7239,N_7734);
and U8216 (N_8216,N_7843,N_7483);
nor U8217 (N_8217,N_7140,N_7822);
xnor U8218 (N_8218,N_7281,N_7345);
and U8219 (N_8219,N_7248,N_7831);
or U8220 (N_8220,N_7449,N_7236);
xor U8221 (N_8221,N_7359,N_7052);
nand U8222 (N_8222,N_7625,N_7896);
and U8223 (N_8223,N_7816,N_7926);
nor U8224 (N_8224,N_7742,N_7933);
nor U8225 (N_8225,N_7944,N_7547);
nor U8226 (N_8226,N_7135,N_7378);
xor U8227 (N_8227,N_7983,N_7260);
and U8228 (N_8228,N_7655,N_7087);
xnor U8229 (N_8229,N_7366,N_7604);
or U8230 (N_8230,N_7174,N_7154);
or U8231 (N_8231,N_7872,N_7899);
and U8232 (N_8232,N_7919,N_7692);
and U8233 (N_8233,N_7290,N_7641);
xor U8234 (N_8234,N_7155,N_7418);
nand U8235 (N_8235,N_7057,N_7898);
nor U8236 (N_8236,N_7650,N_7075);
and U8237 (N_8237,N_7723,N_7985);
nand U8238 (N_8238,N_7417,N_7826);
nand U8239 (N_8239,N_7333,N_7846);
nor U8240 (N_8240,N_7649,N_7793);
xor U8241 (N_8241,N_7714,N_7114);
nand U8242 (N_8242,N_7397,N_7481);
xnor U8243 (N_8243,N_7374,N_7905);
and U8244 (N_8244,N_7390,N_7914);
xor U8245 (N_8245,N_7707,N_7231);
nor U8246 (N_8246,N_7381,N_7160);
nand U8247 (N_8247,N_7564,N_7186);
nand U8248 (N_8248,N_7370,N_7060);
nor U8249 (N_8249,N_7167,N_7022);
xnor U8250 (N_8250,N_7111,N_7623);
or U8251 (N_8251,N_7864,N_7938);
nor U8252 (N_8252,N_7752,N_7876);
nand U8253 (N_8253,N_7361,N_7638);
xnor U8254 (N_8254,N_7036,N_7718);
and U8255 (N_8255,N_7327,N_7699);
and U8256 (N_8256,N_7238,N_7705);
nand U8257 (N_8257,N_7494,N_7709);
nor U8258 (N_8258,N_7485,N_7338);
xnor U8259 (N_8259,N_7741,N_7182);
and U8260 (N_8260,N_7032,N_7520);
xor U8261 (N_8261,N_7627,N_7689);
nand U8262 (N_8262,N_7738,N_7814);
nor U8263 (N_8263,N_7496,N_7809);
and U8264 (N_8264,N_7033,N_7283);
nor U8265 (N_8265,N_7794,N_7321);
and U8266 (N_8266,N_7774,N_7263);
and U8267 (N_8267,N_7133,N_7773);
or U8268 (N_8268,N_7538,N_7583);
nand U8269 (N_8269,N_7866,N_7137);
and U8270 (N_8270,N_7590,N_7570);
xnor U8271 (N_8271,N_7578,N_7255);
or U8272 (N_8272,N_7353,N_7679);
xnor U8273 (N_8273,N_7832,N_7192);
or U8274 (N_8274,N_7184,N_7783);
xnor U8275 (N_8275,N_7319,N_7958);
and U8276 (N_8276,N_7118,N_7434);
nor U8277 (N_8277,N_7587,N_7994);
and U8278 (N_8278,N_7621,N_7344);
xor U8279 (N_8279,N_7166,N_7659);
or U8280 (N_8280,N_7183,N_7304);
nor U8281 (N_8281,N_7868,N_7681);
xnor U8282 (N_8282,N_7907,N_7373);
nor U8283 (N_8283,N_7320,N_7000);
or U8284 (N_8284,N_7720,N_7435);
nor U8285 (N_8285,N_7400,N_7063);
and U8286 (N_8286,N_7672,N_7405);
nand U8287 (N_8287,N_7376,N_7558);
or U8288 (N_8288,N_7993,N_7912);
nand U8289 (N_8289,N_7651,N_7693);
nor U8290 (N_8290,N_7922,N_7207);
and U8291 (N_8291,N_7261,N_7668);
nor U8292 (N_8292,N_7581,N_7839);
nor U8293 (N_8293,N_7665,N_7640);
or U8294 (N_8294,N_7778,N_7375);
xnor U8295 (N_8295,N_7152,N_7974);
and U8296 (N_8296,N_7643,N_7415);
nand U8297 (N_8297,N_7856,N_7408);
xor U8298 (N_8298,N_7429,N_7626);
nand U8299 (N_8299,N_7729,N_7931);
nor U8300 (N_8300,N_7510,N_7393);
xnor U8301 (N_8301,N_7089,N_7923);
nor U8302 (N_8302,N_7365,N_7125);
or U8303 (N_8303,N_7168,N_7458);
nand U8304 (N_8304,N_7364,N_7086);
or U8305 (N_8305,N_7981,N_7817);
or U8306 (N_8306,N_7093,N_7716);
nor U8307 (N_8307,N_7085,N_7941);
nand U8308 (N_8308,N_7132,N_7565);
and U8309 (N_8309,N_7837,N_7696);
xor U8310 (N_8310,N_7951,N_7315);
xnor U8311 (N_8311,N_7529,N_7636);
nor U8312 (N_8312,N_7713,N_7294);
nor U8313 (N_8313,N_7251,N_7095);
and U8314 (N_8314,N_7535,N_7715);
and U8315 (N_8315,N_7946,N_7592);
or U8316 (N_8316,N_7035,N_7939);
and U8317 (N_8317,N_7801,N_7800);
nand U8318 (N_8318,N_7269,N_7770);
xnor U8319 (N_8319,N_7082,N_7947);
xor U8320 (N_8320,N_7276,N_7694);
nand U8321 (N_8321,N_7410,N_7059);
xor U8322 (N_8322,N_7179,N_7791);
xnor U8323 (N_8323,N_7675,N_7937);
xor U8324 (N_8324,N_7531,N_7043);
and U8325 (N_8325,N_7788,N_7163);
and U8326 (N_8326,N_7505,N_7865);
nor U8327 (N_8327,N_7894,N_7497);
nand U8328 (N_8328,N_7855,N_7146);
xnor U8329 (N_8329,N_7190,N_7191);
or U8330 (N_8330,N_7661,N_7445);
and U8331 (N_8331,N_7372,N_7955);
nand U8332 (N_8332,N_7545,N_7414);
nor U8333 (N_8333,N_7084,N_7398);
or U8334 (N_8334,N_7569,N_7195);
or U8335 (N_8335,N_7690,N_7988);
and U8336 (N_8336,N_7267,N_7313);
and U8337 (N_8337,N_7476,N_7042);
nor U8338 (N_8338,N_7663,N_7244);
xnor U8339 (N_8339,N_7479,N_7683);
nand U8340 (N_8340,N_7273,N_7293);
xor U8341 (N_8341,N_7472,N_7228);
nor U8342 (N_8342,N_7235,N_7984);
xnor U8343 (N_8343,N_7628,N_7223);
nor U8344 (N_8344,N_7305,N_7096);
or U8345 (N_8345,N_7823,N_7177);
or U8346 (N_8346,N_7173,N_7635);
nor U8347 (N_8347,N_7383,N_7507);
nor U8348 (N_8348,N_7585,N_7688);
nor U8349 (N_8349,N_7437,N_7772);
xor U8350 (N_8350,N_7722,N_7977);
and U8351 (N_8351,N_7991,N_7213);
or U8352 (N_8352,N_7401,N_7584);
xor U8353 (N_8353,N_7121,N_7172);
xnor U8354 (N_8354,N_7610,N_7906);
nor U8355 (N_8355,N_7711,N_7530);
or U8356 (N_8356,N_7201,N_7330);
nand U8357 (N_8357,N_7380,N_7278);
xor U8358 (N_8358,N_7766,N_7840);
xnor U8359 (N_8359,N_7879,N_7575);
xnor U8360 (N_8360,N_7065,N_7102);
and U8361 (N_8361,N_7264,N_7658);
nor U8362 (N_8362,N_7755,N_7929);
nand U8363 (N_8363,N_7677,N_7296);
nand U8364 (N_8364,N_7157,N_7835);
nor U8365 (N_8365,N_7023,N_7210);
xor U8366 (N_8366,N_7591,N_7219);
nand U8367 (N_8367,N_7249,N_7897);
or U8368 (N_8368,N_7948,N_7441);
xnor U8369 (N_8369,N_7216,N_7678);
nand U8370 (N_8370,N_7367,N_7205);
nor U8371 (N_8371,N_7684,N_7721);
xor U8372 (N_8372,N_7854,N_7044);
and U8373 (N_8373,N_7695,N_7960);
nand U8374 (N_8374,N_7387,N_7334);
nand U8375 (N_8375,N_7326,N_7309);
xor U8376 (N_8376,N_7556,N_7056);
or U8377 (N_8377,N_7385,N_7717);
or U8378 (N_8378,N_7902,N_7893);
xor U8379 (N_8379,N_7966,N_7450);
xnor U8380 (N_8380,N_7574,N_7526);
nand U8381 (N_8381,N_7038,N_7967);
xor U8382 (N_8382,N_7567,N_7395);
nor U8383 (N_8383,N_7067,N_7751);
or U8384 (N_8384,N_7769,N_7990);
and U8385 (N_8385,N_7258,N_7431);
and U8386 (N_8386,N_7489,N_7368);
xor U8387 (N_8387,N_7126,N_7724);
nand U8388 (N_8388,N_7779,N_7849);
or U8389 (N_8389,N_7382,N_7594);
nor U8390 (N_8390,N_7175,N_7842);
nor U8391 (N_8391,N_7432,N_7700);
nor U8392 (N_8392,N_7596,N_7324);
or U8393 (N_8393,N_7762,N_7220);
nand U8394 (N_8394,N_7316,N_7134);
or U8395 (N_8395,N_7613,N_7730);
nand U8396 (N_8396,N_7443,N_7200);
nor U8397 (N_8397,N_7081,N_7622);
and U8398 (N_8398,N_7196,N_7058);
nand U8399 (N_8399,N_7895,N_7422);
nor U8400 (N_8400,N_7233,N_7328);
xor U8401 (N_8401,N_7004,N_7986);
or U8402 (N_8402,N_7277,N_7869);
or U8403 (N_8403,N_7340,N_7561);
nand U8404 (N_8404,N_7493,N_7660);
and U8405 (N_8405,N_7297,N_7252);
xor U8406 (N_8406,N_7851,N_7124);
or U8407 (N_8407,N_7123,N_7284);
xnor U8408 (N_8408,N_7768,N_7624);
xnor U8409 (N_8409,N_7853,N_7518);
and U8410 (N_8410,N_7050,N_7924);
or U8411 (N_8411,N_7885,N_7519);
nand U8412 (N_8412,N_7384,N_7785);
or U8413 (N_8413,N_7227,N_7311);
nor U8414 (N_8414,N_7464,N_7605);
nand U8415 (N_8415,N_7673,N_7618);
and U8416 (N_8416,N_7271,N_7234);
nand U8417 (N_8417,N_7409,N_7015);
xor U8418 (N_8418,N_7391,N_7964);
xor U8419 (N_8419,N_7607,N_7615);
xor U8420 (N_8420,N_7976,N_7444);
nor U8421 (N_8421,N_7202,N_7632);
or U8422 (N_8422,N_7246,N_7808);
nor U8423 (N_8423,N_7928,N_7180);
and U8424 (N_8424,N_7307,N_7229);
or U8425 (N_8425,N_7579,N_7010);
xor U8426 (N_8426,N_7536,N_7480);
or U8427 (N_8427,N_7642,N_7208);
and U8428 (N_8428,N_7028,N_7211);
nand U8429 (N_8429,N_7138,N_7534);
nand U8430 (N_8430,N_7608,N_7848);
nor U8431 (N_8431,N_7820,N_7090);
xnor U8432 (N_8432,N_7858,N_7074);
and U8433 (N_8433,N_7113,N_7159);
and U8434 (N_8434,N_7013,N_7468);
and U8435 (N_8435,N_7589,N_7553);
and U8436 (N_8436,N_7404,N_7091);
and U8437 (N_8437,N_7452,N_7784);
nor U8438 (N_8438,N_7909,N_7222);
or U8439 (N_8439,N_7454,N_7671);
or U8440 (N_8440,N_7073,N_7844);
nor U8441 (N_8441,N_7593,N_7514);
xor U8442 (N_8442,N_7068,N_7634);
and U8443 (N_8443,N_7656,N_7968);
or U8444 (N_8444,N_7164,N_7969);
nor U8445 (N_8445,N_7562,N_7703);
nor U8446 (N_8446,N_7427,N_7609);
nand U8447 (N_8447,N_7083,N_7360);
or U8448 (N_8448,N_7580,N_7595);
or U8449 (N_8449,N_7873,N_7888);
and U8450 (N_8450,N_7469,N_7112);
nor U8451 (N_8451,N_7356,N_7828);
or U8452 (N_8452,N_7270,N_7051);
or U8453 (N_8453,N_7165,N_7775);
or U8454 (N_8454,N_7465,N_7987);
and U8455 (N_8455,N_7424,N_7786);
xor U8456 (N_8456,N_7467,N_7209);
and U8457 (N_8457,N_7149,N_7457);
nor U8458 (N_8458,N_7754,N_7214);
and U8459 (N_8459,N_7078,N_7560);
nor U8460 (N_8460,N_7357,N_7206);
nand U8461 (N_8461,N_7631,N_7576);
or U8462 (N_8462,N_7295,N_7573);
nor U8463 (N_8463,N_7412,N_7419);
or U8464 (N_8464,N_7513,N_7647);
nand U8465 (N_8465,N_7299,N_7903);
xnor U8466 (N_8466,N_7325,N_7460);
and U8467 (N_8467,N_7998,N_7606);
or U8468 (N_8468,N_7303,N_7916);
or U8469 (N_8469,N_7691,N_7379);
nor U8470 (N_8470,N_7127,N_7289);
nor U8471 (N_8471,N_7813,N_7588);
and U8472 (N_8472,N_7421,N_7141);
xor U8473 (N_8473,N_7878,N_7777);
nand U8474 (N_8474,N_7943,N_7224);
nand U8475 (N_8475,N_7282,N_7020);
xnor U8476 (N_8476,N_7572,N_7070);
or U8477 (N_8477,N_7904,N_7079);
nand U8478 (N_8478,N_7442,N_7577);
or U8479 (N_8479,N_7451,N_7687);
xor U8480 (N_8480,N_7221,N_7341);
nand U8481 (N_8481,N_7145,N_7403);
xnor U8482 (N_8482,N_7972,N_7971);
nand U8483 (N_8483,N_7272,N_7150);
nor U8484 (N_8484,N_7566,N_7601);
xor U8485 (N_8485,N_7863,N_7614);
and U8486 (N_8486,N_7265,N_7463);
nor U8487 (N_8487,N_7181,N_7048);
nand U8488 (N_8488,N_7918,N_7523);
and U8489 (N_8489,N_7108,N_7285);
xor U8490 (N_8490,N_7188,N_7629);
xnor U8491 (N_8491,N_7143,N_7540);
nor U8492 (N_8492,N_7728,N_7107);
nand U8493 (N_8493,N_7176,N_7733);
and U8494 (N_8494,N_7029,N_7354);
nor U8495 (N_8495,N_7708,N_7917);
nor U8496 (N_8496,N_7310,N_7105);
and U8497 (N_8497,N_7193,N_7428);
and U8498 (N_8498,N_7110,N_7503);
xnor U8499 (N_8499,N_7240,N_7302);
and U8500 (N_8500,N_7092,N_7970);
xor U8501 (N_8501,N_7800,N_7314);
nand U8502 (N_8502,N_7387,N_7712);
or U8503 (N_8503,N_7533,N_7397);
nor U8504 (N_8504,N_7509,N_7007);
and U8505 (N_8505,N_7354,N_7237);
or U8506 (N_8506,N_7168,N_7751);
nor U8507 (N_8507,N_7153,N_7665);
and U8508 (N_8508,N_7909,N_7512);
nor U8509 (N_8509,N_7834,N_7948);
or U8510 (N_8510,N_7195,N_7161);
and U8511 (N_8511,N_7091,N_7158);
nor U8512 (N_8512,N_7554,N_7772);
nor U8513 (N_8513,N_7689,N_7551);
xor U8514 (N_8514,N_7466,N_7841);
xnor U8515 (N_8515,N_7381,N_7214);
nor U8516 (N_8516,N_7141,N_7637);
xor U8517 (N_8517,N_7659,N_7003);
nand U8518 (N_8518,N_7186,N_7858);
nor U8519 (N_8519,N_7379,N_7863);
xor U8520 (N_8520,N_7752,N_7871);
and U8521 (N_8521,N_7619,N_7756);
xor U8522 (N_8522,N_7673,N_7693);
xor U8523 (N_8523,N_7923,N_7360);
and U8524 (N_8524,N_7554,N_7175);
xnor U8525 (N_8525,N_7173,N_7540);
or U8526 (N_8526,N_7050,N_7310);
nor U8527 (N_8527,N_7581,N_7631);
or U8528 (N_8528,N_7364,N_7713);
nor U8529 (N_8529,N_7752,N_7383);
and U8530 (N_8530,N_7864,N_7696);
nand U8531 (N_8531,N_7392,N_7996);
or U8532 (N_8532,N_7375,N_7135);
or U8533 (N_8533,N_7133,N_7947);
nand U8534 (N_8534,N_7905,N_7499);
or U8535 (N_8535,N_7536,N_7159);
nand U8536 (N_8536,N_7496,N_7996);
and U8537 (N_8537,N_7425,N_7056);
and U8538 (N_8538,N_7988,N_7030);
and U8539 (N_8539,N_7113,N_7093);
xor U8540 (N_8540,N_7177,N_7608);
xor U8541 (N_8541,N_7462,N_7119);
or U8542 (N_8542,N_7936,N_7341);
xnor U8543 (N_8543,N_7335,N_7649);
nor U8544 (N_8544,N_7815,N_7930);
nand U8545 (N_8545,N_7758,N_7411);
xor U8546 (N_8546,N_7458,N_7352);
xor U8547 (N_8547,N_7462,N_7700);
or U8548 (N_8548,N_7256,N_7954);
nand U8549 (N_8549,N_7999,N_7032);
nor U8550 (N_8550,N_7512,N_7714);
xor U8551 (N_8551,N_7822,N_7025);
or U8552 (N_8552,N_7719,N_7098);
nor U8553 (N_8553,N_7724,N_7677);
and U8554 (N_8554,N_7615,N_7557);
xor U8555 (N_8555,N_7418,N_7910);
or U8556 (N_8556,N_7051,N_7565);
xor U8557 (N_8557,N_7108,N_7064);
nor U8558 (N_8558,N_7238,N_7872);
nor U8559 (N_8559,N_7850,N_7860);
and U8560 (N_8560,N_7146,N_7822);
xnor U8561 (N_8561,N_7952,N_7578);
or U8562 (N_8562,N_7728,N_7050);
nor U8563 (N_8563,N_7067,N_7128);
xor U8564 (N_8564,N_7743,N_7290);
xnor U8565 (N_8565,N_7376,N_7369);
or U8566 (N_8566,N_7371,N_7501);
xnor U8567 (N_8567,N_7807,N_7277);
and U8568 (N_8568,N_7995,N_7992);
xnor U8569 (N_8569,N_7031,N_7581);
xor U8570 (N_8570,N_7115,N_7794);
nand U8571 (N_8571,N_7635,N_7575);
nor U8572 (N_8572,N_7082,N_7109);
nor U8573 (N_8573,N_7754,N_7176);
nand U8574 (N_8574,N_7804,N_7102);
nand U8575 (N_8575,N_7288,N_7742);
and U8576 (N_8576,N_7691,N_7771);
nand U8577 (N_8577,N_7909,N_7995);
nand U8578 (N_8578,N_7021,N_7806);
xnor U8579 (N_8579,N_7412,N_7482);
and U8580 (N_8580,N_7923,N_7829);
and U8581 (N_8581,N_7193,N_7313);
and U8582 (N_8582,N_7249,N_7232);
nor U8583 (N_8583,N_7827,N_7407);
nand U8584 (N_8584,N_7949,N_7557);
xor U8585 (N_8585,N_7847,N_7976);
nor U8586 (N_8586,N_7720,N_7193);
and U8587 (N_8587,N_7873,N_7727);
and U8588 (N_8588,N_7875,N_7508);
nand U8589 (N_8589,N_7032,N_7801);
xnor U8590 (N_8590,N_7420,N_7672);
nand U8591 (N_8591,N_7910,N_7413);
nand U8592 (N_8592,N_7096,N_7930);
nor U8593 (N_8593,N_7074,N_7079);
xor U8594 (N_8594,N_7383,N_7555);
and U8595 (N_8595,N_7044,N_7071);
xnor U8596 (N_8596,N_7104,N_7718);
nand U8597 (N_8597,N_7544,N_7166);
or U8598 (N_8598,N_7941,N_7348);
or U8599 (N_8599,N_7231,N_7280);
nor U8600 (N_8600,N_7776,N_7405);
nor U8601 (N_8601,N_7846,N_7701);
xor U8602 (N_8602,N_7965,N_7057);
and U8603 (N_8603,N_7340,N_7550);
nor U8604 (N_8604,N_7438,N_7544);
or U8605 (N_8605,N_7235,N_7346);
nor U8606 (N_8606,N_7619,N_7151);
xnor U8607 (N_8607,N_7442,N_7184);
or U8608 (N_8608,N_7447,N_7801);
or U8609 (N_8609,N_7644,N_7561);
or U8610 (N_8610,N_7061,N_7989);
xnor U8611 (N_8611,N_7834,N_7781);
nand U8612 (N_8612,N_7933,N_7731);
or U8613 (N_8613,N_7397,N_7453);
nor U8614 (N_8614,N_7400,N_7551);
xnor U8615 (N_8615,N_7513,N_7315);
or U8616 (N_8616,N_7491,N_7641);
xor U8617 (N_8617,N_7759,N_7069);
and U8618 (N_8618,N_7481,N_7991);
nand U8619 (N_8619,N_7909,N_7821);
nor U8620 (N_8620,N_7451,N_7112);
or U8621 (N_8621,N_7329,N_7659);
or U8622 (N_8622,N_7797,N_7618);
nor U8623 (N_8623,N_7963,N_7394);
xnor U8624 (N_8624,N_7813,N_7734);
xnor U8625 (N_8625,N_7173,N_7862);
and U8626 (N_8626,N_7450,N_7035);
nor U8627 (N_8627,N_7183,N_7671);
or U8628 (N_8628,N_7963,N_7451);
and U8629 (N_8629,N_7975,N_7898);
xor U8630 (N_8630,N_7046,N_7766);
nor U8631 (N_8631,N_7126,N_7512);
xnor U8632 (N_8632,N_7767,N_7566);
nand U8633 (N_8633,N_7777,N_7327);
nand U8634 (N_8634,N_7952,N_7589);
nor U8635 (N_8635,N_7014,N_7701);
or U8636 (N_8636,N_7512,N_7164);
or U8637 (N_8637,N_7342,N_7464);
and U8638 (N_8638,N_7703,N_7044);
nand U8639 (N_8639,N_7758,N_7070);
nor U8640 (N_8640,N_7800,N_7225);
and U8641 (N_8641,N_7791,N_7939);
or U8642 (N_8642,N_7878,N_7785);
xor U8643 (N_8643,N_7726,N_7696);
xnor U8644 (N_8644,N_7173,N_7488);
xnor U8645 (N_8645,N_7113,N_7428);
xnor U8646 (N_8646,N_7876,N_7352);
nand U8647 (N_8647,N_7136,N_7042);
and U8648 (N_8648,N_7971,N_7593);
xor U8649 (N_8649,N_7272,N_7849);
and U8650 (N_8650,N_7509,N_7202);
or U8651 (N_8651,N_7015,N_7281);
or U8652 (N_8652,N_7490,N_7768);
and U8653 (N_8653,N_7475,N_7190);
nand U8654 (N_8654,N_7061,N_7513);
nand U8655 (N_8655,N_7998,N_7162);
nor U8656 (N_8656,N_7264,N_7010);
xor U8657 (N_8657,N_7646,N_7384);
and U8658 (N_8658,N_7713,N_7513);
and U8659 (N_8659,N_7550,N_7977);
nor U8660 (N_8660,N_7033,N_7223);
nor U8661 (N_8661,N_7229,N_7197);
nand U8662 (N_8662,N_7040,N_7716);
and U8663 (N_8663,N_7873,N_7109);
nor U8664 (N_8664,N_7435,N_7914);
or U8665 (N_8665,N_7637,N_7129);
and U8666 (N_8666,N_7525,N_7061);
nor U8667 (N_8667,N_7634,N_7314);
nand U8668 (N_8668,N_7513,N_7177);
and U8669 (N_8669,N_7341,N_7413);
nand U8670 (N_8670,N_7252,N_7326);
and U8671 (N_8671,N_7360,N_7843);
nor U8672 (N_8672,N_7796,N_7774);
nor U8673 (N_8673,N_7835,N_7141);
nand U8674 (N_8674,N_7654,N_7044);
and U8675 (N_8675,N_7124,N_7729);
nand U8676 (N_8676,N_7979,N_7661);
and U8677 (N_8677,N_7418,N_7411);
nand U8678 (N_8678,N_7530,N_7014);
nor U8679 (N_8679,N_7512,N_7158);
nor U8680 (N_8680,N_7035,N_7690);
nand U8681 (N_8681,N_7753,N_7366);
and U8682 (N_8682,N_7413,N_7205);
or U8683 (N_8683,N_7218,N_7969);
and U8684 (N_8684,N_7514,N_7149);
and U8685 (N_8685,N_7140,N_7474);
and U8686 (N_8686,N_7803,N_7238);
and U8687 (N_8687,N_7023,N_7634);
nand U8688 (N_8688,N_7395,N_7488);
nand U8689 (N_8689,N_7195,N_7001);
or U8690 (N_8690,N_7011,N_7341);
xor U8691 (N_8691,N_7693,N_7280);
xnor U8692 (N_8692,N_7426,N_7271);
nor U8693 (N_8693,N_7546,N_7735);
and U8694 (N_8694,N_7425,N_7899);
or U8695 (N_8695,N_7226,N_7405);
nor U8696 (N_8696,N_7007,N_7726);
xnor U8697 (N_8697,N_7649,N_7329);
nand U8698 (N_8698,N_7725,N_7883);
and U8699 (N_8699,N_7657,N_7404);
nand U8700 (N_8700,N_7750,N_7134);
nand U8701 (N_8701,N_7474,N_7852);
and U8702 (N_8702,N_7213,N_7754);
nor U8703 (N_8703,N_7742,N_7761);
xor U8704 (N_8704,N_7301,N_7636);
nor U8705 (N_8705,N_7089,N_7644);
nand U8706 (N_8706,N_7081,N_7745);
xor U8707 (N_8707,N_7904,N_7418);
nor U8708 (N_8708,N_7371,N_7723);
and U8709 (N_8709,N_7146,N_7643);
nor U8710 (N_8710,N_7160,N_7724);
and U8711 (N_8711,N_7232,N_7158);
nand U8712 (N_8712,N_7518,N_7755);
nor U8713 (N_8713,N_7021,N_7457);
and U8714 (N_8714,N_7755,N_7868);
xor U8715 (N_8715,N_7734,N_7894);
or U8716 (N_8716,N_7355,N_7414);
nand U8717 (N_8717,N_7367,N_7968);
and U8718 (N_8718,N_7805,N_7682);
xor U8719 (N_8719,N_7982,N_7369);
or U8720 (N_8720,N_7675,N_7162);
or U8721 (N_8721,N_7191,N_7736);
xnor U8722 (N_8722,N_7610,N_7314);
nor U8723 (N_8723,N_7956,N_7104);
nor U8724 (N_8724,N_7566,N_7811);
nand U8725 (N_8725,N_7827,N_7061);
xor U8726 (N_8726,N_7612,N_7894);
xnor U8727 (N_8727,N_7954,N_7514);
xnor U8728 (N_8728,N_7544,N_7453);
xor U8729 (N_8729,N_7424,N_7682);
and U8730 (N_8730,N_7851,N_7870);
or U8731 (N_8731,N_7834,N_7235);
nor U8732 (N_8732,N_7953,N_7216);
and U8733 (N_8733,N_7081,N_7918);
nor U8734 (N_8734,N_7413,N_7852);
or U8735 (N_8735,N_7322,N_7407);
nor U8736 (N_8736,N_7305,N_7961);
nand U8737 (N_8737,N_7406,N_7143);
xor U8738 (N_8738,N_7684,N_7364);
nor U8739 (N_8739,N_7575,N_7665);
or U8740 (N_8740,N_7473,N_7480);
nand U8741 (N_8741,N_7874,N_7027);
nand U8742 (N_8742,N_7640,N_7722);
nor U8743 (N_8743,N_7235,N_7901);
nand U8744 (N_8744,N_7402,N_7970);
or U8745 (N_8745,N_7603,N_7107);
nor U8746 (N_8746,N_7299,N_7141);
nand U8747 (N_8747,N_7765,N_7491);
nor U8748 (N_8748,N_7278,N_7384);
or U8749 (N_8749,N_7483,N_7442);
xnor U8750 (N_8750,N_7436,N_7375);
xor U8751 (N_8751,N_7515,N_7268);
xor U8752 (N_8752,N_7321,N_7141);
nand U8753 (N_8753,N_7376,N_7917);
and U8754 (N_8754,N_7216,N_7957);
xnor U8755 (N_8755,N_7371,N_7444);
and U8756 (N_8756,N_7623,N_7124);
or U8757 (N_8757,N_7603,N_7954);
nor U8758 (N_8758,N_7991,N_7312);
nand U8759 (N_8759,N_7639,N_7522);
and U8760 (N_8760,N_7947,N_7181);
xnor U8761 (N_8761,N_7237,N_7633);
or U8762 (N_8762,N_7217,N_7258);
or U8763 (N_8763,N_7579,N_7241);
nor U8764 (N_8764,N_7339,N_7272);
nand U8765 (N_8765,N_7679,N_7002);
or U8766 (N_8766,N_7382,N_7218);
nor U8767 (N_8767,N_7195,N_7851);
nor U8768 (N_8768,N_7144,N_7060);
xor U8769 (N_8769,N_7217,N_7037);
and U8770 (N_8770,N_7250,N_7133);
nand U8771 (N_8771,N_7784,N_7519);
xnor U8772 (N_8772,N_7423,N_7400);
or U8773 (N_8773,N_7565,N_7809);
or U8774 (N_8774,N_7833,N_7814);
or U8775 (N_8775,N_7639,N_7167);
and U8776 (N_8776,N_7728,N_7729);
or U8777 (N_8777,N_7856,N_7924);
xnor U8778 (N_8778,N_7458,N_7175);
xor U8779 (N_8779,N_7489,N_7840);
nand U8780 (N_8780,N_7310,N_7271);
or U8781 (N_8781,N_7553,N_7691);
nor U8782 (N_8782,N_7166,N_7898);
xor U8783 (N_8783,N_7546,N_7766);
xor U8784 (N_8784,N_7980,N_7652);
or U8785 (N_8785,N_7944,N_7930);
nor U8786 (N_8786,N_7554,N_7535);
or U8787 (N_8787,N_7742,N_7698);
or U8788 (N_8788,N_7274,N_7672);
nor U8789 (N_8789,N_7682,N_7634);
and U8790 (N_8790,N_7961,N_7329);
nand U8791 (N_8791,N_7051,N_7084);
nand U8792 (N_8792,N_7634,N_7994);
and U8793 (N_8793,N_7760,N_7859);
or U8794 (N_8794,N_7825,N_7509);
nor U8795 (N_8795,N_7877,N_7907);
nor U8796 (N_8796,N_7983,N_7032);
and U8797 (N_8797,N_7130,N_7643);
xor U8798 (N_8798,N_7626,N_7221);
or U8799 (N_8799,N_7508,N_7970);
xor U8800 (N_8800,N_7049,N_7019);
xnor U8801 (N_8801,N_7095,N_7497);
and U8802 (N_8802,N_7508,N_7941);
xnor U8803 (N_8803,N_7840,N_7253);
xor U8804 (N_8804,N_7455,N_7253);
nor U8805 (N_8805,N_7829,N_7671);
and U8806 (N_8806,N_7702,N_7986);
nor U8807 (N_8807,N_7372,N_7751);
nor U8808 (N_8808,N_7753,N_7885);
or U8809 (N_8809,N_7081,N_7134);
nand U8810 (N_8810,N_7761,N_7026);
xnor U8811 (N_8811,N_7170,N_7245);
xor U8812 (N_8812,N_7766,N_7314);
nand U8813 (N_8813,N_7267,N_7866);
xor U8814 (N_8814,N_7907,N_7306);
nand U8815 (N_8815,N_7331,N_7781);
or U8816 (N_8816,N_7111,N_7174);
nand U8817 (N_8817,N_7892,N_7010);
nor U8818 (N_8818,N_7157,N_7124);
xnor U8819 (N_8819,N_7642,N_7907);
xnor U8820 (N_8820,N_7877,N_7701);
and U8821 (N_8821,N_7991,N_7517);
xnor U8822 (N_8822,N_7796,N_7178);
nor U8823 (N_8823,N_7374,N_7746);
and U8824 (N_8824,N_7299,N_7807);
nand U8825 (N_8825,N_7999,N_7267);
xnor U8826 (N_8826,N_7803,N_7076);
or U8827 (N_8827,N_7616,N_7797);
or U8828 (N_8828,N_7539,N_7346);
xnor U8829 (N_8829,N_7632,N_7777);
nor U8830 (N_8830,N_7389,N_7364);
nand U8831 (N_8831,N_7624,N_7216);
and U8832 (N_8832,N_7858,N_7375);
xor U8833 (N_8833,N_7486,N_7939);
or U8834 (N_8834,N_7759,N_7519);
nand U8835 (N_8835,N_7894,N_7877);
and U8836 (N_8836,N_7667,N_7502);
or U8837 (N_8837,N_7771,N_7966);
and U8838 (N_8838,N_7719,N_7672);
nand U8839 (N_8839,N_7750,N_7523);
xnor U8840 (N_8840,N_7992,N_7347);
xnor U8841 (N_8841,N_7048,N_7128);
and U8842 (N_8842,N_7105,N_7491);
nor U8843 (N_8843,N_7538,N_7585);
xor U8844 (N_8844,N_7062,N_7787);
xnor U8845 (N_8845,N_7061,N_7631);
nand U8846 (N_8846,N_7753,N_7821);
nor U8847 (N_8847,N_7277,N_7872);
or U8848 (N_8848,N_7399,N_7340);
or U8849 (N_8849,N_7745,N_7893);
xor U8850 (N_8850,N_7649,N_7598);
nand U8851 (N_8851,N_7077,N_7756);
xor U8852 (N_8852,N_7522,N_7497);
or U8853 (N_8853,N_7482,N_7201);
and U8854 (N_8854,N_7570,N_7807);
xnor U8855 (N_8855,N_7886,N_7024);
or U8856 (N_8856,N_7544,N_7500);
xnor U8857 (N_8857,N_7421,N_7715);
or U8858 (N_8858,N_7666,N_7452);
and U8859 (N_8859,N_7658,N_7477);
or U8860 (N_8860,N_7718,N_7523);
nor U8861 (N_8861,N_7192,N_7518);
or U8862 (N_8862,N_7943,N_7157);
nand U8863 (N_8863,N_7237,N_7919);
nor U8864 (N_8864,N_7673,N_7918);
and U8865 (N_8865,N_7380,N_7999);
nand U8866 (N_8866,N_7764,N_7611);
nand U8867 (N_8867,N_7424,N_7885);
and U8868 (N_8868,N_7196,N_7408);
or U8869 (N_8869,N_7447,N_7543);
or U8870 (N_8870,N_7076,N_7492);
xor U8871 (N_8871,N_7903,N_7297);
nand U8872 (N_8872,N_7650,N_7291);
and U8873 (N_8873,N_7050,N_7189);
xor U8874 (N_8874,N_7274,N_7181);
nor U8875 (N_8875,N_7425,N_7661);
nor U8876 (N_8876,N_7158,N_7312);
nor U8877 (N_8877,N_7501,N_7911);
nor U8878 (N_8878,N_7152,N_7753);
nand U8879 (N_8879,N_7653,N_7332);
and U8880 (N_8880,N_7181,N_7890);
and U8881 (N_8881,N_7250,N_7420);
or U8882 (N_8882,N_7531,N_7368);
xor U8883 (N_8883,N_7139,N_7690);
or U8884 (N_8884,N_7317,N_7440);
and U8885 (N_8885,N_7931,N_7554);
xor U8886 (N_8886,N_7052,N_7590);
and U8887 (N_8887,N_7827,N_7210);
and U8888 (N_8888,N_7570,N_7589);
and U8889 (N_8889,N_7206,N_7332);
or U8890 (N_8890,N_7781,N_7684);
and U8891 (N_8891,N_7821,N_7163);
nor U8892 (N_8892,N_7105,N_7953);
and U8893 (N_8893,N_7641,N_7168);
nand U8894 (N_8894,N_7061,N_7066);
nand U8895 (N_8895,N_7539,N_7138);
nand U8896 (N_8896,N_7675,N_7293);
xnor U8897 (N_8897,N_7499,N_7161);
or U8898 (N_8898,N_7896,N_7410);
nor U8899 (N_8899,N_7700,N_7627);
nand U8900 (N_8900,N_7066,N_7184);
and U8901 (N_8901,N_7018,N_7063);
nand U8902 (N_8902,N_7632,N_7687);
and U8903 (N_8903,N_7638,N_7275);
and U8904 (N_8904,N_7756,N_7730);
nand U8905 (N_8905,N_7947,N_7835);
nor U8906 (N_8906,N_7571,N_7136);
xnor U8907 (N_8907,N_7926,N_7513);
and U8908 (N_8908,N_7385,N_7626);
and U8909 (N_8909,N_7177,N_7881);
xnor U8910 (N_8910,N_7334,N_7519);
or U8911 (N_8911,N_7478,N_7703);
xnor U8912 (N_8912,N_7013,N_7162);
nor U8913 (N_8913,N_7665,N_7397);
or U8914 (N_8914,N_7760,N_7328);
nand U8915 (N_8915,N_7560,N_7762);
and U8916 (N_8916,N_7590,N_7988);
nor U8917 (N_8917,N_7843,N_7585);
xnor U8918 (N_8918,N_7064,N_7562);
nor U8919 (N_8919,N_7739,N_7331);
xor U8920 (N_8920,N_7216,N_7929);
or U8921 (N_8921,N_7818,N_7775);
or U8922 (N_8922,N_7841,N_7941);
nand U8923 (N_8923,N_7684,N_7220);
or U8924 (N_8924,N_7257,N_7184);
nand U8925 (N_8925,N_7412,N_7522);
nor U8926 (N_8926,N_7142,N_7115);
nand U8927 (N_8927,N_7726,N_7616);
or U8928 (N_8928,N_7599,N_7090);
xnor U8929 (N_8929,N_7449,N_7800);
xnor U8930 (N_8930,N_7860,N_7117);
nor U8931 (N_8931,N_7415,N_7421);
nand U8932 (N_8932,N_7441,N_7795);
nand U8933 (N_8933,N_7452,N_7868);
and U8934 (N_8934,N_7931,N_7012);
and U8935 (N_8935,N_7638,N_7876);
or U8936 (N_8936,N_7533,N_7140);
xor U8937 (N_8937,N_7312,N_7934);
or U8938 (N_8938,N_7438,N_7050);
xor U8939 (N_8939,N_7439,N_7314);
or U8940 (N_8940,N_7098,N_7193);
nand U8941 (N_8941,N_7218,N_7719);
nand U8942 (N_8942,N_7513,N_7851);
or U8943 (N_8943,N_7237,N_7976);
nand U8944 (N_8944,N_7524,N_7065);
nor U8945 (N_8945,N_7077,N_7698);
xor U8946 (N_8946,N_7333,N_7143);
nand U8947 (N_8947,N_7552,N_7245);
nor U8948 (N_8948,N_7654,N_7578);
nand U8949 (N_8949,N_7501,N_7726);
nor U8950 (N_8950,N_7813,N_7536);
xor U8951 (N_8951,N_7724,N_7869);
nand U8952 (N_8952,N_7715,N_7106);
nand U8953 (N_8953,N_7027,N_7293);
or U8954 (N_8954,N_7140,N_7327);
nand U8955 (N_8955,N_7988,N_7438);
and U8956 (N_8956,N_7642,N_7563);
and U8957 (N_8957,N_7841,N_7171);
nand U8958 (N_8958,N_7525,N_7864);
nand U8959 (N_8959,N_7909,N_7167);
or U8960 (N_8960,N_7073,N_7229);
nand U8961 (N_8961,N_7206,N_7718);
xnor U8962 (N_8962,N_7935,N_7513);
nand U8963 (N_8963,N_7304,N_7734);
or U8964 (N_8964,N_7493,N_7655);
and U8965 (N_8965,N_7467,N_7741);
and U8966 (N_8966,N_7474,N_7342);
nor U8967 (N_8967,N_7776,N_7753);
nand U8968 (N_8968,N_7389,N_7910);
nor U8969 (N_8969,N_7978,N_7222);
nor U8970 (N_8970,N_7015,N_7373);
nand U8971 (N_8971,N_7575,N_7361);
or U8972 (N_8972,N_7893,N_7662);
and U8973 (N_8973,N_7952,N_7791);
nor U8974 (N_8974,N_7543,N_7220);
xnor U8975 (N_8975,N_7169,N_7186);
nand U8976 (N_8976,N_7572,N_7011);
or U8977 (N_8977,N_7391,N_7316);
nor U8978 (N_8978,N_7225,N_7410);
nand U8979 (N_8979,N_7968,N_7201);
or U8980 (N_8980,N_7878,N_7989);
or U8981 (N_8981,N_7065,N_7619);
nor U8982 (N_8982,N_7538,N_7151);
xor U8983 (N_8983,N_7125,N_7258);
or U8984 (N_8984,N_7193,N_7117);
and U8985 (N_8985,N_7029,N_7323);
nand U8986 (N_8986,N_7166,N_7569);
xor U8987 (N_8987,N_7031,N_7589);
nor U8988 (N_8988,N_7414,N_7765);
nand U8989 (N_8989,N_7994,N_7905);
nand U8990 (N_8990,N_7989,N_7863);
nand U8991 (N_8991,N_7353,N_7037);
nand U8992 (N_8992,N_7737,N_7250);
and U8993 (N_8993,N_7011,N_7990);
xnor U8994 (N_8994,N_7353,N_7256);
nor U8995 (N_8995,N_7774,N_7143);
nand U8996 (N_8996,N_7584,N_7314);
or U8997 (N_8997,N_7976,N_7919);
or U8998 (N_8998,N_7553,N_7031);
xor U8999 (N_8999,N_7496,N_7118);
and U9000 (N_9000,N_8833,N_8681);
nor U9001 (N_9001,N_8530,N_8045);
nor U9002 (N_9002,N_8840,N_8892);
and U9003 (N_9003,N_8515,N_8697);
xor U9004 (N_9004,N_8660,N_8082);
nand U9005 (N_9005,N_8032,N_8704);
and U9006 (N_9006,N_8441,N_8602);
xor U9007 (N_9007,N_8277,N_8972);
nor U9008 (N_9008,N_8226,N_8984);
nor U9009 (N_9009,N_8264,N_8190);
or U9010 (N_9010,N_8887,N_8049);
or U9011 (N_9011,N_8363,N_8422);
nand U9012 (N_9012,N_8985,N_8702);
xor U9013 (N_9013,N_8987,N_8313);
and U9014 (N_9014,N_8338,N_8362);
and U9015 (N_9015,N_8506,N_8736);
nand U9016 (N_9016,N_8797,N_8755);
xor U9017 (N_9017,N_8393,N_8137);
nand U9018 (N_9018,N_8883,N_8298);
nand U9019 (N_9019,N_8759,N_8606);
and U9020 (N_9020,N_8412,N_8579);
nand U9021 (N_9021,N_8209,N_8097);
and U9022 (N_9022,N_8541,N_8815);
or U9023 (N_9023,N_8976,N_8726);
and U9024 (N_9024,N_8882,N_8732);
and U9025 (N_9025,N_8600,N_8935);
nor U9026 (N_9026,N_8677,N_8199);
or U9027 (N_9027,N_8015,N_8193);
and U9028 (N_9028,N_8788,N_8671);
and U9029 (N_9029,N_8295,N_8496);
nor U9030 (N_9030,N_8562,N_8713);
or U9031 (N_9031,N_8122,N_8529);
nand U9032 (N_9032,N_8867,N_8091);
or U9033 (N_9033,N_8477,N_8276);
or U9034 (N_9034,N_8372,N_8737);
xor U9035 (N_9035,N_8652,N_8722);
xnor U9036 (N_9036,N_8498,N_8554);
nand U9037 (N_9037,N_8905,N_8907);
or U9038 (N_9038,N_8084,N_8922);
and U9039 (N_9039,N_8013,N_8921);
nand U9040 (N_9040,N_8436,N_8272);
or U9041 (N_9041,N_8842,N_8399);
or U9042 (N_9042,N_8818,N_8410);
xor U9043 (N_9043,N_8880,N_8253);
nor U9044 (N_9044,N_8381,N_8742);
nand U9045 (N_9045,N_8693,N_8782);
xor U9046 (N_9046,N_8760,N_8349);
or U9047 (N_9047,N_8160,N_8252);
nand U9048 (N_9048,N_8262,N_8731);
xnor U9049 (N_9049,N_8587,N_8631);
or U9050 (N_9050,N_8617,N_8542);
xnor U9051 (N_9051,N_8208,N_8945);
xor U9052 (N_9052,N_8392,N_8510);
nor U9053 (N_9053,N_8949,N_8453);
and U9054 (N_9054,N_8689,N_8911);
xor U9055 (N_9055,N_8041,N_8430);
xnor U9056 (N_9056,N_8405,N_8023);
xnor U9057 (N_9057,N_8933,N_8938);
nand U9058 (N_9058,N_8896,N_8991);
nand U9059 (N_9059,N_8189,N_8786);
or U9060 (N_9060,N_8157,N_8281);
or U9061 (N_9061,N_8472,N_8042);
and U9062 (N_9062,N_8730,N_8953);
or U9063 (N_9063,N_8265,N_8240);
and U9064 (N_9064,N_8112,N_8879);
and U9065 (N_9065,N_8361,N_8803);
nand U9066 (N_9066,N_8549,N_8270);
nor U9067 (N_9067,N_8229,N_8802);
nand U9068 (N_9068,N_8563,N_8378);
or U9069 (N_9069,N_8512,N_8877);
and U9070 (N_9070,N_8709,N_8646);
nand U9071 (N_9071,N_8806,N_8201);
nor U9072 (N_9072,N_8126,N_8343);
nand U9073 (N_9073,N_8968,N_8364);
nand U9074 (N_9074,N_8409,N_8897);
nand U9075 (N_9075,N_8464,N_8275);
or U9076 (N_9076,N_8036,N_8345);
nand U9077 (N_9077,N_8799,N_8993);
nor U9078 (N_9078,N_8375,N_8571);
nand U9079 (N_9079,N_8639,N_8889);
nand U9080 (N_9080,N_8576,N_8304);
or U9081 (N_9081,N_8266,N_8981);
and U9082 (N_9082,N_8168,N_8028);
nor U9083 (N_9083,N_8152,N_8535);
xnor U9084 (N_9084,N_8117,N_8656);
and U9085 (N_9085,N_8242,N_8643);
nand U9086 (N_9086,N_8902,N_8147);
nor U9087 (N_9087,N_8075,N_8948);
nand U9088 (N_9088,N_8508,N_8793);
nor U9089 (N_9089,N_8690,N_8664);
and U9090 (N_9090,N_8320,N_8163);
nor U9091 (N_9091,N_8403,N_8068);
and U9092 (N_9092,N_8961,N_8413);
nor U9093 (N_9093,N_8143,N_8169);
xnor U9094 (N_9094,N_8145,N_8936);
or U9095 (N_9095,N_8300,N_8625);
nor U9096 (N_9096,N_8521,N_8951);
nand U9097 (N_9097,N_8531,N_8784);
nor U9098 (N_9098,N_8359,N_8288);
and U9099 (N_9099,N_8177,N_8448);
or U9100 (N_9100,N_8766,N_8780);
nand U9101 (N_9101,N_8107,N_8575);
and U9102 (N_9102,N_8460,N_8994);
nor U9103 (N_9103,N_8250,N_8449);
xnor U9104 (N_9104,N_8663,N_8826);
xor U9105 (N_9105,N_8629,N_8746);
or U9106 (N_9106,N_8257,N_8156);
nand U9107 (N_9107,N_8578,N_8283);
or U9108 (N_9108,N_8493,N_8988);
and U9109 (N_9109,N_8110,N_8100);
xnor U9110 (N_9110,N_8206,N_8094);
and U9111 (N_9111,N_8970,N_8928);
nand U9112 (N_9112,N_8260,N_8678);
nand U9113 (N_9113,N_8241,N_8178);
nand U9114 (N_9114,N_8052,N_8767);
xor U9115 (N_9115,N_8705,N_8341);
or U9116 (N_9116,N_8481,N_8164);
or U9117 (N_9117,N_8333,N_8081);
xnor U9118 (N_9118,N_8166,N_8955);
and U9119 (N_9119,N_8845,N_8106);
and U9120 (N_9120,N_8354,N_8995);
and U9121 (N_9121,N_8202,N_8593);
or U9122 (N_9122,N_8975,N_8719);
xor U9123 (N_9123,N_8329,N_8317);
nor U9124 (N_9124,N_8556,N_8454);
xor U9125 (N_9125,N_8829,N_8572);
nand U9126 (N_9126,N_8609,N_8616);
or U9127 (N_9127,N_8757,N_8424);
and U9128 (N_9128,N_8798,N_8247);
or U9129 (N_9129,N_8673,N_8532);
xnor U9130 (N_9130,N_8822,N_8694);
and U9131 (N_9131,N_8305,N_8044);
xor U9132 (N_9132,N_8219,N_8764);
nor U9133 (N_9133,N_8603,N_8059);
or U9134 (N_9134,N_8624,N_8374);
nor U9135 (N_9135,N_8326,N_8947);
nor U9136 (N_9136,N_8109,N_8781);
nor U9137 (N_9137,N_8849,N_8058);
xor U9138 (N_9138,N_8330,N_8514);
and U9139 (N_9139,N_8886,N_8591);
nand U9140 (N_9140,N_8926,N_8653);
nor U9141 (N_9141,N_8239,N_8765);
or U9142 (N_9142,N_8325,N_8724);
nand U9143 (N_9143,N_8334,N_8710);
nor U9144 (N_9144,N_8864,N_8520);
or U9145 (N_9145,N_8397,N_8810);
xnor U9146 (N_9146,N_8061,N_8561);
or U9147 (N_9147,N_8350,N_8367);
nor U9148 (N_9148,N_8387,N_8821);
or U9149 (N_9149,N_8509,N_8093);
nor U9150 (N_9150,N_8158,N_8855);
xnor U9151 (N_9151,N_8973,N_8550);
xor U9152 (N_9152,N_8963,N_8000);
xor U9153 (N_9153,N_8830,N_8360);
nand U9154 (N_9154,N_8753,N_8811);
nand U9155 (N_9155,N_8628,N_8835);
nand U9156 (N_9156,N_8194,N_8141);
nand U9157 (N_9157,N_8473,N_8480);
or U9158 (N_9158,N_8876,N_8407);
nand U9159 (N_9159,N_8284,N_8125);
and U9160 (N_9160,N_8303,N_8621);
and U9161 (N_9161,N_8517,N_8170);
nor U9162 (N_9162,N_8688,N_8212);
and U9163 (N_9163,N_8470,N_8528);
or U9164 (N_9164,N_8459,N_8129);
xor U9165 (N_9165,N_8642,N_8006);
xnor U9166 (N_9166,N_8640,N_8683);
xor U9167 (N_9167,N_8008,N_8072);
and U9168 (N_9168,N_8466,N_8336);
nor U9169 (N_9169,N_8992,N_8200);
xor U9170 (N_9170,N_8622,N_8670);
or U9171 (N_9171,N_8136,N_8069);
nand U9172 (N_9172,N_8655,N_8964);
nand U9173 (N_9173,N_8699,N_8998);
nand U9174 (N_9174,N_8487,N_8831);
xor U9175 (N_9175,N_8862,N_8455);
nor U9176 (N_9176,N_8382,N_8256);
xor U9177 (N_9177,N_8001,N_8733);
and U9178 (N_9178,N_8172,N_8539);
nand U9179 (N_9179,N_8501,N_8982);
xor U9180 (N_9180,N_8344,N_8744);
or U9181 (N_9181,N_8618,N_8014);
xnor U9182 (N_9182,N_8115,N_8033);
nor U9183 (N_9183,N_8930,N_8183);
and U9184 (N_9184,N_8931,N_8144);
nor U9185 (N_9185,N_8977,N_8940);
or U9186 (N_9186,N_8773,N_8997);
xor U9187 (N_9187,N_8890,N_8401);
nand U9188 (N_9188,N_8686,N_8127);
nor U9189 (N_9189,N_8598,N_8148);
and U9190 (N_9190,N_8159,N_8500);
or U9191 (N_9191,N_8687,N_8268);
nor U9192 (N_9192,N_8118,N_8066);
and U9193 (N_9193,N_8906,N_8874);
nor U9194 (N_9194,N_8021,N_8012);
and U9195 (N_9195,N_8577,N_8919);
and U9196 (N_9196,N_8296,N_8195);
nor U9197 (N_9197,N_8096,N_8866);
or U9198 (N_9198,N_8682,N_8340);
xnor U9199 (N_9199,N_8511,N_8259);
and U9200 (N_9200,N_8776,N_8064);
or U9201 (N_9201,N_8099,N_8221);
nand U9202 (N_9202,N_8747,N_8016);
nor U9203 (N_9203,N_8708,N_8139);
or U9204 (N_9204,N_8488,N_8020);
or U9205 (N_9205,N_8585,N_8130);
nor U9206 (N_9206,N_8279,N_8769);
and U9207 (N_9207,N_8071,N_8654);
nor U9208 (N_9208,N_8944,N_8037);
or U9209 (N_9209,N_8030,N_8476);
nor U9210 (N_9210,N_8743,N_8565);
nand U9211 (N_9211,N_8167,N_8232);
xor U9212 (N_9212,N_8376,N_8318);
or U9213 (N_9213,N_8513,N_8003);
or U9214 (N_9214,N_8437,N_8969);
xnor U9215 (N_9215,N_8456,N_8319);
nor U9216 (N_9216,N_8134,N_8471);
or U9217 (N_9217,N_8146,N_8089);
or U9218 (N_9218,N_8322,N_8584);
and U9219 (N_9219,N_8452,N_8294);
nor U9220 (N_9220,N_8872,N_8370);
xnor U9221 (N_9221,N_8280,N_8820);
xor U9222 (N_9222,N_8235,N_8536);
xor U9223 (N_9223,N_8952,N_8924);
nand U9224 (N_9224,N_8943,N_8289);
nand U9225 (N_9225,N_8551,N_8038);
nand U9226 (N_9226,N_8601,N_8332);
xnor U9227 (N_9227,N_8123,N_8179);
xor U9228 (N_9228,N_8827,N_8675);
or U9229 (N_9229,N_8445,N_8132);
or U9230 (N_9230,N_8558,N_8077);
or U9231 (N_9231,N_8626,N_8234);
or U9232 (N_9232,N_8852,N_8634);
and U9233 (N_9233,N_8668,N_8315);
or U9234 (N_9234,N_8751,N_8365);
nor U9235 (N_9235,N_8429,N_8915);
and U9236 (N_9236,N_8224,N_8142);
nand U9237 (N_9237,N_8173,N_8790);
nand U9238 (N_9238,N_8898,N_8323);
nor U9239 (N_9239,N_8222,N_8216);
and U9240 (N_9240,N_8237,N_8560);
or U9241 (N_9241,N_8328,N_8053);
nor U9242 (N_9242,N_8181,N_8062);
or U9243 (N_9243,N_8929,N_8856);
and U9244 (N_9244,N_8665,N_8098);
xnor U9245 (N_9245,N_8388,N_8779);
xor U9246 (N_9246,N_8717,N_8807);
and U9247 (N_9247,N_8958,N_8611);
and U9248 (N_9248,N_8727,N_8908);
and U9249 (N_9249,N_8217,N_8153);
and U9250 (N_9250,N_8980,N_8899);
nor U9251 (N_9251,N_8808,N_8461);
xnor U9252 (N_9252,N_8809,N_8468);
xnor U9253 (N_9253,N_8331,N_8772);
nand U9254 (N_9254,N_8116,N_8881);
nor U9255 (N_9255,N_8739,N_8519);
nor U9256 (N_9256,N_8884,N_8352);
or U9257 (N_9257,N_8901,N_8419);
or U9258 (N_9258,N_8114,N_8762);
xnor U9259 (N_9259,N_8478,N_8925);
nor U9260 (N_9260,N_8150,N_8078);
and U9261 (N_9261,N_8805,N_8604);
and U9262 (N_9262,N_8228,N_8394);
nor U9263 (N_9263,N_8076,N_8040);
xor U9264 (N_9264,N_8548,N_8567);
xor U9265 (N_9265,N_8457,N_8785);
and U9266 (N_9266,N_8770,N_8269);
or U9267 (N_9267,N_8108,N_8263);
or U9268 (N_9268,N_8192,N_8384);
and U9269 (N_9269,N_8927,N_8599);
xor U9270 (N_9270,N_8986,N_8771);
nand U9271 (N_9271,N_8442,N_8421);
xor U9272 (N_9272,N_8543,N_8246);
nand U9273 (N_9273,N_8650,N_8916);
and U9274 (N_9274,N_8087,N_8768);
or U9275 (N_9275,N_8574,N_8836);
nand U9276 (N_9276,N_8745,N_8486);
nand U9277 (N_9277,N_8171,N_8346);
xor U9278 (N_9278,N_8996,N_8339);
and U9279 (N_9279,N_8377,N_8215);
or U9280 (N_9280,N_8051,N_8111);
and U9281 (N_9281,N_8503,N_8698);
or U9282 (N_9282,N_8103,N_8067);
xor U9283 (N_9283,N_8337,N_8187);
and U9284 (N_9284,N_8850,N_8989);
and U9285 (N_9285,N_8716,N_8026);
nor U9286 (N_9286,N_8754,N_8285);
xnor U9287 (N_9287,N_8391,N_8588);
xnor U9288 (N_9288,N_8004,N_8474);
nor U9289 (N_9289,N_8400,N_8395);
nand U9290 (N_9290,N_8196,N_8527);
and U9291 (N_9291,N_8233,N_8796);
xor U9292 (N_9292,N_8297,N_8443);
nor U9293 (N_9293,N_8633,N_8151);
nor U9294 (N_9294,N_8635,N_8846);
xnor U9295 (N_9295,N_8853,N_8065);
xor U9296 (N_9296,N_8203,N_8282);
xor U9297 (N_9297,N_8957,N_8795);
and U9298 (N_9298,N_8789,N_8865);
nand U9299 (N_9299,N_8290,N_8937);
nand U9300 (N_9300,N_8761,N_8465);
nand U9301 (N_9301,N_8416,N_8007);
or U9302 (N_9302,N_8718,N_8844);
xnor U9303 (N_9303,N_8910,N_8031);
or U9304 (N_9304,N_8659,N_8133);
nor U9305 (N_9305,N_8404,N_8914);
or U9306 (N_9306,N_8131,N_8418);
nand U9307 (N_9307,N_8458,N_8197);
xnor U9308 (N_9308,N_8524,N_8291);
and U9309 (N_9309,N_8475,N_8244);
nand U9310 (N_9310,N_8425,N_8909);
and U9311 (N_9311,N_8715,N_8778);
and U9312 (N_9312,N_8314,N_8703);
nor U9313 (N_9313,N_8662,N_8869);
xor U9314 (N_9314,N_8590,N_8547);
nand U9315 (N_9315,N_8396,N_8763);
or U9316 (N_9316,N_8046,N_8965);
xor U9317 (N_9317,N_8706,N_8707);
nor U9318 (N_9318,N_8469,N_8612);
xnor U9319 (N_9319,N_8861,N_8615);
or U9320 (N_9320,N_8095,N_8522);
nor U9321 (N_9321,N_8439,N_8586);
or U9322 (N_9322,N_8573,N_8946);
xnor U9323 (N_9323,N_8557,N_8932);
nor U9324 (N_9324,N_8959,N_8566);
nor U9325 (N_9325,N_8823,N_8638);
nor U9326 (N_9326,N_8005,N_8149);
xnor U9327 (N_9327,N_8495,N_8274);
nand U9328 (N_9328,N_8525,N_8316);
and U9329 (N_9329,N_8348,N_8605);
or U9330 (N_9330,N_8950,N_8630);
or U9331 (N_9331,N_8243,N_8592);
nor U9332 (N_9332,N_8154,N_8426);
or U9333 (N_9333,N_8175,N_8301);
nand U9334 (N_9334,N_8775,N_8278);
and U9335 (N_9335,N_8939,N_8685);
and U9336 (N_9336,N_8523,N_8819);
or U9337 (N_9337,N_8983,N_8534);
nor U9338 (N_9338,N_8356,N_8714);
or U9339 (N_9339,N_8581,N_8614);
and U9340 (N_9340,N_8433,N_8482);
or U9341 (N_9341,N_8728,N_8934);
xnor U9342 (N_9342,N_8923,N_8540);
or U9343 (N_9343,N_8312,N_8182);
nor U9344 (N_9344,N_8119,N_8018);
or U9345 (N_9345,N_8729,N_8701);
xnor U9346 (N_9346,N_8255,N_8641);
nand U9347 (N_9347,N_8351,N_8875);
nand U9348 (N_9348,N_8494,N_8451);
nand U9349 (N_9349,N_8999,N_8083);
nand U9350 (N_9350,N_8787,N_8057);
nor U9351 (N_9351,N_8386,N_8841);
and U9352 (N_9352,N_8347,N_8804);
and U9353 (N_9353,N_8185,N_8894);
and U9354 (N_9354,N_8636,N_8074);
nor U9355 (N_9355,N_8735,N_8680);
nand U9356 (N_9356,N_8105,N_8415);
or U9357 (N_9357,N_8555,N_8627);
and U9358 (N_9358,N_8124,N_8251);
nor U9359 (N_9359,N_8832,N_8582);
nand U9360 (N_9360,N_8029,N_8676);
and U9361 (N_9361,N_8080,N_8311);
xor U9362 (N_9362,N_8792,N_8838);
nor U9363 (N_9363,N_8186,N_8446);
nor U9364 (N_9364,N_8960,N_8647);
nand U9365 (N_9365,N_8380,N_8917);
or U9366 (N_9366,N_8794,N_8408);
xor U9367 (N_9367,N_8249,N_8878);
nor U9368 (N_9368,N_8580,N_8489);
and U9369 (N_9369,N_8204,N_8596);
nor U9370 (N_9370,N_8054,N_8389);
and U9371 (N_9371,N_8533,N_8813);
xor U9372 (N_9372,N_8692,N_8414);
xnor U9373 (N_9373,N_8043,N_8390);
xnor U9374 (N_9374,N_8245,N_8438);
xnor U9375 (N_9375,N_8696,N_8073);
xor U9376 (N_9376,N_8321,N_8420);
nor U9377 (N_9377,N_8490,N_8649);
and U9378 (N_9378,N_8700,N_8752);
or U9379 (N_9379,N_8213,N_8583);
or U9380 (N_9380,N_8373,N_8750);
and U9381 (N_9381,N_8034,N_8292);
and U9382 (N_9382,N_8858,N_8814);
nand U9383 (N_9383,N_8967,N_8777);
xnor U9384 (N_9384,N_8904,N_8411);
and U9385 (N_9385,N_8507,N_8025);
nor U9386 (N_9386,N_8086,N_8227);
and U9387 (N_9387,N_8545,N_8379);
nand U9388 (N_9388,N_8056,N_8637);
and U9389 (N_9389,N_8230,N_8113);
or U9390 (N_9390,N_8758,N_8783);
and U9391 (N_9391,N_8431,N_8258);
and U9392 (N_9392,N_8667,N_8353);
nand U9393 (N_9393,N_8368,N_8238);
xnor U9394 (N_9394,N_8888,N_8335);
xnor U9395 (N_9395,N_8847,N_8463);
nand U9396 (N_9396,N_8302,N_8559);
nand U9397 (N_9397,N_8214,N_8851);
and U9398 (N_9398,N_8155,N_8165);
nor U9399 (N_9399,N_8942,N_8128);
nor U9400 (N_9400,N_8800,N_8047);
and U9401 (N_9401,N_8293,N_8138);
and U9402 (N_9402,N_8564,N_8218);
nand U9403 (N_9403,N_8299,N_8104);
and U9404 (N_9404,N_8063,N_8011);
nor U9405 (N_9405,N_8254,N_8684);
nor U9406 (N_9406,N_8121,N_8184);
and U9407 (N_9407,N_8979,N_8544);
nand U9408 (N_9408,N_8553,N_8180);
or U9409 (N_9409,N_8484,N_8920);
and U9410 (N_9410,N_8161,N_8774);
or U9411 (N_9411,N_8589,N_8843);
xnor U9412 (N_9412,N_8479,N_8220);
nor U9413 (N_9413,N_8824,N_8306);
nor U9414 (N_9414,N_8483,N_8672);
nand U9415 (N_9415,N_8309,N_8900);
and U9416 (N_9416,N_8248,N_8594);
and U9417 (N_9417,N_8691,N_8516);
and U9418 (N_9418,N_8492,N_8749);
or U9419 (N_9419,N_8427,N_8010);
nand U9420 (N_9420,N_8538,N_8828);
and U9421 (N_9421,N_8913,N_8552);
or U9422 (N_9422,N_8027,N_8679);
nor U9423 (N_9423,N_8060,N_8623);
nor U9424 (N_9424,N_8491,N_8055);
and U9425 (N_9425,N_8140,N_8398);
or U9426 (N_9426,N_8120,N_8723);
xnor U9427 (N_9427,N_8569,N_8286);
and U9428 (N_9428,N_8791,N_8342);
nand U9429 (N_9429,N_8327,N_8962);
nor U9430 (N_9430,N_8499,N_8085);
xor U9431 (N_9431,N_8974,N_8871);
nand U9432 (N_9432,N_8174,N_8868);
xor U9433 (N_9433,N_8870,N_8432);
nand U9434 (N_9434,N_8941,N_8608);
and U9435 (N_9435,N_8570,N_8848);
and U9436 (N_9436,N_8504,N_8050);
or U9437 (N_9437,N_8893,N_8261);
nor U9438 (N_9438,N_8462,N_8497);
and U9439 (N_9439,N_8756,N_8669);
xor U9440 (N_9440,N_8834,N_8417);
xor U9441 (N_9441,N_8817,N_8912);
and U9442 (N_9442,N_8816,N_8954);
and U9443 (N_9443,N_8207,N_8369);
and U9444 (N_9444,N_8537,N_8371);
xor U9445 (N_9445,N_8019,N_8444);
and U9446 (N_9446,N_8366,N_8644);
nor U9447 (N_9447,N_8017,N_8648);
nor U9448 (N_9448,N_8518,N_8009);
and U9449 (N_9449,N_8423,N_8188);
and U9450 (N_9450,N_8839,N_8825);
or U9451 (N_9451,N_8674,N_8505);
xnor U9452 (N_9452,N_8355,N_8024);
nor U9453 (N_9453,N_8310,N_8070);
or U9454 (N_9454,N_8734,N_8918);
nor U9455 (N_9455,N_8002,N_8287);
and U9456 (N_9456,N_8198,N_8191);
xor U9457 (N_9457,N_8854,N_8210);
nand U9458 (N_9458,N_8966,N_8610);
and U9459 (N_9459,N_8385,N_8860);
or U9460 (N_9460,N_8978,N_8748);
or U9461 (N_9461,N_8837,N_8712);
and U9462 (N_9462,N_8440,N_8307);
nor U9463 (N_9463,N_8225,N_8273);
nand U9464 (N_9464,N_8236,N_8324);
xor U9465 (N_9465,N_8595,N_8135);
nand U9466 (N_9466,N_8092,N_8101);
nand U9467 (N_9467,N_8205,N_8738);
nor U9468 (N_9468,N_8903,N_8613);
and U9469 (N_9469,N_8741,N_8720);
nand U9470 (N_9470,N_8231,N_8695);
or U9471 (N_9471,N_8873,N_8450);
and U9472 (N_9472,N_8176,N_8485);
and U9473 (N_9473,N_8632,N_8568);
and U9474 (N_9474,N_8645,N_8863);
xnor U9475 (N_9475,N_8526,N_8428);
xor U9476 (N_9476,N_8022,N_8039);
nand U9477 (N_9477,N_8090,N_8435);
nand U9478 (N_9478,N_8035,N_8651);
xor U9479 (N_9479,N_8308,N_8502);
nor U9480 (N_9480,N_8721,N_8358);
xor U9481 (N_9481,N_8857,N_8383);
and U9482 (N_9482,N_8725,N_8162);
nand U9483 (N_9483,N_8546,N_8402);
or U9484 (N_9484,N_8079,N_8447);
or U9485 (N_9485,N_8088,N_8971);
xnor U9486 (N_9486,N_8891,N_8619);
or U9487 (N_9487,N_8223,N_8956);
or U9488 (N_9488,N_8711,N_8434);
nand U9489 (N_9489,N_8658,N_8801);
nor U9490 (N_9490,N_8467,N_8267);
or U9491 (N_9491,N_8885,N_8661);
nor U9492 (N_9492,N_8357,N_8048);
nand U9493 (N_9493,N_8657,N_8597);
xor U9494 (N_9494,N_8895,N_8990);
nand U9495 (N_9495,N_8740,N_8859);
or U9496 (N_9496,N_8607,N_8620);
xnor U9497 (N_9497,N_8812,N_8211);
nor U9498 (N_9498,N_8406,N_8102);
nor U9499 (N_9499,N_8666,N_8271);
or U9500 (N_9500,N_8271,N_8160);
and U9501 (N_9501,N_8596,N_8804);
and U9502 (N_9502,N_8109,N_8775);
xor U9503 (N_9503,N_8872,N_8659);
nor U9504 (N_9504,N_8528,N_8832);
and U9505 (N_9505,N_8539,N_8960);
or U9506 (N_9506,N_8026,N_8771);
or U9507 (N_9507,N_8192,N_8832);
nand U9508 (N_9508,N_8543,N_8467);
or U9509 (N_9509,N_8342,N_8626);
or U9510 (N_9510,N_8529,N_8744);
and U9511 (N_9511,N_8934,N_8420);
or U9512 (N_9512,N_8630,N_8188);
nand U9513 (N_9513,N_8783,N_8965);
or U9514 (N_9514,N_8527,N_8458);
nor U9515 (N_9515,N_8479,N_8961);
or U9516 (N_9516,N_8384,N_8681);
and U9517 (N_9517,N_8212,N_8075);
nor U9518 (N_9518,N_8089,N_8135);
nor U9519 (N_9519,N_8304,N_8277);
nor U9520 (N_9520,N_8823,N_8663);
nor U9521 (N_9521,N_8509,N_8281);
and U9522 (N_9522,N_8809,N_8635);
nor U9523 (N_9523,N_8907,N_8692);
nand U9524 (N_9524,N_8104,N_8623);
or U9525 (N_9525,N_8246,N_8134);
nor U9526 (N_9526,N_8914,N_8411);
and U9527 (N_9527,N_8578,N_8349);
nand U9528 (N_9528,N_8191,N_8987);
nand U9529 (N_9529,N_8638,N_8886);
and U9530 (N_9530,N_8196,N_8192);
xnor U9531 (N_9531,N_8750,N_8855);
nand U9532 (N_9532,N_8763,N_8245);
or U9533 (N_9533,N_8057,N_8437);
nand U9534 (N_9534,N_8601,N_8357);
nand U9535 (N_9535,N_8003,N_8402);
nor U9536 (N_9536,N_8390,N_8355);
and U9537 (N_9537,N_8980,N_8979);
xor U9538 (N_9538,N_8698,N_8010);
xnor U9539 (N_9539,N_8093,N_8655);
xor U9540 (N_9540,N_8028,N_8540);
nand U9541 (N_9541,N_8324,N_8106);
nand U9542 (N_9542,N_8936,N_8807);
xnor U9543 (N_9543,N_8628,N_8553);
nor U9544 (N_9544,N_8145,N_8581);
and U9545 (N_9545,N_8088,N_8499);
xnor U9546 (N_9546,N_8854,N_8466);
or U9547 (N_9547,N_8450,N_8400);
nor U9548 (N_9548,N_8234,N_8897);
or U9549 (N_9549,N_8522,N_8931);
xor U9550 (N_9550,N_8432,N_8489);
nor U9551 (N_9551,N_8207,N_8330);
nor U9552 (N_9552,N_8116,N_8335);
nor U9553 (N_9553,N_8445,N_8919);
and U9554 (N_9554,N_8292,N_8498);
nor U9555 (N_9555,N_8423,N_8432);
and U9556 (N_9556,N_8315,N_8082);
nor U9557 (N_9557,N_8879,N_8794);
nand U9558 (N_9558,N_8275,N_8716);
xnor U9559 (N_9559,N_8005,N_8735);
nor U9560 (N_9560,N_8021,N_8576);
nor U9561 (N_9561,N_8733,N_8134);
or U9562 (N_9562,N_8322,N_8912);
nand U9563 (N_9563,N_8149,N_8626);
nand U9564 (N_9564,N_8155,N_8731);
or U9565 (N_9565,N_8735,N_8625);
and U9566 (N_9566,N_8688,N_8936);
nor U9567 (N_9567,N_8026,N_8013);
or U9568 (N_9568,N_8121,N_8865);
nand U9569 (N_9569,N_8725,N_8503);
and U9570 (N_9570,N_8923,N_8692);
nor U9571 (N_9571,N_8935,N_8293);
or U9572 (N_9572,N_8800,N_8020);
or U9573 (N_9573,N_8955,N_8547);
nor U9574 (N_9574,N_8058,N_8286);
and U9575 (N_9575,N_8426,N_8121);
xnor U9576 (N_9576,N_8371,N_8260);
or U9577 (N_9577,N_8083,N_8050);
xnor U9578 (N_9578,N_8301,N_8108);
and U9579 (N_9579,N_8511,N_8155);
xor U9580 (N_9580,N_8967,N_8571);
nand U9581 (N_9581,N_8163,N_8129);
or U9582 (N_9582,N_8156,N_8728);
nand U9583 (N_9583,N_8598,N_8063);
and U9584 (N_9584,N_8910,N_8208);
xnor U9585 (N_9585,N_8301,N_8718);
xor U9586 (N_9586,N_8302,N_8491);
nor U9587 (N_9587,N_8828,N_8384);
or U9588 (N_9588,N_8051,N_8651);
nor U9589 (N_9589,N_8942,N_8295);
nor U9590 (N_9590,N_8203,N_8288);
nor U9591 (N_9591,N_8887,N_8255);
nor U9592 (N_9592,N_8376,N_8597);
and U9593 (N_9593,N_8932,N_8773);
nand U9594 (N_9594,N_8166,N_8757);
nand U9595 (N_9595,N_8382,N_8329);
nand U9596 (N_9596,N_8349,N_8362);
and U9597 (N_9597,N_8050,N_8806);
xnor U9598 (N_9598,N_8657,N_8492);
nand U9599 (N_9599,N_8859,N_8394);
nand U9600 (N_9600,N_8613,N_8971);
and U9601 (N_9601,N_8777,N_8457);
or U9602 (N_9602,N_8060,N_8114);
and U9603 (N_9603,N_8808,N_8402);
nor U9604 (N_9604,N_8088,N_8575);
xor U9605 (N_9605,N_8564,N_8802);
or U9606 (N_9606,N_8520,N_8242);
or U9607 (N_9607,N_8640,N_8003);
nand U9608 (N_9608,N_8414,N_8608);
xnor U9609 (N_9609,N_8229,N_8556);
nor U9610 (N_9610,N_8321,N_8486);
nand U9611 (N_9611,N_8099,N_8844);
and U9612 (N_9612,N_8950,N_8890);
and U9613 (N_9613,N_8537,N_8348);
or U9614 (N_9614,N_8115,N_8082);
nor U9615 (N_9615,N_8981,N_8825);
xor U9616 (N_9616,N_8364,N_8651);
xor U9617 (N_9617,N_8091,N_8587);
xnor U9618 (N_9618,N_8065,N_8681);
nor U9619 (N_9619,N_8638,N_8509);
or U9620 (N_9620,N_8316,N_8820);
xnor U9621 (N_9621,N_8061,N_8321);
nor U9622 (N_9622,N_8012,N_8631);
or U9623 (N_9623,N_8084,N_8904);
nor U9624 (N_9624,N_8288,N_8061);
or U9625 (N_9625,N_8555,N_8149);
and U9626 (N_9626,N_8619,N_8426);
or U9627 (N_9627,N_8251,N_8346);
xnor U9628 (N_9628,N_8920,N_8520);
xor U9629 (N_9629,N_8186,N_8586);
or U9630 (N_9630,N_8606,N_8291);
xor U9631 (N_9631,N_8521,N_8015);
nor U9632 (N_9632,N_8586,N_8163);
or U9633 (N_9633,N_8486,N_8202);
and U9634 (N_9634,N_8340,N_8325);
or U9635 (N_9635,N_8292,N_8751);
xor U9636 (N_9636,N_8516,N_8393);
xnor U9637 (N_9637,N_8361,N_8122);
nor U9638 (N_9638,N_8667,N_8165);
and U9639 (N_9639,N_8003,N_8976);
or U9640 (N_9640,N_8996,N_8774);
xnor U9641 (N_9641,N_8331,N_8998);
or U9642 (N_9642,N_8223,N_8944);
and U9643 (N_9643,N_8875,N_8091);
nor U9644 (N_9644,N_8227,N_8956);
nor U9645 (N_9645,N_8591,N_8267);
xor U9646 (N_9646,N_8293,N_8783);
nor U9647 (N_9647,N_8473,N_8505);
and U9648 (N_9648,N_8738,N_8286);
nor U9649 (N_9649,N_8542,N_8525);
nand U9650 (N_9650,N_8213,N_8386);
and U9651 (N_9651,N_8651,N_8228);
xor U9652 (N_9652,N_8277,N_8276);
and U9653 (N_9653,N_8954,N_8755);
nand U9654 (N_9654,N_8845,N_8189);
nor U9655 (N_9655,N_8640,N_8002);
and U9656 (N_9656,N_8001,N_8886);
xnor U9657 (N_9657,N_8999,N_8924);
or U9658 (N_9658,N_8922,N_8490);
xor U9659 (N_9659,N_8948,N_8201);
or U9660 (N_9660,N_8647,N_8226);
nor U9661 (N_9661,N_8368,N_8104);
nor U9662 (N_9662,N_8272,N_8937);
nor U9663 (N_9663,N_8017,N_8251);
nor U9664 (N_9664,N_8466,N_8038);
and U9665 (N_9665,N_8692,N_8514);
or U9666 (N_9666,N_8739,N_8121);
xor U9667 (N_9667,N_8735,N_8538);
nor U9668 (N_9668,N_8448,N_8517);
nand U9669 (N_9669,N_8240,N_8808);
nor U9670 (N_9670,N_8534,N_8374);
or U9671 (N_9671,N_8504,N_8410);
xor U9672 (N_9672,N_8230,N_8133);
nor U9673 (N_9673,N_8628,N_8013);
xnor U9674 (N_9674,N_8776,N_8083);
nor U9675 (N_9675,N_8242,N_8458);
nand U9676 (N_9676,N_8143,N_8276);
xor U9677 (N_9677,N_8961,N_8755);
and U9678 (N_9678,N_8275,N_8119);
nor U9679 (N_9679,N_8576,N_8213);
or U9680 (N_9680,N_8158,N_8086);
nor U9681 (N_9681,N_8286,N_8607);
nor U9682 (N_9682,N_8226,N_8372);
xnor U9683 (N_9683,N_8777,N_8308);
and U9684 (N_9684,N_8703,N_8655);
nand U9685 (N_9685,N_8766,N_8059);
and U9686 (N_9686,N_8836,N_8616);
or U9687 (N_9687,N_8316,N_8636);
nand U9688 (N_9688,N_8886,N_8348);
nor U9689 (N_9689,N_8677,N_8905);
xnor U9690 (N_9690,N_8183,N_8544);
and U9691 (N_9691,N_8266,N_8972);
nand U9692 (N_9692,N_8529,N_8397);
nor U9693 (N_9693,N_8930,N_8970);
nand U9694 (N_9694,N_8384,N_8703);
nand U9695 (N_9695,N_8389,N_8639);
or U9696 (N_9696,N_8670,N_8747);
nor U9697 (N_9697,N_8086,N_8108);
nand U9698 (N_9698,N_8261,N_8770);
xor U9699 (N_9699,N_8136,N_8197);
or U9700 (N_9700,N_8110,N_8960);
nor U9701 (N_9701,N_8679,N_8548);
nand U9702 (N_9702,N_8309,N_8474);
or U9703 (N_9703,N_8014,N_8630);
nand U9704 (N_9704,N_8888,N_8245);
and U9705 (N_9705,N_8658,N_8864);
and U9706 (N_9706,N_8008,N_8942);
and U9707 (N_9707,N_8117,N_8795);
xor U9708 (N_9708,N_8774,N_8642);
nor U9709 (N_9709,N_8152,N_8081);
nand U9710 (N_9710,N_8025,N_8048);
and U9711 (N_9711,N_8147,N_8806);
or U9712 (N_9712,N_8025,N_8042);
or U9713 (N_9713,N_8250,N_8458);
or U9714 (N_9714,N_8799,N_8952);
and U9715 (N_9715,N_8232,N_8494);
and U9716 (N_9716,N_8246,N_8113);
and U9717 (N_9717,N_8317,N_8682);
xnor U9718 (N_9718,N_8203,N_8999);
or U9719 (N_9719,N_8838,N_8868);
nand U9720 (N_9720,N_8677,N_8949);
nand U9721 (N_9721,N_8989,N_8219);
and U9722 (N_9722,N_8596,N_8926);
or U9723 (N_9723,N_8628,N_8631);
and U9724 (N_9724,N_8578,N_8866);
nor U9725 (N_9725,N_8930,N_8921);
nand U9726 (N_9726,N_8499,N_8026);
xnor U9727 (N_9727,N_8856,N_8397);
nor U9728 (N_9728,N_8834,N_8074);
nor U9729 (N_9729,N_8772,N_8640);
xnor U9730 (N_9730,N_8317,N_8871);
or U9731 (N_9731,N_8941,N_8119);
or U9732 (N_9732,N_8922,N_8742);
or U9733 (N_9733,N_8379,N_8371);
and U9734 (N_9734,N_8579,N_8912);
or U9735 (N_9735,N_8264,N_8589);
nor U9736 (N_9736,N_8903,N_8394);
and U9737 (N_9737,N_8187,N_8459);
or U9738 (N_9738,N_8265,N_8713);
or U9739 (N_9739,N_8149,N_8365);
and U9740 (N_9740,N_8049,N_8928);
nand U9741 (N_9741,N_8406,N_8314);
xor U9742 (N_9742,N_8800,N_8009);
nor U9743 (N_9743,N_8481,N_8839);
or U9744 (N_9744,N_8722,N_8864);
nor U9745 (N_9745,N_8835,N_8698);
nor U9746 (N_9746,N_8857,N_8585);
and U9747 (N_9747,N_8168,N_8304);
nor U9748 (N_9748,N_8459,N_8282);
xnor U9749 (N_9749,N_8127,N_8544);
and U9750 (N_9750,N_8713,N_8110);
nor U9751 (N_9751,N_8222,N_8711);
and U9752 (N_9752,N_8079,N_8243);
and U9753 (N_9753,N_8861,N_8455);
nand U9754 (N_9754,N_8569,N_8430);
nor U9755 (N_9755,N_8790,N_8004);
nor U9756 (N_9756,N_8145,N_8493);
nor U9757 (N_9757,N_8997,N_8583);
xor U9758 (N_9758,N_8049,N_8573);
nand U9759 (N_9759,N_8380,N_8265);
nor U9760 (N_9760,N_8772,N_8275);
or U9761 (N_9761,N_8372,N_8279);
and U9762 (N_9762,N_8615,N_8246);
or U9763 (N_9763,N_8323,N_8952);
and U9764 (N_9764,N_8624,N_8931);
nor U9765 (N_9765,N_8469,N_8961);
and U9766 (N_9766,N_8471,N_8454);
or U9767 (N_9767,N_8496,N_8807);
nor U9768 (N_9768,N_8824,N_8361);
or U9769 (N_9769,N_8125,N_8408);
or U9770 (N_9770,N_8799,N_8806);
xor U9771 (N_9771,N_8367,N_8978);
nor U9772 (N_9772,N_8935,N_8652);
and U9773 (N_9773,N_8966,N_8103);
or U9774 (N_9774,N_8972,N_8921);
or U9775 (N_9775,N_8164,N_8767);
nor U9776 (N_9776,N_8840,N_8930);
xor U9777 (N_9777,N_8667,N_8047);
and U9778 (N_9778,N_8245,N_8323);
or U9779 (N_9779,N_8668,N_8508);
and U9780 (N_9780,N_8343,N_8564);
xor U9781 (N_9781,N_8389,N_8076);
nand U9782 (N_9782,N_8827,N_8330);
xor U9783 (N_9783,N_8946,N_8732);
nor U9784 (N_9784,N_8425,N_8874);
nor U9785 (N_9785,N_8395,N_8045);
and U9786 (N_9786,N_8116,N_8599);
and U9787 (N_9787,N_8690,N_8138);
nor U9788 (N_9788,N_8642,N_8287);
nand U9789 (N_9789,N_8993,N_8135);
or U9790 (N_9790,N_8755,N_8131);
xor U9791 (N_9791,N_8938,N_8529);
nand U9792 (N_9792,N_8215,N_8567);
and U9793 (N_9793,N_8384,N_8841);
and U9794 (N_9794,N_8665,N_8039);
nand U9795 (N_9795,N_8762,N_8053);
or U9796 (N_9796,N_8978,N_8361);
nor U9797 (N_9797,N_8859,N_8928);
nand U9798 (N_9798,N_8298,N_8760);
and U9799 (N_9799,N_8732,N_8316);
nand U9800 (N_9800,N_8552,N_8824);
and U9801 (N_9801,N_8538,N_8680);
nand U9802 (N_9802,N_8577,N_8431);
and U9803 (N_9803,N_8860,N_8405);
or U9804 (N_9804,N_8093,N_8822);
and U9805 (N_9805,N_8366,N_8038);
or U9806 (N_9806,N_8835,N_8022);
or U9807 (N_9807,N_8455,N_8741);
nand U9808 (N_9808,N_8653,N_8220);
or U9809 (N_9809,N_8235,N_8445);
nand U9810 (N_9810,N_8161,N_8325);
and U9811 (N_9811,N_8563,N_8100);
xnor U9812 (N_9812,N_8088,N_8137);
nand U9813 (N_9813,N_8414,N_8510);
and U9814 (N_9814,N_8184,N_8475);
and U9815 (N_9815,N_8009,N_8027);
nand U9816 (N_9816,N_8126,N_8778);
xnor U9817 (N_9817,N_8436,N_8239);
xnor U9818 (N_9818,N_8442,N_8130);
nand U9819 (N_9819,N_8116,N_8361);
nand U9820 (N_9820,N_8763,N_8357);
nor U9821 (N_9821,N_8605,N_8238);
nand U9822 (N_9822,N_8921,N_8344);
xor U9823 (N_9823,N_8088,N_8918);
nor U9824 (N_9824,N_8895,N_8072);
nor U9825 (N_9825,N_8497,N_8921);
or U9826 (N_9826,N_8986,N_8890);
and U9827 (N_9827,N_8153,N_8091);
and U9828 (N_9828,N_8654,N_8285);
nor U9829 (N_9829,N_8743,N_8726);
or U9830 (N_9830,N_8584,N_8881);
xnor U9831 (N_9831,N_8031,N_8859);
xor U9832 (N_9832,N_8298,N_8258);
or U9833 (N_9833,N_8671,N_8632);
and U9834 (N_9834,N_8438,N_8935);
xor U9835 (N_9835,N_8844,N_8048);
or U9836 (N_9836,N_8195,N_8702);
or U9837 (N_9837,N_8903,N_8759);
xnor U9838 (N_9838,N_8634,N_8892);
xor U9839 (N_9839,N_8877,N_8875);
and U9840 (N_9840,N_8791,N_8693);
nor U9841 (N_9841,N_8932,N_8098);
nand U9842 (N_9842,N_8048,N_8591);
nand U9843 (N_9843,N_8275,N_8857);
xor U9844 (N_9844,N_8472,N_8861);
xor U9845 (N_9845,N_8713,N_8611);
xnor U9846 (N_9846,N_8643,N_8782);
xnor U9847 (N_9847,N_8821,N_8612);
xnor U9848 (N_9848,N_8539,N_8493);
nor U9849 (N_9849,N_8219,N_8402);
or U9850 (N_9850,N_8490,N_8324);
nand U9851 (N_9851,N_8088,N_8514);
nand U9852 (N_9852,N_8445,N_8454);
xor U9853 (N_9853,N_8005,N_8547);
nor U9854 (N_9854,N_8002,N_8911);
nor U9855 (N_9855,N_8017,N_8959);
nor U9856 (N_9856,N_8731,N_8957);
or U9857 (N_9857,N_8973,N_8874);
nand U9858 (N_9858,N_8905,N_8837);
xor U9859 (N_9859,N_8536,N_8058);
or U9860 (N_9860,N_8510,N_8788);
nand U9861 (N_9861,N_8186,N_8094);
or U9862 (N_9862,N_8497,N_8495);
xnor U9863 (N_9863,N_8299,N_8155);
and U9864 (N_9864,N_8187,N_8405);
nor U9865 (N_9865,N_8460,N_8759);
or U9866 (N_9866,N_8550,N_8820);
nand U9867 (N_9867,N_8665,N_8791);
nand U9868 (N_9868,N_8971,N_8412);
or U9869 (N_9869,N_8055,N_8761);
nand U9870 (N_9870,N_8470,N_8477);
nor U9871 (N_9871,N_8779,N_8879);
nor U9872 (N_9872,N_8561,N_8386);
or U9873 (N_9873,N_8412,N_8021);
xnor U9874 (N_9874,N_8331,N_8594);
or U9875 (N_9875,N_8849,N_8421);
nor U9876 (N_9876,N_8144,N_8636);
nand U9877 (N_9877,N_8008,N_8631);
nand U9878 (N_9878,N_8346,N_8841);
nor U9879 (N_9879,N_8184,N_8478);
nand U9880 (N_9880,N_8429,N_8652);
or U9881 (N_9881,N_8595,N_8296);
nor U9882 (N_9882,N_8183,N_8224);
or U9883 (N_9883,N_8655,N_8321);
nand U9884 (N_9884,N_8439,N_8517);
xnor U9885 (N_9885,N_8240,N_8506);
and U9886 (N_9886,N_8420,N_8345);
or U9887 (N_9887,N_8056,N_8505);
or U9888 (N_9888,N_8538,N_8196);
nor U9889 (N_9889,N_8280,N_8255);
xnor U9890 (N_9890,N_8922,N_8776);
and U9891 (N_9891,N_8315,N_8313);
xor U9892 (N_9892,N_8969,N_8508);
or U9893 (N_9893,N_8143,N_8769);
nor U9894 (N_9894,N_8380,N_8272);
or U9895 (N_9895,N_8114,N_8184);
and U9896 (N_9896,N_8404,N_8603);
nor U9897 (N_9897,N_8627,N_8116);
xor U9898 (N_9898,N_8308,N_8930);
and U9899 (N_9899,N_8307,N_8825);
xnor U9900 (N_9900,N_8591,N_8524);
xnor U9901 (N_9901,N_8700,N_8932);
and U9902 (N_9902,N_8335,N_8407);
nand U9903 (N_9903,N_8280,N_8325);
or U9904 (N_9904,N_8627,N_8977);
xor U9905 (N_9905,N_8905,N_8299);
and U9906 (N_9906,N_8802,N_8817);
and U9907 (N_9907,N_8159,N_8552);
nand U9908 (N_9908,N_8751,N_8431);
nor U9909 (N_9909,N_8451,N_8434);
or U9910 (N_9910,N_8656,N_8581);
xor U9911 (N_9911,N_8239,N_8749);
xnor U9912 (N_9912,N_8952,N_8750);
nor U9913 (N_9913,N_8586,N_8164);
and U9914 (N_9914,N_8074,N_8445);
and U9915 (N_9915,N_8194,N_8265);
nand U9916 (N_9916,N_8069,N_8666);
xor U9917 (N_9917,N_8421,N_8477);
nand U9918 (N_9918,N_8265,N_8322);
nor U9919 (N_9919,N_8285,N_8898);
nand U9920 (N_9920,N_8946,N_8652);
xor U9921 (N_9921,N_8191,N_8299);
nand U9922 (N_9922,N_8073,N_8422);
nand U9923 (N_9923,N_8736,N_8256);
and U9924 (N_9924,N_8046,N_8511);
xor U9925 (N_9925,N_8957,N_8017);
xnor U9926 (N_9926,N_8802,N_8562);
or U9927 (N_9927,N_8392,N_8167);
or U9928 (N_9928,N_8109,N_8560);
and U9929 (N_9929,N_8030,N_8118);
or U9930 (N_9930,N_8260,N_8288);
nor U9931 (N_9931,N_8684,N_8901);
nor U9932 (N_9932,N_8022,N_8495);
xor U9933 (N_9933,N_8547,N_8137);
xor U9934 (N_9934,N_8927,N_8798);
nand U9935 (N_9935,N_8674,N_8797);
nand U9936 (N_9936,N_8818,N_8639);
or U9937 (N_9937,N_8225,N_8870);
or U9938 (N_9938,N_8419,N_8489);
xor U9939 (N_9939,N_8688,N_8488);
xnor U9940 (N_9940,N_8876,N_8509);
and U9941 (N_9941,N_8088,N_8793);
or U9942 (N_9942,N_8933,N_8110);
and U9943 (N_9943,N_8826,N_8063);
nand U9944 (N_9944,N_8749,N_8500);
or U9945 (N_9945,N_8954,N_8398);
or U9946 (N_9946,N_8641,N_8224);
nor U9947 (N_9947,N_8628,N_8185);
or U9948 (N_9948,N_8652,N_8368);
or U9949 (N_9949,N_8996,N_8582);
xnor U9950 (N_9950,N_8429,N_8402);
and U9951 (N_9951,N_8180,N_8774);
nand U9952 (N_9952,N_8066,N_8353);
nand U9953 (N_9953,N_8574,N_8356);
or U9954 (N_9954,N_8318,N_8445);
xnor U9955 (N_9955,N_8746,N_8681);
xor U9956 (N_9956,N_8524,N_8700);
xnor U9957 (N_9957,N_8935,N_8723);
nand U9958 (N_9958,N_8632,N_8504);
xor U9959 (N_9959,N_8048,N_8730);
nor U9960 (N_9960,N_8517,N_8312);
nand U9961 (N_9961,N_8052,N_8223);
or U9962 (N_9962,N_8111,N_8739);
and U9963 (N_9963,N_8348,N_8060);
or U9964 (N_9964,N_8781,N_8972);
and U9965 (N_9965,N_8903,N_8571);
xnor U9966 (N_9966,N_8740,N_8621);
xnor U9967 (N_9967,N_8734,N_8503);
nor U9968 (N_9968,N_8070,N_8602);
xnor U9969 (N_9969,N_8855,N_8422);
or U9970 (N_9970,N_8961,N_8594);
and U9971 (N_9971,N_8282,N_8743);
xor U9972 (N_9972,N_8669,N_8134);
nor U9973 (N_9973,N_8419,N_8067);
xnor U9974 (N_9974,N_8466,N_8707);
and U9975 (N_9975,N_8009,N_8103);
or U9976 (N_9976,N_8727,N_8713);
nand U9977 (N_9977,N_8598,N_8139);
nor U9978 (N_9978,N_8810,N_8308);
and U9979 (N_9979,N_8262,N_8847);
or U9980 (N_9980,N_8068,N_8595);
nor U9981 (N_9981,N_8891,N_8309);
nand U9982 (N_9982,N_8513,N_8505);
xnor U9983 (N_9983,N_8056,N_8974);
or U9984 (N_9984,N_8268,N_8409);
nor U9985 (N_9985,N_8926,N_8801);
and U9986 (N_9986,N_8580,N_8300);
xnor U9987 (N_9987,N_8864,N_8088);
nand U9988 (N_9988,N_8613,N_8304);
xnor U9989 (N_9989,N_8836,N_8048);
nand U9990 (N_9990,N_8858,N_8714);
xor U9991 (N_9991,N_8757,N_8315);
xnor U9992 (N_9992,N_8873,N_8944);
nor U9993 (N_9993,N_8173,N_8112);
or U9994 (N_9994,N_8339,N_8134);
and U9995 (N_9995,N_8409,N_8130);
nand U9996 (N_9996,N_8405,N_8989);
and U9997 (N_9997,N_8596,N_8393);
nor U9998 (N_9998,N_8226,N_8218);
and U9999 (N_9999,N_8767,N_8369);
xor U10000 (N_10000,N_9032,N_9215);
xnor U10001 (N_10001,N_9216,N_9457);
and U10002 (N_10002,N_9637,N_9534);
and U10003 (N_10003,N_9532,N_9268);
and U10004 (N_10004,N_9141,N_9337);
and U10005 (N_10005,N_9370,N_9230);
or U10006 (N_10006,N_9279,N_9171);
nor U10007 (N_10007,N_9820,N_9316);
and U10008 (N_10008,N_9516,N_9306);
xor U10009 (N_10009,N_9679,N_9517);
nand U10010 (N_10010,N_9162,N_9385);
or U10011 (N_10011,N_9739,N_9664);
or U10012 (N_10012,N_9289,N_9156);
or U10013 (N_10013,N_9830,N_9834);
nor U10014 (N_10014,N_9020,N_9527);
xor U10015 (N_10015,N_9789,N_9418);
nand U10016 (N_10016,N_9214,N_9336);
and U10017 (N_10017,N_9544,N_9762);
nor U10018 (N_10018,N_9083,N_9939);
nand U10019 (N_10019,N_9573,N_9660);
nor U10020 (N_10020,N_9266,N_9646);
nand U10021 (N_10021,N_9930,N_9982);
or U10022 (N_10022,N_9650,N_9080);
xnor U10023 (N_10023,N_9062,N_9643);
xor U10024 (N_10024,N_9591,N_9614);
nand U10025 (N_10025,N_9757,N_9455);
or U10026 (N_10026,N_9831,N_9025);
and U10027 (N_10027,N_9477,N_9656);
nor U10028 (N_10028,N_9277,N_9489);
and U10029 (N_10029,N_9961,N_9072);
nor U10030 (N_10030,N_9284,N_9401);
or U10031 (N_10031,N_9040,N_9099);
or U10032 (N_10032,N_9552,N_9641);
or U10033 (N_10033,N_9872,N_9602);
xor U10034 (N_10034,N_9240,N_9364);
or U10035 (N_10035,N_9628,N_9124);
nand U10036 (N_10036,N_9330,N_9157);
nor U10037 (N_10037,N_9061,N_9115);
nor U10038 (N_10038,N_9521,N_9538);
and U10039 (N_10039,N_9129,N_9706);
nand U10040 (N_10040,N_9004,N_9555);
nand U10041 (N_10041,N_9949,N_9966);
nor U10042 (N_10042,N_9823,N_9466);
or U10043 (N_10043,N_9267,N_9593);
and U10044 (N_10044,N_9726,N_9222);
or U10045 (N_10045,N_9674,N_9146);
nand U10046 (N_10046,N_9168,N_9339);
xor U10047 (N_10047,N_9935,N_9498);
xnor U10048 (N_10048,N_9962,N_9741);
nor U10049 (N_10049,N_9116,N_9662);
nor U10050 (N_10050,N_9753,N_9668);
xor U10051 (N_10051,N_9568,N_9916);
xnor U10052 (N_10052,N_9788,N_9848);
xor U10053 (N_10053,N_9967,N_9703);
and U10054 (N_10054,N_9533,N_9066);
xnor U10055 (N_10055,N_9127,N_9299);
nor U10056 (N_10056,N_9079,N_9950);
nand U10057 (N_10057,N_9545,N_9885);
or U10058 (N_10058,N_9531,N_9041);
xor U10059 (N_10059,N_9122,N_9599);
and U10060 (N_10060,N_9791,N_9426);
and U10061 (N_10061,N_9526,N_9852);
xnor U10062 (N_10062,N_9932,N_9611);
and U10063 (N_10063,N_9743,N_9972);
and U10064 (N_10064,N_9399,N_9409);
nand U10065 (N_10065,N_9981,N_9003);
and U10066 (N_10066,N_9839,N_9778);
xor U10067 (N_10067,N_9153,N_9280);
nand U10068 (N_10068,N_9394,N_9528);
or U10069 (N_10069,N_9014,N_9001);
or U10070 (N_10070,N_9348,N_9262);
nand U10071 (N_10071,N_9236,N_9804);
xor U10072 (N_10072,N_9749,N_9325);
or U10073 (N_10073,N_9414,N_9824);
nor U10074 (N_10074,N_9524,N_9459);
xnor U10075 (N_10075,N_9577,N_9057);
nand U10076 (N_10076,N_9803,N_9888);
nor U10077 (N_10077,N_9717,N_9081);
xnor U10078 (N_10078,N_9082,N_9601);
nor U10079 (N_10079,N_9630,N_9217);
nand U10080 (N_10080,N_9442,N_9805);
or U10081 (N_10081,N_9126,N_9386);
nand U10082 (N_10082,N_9507,N_9673);
and U10083 (N_10083,N_9011,N_9798);
and U10084 (N_10084,N_9147,N_9863);
nand U10085 (N_10085,N_9782,N_9451);
and U10086 (N_10086,N_9965,N_9075);
nor U10087 (N_10087,N_9607,N_9996);
or U10088 (N_10088,N_9049,N_9000);
and U10089 (N_10089,N_9756,N_9449);
nor U10090 (N_10090,N_9632,N_9132);
nor U10091 (N_10091,N_9832,N_9374);
nand U10092 (N_10092,N_9270,N_9106);
and U10093 (N_10093,N_9197,N_9248);
nand U10094 (N_10094,N_9200,N_9810);
nor U10095 (N_10095,N_9702,N_9826);
and U10096 (N_10096,N_9427,N_9887);
nand U10097 (N_10097,N_9100,N_9398);
nor U10098 (N_10098,N_9112,N_9143);
xor U10099 (N_10099,N_9604,N_9360);
or U10100 (N_10100,N_9612,N_9154);
nand U10101 (N_10101,N_9121,N_9670);
and U10102 (N_10102,N_9219,N_9669);
and U10103 (N_10103,N_9358,N_9985);
xnor U10104 (N_10104,N_9192,N_9086);
nor U10105 (N_10105,N_9909,N_9898);
and U10106 (N_10106,N_9058,N_9980);
nor U10107 (N_10107,N_9689,N_9039);
and U10108 (N_10108,N_9535,N_9028);
xor U10109 (N_10109,N_9381,N_9616);
xnor U10110 (N_10110,N_9755,N_9857);
nor U10111 (N_10111,N_9968,N_9429);
nor U10112 (N_10112,N_9787,N_9882);
or U10113 (N_10113,N_9415,N_9210);
xor U10114 (N_10114,N_9999,N_9559);
xor U10115 (N_10115,N_9110,N_9130);
and U10116 (N_10116,N_9549,N_9505);
nand U10117 (N_10117,N_9204,N_9391);
or U10118 (N_10118,N_9992,N_9564);
or U10119 (N_10119,N_9237,N_9140);
nand U10120 (N_10120,N_9149,N_9499);
and U10121 (N_10121,N_9472,N_9492);
or U10122 (N_10122,N_9111,N_9686);
nand U10123 (N_10123,N_9844,N_9977);
or U10124 (N_10124,N_9841,N_9301);
xnor U10125 (N_10125,N_9493,N_9366);
or U10126 (N_10126,N_9987,N_9379);
and U10127 (N_10127,N_9367,N_9257);
xor U10128 (N_10128,N_9822,N_9501);
xnor U10129 (N_10129,N_9194,N_9595);
and U10130 (N_10130,N_9006,N_9241);
xor U10131 (N_10131,N_9677,N_9118);
nor U10132 (N_10132,N_9588,N_9312);
xor U10133 (N_10133,N_9922,N_9634);
nor U10134 (N_10134,N_9550,N_9658);
nand U10135 (N_10135,N_9676,N_9748);
and U10136 (N_10136,N_9021,N_9818);
or U10137 (N_10137,N_9690,N_9940);
nand U10138 (N_10138,N_9167,N_9902);
or U10139 (N_10139,N_9036,N_9211);
or U10140 (N_10140,N_9581,N_9085);
or U10141 (N_10141,N_9542,N_9186);
or U10142 (N_10142,N_9671,N_9059);
xnor U10143 (N_10143,N_9800,N_9586);
nor U10144 (N_10144,N_9605,N_9024);
nor U10145 (N_10145,N_9868,N_9113);
or U10146 (N_10146,N_9736,N_9187);
nand U10147 (N_10147,N_9227,N_9433);
nand U10148 (N_10148,N_9343,N_9395);
or U10149 (N_10149,N_9165,N_9189);
nand U10150 (N_10150,N_9462,N_9907);
or U10151 (N_10151,N_9514,N_9447);
nor U10152 (N_10152,N_9443,N_9687);
nor U10153 (N_10153,N_9205,N_9889);
xnor U10154 (N_10154,N_9575,N_9722);
nand U10155 (N_10155,N_9948,N_9983);
nor U10156 (N_10156,N_9963,N_9023);
or U10157 (N_10157,N_9496,N_9582);
nor U10158 (N_10158,N_9056,N_9864);
nor U10159 (N_10159,N_9239,N_9037);
or U10160 (N_10160,N_9362,N_9213);
xor U10161 (N_10161,N_9208,N_9342);
nor U10162 (N_10162,N_9875,N_9619);
xor U10163 (N_10163,N_9812,N_9334);
xnor U10164 (N_10164,N_9639,N_9264);
or U10165 (N_10165,N_9302,N_9294);
or U10166 (N_10166,N_9710,N_9566);
or U10167 (N_10167,N_9708,N_9245);
or U10168 (N_10168,N_9166,N_9318);
and U10169 (N_10169,N_9022,N_9924);
or U10170 (N_10170,N_9750,N_9176);
nand U10171 (N_10171,N_9861,N_9728);
and U10172 (N_10172,N_9030,N_9405);
xnor U10173 (N_10173,N_9827,N_9504);
nor U10174 (N_10174,N_9152,N_9995);
or U10175 (N_10175,N_9801,N_9920);
or U10176 (N_10176,N_9840,N_9546);
and U10177 (N_10177,N_9867,N_9624);
and U10178 (N_10178,N_9069,N_9692);
nor U10179 (N_10179,N_9911,N_9589);
nand U10180 (N_10180,N_9793,N_9468);
or U10181 (N_10181,N_9918,N_9071);
or U10182 (N_10182,N_9474,N_9494);
or U10183 (N_10183,N_9644,N_9733);
xor U10184 (N_10184,N_9901,N_9519);
nand U10185 (N_10185,N_9583,N_9636);
or U10186 (N_10186,N_9221,N_9711);
and U10187 (N_10187,N_9631,N_9957);
or U10188 (N_10188,N_9308,N_9955);
or U10189 (N_10189,N_9259,N_9232);
nand U10190 (N_10190,N_9355,N_9365);
nand U10191 (N_10191,N_9328,N_9884);
and U10192 (N_10192,N_9453,N_9483);
and U10193 (N_10193,N_9005,N_9314);
and U10194 (N_10194,N_9393,N_9900);
xor U10195 (N_10195,N_9855,N_9880);
and U10196 (N_10196,N_9562,N_9926);
xor U10197 (N_10197,N_9825,N_9406);
and U10198 (N_10198,N_9376,N_9002);
nor U10199 (N_10199,N_9886,N_9714);
xnor U10200 (N_10200,N_9937,N_9837);
nor U10201 (N_10201,N_9508,N_9307);
and U10202 (N_10202,N_9997,N_9770);
and U10203 (N_10203,N_9138,N_9389);
or U10204 (N_10204,N_9808,N_9073);
nor U10205 (N_10205,N_9169,N_9696);
nand U10206 (N_10206,N_9809,N_9665);
nand U10207 (N_10207,N_9175,N_9027);
xor U10208 (N_10208,N_9285,N_9139);
and U10209 (N_10209,N_9260,N_9251);
xor U10210 (N_10210,N_9422,N_9092);
xnor U10211 (N_10211,N_9145,N_9402);
nand U10212 (N_10212,N_9087,N_9835);
nor U10213 (N_10213,N_9767,N_9290);
xor U10214 (N_10214,N_9917,N_9744);
xnor U10215 (N_10215,N_9529,N_9497);
or U10216 (N_10216,N_9751,N_9009);
and U10217 (N_10217,N_9363,N_9850);
nor U10218 (N_10218,N_9742,N_9719);
xor U10219 (N_10219,N_9682,N_9929);
or U10220 (N_10220,N_9202,N_9699);
xor U10221 (N_10221,N_9263,N_9912);
xor U10222 (N_10222,N_9396,N_9817);
nand U10223 (N_10223,N_9098,N_9209);
xor U10224 (N_10224,N_9947,N_9148);
nor U10225 (N_10225,N_9775,N_9953);
or U10226 (N_10226,N_9090,N_9574);
nor U10227 (N_10227,N_9296,N_9408);
or U10228 (N_10228,N_9046,N_9869);
xnor U10229 (N_10229,N_9522,N_9873);
and U10230 (N_10230,N_9354,N_9101);
xor U10231 (N_10231,N_9648,N_9933);
nor U10232 (N_10232,N_9476,N_9470);
nor U10233 (N_10233,N_9084,N_9018);
nand U10234 (N_10234,N_9029,N_9054);
xor U10235 (N_10235,N_9928,N_9865);
xor U10236 (N_10236,N_9068,N_9849);
or U10237 (N_10237,N_9813,N_9856);
and U10238 (N_10238,N_9510,N_9407);
xnor U10239 (N_10239,N_9876,N_9672);
nor U10240 (N_10240,N_9645,N_9951);
xor U10241 (N_10241,N_9653,N_9554);
xnor U10242 (N_10242,N_9450,N_9471);
and U10243 (N_10243,N_9811,N_9609);
xor U10244 (N_10244,N_9220,N_9077);
and U10245 (N_10245,N_9458,N_9666);
nand U10246 (N_10246,N_9255,N_9740);
nor U10247 (N_10247,N_9525,N_9509);
or U10248 (N_10248,N_9338,N_9874);
nand U10249 (N_10249,N_9400,N_9843);
nand U10250 (N_10250,N_9247,N_9608);
xor U10251 (N_10251,N_9892,N_9109);
and U10252 (N_10252,N_9196,N_9361);
and U10253 (N_10253,N_9125,N_9012);
nand U10254 (N_10254,N_9807,N_9045);
and U10255 (N_10255,N_9883,N_9560);
xor U10256 (N_10256,N_9960,N_9173);
nand U10257 (N_10257,N_9235,N_9585);
or U10258 (N_10258,N_9008,N_9761);
and U10259 (N_10259,N_9369,N_9561);
or U10260 (N_10260,N_9252,N_9944);
nor U10261 (N_10261,N_9322,N_9914);
and U10262 (N_10262,N_9925,N_9891);
or U10263 (N_10263,N_9144,N_9345);
nor U10264 (N_10264,N_9225,N_9231);
nand U10265 (N_10265,N_9033,N_9500);
or U10266 (N_10266,N_9760,N_9557);
xnor U10267 (N_10267,N_9567,N_9410);
nor U10268 (N_10268,N_9439,N_9305);
or U10269 (N_10269,N_9579,N_9321);
xor U10270 (N_10270,N_9539,N_9380);
nor U10271 (N_10271,N_9053,N_9044);
nand U10272 (N_10272,N_9897,N_9715);
xor U10273 (N_10273,N_9076,N_9623);
or U10274 (N_10274,N_9051,N_9303);
nand U10275 (N_10275,N_9160,N_9088);
and U10276 (N_10276,N_9155,N_9661);
nand U10277 (N_10277,N_9731,N_9278);
nand U10278 (N_10278,N_9015,N_9067);
and U10279 (N_10279,N_9486,N_9780);
or U10280 (N_10280,N_9816,N_9543);
nand U10281 (N_10281,N_9368,N_9013);
xor U10282 (N_10282,N_9603,N_9377);
and U10283 (N_10283,N_9357,N_9858);
and U10284 (N_10284,N_9007,N_9319);
and U10285 (N_10285,N_9541,N_9271);
nor U10286 (N_10286,N_9768,N_9667);
nand U10287 (N_10287,N_9317,N_9763);
nand U10288 (N_10288,N_9946,N_9984);
xor U10289 (N_10289,N_9164,N_9732);
or U10290 (N_10290,N_9275,N_9870);
and U10291 (N_10291,N_9383,N_9685);
nor U10292 (N_10292,N_9218,N_9282);
nor U10293 (N_10293,N_9475,N_9070);
nand U10294 (N_10294,N_9713,N_9170);
nor U10295 (N_10295,N_9229,N_9598);
xor U10296 (N_10296,N_9356,N_9765);
nor U10297 (N_10297,N_9064,N_9326);
nor U10298 (N_10298,N_9707,N_9107);
nand U10299 (N_10299,N_9460,N_9615);
nand U10300 (N_10300,N_9244,N_9441);
and U10301 (N_10301,N_9311,N_9847);
and U10302 (N_10302,N_9903,N_9506);
nand U10303 (N_10303,N_9397,N_9161);
or U10304 (N_10304,N_9783,N_9754);
nor U10305 (N_10305,N_9017,N_9547);
nor U10306 (N_10306,N_9384,N_9988);
and U10307 (N_10307,N_9135,N_9102);
or U10308 (N_10308,N_9993,N_9478);
and U10309 (N_10309,N_9969,N_9678);
nand U10310 (N_10310,N_9821,N_9201);
and U10311 (N_10311,N_9291,N_9484);
nor U10312 (N_10312,N_9055,N_9734);
xnor U10313 (N_10313,N_9452,N_9423);
xnor U10314 (N_10314,N_9776,N_9315);
or U10315 (N_10315,N_9952,N_9720);
nand U10316 (N_10316,N_9065,N_9594);
nor U10317 (N_10317,N_9288,N_9473);
and U10318 (N_10318,N_9530,N_9705);
xnor U10319 (N_10319,N_9572,N_9908);
nand U10320 (N_10320,N_9403,N_9324);
nand U10321 (N_10321,N_9404,N_9938);
nor U10322 (N_10322,N_9446,N_9331);
nand U10323 (N_10323,N_9243,N_9089);
nand U10324 (N_10324,N_9375,N_9626);
or U10325 (N_10325,N_9647,N_9919);
xnor U10326 (N_10326,N_9190,N_9137);
nor U10327 (N_10327,N_9688,N_9332);
nand U10328 (N_10328,N_9465,N_9792);
or U10329 (N_10329,N_9224,N_9060);
nor U10330 (N_10330,N_9359,N_9758);
nor U10331 (N_10331,N_9975,N_9899);
and U10332 (N_10332,N_9467,N_9479);
or U10333 (N_10333,N_9640,N_9469);
xor U10334 (N_10334,N_9444,N_9618);
xnor U10335 (N_10335,N_9185,N_9151);
nand U10336 (N_10336,N_9242,N_9620);
nor U10337 (N_10337,N_9590,N_9016);
xnor U10338 (N_10338,N_9651,N_9617);
or U10339 (N_10339,N_9536,N_9906);
xnor U10340 (N_10340,N_9853,N_9895);
and U10341 (N_10341,N_9223,N_9518);
xor U10342 (N_10342,N_9063,N_9413);
xor U10343 (N_10343,N_9698,N_9842);
nor U10344 (N_10344,N_9108,N_9131);
or U10345 (N_10345,N_9276,N_9693);
or U10346 (N_10346,N_9234,N_9382);
xnor U10347 (N_10347,N_9269,N_9851);
nor U10348 (N_10348,N_9724,N_9254);
nor U10349 (N_10349,N_9774,N_9512);
or U10350 (N_10350,N_9096,N_9293);
nor U10351 (N_10351,N_9704,N_9729);
nor U10352 (N_10352,N_9879,N_9463);
and U10353 (N_10353,N_9412,N_9716);
xnor U10354 (N_10354,N_9772,N_9274);
or U10355 (N_10355,N_9281,N_9120);
xnor U10356 (N_10356,N_9571,N_9921);
xnor U10357 (N_10357,N_9198,N_9563);
xnor U10358 (N_10358,N_9785,N_9941);
nand U10359 (N_10359,N_9828,N_9273);
nor U10360 (N_10360,N_9854,N_9158);
or U10361 (N_10361,N_9738,N_9814);
xor U10362 (N_10362,N_9199,N_9600);
or U10363 (N_10363,N_9425,N_9074);
and U10364 (N_10364,N_9034,N_9411);
xnor U10365 (N_10365,N_9495,N_9576);
nor U10366 (N_10366,N_9675,N_9177);
or U10367 (N_10367,N_9352,N_9123);
and U10368 (N_10368,N_9432,N_9959);
or U10369 (N_10369,N_9097,N_9249);
xor U10370 (N_10370,N_9456,N_9635);
or U10371 (N_10371,N_9584,N_9253);
nor U10372 (N_10372,N_9610,N_9511);
and U10373 (N_10373,N_9836,N_9373);
nand U10374 (N_10374,N_9387,N_9936);
nor U10375 (N_10375,N_9435,N_9445);
xnor U10376 (N_10376,N_9727,N_9464);
nand U10377 (N_10377,N_9904,N_9663);
xor U10378 (N_10378,N_9309,N_9652);
or U10379 (N_10379,N_9866,N_9378);
or U10380 (N_10380,N_9700,N_9638);
nand U10381 (N_10381,N_9860,N_9485);
xnor U10382 (N_10382,N_9105,N_9802);
nand U10383 (N_10383,N_9283,N_9746);
xnor U10384 (N_10384,N_9295,N_9250);
and U10385 (N_10385,N_9799,N_9735);
and U10386 (N_10386,N_9759,N_9300);
nand U10387 (N_10387,N_9893,N_9390);
nor U10388 (N_10388,N_9723,N_9553);
or U10389 (N_10389,N_9766,N_9019);
xnor U10390 (N_10390,N_9310,N_9871);
xor U10391 (N_10391,N_9945,N_9298);
nand U10392 (N_10392,N_9419,N_9797);
xor U10393 (N_10393,N_9272,N_9417);
and U10394 (N_10394,N_9915,N_9569);
and U10395 (N_10395,N_9043,N_9942);
or U10396 (N_10396,N_9709,N_9747);
nand U10397 (N_10397,N_9606,N_9313);
or U10398 (N_10398,N_9931,N_9513);
xor U10399 (N_10399,N_9973,N_9480);
nor U10400 (N_10400,N_9998,N_9784);
or U10401 (N_10401,N_9482,N_9565);
and U10402 (N_10402,N_9725,N_9238);
xnor U10403 (N_10403,N_9438,N_9286);
and U10404 (N_10404,N_9371,N_9974);
nor U10405 (N_10405,N_9781,N_9989);
or U10406 (N_10406,N_9461,N_9329);
and U10407 (N_10407,N_9570,N_9683);
or U10408 (N_10408,N_9179,N_9103);
nor U10409 (N_10409,N_9991,N_9431);
xor U10410 (N_10410,N_9420,N_9551);
nand U10411 (N_10411,N_9846,N_9752);
xor U10412 (N_10412,N_9990,N_9958);
and U10413 (N_10413,N_9520,N_9195);
xor U10414 (N_10414,N_9878,N_9031);
xnor U10415 (N_10415,N_9178,N_9351);
and U10416 (N_10416,N_9349,N_9490);
xnor U10417 (N_10417,N_9649,N_9344);
nor U10418 (N_10418,N_9163,N_9764);
nor U10419 (N_10419,N_9035,N_9430);
and U10420 (N_10420,N_9796,N_9592);
and U10421 (N_10421,N_9580,N_9128);
and U10422 (N_10422,N_9174,N_9659);
and U10423 (N_10423,N_9159,N_9424);
and U10424 (N_10424,N_9877,N_9042);
and U10425 (N_10425,N_9633,N_9180);
and U10426 (N_10426,N_9558,N_9721);
nand U10427 (N_10427,N_9540,N_9681);
and U10428 (N_10428,N_9923,N_9502);
xor U10429 (N_10429,N_9881,N_9256);
nor U10430 (N_10430,N_9815,N_9188);
xor U10431 (N_10431,N_9970,N_9333);
nand U10432 (N_10432,N_9182,N_9680);
nand U10433 (N_10433,N_9117,N_9769);
or U10434 (N_10434,N_9979,N_9341);
nand U10435 (N_10435,N_9833,N_9819);
xnor U10436 (N_10436,N_9078,N_9421);
nand U10437 (N_10437,N_9515,N_9095);
or U10438 (N_10438,N_9622,N_9994);
and U10439 (N_10439,N_9206,N_9862);
xnor U10440 (N_10440,N_9448,N_9487);
xor U10441 (N_10441,N_9777,N_9745);
nand U10442 (N_10442,N_9297,N_9434);
xnor U10443 (N_10443,N_9440,N_9050);
xnor U10444 (N_10444,N_9323,N_9790);
or U10445 (N_10445,N_9488,N_9104);
nor U10446 (N_10446,N_9587,N_9910);
and U10447 (N_10447,N_9718,N_9150);
or U10448 (N_10448,N_9954,N_9292);
xor U10449 (N_10449,N_9556,N_9335);
nand U10450 (N_10450,N_9629,N_9228);
and U10451 (N_10451,N_9694,N_9133);
nor U10452 (N_10452,N_9625,N_9786);
nand U10453 (N_10453,N_9094,N_9701);
xor U10454 (N_10454,N_9597,N_9136);
nand U10455 (N_10455,N_9184,N_9657);
nor U10456 (N_10456,N_9026,N_9537);
or U10457 (N_10457,N_9265,N_9596);
xnor U10458 (N_10458,N_9697,N_9010);
or U10459 (N_10459,N_9183,N_9927);
xor U10460 (N_10460,N_9114,N_9737);
xnor U10461 (N_10461,N_9454,N_9890);
nor U10462 (N_10462,N_9428,N_9142);
nand U10463 (N_10463,N_9655,N_9956);
xnor U10464 (N_10464,N_9392,N_9712);
xnor U10465 (N_10465,N_9347,N_9119);
and U10466 (N_10466,N_9048,N_9621);
xor U10467 (N_10467,N_9779,N_9437);
xor U10468 (N_10468,N_9771,N_9986);
nand U10469 (N_10469,N_9327,N_9233);
nor U10470 (N_10470,N_9642,N_9503);
nor U10471 (N_10471,N_9172,N_9052);
and U10472 (N_10472,N_9730,N_9829);
xor U10473 (N_10473,N_9320,N_9181);
and U10474 (N_10474,N_9838,N_9934);
and U10475 (N_10475,N_9246,N_9794);
or U10476 (N_10476,N_9350,N_9481);
xnor U10477 (N_10477,N_9258,N_9943);
or U10478 (N_10478,N_9346,N_9134);
or U10479 (N_10479,N_9795,N_9691);
or U10480 (N_10480,N_9548,N_9896);
or U10481 (N_10481,N_9491,N_9578);
or U10482 (N_10482,N_9340,N_9806);
or U10483 (N_10483,N_9203,N_9191);
or U10484 (N_10484,N_9773,N_9287);
or U10485 (N_10485,N_9684,N_9416);
or U10486 (N_10486,N_9964,N_9845);
or U10487 (N_10487,N_9523,N_9436);
nor U10488 (N_10488,N_9859,N_9894);
or U10489 (N_10489,N_9613,N_9913);
or U10490 (N_10490,N_9091,N_9261);
nand U10491 (N_10491,N_9193,N_9038);
and U10492 (N_10492,N_9226,N_9353);
xor U10493 (N_10493,N_9905,N_9654);
nor U10494 (N_10494,N_9207,N_9627);
nor U10495 (N_10495,N_9388,N_9212);
nand U10496 (N_10496,N_9047,N_9978);
or U10497 (N_10497,N_9695,N_9093);
nand U10498 (N_10498,N_9971,N_9372);
nand U10499 (N_10499,N_9976,N_9304);
nand U10500 (N_10500,N_9888,N_9614);
and U10501 (N_10501,N_9366,N_9383);
nand U10502 (N_10502,N_9363,N_9108);
or U10503 (N_10503,N_9596,N_9869);
and U10504 (N_10504,N_9637,N_9246);
nand U10505 (N_10505,N_9998,N_9671);
nand U10506 (N_10506,N_9087,N_9555);
and U10507 (N_10507,N_9623,N_9262);
or U10508 (N_10508,N_9467,N_9613);
nor U10509 (N_10509,N_9658,N_9449);
nor U10510 (N_10510,N_9600,N_9287);
nor U10511 (N_10511,N_9577,N_9348);
xor U10512 (N_10512,N_9742,N_9879);
and U10513 (N_10513,N_9498,N_9787);
or U10514 (N_10514,N_9609,N_9767);
or U10515 (N_10515,N_9261,N_9079);
and U10516 (N_10516,N_9692,N_9997);
or U10517 (N_10517,N_9839,N_9686);
nor U10518 (N_10518,N_9378,N_9190);
nand U10519 (N_10519,N_9558,N_9519);
nand U10520 (N_10520,N_9608,N_9680);
nor U10521 (N_10521,N_9963,N_9901);
or U10522 (N_10522,N_9184,N_9413);
or U10523 (N_10523,N_9139,N_9962);
or U10524 (N_10524,N_9919,N_9558);
nand U10525 (N_10525,N_9578,N_9254);
nor U10526 (N_10526,N_9942,N_9538);
nand U10527 (N_10527,N_9404,N_9764);
xor U10528 (N_10528,N_9545,N_9025);
nor U10529 (N_10529,N_9145,N_9521);
and U10530 (N_10530,N_9770,N_9273);
nor U10531 (N_10531,N_9918,N_9714);
nand U10532 (N_10532,N_9624,N_9607);
xor U10533 (N_10533,N_9980,N_9557);
or U10534 (N_10534,N_9494,N_9423);
or U10535 (N_10535,N_9357,N_9122);
and U10536 (N_10536,N_9826,N_9708);
nor U10537 (N_10537,N_9484,N_9224);
xor U10538 (N_10538,N_9886,N_9285);
or U10539 (N_10539,N_9816,N_9835);
nand U10540 (N_10540,N_9078,N_9389);
nand U10541 (N_10541,N_9637,N_9016);
or U10542 (N_10542,N_9675,N_9311);
nand U10543 (N_10543,N_9595,N_9164);
or U10544 (N_10544,N_9696,N_9173);
nand U10545 (N_10545,N_9232,N_9741);
or U10546 (N_10546,N_9670,N_9528);
nor U10547 (N_10547,N_9123,N_9156);
and U10548 (N_10548,N_9110,N_9321);
xor U10549 (N_10549,N_9943,N_9440);
nand U10550 (N_10550,N_9693,N_9047);
nand U10551 (N_10551,N_9726,N_9309);
nand U10552 (N_10552,N_9475,N_9872);
and U10553 (N_10553,N_9265,N_9545);
nand U10554 (N_10554,N_9942,N_9779);
and U10555 (N_10555,N_9143,N_9162);
and U10556 (N_10556,N_9767,N_9283);
or U10557 (N_10557,N_9503,N_9886);
xnor U10558 (N_10558,N_9164,N_9646);
nor U10559 (N_10559,N_9013,N_9444);
and U10560 (N_10560,N_9431,N_9940);
and U10561 (N_10561,N_9325,N_9398);
xnor U10562 (N_10562,N_9935,N_9245);
xnor U10563 (N_10563,N_9564,N_9346);
nor U10564 (N_10564,N_9125,N_9442);
or U10565 (N_10565,N_9303,N_9225);
nor U10566 (N_10566,N_9893,N_9961);
nand U10567 (N_10567,N_9844,N_9699);
xor U10568 (N_10568,N_9440,N_9869);
xor U10569 (N_10569,N_9757,N_9574);
and U10570 (N_10570,N_9917,N_9117);
or U10571 (N_10571,N_9396,N_9738);
nand U10572 (N_10572,N_9735,N_9077);
nor U10573 (N_10573,N_9265,N_9312);
nand U10574 (N_10574,N_9047,N_9554);
nand U10575 (N_10575,N_9311,N_9334);
or U10576 (N_10576,N_9280,N_9437);
xnor U10577 (N_10577,N_9629,N_9967);
nand U10578 (N_10578,N_9502,N_9844);
and U10579 (N_10579,N_9628,N_9275);
nor U10580 (N_10580,N_9115,N_9251);
nand U10581 (N_10581,N_9438,N_9451);
or U10582 (N_10582,N_9635,N_9996);
or U10583 (N_10583,N_9326,N_9358);
xnor U10584 (N_10584,N_9243,N_9575);
xnor U10585 (N_10585,N_9561,N_9589);
nand U10586 (N_10586,N_9182,N_9041);
or U10587 (N_10587,N_9343,N_9269);
or U10588 (N_10588,N_9284,N_9079);
xnor U10589 (N_10589,N_9385,N_9313);
xor U10590 (N_10590,N_9002,N_9185);
nor U10591 (N_10591,N_9434,N_9952);
nor U10592 (N_10592,N_9534,N_9270);
nor U10593 (N_10593,N_9700,N_9061);
nand U10594 (N_10594,N_9324,N_9168);
nor U10595 (N_10595,N_9074,N_9444);
nor U10596 (N_10596,N_9957,N_9773);
nor U10597 (N_10597,N_9018,N_9445);
nand U10598 (N_10598,N_9476,N_9916);
or U10599 (N_10599,N_9082,N_9095);
nor U10600 (N_10600,N_9387,N_9399);
and U10601 (N_10601,N_9016,N_9250);
and U10602 (N_10602,N_9673,N_9696);
nand U10603 (N_10603,N_9178,N_9406);
nor U10604 (N_10604,N_9160,N_9023);
xor U10605 (N_10605,N_9125,N_9925);
xnor U10606 (N_10606,N_9073,N_9428);
xor U10607 (N_10607,N_9190,N_9753);
xnor U10608 (N_10608,N_9296,N_9701);
and U10609 (N_10609,N_9286,N_9141);
nor U10610 (N_10610,N_9122,N_9381);
nor U10611 (N_10611,N_9300,N_9803);
xnor U10612 (N_10612,N_9283,N_9364);
or U10613 (N_10613,N_9641,N_9556);
and U10614 (N_10614,N_9730,N_9038);
and U10615 (N_10615,N_9705,N_9164);
xnor U10616 (N_10616,N_9113,N_9797);
and U10617 (N_10617,N_9796,N_9208);
and U10618 (N_10618,N_9190,N_9593);
or U10619 (N_10619,N_9067,N_9237);
nand U10620 (N_10620,N_9107,N_9223);
nand U10621 (N_10621,N_9454,N_9547);
xor U10622 (N_10622,N_9885,N_9554);
xor U10623 (N_10623,N_9343,N_9277);
and U10624 (N_10624,N_9951,N_9926);
nand U10625 (N_10625,N_9149,N_9458);
nor U10626 (N_10626,N_9307,N_9791);
nand U10627 (N_10627,N_9705,N_9249);
nor U10628 (N_10628,N_9451,N_9802);
xor U10629 (N_10629,N_9323,N_9151);
and U10630 (N_10630,N_9492,N_9107);
or U10631 (N_10631,N_9788,N_9005);
nand U10632 (N_10632,N_9870,N_9526);
xnor U10633 (N_10633,N_9992,N_9583);
and U10634 (N_10634,N_9927,N_9114);
and U10635 (N_10635,N_9247,N_9099);
and U10636 (N_10636,N_9885,N_9790);
and U10637 (N_10637,N_9854,N_9372);
nor U10638 (N_10638,N_9788,N_9169);
or U10639 (N_10639,N_9090,N_9699);
xnor U10640 (N_10640,N_9472,N_9175);
or U10641 (N_10641,N_9349,N_9904);
nor U10642 (N_10642,N_9160,N_9469);
nand U10643 (N_10643,N_9243,N_9196);
xnor U10644 (N_10644,N_9945,N_9315);
xor U10645 (N_10645,N_9131,N_9665);
and U10646 (N_10646,N_9726,N_9927);
or U10647 (N_10647,N_9828,N_9680);
and U10648 (N_10648,N_9546,N_9214);
and U10649 (N_10649,N_9855,N_9508);
xor U10650 (N_10650,N_9938,N_9156);
or U10651 (N_10651,N_9407,N_9773);
and U10652 (N_10652,N_9858,N_9023);
and U10653 (N_10653,N_9896,N_9446);
nand U10654 (N_10654,N_9241,N_9168);
and U10655 (N_10655,N_9820,N_9414);
and U10656 (N_10656,N_9306,N_9460);
nor U10657 (N_10657,N_9207,N_9384);
nor U10658 (N_10658,N_9873,N_9680);
xnor U10659 (N_10659,N_9671,N_9538);
nor U10660 (N_10660,N_9239,N_9482);
nor U10661 (N_10661,N_9948,N_9407);
nand U10662 (N_10662,N_9541,N_9756);
and U10663 (N_10663,N_9629,N_9957);
and U10664 (N_10664,N_9734,N_9658);
and U10665 (N_10665,N_9233,N_9518);
xor U10666 (N_10666,N_9400,N_9493);
and U10667 (N_10667,N_9709,N_9149);
nor U10668 (N_10668,N_9809,N_9283);
and U10669 (N_10669,N_9275,N_9431);
and U10670 (N_10670,N_9405,N_9977);
nand U10671 (N_10671,N_9784,N_9735);
and U10672 (N_10672,N_9625,N_9959);
and U10673 (N_10673,N_9049,N_9041);
nor U10674 (N_10674,N_9161,N_9557);
and U10675 (N_10675,N_9132,N_9504);
nor U10676 (N_10676,N_9808,N_9231);
nor U10677 (N_10677,N_9423,N_9247);
nand U10678 (N_10678,N_9649,N_9381);
or U10679 (N_10679,N_9616,N_9215);
and U10680 (N_10680,N_9538,N_9630);
and U10681 (N_10681,N_9018,N_9381);
nor U10682 (N_10682,N_9534,N_9901);
or U10683 (N_10683,N_9779,N_9525);
nor U10684 (N_10684,N_9554,N_9164);
and U10685 (N_10685,N_9656,N_9905);
nor U10686 (N_10686,N_9450,N_9518);
nor U10687 (N_10687,N_9898,N_9346);
or U10688 (N_10688,N_9430,N_9885);
nor U10689 (N_10689,N_9005,N_9211);
xnor U10690 (N_10690,N_9998,N_9917);
xnor U10691 (N_10691,N_9935,N_9529);
or U10692 (N_10692,N_9348,N_9851);
or U10693 (N_10693,N_9176,N_9113);
nor U10694 (N_10694,N_9748,N_9085);
xor U10695 (N_10695,N_9228,N_9185);
nand U10696 (N_10696,N_9000,N_9494);
nor U10697 (N_10697,N_9062,N_9490);
xor U10698 (N_10698,N_9229,N_9065);
xor U10699 (N_10699,N_9538,N_9577);
nand U10700 (N_10700,N_9640,N_9739);
nand U10701 (N_10701,N_9821,N_9017);
xor U10702 (N_10702,N_9711,N_9087);
or U10703 (N_10703,N_9875,N_9447);
nor U10704 (N_10704,N_9402,N_9405);
nor U10705 (N_10705,N_9926,N_9446);
and U10706 (N_10706,N_9189,N_9433);
and U10707 (N_10707,N_9623,N_9617);
xnor U10708 (N_10708,N_9146,N_9984);
nand U10709 (N_10709,N_9493,N_9093);
xnor U10710 (N_10710,N_9874,N_9045);
nand U10711 (N_10711,N_9478,N_9151);
and U10712 (N_10712,N_9248,N_9130);
nand U10713 (N_10713,N_9179,N_9053);
or U10714 (N_10714,N_9946,N_9618);
and U10715 (N_10715,N_9653,N_9725);
or U10716 (N_10716,N_9912,N_9319);
nand U10717 (N_10717,N_9782,N_9918);
and U10718 (N_10718,N_9415,N_9202);
nand U10719 (N_10719,N_9361,N_9695);
and U10720 (N_10720,N_9641,N_9274);
nand U10721 (N_10721,N_9080,N_9562);
nand U10722 (N_10722,N_9768,N_9425);
and U10723 (N_10723,N_9481,N_9062);
xor U10724 (N_10724,N_9418,N_9650);
nor U10725 (N_10725,N_9964,N_9729);
nor U10726 (N_10726,N_9351,N_9265);
and U10727 (N_10727,N_9876,N_9397);
or U10728 (N_10728,N_9061,N_9476);
nor U10729 (N_10729,N_9157,N_9371);
nor U10730 (N_10730,N_9655,N_9508);
and U10731 (N_10731,N_9135,N_9255);
xor U10732 (N_10732,N_9205,N_9933);
nor U10733 (N_10733,N_9234,N_9391);
xnor U10734 (N_10734,N_9118,N_9160);
or U10735 (N_10735,N_9416,N_9491);
or U10736 (N_10736,N_9322,N_9170);
or U10737 (N_10737,N_9457,N_9189);
nand U10738 (N_10738,N_9055,N_9831);
and U10739 (N_10739,N_9406,N_9548);
xor U10740 (N_10740,N_9261,N_9687);
xnor U10741 (N_10741,N_9158,N_9390);
nor U10742 (N_10742,N_9120,N_9509);
and U10743 (N_10743,N_9063,N_9203);
xor U10744 (N_10744,N_9229,N_9687);
xor U10745 (N_10745,N_9997,N_9336);
xor U10746 (N_10746,N_9919,N_9630);
and U10747 (N_10747,N_9216,N_9391);
or U10748 (N_10748,N_9265,N_9045);
nor U10749 (N_10749,N_9969,N_9994);
or U10750 (N_10750,N_9262,N_9797);
or U10751 (N_10751,N_9809,N_9629);
or U10752 (N_10752,N_9297,N_9673);
nor U10753 (N_10753,N_9265,N_9911);
xor U10754 (N_10754,N_9598,N_9634);
or U10755 (N_10755,N_9903,N_9454);
nand U10756 (N_10756,N_9811,N_9487);
xnor U10757 (N_10757,N_9038,N_9506);
or U10758 (N_10758,N_9579,N_9651);
or U10759 (N_10759,N_9113,N_9019);
and U10760 (N_10760,N_9856,N_9275);
nor U10761 (N_10761,N_9681,N_9501);
nor U10762 (N_10762,N_9580,N_9418);
xnor U10763 (N_10763,N_9484,N_9115);
nor U10764 (N_10764,N_9464,N_9052);
nand U10765 (N_10765,N_9192,N_9834);
xor U10766 (N_10766,N_9839,N_9327);
nand U10767 (N_10767,N_9384,N_9045);
nand U10768 (N_10768,N_9260,N_9908);
or U10769 (N_10769,N_9881,N_9271);
nand U10770 (N_10770,N_9220,N_9982);
nand U10771 (N_10771,N_9977,N_9473);
or U10772 (N_10772,N_9827,N_9656);
nand U10773 (N_10773,N_9267,N_9181);
and U10774 (N_10774,N_9309,N_9906);
xnor U10775 (N_10775,N_9472,N_9958);
nor U10776 (N_10776,N_9674,N_9870);
nand U10777 (N_10777,N_9647,N_9532);
nand U10778 (N_10778,N_9887,N_9341);
xnor U10779 (N_10779,N_9850,N_9387);
xnor U10780 (N_10780,N_9544,N_9513);
nand U10781 (N_10781,N_9665,N_9655);
nand U10782 (N_10782,N_9804,N_9762);
xor U10783 (N_10783,N_9015,N_9242);
xnor U10784 (N_10784,N_9527,N_9626);
or U10785 (N_10785,N_9445,N_9290);
nor U10786 (N_10786,N_9383,N_9890);
and U10787 (N_10787,N_9044,N_9245);
nand U10788 (N_10788,N_9772,N_9367);
nor U10789 (N_10789,N_9809,N_9958);
or U10790 (N_10790,N_9832,N_9087);
nor U10791 (N_10791,N_9353,N_9585);
or U10792 (N_10792,N_9345,N_9164);
xnor U10793 (N_10793,N_9881,N_9191);
nand U10794 (N_10794,N_9355,N_9226);
nand U10795 (N_10795,N_9511,N_9530);
and U10796 (N_10796,N_9225,N_9147);
xor U10797 (N_10797,N_9526,N_9466);
nand U10798 (N_10798,N_9228,N_9170);
xor U10799 (N_10799,N_9624,N_9214);
or U10800 (N_10800,N_9223,N_9026);
nand U10801 (N_10801,N_9521,N_9385);
or U10802 (N_10802,N_9196,N_9429);
nor U10803 (N_10803,N_9657,N_9662);
and U10804 (N_10804,N_9394,N_9275);
and U10805 (N_10805,N_9638,N_9503);
nand U10806 (N_10806,N_9600,N_9188);
nand U10807 (N_10807,N_9772,N_9174);
or U10808 (N_10808,N_9593,N_9764);
nor U10809 (N_10809,N_9681,N_9771);
and U10810 (N_10810,N_9934,N_9286);
nor U10811 (N_10811,N_9159,N_9878);
and U10812 (N_10812,N_9080,N_9381);
nor U10813 (N_10813,N_9744,N_9915);
nand U10814 (N_10814,N_9104,N_9061);
and U10815 (N_10815,N_9419,N_9057);
xor U10816 (N_10816,N_9717,N_9181);
nor U10817 (N_10817,N_9374,N_9980);
or U10818 (N_10818,N_9996,N_9477);
xnor U10819 (N_10819,N_9916,N_9475);
nand U10820 (N_10820,N_9266,N_9248);
nor U10821 (N_10821,N_9486,N_9482);
nor U10822 (N_10822,N_9948,N_9863);
nor U10823 (N_10823,N_9660,N_9578);
xor U10824 (N_10824,N_9394,N_9572);
and U10825 (N_10825,N_9943,N_9388);
and U10826 (N_10826,N_9683,N_9261);
nand U10827 (N_10827,N_9627,N_9158);
nor U10828 (N_10828,N_9455,N_9282);
and U10829 (N_10829,N_9270,N_9732);
or U10830 (N_10830,N_9170,N_9640);
nand U10831 (N_10831,N_9556,N_9030);
and U10832 (N_10832,N_9677,N_9760);
or U10833 (N_10833,N_9514,N_9380);
xor U10834 (N_10834,N_9581,N_9202);
or U10835 (N_10835,N_9492,N_9263);
or U10836 (N_10836,N_9068,N_9308);
or U10837 (N_10837,N_9920,N_9403);
xor U10838 (N_10838,N_9657,N_9572);
xnor U10839 (N_10839,N_9132,N_9109);
or U10840 (N_10840,N_9832,N_9422);
nor U10841 (N_10841,N_9030,N_9239);
nor U10842 (N_10842,N_9115,N_9570);
xnor U10843 (N_10843,N_9518,N_9488);
xnor U10844 (N_10844,N_9021,N_9740);
and U10845 (N_10845,N_9985,N_9984);
nor U10846 (N_10846,N_9755,N_9424);
xnor U10847 (N_10847,N_9484,N_9783);
and U10848 (N_10848,N_9888,N_9335);
and U10849 (N_10849,N_9237,N_9983);
and U10850 (N_10850,N_9264,N_9525);
and U10851 (N_10851,N_9516,N_9988);
xnor U10852 (N_10852,N_9123,N_9683);
nor U10853 (N_10853,N_9148,N_9312);
or U10854 (N_10854,N_9762,N_9229);
or U10855 (N_10855,N_9632,N_9700);
nand U10856 (N_10856,N_9668,N_9572);
or U10857 (N_10857,N_9062,N_9181);
nor U10858 (N_10858,N_9197,N_9781);
nand U10859 (N_10859,N_9019,N_9944);
or U10860 (N_10860,N_9951,N_9306);
nand U10861 (N_10861,N_9415,N_9621);
xor U10862 (N_10862,N_9505,N_9928);
nor U10863 (N_10863,N_9176,N_9372);
xnor U10864 (N_10864,N_9568,N_9777);
nand U10865 (N_10865,N_9572,N_9143);
nor U10866 (N_10866,N_9764,N_9524);
or U10867 (N_10867,N_9767,N_9779);
nor U10868 (N_10868,N_9529,N_9048);
nor U10869 (N_10869,N_9771,N_9510);
or U10870 (N_10870,N_9984,N_9617);
xor U10871 (N_10871,N_9935,N_9585);
nand U10872 (N_10872,N_9579,N_9618);
nor U10873 (N_10873,N_9592,N_9794);
nor U10874 (N_10874,N_9524,N_9354);
and U10875 (N_10875,N_9774,N_9265);
or U10876 (N_10876,N_9208,N_9252);
nand U10877 (N_10877,N_9024,N_9146);
xnor U10878 (N_10878,N_9528,N_9295);
and U10879 (N_10879,N_9745,N_9086);
or U10880 (N_10880,N_9725,N_9319);
and U10881 (N_10881,N_9809,N_9995);
xor U10882 (N_10882,N_9098,N_9733);
xnor U10883 (N_10883,N_9916,N_9341);
xnor U10884 (N_10884,N_9106,N_9148);
or U10885 (N_10885,N_9734,N_9356);
nor U10886 (N_10886,N_9690,N_9087);
nand U10887 (N_10887,N_9464,N_9275);
xnor U10888 (N_10888,N_9080,N_9795);
or U10889 (N_10889,N_9249,N_9402);
or U10890 (N_10890,N_9795,N_9541);
nand U10891 (N_10891,N_9820,N_9175);
nor U10892 (N_10892,N_9242,N_9776);
nor U10893 (N_10893,N_9932,N_9170);
xor U10894 (N_10894,N_9546,N_9155);
xor U10895 (N_10895,N_9873,N_9588);
and U10896 (N_10896,N_9190,N_9239);
nand U10897 (N_10897,N_9428,N_9723);
and U10898 (N_10898,N_9985,N_9958);
or U10899 (N_10899,N_9894,N_9358);
or U10900 (N_10900,N_9251,N_9795);
or U10901 (N_10901,N_9959,N_9171);
or U10902 (N_10902,N_9372,N_9388);
xor U10903 (N_10903,N_9394,N_9241);
and U10904 (N_10904,N_9281,N_9024);
nor U10905 (N_10905,N_9004,N_9346);
or U10906 (N_10906,N_9538,N_9755);
and U10907 (N_10907,N_9748,N_9933);
and U10908 (N_10908,N_9008,N_9504);
or U10909 (N_10909,N_9679,N_9073);
nor U10910 (N_10910,N_9034,N_9651);
nor U10911 (N_10911,N_9219,N_9450);
xor U10912 (N_10912,N_9046,N_9852);
nand U10913 (N_10913,N_9510,N_9141);
nand U10914 (N_10914,N_9594,N_9674);
xor U10915 (N_10915,N_9161,N_9892);
nor U10916 (N_10916,N_9468,N_9309);
and U10917 (N_10917,N_9969,N_9024);
or U10918 (N_10918,N_9322,N_9916);
nor U10919 (N_10919,N_9678,N_9881);
nor U10920 (N_10920,N_9261,N_9883);
nand U10921 (N_10921,N_9063,N_9917);
nor U10922 (N_10922,N_9778,N_9718);
xnor U10923 (N_10923,N_9861,N_9739);
nand U10924 (N_10924,N_9362,N_9657);
and U10925 (N_10925,N_9518,N_9227);
nand U10926 (N_10926,N_9073,N_9994);
or U10927 (N_10927,N_9245,N_9620);
nand U10928 (N_10928,N_9197,N_9615);
or U10929 (N_10929,N_9942,N_9061);
or U10930 (N_10930,N_9336,N_9082);
or U10931 (N_10931,N_9086,N_9808);
or U10932 (N_10932,N_9985,N_9418);
nand U10933 (N_10933,N_9066,N_9987);
xor U10934 (N_10934,N_9307,N_9936);
xnor U10935 (N_10935,N_9497,N_9182);
and U10936 (N_10936,N_9742,N_9454);
nor U10937 (N_10937,N_9580,N_9971);
xor U10938 (N_10938,N_9603,N_9433);
nand U10939 (N_10939,N_9568,N_9648);
xnor U10940 (N_10940,N_9349,N_9854);
nor U10941 (N_10941,N_9682,N_9439);
nand U10942 (N_10942,N_9896,N_9493);
nor U10943 (N_10943,N_9668,N_9178);
or U10944 (N_10944,N_9224,N_9790);
and U10945 (N_10945,N_9931,N_9785);
nor U10946 (N_10946,N_9639,N_9268);
and U10947 (N_10947,N_9309,N_9913);
nor U10948 (N_10948,N_9639,N_9089);
or U10949 (N_10949,N_9244,N_9292);
or U10950 (N_10950,N_9298,N_9537);
or U10951 (N_10951,N_9635,N_9231);
nand U10952 (N_10952,N_9146,N_9880);
nand U10953 (N_10953,N_9115,N_9063);
or U10954 (N_10954,N_9961,N_9381);
xnor U10955 (N_10955,N_9669,N_9209);
xnor U10956 (N_10956,N_9804,N_9044);
or U10957 (N_10957,N_9224,N_9513);
nand U10958 (N_10958,N_9053,N_9861);
nor U10959 (N_10959,N_9763,N_9657);
and U10960 (N_10960,N_9592,N_9569);
nor U10961 (N_10961,N_9191,N_9132);
or U10962 (N_10962,N_9941,N_9217);
nor U10963 (N_10963,N_9975,N_9024);
and U10964 (N_10964,N_9332,N_9579);
or U10965 (N_10965,N_9174,N_9890);
xor U10966 (N_10966,N_9258,N_9968);
nand U10967 (N_10967,N_9209,N_9636);
nand U10968 (N_10968,N_9001,N_9316);
nand U10969 (N_10969,N_9262,N_9457);
nor U10970 (N_10970,N_9381,N_9284);
nor U10971 (N_10971,N_9526,N_9156);
xnor U10972 (N_10972,N_9479,N_9117);
or U10973 (N_10973,N_9237,N_9990);
xnor U10974 (N_10974,N_9870,N_9643);
nand U10975 (N_10975,N_9252,N_9075);
and U10976 (N_10976,N_9548,N_9505);
and U10977 (N_10977,N_9858,N_9354);
xnor U10978 (N_10978,N_9891,N_9119);
and U10979 (N_10979,N_9734,N_9841);
and U10980 (N_10980,N_9105,N_9576);
nand U10981 (N_10981,N_9135,N_9684);
and U10982 (N_10982,N_9103,N_9130);
or U10983 (N_10983,N_9410,N_9418);
and U10984 (N_10984,N_9278,N_9391);
and U10985 (N_10985,N_9272,N_9268);
xnor U10986 (N_10986,N_9788,N_9748);
nor U10987 (N_10987,N_9188,N_9603);
nand U10988 (N_10988,N_9956,N_9281);
nor U10989 (N_10989,N_9766,N_9891);
and U10990 (N_10990,N_9569,N_9759);
nor U10991 (N_10991,N_9580,N_9652);
nand U10992 (N_10992,N_9724,N_9936);
xnor U10993 (N_10993,N_9716,N_9956);
nor U10994 (N_10994,N_9717,N_9456);
or U10995 (N_10995,N_9513,N_9856);
nand U10996 (N_10996,N_9653,N_9868);
xor U10997 (N_10997,N_9087,N_9466);
xnor U10998 (N_10998,N_9667,N_9250);
xnor U10999 (N_10999,N_9402,N_9938);
xnor U11000 (N_11000,N_10601,N_10646);
and U11001 (N_11001,N_10648,N_10330);
xnor U11002 (N_11002,N_10293,N_10668);
or U11003 (N_11003,N_10983,N_10764);
nor U11004 (N_11004,N_10962,N_10893);
nand U11005 (N_11005,N_10947,N_10072);
xor U11006 (N_11006,N_10760,N_10027);
nor U11007 (N_11007,N_10345,N_10918);
or U11008 (N_11008,N_10631,N_10123);
and U11009 (N_11009,N_10169,N_10722);
nand U11010 (N_11010,N_10633,N_10076);
or U11011 (N_11011,N_10116,N_10559);
or U11012 (N_11012,N_10925,N_10261);
nand U11013 (N_11013,N_10409,N_10984);
xnor U11014 (N_11014,N_10029,N_10859);
xnor U11015 (N_11015,N_10567,N_10794);
nand U11016 (N_11016,N_10328,N_10767);
or U11017 (N_11017,N_10912,N_10647);
and U11018 (N_11018,N_10299,N_10817);
or U11019 (N_11019,N_10968,N_10804);
nand U11020 (N_11020,N_10250,N_10606);
xnor U11021 (N_11021,N_10142,N_10307);
and U11022 (N_11022,N_10212,N_10678);
or U11023 (N_11023,N_10824,N_10527);
or U11024 (N_11024,N_10177,N_10295);
xor U11025 (N_11025,N_10810,N_10531);
and U11026 (N_11026,N_10480,N_10883);
nand U11027 (N_11027,N_10078,N_10879);
or U11028 (N_11028,N_10946,N_10043);
nor U11029 (N_11029,N_10639,N_10097);
or U11030 (N_11030,N_10613,N_10511);
nor U11031 (N_11031,N_10037,N_10599);
nor U11032 (N_11032,N_10198,N_10755);
or U11033 (N_11033,N_10865,N_10023);
nor U11034 (N_11034,N_10120,N_10706);
xor U11035 (N_11035,N_10199,N_10447);
and U11036 (N_11036,N_10827,N_10541);
nand U11037 (N_11037,N_10329,N_10263);
nor U11038 (N_11038,N_10216,N_10162);
or U11039 (N_11039,N_10287,N_10259);
nor U11040 (N_11040,N_10642,N_10506);
nor U11041 (N_11041,N_10994,N_10269);
xor U11042 (N_11042,N_10791,N_10862);
xnor U11043 (N_11043,N_10666,N_10481);
xor U11044 (N_11044,N_10430,N_10114);
nor U11045 (N_11045,N_10225,N_10474);
or U11046 (N_11046,N_10508,N_10540);
and U11047 (N_11047,N_10267,N_10277);
or U11048 (N_11048,N_10604,N_10429);
and U11049 (N_11049,N_10058,N_10868);
xnor U11050 (N_11050,N_10999,N_10725);
nor U11051 (N_11051,N_10542,N_10008);
xnor U11052 (N_11052,N_10680,N_10244);
and U11053 (N_11053,N_10094,N_10450);
and U11054 (N_11054,N_10135,N_10358);
nor U11055 (N_11055,N_10797,N_10594);
and U11056 (N_11056,N_10363,N_10007);
xor U11057 (N_11057,N_10009,N_10603);
nand U11058 (N_11058,N_10993,N_10738);
xnor U11059 (N_11059,N_10533,N_10718);
nand U11060 (N_11060,N_10995,N_10271);
xor U11061 (N_11061,N_10191,N_10170);
nand U11062 (N_11062,N_10825,N_10987);
or U11063 (N_11063,N_10458,N_10470);
xnor U11064 (N_11064,N_10001,N_10418);
xor U11065 (N_11065,N_10944,N_10514);
or U11066 (N_11066,N_10251,N_10012);
nor U11067 (N_11067,N_10134,N_10843);
or U11068 (N_11068,N_10276,N_10951);
nand U11069 (N_11069,N_10935,N_10252);
or U11070 (N_11070,N_10714,N_10888);
nand U11071 (N_11071,N_10886,N_10332);
and U11072 (N_11072,N_10898,N_10592);
and U11073 (N_11073,N_10716,N_10586);
and U11074 (N_11074,N_10548,N_10917);
nor U11075 (N_11075,N_10851,N_10789);
nand U11076 (N_11076,N_10786,N_10117);
and U11077 (N_11077,N_10090,N_10692);
xor U11078 (N_11078,N_10889,N_10712);
nand U11079 (N_11079,N_10897,N_10530);
nor U11080 (N_11080,N_10923,N_10327);
nand U11081 (N_11081,N_10131,N_10290);
and U11082 (N_11082,N_10873,N_10473);
xor U11083 (N_11083,N_10636,N_10899);
or U11084 (N_11084,N_10776,N_10801);
nor U11085 (N_11085,N_10537,N_10010);
or U11086 (N_11086,N_10071,N_10337);
and U11087 (N_11087,N_10203,N_10294);
nand U11088 (N_11088,N_10301,N_10557);
nor U11089 (N_11089,N_10919,N_10449);
nor U11090 (N_11090,N_10857,N_10763);
nand U11091 (N_11091,N_10839,N_10468);
or U11092 (N_11092,N_10619,N_10482);
nand U11093 (N_11093,N_10448,N_10353);
and U11094 (N_11094,N_10284,N_10502);
nand U11095 (N_11095,N_10781,N_10664);
nand U11096 (N_11096,N_10461,N_10878);
and U11097 (N_11097,N_10655,N_10635);
nor U11098 (N_11098,N_10545,N_10910);
and U11099 (N_11099,N_10414,N_10890);
and U11100 (N_11100,N_10595,N_10772);
or U11101 (N_11101,N_10986,N_10066);
xor U11102 (N_11102,N_10534,N_10156);
xnor U11103 (N_11103,N_10721,N_10036);
nor U11104 (N_11104,N_10675,N_10611);
nor U11105 (N_11105,N_10849,N_10264);
or U11106 (N_11106,N_10629,N_10625);
and U11107 (N_11107,N_10411,N_10615);
nor U11108 (N_11108,N_10281,N_10937);
nand U11109 (N_11109,N_10192,N_10892);
nand U11110 (N_11110,N_10576,N_10671);
xor U11111 (N_11111,N_10719,N_10331);
nand U11112 (N_11112,N_10723,N_10324);
xnor U11113 (N_11113,N_10698,N_10348);
nor U11114 (N_11114,N_10194,N_10869);
nor U11115 (N_11115,N_10350,N_10217);
nor U11116 (N_11116,N_10741,N_10283);
nor U11117 (N_11117,N_10992,N_10355);
and U11118 (N_11118,N_10375,N_10852);
nor U11119 (N_11119,N_10729,N_10174);
nor U11120 (N_11120,N_10863,N_10553);
or U11121 (N_11121,N_10588,N_10507);
xor U11122 (N_11122,N_10376,N_10206);
or U11123 (N_11123,N_10247,N_10197);
and U11124 (N_11124,N_10513,N_10491);
xnor U11125 (N_11125,N_10504,N_10652);
xnor U11126 (N_11126,N_10710,N_10026);
and U11127 (N_11127,N_10128,N_10143);
or U11128 (N_11128,N_10039,N_10459);
nand U11129 (N_11129,N_10093,N_10799);
or U11130 (N_11130,N_10172,N_10150);
xor U11131 (N_11131,N_10018,N_10105);
nand U11132 (N_11132,N_10014,N_10657);
nand U11133 (N_11133,N_10248,N_10386);
or U11134 (N_11134,N_10478,N_10304);
or U11135 (N_11135,N_10193,N_10104);
and U11136 (N_11136,N_10352,N_10979);
nand U11137 (N_11137,N_10069,N_10795);
nor U11138 (N_11138,N_10452,N_10109);
or U11139 (N_11139,N_10052,N_10998);
or U11140 (N_11140,N_10146,N_10147);
xnor U11141 (N_11141,N_10028,N_10616);
nand U11142 (N_11142,N_10361,N_10079);
and U11143 (N_11143,N_10543,N_10630);
nand U11144 (N_11144,N_10273,N_10546);
xor U11145 (N_11145,N_10798,N_10322);
nand U11146 (N_11146,N_10569,N_10050);
xor U11147 (N_11147,N_10469,N_10341);
nor U11148 (N_11148,N_10628,N_10242);
nor U11149 (N_11149,N_10676,N_10720);
nand U11150 (N_11150,N_10550,N_10484);
and U11151 (N_11151,N_10590,N_10187);
and U11152 (N_11152,N_10391,N_10260);
nand U11153 (N_11153,N_10617,N_10634);
or U11154 (N_11154,N_10982,N_10285);
nand U11155 (N_11155,N_10130,N_10920);
nand U11156 (N_11156,N_10171,N_10988);
nor U11157 (N_11157,N_10913,N_10685);
nand U11158 (N_11158,N_10015,N_10864);
or U11159 (N_11159,N_10425,N_10035);
xnor U11160 (N_11160,N_10739,N_10532);
nand U11161 (N_11161,N_10077,N_10451);
or U11162 (N_11162,N_10492,N_10765);
nand U11163 (N_11163,N_10038,N_10748);
and U11164 (N_11164,N_10577,N_10936);
and U11165 (N_11165,N_10231,N_10743);
or U11166 (N_11166,N_10949,N_10821);
nand U11167 (N_11167,N_10997,N_10833);
and U11168 (N_11168,N_10370,N_10049);
xor U11169 (N_11169,N_10288,N_10236);
nand U11170 (N_11170,N_10224,N_10674);
nor U11171 (N_11171,N_10265,N_10965);
nor U11172 (N_11172,N_10940,N_10420);
and U11173 (N_11173,N_10768,N_10214);
or U11174 (N_11174,N_10434,N_10245);
xnor U11175 (N_11175,N_10239,N_10660);
or U11176 (N_11176,N_10040,N_10841);
nor U11177 (N_11177,N_10189,N_10486);
or U11178 (N_11178,N_10963,N_10818);
xnor U11179 (N_11179,N_10319,N_10895);
and U11180 (N_11180,N_10070,N_10046);
nand U11181 (N_11181,N_10784,N_10462);
nor U11182 (N_11182,N_10233,N_10119);
or U11183 (N_11183,N_10702,N_10313);
nand U11184 (N_11184,N_10275,N_10083);
nor U11185 (N_11185,N_10292,N_10339);
or U11186 (N_11186,N_10318,N_10138);
and U11187 (N_11187,N_10455,N_10691);
xor U11188 (N_11188,N_10773,N_10802);
nand U11189 (N_11189,N_10911,N_10783);
nand U11190 (N_11190,N_10905,N_10378);
or U11191 (N_11191,N_10551,N_10842);
or U11192 (N_11192,N_10521,N_10382);
nand U11193 (N_11193,N_10493,N_10445);
xnor U11194 (N_11194,N_10608,N_10432);
and U11195 (N_11195,N_10204,N_10638);
nand U11196 (N_11196,N_10834,N_10344);
xor U11197 (N_11197,N_10145,N_10067);
nand U11198 (N_11198,N_10336,N_10485);
and U11199 (N_11199,N_10106,N_10308);
nand U11200 (N_11200,N_10321,N_10175);
or U11201 (N_11201,N_10368,N_10234);
nor U11202 (N_11202,N_10402,N_10042);
xnor U11203 (N_11203,N_10113,N_10574);
xor U11204 (N_11204,N_10637,N_10747);
nand U11205 (N_11205,N_10844,N_10195);
xnor U11206 (N_11206,N_10373,N_10854);
or U11207 (N_11207,N_10168,N_10465);
xnor U11208 (N_11208,N_10510,N_10367);
nand U11209 (N_11209,N_10778,N_10400);
nand U11210 (N_11210,N_10365,N_10823);
or U11211 (N_11211,N_10315,N_10737);
nor U11212 (N_11212,N_10053,N_10185);
xnor U11213 (N_11213,N_10314,N_10974);
nand U11214 (N_11214,N_10746,N_10446);
nand U11215 (N_11215,N_10082,N_10884);
or U11216 (N_11216,N_10064,N_10412);
and U11217 (N_11217,N_10835,N_10074);
nand U11218 (N_11218,N_10041,N_10441);
nor U11219 (N_11219,N_10300,N_10958);
and U11220 (N_11220,N_10587,N_10305);
or U11221 (N_11221,N_10934,N_10061);
and U11222 (N_11222,N_10153,N_10707);
nor U11223 (N_11223,N_10693,N_10578);
nand U11224 (N_11224,N_10969,N_10564);
nor U11225 (N_11225,N_10101,N_10397);
xor U11226 (N_11226,N_10697,N_10051);
nand U11227 (N_11227,N_10522,N_10356);
and U11228 (N_11228,N_10512,N_10663);
nand U11229 (N_11229,N_10990,N_10938);
nand U11230 (N_11230,N_10600,N_10408);
xor U11231 (N_11231,N_10133,N_10535);
xnor U11232 (N_11232,N_10091,N_10891);
or U11233 (N_11233,N_10605,N_10807);
and U11234 (N_11234,N_10985,N_10715);
or U11235 (N_11235,N_10280,N_10068);
xor U11236 (N_11236,N_10334,N_10607);
or U11237 (N_11237,N_10494,N_10749);
and U11238 (N_11238,N_10243,N_10205);
nor U11239 (N_11239,N_10745,N_10179);
xor U11240 (N_11240,N_10831,N_10479);
xnor U11241 (N_11241,N_10699,N_10812);
nand U11242 (N_11242,N_10930,N_10907);
xor U11243 (N_11243,N_10961,N_10705);
xnor U11244 (N_11244,N_10756,N_10270);
xnor U11245 (N_11245,N_10549,N_10065);
or U11246 (N_11246,N_10048,N_10904);
nand U11247 (N_11247,N_10967,N_10659);
nor U11248 (N_11248,N_10524,N_10387);
and U11249 (N_11249,N_10614,N_10928);
or U11250 (N_11250,N_10152,N_10144);
or U11251 (N_11251,N_10730,N_10796);
and U11252 (N_11252,N_10004,N_10310);
xnor U11253 (N_11253,N_10505,N_10838);
and U11254 (N_11254,N_10347,N_10257);
xnor U11255 (N_11255,N_10673,N_10054);
and U11256 (N_11256,N_10980,N_10098);
and U11257 (N_11257,N_10683,N_10782);
or U11258 (N_11258,N_10771,N_10333);
and U11259 (N_11259,N_10538,N_10686);
or U11260 (N_11260,N_10176,N_10080);
nand U11261 (N_11261,N_10132,N_10346);
nor U11262 (N_11262,N_10845,N_10374);
and U11263 (N_11263,N_10226,N_10896);
nor U11264 (N_11264,N_10256,N_10253);
nand U11265 (N_11265,N_10955,N_10240);
and U11266 (N_11266,N_10742,N_10816);
and U11267 (N_11267,N_10112,N_10774);
nor U11268 (N_11268,N_10490,N_10207);
xnor U11269 (N_11269,N_10581,N_10309);
nor U11270 (N_11270,N_10151,N_10840);
and U11271 (N_11271,N_10621,N_10921);
nor U11272 (N_11272,N_10561,N_10596);
xnor U11273 (N_11273,N_10249,N_10417);
and U11274 (N_11274,N_10927,N_10653);
xor U11275 (N_11275,N_10654,N_10125);
nor U11276 (N_11276,N_10213,N_10326);
xor U11277 (N_11277,N_10424,N_10279);
xor U11278 (N_11278,N_10011,N_10670);
nor U11279 (N_11279,N_10395,N_10853);
and U11280 (N_11280,N_10620,N_10274);
and U11281 (N_11281,N_10343,N_10750);
nor U11282 (N_11282,N_10403,N_10002);
xor U11283 (N_11283,N_10460,N_10832);
xor U11284 (N_11284,N_10566,N_10689);
nor U11285 (N_11285,N_10384,N_10235);
nor U11286 (N_11286,N_10255,N_10882);
and U11287 (N_11287,N_10939,N_10266);
and U11288 (N_11288,N_10929,N_10181);
nand U11289 (N_11289,N_10597,N_10931);
nor U11290 (N_11290,N_10487,N_10149);
and U11291 (N_11291,N_10419,N_10320);
nand U11292 (N_11292,N_10866,N_10973);
xnor U11293 (N_11293,N_10221,N_10354);
nor U11294 (N_11294,N_10338,N_10392);
nor U11295 (N_11295,N_10762,N_10059);
nand U11296 (N_11296,N_10690,N_10111);
and U11297 (N_11297,N_10503,N_10941);
xor U11298 (N_11298,N_10063,N_10602);
and U11299 (N_11299,N_10006,N_10154);
or U11300 (N_11300,N_10383,N_10860);
nor U11301 (N_11301,N_10708,N_10219);
nor U11302 (N_11302,N_10736,N_10020);
or U11303 (N_11303,N_10140,N_10759);
and U11304 (N_11304,N_10959,N_10081);
and U11305 (N_11305,N_10463,N_10871);
nand U11306 (N_11306,N_10095,N_10900);
or U11307 (N_11307,N_10396,N_10836);
nor U11308 (N_11308,N_10410,N_10665);
xor U11309 (N_11309,N_10394,N_10407);
nor U11310 (N_11310,N_10901,N_10751);
or U11311 (N_11311,N_10830,N_10909);
or U11312 (N_11312,N_10573,N_10717);
nand U11313 (N_11313,N_10727,N_10681);
and U11314 (N_11314,N_10682,N_10302);
or U11315 (N_11315,N_10024,N_10454);
nand U11316 (N_11316,N_10389,N_10811);
or U11317 (N_11317,N_10554,N_10388);
or U11318 (N_11318,N_10464,N_10158);
xnor U11319 (N_11319,N_10291,N_10536);
nand U11320 (N_11320,N_10317,N_10627);
nand U11321 (N_11321,N_10585,N_10254);
and U11322 (N_11322,N_10021,N_10489);
or U11323 (N_11323,N_10696,N_10643);
nor U11324 (N_11324,N_10528,N_10335);
or U11325 (N_11325,N_10096,N_10438);
xor U11326 (N_11326,N_10003,N_10115);
nor U11327 (N_11327,N_10060,N_10100);
nor U11328 (N_11328,N_10289,N_10770);
xnor U11329 (N_11329,N_10428,N_10877);
xor U11330 (N_11330,N_10644,N_10754);
nor U11331 (N_11331,N_10806,N_10677);
nor U11332 (N_11332,N_10552,N_10850);
xor U11333 (N_11333,N_10110,N_10467);
xnor U11334 (N_11334,N_10422,N_10572);
and U11335 (N_11335,N_10325,N_10238);
or U11336 (N_11336,N_10735,N_10571);
nor U11337 (N_11337,N_10874,N_10342);
xor U11338 (N_11338,N_10084,N_10870);
and U11339 (N_11339,N_10210,N_10031);
or U11340 (N_11340,N_10672,N_10013);
nand U11341 (N_11341,N_10858,N_10229);
and U11342 (N_11342,N_10045,N_10780);
and U11343 (N_11343,N_10954,N_10583);
and U11344 (N_11344,N_10570,N_10453);
nand U11345 (N_11345,N_10000,N_10731);
nand U11346 (N_11346,N_10829,N_10087);
nor U11347 (N_11347,N_10431,N_10560);
and U11348 (N_11348,N_10433,N_10822);
nand U11349 (N_11349,N_10501,N_10753);
and U11350 (N_11350,N_10519,N_10139);
nor U11351 (N_11351,N_10278,N_10598);
nor U11352 (N_11352,N_10649,N_10016);
and U11353 (N_11353,N_10127,N_10894);
nor U11354 (N_11354,N_10196,N_10443);
nor U11355 (N_11355,N_10201,N_10471);
and U11356 (N_11356,N_10568,N_10475);
and U11357 (N_11357,N_10499,N_10565);
and U11358 (N_11358,N_10498,N_10775);
and U11359 (N_11359,N_10656,N_10034);
nand U11360 (N_11360,N_10591,N_10488);
or U11361 (N_11361,N_10726,N_10711);
or U11362 (N_11362,N_10948,N_10903);
nor U11363 (N_11363,N_10057,N_10136);
xnor U11364 (N_11364,N_10978,N_10401);
nor U11365 (N_11365,N_10377,N_10323);
and U11366 (N_11366,N_10220,N_10785);
xnor U11367 (N_11367,N_10086,N_10662);
nand U11368 (N_11368,N_10349,N_10359);
xnor U11369 (N_11369,N_10525,N_10183);
nor U11370 (N_11370,N_10167,N_10924);
and U11371 (N_11371,N_10357,N_10808);
xor U11372 (N_11372,N_10881,N_10188);
or U11373 (N_11373,N_10157,N_10790);
nor U11374 (N_11374,N_10472,N_10700);
and U11375 (N_11375,N_10209,N_10232);
xor U11376 (N_11376,N_10610,N_10709);
or U11377 (N_11377,N_10173,N_10103);
and U11378 (N_11378,N_10483,N_10286);
or U11379 (N_11379,N_10575,N_10792);
xnor U11380 (N_11380,N_10916,N_10371);
and U11381 (N_11381,N_10427,N_10362);
and U11382 (N_11382,N_10957,N_10972);
nor U11383 (N_11383,N_10159,N_10141);
xor U11384 (N_11384,N_10056,N_10495);
xor U11385 (N_11385,N_10372,N_10062);
nor U11386 (N_11386,N_10661,N_10520);
and U11387 (N_11387,N_10752,N_10529);
nor U11388 (N_11388,N_10073,N_10744);
nor U11389 (N_11389,N_10926,N_10099);
nand U11390 (N_11390,N_10724,N_10230);
nor U11391 (N_11391,N_10178,N_10915);
xnor U11392 (N_11392,N_10970,N_10885);
xor U11393 (N_11393,N_10122,N_10025);
and U11394 (N_11394,N_10404,N_10258);
nand U11395 (N_11395,N_10416,N_10044);
nand U11396 (N_11396,N_10593,N_10163);
or U11397 (N_11397,N_10517,N_10645);
nand U11398 (N_11398,N_10033,N_10089);
nor U11399 (N_11399,N_10624,N_10164);
or U11400 (N_11400,N_10922,N_10847);
or U11401 (N_11401,N_10500,N_10932);
nand U11402 (N_11402,N_10989,N_10728);
and U11403 (N_11403,N_10875,N_10952);
nor U11404 (N_11404,N_10813,N_10953);
nor U11405 (N_11405,N_10369,N_10311);
nor U11406 (N_11406,N_10227,N_10547);
xnor U11407 (N_11407,N_10047,N_10848);
or U11408 (N_11408,N_10766,N_10732);
xnor U11409 (N_11409,N_10148,N_10914);
xnor U11410 (N_11410,N_10055,N_10703);
or U11411 (N_11411,N_10695,N_10757);
xnor U11412 (N_11412,N_10155,N_10075);
or U11413 (N_11413,N_10108,N_10622);
or U11414 (N_11414,N_10618,N_10945);
or U11415 (N_11415,N_10713,N_10184);
xor U11416 (N_11416,N_10684,N_10366);
nand U11417 (N_11417,N_10902,N_10241);
and U11418 (N_11418,N_10558,N_10129);
or U11419 (N_11419,N_10211,N_10861);
nor U11420 (N_11420,N_10223,N_10942);
and U11421 (N_11421,N_10867,N_10005);
and U11422 (N_11422,N_10828,N_10312);
nor U11423 (N_11423,N_10906,N_10996);
and U11424 (N_11424,N_10837,N_10956);
nand U11425 (N_11425,N_10316,N_10518);
and U11426 (N_11426,N_10761,N_10964);
or U11427 (N_11427,N_10436,N_10423);
xnor U11428 (N_11428,N_10161,N_10297);
or U11429 (N_11429,N_10688,N_10124);
xnor U11430 (N_11430,N_10667,N_10439);
xnor U11431 (N_11431,N_10971,N_10640);
nor U11432 (N_11432,N_10805,N_10215);
nor U11433 (N_11433,N_10406,N_10966);
or U11434 (N_11434,N_10539,N_10496);
nand U11435 (N_11435,N_10814,N_10800);
nor U11436 (N_11436,N_10562,N_10121);
xnor U11437 (N_11437,N_10200,N_10019);
and U11438 (N_11438,N_10017,N_10364);
and U11439 (N_11439,N_10415,N_10779);
and U11440 (N_11440,N_10515,N_10815);
nand U11441 (N_11441,N_10202,N_10933);
or U11442 (N_11442,N_10237,N_10222);
nand U11443 (N_11443,N_10880,N_10740);
or U11444 (N_11444,N_10444,N_10580);
and U11445 (N_11445,N_10088,N_10166);
xor U11446 (N_11446,N_10526,N_10268);
nor U11447 (N_11447,N_10820,N_10556);
nand U11448 (N_11448,N_10516,N_10092);
or U11449 (N_11449,N_10632,N_10413);
or U11450 (N_11450,N_10704,N_10421);
nor U11451 (N_11451,N_10032,N_10950);
nand U11452 (N_11452,N_10442,N_10612);
nor U11453 (N_11453,N_10793,N_10650);
nor U11454 (N_11454,N_10544,N_10186);
or U11455 (N_11455,N_10908,N_10380);
xnor U11456 (N_11456,N_10306,N_10609);
or U11457 (N_11457,N_10360,N_10296);
nor U11458 (N_11458,N_10523,N_10399);
nor U11459 (N_11459,N_10509,N_10658);
nor U11460 (N_11460,N_10477,N_10803);
nor U11461 (N_11461,N_10180,N_10426);
or U11462 (N_11462,N_10228,N_10734);
nor U11463 (N_11463,N_10819,N_10437);
or U11464 (N_11464,N_10777,N_10282);
and U11465 (N_11465,N_10435,N_10589);
and U11466 (N_11466,N_10943,N_10218);
xnor U11467 (N_11467,N_10887,N_10769);
nor U11468 (N_11468,N_10246,N_10623);
xor U11469 (N_11469,N_10476,N_10440);
or U11470 (N_11470,N_10669,N_10030);
nor U11471 (N_11471,N_10687,N_10208);
or U11472 (N_11472,N_10876,N_10733);
xor U11473 (N_11473,N_10456,N_10855);
and U11474 (N_11474,N_10582,N_10846);
nor U11475 (N_11475,N_10398,N_10272);
and U11476 (N_11476,N_10118,N_10975);
nand U11477 (N_11477,N_10393,N_10626);
and U11478 (N_11478,N_10679,N_10126);
xnor U11479 (N_11479,N_10137,N_10022);
and U11480 (N_11480,N_10182,N_10351);
xor U11481 (N_11481,N_10701,N_10981);
nand U11482 (N_11482,N_10584,N_10457);
xor U11483 (N_11483,N_10381,N_10390);
nor U11484 (N_11484,N_10107,N_10856);
nand U11485 (N_11485,N_10976,N_10303);
or U11486 (N_11486,N_10160,N_10262);
nand U11487 (N_11487,N_10788,N_10977);
or U11488 (N_11488,N_10298,N_10809);
nor U11489 (N_11489,N_10960,N_10694);
nor U11490 (N_11490,N_10497,N_10872);
and U11491 (N_11491,N_10379,N_10563);
and U11492 (N_11492,N_10466,N_10405);
nor U11493 (N_11493,N_10165,N_10555);
nor U11494 (N_11494,N_10991,N_10579);
nor U11495 (N_11495,N_10190,N_10102);
xor U11496 (N_11496,N_10085,N_10651);
nor U11497 (N_11497,N_10340,N_10758);
nand U11498 (N_11498,N_10787,N_10385);
and U11499 (N_11499,N_10826,N_10641);
nand U11500 (N_11500,N_10361,N_10301);
and U11501 (N_11501,N_10866,N_10353);
xor U11502 (N_11502,N_10287,N_10267);
or U11503 (N_11503,N_10610,N_10841);
xnor U11504 (N_11504,N_10816,N_10713);
nand U11505 (N_11505,N_10826,N_10082);
nand U11506 (N_11506,N_10386,N_10261);
nand U11507 (N_11507,N_10054,N_10375);
nor U11508 (N_11508,N_10968,N_10487);
nand U11509 (N_11509,N_10395,N_10733);
nor U11510 (N_11510,N_10096,N_10374);
nand U11511 (N_11511,N_10412,N_10205);
nand U11512 (N_11512,N_10884,N_10361);
nor U11513 (N_11513,N_10026,N_10900);
xor U11514 (N_11514,N_10048,N_10981);
nand U11515 (N_11515,N_10462,N_10944);
nor U11516 (N_11516,N_10174,N_10664);
or U11517 (N_11517,N_10047,N_10007);
nand U11518 (N_11518,N_10675,N_10061);
nor U11519 (N_11519,N_10896,N_10108);
nand U11520 (N_11520,N_10668,N_10334);
nor U11521 (N_11521,N_10690,N_10020);
xnor U11522 (N_11522,N_10106,N_10160);
and U11523 (N_11523,N_10759,N_10095);
nor U11524 (N_11524,N_10689,N_10357);
or U11525 (N_11525,N_10933,N_10025);
and U11526 (N_11526,N_10171,N_10888);
or U11527 (N_11527,N_10638,N_10636);
and U11528 (N_11528,N_10863,N_10928);
and U11529 (N_11529,N_10330,N_10542);
xor U11530 (N_11530,N_10831,N_10757);
nor U11531 (N_11531,N_10283,N_10068);
nand U11532 (N_11532,N_10317,N_10489);
nor U11533 (N_11533,N_10668,N_10857);
or U11534 (N_11534,N_10943,N_10028);
nor U11535 (N_11535,N_10144,N_10618);
xnor U11536 (N_11536,N_10944,N_10055);
xor U11537 (N_11537,N_10427,N_10738);
xnor U11538 (N_11538,N_10477,N_10564);
nor U11539 (N_11539,N_10215,N_10719);
nand U11540 (N_11540,N_10166,N_10800);
and U11541 (N_11541,N_10914,N_10781);
nand U11542 (N_11542,N_10066,N_10431);
and U11543 (N_11543,N_10931,N_10879);
or U11544 (N_11544,N_10385,N_10974);
nor U11545 (N_11545,N_10702,N_10974);
nor U11546 (N_11546,N_10618,N_10926);
nand U11547 (N_11547,N_10862,N_10932);
nor U11548 (N_11548,N_10059,N_10308);
nor U11549 (N_11549,N_10052,N_10316);
xnor U11550 (N_11550,N_10886,N_10900);
nand U11551 (N_11551,N_10955,N_10519);
and U11552 (N_11552,N_10023,N_10606);
nor U11553 (N_11553,N_10808,N_10885);
xor U11554 (N_11554,N_10528,N_10836);
nand U11555 (N_11555,N_10555,N_10202);
xor U11556 (N_11556,N_10885,N_10124);
and U11557 (N_11557,N_10455,N_10937);
xnor U11558 (N_11558,N_10138,N_10858);
and U11559 (N_11559,N_10852,N_10643);
or U11560 (N_11560,N_10727,N_10215);
and U11561 (N_11561,N_10869,N_10459);
and U11562 (N_11562,N_10044,N_10415);
or U11563 (N_11563,N_10385,N_10457);
nand U11564 (N_11564,N_10588,N_10243);
and U11565 (N_11565,N_10126,N_10969);
nand U11566 (N_11566,N_10570,N_10421);
or U11567 (N_11567,N_10077,N_10791);
and U11568 (N_11568,N_10182,N_10600);
and U11569 (N_11569,N_10673,N_10380);
nor U11570 (N_11570,N_10291,N_10577);
nor U11571 (N_11571,N_10335,N_10969);
nor U11572 (N_11572,N_10206,N_10325);
and U11573 (N_11573,N_10461,N_10127);
xor U11574 (N_11574,N_10747,N_10915);
or U11575 (N_11575,N_10763,N_10092);
nand U11576 (N_11576,N_10672,N_10344);
and U11577 (N_11577,N_10694,N_10767);
nor U11578 (N_11578,N_10571,N_10589);
and U11579 (N_11579,N_10202,N_10503);
nand U11580 (N_11580,N_10149,N_10796);
xor U11581 (N_11581,N_10349,N_10135);
xor U11582 (N_11582,N_10733,N_10350);
or U11583 (N_11583,N_10253,N_10866);
xor U11584 (N_11584,N_10531,N_10929);
nor U11585 (N_11585,N_10279,N_10597);
nand U11586 (N_11586,N_10810,N_10328);
and U11587 (N_11587,N_10074,N_10932);
xor U11588 (N_11588,N_10651,N_10778);
and U11589 (N_11589,N_10596,N_10879);
xnor U11590 (N_11590,N_10978,N_10814);
or U11591 (N_11591,N_10395,N_10471);
and U11592 (N_11592,N_10920,N_10774);
or U11593 (N_11593,N_10107,N_10328);
or U11594 (N_11594,N_10722,N_10606);
nor U11595 (N_11595,N_10959,N_10051);
or U11596 (N_11596,N_10330,N_10627);
nor U11597 (N_11597,N_10675,N_10354);
and U11598 (N_11598,N_10048,N_10635);
nor U11599 (N_11599,N_10291,N_10814);
nor U11600 (N_11600,N_10108,N_10626);
and U11601 (N_11601,N_10766,N_10330);
nor U11602 (N_11602,N_10233,N_10731);
or U11603 (N_11603,N_10971,N_10592);
or U11604 (N_11604,N_10333,N_10269);
and U11605 (N_11605,N_10571,N_10613);
xor U11606 (N_11606,N_10259,N_10748);
and U11607 (N_11607,N_10730,N_10641);
or U11608 (N_11608,N_10347,N_10339);
nand U11609 (N_11609,N_10178,N_10953);
nand U11610 (N_11610,N_10450,N_10627);
nand U11611 (N_11611,N_10808,N_10198);
and U11612 (N_11612,N_10737,N_10253);
or U11613 (N_11613,N_10198,N_10599);
and U11614 (N_11614,N_10766,N_10056);
nand U11615 (N_11615,N_10385,N_10198);
and U11616 (N_11616,N_10844,N_10039);
or U11617 (N_11617,N_10002,N_10086);
nor U11618 (N_11618,N_10430,N_10426);
nor U11619 (N_11619,N_10867,N_10590);
nor U11620 (N_11620,N_10149,N_10402);
or U11621 (N_11621,N_10243,N_10814);
or U11622 (N_11622,N_10566,N_10660);
nand U11623 (N_11623,N_10750,N_10666);
xnor U11624 (N_11624,N_10773,N_10241);
nand U11625 (N_11625,N_10991,N_10775);
nor U11626 (N_11626,N_10162,N_10817);
and U11627 (N_11627,N_10269,N_10273);
nor U11628 (N_11628,N_10662,N_10923);
nor U11629 (N_11629,N_10339,N_10400);
and U11630 (N_11630,N_10889,N_10823);
and U11631 (N_11631,N_10302,N_10522);
nand U11632 (N_11632,N_10895,N_10397);
or U11633 (N_11633,N_10850,N_10551);
nor U11634 (N_11634,N_10746,N_10543);
or U11635 (N_11635,N_10010,N_10469);
and U11636 (N_11636,N_10662,N_10509);
and U11637 (N_11637,N_10800,N_10229);
nand U11638 (N_11638,N_10167,N_10003);
nor U11639 (N_11639,N_10723,N_10231);
xor U11640 (N_11640,N_10067,N_10910);
xor U11641 (N_11641,N_10943,N_10260);
xnor U11642 (N_11642,N_10091,N_10094);
and U11643 (N_11643,N_10419,N_10543);
or U11644 (N_11644,N_10275,N_10038);
nor U11645 (N_11645,N_10697,N_10545);
xor U11646 (N_11646,N_10648,N_10836);
nor U11647 (N_11647,N_10762,N_10405);
and U11648 (N_11648,N_10504,N_10509);
xnor U11649 (N_11649,N_10336,N_10118);
xnor U11650 (N_11650,N_10517,N_10635);
xnor U11651 (N_11651,N_10953,N_10660);
nor U11652 (N_11652,N_10019,N_10238);
or U11653 (N_11653,N_10313,N_10380);
or U11654 (N_11654,N_10843,N_10431);
xor U11655 (N_11655,N_10598,N_10355);
nor U11656 (N_11656,N_10545,N_10234);
xnor U11657 (N_11657,N_10153,N_10915);
xor U11658 (N_11658,N_10943,N_10327);
nor U11659 (N_11659,N_10342,N_10943);
or U11660 (N_11660,N_10713,N_10608);
and U11661 (N_11661,N_10188,N_10656);
and U11662 (N_11662,N_10854,N_10520);
and U11663 (N_11663,N_10411,N_10768);
nor U11664 (N_11664,N_10904,N_10136);
nor U11665 (N_11665,N_10919,N_10075);
nor U11666 (N_11666,N_10907,N_10703);
or U11667 (N_11667,N_10518,N_10938);
xor U11668 (N_11668,N_10841,N_10494);
nor U11669 (N_11669,N_10947,N_10624);
nor U11670 (N_11670,N_10323,N_10815);
nor U11671 (N_11671,N_10146,N_10594);
xor U11672 (N_11672,N_10538,N_10264);
and U11673 (N_11673,N_10453,N_10031);
nor U11674 (N_11674,N_10356,N_10397);
and U11675 (N_11675,N_10050,N_10798);
and U11676 (N_11676,N_10078,N_10843);
and U11677 (N_11677,N_10805,N_10546);
xnor U11678 (N_11678,N_10086,N_10498);
and U11679 (N_11679,N_10431,N_10274);
nand U11680 (N_11680,N_10424,N_10592);
or U11681 (N_11681,N_10149,N_10838);
xnor U11682 (N_11682,N_10606,N_10933);
nor U11683 (N_11683,N_10143,N_10399);
or U11684 (N_11684,N_10832,N_10009);
nor U11685 (N_11685,N_10459,N_10035);
nand U11686 (N_11686,N_10361,N_10830);
and U11687 (N_11687,N_10706,N_10712);
nand U11688 (N_11688,N_10116,N_10086);
nand U11689 (N_11689,N_10427,N_10816);
nor U11690 (N_11690,N_10349,N_10481);
nor U11691 (N_11691,N_10585,N_10298);
and U11692 (N_11692,N_10783,N_10257);
or U11693 (N_11693,N_10117,N_10242);
or U11694 (N_11694,N_10590,N_10615);
or U11695 (N_11695,N_10745,N_10540);
nand U11696 (N_11696,N_10810,N_10730);
and U11697 (N_11697,N_10468,N_10074);
nor U11698 (N_11698,N_10145,N_10283);
xor U11699 (N_11699,N_10999,N_10252);
nor U11700 (N_11700,N_10531,N_10753);
or U11701 (N_11701,N_10842,N_10929);
xor U11702 (N_11702,N_10939,N_10719);
or U11703 (N_11703,N_10224,N_10636);
nor U11704 (N_11704,N_10340,N_10334);
or U11705 (N_11705,N_10946,N_10530);
or U11706 (N_11706,N_10772,N_10776);
nor U11707 (N_11707,N_10822,N_10292);
nand U11708 (N_11708,N_10091,N_10736);
nand U11709 (N_11709,N_10562,N_10415);
or U11710 (N_11710,N_10700,N_10308);
xnor U11711 (N_11711,N_10104,N_10058);
and U11712 (N_11712,N_10565,N_10664);
and U11713 (N_11713,N_10618,N_10466);
xnor U11714 (N_11714,N_10031,N_10544);
nand U11715 (N_11715,N_10749,N_10143);
or U11716 (N_11716,N_10268,N_10583);
and U11717 (N_11717,N_10176,N_10809);
nand U11718 (N_11718,N_10922,N_10219);
nand U11719 (N_11719,N_10790,N_10028);
nor U11720 (N_11720,N_10507,N_10750);
nand U11721 (N_11721,N_10056,N_10259);
or U11722 (N_11722,N_10371,N_10159);
or U11723 (N_11723,N_10232,N_10137);
xor U11724 (N_11724,N_10239,N_10383);
and U11725 (N_11725,N_10322,N_10469);
nor U11726 (N_11726,N_10576,N_10727);
xor U11727 (N_11727,N_10214,N_10560);
and U11728 (N_11728,N_10694,N_10300);
or U11729 (N_11729,N_10486,N_10306);
or U11730 (N_11730,N_10430,N_10660);
and U11731 (N_11731,N_10392,N_10694);
nor U11732 (N_11732,N_10277,N_10692);
nor U11733 (N_11733,N_10101,N_10798);
nor U11734 (N_11734,N_10679,N_10011);
xor U11735 (N_11735,N_10308,N_10713);
xor U11736 (N_11736,N_10099,N_10699);
or U11737 (N_11737,N_10938,N_10586);
nand U11738 (N_11738,N_10052,N_10424);
or U11739 (N_11739,N_10542,N_10551);
xor U11740 (N_11740,N_10070,N_10283);
nand U11741 (N_11741,N_10252,N_10187);
xor U11742 (N_11742,N_10994,N_10772);
nand U11743 (N_11743,N_10315,N_10400);
and U11744 (N_11744,N_10068,N_10683);
nand U11745 (N_11745,N_10437,N_10240);
nand U11746 (N_11746,N_10437,N_10016);
xnor U11747 (N_11747,N_10861,N_10180);
or U11748 (N_11748,N_10356,N_10060);
nor U11749 (N_11749,N_10213,N_10121);
xor U11750 (N_11750,N_10459,N_10804);
nor U11751 (N_11751,N_10784,N_10131);
nor U11752 (N_11752,N_10549,N_10386);
or U11753 (N_11753,N_10043,N_10354);
xor U11754 (N_11754,N_10472,N_10890);
xor U11755 (N_11755,N_10156,N_10282);
nor U11756 (N_11756,N_10855,N_10534);
and U11757 (N_11757,N_10865,N_10382);
nor U11758 (N_11758,N_10479,N_10546);
or U11759 (N_11759,N_10747,N_10706);
xor U11760 (N_11760,N_10547,N_10167);
and U11761 (N_11761,N_10657,N_10691);
nand U11762 (N_11762,N_10226,N_10680);
nor U11763 (N_11763,N_10856,N_10805);
xnor U11764 (N_11764,N_10945,N_10196);
and U11765 (N_11765,N_10118,N_10151);
nand U11766 (N_11766,N_10220,N_10677);
or U11767 (N_11767,N_10326,N_10186);
nand U11768 (N_11768,N_10280,N_10494);
and U11769 (N_11769,N_10460,N_10982);
xor U11770 (N_11770,N_10655,N_10158);
nor U11771 (N_11771,N_10893,N_10963);
and U11772 (N_11772,N_10753,N_10197);
nor U11773 (N_11773,N_10559,N_10485);
or U11774 (N_11774,N_10710,N_10930);
nor U11775 (N_11775,N_10084,N_10175);
nor U11776 (N_11776,N_10609,N_10446);
nor U11777 (N_11777,N_10809,N_10685);
nand U11778 (N_11778,N_10912,N_10259);
xor U11779 (N_11779,N_10153,N_10766);
and U11780 (N_11780,N_10822,N_10933);
or U11781 (N_11781,N_10321,N_10446);
or U11782 (N_11782,N_10243,N_10046);
xor U11783 (N_11783,N_10651,N_10723);
or U11784 (N_11784,N_10847,N_10661);
or U11785 (N_11785,N_10734,N_10917);
nor U11786 (N_11786,N_10757,N_10042);
and U11787 (N_11787,N_10130,N_10760);
nor U11788 (N_11788,N_10109,N_10708);
nand U11789 (N_11789,N_10984,N_10576);
nor U11790 (N_11790,N_10203,N_10381);
xnor U11791 (N_11791,N_10104,N_10567);
xnor U11792 (N_11792,N_10741,N_10838);
xor U11793 (N_11793,N_10992,N_10369);
xnor U11794 (N_11794,N_10196,N_10367);
nor U11795 (N_11795,N_10696,N_10588);
and U11796 (N_11796,N_10745,N_10208);
and U11797 (N_11797,N_10451,N_10006);
or U11798 (N_11798,N_10824,N_10551);
nand U11799 (N_11799,N_10699,N_10886);
xor U11800 (N_11800,N_10379,N_10494);
xor U11801 (N_11801,N_10694,N_10761);
or U11802 (N_11802,N_10284,N_10231);
and U11803 (N_11803,N_10263,N_10137);
nor U11804 (N_11804,N_10092,N_10665);
nand U11805 (N_11805,N_10480,N_10737);
nand U11806 (N_11806,N_10830,N_10069);
xnor U11807 (N_11807,N_10835,N_10185);
nor U11808 (N_11808,N_10943,N_10613);
nor U11809 (N_11809,N_10489,N_10593);
nor U11810 (N_11810,N_10278,N_10704);
or U11811 (N_11811,N_10567,N_10316);
or U11812 (N_11812,N_10780,N_10116);
nand U11813 (N_11813,N_10517,N_10335);
nand U11814 (N_11814,N_10060,N_10279);
xor U11815 (N_11815,N_10374,N_10640);
or U11816 (N_11816,N_10711,N_10447);
xor U11817 (N_11817,N_10701,N_10230);
xnor U11818 (N_11818,N_10102,N_10491);
xor U11819 (N_11819,N_10958,N_10464);
xnor U11820 (N_11820,N_10713,N_10063);
xnor U11821 (N_11821,N_10411,N_10020);
or U11822 (N_11822,N_10576,N_10661);
and U11823 (N_11823,N_10470,N_10640);
nand U11824 (N_11824,N_10918,N_10603);
nand U11825 (N_11825,N_10011,N_10688);
nand U11826 (N_11826,N_10492,N_10516);
and U11827 (N_11827,N_10703,N_10202);
and U11828 (N_11828,N_10076,N_10999);
or U11829 (N_11829,N_10619,N_10545);
nand U11830 (N_11830,N_10038,N_10700);
or U11831 (N_11831,N_10870,N_10270);
or U11832 (N_11832,N_10841,N_10577);
xnor U11833 (N_11833,N_10953,N_10821);
or U11834 (N_11834,N_10610,N_10611);
nor U11835 (N_11835,N_10193,N_10818);
nor U11836 (N_11836,N_10243,N_10394);
and U11837 (N_11837,N_10747,N_10040);
nor U11838 (N_11838,N_10136,N_10063);
nand U11839 (N_11839,N_10796,N_10946);
and U11840 (N_11840,N_10951,N_10642);
or U11841 (N_11841,N_10596,N_10142);
and U11842 (N_11842,N_10157,N_10314);
nor U11843 (N_11843,N_10888,N_10226);
nor U11844 (N_11844,N_10526,N_10181);
or U11845 (N_11845,N_10822,N_10245);
xor U11846 (N_11846,N_10002,N_10566);
xnor U11847 (N_11847,N_10669,N_10186);
nand U11848 (N_11848,N_10753,N_10078);
nor U11849 (N_11849,N_10708,N_10981);
xnor U11850 (N_11850,N_10750,N_10662);
and U11851 (N_11851,N_10289,N_10047);
nor U11852 (N_11852,N_10950,N_10296);
or U11853 (N_11853,N_10086,N_10649);
or U11854 (N_11854,N_10274,N_10832);
or U11855 (N_11855,N_10253,N_10474);
nand U11856 (N_11856,N_10467,N_10478);
nand U11857 (N_11857,N_10373,N_10635);
nor U11858 (N_11858,N_10841,N_10197);
nor U11859 (N_11859,N_10215,N_10480);
nand U11860 (N_11860,N_10344,N_10828);
nand U11861 (N_11861,N_10093,N_10749);
nand U11862 (N_11862,N_10532,N_10563);
and U11863 (N_11863,N_10868,N_10136);
or U11864 (N_11864,N_10298,N_10840);
or U11865 (N_11865,N_10448,N_10698);
and U11866 (N_11866,N_10095,N_10934);
or U11867 (N_11867,N_10986,N_10538);
xor U11868 (N_11868,N_10559,N_10212);
or U11869 (N_11869,N_10347,N_10308);
nor U11870 (N_11870,N_10375,N_10023);
nand U11871 (N_11871,N_10352,N_10318);
or U11872 (N_11872,N_10611,N_10906);
xor U11873 (N_11873,N_10477,N_10904);
xor U11874 (N_11874,N_10912,N_10996);
nand U11875 (N_11875,N_10225,N_10039);
and U11876 (N_11876,N_10047,N_10627);
xor U11877 (N_11877,N_10416,N_10261);
or U11878 (N_11878,N_10218,N_10969);
nor U11879 (N_11879,N_10296,N_10176);
or U11880 (N_11880,N_10851,N_10879);
or U11881 (N_11881,N_10258,N_10164);
and U11882 (N_11882,N_10602,N_10196);
nand U11883 (N_11883,N_10240,N_10540);
nand U11884 (N_11884,N_10868,N_10631);
xor U11885 (N_11885,N_10978,N_10945);
or U11886 (N_11886,N_10111,N_10795);
nor U11887 (N_11887,N_10709,N_10813);
xnor U11888 (N_11888,N_10366,N_10327);
xnor U11889 (N_11889,N_10596,N_10238);
nor U11890 (N_11890,N_10702,N_10844);
xor U11891 (N_11891,N_10279,N_10208);
or U11892 (N_11892,N_10267,N_10644);
and U11893 (N_11893,N_10329,N_10699);
nor U11894 (N_11894,N_10585,N_10069);
or U11895 (N_11895,N_10483,N_10352);
xnor U11896 (N_11896,N_10483,N_10864);
and U11897 (N_11897,N_10159,N_10044);
nor U11898 (N_11898,N_10423,N_10578);
nand U11899 (N_11899,N_10280,N_10299);
nand U11900 (N_11900,N_10032,N_10486);
nor U11901 (N_11901,N_10470,N_10622);
or U11902 (N_11902,N_10340,N_10533);
and U11903 (N_11903,N_10661,N_10325);
nand U11904 (N_11904,N_10890,N_10637);
and U11905 (N_11905,N_10620,N_10790);
nor U11906 (N_11906,N_10372,N_10579);
nand U11907 (N_11907,N_10718,N_10985);
nor U11908 (N_11908,N_10890,N_10908);
nor U11909 (N_11909,N_10201,N_10514);
nand U11910 (N_11910,N_10845,N_10480);
or U11911 (N_11911,N_10083,N_10703);
xnor U11912 (N_11912,N_10007,N_10846);
and U11913 (N_11913,N_10057,N_10912);
or U11914 (N_11914,N_10244,N_10386);
and U11915 (N_11915,N_10745,N_10975);
or U11916 (N_11916,N_10701,N_10244);
nor U11917 (N_11917,N_10208,N_10164);
xnor U11918 (N_11918,N_10168,N_10453);
and U11919 (N_11919,N_10289,N_10400);
and U11920 (N_11920,N_10999,N_10899);
and U11921 (N_11921,N_10316,N_10716);
nand U11922 (N_11922,N_10649,N_10327);
nor U11923 (N_11923,N_10753,N_10769);
nor U11924 (N_11924,N_10123,N_10545);
xor U11925 (N_11925,N_10365,N_10821);
nand U11926 (N_11926,N_10312,N_10228);
xor U11927 (N_11927,N_10079,N_10344);
and U11928 (N_11928,N_10553,N_10022);
nand U11929 (N_11929,N_10344,N_10147);
nand U11930 (N_11930,N_10262,N_10825);
nand U11931 (N_11931,N_10716,N_10515);
nand U11932 (N_11932,N_10551,N_10163);
and U11933 (N_11933,N_10652,N_10408);
or U11934 (N_11934,N_10889,N_10843);
and U11935 (N_11935,N_10873,N_10256);
or U11936 (N_11936,N_10838,N_10863);
nor U11937 (N_11937,N_10926,N_10808);
nor U11938 (N_11938,N_10431,N_10779);
or U11939 (N_11939,N_10642,N_10229);
nand U11940 (N_11940,N_10326,N_10195);
nor U11941 (N_11941,N_10521,N_10596);
and U11942 (N_11942,N_10820,N_10636);
xor U11943 (N_11943,N_10917,N_10815);
and U11944 (N_11944,N_10361,N_10514);
or U11945 (N_11945,N_10754,N_10180);
or U11946 (N_11946,N_10781,N_10314);
xor U11947 (N_11947,N_10648,N_10131);
xnor U11948 (N_11948,N_10721,N_10923);
nand U11949 (N_11949,N_10004,N_10482);
nor U11950 (N_11950,N_10303,N_10709);
xor U11951 (N_11951,N_10365,N_10595);
nor U11952 (N_11952,N_10316,N_10577);
or U11953 (N_11953,N_10372,N_10059);
or U11954 (N_11954,N_10670,N_10033);
and U11955 (N_11955,N_10051,N_10742);
nor U11956 (N_11956,N_10925,N_10541);
nand U11957 (N_11957,N_10022,N_10697);
or U11958 (N_11958,N_10859,N_10887);
and U11959 (N_11959,N_10902,N_10173);
xor U11960 (N_11960,N_10382,N_10266);
and U11961 (N_11961,N_10670,N_10272);
nor U11962 (N_11962,N_10217,N_10301);
or U11963 (N_11963,N_10831,N_10313);
xor U11964 (N_11964,N_10589,N_10259);
nand U11965 (N_11965,N_10734,N_10509);
or U11966 (N_11966,N_10039,N_10297);
or U11967 (N_11967,N_10815,N_10843);
xnor U11968 (N_11968,N_10017,N_10422);
and U11969 (N_11969,N_10765,N_10302);
nor U11970 (N_11970,N_10427,N_10736);
and U11971 (N_11971,N_10121,N_10890);
nand U11972 (N_11972,N_10743,N_10064);
and U11973 (N_11973,N_10630,N_10241);
nand U11974 (N_11974,N_10310,N_10534);
nor U11975 (N_11975,N_10813,N_10280);
and U11976 (N_11976,N_10566,N_10305);
nand U11977 (N_11977,N_10793,N_10792);
or U11978 (N_11978,N_10375,N_10798);
nor U11979 (N_11979,N_10775,N_10196);
xor U11980 (N_11980,N_10165,N_10760);
xor U11981 (N_11981,N_10131,N_10715);
or U11982 (N_11982,N_10857,N_10333);
nor U11983 (N_11983,N_10726,N_10584);
xor U11984 (N_11984,N_10283,N_10859);
or U11985 (N_11985,N_10958,N_10758);
xor U11986 (N_11986,N_10956,N_10754);
or U11987 (N_11987,N_10096,N_10075);
nor U11988 (N_11988,N_10057,N_10157);
or U11989 (N_11989,N_10276,N_10786);
and U11990 (N_11990,N_10487,N_10068);
or U11991 (N_11991,N_10482,N_10651);
and U11992 (N_11992,N_10608,N_10695);
or U11993 (N_11993,N_10296,N_10050);
nor U11994 (N_11994,N_10228,N_10265);
nor U11995 (N_11995,N_10630,N_10009);
xnor U11996 (N_11996,N_10911,N_10353);
nor U11997 (N_11997,N_10951,N_10897);
nand U11998 (N_11998,N_10632,N_10420);
and U11999 (N_11999,N_10081,N_10264);
nand U12000 (N_12000,N_11129,N_11516);
or U12001 (N_12001,N_11075,N_11130);
or U12002 (N_12002,N_11478,N_11855);
xor U12003 (N_12003,N_11676,N_11553);
nand U12004 (N_12004,N_11269,N_11037);
nor U12005 (N_12005,N_11459,N_11126);
or U12006 (N_12006,N_11860,N_11442);
xor U12007 (N_12007,N_11850,N_11343);
nand U12008 (N_12008,N_11755,N_11863);
nand U12009 (N_12009,N_11697,N_11226);
and U12010 (N_12010,N_11603,N_11042);
or U12011 (N_12011,N_11532,N_11745);
xnor U12012 (N_12012,N_11311,N_11172);
and U12013 (N_12013,N_11303,N_11752);
xor U12014 (N_12014,N_11403,N_11367);
nor U12015 (N_12015,N_11954,N_11901);
and U12016 (N_12016,N_11939,N_11610);
or U12017 (N_12017,N_11451,N_11812);
or U12018 (N_12018,N_11998,N_11094);
nor U12019 (N_12019,N_11982,N_11615);
and U12020 (N_12020,N_11190,N_11981);
nand U12021 (N_12021,N_11817,N_11972);
xor U12022 (N_12022,N_11043,N_11496);
nor U12023 (N_12023,N_11884,N_11647);
and U12024 (N_12024,N_11589,N_11994);
and U12025 (N_12025,N_11514,N_11853);
nor U12026 (N_12026,N_11717,N_11005);
or U12027 (N_12027,N_11929,N_11893);
xnor U12028 (N_12028,N_11027,N_11688);
and U12029 (N_12029,N_11297,N_11856);
nand U12030 (N_12030,N_11124,N_11656);
nor U12031 (N_12031,N_11405,N_11221);
nand U12032 (N_12032,N_11302,N_11063);
nor U12033 (N_12033,N_11571,N_11624);
nand U12034 (N_12034,N_11462,N_11675);
or U12035 (N_12035,N_11798,N_11248);
nand U12036 (N_12036,N_11527,N_11876);
and U12037 (N_12037,N_11799,N_11337);
nor U12038 (N_12038,N_11620,N_11086);
and U12039 (N_12039,N_11249,N_11274);
or U12040 (N_12040,N_11414,N_11825);
nand U12041 (N_12041,N_11788,N_11525);
nand U12042 (N_12042,N_11892,N_11563);
and U12043 (N_12043,N_11180,N_11120);
or U12044 (N_12044,N_11200,N_11066);
nor U12045 (N_12045,N_11704,N_11597);
nor U12046 (N_12046,N_11292,N_11594);
and U12047 (N_12047,N_11329,N_11957);
nand U12048 (N_12048,N_11699,N_11879);
nor U12049 (N_12049,N_11339,N_11573);
or U12050 (N_12050,N_11970,N_11355);
and U12051 (N_12051,N_11800,N_11847);
nand U12052 (N_12052,N_11239,N_11194);
nand U12053 (N_12053,N_11169,N_11690);
nor U12054 (N_12054,N_11109,N_11201);
xnor U12055 (N_12055,N_11542,N_11744);
or U12056 (N_12056,N_11902,N_11626);
xor U12057 (N_12057,N_11210,N_11684);
or U12058 (N_12058,N_11625,N_11472);
or U12059 (N_12059,N_11434,N_11653);
and U12060 (N_12060,N_11204,N_11071);
nor U12061 (N_12061,N_11164,N_11051);
and U12062 (N_12062,N_11568,N_11286);
nor U12063 (N_12063,N_11851,N_11163);
and U12064 (N_12064,N_11187,N_11826);
and U12065 (N_12065,N_11551,N_11554);
or U12066 (N_12066,N_11728,N_11609);
or U12067 (N_12067,N_11465,N_11041);
xnor U12068 (N_12068,N_11305,N_11531);
nor U12069 (N_12069,N_11395,N_11336);
nand U12070 (N_12070,N_11999,N_11724);
xnor U12071 (N_12071,N_11579,N_11830);
xnor U12072 (N_12072,N_11099,N_11016);
and U12073 (N_12073,N_11211,N_11369);
and U12074 (N_12074,N_11088,N_11389);
xnor U12075 (N_12075,N_11447,N_11679);
and U12076 (N_12076,N_11060,N_11736);
and U12077 (N_12077,N_11148,N_11548);
nand U12078 (N_12078,N_11661,N_11556);
xnor U12079 (N_12079,N_11960,N_11113);
nand U12080 (N_12080,N_11686,N_11701);
nand U12081 (N_12081,N_11273,N_11419);
nor U12082 (N_12082,N_11272,N_11374);
or U12083 (N_12083,N_11000,N_11522);
and U12084 (N_12084,N_11771,N_11185);
and U12085 (N_12085,N_11460,N_11836);
and U12086 (N_12086,N_11267,N_11456);
nor U12087 (N_12087,N_11485,N_11435);
nand U12088 (N_12088,N_11733,N_11175);
or U12089 (N_12089,N_11035,N_11543);
nor U12090 (N_12090,N_11645,N_11997);
or U12091 (N_12091,N_11846,N_11228);
and U12092 (N_12092,N_11199,N_11168);
or U12093 (N_12093,N_11885,N_11739);
and U12094 (N_12094,N_11810,N_11790);
or U12095 (N_12095,N_11268,N_11011);
nand U12096 (N_12096,N_11084,N_11772);
or U12097 (N_12097,N_11815,N_11494);
nand U12098 (N_12098,N_11700,N_11209);
nor U12099 (N_12099,N_11449,N_11783);
and U12100 (N_12100,N_11466,N_11651);
nor U12101 (N_12101,N_11087,N_11136);
or U12102 (N_12102,N_11284,N_11469);
and U12103 (N_12103,N_11608,N_11483);
or U12104 (N_12104,N_11153,N_11309);
xnor U12105 (N_12105,N_11991,N_11490);
and U12106 (N_12106,N_11517,N_11152);
or U12107 (N_12107,N_11980,N_11667);
nor U12108 (N_12108,N_11695,N_11895);
xnor U12109 (N_12109,N_11677,N_11476);
nor U12110 (N_12110,N_11920,N_11726);
xnor U12111 (N_12111,N_11513,N_11869);
and U12112 (N_12112,N_11505,N_11026);
or U12113 (N_12113,N_11425,N_11538);
xnor U12114 (N_12114,N_11370,N_11737);
nor U12115 (N_12115,N_11816,N_11600);
xor U12116 (N_12116,N_11452,N_11096);
and U12117 (N_12117,N_11471,N_11330);
or U12118 (N_12118,N_11931,N_11149);
or U12119 (N_12119,N_11844,N_11523);
xnor U12120 (N_12120,N_11227,N_11881);
nor U12121 (N_12121,N_11421,N_11214);
xor U12122 (N_12122,N_11952,N_11196);
nand U12123 (N_12123,N_11400,N_11009);
nor U12124 (N_12124,N_11019,N_11077);
nor U12125 (N_12125,N_11362,N_11720);
xnor U12126 (N_12126,N_11347,N_11417);
xnor U12127 (N_12127,N_11663,N_11807);
and U12128 (N_12128,N_11497,N_11680);
nand U12129 (N_12129,N_11006,N_11315);
nand U12130 (N_12130,N_11304,N_11660);
and U12131 (N_12131,N_11251,N_11698);
xnor U12132 (N_12132,N_11072,N_11528);
or U12133 (N_12133,N_11854,N_11406);
xnor U12134 (N_12134,N_11511,N_11154);
or U12135 (N_12135,N_11393,N_11743);
nor U12136 (N_12136,N_11257,N_11010);
and U12137 (N_12137,N_11662,N_11875);
nand U12138 (N_12138,N_11001,N_11508);
xnor U12139 (N_12139,N_11392,N_11404);
nor U12140 (N_12140,N_11433,N_11593);
nor U12141 (N_12141,N_11588,N_11263);
xnor U12142 (N_12142,N_11968,N_11391);
or U12143 (N_12143,N_11454,N_11029);
or U12144 (N_12144,N_11105,N_11107);
nor U12145 (N_12145,N_11580,N_11504);
xor U12146 (N_12146,N_11671,N_11344);
and U12147 (N_12147,N_11123,N_11186);
nand U12148 (N_12148,N_11503,N_11162);
nor U12149 (N_12149,N_11440,N_11781);
xnor U12150 (N_12150,N_11742,N_11232);
and U12151 (N_12151,N_11242,N_11722);
nor U12152 (N_12152,N_11572,N_11606);
or U12153 (N_12153,N_11636,N_11282);
nand U12154 (N_12154,N_11927,N_11719);
and U12155 (N_12155,N_11312,N_11888);
nor U12156 (N_12156,N_11054,N_11020);
nor U12157 (N_12157,N_11166,N_11890);
nor U12158 (N_12158,N_11611,N_11386);
or U12159 (N_12159,N_11539,N_11911);
or U12160 (N_12160,N_11486,N_11537);
or U12161 (N_12161,N_11794,N_11340);
nor U12162 (N_12162,N_11802,N_11371);
nor U12163 (N_12163,N_11703,N_11104);
and U12164 (N_12164,N_11484,N_11382);
xor U12165 (N_12165,N_11354,N_11838);
nor U12166 (N_12166,N_11253,N_11193);
and U12167 (N_12167,N_11837,N_11831);
nand U12168 (N_12168,N_11687,N_11682);
nor U12169 (N_12169,N_11683,N_11295);
xnor U12170 (N_12170,N_11331,N_11081);
or U12171 (N_12171,N_11482,N_11208);
nand U12172 (N_12172,N_11264,N_11373);
xnor U12173 (N_12173,N_11383,N_11832);
nand U12174 (N_12174,N_11155,N_11768);
xor U12175 (N_12175,N_11431,N_11657);
nand U12176 (N_12176,N_11381,N_11464);
xnor U12177 (N_12177,N_11849,N_11119);
and U12178 (N_12178,N_11550,N_11899);
nor U12179 (N_12179,N_11937,N_11649);
nor U12180 (N_12180,N_11940,N_11648);
nor U12181 (N_12181,N_11827,N_11873);
nor U12182 (N_12182,N_11028,N_11987);
xor U12183 (N_12183,N_11364,N_11147);
xnor U12184 (N_12184,N_11509,N_11764);
xor U12185 (N_12185,N_11599,N_11101);
and U12186 (N_12186,N_11506,N_11840);
and U12187 (N_12187,N_11806,N_11252);
and U12188 (N_12188,N_11157,N_11225);
xor U12189 (N_12189,N_11534,N_11928);
or U12190 (N_12190,N_11602,N_11595);
xor U12191 (N_12191,N_11629,N_11756);
xor U12192 (N_12192,N_11188,N_11965);
nand U12193 (N_12193,N_11322,N_11352);
nor U12194 (N_12194,N_11487,N_11491);
and U12195 (N_12195,N_11641,N_11250);
or U12196 (N_12196,N_11023,N_11566);
or U12197 (N_12197,N_11444,N_11897);
xnor U12198 (N_12198,N_11365,N_11195);
nor U12199 (N_12199,N_11247,N_11921);
nor U12200 (N_12200,N_11917,N_11357);
nor U12201 (N_12201,N_11933,N_11499);
xor U12202 (N_12202,N_11488,N_11289);
xor U12203 (N_12203,N_11740,N_11407);
and U12204 (N_12204,N_11241,N_11926);
or U12205 (N_12205,N_11642,N_11622);
xor U12206 (N_12206,N_11723,N_11256);
nor U12207 (N_12207,N_11243,N_11658);
and U12208 (N_12208,N_11942,N_11628);
or U12209 (N_12209,N_11839,N_11348);
xor U12210 (N_12210,N_11995,N_11245);
nand U12211 (N_12211,N_11230,N_11576);
nand U12212 (N_12212,N_11045,N_11067);
and U12213 (N_12213,N_11215,N_11592);
nand U12214 (N_12214,N_11894,N_11567);
nor U12215 (N_12215,N_11399,N_11824);
or U12216 (N_12216,N_11852,N_11012);
and U12217 (N_12217,N_11036,N_11307);
nand U12218 (N_12218,N_11223,N_11398);
and U12219 (N_12219,N_11396,N_11368);
nor U12220 (N_12220,N_11668,N_11716);
or U12221 (N_12221,N_11092,N_11052);
nand U12222 (N_12222,N_11335,N_11582);
or U12223 (N_12223,N_11025,N_11774);
and U12224 (N_12224,N_11468,N_11782);
nand U12225 (N_12225,N_11570,N_11547);
or U12226 (N_12226,N_11654,N_11578);
and U12227 (N_12227,N_11021,N_11596);
nand U12228 (N_12228,N_11453,N_11377);
or U12229 (N_12229,N_11958,N_11590);
and U12230 (N_12230,N_11685,N_11565);
xor U12231 (N_12231,N_11637,N_11635);
or U12232 (N_12232,N_11546,N_11627);
and U12233 (N_12233,N_11358,N_11941);
xnor U12234 (N_12234,N_11379,N_11325);
nand U12235 (N_12235,N_11412,N_11115);
xnor U12236 (N_12236,N_11874,N_11181);
or U12237 (N_12237,N_11681,N_11731);
xor U12238 (N_12238,N_11032,N_11923);
xnor U12239 (N_12239,N_11171,N_11050);
nor U12240 (N_12240,N_11353,N_11135);
nor U12241 (N_12241,N_11288,N_11324);
or U12242 (N_12242,N_11192,N_11328);
nor U12243 (N_12243,N_11944,N_11977);
or U12244 (N_12244,N_11296,N_11408);
nand U12245 (N_12245,N_11865,N_11828);
xor U12246 (N_12246,N_11301,N_11143);
xnor U12247 (N_12247,N_11841,N_11061);
xnor U12248 (N_12248,N_11366,N_11934);
or U12249 (N_12249,N_11448,N_11438);
xnor U12250 (N_12250,N_11420,N_11604);
nor U12251 (N_12251,N_11633,N_11882);
nor U12252 (N_12252,N_11235,N_11631);
or U12253 (N_12253,N_11858,N_11132);
nor U12254 (N_12254,N_11038,N_11614);
nor U12255 (N_12255,N_11057,N_11378);
nand U12256 (N_12256,N_11935,N_11512);
nor U12257 (N_12257,N_11446,N_11947);
nor U12258 (N_12258,N_11963,N_11692);
nor U12259 (N_12259,N_11411,N_11632);
nor U12260 (N_12260,N_11983,N_11138);
xor U12261 (N_12261,N_11308,N_11334);
or U12262 (N_12262,N_11317,N_11813);
and U12263 (N_12263,N_11384,N_11691);
nor U12264 (N_12264,N_11880,N_11765);
nor U12265 (N_12265,N_11069,N_11259);
xnor U12266 (N_12266,N_11584,N_11822);
and U12267 (N_12267,N_11280,N_11422);
nand U12268 (N_12268,N_11988,N_11212);
nand U12269 (N_12269,N_11178,N_11443);
xnor U12270 (N_12270,N_11644,N_11867);
or U12271 (N_12271,N_11290,N_11146);
nand U12272 (N_12272,N_11961,N_11461);
xor U12273 (N_12273,N_11909,N_11956);
nor U12274 (N_12274,N_11903,N_11607);
nor U12275 (N_12275,N_11473,N_11093);
xnor U12276 (N_12276,N_11238,N_11122);
and U12277 (N_12277,N_11213,N_11749);
xor U12278 (N_12278,N_11350,N_11445);
nand U12279 (N_12279,N_11993,N_11669);
or U12280 (N_12280,N_11761,N_11613);
xor U12281 (N_12281,N_11616,N_11712);
and U12282 (N_12282,N_11179,N_11202);
or U12283 (N_12283,N_11076,N_11246);
or U12284 (N_12284,N_11889,N_11634);
or U12285 (N_12285,N_11801,N_11121);
or U12286 (N_12286,N_11769,N_11160);
nand U12287 (N_12287,N_11834,N_11507);
xor U12288 (N_12288,N_11829,N_11887);
or U12289 (N_12289,N_11912,N_11316);
and U12290 (N_12290,N_11457,N_11919);
or U12291 (N_12291,N_11427,N_11332);
nand U12292 (N_12292,N_11306,N_11821);
xnor U12293 (N_12293,N_11666,N_11714);
nand U12294 (N_12294,N_11763,N_11004);
and U12295 (N_12295,N_11612,N_11564);
or U12296 (N_12296,N_11085,N_11672);
nand U12297 (N_12297,N_11842,N_11321);
or U12298 (N_12298,N_11776,N_11702);
nor U12299 (N_12299,N_11750,N_11024);
and U12300 (N_12300,N_11283,N_11189);
xor U12301 (N_12301,N_11299,N_11727);
nor U12302 (N_12302,N_11401,N_11966);
nand U12303 (N_12303,N_11730,N_11904);
xnor U12304 (N_12304,N_11244,N_11964);
xnor U12305 (N_12305,N_11916,N_11500);
or U12306 (N_12306,N_11165,N_11918);
or U12307 (N_12307,N_11835,N_11342);
xnor U12308 (N_12308,N_11985,N_11818);
nor U12309 (N_12309,N_11955,N_11470);
xor U12310 (N_12310,N_11128,N_11530);
or U12311 (N_12311,N_11255,N_11493);
nand U12312 (N_12312,N_11779,N_11770);
nor U12313 (N_12313,N_11229,N_11319);
or U12314 (N_12314,N_11519,N_11545);
xnor U12315 (N_12315,N_11158,N_11533);
or U12316 (N_12316,N_11049,N_11536);
and U12317 (N_12317,N_11693,N_11689);
and U12318 (N_12318,N_11561,N_11930);
and U12319 (N_12319,N_11003,N_11759);
nand U12320 (N_12320,N_11510,N_11908);
or U12321 (N_12321,N_11065,N_11097);
and U12322 (N_12322,N_11915,N_11207);
and U12323 (N_12323,N_11797,N_11619);
and U12324 (N_12324,N_11924,N_11481);
nand U12325 (N_12325,N_11706,N_11914);
nand U12326 (N_12326,N_11555,N_11872);
nor U12327 (N_12327,N_11540,N_11804);
xnor U12328 (N_12328,N_11796,N_11070);
xor U12329 (N_12329,N_11116,N_11809);
and U12330 (N_12330,N_11013,N_11721);
nand U12331 (N_12331,N_11455,N_11877);
or U12332 (N_12332,N_11646,N_11142);
or U12333 (N_12333,N_11559,N_11137);
or U12334 (N_12334,N_11007,N_11711);
or U12335 (N_12335,N_11823,N_11948);
or U12336 (N_12336,N_11707,N_11959);
nor U12337 (N_12337,N_11098,N_11359);
or U12338 (N_12338,N_11375,N_11746);
or U12339 (N_12339,N_11710,N_11762);
and U12340 (N_12340,N_11962,N_11870);
and U12341 (N_12341,N_11022,N_11975);
and U12342 (N_12342,N_11217,N_11585);
nand U12343 (N_12343,N_11133,N_11141);
and U12344 (N_12344,N_11281,N_11574);
nor U12345 (N_12345,N_11333,N_11151);
nor U12346 (N_12346,N_11062,N_11978);
xnor U12347 (N_12347,N_11089,N_11265);
xor U12348 (N_12348,N_11713,N_11953);
xor U12349 (N_12349,N_11560,N_11734);
or U12350 (N_12350,N_11039,N_11118);
or U12351 (N_12351,N_11033,N_11441);
and U12352 (N_12352,N_11906,N_11183);
nor U12353 (N_12353,N_11047,N_11277);
nor U12354 (N_12354,N_11976,N_11883);
nand U12355 (N_12355,N_11520,N_11426);
nor U12356 (N_12356,N_11951,N_11467);
or U12357 (N_12357,N_11878,N_11480);
nor U12358 (N_12358,N_11886,N_11967);
or U12359 (N_12359,N_11298,N_11111);
nand U12360 (N_12360,N_11327,N_11515);
xor U12361 (N_12361,N_11205,N_11413);
nor U12362 (N_12362,N_11673,N_11640);
or U12363 (N_12363,N_11623,N_11231);
and U12364 (N_12364,N_11345,N_11639);
nor U12365 (N_12365,N_11173,N_11795);
and U12366 (N_12366,N_11018,N_11715);
nand U12367 (N_12367,N_11275,N_11936);
or U12368 (N_12368,N_11326,N_11380);
nor U12369 (N_12369,N_11767,N_11922);
and U12370 (N_12370,N_11078,N_11258);
nor U12371 (N_12371,N_11150,N_11385);
nand U12372 (N_12372,N_11650,N_11017);
or U12373 (N_12373,N_11198,N_11862);
or U12374 (N_12374,N_11262,N_11819);
and U12375 (N_12375,N_11415,N_11361);
or U12376 (N_12376,N_11387,N_11323);
nor U12377 (N_12377,N_11581,N_11575);
and U12378 (N_12378,N_11074,N_11705);
xor U12379 (N_12379,N_11738,N_11786);
nand U12380 (N_12380,N_11346,N_11741);
nand U12381 (N_12381,N_11652,N_11820);
and U12382 (N_12382,N_11068,N_11859);
nand U12383 (N_12383,N_11064,N_11218);
or U12384 (N_12384,N_11182,N_11562);
nor U12385 (N_12385,N_11845,N_11605);
and U12386 (N_12386,N_11040,N_11044);
xnor U12387 (N_12387,N_11814,N_11144);
and U12388 (N_12388,N_11110,N_11524);
nor U12389 (N_12389,N_11974,N_11095);
nor U12390 (N_12390,N_11754,N_11082);
and U12391 (N_12391,N_11056,N_11176);
xor U12392 (N_12392,N_11618,N_11973);
and U12393 (N_12393,N_11678,N_11117);
nor U12394 (N_12394,N_11843,N_11785);
xor U12395 (N_12395,N_11898,N_11766);
nand U12396 (N_12396,N_11501,N_11423);
and U12397 (N_12397,N_11100,N_11191);
and U12398 (N_12398,N_11475,N_11233);
xor U12399 (N_12399,N_11803,N_11287);
or U12400 (N_12400,N_11015,N_11552);
and U12401 (N_12401,N_11224,N_11418);
xor U12402 (N_12402,N_11780,N_11986);
or U12403 (N_12403,N_11913,N_11156);
nor U12404 (N_12404,N_11694,N_11479);
nand U12405 (N_12405,N_11108,N_11293);
nor U12406 (N_12406,N_11773,N_11161);
xnor U12407 (N_12407,N_11046,N_11285);
nor U12408 (N_12408,N_11477,N_11617);
xnor U12409 (N_12409,N_11261,N_11318);
and U12410 (N_12410,N_11439,N_11432);
nand U12411 (N_12411,N_11777,N_11498);
and U12412 (N_12412,N_11989,N_11871);
xnor U12413 (N_12413,N_11320,N_11397);
nand U12414 (N_12414,N_11159,N_11197);
nand U12415 (N_12415,N_11518,N_11131);
nor U12416 (N_12416,N_11925,N_11557);
nand U12417 (N_12417,N_11753,N_11276);
or U12418 (N_12418,N_11106,N_11577);
or U12419 (N_12419,N_11938,N_11943);
or U12420 (N_12420,N_11670,N_11450);
and U12421 (N_12421,N_11140,N_11410);
nor U12422 (N_12422,N_11271,N_11778);
xor U12423 (N_12423,N_11436,N_11177);
and U12424 (N_12424,N_11219,N_11260);
nor U12425 (N_12425,N_11489,N_11145);
and U12426 (N_12426,N_11655,N_11587);
or U12427 (N_12427,N_11349,N_11216);
xor U12428 (N_12428,N_11080,N_11059);
nor U12429 (N_12429,N_11313,N_11808);
or U12430 (N_12430,N_11971,N_11748);
nor U12431 (N_12431,N_11341,N_11583);
nand U12432 (N_12432,N_11718,N_11792);
xor U12433 (N_12433,N_11053,N_11206);
xnor U12434 (N_12434,N_11170,N_11729);
nor U12435 (N_12435,N_11279,N_11868);
nor U12436 (N_12436,N_11979,N_11758);
or U12437 (N_12437,N_11725,N_11709);
or U12438 (N_12438,N_11234,N_11791);
or U12439 (N_12439,N_11114,N_11946);
nand U12440 (N_12440,N_11945,N_11861);
or U12441 (N_12441,N_11664,N_11760);
xnor U12442 (N_12442,N_11428,N_11236);
nor U12443 (N_12443,N_11103,N_11388);
and U12444 (N_12444,N_11437,N_11220);
and U12445 (N_12445,N_11900,N_11787);
and U12446 (N_12446,N_11789,N_11544);
and U12447 (N_12447,N_11659,N_11372);
xnor U12448 (N_12448,N_11310,N_11351);
nor U12449 (N_12449,N_11932,N_11905);
nor U12450 (N_12450,N_11237,N_11030);
nor U12451 (N_12451,N_11811,N_11424);
and U12452 (N_12452,N_11535,N_11643);
or U12453 (N_12453,N_11360,N_11990);
nor U12454 (N_12454,N_11134,N_11356);
xnor U12455 (N_12455,N_11254,N_11112);
nand U12456 (N_12456,N_11586,N_11757);
and U12457 (N_12457,N_11996,N_11300);
and U12458 (N_12458,N_11031,N_11314);
xnor U12459 (N_12459,N_11866,N_11429);
nor U12460 (N_12460,N_11984,N_11907);
nand U12461 (N_12461,N_11492,N_11708);
nor U12462 (N_12462,N_11394,N_11058);
and U12463 (N_12463,N_11203,N_11569);
or U12464 (N_12464,N_11174,N_11992);
nor U12465 (N_12465,N_11002,N_11784);
nand U12466 (N_12466,N_11674,N_11950);
xor U12467 (N_12467,N_11240,N_11558);
nand U12468 (N_12468,N_11184,N_11591);
nand U12469 (N_12469,N_11896,N_11949);
and U12470 (N_12470,N_11598,N_11458);
nor U12471 (N_12471,N_11665,N_11502);
or U12472 (N_12472,N_11735,N_11864);
xor U12473 (N_12473,N_11696,N_11541);
xor U12474 (N_12474,N_11222,N_11601);
and U12475 (N_12475,N_11747,N_11416);
xor U12476 (N_12476,N_11521,N_11008);
and U12477 (N_12477,N_11083,N_11529);
nand U12478 (N_12478,N_11751,N_11430);
nand U12479 (N_12479,N_11402,N_11891);
and U12480 (N_12480,N_11055,N_11549);
or U12481 (N_12481,N_11526,N_11630);
and U12482 (N_12482,N_11775,N_11073);
and U12483 (N_12483,N_11266,N_11390);
or U12484 (N_12484,N_11167,N_11376);
nor U12485 (N_12485,N_11409,N_11034);
nand U12486 (N_12486,N_11732,N_11969);
xor U12487 (N_12487,N_11495,N_11833);
or U12488 (N_12488,N_11014,N_11291);
or U12489 (N_12489,N_11910,N_11102);
and U12490 (N_12490,N_11270,N_11848);
and U12491 (N_12491,N_11048,N_11857);
nand U12492 (N_12492,N_11474,N_11638);
and U12493 (N_12493,N_11793,N_11805);
xnor U12494 (N_12494,N_11139,N_11338);
and U12495 (N_12495,N_11125,N_11363);
nand U12496 (N_12496,N_11621,N_11294);
and U12497 (N_12497,N_11091,N_11127);
nand U12498 (N_12498,N_11463,N_11090);
nor U12499 (N_12499,N_11079,N_11278);
nand U12500 (N_12500,N_11329,N_11287);
xnor U12501 (N_12501,N_11588,N_11624);
nor U12502 (N_12502,N_11917,N_11963);
or U12503 (N_12503,N_11853,N_11960);
xnor U12504 (N_12504,N_11583,N_11429);
or U12505 (N_12505,N_11551,N_11409);
and U12506 (N_12506,N_11197,N_11368);
nor U12507 (N_12507,N_11690,N_11119);
xnor U12508 (N_12508,N_11341,N_11962);
nand U12509 (N_12509,N_11291,N_11123);
nand U12510 (N_12510,N_11389,N_11298);
nand U12511 (N_12511,N_11081,N_11366);
nand U12512 (N_12512,N_11192,N_11904);
or U12513 (N_12513,N_11537,N_11748);
and U12514 (N_12514,N_11833,N_11658);
or U12515 (N_12515,N_11645,N_11382);
or U12516 (N_12516,N_11467,N_11087);
or U12517 (N_12517,N_11786,N_11029);
or U12518 (N_12518,N_11216,N_11695);
xor U12519 (N_12519,N_11388,N_11891);
nor U12520 (N_12520,N_11491,N_11070);
nand U12521 (N_12521,N_11315,N_11439);
and U12522 (N_12522,N_11057,N_11570);
xnor U12523 (N_12523,N_11151,N_11423);
or U12524 (N_12524,N_11223,N_11517);
nor U12525 (N_12525,N_11214,N_11043);
or U12526 (N_12526,N_11663,N_11548);
and U12527 (N_12527,N_11982,N_11292);
nor U12528 (N_12528,N_11748,N_11272);
nand U12529 (N_12529,N_11443,N_11495);
nand U12530 (N_12530,N_11636,N_11081);
and U12531 (N_12531,N_11924,N_11454);
nand U12532 (N_12532,N_11657,N_11180);
or U12533 (N_12533,N_11429,N_11257);
nor U12534 (N_12534,N_11896,N_11922);
or U12535 (N_12535,N_11565,N_11166);
xnor U12536 (N_12536,N_11840,N_11601);
nor U12537 (N_12537,N_11927,N_11511);
nand U12538 (N_12538,N_11266,N_11226);
xor U12539 (N_12539,N_11805,N_11235);
and U12540 (N_12540,N_11357,N_11330);
nand U12541 (N_12541,N_11027,N_11524);
nor U12542 (N_12542,N_11496,N_11162);
nand U12543 (N_12543,N_11893,N_11102);
nor U12544 (N_12544,N_11107,N_11993);
xor U12545 (N_12545,N_11411,N_11795);
nor U12546 (N_12546,N_11971,N_11099);
and U12547 (N_12547,N_11342,N_11055);
and U12548 (N_12548,N_11246,N_11534);
nor U12549 (N_12549,N_11551,N_11720);
nor U12550 (N_12550,N_11221,N_11380);
and U12551 (N_12551,N_11016,N_11836);
nand U12552 (N_12552,N_11854,N_11709);
nor U12553 (N_12553,N_11653,N_11494);
or U12554 (N_12554,N_11634,N_11045);
and U12555 (N_12555,N_11243,N_11381);
or U12556 (N_12556,N_11531,N_11775);
nor U12557 (N_12557,N_11047,N_11029);
and U12558 (N_12558,N_11241,N_11956);
xor U12559 (N_12559,N_11263,N_11165);
nand U12560 (N_12560,N_11101,N_11216);
xnor U12561 (N_12561,N_11621,N_11626);
nor U12562 (N_12562,N_11969,N_11235);
nand U12563 (N_12563,N_11186,N_11156);
nor U12564 (N_12564,N_11470,N_11743);
xnor U12565 (N_12565,N_11033,N_11161);
or U12566 (N_12566,N_11546,N_11047);
xor U12567 (N_12567,N_11821,N_11814);
or U12568 (N_12568,N_11464,N_11319);
and U12569 (N_12569,N_11225,N_11198);
or U12570 (N_12570,N_11926,N_11574);
nand U12571 (N_12571,N_11086,N_11636);
nand U12572 (N_12572,N_11968,N_11467);
and U12573 (N_12573,N_11647,N_11872);
xor U12574 (N_12574,N_11488,N_11011);
nor U12575 (N_12575,N_11982,N_11414);
xnor U12576 (N_12576,N_11051,N_11121);
and U12577 (N_12577,N_11187,N_11658);
xor U12578 (N_12578,N_11352,N_11789);
and U12579 (N_12579,N_11083,N_11595);
or U12580 (N_12580,N_11794,N_11290);
xor U12581 (N_12581,N_11300,N_11218);
nand U12582 (N_12582,N_11878,N_11919);
or U12583 (N_12583,N_11967,N_11064);
nand U12584 (N_12584,N_11183,N_11281);
nand U12585 (N_12585,N_11628,N_11490);
and U12586 (N_12586,N_11685,N_11345);
or U12587 (N_12587,N_11056,N_11266);
or U12588 (N_12588,N_11923,N_11294);
nor U12589 (N_12589,N_11197,N_11370);
xor U12590 (N_12590,N_11080,N_11471);
xor U12591 (N_12591,N_11808,N_11141);
nand U12592 (N_12592,N_11494,N_11846);
xnor U12593 (N_12593,N_11404,N_11734);
xnor U12594 (N_12594,N_11982,N_11694);
and U12595 (N_12595,N_11318,N_11526);
xnor U12596 (N_12596,N_11227,N_11840);
nor U12597 (N_12597,N_11825,N_11123);
or U12598 (N_12598,N_11861,N_11969);
nor U12599 (N_12599,N_11508,N_11493);
nor U12600 (N_12600,N_11837,N_11833);
nand U12601 (N_12601,N_11426,N_11026);
xor U12602 (N_12602,N_11294,N_11018);
nand U12603 (N_12603,N_11056,N_11587);
or U12604 (N_12604,N_11775,N_11277);
or U12605 (N_12605,N_11637,N_11684);
nand U12606 (N_12606,N_11164,N_11711);
or U12607 (N_12607,N_11035,N_11347);
nand U12608 (N_12608,N_11841,N_11937);
nor U12609 (N_12609,N_11561,N_11871);
xor U12610 (N_12610,N_11057,N_11636);
xnor U12611 (N_12611,N_11375,N_11126);
nand U12612 (N_12612,N_11203,N_11373);
xor U12613 (N_12613,N_11647,N_11098);
xor U12614 (N_12614,N_11577,N_11764);
and U12615 (N_12615,N_11519,N_11707);
xor U12616 (N_12616,N_11869,N_11321);
nand U12617 (N_12617,N_11513,N_11054);
nor U12618 (N_12618,N_11140,N_11340);
xnor U12619 (N_12619,N_11116,N_11011);
nand U12620 (N_12620,N_11800,N_11382);
nand U12621 (N_12621,N_11006,N_11317);
and U12622 (N_12622,N_11012,N_11843);
and U12623 (N_12623,N_11583,N_11008);
and U12624 (N_12624,N_11557,N_11885);
and U12625 (N_12625,N_11370,N_11435);
nand U12626 (N_12626,N_11273,N_11705);
and U12627 (N_12627,N_11496,N_11748);
xnor U12628 (N_12628,N_11927,N_11696);
nand U12629 (N_12629,N_11036,N_11206);
and U12630 (N_12630,N_11823,N_11543);
nand U12631 (N_12631,N_11868,N_11382);
and U12632 (N_12632,N_11135,N_11122);
nand U12633 (N_12633,N_11711,N_11689);
xnor U12634 (N_12634,N_11009,N_11100);
or U12635 (N_12635,N_11958,N_11348);
or U12636 (N_12636,N_11529,N_11036);
nand U12637 (N_12637,N_11556,N_11537);
nand U12638 (N_12638,N_11492,N_11235);
xnor U12639 (N_12639,N_11135,N_11169);
xnor U12640 (N_12640,N_11276,N_11919);
and U12641 (N_12641,N_11170,N_11399);
nand U12642 (N_12642,N_11598,N_11068);
and U12643 (N_12643,N_11733,N_11263);
nor U12644 (N_12644,N_11036,N_11383);
nor U12645 (N_12645,N_11626,N_11020);
and U12646 (N_12646,N_11368,N_11829);
or U12647 (N_12647,N_11304,N_11281);
xnor U12648 (N_12648,N_11442,N_11491);
nor U12649 (N_12649,N_11114,N_11792);
or U12650 (N_12650,N_11335,N_11883);
xnor U12651 (N_12651,N_11071,N_11915);
or U12652 (N_12652,N_11522,N_11327);
nand U12653 (N_12653,N_11026,N_11039);
or U12654 (N_12654,N_11565,N_11190);
nor U12655 (N_12655,N_11538,N_11273);
or U12656 (N_12656,N_11847,N_11253);
xor U12657 (N_12657,N_11549,N_11081);
nor U12658 (N_12658,N_11794,N_11639);
or U12659 (N_12659,N_11943,N_11862);
xor U12660 (N_12660,N_11201,N_11525);
or U12661 (N_12661,N_11065,N_11200);
xnor U12662 (N_12662,N_11504,N_11015);
nor U12663 (N_12663,N_11805,N_11607);
nand U12664 (N_12664,N_11711,N_11666);
nand U12665 (N_12665,N_11909,N_11642);
nand U12666 (N_12666,N_11106,N_11365);
or U12667 (N_12667,N_11655,N_11241);
and U12668 (N_12668,N_11262,N_11471);
nand U12669 (N_12669,N_11346,N_11946);
nor U12670 (N_12670,N_11263,N_11911);
xor U12671 (N_12671,N_11154,N_11482);
nand U12672 (N_12672,N_11505,N_11352);
nand U12673 (N_12673,N_11699,N_11587);
xor U12674 (N_12674,N_11314,N_11778);
nor U12675 (N_12675,N_11045,N_11883);
nor U12676 (N_12676,N_11351,N_11158);
nor U12677 (N_12677,N_11622,N_11102);
and U12678 (N_12678,N_11895,N_11722);
nand U12679 (N_12679,N_11852,N_11754);
or U12680 (N_12680,N_11475,N_11323);
nand U12681 (N_12681,N_11802,N_11524);
or U12682 (N_12682,N_11879,N_11323);
xor U12683 (N_12683,N_11311,N_11048);
nand U12684 (N_12684,N_11624,N_11094);
xnor U12685 (N_12685,N_11393,N_11689);
and U12686 (N_12686,N_11187,N_11162);
xor U12687 (N_12687,N_11458,N_11234);
xnor U12688 (N_12688,N_11747,N_11120);
or U12689 (N_12689,N_11355,N_11863);
and U12690 (N_12690,N_11813,N_11756);
nor U12691 (N_12691,N_11668,N_11502);
xnor U12692 (N_12692,N_11883,N_11842);
xnor U12693 (N_12693,N_11396,N_11336);
nor U12694 (N_12694,N_11896,N_11493);
nor U12695 (N_12695,N_11430,N_11550);
and U12696 (N_12696,N_11261,N_11002);
nor U12697 (N_12697,N_11570,N_11111);
and U12698 (N_12698,N_11679,N_11487);
and U12699 (N_12699,N_11083,N_11834);
xnor U12700 (N_12700,N_11304,N_11432);
nand U12701 (N_12701,N_11573,N_11910);
xor U12702 (N_12702,N_11974,N_11273);
nor U12703 (N_12703,N_11288,N_11260);
and U12704 (N_12704,N_11109,N_11403);
and U12705 (N_12705,N_11895,N_11803);
xnor U12706 (N_12706,N_11024,N_11194);
or U12707 (N_12707,N_11905,N_11460);
or U12708 (N_12708,N_11284,N_11350);
xor U12709 (N_12709,N_11831,N_11688);
and U12710 (N_12710,N_11176,N_11283);
nand U12711 (N_12711,N_11705,N_11528);
nand U12712 (N_12712,N_11267,N_11808);
or U12713 (N_12713,N_11789,N_11585);
nor U12714 (N_12714,N_11440,N_11587);
xor U12715 (N_12715,N_11662,N_11162);
or U12716 (N_12716,N_11977,N_11913);
nor U12717 (N_12717,N_11117,N_11748);
xnor U12718 (N_12718,N_11056,N_11876);
nor U12719 (N_12719,N_11749,N_11947);
and U12720 (N_12720,N_11767,N_11747);
nor U12721 (N_12721,N_11103,N_11738);
nor U12722 (N_12722,N_11127,N_11986);
nor U12723 (N_12723,N_11824,N_11531);
or U12724 (N_12724,N_11743,N_11827);
xnor U12725 (N_12725,N_11397,N_11470);
xor U12726 (N_12726,N_11041,N_11806);
or U12727 (N_12727,N_11830,N_11994);
xor U12728 (N_12728,N_11025,N_11885);
and U12729 (N_12729,N_11963,N_11166);
xnor U12730 (N_12730,N_11447,N_11987);
nand U12731 (N_12731,N_11516,N_11476);
and U12732 (N_12732,N_11099,N_11659);
nand U12733 (N_12733,N_11206,N_11417);
or U12734 (N_12734,N_11445,N_11582);
nor U12735 (N_12735,N_11671,N_11210);
or U12736 (N_12736,N_11920,N_11916);
nor U12737 (N_12737,N_11149,N_11721);
nand U12738 (N_12738,N_11941,N_11142);
nor U12739 (N_12739,N_11780,N_11111);
nor U12740 (N_12740,N_11698,N_11396);
or U12741 (N_12741,N_11752,N_11401);
and U12742 (N_12742,N_11338,N_11913);
xor U12743 (N_12743,N_11593,N_11173);
xor U12744 (N_12744,N_11845,N_11161);
nor U12745 (N_12745,N_11371,N_11093);
nand U12746 (N_12746,N_11320,N_11841);
or U12747 (N_12747,N_11213,N_11984);
nor U12748 (N_12748,N_11494,N_11949);
nor U12749 (N_12749,N_11134,N_11142);
or U12750 (N_12750,N_11591,N_11508);
xor U12751 (N_12751,N_11432,N_11231);
or U12752 (N_12752,N_11536,N_11662);
nand U12753 (N_12753,N_11622,N_11411);
and U12754 (N_12754,N_11414,N_11467);
nand U12755 (N_12755,N_11191,N_11810);
or U12756 (N_12756,N_11380,N_11546);
xnor U12757 (N_12757,N_11300,N_11049);
nor U12758 (N_12758,N_11459,N_11299);
nand U12759 (N_12759,N_11258,N_11625);
xnor U12760 (N_12760,N_11781,N_11444);
or U12761 (N_12761,N_11288,N_11274);
xor U12762 (N_12762,N_11948,N_11834);
nand U12763 (N_12763,N_11813,N_11931);
and U12764 (N_12764,N_11383,N_11087);
nor U12765 (N_12765,N_11886,N_11725);
xnor U12766 (N_12766,N_11186,N_11686);
or U12767 (N_12767,N_11580,N_11994);
nand U12768 (N_12768,N_11981,N_11069);
xor U12769 (N_12769,N_11633,N_11893);
xnor U12770 (N_12770,N_11603,N_11969);
and U12771 (N_12771,N_11334,N_11170);
nand U12772 (N_12772,N_11185,N_11555);
nor U12773 (N_12773,N_11649,N_11986);
or U12774 (N_12774,N_11034,N_11003);
nor U12775 (N_12775,N_11546,N_11175);
and U12776 (N_12776,N_11874,N_11524);
xor U12777 (N_12777,N_11385,N_11425);
nand U12778 (N_12778,N_11565,N_11039);
nor U12779 (N_12779,N_11140,N_11968);
nand U12780 (N_12780,N_11778,N_11888);
and U12781 (N_12781,N_11186,N_11912);
nor U12782 (N_12782,N_11896,N_11406);
or U12783 (N_12783,N_11477,N_11096);
nand U12784 (N_12784,N_11451,N_11897);
and U12785 (N_12785,N_11842,N_11149);
and U12786 (N_12786,N_11173,N_11110);
xnor U12787 (N_12787,N_11124,N_11706);
xnor U12788 (N_12788,N_11517,N_11673);
xor U12789 (N_12789,N_11661,N_11891);
and U12790 (N_12790,N_11996,N_11016);
nand U12791 (N_12791,N_11170,N_11074);
and U12792 (N_12792,N_11076,N_11548);
xor U12793 (N_12793,N_11313,N_11855);
nor U12794 (N_12794,N_11211,N_11443);
and U12795 (N_12795,N_11289,N_11002);
and U12796 (N_12796,N_11379,N_11351);
nand U12797 (N_12797,N_11361,N_11421);
nand U12798 (N_12798,N_11148,N_11542);
and U12799 (N_12799,N_11691,N_11047);
xor U12800 (N_12800,N_11927,N_11556);
xnor U12801 (N_12801,N_11077,N_11251);
or U12802 (N_12802,N_11671,N_11118);
nor U12803 (N_12803,N_11697,N_11688);
nand U12804 (N_12804,N_11733,N_11034);
nor U12805 (N_12805,N_11751,N_11339);
or U12806 (N_12806,N_11551,N_11107);
xor U12807 (N_12807,N_11105,N_11829);
nor U12808 (N_12808,N_11856,N_11009);
or U12809 (N_12809,N_11251,N_11646);
nand U12810 (N_12810,N_11534,N_11999);
xor U12811 (N_12811,N_11376,N_11236);
or U12812 (N_12812,N_11745,N_11381);
or U12813 (N_12813,N_11632,N_11448);
nand U12814 (N_12814,N_11144,N_11669);
nor U12815 (N_12815,N_11222,N_11132);
nor U12816 (N_12816,N_11726,N_11244);
or U12817 (N_12817,N_11226,N_11950);
or U12818 (N_12818,N_11843,N_11735);
xnor U12819 (N_12819,N_11034,N_11934);
xor U12820 (N_12820,N_11340,N_11824);
xnor U12821 (N_12821,N_11004,N_11103);
or U12822 (N_12822,N_11060,N_11549);
xnor U12823 (N_12823,N_11232,N_11365);
nand U12824 (N_12824,N_11371,N_11936);
nor U12825 (N_12825,N_11859,N_11314);
and U12826 (N_12826,N_11767,N_11107);
nand U12827 (N_12827,N_11737,N_11616);
and U12828 (N_12828,N_11251,N_11741);
xnor U12829 (N_12829,N_11149,N_11361);
and U12830 (N_12830,N_11971,N_11045);
xnor U12831 (N_12831,N_11353,N_11933);
nand U12832 (N_12832,N_11087,N_11147);
nor U12833 (N_12833,N_11909,N_11418);
nand U12834 (N_12834,N_11720,N_11926);
xnor U12835 (N_12835,N_11494,N_11501);
nand U12836 (N_12836,N_11111,N_11019);
nor U12837 (N_12837,N_11053,N_11997);
nand U12838 (N_12838,N_11763,N_11407);
nand U12839 (N_12839,N_11472,N_11275);
and U12840 (N_12840,N_11619,N_11930);
nor U12841 (N_12841,N_11273,N_11709);
or U12842 (N_12842,N_11103,N_11852);
xor U12843 (N_12843,N_11062,N_11750);
and U12844 (N_12844,N_11101,N_11923);
nand U12845 (N_12845,N_11040,N_11905);
nand U12846 (N_12846,N_11074,N_11413);
nor U12847 (N_12847,N_11432,N_11820);
or U12848 (N_12848,N_11165,N_11620);
or U12849 (N_12849,N_11334,N_11282);
nor U12850 (N_12850,N_11131,N_11917);
xor U12851 (N_12851,N_11466,N_11215);
nand U12852 (N_12852,N_11674,N_11245);
and U12853 (N_12853,N_11647,N_11617);
nand U12854 (N_12854,N_11472,N_11808);
xnor U12855 (N_12855,N_11133,N_11314);
or U12856 (N_12856,N_11043,N_11592);
or U12857 (N_12857,N_11985,N_11551);
and U12858 (N_12858,N_11661,N_11757);
xor U12859 (N_12859,N_11063,N_11693);
nand U12860 (N_12860,N_11418,N_11532);
nand U12861 (N_12861,N_11935,N_11640);
nand U12862 (N_12862,N_11097,N_11414);
nor U12863 (N_12863,N_11543,N_11540);
xor U12864 (N_12864,N_11723,N_11423);
or U12865 (N_12865,N_11201,N_11930);
nor U12866 (N_12866,N_11003,N_11057);
nor U12867 (N_12867,N_11911,N_11915);
xor U12868 (N_12868,N_11817,N_11849);
or U12869 (N_12869,N_11162,N_11144);
or U12870 (N_12870,N_11331,N_11787);
and U12871 (N_12871,N_11027,N_11445);
nand U12872 (N_12872,N_11284,N_11425);
xnor U12873 (N_12873,N_11393,N_11804);
xnor U12874 (N_12874,N_11727,N_11237);
or U12875 (N_12875,N_11120,N_11366);
nand U12876 (N_12876,N_11314,N_11115);
nor U12877 (N_12877,N_11822,N_11019);
and U12878 (N_12878,N_11461,N_11336);
xor U12879 (N_12879,N_11430,N_11442);
and U12880 (N_12880,N_11707,N_11068);
and U12881 (N_12881,N_11267,N_11064);
and U12882 (N_12882,N_11435,N_11229);
nor U12883 (N_12883,N_11837,N_11966);
and U12884 (N_12884,N_11048,N_11765);
and U12885 (N_12885,N_11368,N_11009);
nor U12886 (N_12886,N_11332,N_11622);
nor U12887 (N_12887,N_11035,N_11464);
nor U12888 (N_12888,N_11361,N_11958);
nor U12889 (N_12889,N_11462,N_11811);
nand U12890 (N_12890,N_11723,N_11977);
nor U12891 (N_12891,N_11733,N_11792);
or U12892 (N_12892,N_11788,N_11643);
and U12893 (N_12893,N_11356,N_11631);
and U12894 (N_12894,N_11633,N_11351);
nand U12895 (N_12895,N_11706,N_11343);
nor U12896 (N_12896,N_11533,N_11591);
xor U12897 (N_12897,N_11432,N_11714);
nand U12898 (N_12898,N_11271,N_11334);
or U12899 (N_12899,N_11692,N_11103);
and U12900 (N_12900,N_11778,N_11581);
and U12901 (N_12901,N_11874,N_11153);
and U12902 (N_12902,N_11195,N_11936);
xnor U12903 (N_12903,N_11830,N_11304);
or U12904 (N_12904,N_11610,N_11763);
xnor U12905 (N_12905,N_11282,N_11161);
and U12906 (N_12906,N_11598,N_11542);
nor U12907 (N_12907,N_11876,N_11840);
xor U12908 (N_12908,N_11784,N_11883);
xor U12909 (N_12909,N_11900,N_11970);
xor U12910 (N_12910,N_11117,N_11870);
xor U12911 (N_12911,N_11783,N_11143);
xor U12912 (N_12912,N_11656,N_11841);
xor U12913 (N_12913,N_11561,N_11082);
and U12914 (N_12914,N_11808,N_11417);
nor U12915 (N_12915,N_11734,N_11924);
nor U12916 (N_12916,N_11318,N_11572);
or U12917 (N_12917,N_11589,N_11750);
nor U12918 (N_12918,N_11606,N_11318);
and U12919 (N_12919,N_11452,N_11322);
nor U12920 (N_12920,N_11807,N_11432);
nor U12921 (N_12921,N_11208,N_11093);
nand U12922 (N_12922,N_11112,N_11187);
or U12923 (N_12923,N_11473,N_11745);
xor U12924 (N_12924,N_11253,N_11642);
xnor U12925 (N_12925,N_11603,N_11756);
and U12926 (N_12926,N_11846,N_11746);
xnor U12927 (N_12927,N_11880,N_11276);
nand U12928 (N_12928,N_11411,N_11458);
and U12929 (N_12929,N_11581,N_11492);
nand U12930 (N_12930,N_11645,N_11026);
nand U12931 (N_12931,N_11324,N_11166);
and U12932 (N_12932,N_11087,N_11291);
and U12933 (N_12933,N_11216,N_11055);
nand U12934 (N_12934,N_11454,N_11335);
xor U12935 (N_12935,N_11634,N_11187);
xnor U12936 (N_12936,N_11613,N_11201);
nand U12937 (N_12937,N_11932,N_11515);
xor U12938 (N_12938,N_11924,N_11693);
or U12939 (N_12939,N_11857,N_11769);
nand U12940 (N_12940,N_11320,N_11087);
and U12941 (N_12941,N_11898,N_11744);
nand U12942 (N_12942,N_11813,N_11500);
nand U12943 (N_12943,N_11459,N_11969);
or U12944 (N_12944,N_11807,N_11288);
nand U12945 (N_12945,N_11253,N_11817);
nor U12946 (N_12946,N_11737,N_11928);
xor U12947 (N_12947,N_11066,N_11154);
nor U12948 (N_12948,N_11003,N_11244);
nor U12949 (N_12949,N_11973,N_11429);
and U12950 (N_12950,N_11228,N_11039);
and U12951 (N_12951,N_11547,N_11982);
or U12952 (N_12952,N_11217,N_11012);
nand U12953 (N_12953,N_11557,N_11806);
xor U12954 (N_12954,N_11135,N_11563);
and U12955 (N_12955,N_11208,N_11445);
nor U12956 (N_12956,N_11070,N_11115);
or U12957 (N_12957,N_11114,N_11059);
xnor U12958 (N_12958,N_11806,N_11359);
xor U12959 (N_12959,N_11521,N_11330);
xor U12960 (N_12960,N_11939,N_11576);
nor U12961 (N_12961,N_11700,N_11288);
and U12962 (N_12962,N_11823,N_11924);
xor U12963 (N_12963,N_11290,N_11788);
nand U12964 (N_12964,N_11833,N_11728);
and U12965 (N_12965,N_11296,N_11201);
xor U12966 (N_12966,N_11649,N_11531);
nand U12967 (N_12967,N_11615,N_11673);
or U12968 (N_12968,N_11681,N_11821);
xnor U12969 (N_12969,N_11549,N_11535);
xor U12970 (N_12970,N_11101,N_11058);
or U12971 (N_12971,N_11933,N_11028);
or U12972 (N_12972,N_11070,N_11541);
nor U12973 (N_12973,N_11496,N_11818);
or U12974 (N_12974,N_11784,N_11001);
nor U12975 (N_12975,N_11402,N_11229);
or U12976 (N_12976,N_11577,N_11518);
and U12977 (N_12977,N_11467,N_11833);
nand U12978 (N_12978,N_11236,N_11320);
and U12979 (N_12979,N_11156,N_11051);
xnor U12980 (N_12980,N_11987,N_11553);
xnor U12981 (N_12981,N_11270,N_11374);
nor U12982 (N_12982,N_11621,N_11313);
and U12983 (N_12983,N_11586,N_11746);
nor U12984 (N_12984,N_11524,N_11240);
and U12985 (N_12985,N_11658,N_11741);
nor U12986 (N_12986,N_11647,N_11566);
and U12987 (N_12987,N_11485,N_11503);
xor U12988 (N_12988,N_11849,N_11750);
nor U12989 (N_12989,N_11608,N_11997);
and U12990 (N_12990,N_11924,N_11008);
nor U12991 (N_12991,N_11169,N_11039);
and U12992 (N_12992,N_11624,N_11301);
nor U12993 (N_12993,N_11894,N_11941);
and U12994 (N_12994,N_11829,N_11951);
xor U12995 (N_12995,N_11829,N_11068);
or U12996 (N_12996,N_11640,N_11633);
nor U12997 (N_12997,N_11775,N_11457);
nor U12998 (N_12998,N_11408,N_11608);
xor U12999 (N_12999,N_11516,N_11964);
nor U13000 (N_13000,N_12999,N_12079);
nand U13001 (N_13001,N_12879,N_12149);
nand U13002 (N_13002,N_12157,N_12880);
xor U13003 (N_13003,N_12348,N_12610);
nor U13004 (N_13004,N_12775,N_12202);
nor U13005 (N_13005,N_12948,N_12389);
xnor U13006 (N_13006,N_12509,N_12305);
nor U13007 (N_13007,N_12131,N_12877);
xnor U13008 (N_13008,N_12828,N_12307);
nor U13009 (N_13009,N_12361,N_12680);
nor U13010 (N_13010,N_12069,N_12533);
xnor U13011 (N_13011,N_12770,N_12398);
xor U13012 (N_13012,N_12951,N_12074);
xnor U13013 (N_13013,N_12891,N_12747);
or U13014 (N_13014,N_12250,N_12643);
and U13015 (N_13015,N_12303,N_12511);
nor U13016 (N_13016,N_12583,N_12671);
xor U13017 (N_13017,N_12133,N_12184);
and U13018 (N_13018,N_12829,N_12379);
and U13019 (N_13019,N_12797,N_12724);
or U13020 (N_13020,N_12164,N_12431);
and U13021 (N_13021,N_12106,N_12397);
nand U13022 (N_13022,N_12504,N_12189);
nand U13023 (N_13023,N_12753,N_12630);
nand U13024 (N_13024,N_12532,N_12637);
xor U13025 (N_13025,N_12947,N_12661);
or U13026 (N_13026,N_12898,N_12900);
xor U13027 (N_13027,N_12574,N_12371);
or U13028 (N_13028,N_12415,N_12919);
nor U13029 (N_13029,N_12830,N_12567);
or U13030 (N_13030,N_12056,N_12393);
nand U13031 (N_13031,N_12049,N_12417);
or U13032 (N_13032,N_12973,N_12057);
and U13033 (N_13033,N_12743,N_12225);
xnor U13034 (N_13034,N_12104,N_12866);
and U13035 (N_13035,N_12972,N_12076);
xor U13036 (N_13036,N_12542,N_12293);
nor U13037 (N_13037,N_12997,N_12084);
xor U13038 (N_13038,N_12675,N_12683);
nor U13039 (N_13039,N_12242,N_12731);
and U13040 (N_13040,N_12055,N_12781);
xor U13041 (N_13041,N_12722,N_12600);
xnor U13042 (N_13042,N_12782,N_12950);
or U13043 (N_13043,N_12689,N_12012);
and U13044 (N_13044,N_12404,N_12459);
or U13045 (N_13045,N_12000,N_12390);
nand U13046 (N_13046,N_12014,N_12368);
or U13047 (N_13047,N_12153,N_12888);
nor U13048 (N_13048,N_12385,N_12239);
or U13049 (N_13049,N_12614,N_12757);
nand U13050 (N_13050,N_12218,N_12645);
nor U13051 (N_13051,N_12792,N_12452);
or U13052 (N_13052,N_12186,N_12045);
nor U13053 (N_13053,N_12188,N_12495);
and U13054 (N_13054,N_12146,N_12099);
or U13055 (N_13055,N_12941,N_12205);
xnor U13056 (N_13056,N_12867,N_12050);
or U13057 (N_13057,N_12844,N_12840);
xnor U13058 (N_13058,N_12328,N_12791);
and U13059 (N_13059,N_12760,N_12952);
nand U13060 (N_13060,N_12794,N_12875);
nand U13061 (N_13061,N_12489,N_12136);
xnor U13062 (N_13062,N_12020,N_12060);
nor U13063 (N_13063,N_12264,N_12969);
or U13064 (N_13064,N_12581,N_12429);
nand U13065 (N_13065,N_12147,N_12059);
and U13066 (N_13066,N_12981,N_12632);
nor U13067 (N_13067,N_12447,N_12375);
or U13068 (N_13068,N_12652,N_12721);
or U13069 (N_13069,N_12091,N_12514);
or U13070 (N_13070,N_12081,N_12508);
xor U13071 (N_13071,N_12241,N_12887);
nand U13072 (N_13072,N_12024,N_12473);
nor U13073 (N_13073,N_12736,N_12827);
nor U13074 (N_13074,N_12931,N_12923);
and U13075 (N_13075,N_12204,N_12578);
nor U13076 (N_13076,N_12565,N_12088);
and U13077 (N_13077,N_12313,N_12430);
and U13078 (N_13078,N_12247,N_12819);
nand U13079 (N_13079,N_12155,N_12917);
nor U13080 (N_13080,N_12488,N_12213);
or U13081 (N_13081,N_12198,N_12409);
nand U13082 (N_13082,N_12873,N_12309);
xor U13083 (N_13083,N_12737,N_12572);
xor U13084 (N_13084,N_12640,N_12615);
xnor U13085 (N_13085,N_12748,N_12591);
and U13086 (N_13086,N_12436,N_12858);
or U13087 (N_13087,N_12434,N_12786);
nand U13088 (N_13088,N_12622,N_12619);
and U13089 (N_13089,N_12820,N_12347);
xor U13090 (N_13090,N_12221,N_12427);
nor U13091 (N_13091,N_12501,N_12970);
or U13092 (N_13092,N_12051,N_12631);
or U13093 (N_13093,N_12989,N_12296);
or U13094 (N_13094,N_12281,N_12986);
and U13095 (N_13095,N_12550,N_12301);
xnor U13096 (N_13096,N_12647,N_12872);
or U13097 (N_13097,N_12717,N_12428);
and U13098 (N_13098,N_12925,N_12004);
and U13099 (N_13099,N_12359,N_12065);
nor U13100 (N_13100,N_12249,N_12568);
or U13101 (N_13101,N_12119,N_12400);
and U13102 (N_13102,N_12043,N_12124);
xnor U13103 (N_13103,N_12659,N_12603);
xor U13104 (N_13104,N_12723,N_12793);
nand U13105 (N_13105,N_12813,N_12103);
nand U13106 (N_13106,N_12756,N_12895);
and U13107 (N_13107,N_12804,N_12967);
xnor U13108 (N_13108,N_12444,N_12462);
xnor U13109 (N_13109,N_12524,N_12052);
nand U13110 (N_13110,N_12214,N_12573);
and U13111 (N_13111,N_12620,N_12985);
xnor U13112 (N_13112,N_12856,N_12158);
xor U13113 (N_13113,N_12196,N_12818);
nand U13114 (N_13114,N_12073,N_12148);
and U13115 (N_13115,N_12471,N_12372);
nor U13116 (N_13116,N_12850,N_12903);
and U13117 (N_13117,N_12233,N_12208);
xor U13118 (N_13118,N_12211,N_12878);
nand U13119 (N_13119,N_12267,N_12663);
nand U13120 (N_13120,N_12030,N_12773);
nand U13121 (N_13121,N_12714,N_12617);
nand U13122 (N_13122,N_12812,N_12933);
nand U13123 (N_13123,N_12472,N_12984);
or U13124 (N_13124,N_12849,N_12306);
xnor U13125 (N_13125,N_12278,N_12376);
nor U13126 (N_13126,N_12285,N_12682);
nor U13127 (N_13127,N_12512,N_12445);
nor U13128 (N_13128,N_12751,N_12983);
or U13129 (N_13129,N_12602,N_12651);
and U13130 (N_13130,N_12580,N_12121);
nor U13131 (N_13131,N_12499,N_12543);
xor U13132 (N_13132,N_12141,N_12962);
xor U13133 (N_13133,N_12920,N_12235);
or U13134 (N_13134,N_12072,N_12569);
or U13135 (N_13135,N_12621,N_12217);
xnor U13136 (N_13136,N_12808,N_12485);
and U13137 (N_13137,N_12047,N_12064);
nand U13138 (N_13138,N_12996,N_12227);
nor U13139 (N_13139,N_12749,N_12598);
or U13140 (N_13140,N_12126,N_12129);
and U13141 (N_13141,N_12926,N_12082);
nor U13142 (N_13142,N_12102,N_12790);
nor U13143 (N_13143,N_12425,N_12649);
or U13144 (N_13144,N_12505,N_12097);
and U13145 (N_13145,N_12272,N_12800);
nor U13146 (N_13146,N_12350,N_12135);
nor U13147 (N_13147,N_12279,N_12728);
xnor U13148 (N_13148,N_12071,N_12394);
nand U13149 (N_13149,N_12955,N_12381);
and U13150 (N_13150,N_12256,N_12176);
xnor U13151 (N_13151,N_12484,N_12697);
nor U13152 (N_13152,N_12727,N_12107);
nand U13153 (N_13153,N_12953,N_12396);
xnor U13154 (N_13154,N_12443,N_12465);
nor U13155 (N_13155,N_12506,N_12909);
nor U13156 (N_13156,N_12765,N_12206);
or U13157 (N_13157,N_12754,N_12324);
xor U13158 (N_13158,N_12789,N_12946);
nand U13159 (N_13159,N_12526,N_12803);
nor U13160 (N_13160,N_12776,N_12401);
nand U13161 (N_13161,N_12868,N_12657);
xnor U13162 (N_13162,N_12809,N_12384);
xor U13163 (N_13163,N_12283,N_12846);
and U13164 (N_13164,N_12628,N_12266);
nand U13165 (N_13165,N_12788,N_12694);
and U13166 (N_13166,N_12203,N_12650);
and U13167 (N_13167,N_12633,N_12382);
or U13168 (N_13168,N_12594,N_12197);
or U13169 (N_13169,N_12180,N_12624);
or U13170 (N_13170,N_12976,N_12541);
or U13171 (N_13171,N_12134,N_12678);
nor U13172 (N_13172,N_12552,N_12255);
xor U13173 (N_13173,N_12922,N_12251);
xor U13174 (N_13174,N_12492,N_12928);
nor U13175 (N_13175,N_12033,N_12639);
xor U13176 (N_13176,N_12044,N_12294);
and U13177 (N_13177,N_12597,N_12226);
nand U13178 (N_13178,N_12456,N_12168);
and U13179 (N_13179,N_12263,N_12741);
xor U13180 (N_13180,N_12716,N_12886);
xnor U13181 (N_13181,N_12535,N_12245);
nor U13182 (N_13182,N_12921,N_12817);
and U13183 (N_13183,N_12192,N_12345);
or U13184 (N_13184,N_12780,N_12116);
xnor U13185 (N_13185,N_12380,N_12584);
or U13186 (N_13186,N_12383,N_12463);
or U13187 (N_13187,N_12440,N_12496);
nor U13188 (N_13188,N_12178,N_12179);
and U13189 (N_13189,N_12587,N_12668);
xnor U13190 (N_13190,N_12490,N_12191);
xor U13191 (N_13191,N_12352,N_12286);
nor U13192 (N_13192,N_12302,N_12653);
nor U13193 (N_13193,N_12343,N_12193);
xor U13194 (N_13194,N_12699,N_12399);
and U13195 (N_13195,N_12403,N_12287);
xor U13196 (N_13196,N_12712,N_12246);
xor U13197 (N_13197,N_12988,N_12576);
or U13198 (N_13198,N_12240,N_12346);
and U13199 (N_13199,N_12522,N_12876);
or U13200 (N_13200,N_12005,N_12391);
or U13201 (N_13201,N_12304,N_12165);
nor U13202 (N_13202,N_12284,N_12686);
and U13203 (N_13203,N_12563,N_12528);
or U13204 (N_13204,N_12337,N_12118);
nand U13205 (N_13205,N_12290,N_12467);
nand U13206 (N_13206,N_12555,N_12965);
and U13207 (N_13207,N_12627,N_12558);
nor U13208 (N_13208,N_12693,N_12366);
xnor U13209 (N_13209,N_12709,N_12913);
xnor U13210 (N_13210,N_12120,N_12087);
nor U13211 (N_13211,N_12172,N_12853);
and U13212 (N_13212,N_12152,N_12270);
nand U13213 (N_13213,N_12316,N_12023);
nor U13214 (N_13214,N_12957,N_12964);
xnor U13215 (N_13215,N_12314,N_12987);
and U13216 (N_13216,N_12534,N_12130);
or U13217 (N_13217,N_12026,N_12889);
and U13218 (N_13218,N_12423,N_12021);
and U13219 (N_13219,N_12433,N_12171);
and U13220 (N_13220,N_12681,N_12312);
nand U13221 (N_13221,N_12605,N_12642);
or U13222 (N_13222,N_12871,N_12442);
or U13223 (N_13223,N_12016,N_12667);
xnor U13224 (N_13224,N_12612,N_12331);
nor U13225 (N_13225,N_12942,N_12899);
and U13226 (N_13226,N_12935,N_12351);
or U13227 (N_13227,N_12353,N_12274);
xor U13228 (N_13228,N_12322,N_12762);
nor U13229 (N_13229,N_12698,N_12520);
and U13230 (N_13230,N_12494,N_12095);
nor U13231 (N_13231,N_12029,N_12865);
nand U13232 (N_13232,N_12641,N_12507);
xor U13233 (N_13233,N_12660,N_12991);
nor U13234 (N_13234,N_12090,N_12708);
or U13235 (N_13235,N_12582,N_12549);
or U13236 (N_13236,N_12042,N_12703);
xor U13237 (N_13237,N_12785,N_12092);
xnor U13238 (N_13238,N_12609,N_12707);
xor U13239 (N_13239,N_12422,N_12339);
nor U13240 (N_13240,N_12268,N_12862);
nand U13241 (N_13241,N_12822,N_12475);
xor U13242 (N_13242,N_12607,N_12570);
nand U13243 (N_13243,N_12679,N_12861);
nand U13244 (N_13244,N_12897,N_12855);
nand U13245 (N_13245,N_12746,N_12015);
nor U13246 (N_13246,N_12117,N_12860);
nor U13247 (N_13247,N_12706,N_12028);
nor U13248 (N_13248,N_12638,N_12094);
or U13249 (N_13249,N_12655,N_12299);
or U13250 (N_13250,N_12228,N_12990);
nand U13251 (N_13251,N_12273,N_12814);
nand U13252 (N_13252,N_12008,N_12998);
and U13253 (N_13253,N_12160,N_12832);
and U13254 (N_13254,N_12025,N_12618);
or U13255 (N_13255,N_12956,N_12453);
nand U13256 (N_13256,N_12236,N_12478);
nor U13257 (N_13257,N_12695,N_12201);
nand U13258 (N_13258,N_12080,N_12938);
nor U13259 (N_13259,N_12777,N_12636);
and U13260 (N_13260,N_12666,N_12482);
xor U13261 (N_13261,N_12387,N_12177);
or U13262 (N_13262,N_12687,N_12613);
nor U13263 (N_13263,N_12677,N_12579);
xor U13264 (N_13264,N_12733,N_12159);
xnor U13265 (N_13265,N_12450,N_12027);
nor U13266 (N_13266,N_12373,N_12150);
nand U13267 (N_13267,N_12349,N_12342);
and U13268 (N_13268,N_12329,N_12138);
xnor U13269 (N_13269,N_12386,N_12901);
xnor U13270 (N_13270,N_12544,N_12701);
and U13271 (N_13271,N_12115,N_12474);
nand U13272 (N_13272,N_12561,N_12458);
nand U13273 (N_13273,N_12823,N_12061);
nor U13274 (N_13274,N_12330,N_12067);
nor U13275 (N_13275,N_12140,N_12333);
or U13276 (N_13276,N_12959,N_12519);
xnor U13277 (N_13277,N_12019,N_12487);
nor U13278 (N_13278,N_12715,N_12608);
nor U13279 (N_13279,N_12904,N_12257);
nor U13280 (N_13280,N_12571,N_12169);
and U13281 (N_13281,N_12344,N_12013);
nor U13282 (N_13282,N_12711,N_12864);
and U13283 (N_13283,N_12805,N_12289);
and U13284 (N_13284,N_12945,N_12835);
nor U13285 (N_13285,N_12611,N_12843);
xnor U13286 (N_13286,N_12934,N_12658);
nand U13287 (N_13287,N_12363,N_12093);
and U13288 (N_13288,N_12109,N_12908);
and U13289 (N_13289,N_12195,N_12470);
or U13290 (N_13290,N_12362,N_12364);
and U13291 (N_13291,N_12032,N_12455);
xor U13292 (N_13292,N_12662,N_12132);
or U13293 (N_13293,N_12958,N_12317);
and U13294 (N_13294,N_12426,N_12995);
and U13295 (N_13295,N_12838,N_12626);
or U13296 (N_13296,N_12464,N_12419);
nand U13297 (N_13297,N_12261,N_12486);
or U13298 (N_13298,N_12915,N_12960);
nor U13299 (N_13299,N_12085,N_12801);
xor U13300 (N_13300,N_12537,N_12968);
xor U13301 (N_13301,N_12821,N_12625);
or U13302 (N_13302,N_12411,N_12414);
and U13303 (N_13303,N_12599,N_12039);
nand U13304 (N_13304,N_12825,N_12220);
nor U13305 (N_13305,N_12479,N_12408);
or U13306 (N_13306,N_12231,N_12772);
xor U13307 (N_13307,N_12916,N_12105);
or U13308 (N_13308,N_12248,N_12734);
and U13309 (N_13309,N_12367,N_12310);
xor U13310 (N_13310,N_12833,N_12377);
nand U13311 (N_13311,N_12810,N_12575);
nor U13312 (N_13312,N_12112,N_12525);
and U13313 (N_13313,N_12936,N_12167);
nor U13314 (N_13314,N_12066,N_12139);
and U13315 (N_13315,N_12604,N_12518);
nand U13316 (N_13316,N_12837,N_12100);
nor U13317 (N_13317,N_12798,N_12730);
nor U13318 (N_13318,N_12852,N_12654);
or U13319 (N_13319,N_12435,N_12732);
and U13320 (N_13320,N_12282,N_12779);
and U13321 (N_13321,N_12851,N_12321);
or U13322 (N_13322,N_12318,N_12966);
or U13323 (N_13323,N_12114,N_12262);
and U13324 (N_13324,N_12906,N_12767);
nand U13325 (N_13325,N_12229,N_12181);
or U13326 (N_13326,N_12356,N_12592);
or U13327 (N_13327,N_12212,N_12702);
and U13328 (N_13328,N_12726,N_12690);
nor U13329 (N_13329,N_12108,N_12416);
xnor U13330 (N_13330,N_12128,N_12778);
xor U13331 (N_13331,N_12216,N_12038);
nor U13332 (N_13332,N_12295,N_12327);
xnor U13333 (N_13333,N_12360,N_12815);
nor U13334 (N_13334,N_12939,N_12927);
and U13335 (N_13335,N_12766,N_12560);
xnor U13336 (N_13336,N_12980,N_12842);
xor U13337 (N_13337,N_12011,N_12554);
nor U13338 (N_13338,N_12845,N_12841);
nor U13339 (N_13339,N_12127,N_12392);
xnor U13340 (N_13340,N_12672,N_12774);
nor U13341 (N_13341,N_12545,N_12491);
xor U13342 (N_13342,N_12446,N_12665);
nand U13343 (N_13343,N_12924,N_12557);
nand U13344 (N_13344,N_12940,N_12918);
nand U13345 (N_13345,N_12101,N_12145);
nor U13346 (N_13346,N_12993,N_12089);
or U13347 (N_13347,N_12300,N_12311);
nor U13348 (N_13348,N_12824,N_12308);
nand U13349 (N_13349,N_12854,N_12685);
nand U13350 (N_13350,N_12298,N_12523);
and U13351 (N_13351,N_12355,N_12113);
xor U13352 (N_13352,N_12292,N_12476);
and U13353 (N_13353,N_12253,N_12963);
nand U13354 (N_13354,N_12483,N_12863);
xor U13355 (N_13355,N_12735,N_12469);
nand U13356 (N_13356,N_12438,N_12516);
nor U13357 (N_13357,N_12110,N_12811);
nor U13358 (N_13358,N_12215,N_12006);
xnor U13359 (N_13359,N_12468,N_12688);
or U13360 (N_13360,N_12077,N_12288);
xor U13361 (N_13361,N_12338,N_12577);
nand U13362 (N_13362,N_12590,N_12907);
xnor U13363 (N_13363,N_12629,N_12497);
nand U13364 (N_13364,N_12676,N_12031);
or U13365 (N_13365,N_12839,N_12513);
and U13366 (N_13366,N_12378,N_12365);
xnor U13367 (N_13367,N_12161,N_12538);
or U13368 (N_13368,N_12692,N_12949);
and U13369 (N_13369,N_12173,N_12725);
nand U13370 (N_13370,N_12200,N_12596);
nor U13371 (N_13371,N_12498,N_12977);
nand U13372 (N_13372,N_12859,N_12277);
or U13373 (N_13373,N_12884,N_12418);
nand U13374 (N_13374,N_12546,N_12493);
or U13375 (N_13375,N_12644,N_12326);
nand U13376 (N_13376,N_12807,N_12710);
or U13377 (N_13377,N_12902,N_12125);
nor U13378 (N_13378,N_12451,N_12937);
or U13379 (N_13379,N_12847,N_12787);
xor U13380 (N_13380,N_12562,N_12258);
or U13381 (N_13381,N_12063,N_12374);
and U13382 (N_13382,N_12616,N_12199);
nor U13383 (N_13383,N_12530,N_12882);
nand U13384 (N_13384,N_12740,N_12784);
and U13385 (N_13385,N_12003,N_12122);
nand U13386 (N_13386,N_12783,N_12040);
and U13387 (N_13387,N_12664,N_12869);
and U13388 (N_13388,N_12238,N_12589);
nand U13389 (N_13389,N_12078,N_12971);
and U13390 (N_13390,N_12836,N_12515);
xor U13391 (N_13391,N_12883,N_12700);
xnor U13392 (N_13392,N_12232,N_12595);
and U13393 (N_13393,N_12369,N_12761);
xnor U13394 (N_13394,N_12744,N_12466);
and U13395 (N_13395,N_12586,N_12407);
nand U13396 (N_13396,N_12547,N_12075);
and U13397 (N_13397,N_12502,N_12182);
nand U13398 (N_13398,N_12243,N_12357);
xnor U13399 (N_13399,N_12527,N_12460);
or U13400 (N_13400,N_12529,N_12448);
and U13401 (N_13401,N_12244,N_12319);
xor U13402 (N_13402,N_12271,N_12022);
and U13403 (N_13403,N_12291,N_12826);
nor U13404 (N_13404,N_12768,N_12230);
xnor U13405 (N_13405,N_12691,N_12911);
nand U13406 (N_13406,N_12704,N_12635);
or U13407 (N_13407,N_12234,N_12265);
xor U13408 (N_13408,N_12806,N_12062);
and U13409 (N_13409,N_12439,N_12010);
xor U13410 (N_13410,N_12054,N_12332);
and U13411 (N_13411,N_12297,N_12816);
nor U13412 (N_13412,N_12961,N_12564);
or U13413 (N_13413,N_12752,N_12795);
and U13414 (N_13414,N_12222,N_12932);
xor U13415 (N_13415,N_12252,N_12457);
nor U13416 (N_13416,N_12548,N_12481);
nand U13417 (N_13417,N_12914,N_12536);
or U13418 (N_13418,N_12503,N_12750);
or U13419 (N_13419,N_12738,N_12881);
nand U13420 (N_13420,N_12154,N_12718);
xnor U13421 (N_13421,N_12531,N_12943);
nor U13422 (N_13422,N_12796,N_12402);
or U13423 (N_13423,N_12009,N_12035);
xor U13424 (N_13424,N_12269,N_12175);
or U13425 (N_13425,N_12406,N_12183);
and U13426 (N_13426,N_12551,N_12954);
xnor U13427 (N_13427,N_12480,N_12593);
or U13428 (N_13428,N_12994,N_12340);
nor U13429 (N_13429,N_12098,N_12223);
or U13430 (N_13430,N_12151,N_12163);
and U13431 (N_13431,N_12111,N_12068);
or U13432 (N_13432,N_12237,N_12334);
or U13433 (N_13433,N_12510,N_12388);
nand U13434 (N_13434,N_12219,N_12831);
xnor U13435 (N_13435,N_12719,N_12410);
or U13436 (N_13436,N_12207,N_12713);
nor U13437 (N_13437,N_12001,N_12017);
and U13438 (N_13438,N_12421,N_12684);
and U13439 (N_13439,N_12894,N_12764);
and U13440 (N_13440,N_12979,N_12566);
nor U13441 (N_13441,N_12500,N_12556);
and U13442 (N_13442,N_12771,N_12975);
xnor U13443 (N_13443,N_12323,N_12018);
xor U13444 (N_13444,N_12280,N_12669);
nand U13445 (N_13445,N_12978,N_12058);
nand U13446 (N_13446,N_12174,N_12162);
nand U13447 (N_13447,N_12194,N_12315);
nor U13448 (N_13448,N_12086,N_12540);
xor U13449 (N_13449,N_12893,N_12930);
and U13450 (N_13450,N_12769,N_12673);
and U13451 (N_13451,N_12896,N_12123);
and U13452 (N_13452,N_12929,N_12053);
or U13453 (N_13453,N_12041,N_12992);
nor U13454 (N_13454,N_12170,N_12424);
xor U13455 (N_13455,N_12190,N_12848);
nor U13456 (N_13456,N_12646,N_12910);
and U13457 (N_13457,N_12432,N_12634);
nor U13458 (N_13458,N_12354,N_12370);
and U13459 (N_13459,N_12517,N_12857);
nand U13460 (N_13460,N_12729,N_12674);
nand U13461 (N_13461,N_12623,N_12143);
xnor U13462 (N_13462,N_12083,N_12890);
and U13463 (N_13463,N_12648,N_12696);
xor U13464 (N_13464,N_12007,N_12905);
nand U13465 (N_13465,N_12585,N_12912);
or U13466 (N_13466,N_12395,N_12254);
xnor U13467 (N_13467,N_12588,N_12210);
or U13468 (N_13468,N_12036,N_12553);
and U13469 (N_13469,N_12763,N_12670);
nand U13470 (N_13470,N_12046,N_12437);
or U13471 (N_13471,N_12834,N_12870);
or U13472 (N_13472,N_12720,N_12166);
nand U13473 (N_13473,N_12974,N_12209);
nor U13474 (N_13474,N_12144,N_12799);
nor U13475 (N_13475,N_12521,N_12096);
and U13476 (N_13476,N_12325,N_12874);
xnor U13477 (N_13477,N_12802,N_12705);
nand U13478 (N_13478,N_12758,N_12002);
and U13479 (N_13479,N_12260,N_12156);
and U13480 (N_13480,N_12259,N_12405);
xnor U13481 (N_13481,N_12137,N_12413);
nor U13482 (N_13482,N_12944,N_12441);
and U13483 (N_13483,N_12412,N_12070);
nand U13484 (N_13484,N_12656,N_12982);
xor U13485 (N_13485,N_12454,N_12187);
nor U13486 (N_13486,N_12224,N_12606);
or U13487 (N_13487,N_12739,N_12601);
nor U13488 (N_13488,N_12759,N_12276);
or U13489 (N_13489,N_12745,N_12420);
xor U13490 (N_13490,N_12449,N_12892);
and U13491 (N_13491,N_12755,N_12559);
and U13492 (N_13492,N_12358,N_12034);
nand U13493 (N_13493,N_12885,N_12048);
and U13494 (N_13494,N_12142,N_12275);
nand U13495 (N_13495,N_12185,N_12320);
nor U13496 (N_13496,N_12335,N_12336);
or U13497 (N_13497,N_12341,N_12461);
nand U13498 (N_13498,N_12539,N_12037);
or U13499 (N_13499,N_12477,N_12742);
nand U13500 (N_13500,N_12644,N_12155);
or U13501 (N_13501,N_12467,N_12835);
nand U13502 (N_13502,N_12151,N_12458);
or U13503 (N_13503,N_12168,N_12992);
and U13504 (N_13504,N_12571,N_12044);
and U13505 (N_13505,N_12974,N_12738);
and U13506 (N_13506,N_12507,N_12074);
and U13507 (N_13507,N_12025,N_12111);
nor U13508 (N_13508,N_12932,N_12600);
or U13509 (N_13509,N_12300,N_12987);
nand U13510 (N_13510,N_12177,N_12812);
nand U13511 (N_13511,N_12403,N_12412);
and U13512 (N_13512,N_12598,N_12377);
nand U13513 (N_13513,N_12116,N_12456);
and U13514 (N_13514,N_12351,N_12079);
xnor U13515 (N_13515,N_12786,N_12625);
and U13516 (N_13516,N_12677,N_12415);
or U13517 (N_13517,N_12442,N_12855);
and U13518 (N_13518,N_12697,N_12563);
xnor U13519 (N_13519,N_12481,N_12599);
nand U13520 (N_13520,N_12873,N_12030);
xnor U13521 (N_13521,N_12710,N_12385);
nor U13522 (N_13522,N_12978,N_12680);
nor U13523 (N_13523,N_12347,N_12759);
and U13524 (N_13524,N_12709,N_12769);
nand U13525 (N_13525,N_12046,N_12361);
or U13526 (N_13526,N_12821,N_12998);
or U13527 (N_13527,N_12947,N_12922);
xnor U13528 (N_13528,N_12989,N_12271);
xnor U13529 (N_13529,N_12906,N_12529);
or U13530 (N_13530,N_12680,N_12678);
nor U13531 (N_13531,N_12990,N_12934);
nand U13532 (N_13532,N_12882,N_12685);
or U13533 (N_13533,N_12342,N_12294);
or U13534 (N_13534,N_12929,N_12868);
or U13535 (N_13535,N_12713,N_12258);
nor U13536 (N_13536,N_12074,N_12891);
nor U13537 (N_13537,N_12208,N_12859);
nand U13538 (N_13538,N_12326,N_12184);
nor U13539 (N_13539,N_12046,N_12857);
or U13540 (N_13540,N_12808,N_12857);
nor U13541 (N_13541,N_12561,N_12055);
xnor U13542 (N_13542,N_12615,N_12076);
or U13543 (N_13543,N_12619,N_12746);
and U13544 (N_13544,N_12074,N_12381);
nand U13545 (N_13545,N_12689,N_12424);
or U13546 (N_13546,N_12925,N_12047);
xnor U13547 (N_13547,N_12420,N_12293);
nand U13548 (N_13548,N_12796,N_12378);
xor U13549 (N_13549,N_12362,N_12915);
nor U13550 (N_13550,N_12874,N_12988);
and U13551 (N_13551,N_12843,N_12652);
xor U13552 (N_13552,N_12119,N_12048);
nor U13553 (N_13553,N_12773,N_12668);
nand U13554 (N_13554,N_12684,N_12367);
nor U13555 (N_13555,N_12808,N_12886);
xor U13556 (N_13556,N_12841,N_12511);
xnor U13557 (N_13557,N_12459,N_12278);
and U13558 (N_13558,N_12391,N_12022);
and U13559 (N_13559,N_12046,N_12234);
nor U13560 (N_13560,N_12816,N_12911);
nor U13561 (N_13561,N_12038,N_12016);
nand U13562 (N_13562,N_12528,N_12783);
or U13563 (N_13563,N_12960,N_12217);
nor U13564 (N_13564,N_12305,N_12645);
or U13565 (N_13565,N_12347,N_12017);
and U13566 (N_13566,N_12794,N_12430);
xor U13567 (N_13567,N_12164,N_12651);
nand U13568 (N_13568,N_12588,N_12497);
nor U13569 (N_13569,N_12297,N_12459);
nor U13570 (N_13570,N_12739,N_12705);
nand U13571 (N_13571,N_12148,N_12588);
nand U13572 (N_13572,N_12899,N_12276);
xnor U13573 (N_13573,N_12730,N_12672);
or U13574 (N_13574,N_12211,N_12476);
xnor U13575 (N_13575,N_12382,N_12435);
nand U13576 (N_13576,N_12311,N_12284);
nand U13577 (N_13577,N_12261,N_12637);
and U13578 (N_13578,N_12374,N_12575);
and U13579 (N_13579,N_12019,N_12550);
and U13580 (N_13580,N_12871,N_12466);
or U13581 (N_13581,N_12346,N_12530);
nor U13582 (N_13582,N_12979,N_12160);
or U13583 (N_13583,N_12631,N_12728);
xor U13584 (N_13584,N_12722,N_12905);
nor U13585 (N_13585,N_12728,N_12375);
or U13586 (N_13586,N_12100,N_12275);
nand U13587 (N_13587,N_12001,N_12340);
and U13588 (N_13588,N_12559,N_12737);
or U13589 (N_13589,N_12603,N_12965);
or U13590 (N_13590,N_12921,N_12811);
xor U13591 (N_13591,N_12738,N_12473);
or U13592 (N_13592,N_12005,N_12986);
nor U13593 (N_13593,N_12671,N_12668);
or U13594 (N_13594,N_12724,N_12646);
and U13595 (N_13595,N_12483,N_12391);
or U13596 (N_13596,N_12118,N_12201);
nand U13597 (N_13597,N_12982,N_12319);
nor U13598 (N_13598,N_12567,N_12420);
nor U13599 (N_13599,N_12604,N_12254);
and U13600 (N_13600,N_12138,N_12671);
or U13601 (N_13601,N_12458,N_12650);
xnor U13602 (N_13602,N_12979,N_12178);
nand U13603 (N_13603,N_12709,N_12737);
xor U13604 (N_13604,N_12439,N_12771);
xnor U13605 (N_13605,N_12015,N_12796);
xor U13606 (N_13606,N_12351,N_12938);
and U13607 (N_13607,N_12547,N_12182);
or U13608 (N_13608,N_12888,N_12581);
nand U13609 (N_13609,N_12402,N_12444);
or U13610 (N_13610,N_12173,N_12660);
xnor U13611 (N_13611,N_12053,N_12637);
nand U13612 (N_13612,N_12104,N_12647);
or U13613 (N_13613,N_12534,N_12383);
and U13614 (N_13614,N_12643,N_12681);
nand U13615 (N_13615,N_12985,N_12470);
nor U13616 (N_13616,N_12526,N_12456);
xor U13617 (N_13617,N_12950,N_12952);
nand U13618 (N_13618,N_12946,N_12640);
xnor U13619 (N_13619,N_12125,N_12890);
or U13620 (N_13620,N_12858,N_12027);
nor U13621 (N_13621,N_12801,N_12753);
xor U13622 (N_13622,N_12239,N_12944);
and U13623 (N_13623,N_12246,N_12301);
nor U13624 (N_13624,N_12226,N_12444);
or U13625 (N_13625,N_12145,N_12038);
xor U13626 (N_13626,N_12583,N_12385);
nor U13627 (N_13627,N_12978,N_12309);
nand U13628 (N_13628,N_12233,N_12521);
and U13629 (N_13629,N_12590,N_12976);
and U13630 (N_13630,N_12695,N_12678);
or U13631 (N_13631,N_12718,N_12981);
or U13632 (N_13632,N_12175,N_12423);
nand U13633 (N_13633,N_12300,N_12273);
and U13634 (N_13634,N_12711,N_12080);
and U13635 (N_13635,N_12474,N_12809);
nor U13636 (N_13636,N_12931,N_12155);
xor U13637 (N_13637,N_12888,N_12565);
and U13638 (N_13638,N_12387,N_12115);
xor U13639 (N_13639,N_12814,N_12709);
nor U13640 (N_13640,N_12230,N_12103);
nand U13641 (N_13641,N_12190,N_12889);
and U13642 (N_13642,N_12617,N_12306);
nand U13643 (N_13643,N_12845,N_12325);
xnor U13644 (N_13644,N_12101,N_12525);
nand U13645 (N_13645,N_12680,N_12120);
xnor U13646 (N_13646,N_12018,N_12191);
and U13647 (N_13647,N_12306,N_12068);
and U13648 (N_13648,N_12010,N_12729);
or U13649 (N_13649,N_12957,N_12986);
nand U13650 (N_13650,N_12450,N_12011);
and U13651 (N_13651,N_12836,N_12368);
xor U13652 (N_13652,N_12276,N_12369);
xor U13653 (N_13653,N_12132,N_12609);
xor U13654 (N_13654,N_12862,N_12077);
nor U13655 (N_13655,N_12836,N_12385);
or U13656 (N_13656,N_12611,N_12388);
nand U13657 (N_13657,N_12292,N_12253);
nor U13658 (N_13658,N_12995,N_12876);
nand U13659 (N_13659,N_12487,N_12977);
or U13660 (N_13660,N_12602,N_12940);
nor U13661 (N_13661,N_12190,N_12105);
and U13662 (N_13662,N_12598,N_12496);
nand U13663 (N_13663,N_12652,N_12818);
and U13664 (N_13664,N_12628,N_12934);
or U13665 (N_13665,N_12649,N_12801);
xnor U13666 (N_13666,N_12033,N_12490);
nor U13667 (N_13667,N_12351,N_12173);
and U13668 (N_13668,N_12309,N_12398);
and U13669 (N_13669,N_12348,N_12185);
or U13670 (N_13670,N_12986,N_12546);
xnor U13671 (N_13671,N_12489,N_12725);
nand U13672 (N_13672,N_12029,N_12018);
and U13673 (N_13673,N_12480,N_12230);
or U13674 (N_13674,N_12984,N_12536);
xnor U13675 (N_13675,N_12842,N_12259);
xnor U13676 (N_13676,N_12495,N_12511);
or U13677 (N_13677,N_12867,N_12096);
nand U13678 (N_13678,N_12311,N_12948);
and U13679 (N_13679,N_12443,N_12095);
nor U13680 (N_13680,N_12960,N_12712);
nand U13681 (N_13681,N_12930,N_12255);
or U13682 (N_13682,N_12929,N_12700);
and U13683 (N_13683,N_12503,N_12133);
nor U13684 (N_13684,N_12724,N_12769);
nor U13685 (N_13685,N_12468,N_12103);
and U13686 (N_13686,N_12601,N_12607);
or U13687 (N_13687,N_12949,N_12200);
nand U13688 (N_13688,N_12590,N_12179);
nand U13689 (N_13689,N_12013,N_12522);
xor U13690 (N_13690,N_12576,N_12956);
xor U13691 (N_13691,N_12711,N_12402);
or U13692 (N_13692,N_12685,N_12835);
xnor U13693 (N_13693,N_12977,N_12466);
xnor U13694 (N_13694,N_12171,N_12001);
xor U13695 (N_13695,N_12175,N_12115);
and U13696 (N_13696,N_12728,N_12298);
or U13697 (N_13697,N_12467,N_12999);
nor U13698 (N_13698,N_12847,N_12271);
or U13699 (N_13699,N_12999,N_12414);
and U13700 (N_13700,N_12722,N_12376);
and U13701 (N_13701,N_12931,N_12335);
nand U13702 (N_13702,N_12136,N_12353);
nand U13703 (N_13703,N_12659,N_12733);
or U13704 (N_13704,N_12967,N_12115);
nand U13705 (N_13705,N_12421,N_12276);
and U13706 (N_13706,N_12717,N_12443);
or U13707 (N_13707,N_12380,N_12596);
or U13708 (N_13708,N_12549,N_12909);
nand U13709 (N_13709,N_12219,N_12859);
nand U13710 (N_13710,N_12971,N_12570);
or U13711 (N_13711,N_12163,N_12241);
nor U13712 (N_13712,N_12885,N_12024);
xnor U13713 (N_13713,N_12530,N_12433);
xor U13714 (N_13714,N_12457,N_12098);
nand U13715 (N_13715,N_12982,N_12818);
xnor U13716 (N_13716,N_12118,N_12328);
nand U13717 (N_13717,N_12754,N_12436);
and U13718 (N_13718,N_12442,N_12494);
nand U13719 (N_13719,N_12427,N_12508);
nand U13720 (N_13720,N_12242,N_12862);
or U13721 (N_13721,N_12972,N_12306);
and U13722 (N_13722,N_12331,N_12428);
and U13723 (N_13723,N_12432,N_12341);
or U13724 (N_13724,N_12456,N_12140);
xor U13725 (N_13725,N_12739,N_12697);
xor U13726 (N_13726,N_12939,N_12869);
nand U13727 (N_13727,N_12413,N_12940);
or U13728 (N_13728,N_12819,N_12589);
nand U13729 (N_13729,N_12677,N_12187);
and U13730 (N_13730,N_12774,N_12155);
and U13731 (N_13731,N_12397,N_12874);
or U13732 (N_13732,N_12594,N_12270);
nand U13733 (N_13733,N_12744,N_12900);
nand U13734 (N_13734,N_12781,N_12024);
or U13735 (N_13735,N_12796,N_12762);
nand U13736 (N_13736,N_12378,N_12942);
nand U13737 (N_13737,N_12116,N_12318);
or U13738 (N_13738,N_12222,N_12448);
nand U13739 (N_13739,N_12901,N_12205);
xnor U13740 (N_13740,N_12512,N_12199);
nor U13741 (N_13741,N_12126,N_12444);
or U13742 (N_13742,N_12510,N_12679);
and U13743 (N_13743,N_12313,N_12519);
and U13744 (N_13744,N_12247,N_12998);
xnor U13745 (N_13745,N_12161,N_12171);
xor U13746 (N_13746,N_12336,N_12450);
and U13747 (N_13747,N_12744,N_12115);
and U13748 (N_13748,N_12121,N_12866);
nand U13749 (N_13749,N_12946,N_12124);
nand U13750 (N_13750,N_12802,N_12743);
and U13751 (N_13751,N_12939,N_12872);
xnor U13752 (N_13752,N_12921,N_12942);
or U13753 (N_13753,N_12018,N_12875);
nor U13754 (N_13754,N_12977,N_12863);
and U13755 (N_13755,N_12441,N_12339);
xor U13756 (N_13756,N_12165,N_12907);
or U13757 (N_13757,N_12367,N_12143);
nand U13758 (N_13758,N_12780,N_12698);
nor U13759 (N_13759,N_12055,N_12308);
and U13760 (N_13760,N_12235,N_12777);
xnor U13761 (N_13761,N_12491,N_12412);
or U13762 (N_13762,N_12457,N_12007);
xnor U13763 (N_13763,N_12387,N_12576);
nand U13764 (N_13764,N_12473,N_12285);
xnor U13765 (N_13765,N_12341,N_12120);
xor U13766 (N_13766,N_12156,N_12281);
nor U13767 (N_13767,N_12585,N_12645);
xor U13768 (N_13768,N_12908,N_12747);
and U13769 (N_13769,N_12331,N_12161);
or U13770 (N_13770,N_12620,N_12137);
nand U13771 (N_13771,N_12995,N_12062);
xor U13772 (N_13772,N_12915,N_12280);
and U13773 (N_13773,N_12766,N_12285);
nand U13774 (N_13774,N_12864,N_12663);
nand U13775 (N_13775,N_12041,N_12201);
and U13776 (N_13776,N_12892,N_12192);
and U13777 (N_13777,N_12745,N_12077);
xor U13778 (N_13778,N_12158,N_12417);
or U13779 (N_13779,N_12247,N_12771);
xor U13780 (N_13780,N_12755,N_12555);
nand U13781 (N_13781,N_12604,N_12711);
nand U13782 (N_13782,N_12601,N_12989);
and U13783 (N_13783,N_12855,N_12291);
and U13784 (N_13784,N_12838,N_12453);
nand U13785 (N_13785,N_12959,N_12003);
or U13786 (N_13786,N_12666,N_12871);
nor U13787 (N_13787,N_12948,N_12489);
or U13788 (N_13788,N_12260,N_12162);
nand U13789 (N_13789,N_12401,N_12988);
nor U13790 (N_13790,N_12675,N_12005);
nand U13791 (N_13791,N_12603,N_12552);
nor U13792 (N_13792,N_12525,N_12702);
or U13793 (N_13793,N_12684,N_12858);
xor U13794 (N_13794,N_12798,N_12477);
nand U13795 (N_13795,N_12203,N_12154);
or U13796 (N_13796,N_12650,N_12201);
and U13797 (N_13797,N_12186,N_12184);
or U13798 (N_13798,N_12860,N_12078);
or U13799 (N_13799,N_12848,N_12113);
nand U13800 (N_13800,N_12712,N_12720);
or U13801 (N_13801,N_12163,N_12862);
xor U13802 (N_13802,N_12257,N_12614);
nand U13803 (N_13803,N_12383,N_12051);
or U13804 (N_13804,N_12985,N_12846);
or U13805 (N_13805,N_12763,N_12329);
nor U13806 (N_13806,N_12579,N_12803);
nand U13807 (N_13807,N_12716,N_12504);
xnor U13808 (N_13808,N_12433,N_12546);
nand U13809 (N_13809,N_12947,N_12574);
nor U13810 (N_13810,N_12290,N_12175);
and U13811 (N_13811,N_12055,N_12687);
nand U13812 (N_13812,N_12084,N_12110);
nor U13813 (N_13813,N_12098,N_12762);
and U13814 (N_13814,N_12884,N_12645);
and U13815 (N_13815,N_12373,N_12279);
nand U13816 (N_13816,N_12655,N_12430);
xnor U13817 (N_13817,N_12478,N_12722);
nor U13818 (N_13818,N_12565,N_12286);
xor U13819 (N_13819,N_12720,N_12068);
or U13820 (N_13820,N_12327,N_12608);
xor U13821 (N_13821,N_12275,N_12492);
and U13822 (N_13822,N_12350,N_12844);
nand U13823 (N_13823,N_12868,N_12429);
and U13824 (N_13824,N_12427,N_12809);
xnor U13825 (N_13825,N_12126,N_12933);
xor U13826 (N_13826,N_12389,N_12588);
xor U13827 (N_13827,N_12917,N_12314);
or U13828 (N_13828,N_12129,N_12637);
and U13829 (N_13829,N_12822,N_12839);
xnor U13830 (N_13830,N_12002,N_12466);
nand U13831 (N_13831,N_12437,N_12068);
xor U13832 (N_13832,N_12859,N_12558);
xnor U13833 (N_13833,N_12182,N_12929);
nand U13834 (N_13834,N_12922,N_12568);
or U13835 (N_13835,N_12238,N_12895);
nor U13836 (N_13836,N_12413,N_12833);
or U13837 (N_13837,N_12723,N_12556);
nor U13838 (N_13838,N_12448,N_12994);
nor U13839 (N_13839,N_12973,N_12888);
xor U13840 (N_13840,N_12446,N_12174);
and U13841 (N_13841,N_12571,N_12770);
nand U13842 (N_13842,N_12510,N_12061);
and U13843 (N_13843,N_12824,N_12020);
nor U13844 (N_13844,N_12046,N_12271);
nand U13845 (N_13845,N_12029,N_12779);
and U13846 (N_13846,N_12437,N_12022);
nor U13847 (N_13847,N_12096,N_12061);
or U13848 (N_13848,N_12116,N_12753);
xnor U13849 (N_13849,N_12240,N_12677);
nor U13850 (N_13850,N_12582,N_12253);
nor U13851 (N_13851,N_12881,N_12403);
nor U13852 (N_13852,N_12411,N_12715);
nor U13853 (N_13853,N_12746,N_12665);
or U13854 (N_13854,N_12281,N_12480);
or U13855 (N_13855,N_12074,N_12374);
or U13856 (N_13856,N_12277,N_12075);
nand U13857 (N_13857,N_12278,N_12979);
xnor U13858 (N_13858,N_12622,N_12282);
nand U13859 (N_13859,N_12198,N_12499);
xor U13860 (N_13860,N_12700,N_12202);
and U13861 (N_13861,N_12954,N_12529);
or U13862 (N_13862,N_12891,N_12180);
nand U13863 (N_13863,N_12412,N_12687);
and U13864 (N_13864,N_12353,N_12797);
nand U13865 (N_13865,N_12722,N_12883);
and U13866 (N_13866,N_12918,N_12350);
xnor U13867 (N_13867,N_12343,N_12529);
nor U13868 (N_13868,N_12874,N_12843);
xnor U13869 (N_13869,N_12224,N_12165);
and U13870 (N_13870,N_12149,N_12664);
or U13871 (N_13871,N_12672,N_12331);
and U13872 (N_13872,N_12716,N_12124);
nor U13873 (N_13873,N_12057,N_12993);
nor U13874 (N_13874,N_12741,N_12837);
and U13875 (N_13875,N_12161,N_12157);
xnor U13876 (N_13876,N_12852,N_12184);
or U13877 (N_13877,N_12748,N_12844);
nor U13878 (N_13878,N_12257,N_12413);
or U13879 (N_13879,N_12140,N_12466);
nand U13880 (N_13880,N_12084,N_12180);
nand U13881 (N_13881,N_12449,N_12181);
and U13882 (N_13882,N_12113,N_12024);
xor U13883 (N_13883,N_12497,N_12150);
or U13884 (N_13884,N_12088,N_12855);
xor U13885 (N_13885,N_12155,N_12674);
and U13886 (N_13886,N_12674,N_12613);
nand U13887 (N_13887,N_12830,N_12595);
xnor U13888 (N_13888,N_12092,N_12705);
nand U13889 (N_13889,N_12489,N_12727);
nand U13890 (N_13890,N_12603,N_12664);
nor U13891 (N_13891,N_12944,N_12618);
nor U13892 (N_13892,N_12585,N_12056);
and U13893 (N_13893,N_12315,N_12941);
nand U13894 (N_13894,N_12005,N_12543);
and U13895 (N_13895,N_12244,N_12817);
nand U13896 (N_13896,N_12163,N_12963);
xnor U13897 (N_13897,N_12782,N_12748);
nor U13898 (N_13898,N_12109,N_12661);
and U13899 (N_13899,N_12349,N_12594);
or U13900 (N_13900,N_12905,N_12613);
and U13901 (N_13901,N_12898,N_12837);
xnor U13902 (N_13902,N_12787,N_12033);
and U13903 (N_13903,N_12303,N_12126);
and U13904 (N_13904,N_12618,N_12396);
and U13905 (N_13905,N_12452,N_12494);
xor U13906 (N_13906,N_12845,N_12225);
nor U13907 (N_13907,N_12940,N_12255);
xnor U13908 (N_13908,N_12863,N_12405);
and U13909 (N_13909,N_12774,N_12870);
or U13910 (N_13910,N_12021,N_12016);
xnor U13911 (N_13911,N_12322,N_12347);
and U13912 (N_13912,N_12599,N_12687);
nor U13913 (N_13913,N_12341,N_12865);
and U13914 (N_13914,N_12552,N_12373);
nor U13915 (N_13915,N_12144,N_12982);
nand U13916 (N_13916,N_12418,N_12167);
and U13917 (N_13917,N_12926,N_12178);
and U13918 (N_13918,N_12562,N_12464);
nor U13919 (N_13919,N_12188,N_12613);
or U13920 (N_13920,N_12077,N_12572);
or U13921 (N_13921,N_12647,N_12911);
nand U13922 (N_13922,N_12819,N_12935);
or U13923 (N_13923,N_12842,N_12683);
and U13924 (N_13924,N_12746,N_12921);
xnor U13925 (N_13925,N_12004,N_12708);
nand U13926 (N_13926,N_12967,N_12883);
nor U13927 (N_13927,N_12601,N_12535);
xor U13928 (N_13928,N_12835,N_12142);
and U13929 (N_13929,N_12868,N_12123);
or U13930 (N_13930,N_12019,N_12355);
nor U13931 (N_13931,N_12653,N_12149);
nand U13932 (N_13932,N_12911,N_12165);
and U13933 (N_13933,N_12320,N_12073);
xor U13934 (N_13934,N_12313,N_12889);
nand U13935 (N_13935,N_12983,N_12824);
and U13936 (N_13936,N_12862,N_12960);
nand U13937 (N_13937,N_12144,N_12085);
nand U13938 (N_13938,N_12784,N_12350);
xor U13939 (N_13939,N_12962,N_12503);
and U13940 (N_13940,N_12154,N_12593);
and U13941 (N_13941,N_12003,N_12503);
or U13942 (N_13942,N_12380,N_12933);
nor U13943 (N_13943,N_12554,N_12411);
and U13944 (N_13944,N_12172,N_12476);
nand U13945 (N_13945,N_12978,N_12474);
and U13946 (N_13946,N_12794,N_12114);
nor U13947 (N_13947,N_12602,N_12354);
xor U13948 (N_13948,N_12970,N_12453);
xnor U13949 (N_13949,N_12099,N_12420);
nand U13950 (N_13950,N_12363,N_12039);
and U13951 (N_13951,N_12567,N_12480);
nor U13952 (N_13952,N_12947,N_12288);
xnor U13953 (N_13953,N_12202,N_12756);
xor U13954 (N_13954,N_12973,N_12511);
or U13955 (N_13955,N_12433,N_12559);
nor U13956 (N_13956,N_12169,N_12822);
xor U13957 (N_13957,N_12118,N_12442);
or U13958 (N_13958,N_12047,N_12183);
and U13959 (N_13959,N_12184,N_12383);
xnor U13960 (N_13960,N_12432,N_12281);
nand U13961 (N_13961,N_12501,N_12506);
and U13962 (N_13962,N_12079,N_12398);
or U13963 (N_13963,N_12119,N_12622);
and U13964 (N_13964,N_12063,N_12671);
nor U13965 (N_13965,N_12680,N_12173);
nand U13966 (N_13966,N_12094,N_12359);
nand U13967 (N_13967,N_12247,N_12305);
nand U13968 (N_13968,N_12403,N_12849);
nand U13969 (N_13969,N_12339,N_12017);
nand U13970 (N_13970,N_12439,N_12751);
or U13971 (N_13971,N_12357,N_12633);
nand U13972 (N_13972,N_12031,N_12767);
nand U13973 (N_13973,N_12029,N_12775);
nor U13974 (N_13974,N_12541,N_12222);
and U13975 (N_13975,N_12385,N_12699);
xor U13976 (N_13976,N_12826,N_12724);
nand U13977 (N_13977,N_12117,N_12328);
or U13978 (N_13978,N_12885,N_12834);
nor U13979 (N_13979,N_12815,N_12436);
nor U13980 (N_13980,N_12622,N_12331);
nor U13981 (N_13981,N_12574,N_12997);
nand U13982 (N_13982,N_12713,N_12577);
nor U13983 (N_13983,N_12202,N_12736);
nor U13984 (N_13984,N_12356,N_12494);
nand U13985 (N_13985,N_12221,N_12047);
and U13986 (N_13986,N_12564,N_12766);
xor U13987 (N_13987,N_12609,N_12619);
xnor U13988 (N_13988,N_12773,N_12670);
nor U13989 (N_13989,N_12692,N_12327);
xnor U13990 (N_13990,N_12445,N_12917);
or U13991 (N_13991,N_12409,N_12897);
nand U13992 (N_13992,N_12687,N_12607);
nand U13993 (N_13993,N_12958,N_12903);
nor U13994 (N_13994,N_12291,N_12591);
nand U13995 (N_13995,N_12952,N_12988);
nand U13996 (N_13996,N_12688,N_12832);
or U13997 (N_13997,N_12362,N_12230);
nand U13998 (N_13998,N_12130,N_12110);
nor U13999 (N_13999,N_12336,N_12115);
and U14000 (N_14000,N_13868,N_13967);
and U14001 (N_14001,N_13039,N_13140);
and U14002 (N_14002,N_13564,N_13435);
xor U14003 (N_14003,N_13160,N_13365);
or U14004 (N_14004,N_13956,N_13811);
nor U14005 (N_14005,N_13580,N_13534);
and U14006 (N_14006,N_13567,N_13029);
xor U14007 (N_14007,N_13621,N_13082);
and U14008 (N_14008,N_13429,N_13581);
or U14009 (N_14009,N_13069,N_13838);
nand U14010 (N_14010,N_13068,N_13458);
and U14011 (N_14011,N_13338,N_13497);
xor U14012 (N_14012,N_13561,N_13477);
xor U14013 (N_14013,N_13236,N_13329);
or U14014 (N_14014,N_13305,N_13856);
nand U14015 (N_14015,N_13638,N_13326);
or U14016 (N_14016,N_13512,N_13387);
xor U14017 (N_14017,N_13414,N_13912);
nor U14018 (N_14018,N_13297,N_13415);
nor U14019 (N_14019,N_13559,N_13055);
nand U14020 (N_14020,N_13404,N_13177);
nand U14021 (N_14021,N_13438,N_13010);
nor U14022 (N_14022,N_13363,N_13593);
or U14023 (N_14023,N_13900,N_13149);
nor U14024 (N_14024,N_13601,N_13257);
nand U14025 (N_14025,N_13196,N_13301);
nor U14026 (N_14026,N_13883,N_13375);
nand U14027 (N_14027,N_13949,N_13131);
or U14028 (N_14028,N_13396,N_13841);
nand U14029 (N_14029,N_13430,N_13507);
or U14030 (N_14030,N_13065,N_13427);
xnor U14031 (N_14031,N_13339,N_13631);
nor U14032 (N_14032,N_13061,N_13416);
nor U14033 (N_14033,N_13393,N_13103);
xor U14034 (N_14034,N_13522,N_13848);
xnor U14035 (N_14035,N_13726,N_13732);
xnor U14036 (N_14036,N_13734,N_13645);
or U14037 (N_14037,N_13144,N_13366);
nor U14038 (N_14038,N_13816,N_13007);
nand U14039 (N_14039,N_13179,N_13235);
xnor U14040 (N_14040,N_13148,N_13186);
xnor U14041 (N_14041,N_13536,N_13907);
xor U14042 (N_14042,N_13939,N_13314);
or U14043 (N_14043,N_13048,N_13440);
or U14044 (N_14044,N_13938,N_13716);
nand U14045 (N_14045,N_13964,N_13112);
or U14046 (N_14046,N_13209,N_13199);
xnor U14047 (N_14047,N_13099,N_13596);
or U14048 (N_14048,N_13192,N_13860);
or U14049 (N_14049,N_13303,N_13268);
nor U14050 (N_14050,N_13422,N_13506);
or U14051 (N_14051,N_13897,N_13359);
or U14052 (N_14052,N_13189,N_13764);
or U14053 (N_14053,N_13398,N_13541);
or U14054 (N_14054,N_13434,N_13740);
nand U14055 (N_14055,N_13976,N_13935);
or U14056 (N_14056,N_13532,N_13118);
nand U14057 (N_14057,N_13827,N_13796);
or U14058 (N_14058,N_13977,N_13970);
nand U14059 (N_14059,N_13328,N_13805);
and U14060 (N_14060,N_13143,N_13552);
or U14061 (N_14061,N_13558,N_13606);
nor U14062 (N_14062,N_13218,N_13470);
nor U14063 (N_14063,N_13091,N_13480);
nor U14064 (N_14064,N_13300,N_13521);
nand U14065 (N_14065,N_13624,N_13701);
and U14066 (N_14066,N_13000,N_13687);
nor U14067 (N_14067,N_13066,N_13159);
nand U14068 (N_14068,N_13643,N_13498);
nor U14069 (N_14069,N_13439,N_13028);
nor U14070 (N_14070,N_13667,N_13685);
nand U14071 (N_14071,N_13854,N_13153);
and U14072 (N_14072,N_13200,N_13490);
xnor U14073 (N_14073,N_13244,N_13336);
and U14074 (N_14074,N_13281,N_13736);
or U14075 (N_14075,N_13808,N_13527);
xor U14076 (N_14076,N_13382,N_13250);
and U14077 (N_14077,N_13731,N_13261);
nor U14078 (N_14078,N_13745,N_13707);
and U14079 (N_14079,N_13931,N_13096);
nand U14080 (N_14080,N_13960,N_13651);
and U14081 (N_14081,N_13571,N_13446);
nand U14082 (N_14082,N_13230,N_13557);
and U14083 (N_14083,N_13934,N_13425);
or U14084 (N_14084,N_13830,N_13377);
xor U14085 (N_14085,N_13990,N_13284);
nor U14086 (N_14086,N_13248,N_13290);
or U14087 (N_14087,N_13993,N_13341);
and U14088 (N_14088,N_13587,N_13744);
xor U14089 (N_14089,N_13699,N_13962);
xor U14090 (N_14090,N_13482,N_13285);
and U14091 (N_14091,N_13892,N_13602);
or U14092 (N_14092,N_13881,N_13979);
and U14093 (N_14093,N_13893,N_13968);
or U14094 (N_14094,N_13975,N_13465);
nand U14095 (N_14095,N_13421,N_13031);
or U14096 (N_14096,N_13831,N_13171);
nand U14097 (N_14097,N_13861,N_13533);
nor U14098 (N_14098,N_13198,N_13663);
and U14099 (N_14099,N_13965,N_13972);
xor U14100 (N_14100,N_13157,N_13346);
nand U14101 (N_14101,N_13100,N_13319);
nand U14102 (N_14102,N_13666,N_13870);
nor U14103 (N_14103,N_13670,N_13635);
xnor U14104 (N_14104,N_13193,N_13455);
xnor U14105 (N_14105,N_13879,N_13202);
xor U14106 (N_14106,N_13494,N_13582);
nor U14107 (N_14107,N_13272,N_13683);
xnor U14108 (N_14108,N_13735,N_13703);
or U14109 (N_14109,N_13087,N_13604);
nand U14110 (N_14110,N_13768,N_13927);
xor U14111 (N_14111,N_13542,N_13511);
and U14112 (N_14112,N_13992,N_13971);
xnor U14113 (N_14113,N_13226,N_13932);
xor U14114 (N_14114,N_13344,N_13400);
nand U14115 (N_14115,N_13043,N_13672);
nand U14116 (N_14116,N_13980,N_13008);
xnor U14117 (N_14117,N_13508,N_13334);
and U14118 (N_14118,N_13361,N_13570);
or U14119 (N_14119,N_13201,N_13169);
nor U14120 (N_14120,N_13929,N_13839);
xnor U14121 (N_14121,N_13545,N_13933);
nor U14122 (N_14122,N_13682,N_13517);
and U14123 (N_14123,N_13943,N_13655);
nand U14124 (N_14124,N_13443,N_13516);
xnor U14125 (N_14125,N_13484,N_13013);
nand U14126 (N_14126,N_13018,N_13674);
nand U14127 (N_14127,N_13969,N_13546);
or U14128 (N_14128,N_13575,N_13504);
nand U14129 (N_14129,N_13080,N_13766);
nand U14130 (N_14130,N_13821,N_13036);
nor U14131 (N_14131,N_13114,N_13260);
or U14132 (N_14132,N_13899,N_13024);
xnor U14133 (N_14133,N_13001,N_13307);
xor U14134 (N_14134,N_13941,N_13801);
nor U14135 (N_14135,N_13865,N_13641);
nor U14136 (N_14136,N_13763,N_13875);
nor U14137 (N_14137,N_13926,N_13626);
xor U14138 (N_14138,N_13151,N_13106);
xnor U14139 (N_14139,N_13468,N_13316);
nor U14140 (N_14140,N_13167,N_13973);
xor U14141 (N_14141,N_13137,N_13524);
or U14142 (N_14142,N_13397,N_13921);
xor U14143 (N_14143,N_13788,N_13798);
or U14144 (N_14144,N_13963,N_13503);
and U14145 (N_14145,N_13660,N_13249);
or U14146 (N_14146,N_13864,N_13646);
or U14147 (N_14147,N_13806,N_13640);
xnor U14148 (N_14148,N_13676,N_13991);
nor U14149 (N_14149,N_13915,N_13647);
and U14150 (N_14150,N_13882,N_13610);
xor U14151 (N_14151,N_13355,N_13771);
and U14152 (N_14152,N_13364,N_13077);
nor U14153 (N_14153,N_13350,N_13042);
nand U14154 (N_14154,N_13231,N_13928);
nor U14155 (N_14155,N_13324,N_13951);
xor U14156 (N_14156,N_13020,N_13320);
nor U14157 (N_14157,N_13576,N_13616);
nor U14158 (N_14158,N_13110,N_13239);
or U14159 (N_14159,N_13653,N_13862);
nand U14160 (N_14160,N_13431,N_13697);
nor U14161 (N_14161,N_13543,N_13608);
xnor U14162 (N_14162,N_13067,N_13502);
nor U14163 (N_14163,N_13011,N_13003);
or U14164 (N_14164,N_13267,N_13483);
nor U14165 (N_14165,N_13183,N_13277);
nand U14166 (N_14166,N_13617,N_13051);
or U14167 (N_14167,N_13254,N_13588);
nand U14168 (N_14168,N_13733,N_13259);
and U14169 (N_14169,N_13591,N_13221);
and U14170 (N_14170,N_13781,N_13867);
and U14171 (N_14171,N_13690,N_13479);
or U14172 (N_14172,N_13327,N_13182);
nand U14173 (N_14173,N_13444,N_13211);
nor U14174 (N_14174,N_13367,N_13126);
nor U14175 (N_14175,N_13419,N_13911);
nand U14176 (N_14176,N_13717,N_13692);
or U14177 (N_14177,N_13460,N_13715);
or U14178 (N_14178,N_13563,N_13293);
nand U14179 (N_14179,N_13292,N_13168);
or U14180 (N_14180,N_13037,N_13729);
nand U14181 (N_14181,N_13813,N_13252);
xor U14182 (N_14182,N_13850,N_13820);
and U14183 (N_14183,N_13513,N_13652);
xor U14184 (N_14184,N_13358,N_13026);
nor U14185 (N_14185,N_13548,N_13578);
xor U14186 (N_14186,N_13410,N_13266);
nand U14187 (N_14187,N_13150,N_13019);
xnor U14188 (N_14188,N_13695,N_13306);
nand U14189 (N_14189,N_13311,N_13680);
or U14190 (N_14190,N_13691,N_13442);
xnor U14191 (N_14191,N_13214,N_13485);
and U14192 (N_14192,N_13313,N_13174);
and U14193 (N_14193,N_13714,N_13902);
and U14194 (N_14194,N_13905,N_13343);
xor U14195 (N_14195,N_13573,N_13718);
nor U14196 (N_14196,N_13073,N_13467);
and U14197 (N_14197,N_13185,N_13197);
xnor U14198 (N_14198,N_13023,N_13913);
nor U14199 (N_14199,N_13722,N_13823);
xnor U14200 (N_14200,N_13079,N_13255);
nor U14201 (N_14201,N_13594,N_13510);
and U14202 (N_14202,N_13794,N_13920);
xnor U14203 (N_14203,N_13111,N_13321);
xnor U14204 (N_14204,N_13188,N_13923);
nor U14205 (N_14205,N_13749,N_13030);
xnor U14206 (N_14206,N_13139,N_13476);
or U14207 (N_14207,N_13609,N_13296);
and U14208 (N_14208,N_13166,N_13471);
nor U14209 (N_14209,N_13611,N_13180);
nand U14210 (N_14210,N_13946,N_13352);
nor U14211 (N_14211,N_13090,N_13402);
and U14212 (N_14212,N_13605,N_13147);
nor U14213 (N_14213,N_13988,N_13287);
nor U14214 (N_14214,N_13787,N_13017);
xor U14215 (N_14215,N_13793,N_13345);
or U14216 (N_14216,N_13424,N_13800);
xor U14217 (N_14217,N_13280,N_13368);
and U14218 (N_14218,N_13819,N_13241);
nor U14219 (N_14219,N_13961,N_13413);
or U14220 (N_14220,N_13756,N_13493);
and U14221 (N_14221,N_13256,N_13299);
xor U14222 (N_14222,N_13728,N_13629);
xnor U14223 (N_14223,N_13496,N_13906);
or U14224 (N_14224,N_13032,N_13776);
nand U14225 (N_14225,N_13176,N_13360);
xnor U14226 (N_14226,N_13620,N_13987);
nand U14227 (N_14227,N_13273,N_13531);
nand U14228 (N_14228,N_13187,N_13644);
and U14229 (N_14229,N_13549,N_13041);
xor U14230 (N_14230,N_13371,N_13084);
nand U14231 (N_14231,N_13837,N_13812);
nand U14232 (N_14232,N_13857,N_13308);
and U14233 (N_14233,N_13288,N_13136);
xnor U14234 (N_14234,N_13799,N_13262);
or U14235 (N_14235,N_13206,N_13050);
or U14236 (N_14236,N_13062,N_13283);
or U14237 (N_14237,N_13121,N_13642);
xor U14238 (N_14238,N_13705,N_13163);
xor U14239 (N_14239,N_13228,N_13386);
nor U14240 (N_14240,N_13165,N_13803);
xor U14241 (N_14241,N_13625,N_13270);
or U14242 (N_14242,N_13599,N_13027);
nand U14243 (N_14243,N_13782,N_13618);
nand U14244 (N_14244,N_13098,N_13779);
and U14245 (N_14245,N_13145,N_13903);
or U14246 (N_14246,N_13488,N_13790);
nand U14247 (N_14247,N_13922,N_13072);
and U14248 (N_14248,N_13770,N_13217);
nor U14249 (N_14249,N_13040,N_13322);
and U14250 (N_14250,N_13785,N_13562);
nor U14251 (N_14251,N_13886,N_13381);
nor U14252 (N_14252,N_13727,N_13401);
nand U14253 (N_14253,N_13457,N_13614);
nor U14254 (N_14254,N_13983,N_13526);
nor U14255 (N_14255,N_13632,N_13373);
nand U14256 (N_14256,N_13792,N_13279);
nor U14257 (N_14257,N_13528,N_13223);
nor U14258 (N_14258,N_13950,N_13627);
and U14259 (N_14259,N_13464,N_13958);
xnor U14260 (N_14260,N_13135,N_13658);
and U14261 (N_14261,N_13021,N_13351);
and U14262 (N_14262,N_13170,N_13725);
nor U14263 (N_14263,N_13432,N_13994);
xor U14264 (N_14264,N_13234,N_13751);
nand U14265 (N_14265,N_13298,N_13407);
nand U14266 (N_14266,N_13577,N_13895);
xnor U14267 (N_14267,N_13639,N_13681);
nand U14268 (N_14268,N_13203,N_13125);
xor U14269 (N_14269,N_13849,N_13896);
nand U14270 (N_14270,N_13124,N_13156);
nand U14271 (N_14271,N_13275,N_13889);
xor U14272 (N_14272,N_13797,N_13761);
or U14273 (N_14273,N_13141,N_13450);
or U14274 (N_14274,N_13678,N_13649);
or U14275 (N_14275,N_13105,N_13089);
xnor U14276 (N_14276,N_13569,N_13673);
and U14277 (N_14277,N_13686,N_13172);
or U14278 (N_14278,N_13677,N_13843);
nor U14279 (N_14279,N_13748,N_13216);
xor U14280 (N_14280,N_13721,N_13757);
xor U14281 (N_14281,N_13544,N_13737);
or U14282 (N_14282,N_13108,N_13671);
nor U14283 (N_14283,N_13006,N_13064);
xnor U14284 (N_14284,N_13773,N_13370);
nand U14285 (N_14285,N_13815,N_13357);
and U14286 (N_14286,N_13826,N_13974);
nand U14287 (N_14287,N_13762,N_13390);
nand U14288 (N_14288,N_13847,N_13403);
xnor U14289 (N_14289,N_13989,N_13910);
xor U14290 (N_14290,N_13063,N_13132);
nor U14291 (N_14291,N_13173,N_13804);
and U14292 (N_14292,N_13774,N_13161);
or U14293 (N_14293,N_13904,N_13583);
and U14294 (N_14294,N_13878,N_13128);
and U14295 (N_14295,N_13858,N_13122);
or U14296 (N_14296,N_13219,N_13780);
nand U14297 (N_14297,N_13754,N_13117);
nor U14298 (N_14298,N_13984,N_13955);
nor U14299 (N_14299,N_13784,N_13380);
nand U14300 (N_14300,N_13679,N_13835);
or U14301 (N_14301,N_13750,N_13769);
nand U14302 (N_14302,N_13713,N_13809);
or U14303 (N_14303,N_13081,N_13999);
xnor U14304 (N_14304,N_13129,N_13551);
and U14305 (N_14305,N_13636,N_13675);
nand U14306 (N_14306,N_13709,N_13693);
xnor U14307 (N_14307,N_13225,N_13501);
nor U14308 (N_14308,N_13842,N_13489);
or U14309 (N_14309,N_13741,N_13391);
nor U14310 (N_14310,N_13918,N_13840);
xor U14311 (N_14311,N_13786,N_13207);
and U14312 (N_14312,N_13925,N_13312);
or U14313 (N_14313,N_13613,N_13901);
nor U14314 (N_14314,N_13395,N_13592);
or U14315 (N_14315,N_13948,N_13474);
and U14316 (N_14316,N_13509,N_13863);
and U14317 (N_14317,N_13116,N_13995);
and U14318 (N_14318,N_13997,N_13333);
and U14319 (N_14319,N_13451,N_13190);
and U14320 (N_14320,N_13238,N_13874);
nor U14321 (N_14321,N_13331,N_13409);
nand U14322 (N_14322,N_13940,N_13550);
nand U14323 (N_14323,N_13585,N_13224);
or U14324 (N_14324,N_13520,N_13689);
and U14325 (N_14325,N_13227,N_13565);
and U14326 (N_14326,N_13323,N_13612);
xor U14327 (N_14327,N_13454,N_13572);
xor U14328 (N_14328,N_13095,N_13747);
and U14329 (N_14329,N_13109,N_13383);
xnor U14330 (N_14330,N_13579,N_13406);
nor U14331 (N_14331,N_13466,N_13120);
nor U14332 (N_14332,N_13500,N_13828);
xor U14333 (N_14333,N_13852,N_13832);
nand U14334 (N_14334,N_13184,N_13978);
nand U14335 (N_14335,N_13589,N_13146);
nand U14336 (N_14336,N_13758,N_13208);
xor U14337 (N_14337,N_13392,N_13362);
nor U14338 (N_14338,N_13834,N_13891);
nor U14339 (N_14339,N_13034,N_13046);
nor U14340 (N_14340,N_13447,N_13634);
or U14341 (N_14341,N_13514,N_13047);
nor U14342 (N_14342,N_13659,N_13093);
nand U14343 (N_14343,N_13487,N_13560);
nand U14344 (N_14344,N_13282,N_13515);
xnor U14345 (N_14345,N_13668,N_13452);
nor U14346 (N_14346,N_13818,N_13075);
nor U14347 (N_14347,N_13724,N_13518);
nor U14348 (N_14348,N_13278,N_13265);
xnor U14349 (N_14349,N_13795,N_13271);
or U14350 (N_14350,N_13428,N_13952);
xor U14351 (N_14351,N_13142,N_13720);
or U14352 (N_14352,N_13154,N_13730);
xnor U14353 (N_14353,N_13083,N_13449);
nand U14354 (N_14354,N_13092,N_13872);
or U14355 (N_14355,N_13783,N_13240);
nor U14356 (N_14356,N_13535,N_13930);
or U14357 (N_14357,N_13855,N_13369);
or U14358 (N_14358,N_13085,N_13309);
nor U14359 (N_14359,N_13702,N_13162);
or U14360 (N_14360,N_13059,N_13937);
or U14361 (N_14361,N_13547,N_13824);
and U14362 (N_14362,N_13752,N_13453);
xnor U14363 (N_14363,N_13302,N_13742);
and U14364 (N_14364,N_13719,N_13388);
nand U14365 (N_14365,N_13982,N_13251);
and U14366 (N_14366,N_13802,N_13127);
xnor U14367 (N_14367,N_13845,N_13539);
or U14368 (N_14368,N_13775,N_13945);
and U14369 (N_14369,N_13708,N_13492);
or U14370 (N_14370,N_13853,N_13335);
and U14371 (N_14371,N_13372,N_13330);
nand U14372 (N_14372,N_13405,N_13071);
xnor U14373 (N_14373,N_13657,N_13220);
or U14374 (N_14374,N_13789,N_13760);
xor U14375 (N_14375,N_13505,N_13423);
nor U14376 (N_14376,N_13684,N_13204);
nor U14377 (N_14377,N_13871,N_13134);
xnor U14378 (N_14378,N_13607,N_13035);
xor U14379 (N_14379,N_13374,N_13191);
xnor U14380 (N_14380,N_13101,N_13130);
or U14381 (N_14381,N_13195,N_13253);
nand U14382 (N_14382,N_13461,N_13807);
nor U14383 (N_14383,N_13650,N_13002);
or U14384 (N_14384,N_13817,N_13499);
and U14385 (N_14385,N_13998,N_13337);
or U14386 (N_14386,N_13243,N_13033);
nand U14387 (N_14387,N_13877,N_13175);
nor U14388 (N_14388,N_13615,N_13245);
or U14389 (N_14389,N_13222,N_13537);
nor U14390 (N_14390,N_13595,N_13833);
nand U14391 (N_14391,N_13586,N_13056);
nor U14392 (N_14392,N_13481,N_13078);
xnor U14393 (N_14393,N_13060,N_13022);
nand U14394 (N_14394,N_13264,N_13349);
or U14395 (N_14395,N_13590,N_13661);
nand U14396 (N_14396,N_13304,N_13986);
xnor U14397 (N_14397,N_13574,N_13418);
or U14398 (N_14398,N_13389,N_13158);
and U14399 (N_14399,N_13584,N_13263);
or U14400 (N_14400,N_13669,N_13530);
and U14401 (N_14401,N_13469,N_13908);
xor U14402 (N_14402,N_13985,N_13884);
or U14403 (N_14403,N_13025,N_13665);
or U14404 (N_14404,N_13437,N_13996);
or U14405 (N_14405,N_13767,N_13045);
xor U14406 (N_14406,N_13623,N_13814);
nand U14407 (N_14407,N_13354,N_13472);
or U14408 (N_14408,N_13957,N_13825);
and U14409 (N_14409,N_13894,N_13164);
nand U14410 (N_14410,N_13523,N_13851);
nand U14411 (N_14411,N_13739,N_13212);
and U14412 (N_14412,N_13286,N_13866);
xor U14413 (N_14413,N_13755,N_13213);
and U14414 (N_14414,N_13917,N_13876);
nand U14415 (N_14415,N_13556,N_13919);
nand U14416 (N_14416,N_13529,N_13538);
nor U14417 (N_14417,N_13005,N_13981);
or U14418 (N_14418,N_13597,N_13294);
nand U14419 (N_14419,N_13412,N_13936);
nand U14420 (N_14420,N_13743,N_13696);
and U14421 (N_14421,N_13274,N_13791);
or U14422 (N_14422,N_13869,N_13247);
nand U14423 (N_14423,N_13016,N_13553);
xor U14424 (N_14424,N_13568,N_13246);
or U14425 (N_14425,N_13654,N_13598);
or U14426 (N_14426,N_13094,N_13276);
nor U14427 (N_14427,N_13408,N_13347);
nand U14428 (N_14428,N_13317,N_13233);
nor U14429 (N_14429,N_13829,N_13566);
xor U14430 (N_14430,N_13258,N_13074);
nor U14431 (N_14431,N_13778,N_13325);
nor U14432 (N_14432,N_13014,N_13097);
or U14433 (N_14433,N_13698,N_13229);
xor U14434 (N_14434,N_13420,N_13107);
nor U14435 (N_14435,N_13310,N_13916);
nand U14436 (N_14436,N_13909,N_13953);
nor U14437 (N_14437,N_13711,N_13712);
xnor U14438 (N_14438,N_13318,N_13822);
and U14439 (N_14439,N_13242,N_13890);
or U14440 (N_14440,N_13104,N_13656);
nand U14441 (N_14441,N_13070,N_13810);
or U14442 (N_14442,N_13436,N_13630);
xnor U14443 (N_14443,N_13295,N_13012);
and U14444 (N_14444,N_13898,N_13269);
and U14445 (N_14445,N_13633,N_13688);
and U14446 (N_14446,N_13205,N_13888);
xor U14447 (N_14447,N_13411,N_13628);
nand U14448 (N_14448,N_13215,N_13088);
or U14449 (N_14449,N_13765,N_13340);
xor U14450 (N_14450,N_13947,N_13704);
xor U14451 (N_14451,N_13194,N_13119);
xor U14452 (N_14452,N_13706,N_13049);
nor U14453 (N_14453,N_13057,N_13753);
and U14454 (N_14454,N_13417,N_13746);
nand U14455 (N_14455,N_13426,N_13448);
nand U14456 (N_14456,N_13459,N_13475);
xnor U14457 (N_14457,N_13723,N_13959);
or U14458 (N_14458,N_13495,N_13473);
nand U14459 (N_14459,N_13378,N_13237);
nor U14460 (N_14460,N_13015,N_13846);
nand U14461 (N_14461,N_13954,N_13738);
or U14462 (N_14462,N_13619,N_13491);
and U14463 (N_14463,N_13859,N_13942);
or U14464 (N_14464,N_13445,N_13873);
nand U14465 (N_14465,N_13054,N_13966);
nor U14466 (N_14466,N_13836,N_13885);
nor U14467 (N_14467,N_13210,N_13053);
nor U14468 (N_14468,N_13662,N_13777);
xor U14469 (N_14469,N_13133,N_13710);
or U14470 (N_14470,N_13944,N_13622);
and U14471 (N_14471,N_13555,N_13044);
xor U14472 (N_14472,N_13887,N_13058);
nand U14473 (N_14473,N_13759,N_13356);
nor U14474 (N_14474,N_13463,N_13115);
nor U14475 (N_14475,N_13462,N_13181);
nor U14476 (N_14476,N_13384,N_13554);
nand U14477 (N_14477,N_13441,N_13376);
xor U14478 (N_14478,N_13700,N_13694);
or U14479 (N_14479,N_13844,N_13332);
nor U14480 (N_14480,N_13603,N_13433);
xnor U14481 (N_14481,N_13289,N_13102);
nor U14482 (N_14482,N_13664,N_13648);
or U14483 (N_14483,N_13152,N_13379);
and U14484 (N_14484,N_13772,N_13637);
xor U14485 (N_14485,N_13004,N_13155);
nand U14486 (N_14486,N_13394,N_13385);
nand U14487 (N_14487,N_13315,N_13038);
nor U14488 (N_14488,N_13353,N_13525);
nand U14489 (N_14489,N_13086,N_13342);
and U14490 (N_14490,N_13123,N_13052);
or U14491 (N_14491,N_13113,N_13009);
and U14492 (N_14492,N_13348,N_13540);
nor U14493 (N_14493,N_13178,N_13399);
nand U14494 (N_14494,N_13138,N_13232);
and U14495 (N_14495,N_13924,N_13076);
or U14496 (N_14496,N_13600,N_13914);
xnor U14497 (N_14497,N_13456,N_13519);
nand U14498 (N_14498,N_13291,N_13486);
or U14499 (N_14499,N_13478,N_13880);
or U14500 (N_14500,N_13196,N_13727);
nor U14501 (N_14501,N_13885,N_13141);
nor U14502 (N_14502,N_13854,N_13109);
nand U14503 (N_14503,N_13199,N_13767);
or U14504 (N_14504,N_13696,N_13999);
and U14505 (N_14505,N_13907,N_13365);
xnor U14506 (N_14506,N_13182,N_13181);
or U14507 (N_14507,N_13568,N_13418);
or U14508 (N_14508,N_13823,N_13701);
nand U14509 (N_14509,N_13500,N_13936);
or U14510 (N_14510,N_13665,N_13122);
xnor U14511 (N_14511,N_13703,N_13305);
or U14512 (N_14512,N_13379,N_13544);
nor U14513 (N_14513,N_13035,N_13820);
xor U14514 (N_14514,N_13932,N_13479);
nand U14515 (N_14515,N_13397,N_13312);
nor U14516 (N_14516,N_13455,N_13221);
nand U14517 (N_14517,N_13259,N_13347);
nor U14518 (N_14518,N_13099,N_13101);
and U14519 (N_14519,N_13596,N_13773);
xnor U14520 (N_14520,N_13326,N_13521);
and U14521 (N_14521,N_13368,N_13008);
nor U14522 (N_14522,N_13295,N_13740);
or U14523 (N_14523,N_13017,N_13993);
xnor U14524 (N_14524,N_13358,N_13873);
nand U14525 (N_14525,N_13199,N_13002);
or U14526 (N_14526,N_13612,N_13235);
or U14527 (N_14527,N_13742,N_13342);
and U14528 (N_14528,N_13324,N_13865);
or U14529 (N_14529,N_13243,N_13159);
xnor U14530 (N_14530,N_13040,N_13419);
nor U14531 (N_14531,N_13358,N_13014);
nand U14532 (N_14532,N_13829,N_13076);
xnor U14533 (N_14533,N_13724,N_13201);
or U14534 (N_14534,N_13141,N_13076);
nor U14535 (N_14535,N_13333,N_13844);
nand U14536 (N_14536,N_13525,N_13195);
or U14537 (N_14537,N_13960,N_13091);
and U14538 (N_14538,N_13484,N_13768);
nand U14539 (N_14539,N_13107,N_13859);
nor U14540 (N_14540,N_13534,N_13240);
nand U14541 (N_14541,N_13259,N_13026);
nor U14542 (N_14542,N_13809,N_13331);
nor U14543 (N_14543,N_13358,N_13235);
or U14544 (N_14544,N_13510,N_13806);
nand U14545 (N_14545,N_13265,N_13071);
or U14546 (N_14546,N_13759,N_13484);
nor U14547 (N_14547,N_13817,N_13559);
nor U14548 (N_14548,N_13255,N_13671);
and U14549 (N_14549,N_13630,N_13660);
nor U14550 (N_14550,N_13990,N_13155);
nand U14551 (N_14551,N_13269,N_13983);
nand U14552 (N_14552,N_13359,N_13414);
xnor U14553 (N_14553,N_13841,N_13776);
or U14554 (N_14554,N_13951,N_13419);
nor U14555 (N_14555,N_13581,N_13333);
nand U14556 (N_14556,N_13928,N_13562);
nor U14557 (N_14557,N_13296,N_13042);
xnor U14558 (N_14558,N_13352,N_13754);
nor U14559 (N_14559,N_13075,N_13663);
and U14560 (N_14560,N_13053,N_13264);
nor U14561 (N_14561,N_13304,N_13083);
xnor U14562 (N_14562,N_13749,N_13741);
and U14563 (N_14563,N_13957,N_13349);
xnor U14564 (N_14564,N_13632,N_13905);
nor U14565 (N_14565,N_13006,N_13024);
and U14566 (N_14566,N_13622,N_13236);
xnor U14567 (N_14567,N_13091,N_13313);
nand U14568 (N_14568,N_13054,N_13020);
nand U14569 (N_14569,N_13156,N_13056);
xor U14570 (N_14570,N_13891,N_13051);
and U14571 (N_14571,N_13591,N_13401);
and U14572 (N_14572,N_13768,N_13556);
xor U14573 (N_14573,N_13446,N_13898);
or U14574 (N_14574,N_13126,N_13037);
xnor U14575 (N_14575,N_13613,N_13049);
or U14576 (N_14576,N_13627,N_13076);
and U14577 (N_14577,N_13037,N_13071);
xor U14578 (N_14578,N_13052,N_13669);
and U14579 (N_14579,N_13134,N_13238);
nand U14580 (N_14580,N_13592,N_13761);
xnor U14581 (N_14581,N_13323,N_13165);
and U14582 (N_14582,N_13399,N_13417);
nand U14583 (N_14583,N_13751,N_13976);
xor U14584 (N_14584,N_13176,N_13236);
or U14585 (N_14585,N_13240,N_13866);
and U14586 (N_14586,N_13167,N_13926);
xnor U14587 (N_14587,N_13744,N_13953);
xor U14588 (N_14588,N_13868,N_13957);
nor U14589 (N_14589,N_13864,N_13329);
xor U14590 (N_14590,N_13161,N_13077);
nor U14591 (N_14591,N_13501,N_13803);
or U14592 (N_14592,N_13109,N_13839);
nand U14593 (N_14593,N_13369,N_13270);
xnor U14594 (N_14594,N_13525,N_13755);
or U14595 (N_14595,N_13457,N_13937);
xnor U14596 (N_14596,N_13048,N_13694);
or U14597 (N_14597,N_13593,N_13786);
nor U14598 (N_14598,N_13898,N_13173);
nor U14599 (N_14599,N_13363,N_13985);
nand U14600 (N_14600,N_13906,N_13759);
xor U14601 (N_14601,N_13483,N_13106);
xor U14602 (N_14602,N_13426,N_13670);
and U14603 (N_14603,N_13445,N_13482);
or U14604 (N_14604,N_13872,N_13190);
nand U14605 (N_14605,N_13978,N_13228);
and U14606 (N_14606,N_13947,N_13562);
and U14607 (N_14607,N_13866,N_13205);
nand U14608 (N_14608,N_13013,N_13933);
nand U14609 (N_14609,N_13564,N_13292);
xnor U14610 (N_14610,N_13748,N_13064);
nor U14611 (N_14611,N_13583,N_13100);
nand U14612 (N_14612,N_13413,N_13998);
nand U14613 (N_14613,N_13352,N_13853);
or U14614 (N_14614,N_13672,N_13158);
nor U14615 (N_14615,N_13835,N_13284);
nand U14616 (N_14616,N_13667,N_13073);
and U14617 (N_14617,N_13607,N_13371);
nor U14618 (N_14618,N_13232,N_13403);
xnor U14619 (N_14619,N_13217,N_13079);
or U14620 (N_14620,N_13989,N_13274);
and U14621 (N_14621,N_13077,N_13010);
and U14622 (N_14622,N_13516,N_13779);
xnor U14623 (N_14623,N_13608,N_13045);
nand U14624 (N_14624,N_13743,N_13317);
xnor U14625 (N_14625,N_13388,N_13515);
and U14626 (N_14626,N_13421,N_13114);
or U14627 (N_14627,N_13395,N_13276);
xor U14628 (N_14628,N_13854,N_13396);
nand U14629 (N_14629,N_13154,N_13365);
and U14630 (N_14630,N_13902,N_13756);
xor U14631 (N_14631,N_13026,N_13565);
and U14632 (N_14632,N_13154,N_13053);
xor U14633 (N_14633,N_13328,N_13031);
and U14634 (N_14634,N_13314,N_13854);
nor U14635 (N_14635,N_13236,N_13898);
xor U14636 (N_14636,N_13947,N_13064);
or U14637 (N_14637,N_13610,N_13181);
or U14638 (N_14638,N_13023,N_13806);
nand U14639 (N_14639,N_13080,N_13901);
xor U14640 (N_14640,N_13627,N_13679);
nand U14641 (N_14641,N_13678,N_13585);
xor U14642 (N_14642,N_13438,N_13425);
or U14643 (N_14643,N_13572,N_13037);
xnor U14644 (N_14644,N_13808,N_13662);
or U14645 (N_14645,N_13607,N_13865);
nand U14646 (N_14646,N_13569,N_13141);
nand U14647 (N_14647,N_13044,N_13861);
and U14648 (N_14648,N_13874,N_13339);
or U14649 (N_14649,N_13945,N_13212);
or U14650 (N_14650,N_13989,N_13911);
xor U14651 (N_14651,N_13724,N_13777);
nand U14652 (N_14652,N_13456,N_13336);
xor U14653 (N_14653,N_13808,N_13811);
or U14654 (N_14654,N_13198,N_13214);
xor U14655 (N_14655,N_13240,N_13905);
and U14656 (N_14656,N_13826,N_13316);
nor U14657 (N_14657,N_13440,N_13446);
xor U14658 (N_14658,N_13743,N_13950);
xor U14659 (N_14659,N_13912,N_13944);
xnor U14660 (N_14660,N_13304,N_13854);
or U14661 (N_14661,N_13247,N_13911);
nor U14662 (N_14662,N_13290,N_13845);
and U14663 (N_14663,N_13756,N_13002);
or U14664 (N_14664,N_13429,N_13852);
nand U14665 (N_14665,N_13188,N_13016);
xnor U14666 (N_14666,N_13096,N_13732);
xnor U14667 (N_14667,N_13638,N_13837);
or U14668 (N_14668,N_13649,N_13114);
nand U14669 (N_14669,N_13066,N_13907);
nand U14670 (N_14670,N_13737,N_13927);
nand U14671 (N_14671,N_13782,N_13547);
nor U14672 (N_14672,N_13589,N_13297);
or U14673 (N_14673,N_13624,N_13885);
or U14674 (N_14674,N_13483,N_13663);
and U14675 (N_14675,N_13592,N_13151);
nor U14676 (N_14676,N_13767,N_13280);
or U14677 (N_14677,N_13043,N_13589);
xnor U14678 (N_14678,N_13170,N_13445);
xor U14679 (N_14679,N_13304,N_13858);
xor U14680 (N_14680,N_13399,N_13412);
or U14681 (N_14681,N_13944,N_13465);
or U14682 (N_14682,N_13924,N_13970);
nor U14683 (N_14683,N_13064,N_13166);
or U14684 (N_14684,N_13467,N_13162);
xor U14685 (N_14685,N_13406,N_13904);
or U14686 (N_14686,N_13707,N_13612);
xnor U14687 (N_14687,N_13972,N_13821);
nor U14688 (N_14688,N_13445,N_13566);
or U14689 (N_14689,N_13300,N_13914);
and U14690 (N_14690,N_13672,N_13506);
xnor U14691 (N_14691,N_13065,N_13335);
nand U14692 (N_14692,N_13448,N_13514);
and U14693 (N_14693,N_13266,N_13461);
and U14694 (N_14694,N_13082,N_13672);
or U14695 (N_14695,N_13781,N_13416);
xnor U14696 (N_14696,N_13825,N_13838);
and U14697 (N_14697,N_13472,N_13923);
and U14698 (N_14698,N_13539,N_13163);
and U14699 (N_14699,N_13575,N_13227);
nand U14700 (N_14700,N_13249,N_13850);
nand U14701 (N_14701,N_13304,N_13555);
nand U14702 (N_14702,N_13742,N_13032);
nor U14703 (N_14703,N_13574,N_13086);
xnor U14704 (N_14704,N_13268,N_13110);
xnor U14705 (N_14705,N_13104,N_13633);
xor U14706 (N_14706,N_13154,N_13575);
nand U14707 (N_14707,N_13918,N_13249);
nor U14708 (N_14708,N_13036,N_13798);
nor U14709 (N_14709,N_13150,N_13281);
xor U14710 (N_14710,N_13958,N_13396);
or U14711 (N_14711,N_13019,N_13941);
nor U14712 (N_14712,N_13179,N_13803);
nor U14713 (N_14713,N_13461,N_13588);
nor U14714 (N_14714,N_13226,N_13690);
xor U14715 (N_14715,N_13089,N_13822);
nand U14716 (N_14716,N_13596,N_13944);
nor U14717 (N_14717,N_13042,N_13859);
nor U14718 (N_14718,N_13303,N_13018);
nand U14719 (N_14719,N_13736,N_13810);
and U14720 (N_14720,N_13303,N_13889);
nor U14721 (N_14721,N_13979,N_13659);
nand U14722 (N_14722,N_13754,N_13832);
nand U14723 (N_14723,N_13890,N_13531);
xor U14724 (N_14724,N_13198,N_13046);
nor U14725 (N_14725,N_13210,N_13019);
xor U14726 (N_14726,N_13501,N_13136);
nand U14727 (N_14727,N_13184,N_13180);
and U14728 (N_14728,N_13871,N_13857);
nor U14729 (N_14729,N_13329,N_13219);
xor U14730 (N_14730,N_13338,N_13014);
or U14731 (N_14731,N_13116,N_13853);
or U14732 (N_14732,N_13227,N_13005);
nand U14733 (N_14733,N_13476,N_13851);
xnor U14734 (N_14734,N_13796,N_13323);
xor U14735 (N_14735,N_13095,N_13776);
or U14736 (N_14736,N_13863,N_13319);
nand U14737 (N_14737,N_13335,N_13574);
or U14738 (N_14738,N_13273,N_13511);
and U14739 (N_14739,N_13628,N_13159);
or U14740 (N_14740,N_13434,N_13478);
xor U14741 (N_14741,N_13335,N_13314);
nand U14742 (N_14742,N_13721,N_13910);
and U14743 (N_14743,N_13988,N_13983);
and U14744 (N_14744,N_13396,N_13428);
nand U14745 (N_14745,N_13553,N_13667);
xnor U14746 (N_14746,N_13587,N_13444);
or U14747 (N_14747,N_13616,N_13029);
and U14748 (N_14748,N_13843,N_13344);
nand U14749 (N_14749,N_13410,N_13932);
nand U14750 (N_14750,N_13739,N_13810);
xor U14751 (N_14751,N_13669,N_13208);
or U14752 (N_14752,N_13246,N_13022);
and U14753 (N_14753,N_13083,N_13849);
nor U14754 (N_14754,N_13293,N_13909);
nor U14755 (N_14755,N_13540,N_13732);
xor U14756 (N_14756,N_13839,N_13089);
xnor U14757 (N_14757,N_13537,N_13360);
nor U14758 (N_14758,N_13224,N_13657);
nor U14759 (N_14759,N_13985,N_13317);
or U14760 (N_14760,N_13674,N_13617);
xnor U14761 (N_14761,N_13799,N_13111);
or U14762 (N_14762,N_13948,N_13888);
or U14763 (N_14763,N_13188,N_13507);
nand U14764 (N_14764,N_13960,N_13848);
and U14765 (N_14765,N_13446,N_13411);
or U14766 (N_14766,N_13797,N_13978);
and U14767 (N_14767,N_13809,N_13710);
nor U14768 (N_14768,N_13564,N_13613);
and U14769 (N_14769,N_13119,N_13548);
nand U14770 (N_14770,N_13655,N_13490);
xnor U14771 (N_14771,N_13695,N_13410);
nand U14772 (N_14772,N_13462,N_13432);
or U14773 (N_14773,N_13486,N_13192);
and U14774 (N_14774,N_13610,N_13494);
nor U14775 (N_14775,N_13377,N_13682);
xor U14776 (N_14776,N_13788,N_13512);
nor U14777 (N_14777,N_13767,N_13014);
and U14778 (N_14778,N_13292,N_13440);
nor U14779 (N_14779,N_13075,N_13143);
or U14780 (N_14780,N_13804,N_13558);
xor U14781 (N_14781,N_13925,N_13919);
xnor U14782 (N_14782,N_13330,N_13244);
and U14783 (N_14783,N_13575,N_13980);
xor U14784 (N_14784,N_13569,N_13667);
nand U14785 (N_14785,N_13789,N_13433);
nand U14786 (N_14786,N_13537,N_13716);
and U14787 (N_14787,N_13236,N_13118);
nand U14788 (N_14788,N_13714,N_13219);
nand U14789 (N_14789,N_13152,N_13323);
and U14790 (N_14790,N_13278,N_13812);
xnor U14791 (N_14791,N_13240,N_13479);
and U14792 (N_14792,N_13600,N_13714);
xnor U14793 (N_14793,N_13324,N_13089);
xnor U14794 (N_14794,N_13302,N_13866);
nand U14795 (N_14795,N_13987,N_13415);
and U14796 (N_14796,N_13655,N_13590);
or U14797 (N_14797,N_13962,N_13226);
or U14798 (N_14798,N_13965,N_13763);
and U14799 (N_14799,N_13897,N_13355);
or U14800 (N_14800,N_13373,N_13512);
nor U14801 (N_14801,N_13401,N_13751);
and U14802 (N_14802,N_13544,N_13818);
nand U14803 (N_14803,N_13286,N_13000);
xnor U14804 (N_14804,N_13366,N_13915);
nor U14805 (N_14805,N_13670,N_13201);
and U14806 (N_14806,N_13226,N_13197);
nor U14807 (N_14807,N_13766,N_13349);
nand U14808 (N_14808,N_13651,N_13607);
xor U14809 (N_14809,N_13434,N_13553);
xnor U14810 (N_14810,N_13968,N_13729);
or U14811 (N_14811,N_13765,N_13837);
nor U14812 (N_14812,N_13887,N_13045);
nor U14813 (N_14813,N_13055,N_13784);
nor U14814 (N_14814,N_13808,N_13513);
nand U14815 (N_14815,N_13805,N_13550);
xor U14816 (N_14816,N_13634,N_13275);
xor U14817 (N_14817,N_13088,N_13470);
xnor U14818 (N_14818,N_13593,N_13604);
or U14819 (N_14819,N_13453,N_13313);
nand U14820 (N_14820,N_13802,N_13587);
and U14821 (N_14821,N_13322,N_13391);
nand U14822 (N_14822,N_13074,N_13417);
xnor U14823 (N_14823,N_13021,N_13187);
nor U14824 (N_14824,N_13499,N_13067);
or U14825 (N_14825,N_13565,N_13130);
or U14826 (N_14826,N_13656,N_13320);
nor U14827 (N_14827,N_13906,N_13242);
or U14828 (N_14828,N_13574,N_13092);
and U14829 (N_14829,N_13099,N_13074);
nor U14830 (N_14830,N_13268,N_13605);
nand U14831 (N_14831,N_13635,N_13728);
xnor U14832 (N_14832,N_13838,N_13421);
nand U14833 (N_14833,N_13183,N_13044);
or U14834 (N_14834,N_13771,N_13084);
or U14835 (N_14835,N_13886,N_13191);
xnor U14836 (N_14836,N_13953,N_13859);
xnor U14837 (N_14837,N_13494,N_13031);
xor U14838 (N_14838,N_13542,N_13449);
or U14839 (N_14839,N_13967,N_13121);
xor U14840 (N_14840,N_13560,N_13658);
nand U14841 (N_14841,N_13811,N_13066);
nor U14842 (N_14842,N_13301,N_13948);
nand U14843 (N_14843,N_13271,N_13354);
nor U14844 (N_14844,N_13503,N_13259);
xor U14845 (N_14845,N_13292,N_13616);
and U14846 (N_14846,N_13187,N_13226);
nand U14847 (N_14847,N_13534,N_13925);
and U14848 (N_14848,N_13624,N_13344);
or U14849 (N_14849,N_13210,N_13244);
and U14850 (N_14850,N_13335,N_13654);
nor U14851 (N_14851,N_13254,N_13226);
nor U14852 (N_14852,N_13317,N_13877);
and U14853 (N_14853,N_13175,N_13579);
xor U14854 (N_14854,N_13052,N_13258);
nor U14855 (N_14855,N_13019,N_13825);
nand U14856 (N_14856,N_13349,N_13560);
xnor U14857 (N_14857,N_13364,N_13960);
and U14858 (N_14858,N_13834,N_13730);
nand U14859 (N_14859,N_13236,N_13318);
or U14860 (N_14860,N_13097,N_13385);
nor U14861 (N_14861,N_13756,N_13813);
nor U14862 (N_14862,N_13064,N_13228);
nor U14863 (N_14863,N_13188,N_13664);
and U14864 (N_14864,N_13495,N_13404);
nand U14865 (N_14865,N_13180,N_13473);
nor U14866 (N_14866,N_13588,N_13563);
nor U14867 (N_14867,N_13685,N_13639);
xnor U14868 (N_14868,N_13967,N_13978);
and U14869 (N_14869,N_13956,N_13081);
or U14870 (N_14870,N_13155,N_13593);
and U14871 (N_14871,N_13442,N_13252);
nand U14872 (N_14872,N_13603,N_13482);
xnor U14873 (N_14873,N_13243,N_13209);
nand U14874 (N_14874,N_13992,N_13327);
and U14875 (N_14875,N_13319,N_13259);
or U14876 (N_14876,N_13528,N_13542);
nor U14877 (N_14877,N_13055,N_13897);
nor U14878 (N_14878,N_13663,N_13402);
and U14879 (N_14879,N_13080,N_13072);
and U14880 (N_14880,N_13569,N_13811);
and U14881 (N_14881,N_13811,N_13517);
or U14882 (N_14882,N_13677,N_13520);
nor U14883 (N_14883,N_13324,N_13536);
nand U14884 (N_14884,N_13417,N_13837);
and U14885 (N_14885,N_13808,N_13524);
or U14886 (N_14886,N_13864,N_13765);
nand U14887 (N_14887,N_13912,N_13652);
nor U14888 (N_14888,N_13315,N_13260);
and U14889 (N_14889,N_13769,N_13733);
xor U14890 (N_14890,N_13319,N_13626);
nand U14891 (N_14891,N_13128,N_13484);
xnor U14892 (N_14892,N_13045,N_13376);
xnor U14893 (N_14893,N_13994,N_13887);
and U14894 (N_14894,N_13028,N_13914);
xnor U14895 (N_14895,N_13280,N_13740);
nand U14896 (N_14896,N_13295,N_13054);
nor U14897 (N_14897,N_13384,N_13976);
xor U14898 (N_14898,N_13488,N_13791);
or U14899 (N_14899,N_13566,N_13798);
nor U14900 (N_14900,N_13613,N_13269);
xor U14901 (N_14901,N_13636,N_13449);
xor U14902 (N_14902,N_13943,N_13739);
nor U14903 (N_14903,N_13119,N_13713);
or U14904 (N_14904,N_13889,N_13327);
and U14905 (N_14905,N_13544,N_13205);
xnor U14906 (N_14906,N_13705,N_13129);
or U14907 (N_14907,N_13625,N_13264);
nand U14908 (N_14908,N_13839,N_13071);
and U14909 (N_14909,N_13364,N_13828);
xnor U14910 (N_14910,N_13284,N_13267);
xnor U14911 (N_14911,N_13585,N_13057);
or U14912 (N_14912,N_13431,N_13714);
nand U14913 (N_14913,N_13770,N_13509);
nor U14914 (N_14914,N_13985,N_13938);
or U14915 (N_14915,N_13380,N_13086);
or U14916 (N_14916,N_13237,N_13505);
xor U14917 (N_14917,N_13364,N_13930);
nor U14918 (N_14918,N_13661,N_13867);
or U14919 (N_14919,N_13322,N_13932);
nand U14920 (N_14920,N_13276,N_13299);
or U14921 (N_14921,N_13043,N_13056);
or U14922 (N_14922,N_13689,N_13425);
nor U14923 (N_14923,N_13806,N_13734);
xor U14924 (N_14924,N_13744,N_13591);
and U14925 (N_14925,N_13686,N_13472);
or U14926 (N_14926,N_13722,N_13707);
or U14927 (N_14927,N_13097,N_13883);
or U14928 (N_14928,N_13996,N_13160);
or U14929 (N_14929,N_13266,N_13575);
xor U14930 (N_14930,N_13966,N_13236);
nor U14931 (N_14931,N_13339,N_13586);
nand U14932 (N_14932,N_13531,N_13724);
or U14933 (N_14933,N_13341,N_13412);
or U14934 (N_14934,N_13085,N_13638);
nand U14935 (N_14935,N_13093,N_13867);
nand U14936 (N_14936,N_13592,N_13955);
or U14937 (N_14937,N_13546,N_13166);
nor U14938 (N_14938,N_13332,N_13969);
and U14939 (N_14939,N_13074,N_13968);
nand U14940 (N_14940,N_13638,N_13569);
or U14941 (N_14941,N_13049,N_13347);
xor U14942 (N_14942,N_13520,N_13903);
nor U14943 (N_14943,N_13620,N_13426);
xor U14944 (N_14944,N_13492,N_13400);
nand U14945 (N_14945,N_13859,N_13261);
or U14946 (N_14946,N_13977,N_13689);
and U14947 (N_14947,N_13179,N_13584);
or U14948 (N_14948,N_13487,N_13164);
and U14949 (N_14949,N_13561,N_13519);
or U14950 (N_14950,N_13545,N_13825);
or U14951 (N_14951,N_13567,N_13697);
xnor U14952 (N_14952,N_13709,N_13932);
nand U14953 (N_14953,N_13714,N_13294);
or U14954 (N_14954,N_13524,N_13010);
and U14955 (N_14955,N_13635,N_13485);
xnor U14956 (N_14956,N_13784,N_13800);
xnor U14957 (N_14957,N_13134,N_13118);
or U14958 (N_14958,N_13294,N_13434);
or U14959 (N_14959,N_13338,N_13835);
xnor U14960 (N_14960,N_13286,N_13277);
and U14961 (N_14961,N_13922,N_13964);
or U14962 (N_14962,N_13917,N_13122);
and U14963 (N_14963,N_13117,N_13615);
or U14964 (N_14964,N_13412,N_13334);
and U14965 (N_14965,N_13471,N_13878);
or U14966 (N_14966,N_13064,N_13148);
xnor U14967 (N_14967,N_13904,N_13010);
nor U14968 (N_14968,N_13380,N_13739);
or U14969 (N_14969,N_13456,N_13900);
nor U14970 (N_14970,N_13621,N_13076);
nor U14971 (N_14971,N_13916,N_13792);
nor U14972 (N_14972,N_13663,N_13744);
or U14973 (N_14973,N_13055,N_13752);
or U14974 (N_14974,N_13088,N_13975);
nor U14975 (N_14975,N_13624,N_13967);
or U14976 (N_14976,N_13171,N_13235);
xnor U14977 (N_14977,N_13525,N_13057);
or U14978 (N_14978,N_13123,N_13738);
and U14979 (N_14979,N_13347,N_13884);
and U14980 (N_14980,N_13500,N_13097);
and U14981 (N_14981,N_13636,N_13493);
or U14982 (N_14982,N_13615,N_13703);
nand U14983 (N_14983,N_13840,N_13390);
and U14984 (N_14984,N_13940,N_13116);
and U14985 (N_14985,N_13260,N_13719);
and U14986 (N_14986,N_13702,N_13816);
nand U14987 (N_14987,N_13813,N_13880);
nor U14988 (N_14988,N_13488,N_13406);
and U14989 (N_14989,N_13080,N_13679);
xor U14990 (N_14990,N_13321,N_13866);
nand U14991 (N_14991,N_13655,N_13450);
nand U14992 (N_14992,N_13863,N_13239);
nand U14993 (N_14993,N_13939,N_13088);
xor U14994 (N_14994,N_13918,N_13773);
and U14995 (N_14995,N_13613,N_13741);
or U14996 (N_14996,N_13365,N_13436);
and U14997 (N_14997,N_13681,N_13579);
nor U14998 (N_14998,N_13613,N_13981);
xnor U14999 (N_14999,N_13949,N_13960);
and U15000 (N_15000,N_14063,N_14817);
xor U15001 (N_15001,N_14225,N_14428);
or U15002 (N_15002,N_14681,N_14667);
xor U15003 (N_15003,N_14289,N_14677);
or U15004 (N_15004,N_14334,N_14566);
and U15005 (N_15005,N_14854,N_14673);
nand U15006 (N_15006,N_14570,N_14174);
nor U15007 (N_15007,N_14018,N_14723);
nor U15008 (N_15008,N_14203,N_14163);
nand U15009 (N_15009,N_14499,N_14037);
or U15010 (N_15010,N_14722,N_14030);
nor U15011 (N_15011,N_14493,N_14537);
xnor U15012 (N_15012,N_14699,N_14130);
and U15013 (N_15013,N_14865,N_14369);
xnor U15014 (N_15014,N_14015,N_14983);
nand U15015 (N_15015,N_14489,N_14841);
nor U15016 (N_15016,N_14919,N_14059);
nor U15017 (N_15017,N_14338,N_14964);
and U15018 (N_15018,N_14974,N_14832);
and U15019 (N_15019,N_14367,N_14294);
and U15020 (N_15020,N_14523,N_14134);
and U15021 (N_15021,N_14265,N_14813);
and U15022 (N_15022,N_14268,N_14549);
nor U15023 (N_15023,N_14179,N_14125);
nor U15024 (N_15024,N_14404,N_14229);
nand U15025 (N_15025,N_14167,N_14575);
nor U15026 (N_15026,N_14906,N_14024);
nor U15027 (N_15027,N_14871,N_14506);
xnor U15028 (N_15028,N_14756,N_14312);
nor U15029 (N_15029,N_14823,N_14718);
nor U15030 (N_15030,N_14736,N_14226);
and U15031 (N_15031,N_14313,N_14425);
and U15032 (N_15032,N_14810,N_14465);
and U15033 (N_15033,N_14302,N_14033);
xnor U15034 (N_15034,N_14942,N_14686);
xor U15035 (N_15035,N_14494,N_14145);
nand U15036 (N_15036,N_14066,N_14941);
nor U15037 (N_15037,N_14212,N_14878);
xnor U15038 (N_15038,N_14251,N_14990);
and U15039 (N_15039,N_14855,N_14335);
and U15040 (N_15040,N_14726,N_14547);
xor U15041 (N_15041,N_14784,N_14044);
nand U15042 (N_15042,N_14808,N_14288);
or U15043 (N_15043,N_14508,N_14740);
or U15044 (N_15044,N_14580,N_14440);
nand U15045 (N_15045,N_14462,N_14490);
and U15046 (N_15046,N_14514,N_14504);
nor U15047 (N_15047,N_14303,N_14096);
xnor U15048 (N_15048,N_14023,N_14086);
xnor U15049 (N_15049,N_14257,N_14640);
nand U15050 (N_15050,N_14856,N_14183);
and U15051 (N_15051,N_14616,N_14770);
nand U15052 (N_15052,N_14707,N_14912);
or U15053 (N_15053,N_14531,N_14910);
xnor U15054 (N_15054,N_14131,N_14778);
xor U15055 (N_15055,N_14725,N_14399);
or U15056 (N_15056,N_14711,N_14219);
nor U15057 (N_15057,N_14204,N_14483);
or U15058 (N_15058,N_14842,N_14947);
xor U15059 (N_15059,N_14684,N_14755);
xnor U15060 (N_15060,N_14004,N_14469);
nand U15061 (N_15061,N_14792,N_14058);
xnor U15062 (N_15062,N_14486,N_14546);
or U15063 (N_15063,N_14074,N_14510);
or U15064 (N_15064,N_14576,N_14780);
or U15065 (N_15065,N_14588,N_14704);
or U15066 (N_15066,N_14263,N_14152);
or U15067 (N_15067,N_14785,N_14326);
nor U15068 (N_15068,N_14835,N_14993);
xnor U15069 (N_15069,N_14497,N_14168);
nor U15070 (N_15070,N_14047,N_14700);
nor U15071 (N_15071,N_14060,N_14877);
and U15072 (N_15072,N_14897,N_14655);
nand U15073 (N_15073,N_14414,N_14337);
xnor U15074 (N_15074,N_14963,N_14986);
xor U15075 (N_15075,N_14881,N_14850);
xor U15076 (N_15076,N_14473,N_14480);
and U15077 (N_15077,N_14559,N_14091);
xor U15078 (N_15078,N_14991,N_14773);
and U15079 (N_15079,N_14371,N_14109);
and U15080 (N_15080,N_14861,N_14393);
or U15081 (N_15081,N_14614,N_14811);
xnor U15082 (N_15082,N_14485,N_14396);
nor U15083 (N_15083,N_14360,N_14935);
xnor U15084 (N_15084,N_14847,N_14264);
xnor U15085 (N_15085,N_14410,N_14612);
xor U15086 (N_15086,N_14278,N_14413);
and U15087 (N_15087,N_14498,N_14636);
xor U15088 (N_15088,N_14409,N_14100);
and U15089 (N_15089,N_14142,N_14228);
or U15090 (N_15090,N_14971,N_14162);
nor U15091 (N_15091,N_14247,N_14594);
xnor U15092 (N_15092,N_14237,N_14451);
and U15093 (N_15093,N_14597,N_14643);
or U15094 (N_15094,N_14442,N_14888);
nand U15095 (N_15095,N_14260,N_14821);
and U15096 (N_15096,N_14186,N_14794);
nand U15097 (N_15097,N_14793,N_14014);
nor U15098 (N_15098,N_14296,N_14077);
nand U15099 (N_15099,N_14149,N_14022);
nand U15100 (N_15100,N_14800,N_14574);
nand U15101 (N_15101,N_14582,N_14513);
nor U15102 (N_15102,N_14315,N_14977);
xnor U15103 (N_15103,N_14545,N_14875);
or U15104 (N_15104,N_14757,N_14447);
nor U15105 (N_15105,N_14457,N_14620);
or U15106 (N_15106,N_14759,N_14764);
or U15107 (N_15107,N_14600,N_14089);
nand U15108 (N_15108,N_14628,N_14309);
or U15109 (N_15109,N_14439,N_14158);
or U15110 (N_15110,N_14114,N_14899);
or U15111 (N_15111,N_14141,N_14467);
xor U15112 (N_15112,N_14061,N_14266);
or U15113 (N_15113,N_14662,N_14631);
xor U15114 (N_15114,N_14085,N_14807);
nand U15115 (N_15115,N_14836,N_14040);
nor U15116 (N_15116,N_14767,N_14311);
nor U15117 (N_15117,N_14664,N_14689);
and U15118 (N_15118,N_14528,N_14925);
xor U15119 (N_15119,N_14761,N_14511);
and U15120 (N_15120,N_14530,N_14132);
nor U15121 (N_15121,N_14564,N_14048);
nor U15122 (N_15122,N_14978,N_14332);
or U15123 (N_15123,N_14739,N_14779);
nand U15124 (N_15124,N_14996,N_14441);
xnor U15125 (N_15125,N_14950,N_14992);
xor U15126 (N_15126,N_14316,N_14801);
or U15127 (N_15127,N_14960,N_14953);
nor U15128 (N_15128,N_14437,N_14999);
and U15129 (N_15129,N_14384,N_14862);
nor U15130 (N_15130,N_14049,N_14284);
nand U15131 (N_15131,N_14064,N_14633);
xor U15132 (N_15132,N_14035,N_14571);
and U15133 (N_15133,N_14324,N_14635);
nand U15134 (N_15134,N_14774,N_14129);
or U15135 (N_15135,N_14914,N_14894);
nor U15136 (N_15136,N_14233,N_14694);
and U15137 (N_15137,N_14293,N_14328);
nor U15138 (N_15138,N_14201,N_14540);
and U15139 (N_15139,N_14395,N_14533);
or U15140 (N_15140,N_14331,N_14080);
nand U15141 (N_15141,N_14325,N_14011);
or U15142 (N_15142,N_14522,N_14177);
nor U15143 (N_15143,N_14563,N_14913);
nand U15144 (N_15144,N_14814,N_14777);
or U15145 (N_15145,N_14353,N_14206);
xor U15146 (N_15146,N_14949,N_14221);
nand U15147 (N_15147,N_14669,N_14834);
nand U15148 (N_15148,N_14924,N_14702);
nand U15149 (N_15149,N_14269,N_14660);
or U15150 (N_15150,N_14381,N_14067);
and U15151 (N_15151,N_14378,N_14933);
nor U15152 (N_15152,N_14363,N_14138);
or U15153 (N_15153,N_14173,N_14867);
and U15154 (N_15154,N_14944,N_14827);
and U15155 (N_15155,N_14954,N_14195);
and U15156 (N_15156,N_14502,N_14976);
nor U15157 (N_15157,N_14215,N_14329);
and U15158 (N_15158,N_14534,N_14587);
and U15159 (N_15159,N_14280,N_14029);
xor U15160 (N_15160,N_14223,N_14333);
or U15161 (N_15161,N_14122,N_14435);
xnor U15162 (N_15162,N_14728,N_14691);
or U15163 (N_15163,N_14320,N_14405);
and U15164 (N_15164,N_14420,N_14246);
xor U15165 (N_15165,N_14830,N_14401);
nor U15166 (N_15166,N_14422,N_14354);
nand U15167 (N_15167,N_14751,N_14426);
xnor U15168 (N_15168,N_14359,N_14261);
or U15169 (N_15169,N_14290,N_14883);
or U15170 (N_15170,N_14147,N_14690);
xor U15171 (N_15171,N_14683,N_14368);
nand U15172 (N_15172,N_14292,N_14961);
nand U15173 (N_15173,N_14222,N_14281);
xor U15174 (N_15174,N_14169,N_14904);
nand U15175 (N_15175,N_14985,N_14989);
and U15176 (N_15176,N_14937,N_14624);
or U15177 (N_15177,N_14357,N_14565);
and U15178 (N_15178,N_14110,N_14535);
nor U15179 (N_15179,N_14042,N_14666);
nand U15180 (N_15180,N_14885,N_14271);
or U15181 (N_15181,N_14592,N_14972);
xnor U15182 (N_15182,N_14833,N_14382);
xnor U15183 (N_15183,N_14584,N_14407);
xnor U15184 (N_15184,N_14788,N_14460);
and U15185 (N_15185,N_14803,N_14596);
nor U15186 (N_15186,N_14967,N_14027);
or U15187 (N_15187,N_14816,N_14242);
xor U15188 (N_15188,N_14458,N_14424);
nor U15189 (N_15189,N_14958,N_14340);
nand U15190 (N_15190,N_14717,N_14892);
nor U15191 (N_15191,N_14589,N_14495);
and U15192 (N_15192,N_14306,N_14386);
and U15193 (N_15193,N_14345,N_14065);
nor U15194 (N_15194,N_14644,N_14105);
nor U15195 (N_15195,N_14283,N_14321);
nor U15196 (N_15196,N_14491,N_14270);
and U15197 (N_15197,N_14455,N_14527);
or U15198 (N_15198,N_14391,N_14276);
nor U15199 (N_15199,N_14599,N_14078);
nor U15200 (N_15200,N_14202,N_14026);
and U15201 (N_15201,N_14446,N_14581);
nor U15202 (N_15202,N_14475,N_14039);
and U15203 (N_15203,N_14092,N_14081);
nand U15204 (N_15204,N_14626,N_14632);
nor U15205 (N_15205,N_14595,N_14846);
or U15206 (N_15206,N_14744,N_14118);
or U15207 (N_15207,N_14826,N_14239);
xnor U15208 (N_15208,N_14532,N_14705);
nand U15209 (N_15209,N_14526,N_14747);
xor U15210 (N_15210,N_14638,N_14782);
nand U15211 (N_15211,N_14796,N_14103);
nand U15212 (N_15212,N_14610,N_14444);
nand U15213 (N_15213,N_14402,N_14973);
and U15214 (N_15214,N_14873,N_14697);
and U15215 (N_15215,N_14210,N_14795);
xnor U15216 (N_15216,N_14998,N_14661);
nor U15217 (N_15217,N_14901,N_14071);
nor U15218 (N_15218,N_14938,N_14746);
nor U15219 (N_15219,N_14358,N_14880);
nand U15220 (N_15220,N_14959,N_14503);
nand U15221 (N_15221,N_14791,N_14005);
nand U15222 (N_15222,N_14300,N_14126);
or U15223 (N_15223,N_14012,N_14923);
and U15224 (N_15224,N_14706,N_14038);
xor U15225 (N_15225,N_14182,N_14646);
nand U15226 (N_15226,N_14196,N_14211);
or U15227 (N_15227,N_14872,N_14905);
nor U15228 (N_15228,N_14552,N_14472);
and U15229 (N_15229,N_14561,N_14124);
nor U15230 (N_15230,N_14094,N_14139);
and U15231 (N_15231,N_14488,N_14088);
or U15232 (N_15232,N_14554,N_14648);
and U15233 (N_15233,N_14945,N_14322);
nand U15234 (N_15234,N_14448,N_14682);
nand U15235 (N_15235,N_14715,N_14275);
xnor U15236 (N_15236,N_14106,N_14693);
or U15237 (N_15237,N_14886,N_14829);
and U15238 (N_15238,N_14539,N_14956);
or U15239 (N_15239,N_14095,N_14299);
and U15240 (N_15240,N_14887,N_14376);
nand U15241 (N_15241,N_14607,N_14234);
nor U15242 (N_15242,N_14374,N_14957);
and U15243 (N_15243,N_14768,N_14282);
xor U15244 (N_15244,N_14084,N_14613);
nor U15245 (N_15245,N_14674,N_14820);
nor U15246 (N_15246,N_14752,N_14787);
or U15247 (N_15247,N_14603,N_14590);
nor U15248 (N_15248,N_14433,N_14562);
nor U15249 (N_15249,N_14216,N_14262);
nand U15250 (N_15250,N_14193,N_14789);
and U15251 (N_15251,N_14364,N_14013);
or U15252 (N_15252,N_14805,N_14192);
and U15253 (N_15253,N_14454,N_14450);
nand U15254 (N_15254,N_14979,N_14250);
and U15255 (N_15255,N_14623,N_14733);
and U15256 (N_15256,N_14043,N_14327);
nor U15257 (N_15257,N_14572,N_14471);
nand U15258 (N_15258,N_14180,N_14891);
xor U15259 (N_15259,N_14474,N_14776);
nor U15260 (N_15260,N_14825,N_14484);
xnor U15261 (N_15261,N_14670,N_14150);
xnor U15262 (N_15262,N_14161,N_14255);
or U15263 (N_15263,N_14054,N_14918);
nor U15264 (N_15264,N_14224,N_14797);
or U15265 (N_15265,N_14927,N_14555);
xnor U15266 (N_15266,N_14235,N_14273);
nand U15267 (N_15267,N_14199,N_14343);
or U15268 (N_15268,N_14968,N_14931);
and U15269 (N_15269,N_14082,N_14737);
nand U15270 (N_15270,N_14955,N_14758);
or U15271 (N_15271,N_14893,N_14853);
nand U15272 (N_15272,N_14198,N_14240);
nor U15273 (N_15273,N_14621,N_14241);
xnor U15274 (N_15274,N_14839,N_14112);
or U15275 (N_15275,N_14415,N_14146);
nand U15276 (N_15276,N_14852,N_14618);
and U15277 (N_15277,N_14922,N_14698);
and U15278 (N_15278,N_14160,N_14121);
nand U15279 (N_15279,N_14016,N_14187);
xnor U15280 (N_15280,N_14009,N_14557);
and U15281 (N_15281,N_14649,N_14287);
or U15282 (N_15282,N_14731,N_14297);
xnor U15283 (N_15283,N_14479,N_14890);
xor U15284 (N_15284,N_14107,N_14962);
or U15285 (N_15285,N_14809,N_14041);
or U15286 (N_15286,N_14341,N_14806);
or U15287 (N_15287,N_14858,N_14524);
nand U15288 (N_15288,N_14032,N_14934);
xor U15289 (N_15289,N_14988,N_14220);
xnor U15290 (N_15290,N_14815,N_14857);
nand U15291 (N_15291,N_14243,N_14166);
or U15292 (N_15292,N_14911,N_14099);
and U15293 (N_15293,N_14267,N_14553);
or U15294 (N_15294,N_14431,N_14845);
nand U15295 (N_15295,N_14445,N_14463);
and U15296 (N_15296,N_14020,N_14676);
xor U15297 (N_15297,N_14002,N_14837);
and U15298 (N_15298,N_14679,N_14710);
and U15299 (N_15299,N_14654,N_14743);
xor U15300 (N_15300,N_14144,N_14548);
and U15301 (N_15301,N_14019,N_14487);
and U15302 (N_15302,N_14675,N_14558);
nor U15303 (N_15303,N_14466,N_14969);
nor U15304 (N_15304,N_14790,N_14647);
xor U15305 (N_15305,N_14310,N_14585);
nand U15306 (N_15306,N_14917,N_14951);
nand U15307 (N_15307,N_14766,N_14799);
xor U15308 (N_15308,N_14373,N_14028);
or U15309 (N_15309,N_14007,N_14754);
or U15310 (N_15310,N_14884,N_14671);
nand U15311 (N_15311,N_14197,N_14400);
xnor U15312 (N_15312,N_14056,N_14984);
xnor U15313 (N_15313,N_14076,N_14176);
xnor U15314 (N_15314,N_14509,N_14102);
nand U15315 (N_15315,N_14209,N_14762);
xnor U15316 (N_15316,N_14365,N_14849);
nand U15317 (N_15317,N_14477,N_14939);
nand U15318 (N_15318,N_14380,N_14178);
nand U15319 (N_15319,N_14135,N_14098);
and U15320 (N_15320,N_14323,N_14031);
or U15321 (N_15321,N_14238,N_14025);
or U15322 (N_15322,N_14344,N_14568);
nand U15323 (N_15323,N_14645,N_14516);
nand U15324 (N_15324,N_14070,N_14903);
nand U15325 (N_15325,N_14665,N_14189);
and U15326 (N_15326,N_14943,N_14653);
nor U15327 (N_15327,N_14436,N_14254);
nand U15328 (N_15328,N_14525,N_14231);
xnor U15329 (N_15329,N_14184,N_14148);
xor U15330 (N_15330,N_14119,N_14214);
nor U15331 (N_15331,N_14248,N_14501);
and U15332 (N_15332,N_14538,N_14355);
nor U15333 (N_15333,N_14601,N_14639);
nor U15334 (N_15334,N_14900,N_14657);
xnor U15335 (N_15335,N_14902,N_14512);
and U15336 (N_15336,N_14609,N_14295);
nand U15337 (N_15337,N_14137,N_14108);
nor U15338 (N_15338,N_14518,N_14742);
nor U15339 (N_15339,N_14379,N_14567);
nand U15340 (N_15340,N_14748,N_14430);
xor U15341 (N_15341,N_14980,N_14113);
nand U15342 (N_15342,N_14185,N_14034);
and U15343 (N_15343,N_14529,N_14920);
nand U15344 (N_15344,N_14330,N_14763);
xor U15345 (N_15345,N_14087,N_14213);
xor U15346 (N_15346,N_14370,N_14408);
nand U15347 (N_15347,N_14046,N_14274);
or U15348 (N_15348,N_14619,N_14432);
and U15349 (N_15349,N_14895,N_14928);
nor U15350 (N_15350,N_14304,N_14760);
xor U15351 (N_15351,N_14236,N_14127);
and U15352 (N_15352,N_14286,N_14712);
nor U15353 (N_15353,N_14277,N_14175);
and U15354 (N_15354,N_14285,N_14492);
and U15355 (N_15355,N_14542,N_14200);
nand U15356 (N_15356,N_14840,N_14190);
and U15357 (N_15357,N_14519,N_14716);
and U15358 (N_15358,N_14366,N_14882);
xor U15359 (N_15359,N_14641,N_14642);
and U15360 (N_15360,N_14423,N_14083);
and U15361 (N_15361,N_14753,N_14615);
nand U15362 (N_15362,N_14703,N_14772);
or U15363 (N_15363,N_14948,N_14403);
and U15364 (N_15364,N_14769,N_14627);
xnor U15365 (N_15365,N_14520,N_14157);
nor U15366 (N_15366,N_14385,N_14397);
and U15367 (N_15367,N_14732,N_14181);
xnor U15368 (N_15368,N_14605,N_14936);
nand U15369 (N_15369,N_14630,N_14003);
or U15370 (N_15370,N_14573,N_14001);
and U15371 (N_15371,N_14940,N_14678);
or U15372 (N_15372,N_14656,N_14586);
or U15373 (N_15373,N_14713,N_14604);
nand U15374 (N_15374,N_14258,N_14804);
nor U15375 (N_15375,N_14298,N_14045);
or U15376 (N_15376,N_14449,N_14577);
xor U15377 (N_15377,N_14392,N_14377);
and U15378 (N_15378,N_14541,N_14591);
nor U15379 (N_15379,N_14232,N_14230);
nor U15380 (N_15380,N_14123,N_14155);
or U15381 (N_15381,N_14342,N_14593);
xor U15382 (N_15382,N_14916,N_14482);
xor U15383 (N_15383,N_14500,N_14383);
and U15384 (N_15384,N_14637,N_14771);
nand U15385 (N_15385,N_14543,N_14116);
nand U15386 (N_15386,N_14120,N_14907);
and U15387 (N_15387,N_14569,N_14617);
or U15388 (N_15388,N_14349,N_14348);
xor U15389 (N_15389,N_14658,N_14418);
or U15390 (N_15390,N_14997,N_14687);
xor U15391 (N_15391,N_14932,N_14843);
nand U15392 (N_15392,N_14714,N_14244);
and U15393 (N_15393,N_14352,N_14438);
and U15394 (N_15394,N_14140,N_14217);
or U15395 (N_15395,N_14339,N_14093);
xnor U15396 (N_15396,N_14164,N_14889);
and U15397 (N_15397,N_14090,N_14291);
nor U15398 (N_15398,N_14079,N_14165);
or U15399 (N_15399,N_14798,N_14578);
xnor U15400 (N_15400,N_14870,N_14000);
or U15401 (N_15401,N_14069,N_14136);
or U15402 (N_15402,N_14611,N_14053);
xor U15403 (N_15403,N_14476,N_14926);
nor U15404 (N_15404,N_14468,N_14478);
nor U15405 (N_15405,N_14429,N_14253);
nor U15406 (N_15406,N_14844,N_14055);
xnor U15407 (N_15407,N_14864,N_14218);
nand U15408 (N_15408,N_14470,N_14659);
xnor U15409 (N_15409,N_14859,N_14551);
nor U15410 (N_15410,N_14245,N_14249);
xor U15411 (N_15411,N_14411,N_14724);
or U15412 (N_15412,N_14072,N_14781);
nor U15413 (N_15413,N_14598,N_14464);
nor U15414 (N_15414,N_14427,N_14734);
nor U15415 (N_15415,N_14879,N_14629);
or U15416 (N_15416,N_14831,N_14663);
nor U15417 (N_15417,N_14461,N_14719);
nor U15418 (N_15418,N_14898,N_14372);
xnor U15419 (N_15419,N_14314,N_14317);
nor U15420 (N_15420,N_14159,N_14556);
nand U15421 (N_15421,N_14434,N_14394);
nor U15422 (N_15422,N_14730,N_14579);
and U15423 (N_15423,N_14036,N_14692);
nand U15424 (N_15424,N_14838,N_14672);
xnor U15425 (N_15425,N_14406,N_14075);
nand U15426 (N_15426,N_14207,N_14205);
nand U15427 (N_15427,N_14720,N_14729);
and U15428 (N_15428,N_14822,N_14507);
nor U15429 (N_15429,N_14668,N_14921);
nor U15430 (N_15430,N_14868,N_14874);
xor U15431 (N_15431,N_14010,N_14481);
nand U15432 (N_15432,N_14975,N_14008);
nor U15433 (N_15433,N_14828,N_14459);
and U15434 (N_15434,N_14443,N_14505);
nor U15435 (N_15435,N_14583,N_14802);
or U15436 (N_15436,N_14930,N_14863);
nor U15437 (N_15437,N_14111,N_14104);
xnor U15438 (N_15438,N_14848,N_14021);
xor U15439 (N_15439,N_14361,N_14709);
nor U15440 (N_15440,N_14272,N_14909);
xnor U15441 (N_15441,N_14966,N_14151);
and U15442 (N_15442,N_14695,N_14786);
nand U15443 (N_15443,N_14970,N_14143);
nor U15444 (N_15444,N_14908,N_14735);
nor U15445 (N_15445,N_14651,N_14521);
or U15446 (N_15446,N_14896,N_14252);
and U15447 (N_15447,N_14952,N_14319);
and U15448 (N_15448,N_14398,N_14696);
and U15449 (N_15449,N_14775,N_14188);
nand U15450 (N_15450,N_14208,N_14456);
or U15451 (N_15451,N_14750,N_14765);
and U15452 (N_15452,N_14006,N_14634);
nor U15453 (N_15453,N_14279,N_14387);
nand U15454 (N_15454,N_14101,N_14305);
or U15455 (N_15455,N_14417,N_14602);
nand U15456 (N_15456,N_14708,N_14362);
or U15457 (N_15457,N_14741,N_14133);
or U15458 (N_15458,N_14680,N_14171);
and U15459 (N_15459,N_14301,N_14606);
or U15460 (N_15460,N_14356,N_14388);
nand U15461 (N_15461,N_14307,N_14981);
nor U15462 (N_15462,N_14625,N_14117);
and U15463 (N_15463,N_14749,N_14869);
or U15464 (N_15464,N_14191,N_14550);
xor U15465 (N_15465,N_14259,N_14824);
and U15466 (N_15466,N_14153,N_14866);
xnor U15467 (N_15467,N_14375,N_14812);
nor U15468 (N_15468,N_14051,N_14544);
and U15469 (N_15469,N_14688,N_14536);
xnor U15470 (N_15470,N_14622,N_14738);
or U15471 (N_15471,N_14745,N_14496);
nor U15472 (N_15472,N_14721,N_14982);
and U15473 (N_15473,N_14389,N_14073);
nor U15474 (N_15474,N_14347,N_14929);
nor U15475 (N_15475,N_14128,N_14650);
and U15476 (N_15476,N_14987,N_14308);
xnor U15477 (N_15477,N_14685,N_14156);
and U15478 (N_15478,N_14346,N_14115);
and U15479 (N_15479,N_14412,N_14517);
nor U15480 (N_15480,N_14818,N_14860);
xnor U15481 (N_15481,N_14727,N_14915);
and U15482 (N_15482,N_14336,N_14416);
xor U15483 (N_15483,N_14256,N_14608);
nor U15484 (N_15484,N_14154,N_14318);
nor U15485 (N_15485,N_14946,N_14351);
or U15486 (N_15486,N_14453,N_14851);
and U15487 (N_15487,N_14194,N_14419);
xor U15488 (N_15488,N_14652,N_14515);
nand U15489 (N_15489,N_14050,N_14052);
nand U15490 (N_15490,N_14819,N_14390);
nand U15491 (N_15491,N_14017,N_14994);
and U15492 (N_15492,N_14068,N_14965);
nand U15493 (N_15493,N_14421,N_14057);
or U15494 (N_15494,N_14995,N_14560);
xnor U15495 (N_15495,N_14170,N_14172);
xor U15496 (N_15496,N_14783,N_14227);
nor U15497 (N_15497,N_14097,N_14876);
nand U15498 (N_15498,N_14062,N_14350);
nand U15499 (N_15499,N_14701,N_14452);
xnor U15500 (N_15500,N_14835,N_14263);
nor U15501 (N_15501,N_14331,N_14556);
xor U15502 (N_15502,N_14176,N_14543);
nand U15503 (N_15503,N_14157,N_14326);
xnor U15504 (N_15504,N_14740,N_14729);
xnor U15505 (N_15505,N_14506,N_14321);
nand U15506 (N_15506,N_14619,N_14021);
or U15507 (N_15507,N_14480,N_14965);
nor U15508 (N_15508,N_14524,N_14364);
and U15509 (N_15509,N_14605,N_14599);
nand U15510 (N_15510,N_14523,N_14962);
nor U15511 (N_15511,N_14871,N_14185);
and U15512 (N_15512,N_14759,N_14424);
nor U15513 (N_15513,N_14562,N_14559);
nor U15514 (N_15514,N_14025,N_14764);
or U15515 (N_15515,N_14139,N_14778);
and U15516 (N_15516,N_14164,N_14089);
nor U15517 (N_15517,N_14065,N_14246);
and U15518 (N_15518,N_14013,N_14508);
nor U15519 (N_15519,N_14973,N_14978);
nor U15520 (N_15520,N_14864,N_14971);
xnor U15521 (N_15521,N_14931,N_14745);
nor U15522 (N_15522,N_14003,N_14492);
and U15523 (N_15523,N_14671,N_14713);
nor U15524 (N_15524,N_14791,N_14242);
nor U15525 (N_15525,N_14529,N_14116);
nor U15526 (N_15526,N_14117,N_14514);
or U15527 (N_15527,N_14139,N_14769);
xor U15528 (N_15528,N_14120,N_14402);
xor U15529 (N_15529,N_14425,N_14448);
xor U15530 (N_15530,N_14187,N_14050);
nand U15531 (N_15531,N_14073,N_14914);
nand U15532 (N_15532,N_14624,N_14568);
nor U15533 (N_15533,N_14824,N_14059);
or U15534 (N_15534,N_14035,N_14140);
xor U15535 (N_15535,N_14831,N_14636);
nand U15536 (N_15536,N_14594,N_14769);
or U15537 (N_15537,N_14533,N_14990);
xnor U15538 (N_15538,N_14758,N_14732);
xor U15539 (N_15539,N_14544,N_14217);
nor U15540 (N_15540,N_14425,N_14526);
or U15541 (N_15541,N_14854,N_14732);
nor U15542 (N_15542,N_14525,N_14779);
or U15543 (N_15543,N_14845,N_14052);
nand U15544 (N_15544,N_14066,N_14210);
and U15545 (N_15545,N_14558,N_14950);
or U15546 (N_15546,N_14428,N_14723);
nor U15547 (N_15547,N_14533,N_14633);
or U15548 (N_15548,N_14148,N_14880);
or U15549 (N_15549,N_14169,N_14264);
xnor U15550 (N_15550,N_14787,N_14591);
nor U15551 (N_15551,N_14282,N_14359);
nor U15552 (N_15552,N_14626,N_14835);
nor U15553 (N_15553,N_14945,N_14271);
nor U15554 (N_15554,N_14022,N_14517);
nand U15555 (N_15555,N_14665,N_14623);
or U15556 (N_15556,N_14712,N_14117);
xor U15557 (N_15557,N_14515,N_14083);
nor U15558 (N_15558,N_14802,N_14000);
nand U15559 (N_15559,N_14948,N_14116);
or U15560 (N_15560,N_14907,N_14013);
or U15561 (N_15561,N_14452,N_14650);
nand U15562 (N_15562,N_14860,N_14833);
and U15563 (N_15563,N_14001,N_14325);
nand U15564 (N_15564,N_14922,N_14963);
nand U15565 (N_15565,N_14124,N_14401);
or U15566 (N_15566,N_14589,N_14017);
and U15567 (N_15567,N_14017,N_14228);
nor U15568 (N_15568,N_14961,N_14383);
nand U15569 (N_15569,N_14167,N_14215);
xnor U15570 (N_15570,N_14368,N_14949);
and U15571 (N_15571,N_14866,N_14701);
nor U15572 (N_15572,N_14277,N_14051);
or U15573 (N_15573,N_14378,N_14806);
or U15574 (N_15574,N_14862,N_14871);
or U15575 (N_15575,N_14420,N_14442);
nand U15576 (N_15576,N_14789,N_14182);
nor U15577 (N_15577,N_14010,N_14702);
nand U15578 (N_15578,N_14931,N_14929);
or U15579 (N_15579,N_14571,N_14022);
nor U15580 (N_15580,N_14676,N_14851);
and U15581 (N_15581,N_14888,N_14355);
nor U15582 (N_15582,N_14638,N_14806);
and U15583 (N_15583,N_14224,N_14677);
and U15584 (N_15584,N_14657,N_14871);
xnor U15585 (N_15585,N_14536,N_14056);
xor U15586 (N_15586,N_14890,N_14711);
xor U15587 (N_15587,N_14420,N_14516);
and U15588 (N_15588,N_14961,N_14441);
or U15589 (N_15589,N_14975,N_14844);
nor U15590 (N_15590,N_14431,N_14944);
xnor U15591 (N_15591,N_14221,N_14441);
or U15592 (N_15592,N_14921,N_14676);
or U15593 (N_15593,N_14810,N_14081);
nor U15594 (N_15594,N_14289,N_14944);
nand U15595 (N_15595,N_14482,N_14819);
and U15596 (N_15596,N_14044,N_14465);
nor U15597 (N_15597,N_14863,N_14492);
and U15598 (N_15598,N_14977,N_14890);
nor U15599 (N_15599,N_14873,N_14990);
or U15600 (N_15600,N_14573,N_14833);
or U15601 (N_15601,N_14159,N_14455);
xor U15602 (N_15602,N_14630,N_14286);
nand U15603 (N_15603,N_14109,N_14470);
or U15604 (N_15604,N_14109,N_14749);
xor U15605 (N_15605,N_14213,N_14957);
nor U15606 (N_15606,N_14177,N_14206);
nand U15607 (N_15607,N_14675,N_14475);
nor U15608 (N_15608,N_14700,N_14582);
and U15609 (N_15609,N_14791,N_14763);
nor U15610 (N_15610,N_14952,N_14941);
and U15611 (N_15611,N_14150,N_14509);
and U15612 (N_15612,N_14448,N_14047);
nor U15613 (N_15613,N_14185,N_14681);
and U15614 (N_15614,N_14027,N_14238);
or U15615 (N_15615,N_14391,N_14393);
xnor U15616 (N_15616,N_14924,N_14331);
nor U15617 (N_15617,N_14065,N_14757);
xor U15618 (N_15618,N_14710,N_14052);
or U15619 (N_15619,N_14384,N_14892);
xnor U15620 (N_15620,N_14981,N_14341);
xnor U15621 (N_15621,N_14445,N_14759);
and U15622 (N_15622,N_14549,N_14542);
nand U15623 (N_15623,N_14974,N_14647);
nor U15624 (N_15624,N_14441,N_14036);
nor U15625 (N_15625,N_14943,N_14356);
nor U15626 (N_15626,N_14838,N_14331);
or U15627 (N_15627,N_14850,N_14637);
nand U15628 (N_15628,N_14030,N_14535);
nor U15629 (N_15629,N_14593,N_14343);
or U15630 (N_15630,N_14225,N_14568);
xnor U15631 (N_15631,N_14952,N_14491);
xor U15632 (N_15632,N_14566,N_14234);
xnor U15633 (N_15633,N_14216,N_14290);
or U15634 (N_15634,N_14215,N_14044);
nor U15635 (N_15635,N_14063,N_14417);
or U15636 (N_15636,N_14516,N_14273);
nor U15637 (N_15637,N_14874,N_14499);
nor U15638 (N_15638,N_14557,N_14466);
xor U15639 (N_15639,N_14691,N_14842);
nor U15640 (N_15640,N_14850,N_14103);
nor U15641 (N_15641,N_14629,N_14714);
and U15642 (N_15642,N_14506,N_14207);
nor U15643 (N_15643,N_14319,N_14499);
and U15644 (N_15644,N_14715,N_14495);
nor U15645 (N_15645,N_14042,N_14690);
xnor U15646 (N_15646,N_14379,N_14092);
or U15647 (N_15647,N_14099,N_14174);
and U15648 (N_15648,N_14884,N_14417);
and U15649 (N_15649,N_14495,N_14660);
xor U15650 (N_15650,N_14764,N_14969);
nand U15651 (N_15651,N_14662,N_14658);
xor U15652 (N_15652,N_14712,N_14423);
xnor U15653 (N_15653,N_14422,N_14399);
and U15654 (N_15654,N_14080,N_14947);
and U15655 (N_15655,N_14368,N_14314);
and U15656 (N_15656,N_14563,N_14934);
nand U15657 (N_15657,N_14911,N_14265);
nand U15658 (N_15658,N_14542,N_14272);
and U15659 (N_15659,N_14246,N_14291);
xor U15660 (N_15660,N_14540,N_14010);
nand U15661 (N_15661,N_14605,N_14300);
and U15662 (N_15662,N_14142,N_14003);
nor U15663 (N_15663,N_14318,N_14162);
and U15664 (N_15664,N_14577,N_14865);
and U15665 (N_15665,N_14061,N_14210);
xnor U15666 (N_15666,N_14046,N_14463);
nand U15667 (N_15667,N_14528,N_14437);
xor U15668 (N_15668,N_14838,N_14425);
or U15669 (N_15669,N_14946,N_14544);
nor U15670 (N_15670,N_14494,N_14390);
xnor U15671 (N_15671,N_14634,N_14825);
xnor U15672 (N_15672,N_14518,N_14570);
or U15673 (N_15673,N_14756,N_14438);
nand U15674 (N_15674,N_14059,N_14315);
and U15675 (N_15675,N_14674,N_14438);
nand U15676 (N_15676,N_14862,N_14783);
nor U15677 (N_15677,N_14242,N_14480);
or U15678 (N_15678,N_14504,N_14231);
nand U15679 (N_15679,N_14038,N_14958);
xor U15680 (N_15680,N_14168,N_14198);
nor U15681 (N_15681,N_14223,N_14511);
nor U15682 (N_15682,N_14587,N_14539);
nand U15683 (N_15683,N_14421,N_14422);
xor U15684 (N_15684,N_14577,N_14221);
or U15685 (N_15685,N_14780,N_14740);
nor U15686 (N_15686,N_14132,N_14117);
nand U15687 (N_15687,N_14744,N_14753);
and U15688 (N_15688,N_14492,N_14233);
and U15689 (N_15689,N_14355,N_14592);
xor U15690 (N_15690,N_14120,N_14129);
xor U15691 (N_15691,N_14568,N_14606);
nand U15692 (N_15692,N_14379,N_14869);
or U15693 (N_15693,N_14425,N_14386);
and U15694 (N_15694,N_14304,N_14347);
nand U15695 (N_15695,N_14979,N_14700);
nor U15696 (N_15696,N_14972,N_14526);
and U15697 (N_15697,N_14290,N_14470);
nand U15698 (N_15698,N_14065,N_14708);
nand U15699 (N_15699,N_14491,N_14211);
nor U15700 (N_15700,N_14573,N_14951);
or U15701 (N_15701,N_14837,N_14701);
nand U15702 (N_15702,N_14193,N_14512);
or U15703 (N_15703,N_14101,N_14287);
nand U15704 (N_15704,N_14523,N_14577);
nor U15705 (N_15705,N_14321,N_14004);
nand U15706 (N_15706,N_14011,N_14197);
nand U15707 (N_15707,N_14989,N_14728);
and U15708 (N_15708,N_14692,N_14287);
or U15709 (N_15709,N_14513,N_14912);
or U15710 (N_15710,N_14940,N_14491);
nand U15711 (N_15711,N_14844,N_14565);
xor U15712 (N_15712,N_14987,N_14667);
nor U15713 (N_15713,N_14060,N_14010);
and U15714 (N_15714,N_14135,N_14651);
or U15715 (N_15715,N_14970,N_14212);
or U15716 (N_15716,N_14411,N_14386);
and U15717 (N_15717,N_14768,N_14186);
nor U15718 (N_15718,N_14511,N_14902);
or U15719 (N_15719,N_14500,N_14812);
nor U15720 (N_15720,N_14804,N_14296);
or U15721 (N_15721,N_14852,N_14080);
nand U15722 (N_15722,N_14700,N_14828);
and U15723 (N_15723,N_14236,N_14256);
or U15724 (N_15724,N_14915,N_14883);
nor U15725 (N_15725,N_14847,N_14645);
xnor U15726 (N_15726,N_14538,N_14918);
nand U15727 (N_15727,N_14701,N_14225);
xnor U15728 (N_15728,N_14544,N_14301);
nand U15729 (N_15729,N_14999,N_14396);
xor U15730 (N_15730,N_14383,N_14384);
and U15731 (N_15731,N_14271,N_14566);
xnor U15732 (N_15732,N_14801,N_14526);
or U15733 (N_15733,N_14887,N_14722);
or U15734 (N_15734,N_14663,N_14428);
nor U15735 (N_15735,N_14675,N_14545);
xor U15736 (N_15736,N_14973,N_14948);
xor U15737 (N_15737,N_14660,N_14626);
or U15738 (N_15738,N_14859,N_14766);
and U15739 (N_15739,N_14152,N_14641);
or U15740 (N_15740,N_14060,N_14384);
or U15741 (N_15741,N_14581,N_14317);
or U15742 (N_15742,N_14627,N_14382);
or U15743 (N_15743,N_14102,N_14959);
nand U15744 (N_15744,N_14526,N_14719);
xor U15745 (N_15745,N_14158,N_14031);
nand U15746 (N_15746,N_14309,N_14831);
nor U15747 (N_15747,N_14975,N_14227);
xnor U15748 (N_15748,N_14734,N_14174);
nand U15749 (N_15749,N_14979,N_14216);
and U15750 (N_15750,N_14825,N_14242);
xor U15751 (N_15751,N_14069,N_14846);
and U15752 (N_15752,N_14856,N_14008);
nor U15753 (N_15753,N_14675,N_14044);
nor U15754 (N_15754,N_14984,N_14244);
nor U15755 (N_15755,N_14697,N_14900);
xnor U15756 (N_15756,N_14030,N_14951);
nor U15757 (N_15757,N_14114,N_14641);
nand U15758 (N_15758,N_14514,N_14758);
and U15759 (N_15759,N_14809,N_14493);
or U15760 (N_15760,N_14221,N_14550);
nor U15761 (N_15761,N_14982,N_14378);
and U15762 (N_15762,N_14648,N_14821);
nand U15763 (N_15763,N_14316,N_14879);
nand U15764 (N_15764,N_14653,N_14985);
nor U15765 (N_15765,N_14753,N_14009);
and U15766 (N_15766,N_14684,N_14603);
nand U15767 (N_15767,N_14047,N_14044);
nand U15768 (N_15768,N_14246,N_14628);
xnor U15769 (N_15769,N_14222,N_14935);
or U15770 (N_15770,N_14129,N_14476);
xor U15771 (N_15771,N_14895,N_14786);
xnor U15772 (N_15772,N_14761,N_14353);
and U15773 (N_15773,N_14654,N_14628);
xnor U15774 (N_15774,N_14915,N_14289);
and U15775 (N_15775,N_14237,N_14236);
or U15776 (N_15776,N_14775,N_14685);
nand U15777 (N_15777,N_14967,N_14656);
xnor U15778 (N_15778,N_14214,N_14353);
xnor U15779 (N_15779,N_14763,N_14913);
xnor U15780 (N_15780,N_14696,N_14419);
nor U15781 (N_15781,N_14654,N_14227);
xnor U15782 (N_15782,N_14715,N_14020);
or U15783 (N_15783,N_14007,N_14353);
nor U15784 (N_15784,N_14328,N_14452);
or U15785 (N_15785,N_14026,N_14906);
nor U15786 (N_15786,N_14188,N_14967);
and U15787 (N_15787,N_14946,N_14120);
nand U15788 (N_15788,N_14043,N_14570);
or U15789 (N_15789,N_14520,N_14656);
xnor U15790 (N_15790,N_14099,N_14860);
nor U15791 (N_15791,N_14188,N_14839);
nand U15792 (N_15792,N_14444,N_14411);
or U15793 (N_15793,N_14861,N_14258);
nor U15794 (N_15794,N_14355,N_14787);
nand U15795 (N_15795,N_14966,N_14157);
and U15796 (N_15796,N_14161,N_14091);
or U15797 (N_15797,N_14977,N_14436);
nand U15798 (N_15798,N_14137,N_14648);
nand U15799 (N_15799,N_14840,N_14272);
nor U15800 (N_15800,N_14679,N_14659);
and U15801 (N_15801,N_14282,N_14426);
nor U15802 (N_15802,N_14190,N_14181);
or U15803 (N_15803,N_14399,N_14050);
nand U15804 (N_15804,N_14440,N_14390);
and U15805 (N_15805,N_14897,N_14336);
nor U15806 (N_15806,N_14384,N_14361);
xnor U15807 (N_15807,N_14815,N_14230);
or U15808 (N_15808,N_14250,N_14875);
nor U15809 (N_15809,N_14784,N_14938);
nor U15810 (N_15810,N_14462,N_14249);
and U15811 (N_15811,N_14876,N_14103);
xor U15812 (N_15812,N_14660,N_14937);
xor U15813 (N_15813,N_14773,N_14855);
and U15814 (N_15814,N_14686,N_14124);
and U15815 (N_15815,N_14715,N_14832);
nand U15816 (N_15816,N_14650,N_14471);
nand U15817 (N_15817,N_14521,N_14745);
xor U15818 (N_15818,N_14484,N_14246);
xnor U15819 (N_15819,N_14766,N_14550);
xnor U15820 (N_15820,N_14818,N_14891);
xnor U15821 (N_15821,N_14004,N_14902);
nor U15822 (N_15822,N_14786,N_14182);
and U15823 (N_15823,N_14358,N_14298);
nor U15824 (N_15824,N_14479,N_14719);
nor U15825 (N_15825,N_14617,N_14242);
or U15826 (N_15826,N_14951,N_14005);
and U15827 (N_15827,N_14039,N_14676);
or U15828 (N_15828,N_14736,N_14855);
xor U15829 (N_15829,N_14995,N_14737);
or U15830 (N_15830,N_14978,N_14243);
nor U15831 (N_15831,N_14393,N_14562);
nand U15832 (N_15832,N_14189,N_14051);
nand U15833 (N_15833,N_14555,N_14198);
xor U15834 (N_15834,N_14203,N_14747);
and U15835 (N_15835,N_14626,N_14338);
nand U15836 (N_15836,N_14659,N_14445);
nand U15837 (N_15837,N_14024,N_14447);
or U15838 (N_15838,N_14896,N_14670);
nand U15839 (N_15839,N_14684,N_14119);
nor U15840 (N_15840,N_14158,N_14963);
or U15841 (N_15841,N_14610,N_14333);
nand U15842 (N_15842,N_14507,N_14829);
xor U15843 (N_15843,N_14538,N_14828);
nor U15844 (N_15844,N_14431,N_14411);
or U15845 (N_15845,N_14699,N_14440);
and U15846 (N_15846,N_14613,N_14245);
xnor U15847 (N_15847,N_14174,N_14880);
nand U15848 (N_15848,N_14201,N_14976);
or U15849 (N_15849,N_14659,N_14668);
nor U15850 (N_15850,N_14042,N_14440);
nand U15851 (N_15851,N_14414,N_14761);
nand U15852 (N_15852,N_14652,N_14164);
or U15853 (N_15853,N_14240,N_14134);
and U15854 (N_15854,N_14204,N_14232);
nor U15855 (N_15855,N_14412,N_14861);
or U15856 (N_15856,N_14017,N_14279);
and U15857 (N_15857,N_14255,N_14026);
and U15858 (N_15858,N_14098,N_14250);
xnor U15859 (N_15859,N_14140,N_14464);
nand U15860 (N_15860,N_14774,N_14249);
or U15861 (N_15861,N_14297,N_14726);
nor U15862 (N_15862,N_14767,N_14131);
and U15863 (N_15863,N_14658,N_14164);
or U15864 (N_15864,N_14926,N_14496);
xor U15865 (N_15865,N_14846,N_14633);
nand U15866 (N_15866,N_14249,N_14076);
nor U15867 (N_15867,N_14165,N_14753);
nand U15868 (N_15868,N_14645,N_14027);
nor U15869 (N_15869,N_14034,N_14700);
or U15870 (N_15870,N_14504,N_14940);
or U15871 (N_15871,N_14577,N_14106);
xnor U15872 (N_15872,N_14017,N_14428);
nand U15873 (N_15873,N_14984,N_14976);
nand U15874 (N_15874,N_14374,N_14089);
xor U15875 (N_15875,N_14007,N_14049);
and U15876 (N_15876,N_14334,N_14874);
and U15877 (N_15877,N_14226,N_14870);
nor U15878 (N_15878,N_14779,N_14265);
nor U15879 (N_15879,N_14951,N_14287);
and U15880 (N_15880,N_14437,N_14698);
xor U15881 (N_15881,N_14704,N_14515);
and U15882 (N_15882,N_14215,N_14266);
or U15883 (N_15883,N_14638,N_14568);
xnor U15884 (N_15884,N_14133,N_14067);
xnor U15885 (N_15885,N_14969,N_14234);
nand U15886 (N_15886,N_14657,N_14441);
or U15887 (N_15887,N_14783,N_14835);
and U15888 (N_15888,N_14363,N_14974);
xnor U15889 (N_15889,N_14416,N_14504);
or U15890 (N_15890,N_14194,N_14975);
xor U15891 (N_15891,N_14046,N_14649);
nand U15892 (N_15892,N_14344,N_14517);
and U15893 (N_15893,N_14586,N_14975);
and U15894 (N_15894,N_14749,N_14452);
nor U15895 (N_15895,N_14022,N_14135);
nand U15896 (N_15896,N_14633,N_14196);
and U15897 (N_15897,N_14790,N_14123);
or U15898 (N_15898,N_14495,N_14391);
or U15899 (N_15899,N_14995,N_14103);
nor U15900 (N_15900,N_14393,N_14421);
or U15901 (N_15901,N_14066,N_14848);
xnor U15902 (N_15902,N_14386,N_14671);
and U15903 (N_15903,N_14084,N_14478);
nand U15904 (N_15904,N_14567,N_14790);
and U15905 (N_15905,N_14047,N_14137);
or U15906 (N_15906,N_14813,N_14333);
nor U15907 (N_15907,N_14435,N_14430);
or U15908 (N_15908,N_14263,N_14968);
or U15909 (N_15909,N_14396,N_14581);
and U15910 (N_15910,N_14944,N_14554);
or U15911 (N_15911,N_14210,N_14537);
nand U15912 (N_15912,N_14974,N_14315);
xnor U15913 (N_15913,N_14177,N_14551);
and U15914 (N_15914,N_14222,N_14358);
and U15915 (N_15915,N_14718,N_14510);
nor U15916 (N_15916,N_14599,N_14723);
nand U15917 (N_15917,N_14675,N_14743);
nand U15918 (N_15918,N_14424,N_14757);
xnor U15919 (N_15919,N_14937,N_14382);
xnor U15920 (N_15920,N_14257,N_14230);
and U15921 (N_15921,N_14461,N_14157);
nand U15922 (N_15922,N_14067,N_14377);
and U15923 (N_15923,N_14731,N_14631);
xnor U15924 (N_15924,N_14774,N_14456);
nor U15925 (N_15925,N_14877,N_14313);
xnor U15926 (N_15926,N_14474,N_14350);
or U15927 (N_15927,N_14278,N_14351);
nor U15928 (N_15928,N_14254,N_14417);
and U15929 (N_15929,N_14288,N_14838);
or U15930 (N_15930,N_14252,N_14167);
xor U15931 (N_15931,N_14612,N_14867);
nand U15932 (N_15932,N_14471,N_14390);
and U15933 (N_15933,N_14746,N_14508);
and U15934 (N_15934,N_14657,N_14872);
xor U15935 (N_15935,N_14500,N_14134);
nor U15936 (N_15936,N_14902,N_14553);
and U15937 (N_15937,N_14018,N_14677);
xor U15938 (N_15938,N_14708,N_14605);
nand U15939 (N_15939,N_14598,N_14067);
or U15940 (N_15940,N_14302,N_14062);
nand U15941 (N_15941,N_14937,N_14928);
and U15942 (N_15942,N_14489,N_14260);
xnor U15943 (N_15943,N_14033,N_14623);
nand U15944 (N_15944,N_14516,N_14893);
and U15945 (N_15945,N_14452,N_14305);
and U15946 (N_15946,N_14413,N_14350);
xor U15947 (N_15947,N_14771,N_14639);
xor U15948 (N_15948,N_14703,N_14473);
or U15949 (N_15949,N_14127,N_14440);
or U15950 (N_15950,N_14629,N_14911);
and U15951 (N_15951,N_14077,N_14845);
or U15952 (N_15952,N_14236,N_14830);
xor U15953 (N_15953,N_14396,N_14426);
nand U15954 (N_15954,N_14068,N_14373);
nor U15955 (N_15955,N_14203,N_14708);
xnor U15956 (N_15956,N_14738,N_14641);
nor U15957 (N_15957,N_14539,N_14460);
and U15958 (N_15958,N_14879,N_14426);
nor U15959 (N_15959,N_14825,N_14804);
xor U15960 (N_15960,N_14192,N_14334);
xnor U15961 (N_15961,N_14592,N_14066);
nand U15962 (N_15962,N_14907,N_14027);
or U15963 (N_15963,N_14614,N_14086);
and U15964 (N_15964,N_14548,N_14033);
nand U15965 (N_15965,N_14503,N_14822);
and U15966 (N_15966,N_14113,N_14782);
nand U15967 (N_15967,N_14500,N_14370);
nand U15968 (N_15968,N_14546,N_14909);
or U15969 (N_15969,N_14550,N_14990);
and U15970 (N_15970,N_14669,N_14849);
and U15971 (N_15971,N_14125,N_14311);
nand U15972 (N_15972,N_14165,N_14780);
nand U15973 (N_15973,N_14650,N_14953);
nor U15974 (N_15974,N_14272,N_14059);
and U15975 (N_15975,N_14010,N_14177);
or U15976 (N_15976,N_14335,N_14190);
or U15977 (N_15977,N_14765,N_14193);
nor U15978 (N_15978,N_14082,N_14614);
xnor U15979 (N_15979,N_14214,N_14746);
nor U15980 (N_15980,N_14151,N_14810);
and U15981 (N_15981,N_14833,N_14908);
and U15982 (N_15982,N_14934,N_14154);
nor U15983 (N_15983,N_14768,N_14973);
or U15984 (N_15984,N_14383,N_14499);
and U15985 (N_15985,N_14607,N_14400);
and U15986 (N_15986,N_14533,N_14768);
or U15987 (N_15987,N_14758,N_14426);
nand U15988 (N_15988,N_14816,N_14999);
and U15989 (N_15989,N_14334,N_14424);
nand U15990 (N_15990,N_14272,N_14814);
nor U15991 (N_15991,N_14073,N_14452);
and U15992 (N_15992,N_14371,N_14877);
xnor U15993 (N_15993,N_14984,N_14943);
nor U15994 (N_15994,N_14638,N_14813);
nor U15995 (N_15995,N_14590,N_14772);
and U15996 (N_15996,N_14654,N_14019);
nand U15997 (N_15997,N_14328,N_14012);
nor U15998 (N_15998,N_14457,N_14279);
or U15999 (N_15999,N_14784,N_14485);
and U16000 (N_16000,N_15057,N_15110);
and U16001 (N_16001,N_15692,N_15915);
nand U16002 (N_16002,N_15631,N_15369);
nor U16003 (N_16003,N_15682,N_15332);
nand U16004 (N_16004,N_15395,N_15404);
and U16005 (N_16005,N_15483,N_15989);
nand U16006 (N_16006,N_15446,N_15724);
nor U16007 (N_16007,N_15664,N_15531);
xnor U16008 (N_16008,N_15272,N_15454);
or U16009 (N_16009,N_15412,N_15835);
or U16010 (N_16010,N_15971,N_15829);
nor U16011 (N_16011,N_15242,N_15154);
and U16012 (N_16012,N_15963,N_15824);
nand U16013 (N_16013,N_15775,N_15912);
nor U16014 (N_16014,N_15252,N_15716);
nand U16015 (N_16015,N_15072,N_15473);
and U16016 (N_16016,N_15778,N_15799);
and U16017 (N_16017,N_15656,N_15800);
xor U16018 (N_16018,N_15334,N_15819);
and U16019 (N_16019,N_15816,N_15795);
nor U16020 (N_16020,N_15425,N_15314);
xnor U16021 (N_16021,N_15893,N_15530);
xnor U16022 (N_16022,N_15373,N_15432);
nor U16023 (N_16023,N_15234,N_15321);
nor U16024 (N_16024,N_15734,N_15186);
nor U16025 (N_16025,N_15102,N_15889);
nor U16026 (N_16026,N_15222,N_15270);
nand U16027 (N_16027,N_15316,N_15838);
nand U16028 (N_16028,N_15653,N_15050);
and U16029 (N_16029,N_15673,N_15054);
nor U16030 (N_16030,N_15268,N_15694);
xnor U16031 (N_16031,N_15043,N_15220);
or U16032 (N_16032,N_15020,N_15198);
and U16033 (N_16033,N_15136,N_15307);
and U16034 (N_16034,N_15698,N_15188);
nand U16035 (N_16035,N_15468,N_15419);
xor U16036 (N_16036,N_15150,N_15637);
xor U16037 (N_16037,N_15986,N_15052);
and U16038 (N_16038,N_15004,N_15133);
and U16039 (N_16039,N_15727,N_15037);
nor U16040 (N_16040,N_15084,N_15647);
nand U16041 (N_16041,N_15710,N_15558);
and U16042 (N_16042,N_15559,N_15488);
xnor U16043 (N_16043,N_15783,N_15494);
or U16044 (N_16044,N_15461,N_15400);
nand U16045 (N_16045,N_15933,N_15143);
and U16046 (N_16046,N_15648,N_15585);
nand U16047 (N_16047,N_15093,N_15833);
nand U16048 (N_16048,N_15191,N_15094);
nand U16049 (N_16049,N_15810,N_15665);
nor U16050 (N_16050,N_15815,N_15428);
nand U16051 (N_16051,N_15828,N_15845);
or U16052 (N_16052,N_15212,N_15658);
nand U16053 (N_16053,N_15927,N_15705);
or U16054 (N_16054,N_15958,N_15359);
and U16055 (N_16055,N_15463,N_15011);
xnor U16056 (N_16056,N_15625,N_15184);
nand U16057 (N_16057,N_15496,N_15257);
xor U16058 (N_16058,N_15134,N_15693);
nor U16059 (N_16059,N_15346,N_15604);
xnor U16060 (N_16060,N_15153,N_15563);
nand U16061 (N_16061,N_15495,N_15409);
xnor U16062 (N_16062,N_15672,N_15993);
xnor U16063 (N_16063,N_15229,N_15621);
or U16064 (N_16064,N_15854,N_15343);
or U16065 (N_16065,N_15196,N_15612);
nor U16066 (N_16066,N_15211,N_15539);
or U16067 (N_16067,N_15051,N_15950);
xnor U16068 (N_16068,N_15367,N_15821);
and U16069 (N_16069,N_15437,N_15561);
or U16070 (N_16070,N_15008,N_15453);
or U16071 (N_16071,N_15183,N_15452);
nand U16072 (N_16072,N_15796,N_15396);
xnor U16073 (N_16073,N_15205,N_15758);
and U16074 (N_16074,N_15661,N_15840);
nand U16075 (N_16075,N_15119,N_15903);
nand U16076 (N_16076,N_15472,N_15328);
nand U16077 (N_16077,N_15597,N_15600);
xnor U16078 (N_16078,N_15309,N_15240);
xnor U16079 (N_16079,N_15269,N_15278);
xnor U16080 (N_16080,N_15598,N_15231);
nor U16081 (N_16081,N_15577,N_15053);
and U16082 (N_16082,N_15784,N_15503);
and U16083 (N_16083,N_15152,N_15027);
nand U16084 (N_16084,N_15471,N_15589);
xnor U16085 (N_16085,N_15139,N_15075);
nor U16086 (N_16086,N_15751,N_15519);
nand U16087 (N_16087,N_15703,N_15267);
nor U16088 (N_16088,N_15813,N_15723);
and U16089 (N_16089,N_15929,N_15258);
xnor U16090 (N_16090,N_15263,N_15785);
nand U16091 (N_16091,N_15545,N_15326);
nor U16092 (N_16092,N_15535,N_15361);
nor U16093 (N_16093,N_15081,N_15206);
or U16094 (N_16094,N_15408,N_15555);
xor U16095 (N_16095,N_15970,N_15961);
xor U16096 (N_16096,N_15031,N_15049);
and U16097 (N_16097,N_15937,N_15747);
and U16098 (N_16098,N_15599,N_15039);
xnor U16099 (N_16099,N_15763,N_15801);
and U16100 (N_16100,N_15552,N_15217);
or U16101 (N_16101,N_15615,N_15485);
nor U16102 (N_16102,N_15650,N_15940);
and U16103 (N_16103,N_15025,N_15624);
nand U16104 (N_16104,N_15034,N_15877);
nor U16105 (N_16105,N_15317,N_15932);
xor U16106 (N_16106,N_15200,N_15870);
and U16107 (N_16107,N_15358,N_15863);
nand U16108 (N_16108,N_15881,N_15144);
and U16109 (N_16109,N_15297,N_15247);
and U16110 (N_16110,N_15406,N_15195);
and U16111 (N_16111,N_15706,N_15233);
nor U16112 (N_16112,N_15931,N_15728);
and U16113 (N_16113,N_15606,N_15001);
xnor U16114 (N_16114,N_15410,N_15869);
nand U16115 (N_16115,N_15323,N_15246);
nand U16116 (N_16116,N_15187,N_15762);
nor U16117 (N_16117,N_15477,N_15510);
or U16118 (N_16118,N_15098,N_15103);
xor U16119 (N_16119,N_15383,N_15900);
or U16120 (N_16120,N_15504,N_15430);
nand U16121 (N_16121,N_15882,N_15590);
nor U16122 (N_16122,N_15807,N_15118);
nor U16123 (N_16123,N_15844,N_15888);
nand U16124 (N_16124,N_15935,N_15142);
nor U16125 (N_16125,N_15106,N_15921);
nor U16126 (N_16126,N_15774,N_15507);
or U16127 (N_16127,N_15666,N_15542);
nand U16128 (N_16128,N_15586,N_15274);
or U16129 (N_16129,N_15111,N_15887);
or U16130 (N_16130,N_15365,N_15038);
and U16131 (N_16131,N_15942,N_15722);
nor U16132 (N_16132,N_15370,N_15294);
xnor U16133 (N_16133,N_15667,N_15540);
xnor U16134 (N_16134,N_15148,N_15424);
xnor U16135 (N_16135,N_15161,N_15416);
and U16136 (N_16136,N_15414,N_15431);
nand U16137 (N_16137,N_15726,N_15130);
xnor U16138 (N_16138,N_15831,N_15567);
nand U16139 (N_16139,N_15415,N_15515);
and U16140 (N_16140,N_15413,N_15898);
and U16141 (N_16141,N_15080,N_15964);
nor U16142 (N_16142,N_15256,N_15547);
nor U16143 (N_16143,N_15078,N_15646);
nand U16144 (N_16144,N_15201,N_15391);
or U16145 (N_16145,N_15591,N_15059);
and U16146 (N_16146,N_15099,N_15875);
nand U16147 (N_16147,N_15861,N_15509);
and U16148 (N_16148,N_15501,N_15614);
nor U16149 (N_16149,N_15228,N_15768);
xnor U16150 (N_16150,N_15864,N_15032);
and U16151 (N_16151,N_15909,N_15982);
xor U16152 (N_16152,N_15732,N_15850);
nor U16153 (N_16153,N_15162,N_15164);
xor U16154 (N_16154,N_15980,N_15021);
nor U16155 (N_16155,N_15189,N_15392);
and U16156 (N_16156,N_15923,N_15947);
xor U16157 (N_16157,N_15737,N_15660);
xor U16158 (N_16158,N_15145,N_15534);
nor U16159 (N_16159,N_15681,N_15438);
or U16160 (N_16160,N_15124,N_15549);
or U16161 (N_16161,N_15680,N_15434);
nor U16162 (N_16162,N_15907,N_15802);
nor U16163 (N_16163,N_15207,N_15042);
nand U16164 (N_16164,N_15114,N_15825);
or U16165 (N_16165,N_15457,N_15679);
nor U16166 (N_16166,N_15718,N_15123);
nand U16167 (N_16167,N_15283,N_15969);
nor U16168 (N_16168,N_15526,N_15752);
and U16169 (N_16169,N_15513,N_15429);
xnor U16170 (N_16170,N_15305,N_15376);
and U16171 (N_16171,N_15822,N_15371);
nand U16172 (N_16172,N_15797,N_15943);
and U16173 (N_16173,N_15366,N_15115);
xor U16174 (N_16174,N_15886,N_15765);
xnor U16175 (N_16175,N_15462,N_15834);
nand U16176 (N_16176,N_15467,N_15704);
nor U16177 (N_16177,N_15872,N_15922);
nand U16178 (N_16178,N_15028,N_15556);
and U16179 (N_16179,N_15421,N_15553);
and U16180 (N_16180,N_15223,N_15451);
xnor U16181 (N_16181,N_15730,N_15325);
or U16182 (N_16182,N_15108,N_15551);
xor U16183 (N_16183,N_15192,N_15753);
xor U16184 (N_16184,N_15262,N_15261);
or U16185 (N_16185,N_15065,N_15310);
nand U16186 (N_16186,N_15230,N_15977);
xnor U16187 (N_16187,N_15487,N_15712);
nor U16188 (N_16188,N_15448,N_15185);
or U16189 (N_16189,N_15444,N_15165);
and U16190 (N_16190,N_15180,N_15683);
nand U16191 (N_16191,N_15689,N_15280);
xnor U16192 (N_16192,N_15327,N_15235);
nor U16193 (N_16193,N_15125,N_15006);
nor U16194 (N_16194,N_15388,N_15630);
nand U16195 (N_16195,N_15351,N_15350);
or U16196 (N_16196,N_15700,N_15178);
and U16197 (N_16197,N_15286,N_15436);
nor U16198 (N_16198,N_15092,N_15901);
and U16199 (N_16199,N_15197,N_15936);
nand U16200 (N_16200,N_15445,N_15867);
and U16201 (N_16201,N_15750,N_15380);
nor U16202 (N_16202,N_15804,N_15973);
or U16203 (N_16203,N_15817,N_15622);
or U16204 (N_16204,N_15739,N_15464);
and U16205 (N_16205,N_15127,N_15789);
nor U16206 (N_16206,N_15173,N_15635);
and U16207 (N_16207,N_15167,N_15896);
xor U16208 (N_16208,N_15465,N_15910);
nor U16209 (N_16209,N_15215,N_15160);
nor U16210 (N_16210,N_15459,N_15492);
xnor U16211 (N_16211,N_15984,N_15097);
and U16212 (N_16212,N_15814,N_15209);
nand U16213 (N_16213,N_15318,N_15190);
nand U16214 (N_16214,N_15299,N_15685);
nor U16215 (N_16215,N_15930,N_15754);
nor U16216 (N_16216,N_15955,N_15422);
nor U16217 (N_16217,N_15911,N_15619);
and U16218 (N_16218,N_15405,N_15095);
or U16219 (N_16219,N_15389,N_15067);
and U16220 (N_16220,N_15315,N_15493);
or U16221 (N_16221,N_15121,N_15548);
and U16222 (N_16222,N_15866,N_15290);
xor U16223 (N_16223,N_15780,N_15251);
xor U16224 (N_16224,N_15588,N_15623);
nand U16225 (N_16225,N_15663,N_15874);
and U16226 (N_16226,N_15998,N_15036);
and U16227 (N_16227,N_15808,N_15276);
nand U16228 (N_16228,N_15518,N_15009);
and U16229 (N_16229,N_15891,N_15523);
nor U16230 (N_16230,N_15557,N_15435);
or U16231 (N_16231,N_15618,N_15224);
and U16232 (N_16232,N_15544,N_15571);
or U16233 (N_16233,N_15498,N_15846);
nor U16234 (N_16234,N_15678,N_15480);
nor U16235 (N_16235,N_15959,N_15460);
or U16236 (N_16236,N_15066,N_15331);
xor U16237 (N_16237,N_15729,N_15566);
nand U16238 (N_16238,N_15071,N_15573);
xor U16239 (N_16239,N_15720,N_15827);
and U16240 (N_16240,N_15879,N_15628);
xnor U16241 (N_16241,N_15293,N_15745);
and U16242 (N_16242,N_15607,N_15669);
nand U16243 (N_16243,N_15756,N_15988);
xor U16244 (N_16244,N_15748,N_15354);
and U16245 (N_16245,N_15735,N_15281);
nor U16246 (N_16246,N_15525,N_15776);
xnor U16247 (N_16247,N_15805,N_15478);
xnor U16248 (N_16248,N_15203,N_15104);
or U16249 (N_16249,N_15868,N_15760);
nand U16250 (N_16250,N_15643,N_15733);
nand U16251 (N_16251,N_15061,N_15981);
nand U16252 (N_16252,N_15311,N_15949);
nor U16253 (N_16253,N_15426,N_15449);
or U16254 (N_16254,N_15347,N_15100);
nand U16255 (N_16255,N_15122,N_15965);
or U16256 (N_16256,N_15137,N_15960);
nand U16257 (N_16257,N_15368,N_15766);
nor U16258 (N_16258,N_15594,N_15506);
nand U16259 (N_16259,N_15096,N_15255);
nor U16260 (N_16260,N_15237,N_15356);
or U16261 (N_16261,N_15968,N_15069);
nor U16262 (N_16262,N_15632,N_15338);
nand U16263 (N_16263,N_15301,N_15684);
or U16264 (N_16264,N_15996,N_15013);
nor U16265 (N_16265,N_15849,N_15285);
nor U16266 (N_16266,N_15742,N_15441);
nor U16267 (N_16267,N_15583,N_15402);
or U16268 (N_16268,N_15300,N_15966);
nor U16269 (N_16269,N_15895,N_15107);
nor U16270 (N_16270,N_15344,N_15670);
nor U16271 (N_16271,N_15994,N_15364);
and U16272 (N_16272,N_15490,N_15469);
xor U16273 (N_16273,N_15399,N_15719);
nand U16274 (N_16274,N_15481,N_15403);
and U16275 (N_16275,N_15759,N_15482);
nor U16276 (N_16276,N_15517,N_15091);
xnor U16277 (N_16277,N_15083,N_15638);
and U16278 (N_16278,N_15582,N_15138);
nor U16279 (N_16279,N_15826,N_15873);
nand U16280 (N_16280,N_15339,N_15226);
nand U16281 (N_16281,N_15499,N_15668);
nor U16282 (N_16282,N_15639,N_15738);
xnor U16283 (N_16283,N_15836,N_15537);
and U16284 (N_16284,N_15883,N_15362);
nor U16285 (N_16285,N_15843,N_15128);
xnor U16286 (N_16286,N_15047,N_15131);
nor U16287 (N_16287,N_15767,N_15238);
and U16288 (N_16288,N_15857,N_15502);
and U16289 (N_16289,N_15852,N_15956);
nand U16290 (N_16290,N_15676,N_15112);
xnor U16291 (N_16291,N_15120,N_15374);
nor U16292 (N_16292,N_15687,N_15079);
xnor U16293 (N_16293,N_15791,N_15035);
xor U16294 (N_16294,N_15533,N_15790);
or U16295 (N_16295,N_15713,N_15254);
or U16296 (N_16296,N_15897,N_15295);
nand U16297 (N_16297,N_15662,N_15610);
or U16298 (N_16298,N_15208,N_15860);
or U16299 (N_16299,N_15992,N_15626);
nand U16300 (N_16300,N_15524,N_15798);
xnor U16301 (N_16301,N_15884,N_15902);
nand U16302 (N_16302,N_15249,N_15474);
nor U16303 (N_16303,N_15497,N_15236);
nor U16304 (N_16304,N_15045,N_15945);
and U16305 (N_16305,N_15709,N_15906);
and U16306 (N_16306,N_15129,N_15363);
and U16307 (N_16307,N_15905,N_15644);
nor U16308 (N_16308,N_15440,N_15529);
xnor U16309 (N_16309,N_15641,N_15491);
xnor U16310 (N_16310,N_15764,N_15918);
nor U16311 (N_16311,N_15455,N_15948);
nand U16312 (N_16312,N_15926,N_15890);
and U16313 (N_16313,N_15014,N_15450);
nand U16314 (N_16314,N_15155,N_15859);
nor U16315 (N_16315,N_15608,N_15749);
or U16316 (N_16316,N_15357,N_15755);
xnor U16317 (N_16317,N_15611,N_15407);
nand U16318 (N_16318,N_15972,N_15026);
xnor U16319 (N_16319,N_15175,N_15593);
xor U16320 (N_16320,N_15077,N_15194);
nand U16321 (N_16321,N_15627,N_15292);
nor U16322 (N_16322,N_15584,N_15166);
and U16323 (N_16323,N_15018,N_15983);
and U16324 (N_16324,N_15736,N_15904);
and U16325 (N_16325,N_15287,N_15041);
xor U16326 (N_16326,N_15411,N_15925);
nand U16327 (N_16327,N_15439,N_15924);
and U16328 (N_16328,N_15782,N_15731);
nor U16329 (N_16329,N_15997,N_15058);
or U16330 (N_16330,N_15550,N_15076);
nor U16331 (N_16331,N_15617,N_15337);
xnor U16332 (N_16332,N_15105,N_15174);
or U16333 (N_16333,N_15353,N_15033);
or U16334 (N_16334,N_15177,N_15382);
nand U16335 (N_16335,N_15914,N_15913);
or U16336 (N_16336,N_15385,N_15330);
nand U16337 (N_16337,N_15141,N_15587);
nand U16338 (N_16338,N_15387,N_15862);
and U16339 (N_16339,N_15946,N_15987);
xor U16340 (N_16340,N_15516,N_15740);
xor U16341 (N_16341,N_15288,N_15398);
and U16342 (N_16342,N_15596,N_15851);
and U16343 (N_16343,N_15158,N_15048);
nand U16344 (N_16344,N_15579,N_15642);
xor U16345 (N_16345,N_15086,N_15847);
or U16346 (N_16346,N_15458,N_15225);
and U16347 (N_16347,N_15349,N_15788);
or U16348 (N_16348,N_15417,N_15401);
or U16349 (N_16349,N_15541,N_15885);
nor U16350 (N_16350,N_15320,N_15620);
nand U16351 (N_16351,N_15696,N_15447);
nand U16352 (N_16352,N_15830,N_15919);
and U16353 (N_16353,N_15470,N_15007);
or U16354 (N_16354,N_15794,N_15109);
nand U16355 (N_16355,N_15147,N_15022);
xor U16356 (N_16356,N_15172,N_15976);
xnor U16357 (N_16357,N_15303,N_15538);
nor U16358 (N_16358,N_15871,N_15313);
nor U16359 (N_16359,N_15773,N_15779);
nand U16360 (N_16360,N_15721,N_15677);
nand U16361 (N_16361,N_15146,N_15312);
and U16362 (N_16362,N_15999,N_15319);
or U16363 (N_16363,N_15671,N_15938);
nor U16364 (N_16364,N_15466,N_15360);
or U16365 (N_16365,N_15974,N_15170);
or U16366 (N_16366,N_15811,N_15675);
nor U16367 (N_16367,N_15786,N_15015);
xor U16368 (N_16368,N_15690,N_15711);
xnor U16369 (N_16369,N_15304,N_15030);
xnor U16370 (N_16370,N_15633,N_15341);
xnor U16371 (N_16371,N_15159,N_15275);
nand U16372 (N_16372,N_15335,N_15543);
and U16373 (N_16373,N_15378,N_15219);
nor U16374 (N_16374,N_15908,N_15652);
or U16375 (N_16375,N_15717,N_15241);
xor U16376 (N_16376,N_15651,N_15302);
or U16377 (N_16377,N_15560,N_15839);
or U16378 (N_16378,N_15342,N_15757);
and U16379 (N_16379,N_15044,N_15595);
nand U16380 (N_16380,N_15605,N_15239);
or U16381 (N_16381,N_15602,N_15204);
or U16382 (N_16382,N_15232,N_15005);
nand U16383 (N_16383,N_15761,N_15010);
or U16384 (N_16384,N_15592,N_15135);
xor U16385 (N_16385,N_15837,N_15634);
and U16386 (N_16386,N_15536,N_15616);
and U16387 (N_16387,N_15126,N_15771);
and U16388 (N_16388,N_15149,N_15939);
or U16389 (N_16389,N_15772,N_15393);
nand U16390 (N_16390,N_15169,N_15024);
nor U16391 (N_16391,N_15580,N_15306);
or U16392 (N_16392,N_15777,N_15348);
xnor U16393 (N_16393,N_15101,N_15132);
and U16394 (N_16394,N_15016,N_15390);
nor U16395 (N_16395,N_15420,N_15140);
or U16396 (N_16396,N_15744,N_15995);
nand U16397 (N_16397,N_15565,N_15266);
nor U16398 (N_16398,N_15019,N_15087);
or U16399 (N_16399,N_15842,N_15714);
or U16400 (N_16400,N_15029,N_15521);
nor U16401 (N_16401,N_15832,N_15090);
and U16402 (N_16402,N_15823,N_15952);
nand U16403 (N_16403,N_15284,N_15377);
nand U16404 (N_16404,N_15532,N_15271);
nand U16405 (N_16405,N_15527,N_15576);
nand U16406 (N_16406,N_15500,N_15578);
xnor U16407 (N_16407,N_15916,N_15291);
nor U16408 (N_16408,N_15182,N_15193);
and U16409 (N_16409,N_15741,N_15277);
and U16410 (N_16410,N_15333,N_15117);
nor U16411 (N_16411,N_15990,N_15978);
nor U16412 (N_16412,N_15528,N_15725);
and U16413 (N_16413,N_15688,N_15944);
xnor U16414 (N_16414,N_15645,N_15227);
or U16415 (N_16415,N_15967,N_15522);
or U16416 (N_16416,N_15848,N_15433);
and U16417 (N_16417,N_15324,N_15442);
nand U16418 (N_16418,N_15085,N_15427);
nor U16419 (N_16419,N_15418,N_15171);
or U16420 (N_16420,N_15296,N_15699);
nor U16421 (N_16421,N_15562,N_15329);
nor U16422 (N_16422,N_15655,N_15384);
nand U16423 (N_16423,N_15787,N_15456);
nor U16424 (N_16424,N_15248,N_15002);
xnor U16425 (N_16425,N_15017,N_15476);
nand U16426 (N_16426,N_15259,N_15064);
or U16427 (N_16427,N_15218,N_15708);
xnor U16428 (N_16428,N_15214,N_15489);
or U16429 (N_16429,N_15055,N_15156);
nor U16430 (N_16430,N_15962,N_15264);
nor U16431 (N_16431,N_15336,N_15023);
xor U16432 (N_16432,N_15572,N_15697);
nand U16433 (N_16433,N_15088,N_15063);
xnor U16434 (N_16434,N_15954,N_15957);
nor U16435 (N_16435,N_15289,N_15279);
nand U16436 (N_16436,N_15878,N_15659);
nor U16437 (N_16437,N_15941,N_15820);
nor U16438 (N_16438,N_15743,N_15570);
xnor U16439 (N_16439,N_15221,N_15340);
xor U16440 (N_16440,N_15654,N_15253);
xnor U16441 (N_16441,N_15265,N_15701);
and U16442 (N_16442,N_15116,N_15928);
nor U16443 (N_16443,N_15951,N_15818);
or U16444 (N_16444,N_15674,N_15769);
xor U16445 (N_16445,N_15899,N_15979);
and U16446 (N_16446,N_15073,N_15479);
nor U16447 (N_16447,N_15691,N_15089);
or U16448 (N_16448,N_15991,N_15636);
nand U16449 (N_16449,N_15486,N_15355);
nor U16450 (N_16450,N_15702,N_15372);
xnor U16451 (N_16451,N_15056,N_15640);
nand U16452 (N_16452,N_15520,N_15345);
xor U16453 (N_16453,N_15746,N_15574);
or U16454 (N_16454,N_15803,N_15375);
xnor U16455 (N_16455,N_15397,N_15841);
and U16456 (N_16456,N_15003,N_15381);
xor U16457 (N_16457,N_15386,N_15322);
nand U16458 (N_16458,N_15423,N_15202);
or U16459 (N_16459,N_15512,N_15216);
nand U16460 (N_16460,N_15157,N_15012);
nor U16461 (N_16461,N_15603,N_15809);
or U16462 (N_16462,N_15853,N_15657);
nor U16463 (N_16463,N_15505,N_15770);
nand U16464 (N_16464,N_15113,N_15715);
and U16465 (N_16465,N_15394,N_15273);
and U16466 (N_16466,N_15975,N_15168);
and U16467 (N_16467,N_15514,N_15298);
xor U16468 (N_16468,N_15686,N_15151);
or U16469 (N_16469,N_15876,N_15199);
nor U16470 (N_16470,N_15554,N_15581);
nor U16471 (N_16471,N_15250,N_15781);
and U16472 (N_16472,N_15181,N_15568);
nand U16473 (N_16473,N_15985,N_15892);
nand U16474 (N_16474,N_15244,N_15649);
or U16475 (N_16475,N_15856,N_15060);
nor U16476 (N_16476,N_15858,N_15601);
and U16477 (N_16477,N_15613,N_15046);
nand U16478 (N_16478,N_15920,N_15179);
or U16479 (N_16479,N_15934,N_15210);
nor U16480 (N_16480,N_15484,N_15569);
and U16481 (N_16481,N_15308,N_15880);
xor U16482 (N_16482,N_15792,N_15917);
or U16483 (N_16483,N_15243,N_15575);
xnor U16484 (N_16484,N_15260,N_15855);
xnor U16485 (N_16485,N_15082,N_15475);
or U16486 (N_16486,N_15163,N_15707);
xnor U16487 (N_16487,N_15245,N_15213);
xor U16488 (N_16488,N_15070,N_15443);
or U16489 (N_16489,N_15865,N_15609);
nand U16490 (N_16490,N_15806,N_15629);
nor U16491 (N_16491,N_15068,N_15953);
or U16492 (N_16492,N_15379,N_15564);
or U16493 (N_16493,N_15074,N_15352);
nand U16494 (N_16494,N_15000,N_15282);
and U16495 (N_16495,N_15546,N_15511);
nor U16496 (N_16496,N_15894,N_15062);
and U16497 (N_16497,N_15793,N_15176);
or U16498 (N_16498,N_15695,N_15812);
nand U16499 (N_16499,N_15040,N_15508);
or U16500 (N_16500,N_15103,N_15978);
or U16501 (N_16501,N_15123,N_15759);
and U16502 (N_16502,N_15548,N_15648);
nand U16503 (N_16503,N_15470,N_15453);
nor U16504 (N_16504,N_15153,N_15231);
nor U16505 (N_16505,N_15575,N_15521);
nor U16506 (N_16506,N_15294,N_15101);
or U16507 (N_16507,N_15998,N_15260);
or U16508 (N_16508,N_15009,N_15797);
and U16509 (N_16509,N_15963,N_15196);
xnor U16510 (N_16510,N_15359,N_15530);
or U16511 (N_16511,N_15200,N_15865);
nand U16512 (N_16512,N_15569,N_15781);
nor U16513 (N_16513,N_15466,N_15823);
xnor U16514 (N_16514,N_15692,N_15799);
xor U16515 (N_16515,N_15411,N_15975);
nand U16516 (N_16516,N_15423,N_15759);
and U16517 (N_16517,N_15793,N_15694);
nand U16518 (N_16518,N_15521,N_15390);
nand U16519 (N_16519,N_15469,N_15619);
and U16520 (N_16520,N_15066,N_15085);
nor U16521 (N_16521,N_15948,N_15520);
nor U16522 (N_16522,N_15432,N_15595);
xor U16523 (N_16523,N_15283,N_15211);
nand U16524 (N_16524,N_15021,N_15738);
xnor U16525 (N_16525,N_15543,N_15848);
nor U16526 (N_16526,N_15199,N_15256);
nor U16527 (N_16527,N_15617,N_15161);
xor U16528 (N_16528,N_15794,N_15480);
xor U16529 (N_16529,N_15404,N_15970);
nor U16530 (N_16530,N_15714,N_15418);
and U16531 (N_16531,N_15662,N_15612);
nor U16532 (N_16532,N_15573,N_15371);
and U16533 (N_16533,N_15371,N_15929);
nor U16534 (N_16534,N_15998,N_15153);
and U16535 (N_16535,N_15450,N_15884);
xor U16536 (N_16536,N_15251,N_15049);
nor U16537 (N_16537,N_15565,N_15729);
nor U16538 (N_16538,N_15426,N_15283);
and U16539 (N_16539,N_15397,N_15280);
nand U16540 (N_16540,N_15200,N_15197);
and U16541 (N_16541,N_15693,N_15954);
and U16542 (N_16542,N_15404,N_15266);
nor U16543 (N_16543,N_15814,N_15669);
xnor U16544 (N_16544,N_15669,N_15642);
xor U16545 (N_16545,N_15023,N_15819);
xnor U16546 (N_16546,N_15588,N_15284);
nand U16547 (N_16547,N_15842,N_15047);
xor U16548 (N_16548,N_15866,N_15893);
nand U16549 (N_16549,N_15558,N_15517);
or U16550 (N_16550,N_15066,N_15968);
nor U16551 (N_16551,N_15330,N_15849);
or U16552 (N_16552,N_15048,N_15529);
and U16553 (N_16553,N_15350,N_15806);
nand U16554 (N_16554,N_15828,N_15257);
xnor U16555 (N_16555,N_15675,N_15526);
and U16556 (N_16556,N_15783,N_15798);
or U16557 (N_16557,N_15709,N_15998);
nor U16558 (N_16558,N_15867,N_15420);
nor U16559 (N_16559,N_15604,N_15300);
nor U16560 (N_16560,N_15304,N_15886);
nor U16561 (N_16561,N_15960,N_15741);
or U16562 (N_16562,N_15382,N_15215);
nor U16563 (N_16563,N_15042,N_15863);
nor U16564 (N_16564,N_15902,N_15638);
and U16565 (N_16565,N_15682,N_15564);
or U16566 (N_16566,N_15494,N_15210);
or U16567 (N_16567,N_15483,N_15550);
or U16568 (N_16568,N_15536,N_15777);
nor U16569 (N_16569,N_15916,N_15938);
nand U16570 (N_16570,N_15396,N_15713);
or U16571 (N_16571,N_15207,N_15444);
and U16572 (N_16572,N_15464,N_15983);
and U16573 (N_16573,N_15235,N_15936);
nand U16574 (N_16574,N_15119,N_15271);
and U16575 (N_16575,N_15083,N_15022);
and U16576 (N_16576,N_15169,N_15492);
or U16577 (N_16577,N_15255,N_15919);
xnor U16578 (N_16578,N_15522,N_15885);
nand U16579 (N_16579,N_15264,N_15308);
xor U16580 (N_16580,N_15653,N_15220);
xnor U16581 (N_16581,N_15340,N_15909);
and U16582 (N_16582,N_15018,N_15944);
nor U16583 (N_16583,N_15013,N_15116);
or U16584 (N_16584,N_15833,N_15324);
or U16585 (N_16585,N_15946,N_15836);
xor U16586 (N_16586,N_15093,N_15750);
xnor U16587 (N_16587,N_15874,N_15350);
and U16588 (N_16588,N_15680,N_15554);
nor U16589 (N_16589,N_15351,N_15221);
nor U16590 (N_16590,N_15618,N_15085);
nor U16591 (N_16591,N_15319,N_15566);
and U16592 (N_16592,N_15233,N_15444);
and U16593 (N_16593,N_15418,N_15498);
nand U16594 (N_16594,N_15472,N_15700);
and U16595 (N_16595,N_15065,N_15608);
or U16596 (N_16596,N_15808,N_15524);
and U16597 (N_16597,N_15946,N_15041);
or U16598 (N_16598,N_15760,N_15969);
or U16599 (N_16599,N_15301,N_15501);
nand U16600 (N_16600,N_15997,N_15468);
and U16601 (N_16601,N_15238,N_15184);
and U16602 (N_16602,N_15629,N_15264);
xnor U16603 (N_16603,N_15511,N_15706);
nand U16604 (N_16604,N_15171,N_15051);
nor U16605 (N_16605,N_15388,N_15613);
or U16606 (N_16606,N_15695,N_15551);
xnor U16607 (N_16607,N_15268,N_15681);
nor U16608 (N_16608,N_15569,N_15389);
nor U16609 (N_16609,N_15039,N_15132);
xnor U16610 (N_16610,N_15570,N_15018);
nand U16611 (N_16611,N_15364,N_15593);
and U16612 (N_16612,N_15334,N_15040);
nor U16613 (N_16613,N_15297,N_15906);
or U16614 (N_16614,N_15068,N_15728);
nor U16615 (N_16615,N_15114,N_15975);
xor U16616 (N_16616,N_15340,N_15589);
nand U16617 (N_16617,N_15391,N_15290);
and U16618 (N_16618,N_15301,N_15005);
and U16619 (N_16619,N_15969,N_15082);
or U16620 (N_16620,N_15433,N_15197);
nor U16621 (N_16621,N_15520,N_15790);
or U16622 (N_16622,N_15267,N_15069);
xor U16623 (N_16623,N_15936,N_15480);
nand U16624 (N_16624,N_15638,N_15569);
or U16625 (N_16625,N_15303,N_15913);
and U16626 (N_16626,N_15950,N_15671);
nand U16627 (N_16627,N_15965,N_15488);
nor U16628 (N_16628,N_15242,N_15542);
and U16629 (N_16629,N_15044,N_15923);
xor U16630 (N_16630,N_15984,N_15837);
nand U16631 (N_16631,N_15405,N_15972);
nor U16632 (N_16632,N_15808,N_15865);
or U16633 (N_16633,N_15817,N_15465);
nor U16634 (N_16634,N_15715,N_15892);
and U16635 (N_16635,N_15349,N_15886);
nor U16636 (N_16636,N_15048,N_15949);
and U16637 (N_16637,N_15782,N_15544);
nand U16638 (N_16638,N_15298,N_15447);
nand U16639 (N_16639,N_15930,N_15097);
xor U16640 (N_16640,N_15366,N_15918);
and U16641 (N_16641,N_15833,N_15819);
and U16642 (N_16642,N_15448,N_15989);
xnor U16643 (N_16643,N_15004,N_15593);
or U16644 (N_16644,N_15863,N_15953);
nor U16645 (N_16645,N_15728,N_15898);
nand U16646 (N_16646,N_15906,N_15630);
or U16647 (N_16647,N_15808,N_15758);
and U16648 (N_16648,N_15342,N_15248);
and U16649 (N_16649,N_15634,N_15650);
nand U16650 (N_16650,N_15831,N_15143);
nor U16651 (N_16651,N_15654,N_15836);
nor U16652 (N_16652,N_15057,N_15218);
or U16653 (N_16653,N_15102,N_15814);
xnor U16654 (N_16654,N_15793,N_15096);
nor U16655 (N_16655,N_15150,N_15640);
nor U16656 (N_16656,N_15596,N_15297);
or U16657 (N_16657,N_15248,N_15508);
and U16658 (N_16658,N_15755,N_15480);
and U16659 (N_16659,N_15027,N_15612);
or U16660 (N_16660,N_15386,N_15018);
nand U16661 (N_16661,N_15416,N_15846);
xnor U16662 (N_16662,N_15936,N_15064);
xor U16663 (N_16663,N_15180,N_15385);
nor U16664 (N_16664,N_15710,N_15394);
or U16665 (N_16665,N_15695,N_15610);
nand U16666 (N_16666,N_15871,N_15269);
nor U16667 (N_16667,N_15454,N_15294);
xor U16668 (N_16668,N_15945,N_15249);
nor U16669 (N_16669,N_15179,N_15527);
and U16670 (N_16670,N_15943,N_15374);
and U16671 (N_16671,N_15352,N_15598);
and U16672 (N_16672,N_15633,N_15818);
or U16673 (N_16673,N_15332,N_15669);
nor U16674 (N_16674,N_15180,N_15478);
and U16675 (N_16675,N_15766,N_15791);
nand U16676 (N_16676,N_15858,N_15646);
and U16677 (N_16677,N_15345,N_15859);
and U16678 (N_16678,N_15574,N_15265);
nor U16679 (N_16679,N_15031,N_15412);
nor U16680 (N_16680,N_15502,N_15969);
nand U16681 (N_16681,N_15148,N_15057);
and U16682 (N_16682,N_15943,N_15800);
nand U16683 (N_16683,N_15423,N_15637);
or U16684 (N_16684,N_15129,N_15517);
xor U16685 (N_16685,N_15302,N_15327);
and U16686 (N_16686,N_15316,N_15259);
and U16687 (N_16687,N_15471,N_15939);
xor U16688 (N_16688,N_15745,N_15838);
and U16689 (N_16689,N_15182,N_15924);
xor U16690 (N_16690,N_15012,N_15719);
and U16691 (N_16691,N_15397,N_15265);
nor U16692 (N_16692,N_15331,N_15266);
and U16693 (N_16693,N_15373,N_15310);
or U16694 (N_16694,N_15439,N_15524);
xnor U16695 (N_16695,N_15054,N_15482);
nor U16696 (N_16696,N_15275,N_15858);
nor U16697 (N_16697,N_15789,N_15497);
nand U16698 (N_16698,N_15496,N_15296);
nand U16699 (N_16699,N_15868,N_15899);
or U16700 (N_16700,N_15407,N_15724);
nor U16701 (N_16701,N_15484,N_15868);
or U16702 (N_16702,N_15223,N_15575);
nor U16703 (N_16703,N_15773,N_15046);
or U16704 (N_16704,N_15480,N_15868);
nand U16705 (N_16705,N_15153,N_15736);
xor U16706 (N_16706,N_15772,N_15445);
and U16707 (N_16707,N_15830,N_15424);
nand U16708 (N_16708,N_15803,N_15832);
and U16709 (N_16709,N_15075,N_15302);
nand U16710 (N_16710,N_15538,N_15656);
nand U16711 (N_16711,N_15752,N_15612);
and U16712 (N_16712,N_15542,N_15630);
nand U16713 (N_16713,N_15504,N_15177);
nor U16714 (N_16714,N_15219,N_15457);
xnor U16715 (N_16715,N_15609,N_15336);
nor U16716 (N_16716,N_15753,N_15625);
nand U16717 (N_16717,N_15450,N_15897);
nand U16718 (N_16718,N_15584,N_15476);
nand U16719 (N_16719,N_15300,N_15871);
nor U16720 (N_16720,N_15706,N_15342);
or U16721 (N_16721,N_15043,N_15202);
nor U16722 (N_16722,N_15847,N_15881);
nor U16723 (N_16723,N_15344,N_15951);
xnor U16724 (N_16724,N_15496,N_15588);
nand U16725 (N_16725,N_15631,N_15026);
nand U16726 (N_16726,N_15095,N_15274);
or U16727 (N_16727,N_15319,N_15092);
or U16728 (N_16728,N_15603,N_15075);
nand U16729 (N_16729,N_15730,N_15690);
nand U16730 (N_16730,N_15914,N_15011);
nor U16731 (N_16731,N_15325,N_15896);
nand U16732 (N_16732,N_15744,N_15038);
nand U16733 (N_16733,N_15076,N_15123);
nor U16734 (N_16734,N_15734,N_15642);
nor U16735 (N_16735,N_15190,N_15720);
and U16736 (N_16736,N_15886,N_15162);
nand U16737 (N_16737,N_15393,N_15229);
nand U16738 (N_16738,N_15462,N_15302);
nor U16739 (N_16739,N_15179,N_15105);
xor U16740 (N_16740,N_15311,N_15102);
xnor U16741 (N_16741,N_15118,N_15709);
nand U16742 (N_16742,N_15883,N_15989);
nand U16743 (N_16743,N_15135,N_15588);
or U16744 (N_16744,N_15158,N_15588);
nor U16745 (N_16745,N_15611,N_15597);
xor U16746 (N_16746,N_15252,N_15051);
xnor U16747 (N_16747,N_15802,N_15888);
and U16748 (N_16748,N_15127,N_15088);
and U16749 (N_16749,N_15830,N_15543);
and U16750 (N_16750,N_15391,N_15897);
xnor U16751 (N_16751,N_15129,N_15154);
or U16752 (N_16752,N_15045,N_15385);
nand U16753 (N_16753,N_15008,N_15749);
nand U16754 (N_16754,N_15233,N_15111);
xor U16755 (N_16755,N_15787,N_15268);
xnor U16756 (N_16756,N_15465,N_15034);
nand U16757 (N_16757,N_15176,N_15923);
nor U16758 (N_16758,N_15225,N_15582);
or U16759 (N_16759,N_15402,N_15225);
or U16760 (N_16760,N_15596,N_15739);
xnor U16761 (N_16761,N_15297,N_15980);
xor U16762 (N_16762,N_15906,N_15553);
and U16763 (N_16763,N_15159,N_15481);
nand U16764 (N_16764,N_15874,N_15841);
xnor U16765 (N_16765,N_15727,N_15685);
xnor U16766 (N_16766,N_15767,N_15126);
and U16767 (N_16767,N_15900,N_15084);
nor U16768 (N_16768,N_15609,N_15207);
nand U16769 (N_16769,N_15435,N_15086);
or U16770 (N_16770,N_15058,N_15714);
nand U16771 (N_16771,N_15196,N_15921);
xnor U16772 (N_16772,N_15639,N_15743);
nor U16773 (N_16773,N_15741,N_15547);
nand U16774 (N_16774,N_15274,N_15744);
xnor U16775 (N_16775,N_15438,N_15163);
xnor U16776 (N_16776,N_15512,N_15694);
or U16777 (N_16777,N_15034,N_15481);
nor U16778 (N_16778,N_15930,N_15809);
nor U16779 (N_16779,N_15678,N_15761);
xor U16780 (N_16780,N_15035,N_15829);
and U16781 (N_16781,N_15592,N_15691);
xor U16782 (N_16782,N_15609,N_15356);
nand U16783 (N_16783,N_15540,N_15168);
and U16784 (N_16784,N_15968,N_15311);
xor U16785 (N_16785,N_15563,N_15241);
nand U16786 (N_16786,N_15006,N_15840);
nand U16787 (N_16787,N_15701,N_15416);
and U16788 (N_16788,N_15016,N_15221);
and U16789 (N_16789,N_15291,N_15584);
xor U16790 (N_16790,N_15978,N_15788);
or U16791 (N_16791,N_15075,N_15256);
xor U16792 (N_16792,N_15483,N_15015);
nand U16793 (N_16793,N_15073,N_15565);
nor U16794 (N_16794,N_15707,N_15860);
xor U16795 (N_16795,N_15779,N_15890);
nand U16796 (N_16796,N_15268,N_15111);
nand U16797 (N_16797,N_15710,N_15306);
and U16798 (N_16798,N_15217,N_15119);
and U16799 (N_16799,N_15699,N_15270);
nor U16800 (N_16800,N_15324,N_15347);
nor U16801 (N_16801,N_15851,N_15145);
or U16802 (N_16802,N_15240,N_15605);
nor U16803 (N_16803,N_15049,N_15819);
or U16804 (N_16804,N_15553,N_15848);
nor U16805 (N_16805,N_15342,N_15705);
and U16806 (N_16806,N_15478,N_15883);
or U16807 (N_16807,N_15622,N_15765);
nor U16808 (N_16808,N_15725,N_15949);
nor U16809 (N_16809,N_15613,N_15990);
nand U16810 (N_16810,N_15030,N_15097);
xor U16811 (N_16811,N_15334,N_15898);
nor U16812 (N_16812,N_15693,N_15714);
and U16813 (N_16813,N_15660,N_15691);
and U16814 (N_16814,N_15372,N_15300);
and U16815 (N_16815,N_15155,N_15551);
or U16816 (N_16816,N_15666,N_15002);
nor U16817 (N_16817,N_15877,N_15529);
nand U16818 (N_16818,N_15736,N_15156);
and U16819 (N_16819,N_15177,N_15009);
xnor U16820 (N_16820,N_15947,N_15100);
nor U16821 (N_16821,N_15307,N_15891);
and U16822 (N_16822,N_15667,N_15098);
nand U16823 (N_16823,N_15831,N_15250);
nand U16824 (N_16824,N_15484,N_15220);
and U16825 (N_16825,N_15753,N_15649);
or U16826 (N_16826,N_15818,N_15447);
nand U16827 (N_16827,N_15184,N_15622);
xnor U16828 (N_16828,N_15187,N_15678);
and U16829 (N_16829,N_15519,N_15703);
and U16830 (N_16830,N_15092,N_15469);
nand U16831 (N_16831,N_15107,N_15148);
nor U16832 (N_16832,N_15557,N_15645);
or U16833 (N_16833,N_15920,N_15826);
and U16834 (N_16834,N_15382,N_15575);
nor U16835 (N_16835,N_15203,N_15806);
and U16836 (N_16836,N_15949,N_15285);
nor U16837 (N_16837,N_15581,N_15037);
xnor U16838 (N_16838,N_15927,N_15348);
and U16839 (N_16839,N_15031,N_15475);
xor U16840 (N_16840,N_15472,N_15789);
or U16841 (N_16841,N_15441,N_15764);
or U16842 (N_16842,N_15607,N_15379);
nor U16843 (N_16843,N_15084,N_15322);
and U16844 (N_16844,N_15947,N_15391);
nor U16845 (N_16845,N_15448,N_15297);
and U16846 (N_16846,N_15032,N_15050);
xor U16847 (N_16847,N_15587,N_15768);
and U16848 (N_16848,N_15186,N_15110);
xor U16849 (N_16849,N_15920,N_15631);
or U16850 (N_16850,N_15398,N_15306);
nor U16851 (N_16851,N_15702,N_15440);
nand U16852 (N_16852,N_15603,N_15769);
and U16853 (N_16853,N_15017,N_15431);
nand U16854 (N_16854,N_15455,N_15047);
or U16855 (N_16855,N_15342,N_15736);
xnor U16856 (N_16856,N_15176,N_15464);
and U16857 (N_16857,N_15441,N_15191);
xnor U16858 (N_16858,N_15766,N_15730);
or U16859 (N_16859,N_15136,N_15508);
nor U16860 (N_16860,N_15965,N_15864);
xnor U16861 (N_16861,N_15833,N_15065);
nand U16862 (N_16862,N_15404,N_15084);
xor U16863 (N_16863,N_15235,N_15643);
nor U16864 (N_16864,N_15185,N_15918);
and U16865 (N_16865,N_15060,N_15371);
and U16866 (N_16866,N_15306,N_15242);
xnor U16867 (N_16867,N_15842,N_15987);
or U16868 (N_16868,N_15136,N_15799);
nor U16869 (N_16869,N_15687,N_15180);
and U16870 (N_16870,N_15807,N_15891);
and U16871 (N_16871,N_15239,N_15873);
or U16872 (N_16872,N_15345,N_15327);
nand U16873 (N_16873,N_15654,N_15977);
nor U16874 (N_16874,N_15151,N_15871);
nor U16875 (N_16875,N_15575,N_15333);
or U16876 (N_16876,N_15438,N_15596);
xnor U16877 (N_16877,N_15595,N_15392);
nor U16878 (N_16878,N_15863,N_15709);
xor U16879 (N_16879,N_15840,N_15656);
xnor U16880 (N_16880,N_15867,N_15466);
or U16881 (N_16881,N_15016,N_15015);
nor U16882 (N_16882,N_15000,N_15079);
nor U16883 (N_16883,N_15019,N_15665);
and U16884 (N_16884,N_15749,N_15263);
xor U16885 (N_16885,N_15984,N_15241);
xor U16886 (N_16886,N_15384,N_15690);
and U16887 (N_16887,N_15773,N_15668);
or U16888 (N_16888,N_15615,N_15758);
nor U16889 (N_16889,N_15427,N_15682);
nor U16890 (N_16890,N_15595,N_15257);
or U16891 (N_16891,N_15451,N_15415);
xnor U16892 (N_16892,N_15881,N_15139);
and U16893 (N_16893,N_15149,N_15296);
and U16894 (N_16894,N_15659,N_15349);
nand U16895 (N_16895,N_15631,N_15226);
and U16896 (N_16896,N_15383,N_15610);
or U16897 (N_16897,N_15758,N_15221);
xnor U16898 (N_16898,N_15879,N_15245);
xnor U16899 (N_16899,N_15886,N_15556);
or U16900 (N_16900,N_15565,N_15518);
and U16901 (N_16901,N_15353,N_15180);
nand U16902 (N_16902,N_15779,N_15111);
nand U16903 (N_16903,N_15695,N_15996);
nor U16904 (N_16904,N_15447,N_15415);
xnor U16905 (N_16905,N_15633,N_15647);
nand U16906 (N_16906,N_15447,N_15145);
or U16907 (N_16907,N_15246,N_15265);
nor U16908 (N_16908,N_15020,N_15564);
and U16909 (N_16909,N_15182,N_15975);
nand U16910 (N_16910,N_15117,N_15908);
or U16911 (N_16911,N_15621,N_15113);
xor U16912 (N_16912,N_15531,N_15914);
or U16913 (N_16913,N_15886,N_15249);
or U16914 (N_16914,N_15956,N_15870);
or U16915 (N_16915,N_15369,N_15786);
and U16916 (N_16916,N_15138,N_15763);
and U16917 (N_16917,N_15861,N_15746);
and U16918 (N_16918,N_15349,N_15586);
xnor U16919 (N_16919,N_15373,N_15238);
xnor U16920 (N_16920,N_15109,N_15049);
nor U16921 (N_16921,N_15626,N_15245);
or U16922 (N_16922,N_15058,N_15548);
and U16923 (N_16923,N_15161,N_15312);
nor U16924 (N_16924,N_15652,N_15086);
and U16925 (N_16925,N_15906,N_15510);
xnor U16926 (N_16926,N_15769,N_15330);
xnor U16927 (N_16927,N_15449,N_15268);
and U16928 (N_16928,N_15370,N_15574);
and U16929 (N_16929,N_15971,N_15820);
nand U16930 (N_16930,N_15736,N_15339);
nor U16931 (N_16931,N_15562,N_15595);
nor U16932 (N_16932,N_15200,N_15059);
and U16933 (N_16933,N_15924,N_15038);
nand U16934 (N_16934,N_15292,N_15267);
xor U16935 (N_16935,N_15523,N_15788);
or U16936 (N_16936,N_15906,N_15236);
nand U16937 (N_16937,N_15166,N_15809);
nor U16938 (N_16938,N_15412,N_15099);
and U16939 (N_16939,N_15973,N_15856);
and U16940 (N_16940,N_15288,N_15500);
nand U16941 (N_16941,N_15070,N_15646);
or U16942 (N_16942,N_15659,N_15523);
nor U16943 (N_16943,N_15037,N_15428);
and U16944 (N_16944,N_15613,N_15030);
xor U16945 (N_16945,N_15480,N_15676);
nor U16946 (N_16946,N_15696,N_15908);
nor U16947 (N_16947,N_15925,N_15383);
nor U16948 (N_16948,N_15753,N_15426);
and U16949 (N_16949,N_15071,N_15330);
nor U16950 (N_16950,N_15249,N_15696);
and U16951 (N_16951,N_15175,N_15078);
xor U16952 (N_16952,N_15975,N_15539);
xor U16953 (N_16953,N_15110,N_15279);
xnor U16954 (N_16954,N_15672,N_15378);
nand U16955 (N_16955,N_15067,N_15710);
and U16956 (N_16956,N_15753,N_15148);
xnor U16957 (N_16957,N_15253,N_15842);
and U16958 (N_16958,N_15330,N_15062);
nand U16959 (N_16959,N_15083,N_15621);
or U16960 (N_16960,N_15362,N_15772);
and U16961 (N_16961,N_15557,N_15189);
nor U16962 (N_16962,N_15072,N_15577);
and U16963 (N_16963,N_15845,N_15488);
or U16964 (N_16964,N_15765,N_15483);
nor U16965 (N_16965,N_15911,N_15279);
nor U16966 (N_16966,N_15889,N_15044);
nand U16967 (N_16967,N_15935,N_15416);
or U16968 (N_16968,N_15168,N_15487);
nor U16969 (N_16969,N_15012,N_15044);
nor U16970 (N_16970,N_15215,N_15466);
nor U16971 (N_16971,N_15722,N_15352);
and U16972 (N_16972,N_15608,N_15939);
nand U16973 (N_16973,N_15660,N_15916);
nand U16974 (N_16974,N_15514,N_15589);
and U16975 (N_16975,N_15830,N_15044);
xnor U16976 (N_16976,N_15764,N_15477);
xnor U16977 (N_16977,N_15499,N_15179);
nand U16978 (N_16978,N_15987,N_15701);
nor U16979 (N_16979,N_15954,N_15031);
xnor U16980 (N_16980,N_15512,N_15197);
xor U16981 (N_16981,N_15479,N_15521);
nor U16982 (N_16982,N_15970,N_15148);
nor U16983 (N_16983,N_15321,N_15520);
nand U16984 (N_16984,N_15049,N_15033);
and U16985 (N_16985,N_15454,N_15884);
xor U16986 (N_16986,N_15736,N_15627);
and U16987 (N_16987,N_15601,N_15520);
or U16988 (N_16988,N_15004,N_15677);
xnor U16989 (N_16989,N_15371,N_15530);
nand U16990 (N_16990,N_15565,N_15165);
nand U16991 (N_16991,N_15787,N_15217);
nor U16992 (N_16992,N_15088,N_15124);
or U16993 (N_16993,N_15762,N_15085);
nand U16994 (N_16994,N_15757,N_15403);
and U16995 (N_16995,N_15680,N_15062);
nand U16996 (N_16996,N_15672,N_15963);
and U16997 (N_16997,N_15102,N_15907);
or U16998 (N_16998,N_15686,N_15860);
and U16999 (N_16999,N_15031,N_15411);
nor U17000 (N_17000,N_16614,N_16787);
nand U17001 (N_17001,N_16006,N_16689);
and U17002 (N_17002,N_16041,N_16658);
xor U17003 (N_17003,N_16551,N_16494);
nand U17004 (N_17004,N_16742,N_16423);
nor U17005 (N_17005,N_16532,N_16229);
xor U17006 (N_17006,N_16149,N_16996);
or U17007 (N_17007,N_16783,N_16236);
or U17008 (N_17008,N_16831,N_16034);
xnor U17009 (N_17009,N_16398,N_16472);
nor U17010 (N_17010,N_16365,N_16426);
nor U17011 (N_17011,N_16972,N_16453);
nand U17012 (N_17012,N_16240,N_16355);
nor U17013 (N_17013,N_16058,N_16683);
nor U17014 (N_17014,N_16827,N_16456);
nand U17015 (N_17015,N_16161,N_16022);
nand U17016 (N_17016,N_16618,N_16698);
xor U17017 (N_17017,N_16412,N_16239);
nor U17018 (N_17018,N_16293,N_16526);
nor U17019 (N_17019,N_16891,N_16910);
and U17020 (N_17020,N_16476,N_16554);
or U17021 (N_17021,N_16726,N_16748);
and U17022 (N_17022,N_16096,N_16973);
and U17023 (N_17023,N_16755,N_16182);
and U17024 (N_17024,N_16263,N_16319);
and U17025 (N_17025,N_16521,N_16792);
and U17026 (N_17026,N_16789,N_16055);
xor U17027 (N_17027,N_16357,N_16193);
xnor U17028 (N_17028,N_16143,N_16128);
and U17029 (N_17029,N_16611,N_16375);
nand U17030 (N_17030,N_16490,N_16231);
nor U17031 (N_17031,N_16397,N_16807);
or U17032 (N_17032,N_16601,N_16281);
nand U17033 (N_17033,N_16282,N_16926);
or U17034 (N_17034,N_16109,N_16673);
xor U17035 (N_17035,N_16606,N_16038);
nor U17036 (N_17036,N_16104,N_16648);
xor U17037 (N_17037,N_16892,N_16847);
and U17038 (N_17038,N_16978,N_16919);
and U17039 (N_17039,N_16021,N_16353);
nand U17040 (N_17040,N_16334,N_16562);
nand U17041 (N_17041,N_16053,N_16284);
or U17042 (N_17042,N_16155,N_16123);
nor U17043 (N_17043,N_16524,N_16958);
or U17044 (N_17044,N_16001,N_16003);
and U17045 (N_17045,N_16565,N_16546);
nor U17046 (N_17046,N_16424,N_16617);
nand U17047 (N_17047,N_16641,N_16632);
xnor U17048 (N_17048,N_16868,N_16794);
nand U17049 (N_17049,N_16198,N_16124);
nand U17050 (N_17050,N_16216,N_16060);
or U17051 (N_17051,N_16441,N_16206);
xnor U17052 (N_17052,N_16194,N_16429);
nand U17053 (N_17053,N_16406,N_16242);
and U17054 (N_17054,N_16176,N_16695);
nand U17055 (N_17055,N_16802,N_16044);
xor U17056 (N_17056,N_16579,N_16739);
nand U17057 (N_17057,N_16483,N_16099);
and U17058 (N_17058,N_16049,N_16657);
or U17059 (N_17059,N_16960,N_16437);
xnor U17060 (N_17060,N_16866,N_16713);
xor U17061 (N_17061,N_16577,N_16699);
and U17062 (N_17062,N_16414,N_16328);
xnor U17063 (N_17063,N_16697,N_16095);
or U17064 (N_17064,N_16707,N_16090);
nand U17065 (N_17065,N_16955,N_16782);
and U17066 (N_17066,N_16582,N_16300);
and U17067 (N_17067,N_16708,N_16151);
nand U17068 (N_17068,N_16164,N_16363);
xor U17069 (N_17069,N_16788,N_16106);
nand U17070 (N_17070,N_16184,N_16439);
and U17071 (N_17071,N_16549,N_16311);
xor U17072 (N_17072,N_16081,N_16781);
nand U17073 (N_17073,N_16988,N_16816);
nand U17074 (N_17074,N_16047,N_16480);
nor U17075 (N_17075,N_16643,N_16608);
nand U17076 (N_17076,N_16896,N_16421);
or U17077 (N_17077,N_16276,N_16378);
nand U17078 (N_17078,N_16301,N_16612);
nor U17079 (N_17079,N_16759,N_16347);
and U17080 (N_17080,N_16110,N_16032);
or U17081 (N_17081,N_16872,N_16852);
nor U17082 (N_17082,N_16559,N_16993);
or U17083 (N_17083,N_16920,N_16595);
or U17084 (N_17084,N_16323,N_16101);
xnor U17085 (N_17085,N_16909,N_16541);
and U17086 (N_17086,N_16146,N_16189);
and U17087 (N_17087,N_16438,N_16992);
and U17088 (N_17088,N_16083,N_16070);
xor U17089 (N_17089,N_16877,N_16144);
xnor U17090 (N_17090,N_16817,N_16492);
xnor U17091 (N_17091,N_16298,N_16237);
xor U17092 (N_17092,N_16479,N_16934);
or U17093 (N_17093,N_16224,N_16039);
nor U17094 (N_17094,N_16533,N_16043);
or U17095 (N_17095,N_16740,N_16840);
xnor U17096 (N_17096,N_16839,N_16418);
nor U17097 (N_17097,N_16609,N_16289);
or U17098 (N_17098,N_16523,N_16454);
nand U17099 (N_17099,N_16115,N_16979);
xnor U17100 (N_17100,N_16768,N_16359);
xor U17101 (N_17101,N_16766,N_16447);
nor U17102 (N_17102,N_16922,N_16361);
and U17103 (N_17103,N_16091,N_16348);
xnor U17104 (N_17104,N_16837,N_16136);
xnor U17105 (N_17105,N_16159,N_16141);
xor U17106 (N_17106,N_16848,N_16331);
nor U17107 (N_17107,N_16496,N_16858);
and U17108 (N_17108,N_16644,N_16808);
or U17109 (N_17109,N_16202,N_16667);
and U17110 (N_17110,N_16720,N_16269);
nor U17111 (N_17111,N_16989,N_16287);
nor U17112 (N_17112,N_16659,N_16615);
nand U17113 (N_17113,N_16380,N_16525);
or U17114 (N_17114,N_16349,N_16645);
xor U17115 (N_17115,N_16956,N_16649);
xnor U17116 (N_17116,N_16529,N_16628);
nand U17117 (N_17117,N_16168,N_16745);
and U17118 (N_17118,N_16844,N_16717);
xor U17119 (N_17119,N_16514,N_16336);
or U17120 (N_17120,N_16002,N_16320);
or U17121 (N_17121,N_16261,N_16374);
nand U17122 (N_17122,N_16340,N_16025);
nand U17123 (N_17123,N_16431,N_16660);
xnor U17124 (N_17124,N_16828,N_16969);
nor U17125 (N_17125,N_16527,N_16854);
and U17126 (N_17126,N_16100,N_16207);
and U17127 (N_17127,N_16801,N_16586);
xnor U17128 (N_17128,N_16345,N_16493);
nand U17129 (N_17129,N_16581,N_16140);
and U17130 (N_17130,N_16701,N_16381);
or U17131 (N_17131,N_16646,N_16252);
and U17132 (N_17132,N_16329,N_16324);
or U17133 (N_17133,N_16332,N_16052);
nand U17134 (N_17134,N_16898,N_16593);
nand U17135 (N_17135,N_16631,N_16871);
nand U17136 (N_17136,N_16256,N_16571);
nand U17137 (N_17137,N_16846,N_16142);
nor U17138 (N_17138,N_16157,N_16450);
nor U17139 (N_17139,N_16834,N_16440);
nand U17140 (N_17140,N_16260,N_16211);
nand U17141 (N_17141,N_16605,N_16238);
or U17142 (N_17142,N_16602,N_16102);
nor U17143 (N_17143,N_16603,N_16045);
nor U17144 (N_17144,N_16634,N_16026);
xnor U17145 (N_17145,N_16089,N_16566);
xnor U17146 (N_17146,N_16208,N_16983);
xnor U17147 (N_17147,N_16018,N_16997);
or U17148 (N_17148,N_16550,N_16400);
nand U17149 (N_17149,N_16607,N_16675);
or U17150 (N_17150,N_16062,N_16501);
nor U17151 (N_17151,N_16690,N_16432);
and U17152 (N_17152,N_16651,N_16243);
xnor U17153 (N_17153,N_16841,N_16280);
and U17154 (N_17154,N_16448,N_16927);
or U17155 (N_17155,N_16502,N_16405);
nand U17156 (N_17156,N_16384,N_16545);
nand U17157 (N_17157,N_16779,N_16982);
and U17158 (N_17158,N_16196,N_16829);
and U17159 (N_17159,N_16351,N_16767);
and U17160 (N_17160,N_16725,N_16153);
xor U17161 (N_17161,N_16417,N_16823);
xnor U17162 (N_17162,N_16466,N_16272);
or U17163 (N_17163,N_16731,N_16874);
and U17164 (N_17164,N_16761,N_16408);
nand U17165 (N_17165,N_16033,N_16346);
and U17166 (N_17166,N_16171,N_16227);
xor U17167 (N_17167,N_16650,N_16880);
xnor U17168 (N_17168,N_16422,N_16599);
nor U17169 (N_17169,N_16691,N_16360);
and U17170 (N_17170,N_16195,N_16499);
nor U17171 (N_17171,N_16201,N_16127);
and U17172 (N_17172,N_16084,N_16010);
nand U17173 (N_17173,N_16463,N_16553);
nand U17174 (N_17174,N_16247,N_16183);
nor U17175 (N_17175,N_16434,N_16772);
or U17176 (N_17176,N_16040,N_16913);
xnor U17177 (N_17177,N_16968,N_16536);
nand U17178 (N_17178,N_16179,N_16073);
nand U17179 (N_17179,N_16705,N_16976);
and U17180 (N_17180,N_16461,N_16019);
nor U17181 (N_17181,N_16413,N_16322);
nand U17182 (N_17182,N_16174,N_16574);
and U17183 (N_17183,N_16672,N_16160);
and U17184 (N_17184,N_16403,N_16604);
nand U17185 (N_17185,N_16538,N_16662);
nor U17186 (N_17186,N_16824,N_16732);
and U17187 (N_17187,N_16585,N_16966);
and U17188 (N_17188,N_16503,N_16226);
nand U17189 (N_17189,N_16693,N_16539);
xnor U17190 (N_17190,N_16330,N_16275);
nor U17191 (N_17191,N_16763,N_16621);
xnor U17192 (N_17192,N_16152,N_16815);
xor U17193 (N_17193,N_16148,N_16017);
or U17194 (N_17194,N_16244,N_16568);
nand U17195 (N_17195,N_16561,N_16520);
nor U17196 (N_17196,N_16946,N_16914);
xnor U17197 (N_17197,N_16477,N_16303);
nand U17198 (N_17198,N_16271,N_16886);
or U17199 (N_17199,N_16364,N_16046);
xor U17200 (N_17200,N_16462,N_16647);
nor U17201 (N_17201,N_16430,N_16487);
nand U17202 (N_17202,N_16702,N_16354);
nand U17203 (N_17203,N_16669,N_16250);
or U17204 (N_17204,N_16778,N_16812);
and U17205 (N_17205,N_16481,N_16861);
xnor U17206 (N_17206,N_16011,N_16087);
nand U17207 (N_17207,N_16757,N_16257);
and U17208 (N_17208,N_16210,N_16388);
nor U17209 (N_17209,N_16826,N_16212);
nor U17210 (N_17210,N_16995,N_16362);
nand U17211 (N_17211,N_16775,N_16467);
nor U17212 (N_17212,N_16875,N_16939);
and U17213 (N_17213,N_16190,N_16664);
and U17214 (N_17214,N_16930,N_16205);
and U17215 (N_17215,N_16048,N_16556);
xor U17216 (N_17216,N_16843,N_16059);
xor U17217 (N_17217,N_16855,N_16037);
nand U17218 (N_17218,N_16111,N_16679);
nand U17219 (N_17219,N_16396,N_16986);
and U17220 (N_17220,N_16513,N_16508);
nor U17221 (N_17221,N_16416,N_16098);
nor U17222 (N_17222,N_16971,N_16235);
and U17223 (N_17223,N_16548,N_16806);
or U17224 (N_17224,N_16704,N_16825);
and U17225 (N_17225,N_16068,N_16729);
and U17226 (N_17226,N_16984,N_16470);
nand U17227 (N_17227,N_16942,N_16510);
xnor U17228 (N_17228,N_16784,N_16580);
nand U17229 (N_17229,N_16884,N_16786);
or U17230 (N_17230,N_16390,N_16031);
nand U17231 (N_17231,N_16356,N_16093);
nor U17232 (N_17232,N_16627,N_16012);
nand U17233 (N_17233,N_16793,N_16959);
or U17234 (N_17234,N_16655,N_16722);
nor U17235 (N_17235,N_16935,N_16389);
nand U17236 (N_17236,N_16560,N_16718);
nor U17237 (N_17237,N_16150,N_16665);
or U17238 (N_17238,N_16035,N_16445);
or U17239 (N_17239,N_16819,N_16619);
and U17240 (N_17240,N_16915,N_16994);
or U17241 (N_17241,N_16371,N_16684);
nor U17242 (N_17242,N_16485,N_16878);
nand U17243 (N_17243,N_16107,N_16326);
nor U17244 (N_17244,N_16528,N_16741);
or U17245 (N_17245,N_16799,N_16625);
and U17246 (N_17246,N_16482,N_16180);
and U17247 (N_17247,N_16113,N_16377);
and U17248 (N_17248,N_16590,N_16974);
nand U17249 (N_17249,N_16573,N_16004);
or U17250 (N_17250,N_16009,N_16902);
xnor U17251 (N_17251,N_16457,N_16333);
or U17252 (N_17252,N_16682,N_16917);
nand U17253 (N_17253,N_16557,N_16967);
or U17254 (N_17254,N_16126,N_16344);
or U17255 (N_17255,N_16308,N_16167);
nand U17256 (N_17256,N_16760,N_16097);
and U17257 (N_17257,N_16292,N_16255);
xnor U17258 (N_17258,N_16652,N_16187);
and U17259 (N_17259,N_16894,N_16169);
nand U17260 (N_17260,N_16663,N_16596);
and U17261 (N_17261,N_16882,N_16678);
nand U17262 (N_17262,N_16248,N_16680);
nor U17263 (N_17263,N_16616,N_16558);
xor U17264 (N_17264,N_16249,N_16077);
nand U17265 (N_17265,N_16838,N_16177);
xnor U17266 (N_17266,N_16042,N_16399);
nor U17267 (N_17267,N_16088,N_16297);
nand U17268 (N_17268,N_16563,N_16957);
nor U17269 (N_17269,N_16512,N_16259);
and U17270 (N_17270,N_16232,N_16352);
nor U17271 (N_17271,N_16270,N_16449);
nor U17272 (N_17272,N_16137,N_16842);
nor U17273 (N_17273,N_16591,N_16468);
nand U17274 (N_17274,N_16005,N_16488);
or U17275 (N_17275,N_16130,N_16306);
xor U17276 (N_17276,N_16063,N_16370);
or U17277 (N_17277,N_16507,N_16509);
and U17278 (N_17278,N_16519,N_16633);
nand U17279 (N_17279,N_16134,N_16753);
xnor U17280 (N_17280,N_16600,N_16258);
or U17281 (N_17281,N_16085,N_16000);
nand U17282 (N_17282,N_16350,N_16119);
nor U17283 (N_17283,N_16419,N_16762);
nor U17284 (N_17284,N_16908,N_16268);
nor U17285 (N_17285,N_16233,N_16941);
nand U17286 (N_17286,N_16901,N_16204);
and U17287 (N_17287,N_16635,N_16471);
nor U17288 (N_17288,N_16728,N_16575);
xnor U17289 (N_17289,N_16511,N_16221);
xnor U17290 (N_17290,N_16961,N_16544);
nand U17291 (N_17291,N_16309,N_16415);
and U17292 (N_17292,N_16339,N_16670);
nor U17293 (N_17293,N_16687,N_16620);
nor U17294 (N_17294,N_16990,N_16358);
and U17295 (N_17295,N_16810,N_16945);
or U17296 (N_17296,N_16938,N_16727);
nor U17297 (N_17297,N_16870,N_16862);
or U17298 (N_17298,N_16262,N_16069);
nand U17299 (N_17299,N_16342,N_16302);
or U17300 (N_17300,N_16218,N_16064);
xor U17301 (N_17301,N_16923,N_16188);
nand U17302 (N_17302,N_16800,N_16750);
nand U17303 (N_17303,N_16474,N_16335);
and U17304 (N_17304,N_16873,N_16112);
or U17305 (N_17305,N_16899,N_16305);
or U17306 (N_17306,N_16066,N_16131);
xnor U17307 (N_17307,N_16315,N_16776);
nand U17308 (N_17308,N_16500,N_16020);
nor U17309 (N_17309,N_16931,N_16120);
nand U17310 (N_17310,N_16288,N_16746);
or U17311 (N_17311,N_16790,N_16505);
xnor U17312 (N_17312,N_16312,N_16234);
or U17313 (N_17313,N_16598,N_16116);
nor U17314 (N_17314,N_16572,N_16597);
xnor U17315 (N_17315,N_16343,N_16516);
nor U17316 (N_17316,N_16253,N_16953);
nor U17317 (N_17317,N_16949,N_16166);
and U17318 (N_17318,N_16879,N_16444);
nand U17319 (N_17319,N_16264,N_16932);
xnor U17320 (N_17320,N_16830,N_16299);
xor U17321 (N_17321,N_16637,N_16805);
and U17322 (N_17322,N_16464,N_16578);
xor U17323 (N_17323,N_16853,N_16251);
nor U17324 (N_17324,N_16186,N_16962);
nand U17325 (N_17325,N_16950,N_16735);
xnor U17326 (N_17326,N_16576,N_16024);
xnor U17327 (N_17327,N_16747,N_16079);
and U17328 (N_17328,N_16266,N_16197);
nor U17329 (N_17329,N_16715,N_16696);
and U17330 (N_17330,N_16530,N_16008);
nor U17331 (N_17331,N_16537,N_16890);
nor U17332 (N_17332,N_16056,N_16372);
xnor U17333 (N_17333,N_16991,N_16425);
nor U17334 (N_17334,N_16905,N_16642);
or U17335 (N_17335,N_16803,N_16132);
and U17336 (N_17336,N_16451,N_16475);
and U17337 (N_17337,N_16980,N_16952);
xnor U17338 (N_17338,N_16223,N_16283);
nor U17339 (N_17339,N_16987,N_16241);
and U17340 (N_17340,N_16809,N_16749);
or U17341 (N_17341,N_16518,N_16681);
nand U17342 (N_17342,N_16065,N_16495);
or U17343 (N_17343,N_16916,N_16622);
or U17344 (N_17344,N_16859,N_16314);
nand U17345 (N_17345,N_16654,N_16970);
xnor U17346 (N_17346,N_16080,N_16626);
or U17347 (N_17347,N_16692,N_16321);
nand U17348 (N_17348,N_16856,N_16404);
xnor U17349 (N_17349,N_16129,N_16277);
nand U17350 (N_17350,N_16703,N_16737);
xor U17351 (N_17351,N_16118,N_16947);
or U17352 (N_17352,N_16981,N_16821);
xnor U17353 (N_17353,N_16147,N_16677);
nor U17354 (N_17354,N_16057,N_16436);
xor U17355 (N_17355,N_16963,N_16733);
or U17356 (N_17356,N_16156,N_16818);
nand U17357 (N_17357,N_16555,N_16433);
or U17358 (N_17358,N_16610,N_16900);
and U17359 (N_17359,N_16791,N_16588);
or U17360 (N_17360,N_16710,N_16214);
nor U17361 (N_17361,N_16219,N_16700);
and U17362 (N_17362,N_16936,N_16893);
xnor U17363 (N_17363,N_16304,N_16460);
and U17364 (N_17364,N_16086,N_16246);
or U17365 (N_17365,N_16379,N_16163);
or U17366 (N_17366,N_16797,N_16285);
or U17367 (N_17367,N_16613,N_16181);
nand U17368 (N_17368,N_16709,N_16845);
or U17369 (N_17369,N_16676,N_16921);
or U17370 (N_17370,N_16674,N_16016);
and U17371 (N_17371,N_16583,N_16410);
nand U17372 (N_17372,N_16051,N_16316);
xor U17373 (N_17373,N_16473,N_16832);
xor U17374 (N_17374,N_16686,N_16133);
xor U17375 (N_17375,N_16985,N_16220);
and U17376 (N_17376,N_16754,N_16835);
nand U17377 (N_17377,N_16764,N_16883);
nor U17378 (N_17378,N_16145,N_16925);
or U17379 (N_17379,N_16795,N_16724);
nor U17380 (N_17380,N_16567,N_16712);
xnor U17381 (N_17381,N_16318,N_16640);
and U17382 (N_17382,N_16478,N_16999);
and U17383 (N_17383,N_16851,N_16804);
and U17384 (N_17384,N_16706,N_16769);
nor U17385 (N_17385,N_16552,N_16094);
or U17386 (N_17386,N_16564,N_16185);
xnor U17387 (N_17387,N_16369,N_16225);
and U17388 (N_17388,N_16428,N_16023);
xor U17389 (N_17389,N_16814,N_16624);
and U17390 (N_17390,N_16940,N_16903);
xnor U17391 (N_17391,N_16716,N_16907);
xor U17392 (N_17392,N_16267,N_16636);
nand U17393 (N_17393,N_16623,N_16629);
nor U17394 (N_17394,N_16944,N_16833);
nand U17395 (N_17395,N_16217,N_16078);
and U17396 (N_17396,N_16744,N_16569);
or U17397 (N_17397,N_16535,N_16730);
and U17398 (N_17398,N_16376,N_16867);
and U17399 (N_17399,N_16777,N_16443);
nor U17400 (N_17400,N_16489,N_16639);
nor U17401 (N_17401,N_16402,N_16796);
xor U17402 (N_17402,N_16054,N_16050);
xor U17403 (N_17403,N_16459,N_16638);
or U17404 (N_17404,N_16027,N_16072);
xor U17405 (N_17405,N_16173,N_16765);
or U17406 (N_17406,N_16310,N_16743);
nor U17407 (N_17407,N_16469,N_16170);
or U17408 (N_17408,N_16279,N_16911);
xor U17409 (N_17409,N_16121,N_16082);
and U17410 (N_17410,N_16391,N_16209);
nand U17411 (N_17411,N_16685,N_16162);
nand U17412 (N_17412,N_16394,N_16964);
nor U17413 (N_17413,N_16774,N_16547);
and U17414 (N_17414,N_16455,N_16497);
nand U17415 (N_17415,N_16135,N_16076);
nor U17416 (N_17416,N_16138,N_16849);
nand U17417 (N_17417,N_16446,N_16007);
xnor U17418 (N_17418,N_16154,N_16864);
or U17419 (N_17419,N_16028,N_16484);
xor U17420 (N_17420,N_16758,N_16465);
nand U17421 (N_17421,N_16785,N_16714);
and U17422 (N_17422,N_16688,N_16943);
nand U17423 (N_17423,N_16515,N_16367);
nor U17424 (N_17424,N_16965,N_16029);
nor U17425 (N_17425,N_16172,N_16392);
xor U17426 (N_17426,N_16030,N_16036);
nand U17427 (N_17427,N_16881,N_16977);
xnor U17428 (N_17428,N_16387,N_16014);
xnor U17429 (N_17429,N_16230,N_16850);
and U17430 (N_17430,N_16200,N_16103);
nor U17431 (N_17431,N_16570,N_16904);
xor U17432 (N_17432,N_16929,N_16278);
or U17433 (N_17433,N_16504,N_16420);
or U17434 (N_17434,N_16592,N_16383);
nand U17435 (N_17435,N_16286,N_16114);
and U17436 (N_17436,N_16887,N_16906);
nand U17437 (N_17437,N_16307,N_16395);
xor U17438 (N_17438,N_16951,N_16125);
and U17439 (N_17439,N_16452,N_16860);
nor U17440 (N_17440,N_16928,N_16071);
nor U17441 (N_17441,N_16092,N_16671);
xor U17442 (N_17442,N_16015,N_16998);
nand U17443 (N_17443,N_16409,N_16813);
or U17444 (N_17444,N_16175,N_16338);
and U17445 (N_17445,N_16222,N_16857);
nand U17446 (N_17446,N_16393,N_16117);
or U17447 (N_17447,N_16780,N_16427);
nor U17448 (N_17448,N_16245,N_16290);
nand U17449 (N_17449,N_16954,N_16442);
nor U17450 (N_17450,N_16666,N_16254);
and U17451 (N_17451,N_16317,N_16836);
xnor U17452 (N_17452,N_16401,N_16061);
xnor U17453 (N_17453,N_16506,N_16313);
nand U17454 (N_17454,N_16368,N_16458);
xnor U17455 (N_17455,N_16948,N_16542);
nor U17456 (N_17456,N_16594,N_16863);
nand U17457 (N_17457,N_16865,N_16820);
nand U17458 (N_17458,N_16165,N_16752);
nor U17459 (N_17459,N_16719,N_16734);
nor U17460 (N_17460,N_16888,N_16296);
and U17461 (N_17461,N_16178,N_16486);
and U17462 (N_17462,N_16325,N_16668);
xnor U17463 (N_17463,N_16265,N_16215);
nor U17464 (N_17464,N_16918,N_16924);
xor U17465 (N_17465,N_16773,N_16738);
and U17466 (N_17466,N_16411,N_16543);
and U17467 (N_17467,N_16771,N_16937);
nor U17468 (N_17468,N_16721,N_16382);
nor U17469 (N_17469,N_16736,N_16751);
xor U17470 (N_17470,N_16341,N_16897);
xnor U17471 (N_17471,N_16199,N_16491);
nand U17472 (N_17472,N_16584,N_16435);
nand U17473 (N_17473,N_16274,N_16522);
nand U17474 (N_17474,N_16694,N_16661);
xnor U17475 (N_17475,N_16108,N_16013);
or U17476 (N_17476,N_16386,N_16770);
nor U17477 (N_17477,N_16723,N_16074);
and U17478 (N_17478,N_16531,N_16366);
and U17479 (N_17479,N_16822,N_16373);
and U17480 (N_17480,N_16811,N_16407);
or U17481 (N_17481,N_16975,N_16191);
xnor U17482 (N_17482,N_16105,N_16385);
xnor U17483 (N_17483,N_16889,N_16885);
or U17484 (N_17484,N_16139,N_16273);
nand U17485 (N_17485,N_16540,N_16517);
nor U17486 (N_17486,N_16075,N_16295);
nand U17487 (N_17487,N_16912,N_16213);
and U17488 (N_17488,N_16203,N_16933);
nor U17489 (N_17489,N_16756,N_16192);
xnor U17490 (N_17490,N_16587,N_16656);
xor U17491 (N_17491,N_16876,N_16327);
and U17492 (N_17492,N_16337,N_16630);
xnor U17493 (N_17493,N_16291,N_16158);
nand U17494 (N_17494,N_16653,N_16711);
nand U17495 (N_17495,N_16798,N_16589);
or U17496 (N_17496,N_16895,N_16498);
nand U17497 (N_17497,N_16869,N_16067);
nand U17498 (N_17498,N_16122,N_16228);
and U17499 (N_17499,N_16294,N_16534);
or U17500 (N_17500,N_16588,N_16535);
nand U17501 (N_17501,N_16073,N_16814);
xnor U17502 (N_17502,N_16480,N_16870);
xnor U17503 (N_17503,N_16824,N_16203);
xnor U17504 (N_17504,N_16878,N_16833);
nand U17505 (N_17505,N_16871,N_16318);
nor U17506 (N_17506,N_16216,N_16378);
xor U17507 (N_17507,N_16154,N_16914);
xnor U17508 (N_17508,N_16883,N_16673);
xor U17509 (N_17509,N_16959,N_16227);
xor U17510 (N_17510,N_16565,N_16383);
or U17511 (N_17511,N_16266,N_16814);
xor U17512 (N_17512,N_16705,N_16003);
nand U17513 (N_17513,N_16383,N_16547);
nor U17514 (N_17514,N_16055,N_16317);
or U17515 (N_17515,N_16921,N_16493);
nor U17516 (N_17516,N_16157,N_16206);
nand U17517 (N_17517,N_16882,N_16788);
or U17518 (N_17518,N_16997,N_16315);
nor U17519 (N_17519,N_16370,N_16164);
nor U17520 (N_17520,N_16667,N_16170);
xnor U17521 (N_17521,N_16718,N_16413);
nor U17522 (N_17522,N_16840,N_16450);
xor U17523 (N_17523,N_16847,N_16233);
xnor U17524 (N_17524,N_16228,N_16762);
xnor U17525 (N_17525,N_16854,N_16503);
nand U17526 (N_17526,N_16568,N_16517);
nor U17527 (N_17527,N_16464,N_16524);
or U17528 (N_17528,N_16236,N_16566);
nand U17529 (N_17529,N_16545,N_16933);
xor U17530 (N_17530,N_16941,N_16930);
and U17531 (N_17531,N_16824,N_16196);
or U17532 (N_17532,N_16213,N_16920);
or U17533 (N_17533,N_16320,N_16112);
xnor U17534 (N_17534,N_16627,N_16454);
nor U17535 (N_17535,N_16527,N_16743);
nand U17536 (N_17536,N_16117,N_16455);
nor U17537 (N_17537,N_16507,N_16742);
nor U17538 (N_17538,N_16548,N_16240);
and U17539 (N_17539,N_16563,N_16605);
xnor U17540 (N_17540,N_16794,N_16370);
nor U17541 (N_17541,N_16297,N_16387);
or U17542 (N_17542,N_16766,N_16035);
nor U17543 (N_17543,N_16481,N_16194);
and U17544 (N_17544,N_16872,N_16053);
nor U17545 (N_17545,N_16370,N_16811);
or U17546 (N_17546,N_16060,N_16680);
and U17547 (N_17547,N_16027,N_16536);
and U17548 (N_17548,N_16873,N_16991);
or U17549 (N_17549,N_16827,N_16670);
nor U17550 (N_17550,N_16162,N_16712);
xnor U17551 (N_17551,N_16035,N_16648);
xor U17552 (N_17552,N_16387,N_16391);
and U17553 (N_17553,N_16907,N_16310);
and U17554 (N_17554,N_16578,N_16266);
nand U17555 (N_17555,N_16880,N_16022);
xor U17556 (N_17556,N_16613,N_16311);
and U17557 (N_17557,N_16803,N_16507);
or U17558 (N_17558,N_16366,N_16637);
nand U17559 (N_17559,N_16477,N_16606);
nor U17560 (N_17560,N_16081,N_16359);
xnor U17561 (N_17561,N_16883,N_16683);
xor U17562 (N_17562,N_16960,N_16525);
nand U17563 (N_17563,N_16393,N_16722);
or U17564 (N_17564,N_16475,N_16621);
or U17565 (N_17565,N_16481,N_16620);
and U17566 (N_17566,N_16554,N_16567);
and U17567 (N_17567,N_16290,N_16996);
nor U17568 (N_17568,N_16363,N_16347);
and U17569 (N_17569,N_16685,N_16290);
nor U17570 (N_17570,N_16397,N_16231);
and U17571 (N_17571,N_16207,N_16676);
or U17572 (N_17572,N_16936,N_16151);
xnor U17573 (N_17573,N_16903,N_16914);
nor U17574 (N_17574,N_16529,N_16773);
nand U17575 (N_17575,N_16261,N_16712);
or U17576 (N_17576,N_16303,N_16214);
xnor U17577 (N_17577,N_16980,N_16439);
xnor U17578 (N_17578,N_16990,N_16762);
and U17579 (N_17579,N_16085,N_16552);
or U17580 (N_17580,N_16158,N_16181);
and U17581 (N_17581,N_16728,N_16227);
or U17582 (N_17582,N_16164,N_16530);
xor U17583 (N_17583,N_16501,N_16966);
xor U17584 (N_17584,N_16063,N_16572);
xnor U17585 (N_17585,N_16785,N_16018);
or U17586 (N_17586,N_16642,N_16574);
nand U17587 (N_17587,N_16798,N_16150);
nor U17588 (N_17588,N_16965,N_16607);
nor U17589 (N_17589,N_16509,N_16809);
nor U17590 (N_17590,N_16019,N_16399);
nor U17591 (N_17591,N_16918,N_16780);
or U17592 (N_17592,N_16413,N_16488);
nand U17593 (N_17593,N_16801,N_16722);
nand U17594 (N_17594,N_16518,N_16991);
nand U17595 (N_17595,N_16786,N_16391);
or U17596 (N_17596,N_16859,N_16709);
nor U17597 (N_17597,N_16761,N_16805);
nand U17598 (N_17598,N_16789,N_16873);
xnor U17599 (N_17599,N_16447,N_16801);
or U17600 (N_17600,N_16562,N_16194);
xnor U17601 (N_17601,N_16867,N_16361);
or U17602 (N_17602,N_16910,N_16622);
nor U17603 (N_17603,N_16535,N_16621);
and U17604 (N_17604,N_16602,N_16027);
and U17605 (N_17605,N_16741,N_16974);
nor U17606 (N_17606,N_16745,N_16979);
nor U17607 (N_17607,N_16735,N_16780);
nor U17608 (N_17608,N_16808,N_16190);
xor U17609 (N_17609,N_16788,N_16152);
nand U17610 (N_17610,N_16420,N_16928);
nand U17611 (N_17611,N_16761,N_16332);
and U17612 (N_17612,N_16483,N_16307);
xnor U17613 (N_17613,N_16526,N_16368);
xnor U17614 (N_17614,N_16965,N_16479);
or U17615 (N_17615,N_16511,N_16809);
and U17616 (N_17616,N_16607,N_16645);
nor U17617 (N_17617,N_16233,N_16100);
or U17618 (N_17618,N_16268,N_16558);
nor U17619 (N_17619,N_16904,N_16542);
nor U17620 (N_17620,N_16198,N_16809);
nor U17621 (N_17621,N_16040,N_16085);
and U17622 (N_17622,N_16863,N_16826);
nor U17623 (N_17623,N_16890,N_16798);
or U17624 (N_17624,N_16143,N_16970);
or U17625 (N_17625,N_16713,N_16071);
xor U17626 (N_17626,N_16983,N_16164);
nand U17627 (N_17627,N_16178,N_16078);
nor U17628 (N_17628,N_16447,N_16138);
nor U17629 (N_17629,N_16646,N_16618);
xor U17630 (N_17630,N_16342,N_16566);
nor U17631 (N_17631,N_16240,N_16411);
or U17632 (N_17632,N_16761,N_16765);
xor U17633 (N_17633,N_16802,N_16436);
nor U17634 (N_17634,N_16668,N_16339);
nor U17635 (N_17635,N_16620,N_16362);
xor U17636 (N_17636,N_16828,N_16403);
nand U17637 (N_17637,N_16881,N_16869);
xor U17638 (N_17638,N_16263,N_16633);
or U17639 (N_17639,N_16330,N_16593);
and U17640 (N_17640,N_16091,N_16448);
nor U17641 (N_17641,N_16277,N_16806);
or U17642 (N_17642,N_16713,N_16273);
and U17643 (N_17643,N_16547,N_16203);
xor U17644 (N_17644,N_16860,N_16360);
or U17645 (N_17645,N_16683,N_16940);
nor U17646 (N_17646,N_16453,N_16497);
nand U17647 (N_17647,N_16788,N_16984);
nor U17648 (N_17648,N_16023,N_16072);
nand U17649 (N_17649,N_16600,N_16693);
and U17650 (N_17650,N_16152,N_16432);
nand U17651 (N_17651,N_16910,N_16028);
xnor U17652 (N_17652,N_16026,N_16118);
nand U17653 (N_17653,N_16049,N_16892);
nor U17654 (N_17654,N_16216,N_16588);
xnor U17655 (N_17655,N_16600,N_16356);
nand U17656 (N_17656,N_16622,N_16797);
nor U17657 (N_17657,N_16218,N_16936);
and U17658 (N_17658,N_16368,N_16589);
nor U17659 (N_17659,N_16283,N_16973);
nor U17660 (N_17660,N_16685,N_16338);
xnor U17661 (N_17661,N_16459,N_16912);
or U17662 (N_17662,N_16591,N_16180);
or U17663 (N_17663,N_16585,N_16735);
xnor U17664 (N_17664,N_16605,N_16210);
xor U17665 (N_17665,N_16311,N_16124);
xnor U17666 (N_17666,N_16265,N_16820);
nor U17667 (N_17667,N_16829,N_16915);
xnor U17668 (N_17668,N_16396,N_16186);
and U17669 (N_17669,N_16822,N_16297);
or U17670 (N_17670,N_16187,N_16060);
nor U17671 (N_17671,N_16518,N_16830);
or U17672 (N_17672,N_16847,N_16948);
nor U17673 (N_17673,N_16094,N_16158);
nand U17674 (N_17674,N_16223,N_16147);
or U17675 (N_17675,N_16128,N_16382);
or U17676 (N_17676,N_16199,N_16276);
and U17677 (N_17677,N_16941,N_16798);
xor U17678 (N_17678,N_16730,N_16136);
nand U17679 (N_17679,N_16873,N_16540);
nand U17680 (N_17680,N_16560,N_16703);
nand U17681 (N_17681,N_16753,N_16808);
and U17682 (N_17682,N_16098,N_16178);
and U17683 (N_17683,N_16478,N_16415);
nand U17684 (N_17684,N_16200,N_16692);
xor U17685 (N_17685,N_16782,N_16656);
or U17686 (N_17686,N_16269,N_16037);
nand U17687 (N_17687,N_16175,N_16885);
xor U17688 (N_17688,N_16406,N_16771);
or U17689 (N_17689,N_16046,N_16983);
and U17690 (N_17690,N_16781,N_16349);
nand U17691 (N_17691,N_16730,N_16124);
nor U17692 (N_17692,N_16256,N_16309);
nor U17693 (N_17693,N_16212,N_16701);
xnor U17694 (N_17694,N_16163,N_16289);
and U17695 (N_17695,N_16194,N_16563);
nand U17696 (N_17696,N_16297,N_16256);
or U17697 (N_17697,N_16988,N_16652);
nand U17698 (N_17698,N_16394,N_16670);
or U17699 (N_17699,N_16345,N_16620);
and U17700 (N_17700,N_16078,N_16050);
xnor U17701 (N_17701,N_16488,N_16490);
nand U17702 (N_17702,N_16039,N_16477);
or U17703 (N_17703,N_16161,N_16277);
nand U17704 (N_17704,N_16474,N_16084);
nand U17705 (N_17705,N_16843,N_16733);
nand U17706 (N_17706,N_16146,N_16240);
and U17707 (N_17707,N_16387,N_16639);
and U17708 (N_17708,N_16111,N_16611);
nor U17709 (N_17709,N_16912,N_16295);
xnor U17710 (N_17710,N_16950,N_16707);
or U17711 (N_17711,N_16839,N_16187);
or U17712 (N_17712,N_16056,N_16319);
xnor U17713 (N_17713,N_16358,N_16475);
xnor U17714 (N_17714,N_16400,N_16001);
nand U17715 (N_17715,N_16377,N_16666);
nand U17716 (N_17716,N_16083,N_16295);
xor U17717 (N_17717,N_16827,N_16050);
xor U17718 (N_17718,N_16013,N_16445);
or U17719 (N_17719,N_16823,N_16361);
nand U17720 (N_17720,N_16778,N_16566);
nand U17721 (N_17721,N_16601,N_16623);
and U17722 (N_17722,N_16303,N_16404);
nor U17723 (N_17723,N_16816,N_16211);
or U17724 (N_17724,N_16159,N_16300);
xor U17725 (N_17725,N_16760,N_16976);
nand U17726 (N_17726,N_16492,N_16761);
or U17727 (N_17727,N_16587,N_16335);
and U17728 (N_17728,N_16360,N_16068);
nor U17729 (N_17729,N_16932,N_16205);
nand U17730 (N_17730,N_16964,N_16532);
and U17731 (N_17731,N_16558,N_16135);
xnor U17732 (N_17732,N_16876,N_16307);
or U17733 (N_17733,N_16490,N_16856);
nor U17734 (N_17734,N_16250,N_16921);
and U17735 (N_17735,N_16121,N_16178);
nor U17736 (N_17736,N_16861,N_16789);
xor U17737 (N_17737,N_16526,N_16484);
and U17738 (N_17738,N_16465,N_16150);
and U17739 (N_17739,N_16618,N_16238);
nor U17740 (N_17740,N_16459,N_16615);
or U17741 (N_17741,N_16077,N_16113);
nor U17742 (N_17742,N_16768,N_16760);
and U17743 (N_17743,N_16694,N_16718);
xnor U17744 (N_17744,N_16161,N_16576);
nand U17745 (N_17745,N_16985,N_16755);
nor U17746 (N_17746,N_16353,N_16606);
or U17747 (N_17747,N_16538,N_16791);
xor U17748 (N_17748,N_16565,N_16589);
nor U17749 (N_17749,N_16431,N_16783);
nor U17750 (N_17750,N_16481,N_16723);
and U17751 (N_17751,N_16557,N_16932);
or U17752 (N_17752,N_16532,N_16464);
or U17753 (N_17753,N_16007,N_16723);
nand U17754 (N_17754,N_16423,N_16897);
nand U17755 (N_17755,N_16320,N_16660);
and U17756 (N_17756,N_16965,N_16293);
nand U17757 (N_17757,N_16069,N_16581);
xor U17758 (N_17758,N_16984,N_16475);
nand U17759 (N_17759,N_16088,N_16070);
xor U17760 (N_17760,N_16096,N_16953);
and U17761 (N_17761,N_16621,N_16772);
and U17762 (N_17762,N_16964,N_16103);
and U17763 (N_17763,N_16657,N_16140);
and U17764 (N_17764,N_16454,N_16595);
and U17765 (N_17765,N_16104,N_16812);
or U17766 (N_17766,N_16697,N_16917);
or U17767 (N_17767,N_16328,N_16865);
and U17768 (N_17768,N_16903,N_16135);
nor U17769 (N_17769,N_16604,N_16415);
or U17770 (N_17770,N_16326,N_16598);
or U17771 (N_17771,N_16336,N_16998);
or U17772 (N_17772,N_16857,N_16703);
nand U17773 (N_17773,N_16515,N_16443);
nand U17774 (N_17774,N_16386,N_16627);
nor U17775 (N_17775,N_16919,N_16015);
or U17776 (N_17776,N_16071,N_16602);
or U17777 (N_17777,N_16173,N_16940);
nand U17778 (N_17778,N_16721,N_16272);
nand U17779 (N_17779,N_16252,N_16526);
and U17780 (N_17780,N_16041,N_16801);
xor U17781 (N_17781,N_16409,N_16314);
and U17782 (N_17782,N_16575,N_16646);
nor U17783 (N_17783,N_16010,N_16296);
or U17784 (N_17784,N_16676,N_16870);
nand U17785 (N_17785,N_16417,N_16112);
and U17786 (N_17786,N_16679,N_16615);
nand U17787 (N_17787,N_16152,N_16208);
nor U17788 (N_17788,N_16272,N_16808);
xor U17789 (N_17789,N_16351,N_16842);
nand U17790 (N_17790,N_16049,N_16500);
and U17791 (N_17791,N_16164,N_16536);
or U17792 (N_17792,N_16853,N_16056);
nand U17793 (N_17793,N_16123,N_16609);
and U17794 (N_17794,N_16674,N_16822);
nor U17795 (N_17795,N_16419,N_16820);
nand U17796 (N_17796,N_16877,N_16003);
or U17797 (N_17797,N_16623,N_16599);
nor U17798 (N_17798,N_16912,N_16547);
and U17799 (N_17799,N_16046,N_16146);
xnor U17800 (N_17800,N_16838,N_16405);
or U17801 (N_17801,N_16251,N_16143);
nand U17802 (N_17802,N_16184,N_16097);
nand U17803 (N_17803,N_16131,N_16231);
and U17804 (N_17804,N_16003,N_16731);
xor U17805 (N_17805,N_16562,N_16892);
nand U17806 (N_17806,N_16835,N_16139);
nand U17807 (N_17807,N_16899,N_16214);
nand U17808 (N_17808,N_16755,N_16650);
nand U17809 (N_17809,N_16941,N_16291);
or U17810 (N_17810,N_16412,N_16570);
xor U17811 (N_17811,N_16220,N_16982);
xnor U17812 (N_17812,N_16475,N_16057);
or U17813 (N_17813,N_16450,N_16292);
nand U17814 (N_17814,N_16219,N_16824);
and U17815 (N_17815,N_16580,N_16788);
and U17816 (N_17816,N_16079,N_16528);
or U17817 (N_17817,N_16240,N_16119);
and U17818 (N_17818,N_16370,N_16987);
nor U17819 (N_17819,N_16307,N_16221);
nor U17820 (N_17820,N_16733,N_16134);
nor U17821 (N_17821,N_16573,N_16505);
xnor U17822 (N_17822,N_16465,N_16496);
nand U17823 (N_17823,N_16400,N_16506);
nand U17824 (N_17824,N_16619,N_16521);
xor U17825 (N_17825,N_16392,N_16542);
nand U17826 (N_17826,N_16938,N_16693);
xnor U17827 (N_17827,N_16246,N_16932);
xor U17828 (N_17828,N_16417,N_16846);
nor U17829 (N_17829,N_16012,N_16409);
nand U17830 (N_17830,N_16424,N_16448);
and U17831 (N_17831,N_16274,N_16131);
or U17832 (N_17832,N_16189,N_16317);
xor U17833 (N_17833,N_16330,N_16506);
nand U17834 (N_17834,N_16428,N_16057);
nor U17835 (N_17835,N_16543,N_16805);
nand U17836 (N_17836,N_16790,N_16716);
xnor U17837 (N_17837,N_16972,N_16293);
nand U17838 (N_17838,N_16032,N_16440);
xor U17839 (N_17839,N_16770,N_16926);
xor U17840 (N_17840,N_16359,N_16538);
and U17841 (N_17841,N_16666,N_16639);
and U17842 (N_17842,N_16749,N_16881);
nor U17843 (N_17843,N_16383,N_16293);
nor U17844 (N_17844,N_16575,N_16788);
and U17845 (N_17845,N_16793,N_16651);
nor U17846 (N_17846,N_16212,N_16382);
nor U17847 (N_17847,N_16555,N_16908);
nor U17848 (N_17848,N_16174,N_16766);
nand U17849 (N_17849,N_16713,N_16487);
or U17850 (N_17850,N_16949,N_16896);
nor U17851 (N_17851,N_16221,N_16226);
nor U17852 (N_17852,N_16249,N_16846);
or U17853 (N_17853,N_16601,N_16545);
xor U17854 (N_17854,N_16503,N_16758);
or U17855 (N_17855,N_16048,N_16123);
and U17856 (N_17856,N_16126,N_16090);
or U17857 (N_17857,N_16688,N_16992);
xor U17858 (N_17858,N_16824,N_16589);
or U17859 (N_17859,N_16697,N_16401);
xnor U17860 (N_17860,N_16448,N_16005);
nor U17861 (N_17861,N_16024,N_16399);
or U17862 (N_17862,N_16083,N_16335);
and U17863 (N_17863,N_16487,N_16681);
or U17864 (N_17864,N_16244,N_16302);
nand U17865 (N_17865,N_16210,N_16632);
xnor U17866 (N_17866,N_16068,N_16728);
and U17867 (N_17867,N_16928,N_16183);
nor U17868 (N_17868,N_16747,N_16601);
nor U17869 (N_17869,N_16954,N_16976);
nor U17870 (N_17870,N_16980,N_16641);
xnor U17871 (N_17871,N_16657,N_16906);
or U17872 (N_17872,N_16777,N_16742);
nand U17873 (N_17873,N_16888,N_16500);
or U17874 (N_17874,N_16994,N_16162);
xor U17875 (N_17875,N_16139,N_16239);
and U17876 (N_17876,N_16367,N_16784);
xor U17877 (N_17877,N_16943,N_16410);
xor U17878 (N_17878,N_16737,N_16994);
nand U17879 (N_17879,N_16963,N_16812);
xnor U17880 (N_17880,N_16722,N_16273);
nor U17881 (N_17881,N_16738,N_16794);
or U17882 (N_17882,N_16347,N_16470);
or U17883 (N_17883,N_16857,N_16476);
nor U17884 (N_17884,N_16931,N_16698);
and U17885 (N_17885,N_16260,N_16476);
and U17886 (N_17886,N_16509,N_16675);
xnor U17887 (N_17887,N_16039,N_16155);
and U17888 (N_17888,N_16022,N_16705);
nor U17889 (N_17889,N_16765,N_16366);
or U17890 (N_17890,N_16545,N_16694);
xnor U17891 (N_17891,N_16180,N_16789);
xor U17892 (N_17892,N_16962,N_16152);
nand U17893 (N_17893,N_16316,N_16201);
and U17894 (N_17894,N_16720,N_16575);
and U17895 (N_17895,N_16305,N_16673);
nor U17896 (N_17896,N_16214,N_16618);
nor U17897 (N_17897,N_16969,N_16726);
and U17898 (N_17898,N_16657,N_16370);
xnor U17899 (N_17899,N_16611,N_16201);
nand U17900 (N_17900,N_16006,N_16853);
nor U17901 (N_17901,N_16857,N_16716);
xor U17902 (N_17902,N_16887,N_16537);
nand U17903 (N_17903,N_16553,N_16879);
xor U17904 (N_17904,N_16394,N_16140);
nand U17905 (N_17905,N_16780,N_16720);
or U17906 (N_17906,N_16081,N_16654);
and U17907 (N_17907,N_16677,N_16590);
or U17908 (N_17908,N_16401,N_16142);
or U17909 (N_17909,N_16437,N_16862);
nor U17910 (N_17910,N_16986,N_16150);
and U17911 (N_17911,N_16145,N_16797);
and U17912 (N_17912,N_16749,N_16486);
xnor U17913 (N_17913,N_16125,N_16290);
xnor U17914 (N_17914,N_16036,N_16701);
nor U17915 (N_17915,N_16667,N_16759);
nor U17916 (N_17916,N_16603,N_16043);
xnor U17917 (N_17917,N_16904,N_16948);
nor U17918 (N_17918,N_16942,N_16098);
nand U17919 (N_17919,N_16356,N_16026);
nor U17920 (N_17920,N_16463,N_16879);
and U17921 (N_17921,N_16410,N_16721);
nor U17922 (N_17922,N_16835,N_16863);
or U17923 (N_17923,N_16894,N_16158);
nand U17924 (N_17924,N_16782,N_16658);
or U17925 (N_17925,N_16730,N_16117);
or U17926 (N_17926,N_16041,N_16012);
or U17927 (N_17927,N_16045,N_16413);
xor U17928 (N_17928,N_16189,N_16119);
nand U17929 (N_17929,N_16384,N_16037);
nand U17930 (N_17930,N_16936,N_16258);
and U17931 (N_17931,N_16944,N_16375);
xor U17932 (N_17932,N_16213,N_16337);
or U17933 (N_17933,N_16674,N_16777);
nand U17934 (N_17934,N_16553,N_16139);
and U17935 (N_17935,N_16768,N_16291);
xor U17936 (N_17936,N_16965,N_16816);
and U17937 (N_17937,N_16251,N_16090);
or U17938 (N_17938,N_16186,N_16518);
or U17939 (N_17939,N_16519,N_16824);
or U17940 (N_17940,N_16254,N_16342);
nor U17941 (N_17941,N_16763,N_16087);
nor U17942 (N_17942,N_16593,N_16533);
nor U17943 (N_17943,N_16545,N_16036);
or U17944 (N_17944,N_16468,N_16340);
nand U17945 (N_17945,N_16138,N_16857);
nand U17946 (N_17946,N_16175,N_16609);
xnor U17947 (N_17947,N_16870,N_16080);
xnor U17948 (N_17948,N_16886,N_16049);
nor U17949 (N_17949,N_16338,N_16208);
nor U17950 (N_17950,N_16413,N_16077);
or U17951 (N_17951,N_16192,N_16224);
and U17952 (N_17952,N_16598,N_16673);
or U17953 (N_17953,N_16279,N_16811);
and U17954 (N_17954,N_16729,N_16120);
xnor U17955 (N_17955,N_16372,N_16516);
nand U17956 (N_17956,N_16251,N_16478);
or U17957 (N_17957,N_16930,N_16676);
nand U17958 (N_17958,N_16214,N_16582);
or U17959 (N_17959,N_16174,N_16081);
and U17960 (N_17960,N_16136,N_16530);
and U17961 (N_17961,N_16220,N_16069);
nand U17962 (N_17962,N_16126,N_16846);
nand U17963 (N_17963,N_16955,N_16571);
xnor U17964 (N_17964,N_16674,N_16998);
or U17965 (N_17965,N_16287,N_16758);
nand U17966 (N_17966,N_16082,N_16615);
xnor U17967 (N_17967,N_16482,N_16785);
nand U17968 (N_17968,N_16491,N_16967);
and U17969 (N_17969,N_16885,N_16794);
nor U17970 (N_17970,N_16656,N_16416);
and U17971 (N_17971,N_16131,N_16840);
and U17972 (N_17972,N_16134,N_16220);
and U17973 (N_17973,N_16994,N_16215);
xnor U17974 (N_17974,N_16535,N_16305);
and U17975 (N_17975,N_16545,N_16284);
nor U17976 (N_17976,N_16459,N_16026);
or U17977 (N_17977,N_16407,N_16905);
nor U17978 (N_17978,N_16252,N_16299);
nor U17979 (N_17979,N_16353,N_16455);
and U17980 (N_17980,N_16667,N_16694);
nor U17981 (N_17981,N_16747,N_16439);
nor U17982 (N_17982,N_16809,N_16674);
nor U17983 (N_17983,N_16024,N_16359);
and U17984 (N_17984,N_16298,N_16418);
or U17985 (N_17985,N_16086,N_16785);
nand U17986 (N_17986,N_16218,N_16861);
nor U17987 (N_17987,N_16726,N_16001);
nand U17988 (N_17988,N_16623,N_16540);
nor U17989 (N_17989,N_16270,N_16269);
nand U17990 (N_17990,N_16471,N_16192);
xnor U17991 (N_17991,N_16325,N_16690);
and U17992 (N_17992,N_16245,N_16405);
nor U17993 (N_17993,N_16218,N_16876);
or U17994 (N_17994,N_16406,N_16230);
or U17995 (N_17995,N_16232,N_16481);
nand U17996 (N_17996,N_16199,N_16632);
xor U17997 (N_17997,N_16961,N_16879);
or U17998 (N_17998,N_16370,N_16749);
xor U17999 (N_17999,N_16956,N_16643);
or U18000 (N_18000,N_17795,N_17418);
nand U18001 (N_18001,N_17267,N_17737);
nand U18002 (N_18002,N_17659,N_17598);
xnor U18003 (N_18003,N_17024,N_17180);
or U18004 (N_18004,N_17684,N_17751);
xor U18005 (N_18005,N_17389,N_17981);
and U18006 (N_18006,N_17170,N_17300);
xor U18007 (N_18007,N_17029,N_17532);
or U18008 (N_18008,N_17668,N_17816);
or U18009 (N_18009,N_17345,N_17327);
xor U18010 (N_18010,N_17958,N_17604);
xor U18011 (N_18011,N_17133,N_17447);
and U18012 (N_18012,N_17768,N_17815);
and U18013 (N_18013,N_17543,N_17064);
xor U18014 (N_18014,N_17434,N_17211);
nor U18015 (N_18015,N_17017,N_17626);
nand U18016 (N_18016,N_17836,N_17929);
and U18017 (N_18017,N_17946,N_17335);
nor U18018 (N_18018,N_17473,N_17496);
nand U18019 (N_18019,N_17182,N_17476);
or U18020 (N_18020,N_17558,N_17348);
nor U18021 (N_18021,N_17288,N_17315);
xnor U18022 (N_18022,N_17819,N_17384);
xor U18023 (N_18023,N_17743,N_17408);
and U18024 (N_18024,N_17048,N_17678);
and U18025 (N_18025,N_17577,N_17665);
nand U18026 (N_18026,N_17534,N_17968);
and U18027 (N_18027,N_17754,N_17618);
or U18028 (N_18028,N_17468,N_17154);
xnor U18029 (N_18029,N_17655,N_17038);
and U18030 (N_18030,N_17292,N_17372);
xor U18031 (N_18031,N_17892,N_17999);
and U18032 (N_18032,N_17583,N_17144);
or U18033 (N_18033,N_17673,N_17839);
or U18034 (N_18034,N_17564,N_17756);
nor U18035 (N_18035,N_17371,N_17844);
nand U18036 (N_18036,N_17205,N_17251);
nand U18037 (N_18037,N_17685,N_17068);
or U18038 (N_18038,N_17420,N_17190);
nand U18039 (N_18039,N_17824,N_17651);
and U18040 (N_18040,N_17452,N_17414);
nor U18041 (N_18041,N_17863,N_17099);
nand U18042 (N_18042,N_17279,N_17118);
xor U18043 (N_18043,N_17823,N_17439);
nor U18044 (N_18044,N_17570,N_17609);
and U18045 (N_18045,N_17898,N_17601);
nand U18046 (N_18046,N_17882,N_17484);
xnor U18047 (N_18047,N_17472,N_17977);
nand U18048 (N_18048,N_17829,N_17429);
nand U18049 (N_18049,N_17368,N_17074);
nand U18050 (N_18050,N_17198,N_17639);
and U18051 (N_18051,N_17049,N_17831);
and U18052 (N_18052,N_17440,N_17835);
nand U18053 (N_18053,N_17553,N_17615);
nor U18054 (N_18054,N_17683,N_17840);
or U18055 (N_18055,N_17467,N_17041);
nand U18056 (N_18056,N_17766,N_17202);
xor U18057 (N_18057,N_17719,N_17297);
nand U18058 (N_18058,N_17638,N_17812);
xor U18059 (N_18059,N_17291,N_17217);
xor U18060 (N_18060,N_17309,N_17396);
or U18061 (N_18061,N_17722,N_17358);
xor U18062 (N_18062,N_17456,N_17713);
nand U18063 (N_18063,N_17301,N_17088);
and U18064 (N_18064,N_17866,N_17505);
nand U18065 (N_18065,N_17984,N_17117);
nand U18066 (N_18066,N_17031,N_17412);
nor U18067 (N_18067,N_17983,N_17256);
or U18068 (N_18068,N_17858,N_17216);
xnor U18069 (N_18069,N_17919,N_17698);
nor U18070 (N_18070,N_17725,N_17193);
nand U18071 (N_18071,N_17243,N_17969);
nand U18072 (N_18072,N_17654,N_17524);
and U18073 (N_18073,N_17895,N_17822);
or U18074 (N_18074,N_17040,N_17612);
nor U18075 (N_18075,N_17717,N_17623);
and U18076 (N_18076,N_17188,N_17443);
nand U18077 (N_18077,N_17788,N_17540);
or U18078 (N_18078,N_17887,N_17421);
and U18079 (N_18079,N_17093,N_17430);
xnor U18080 (N_18080,N_17491,N_17886);
or U18081 (N_18081,N_17156,N_17985);
or U18082 (N_18082,N_17407,N_17149);
or U18083 (N_18083,N_17060,N_17459);
nor U18084 (N_18084,N_17030,N_17463);
and U18085 (N_18085,N_17912,N_17298);
or U18086 (N_18086,N_17095,N_17584);
or U18087 (N_18087,N_17246,N_17232);
nor U18088 (N_18088,N_17356,N_17383);
or U18089 (N_18089,N_17634,N_17566);
nand U18090 (N_18090,N_17089,N_17973);
and U18091 (N_18091,N_17446,N_17571);
nand U18092 (N_18092,N_17970,N_17747);
nor U18093 (N_18093,N_17954,N_17873);
and U18094 (N_18094,N_17228,N_17167);
nor U18095 (N_18095,N_17411,N_17113);
nand U18096 (N_18096,N_17672,N_17303);
xnor U18097 (N_18097,N_17793,N_17735);
nor U18098 (N_18098,N_17141,N_17019);
or U18099 (N_18099,N_17640,N_17596);
xnor U18100 (N_18100,N_17227,N_17398);
nand U18101 (N_18101,N_17575,N_17902);
nor U18102 (N_18102,N_17096,N_17478);
or U18103 (N_18103,N_17481,N_17535);
xnor U18104 (N_18104,N_17953,N_17022);
or U18105 (N_18105,N_17004,N_17294);
nand U18106 (N_18106,N_17830,N_17888);
and U18107 (N_18107,N_17183,N_17350);
xor U18108 (N_18108,N_17857,N_17222);
nor U18109 (N_18109,N_17842,N_17001);
nand U18110 (N_18110,N_17045,N_17950);
nand U18111 (N_18111,N_17242,N_17197);
or U18112 (N_18112,N_17426,N_17894);
xnor U18113 (N_18113,N_17807,N_17305);
xor U18114 (N_18114,N_17871,N_17633);
xnor U18115 (N_18115,N_17774,N_17081);
xor U18116 (N_18116,N_17400,N_17192);
xnor U18117 (N_18117,N_17619,N_17658);
and U18118 (N_18118,N_17903,N_17367);
xor U18119 (N_18119,N_17287,N_17313);
nor U18120 (N_18120,N_17280,N_17083);
nor U18121 (N_18121,N_17401,N_17957);
nor U18122 (N_18122,N_17622,N_17994);
and U18123 (N_18123,N_17181,N_17206);
xor U18124 (N_18124,N_17416,N_17550);
xnor U18125 (N_18125,N_17111,N_17592);
nor U18126 (N_18126,N_17843,N_17562);
nand U18127 (N_18127,N_17506,N_17925);
nand U18128 (N_18128,N_17996,N_17764);
xnor U18129 (N_18129,N_17731,N_17784);
nor U18130 (N_18130,N_17585,N_17054);
or U18131 (N_18131,N_17589,N_17938);
nor U18132 (N_18132,N_17509,N_17299);
and U18133 (N_18133,N_17779,N_17025);
nand U18134 (N_18134,N_17475,N_17670);
and U18135 (N_18135,N_17492,N_17131);
and U18136 (N_18136,N_17771,N_17179);
xor U18137 (N_18137,N_17091,N_17221);
or U18138 (N_18138,N_17399,N_17801);
or U18139 (N_18139,N_17069,N_17600);
nand U18140 (N_18140,N_17811,N_17745);
xor U18141 (N_18141,N_17362,N_17514);
nand U18142 (N_18142,N_17098,N_17490);
and U18143 (N_18143,N_17168,N_17960);
nand U18144 (N_18144,N_17470,N_17861);
nand U18145 (N_18145,N_17911,N_17927);
nor U18146 (N_18146,N_17705,N_17359);
or U18147 (N_18147,N_17333,N_17923);
or U18148 (N_18148,N_17748,N_17184);
and U18149 (N_18149,N_17752,N_17310);
nand U18150 (N_18150,N_17453,N_17220);
nand U18151 (N_18151,N_17869,N_17775);
nor U18152 (N_18152,N_17907,N_17449);
and U18153 (N_18153,N_17765,N_17942);
nor U18154 (N_18154,N_17715,N_17218);
nand U18155 (N_18155,N_17365,N_17254);
nand U18156 (N_18156,N_17145,N_17132);
nand U18157 (N_18157,N_17219,N_17349);
or U18158 (N_18158,N_17855,N_17163);
and U18159 (N_18159,N_17507,N_17109);
xor U18160 (N_18160,N_17250,N_17917);
or U18161 (N_18161,N_17777,N_17647);
and U18162 (N_18162,N_17944,N_17661);
xnor U18163 (N_18163,N_17516,N_17720);
and U18164 (N_18164,N_17390,N_17353);
nand U18165 (N_18165,N_17458,N_17671);
or U18166 (N_18166,N_17201,N_17935);
nand U18167 (N_18167,N_17238,N_17212);
nor U18168 (N_18168,N_17194,N_17203);
nand U18169 (N_18169,N_17293,N_17786);
nand U18170 (N_18170,N_17070,N_17990);
xnor U18171 (N_18171,N_17397,N_17853);
xor U18172 (N_18172,N_17065,N_17549);
xor U18173 (N_18173,N_17572,N_17770);
nand U18174 (N_18174,N_17539,N_17248);
nand U18175 (N_18175,N_17679,N_17931);
xnor U18176 (N_18176,N_17005,N_17579);
or U18177 (N_18177,N_17432,N_17738);
nor U18178 (N_18178,N_17974,N_17693);
nor U18179 (N_18179,N_17965,N_17493);
or U18180 (N_18180,N_17860,N_17536);
or U18181 (N_18181,N_17110,N_17186);
or U18182 (N_18182,N_17239,N_17595);
or U18183 (N_18183,N_17057,N_17259);
nor U18184 (N_18184,N_17424,N_17688);
and U18185 (N_18185,N_17850,N_17379);
xnor U18186 (N_18186,N_17906,N_17084);
or U18187 (N_18187,N_17320,N_17605);
or U18188 (N_18188,N_17272,N_17834);
nand U18189 (N_18189,N_17208,N_17791);
xor U18190 (N_18190,N_17522,N_17382);
and U18191 (N_18191,N_17845,N_17213);
nor U18192 (N_18192,N_17402,N_17728);
nor U18193 (N_18193,N_17616,N_17485);
nand U18194 (N_18194,N_17494,N_17195);
xnor U18195 (N_18195,N_17023,N_17997);
and U18196 (N_18196,N_17075,N_17486);
xor U18197 (N_18197,N_17727,N_17501);
xor U18198 (N_18198,N_17643,N_17018);
or U18199 (N_18199,N_17142,N_17645);
xor U18200 (N_18200,N_17657,N_17723);
nand U18201 (N_18201,N_17112,N_17909);
nor U18202 (N_18202,N_17530,N_17531);
nor U18203 (N_18203,N_17941,N_17404);
and U18204 (N_18204,N_17975,N_17231);
or U18205 (N_18205,N_17551,N_17258);
nor U18206 (N_18206,N_17581,N_17094);
nand U18207 (N_18207,N_17159,N_17701);
and U18208 (N_18208,N_17405,N_17007);
nand U18209 (N_18209,N_17307,N_17079);
and U18210 (N_18210,N_17161,N_17085);
xor U18211 (N_18211,N_17972,N_17235);
nand U18212 (N_18212,N_17155,N_17104);
or U18213 (N_18213,N_17918,N_17338);
nand U18214 (N_18214,N_17285,N_17361);
xnor U18215 (N_18215,N_17515,N_17381);
or U18216 (N_18216,N_17846,N_17826);
and U18217 (N_18217,N_17189,N_17244);
and U18218 (N_18218,N_17533,N_17794);
xnor U18219 (N_18219,N_17905,N_17891);
nor U18220 (N_18220,N_17976,N_17696);
and U18221 (N_18221,N_17257,N_17116);
nand U18222 (N_18222,N_17528,N_17234);
xor U18223 (N_18223,N_17063,N_17062);
nor U18224 (N_18224,N_17477,N_17785);
or U18225 (N_18225,N_17363,N_17989);
xnor U18226 (N_18226,N_17465,N_17781);
nand U18227 (N_18227,N_17847,N_17332);
nand U18228 (N_18228,N_17016,N_17707);
nand U18229 (N_18229,N_17395,N_17008);
and U18230 (N_18230,N_17474,N_17597);
nand U18231 (N_18231,N_17580,N_17151);
nor U18232 (N_18232,N_17527,N_17755);
or U18233 (N_18233,N_17431,N_17245);
or U18234 (N_18234,N_17469,N_17862);
or U18235 (N_18235,N_17560,N_17012);
nand U18236 (N_18236,N_17716,N_17662);
nor U18237 (N_18237,N_17236,N_17224);
nor U18238 (N_18238,N_17865,N_17277);
and U18239 (N_18239,N_17854,N_17427);
xor U18240 (N_18240,N_17173,N_17798);
nor U18241 (N_18241,N_17302,N_17417);
and U18242 (N_18242,N_17077,N_17805);
nor U18243 (N_18243,N_17614,N_17312);
nor U18244 (N_18244,N_17122,N_17052);
and U18245 (N_18245,N_17573,N_17675);
nand U18246 (N_18246,N_17175,N_17588);
and U18247 (N_18247,N_17541,N_17460);
xor U18248 (N_18248,N_17963,N_17454);
and U18249 (N_18249,N_17875,N_17870);
nor U18250 (N_18250,N_17995,N_17964);
xnor U18251 (N_18251,N_17620,N_17388);
xor U18252 (N_18252,N_17502,N_17209);
nand U18253 (N_18253,N_17810,N_17799);
nand U18254 (N_18254,N_17603,N_17730);
nand U18255 (N_18255,N_17746,N_17521);
nor U18256 (N_18256,N_17889,N_17694);
nor U18257 (N_18257,N_17726,N_17264);
nor U18258 (N_18258,N_17613,N_17967);
nor U18259 (N_18259,N_17508,N_17269);
xnor U18260 (N_18260,N_17073,N_17067);
and U18261 (N_18261,N_17833,N_17165);
xor U18262 (N_18262,N_17920,N_17102);
or U18263 (N_18263,N_17952,N_17817);
nand U18264 (N_18264,N_17899,N_17268);
or U18265 (N_18265,N_17761,N_17656);
or U18266 (N_18266,N_17124,N_17796);
and U18267 (N_18267,N_17255,N_17178);
xor U18268 (N_18268,N_17107,N_17028);
or U18269 (N_18269,N_17130,N_17199);
or U18270 (N_18270,N_17304,N_17003);
nor U18271 (N_18271,N_17223,N_17901);
and U18272 (N_18272,N_17108,N_17495);
nor U18273 (N_18273,N_17837,N_17628);
or U18274 (N_18274,N_17410,N_17733);
or U18275 (N_18275,N_17624,N_17461);
or U18276 (N_18276,N_17741,N_17924);
nor U18277 (N_18277,N_17136,N_17782);
nand U18278 (N_18278,N_17642,N_17394);
nor U18279 (N_18279,N_17103,N_17922);
nor U18280 (N_18280,N_17436,N_17006);
xor U18281 (N_18281,N_17526,N_17387);
or U18282 (N_18282,N_17351,N_17939);
and U18283 (N_18283,N_17867,N_17275);
or U18284 (N_18284,N_17347,N_17059);
xnor U18285 (N_18285,N_17753,N_17593);
nor U18286 (N_18286,N_17152,N_17135);
or U18287 (N_18287,N_17169,N_17690);
or U18288 (N_18288,N_17649,N_17709);
nand U18289 (N_18289,N_17599,N_17425);
nor U18290 (N_18290,N_17086,N_17364);
nor U18291 (N_18291,N_17352,N_17369);
or U18292 (N_18292,N_17660,N_17825);
or U18293 (N_18293,N_17247,N_17637);
xor U18294 (N_18294,N_17841,N_17319);
or U18295 (N_18295,N_17594,N_17732);
nand U18296 (N_18296,N_17215,N_17119);
and U18297 (N_18297,N_17139,N_17955);
nand U18298 (N_18298,N_17366,N_17316);
nand U18299 (N_18299,N_17207,N_17937);
nor U18300 (N_18300,N_17676,N_17480);
nand U18301 (N_18301,N_17525,N_17790);
or U18302 (N_18302,N_17324,N_17653);
xor U18303 (N_18303,N_17047,N_17128);
and U18304 (N_18304,N_17314,N_17226);
xor U18305 (N_18305,N_17097,N_17483);
xor U18306 (N_18306,N_17036,N_17699);
nor U18307 (N_18307,N_17802,N_17078);
and U18308 (N_18308,N_17692,N_17806);
nand U18309 (N_18309,N_17877,N_17773);
or U18310 (N_18310,N_17883,N_17538);
nor U18311 (N_18311,N_17544,N_17511);
xor U18312 (N_18312,N_17772,N_17471);
or U18313 (N_18313,N_17433,N_17545);
xnor U18314 (N_18314,N_17874,N_17058);
nand U18315 (N_18315,N_17704,N_17286);
or U18316 (N_18316,N_17951,N_17961);
and U18317 (N_18317,N_17187,N_17042);
and U18318 (N_18318,N_17233,N_17926);
xnor U18319 (N_18319,N_17191,N_17711);
and U18320 (N_18320,N_17334,N_17503);
nor U18321 (N_18321,N_17933,N_17237);
and U18322 (N_18322,N_17921,N_17444);
xor U18323 (N_18323,N_17712,N_17991);
nor U18324 (N_18324,N_17547,N_17736);
or U18325 (N_18325,N_17032,N_17512);
xnor U18326 (N_18326,N_17749,N_17852);
nand U18327 (N_18327,N_17105,N_17342);
nor U18328 (N_18328,N_17225,N_17900);
and U18329 (N_18329,N_17355,N_17380);
nand U18330 (N_18330,N_17621,N_17998);
nor U18331 (N_18331,N_17610,N_17498);
or U18332 (N_18332,N_17176,N_17703);
nor U18333 (N_18333,N_17804,N_17100);
xor U18334 (N_18334,N_17520,N_17166);
xor U18335 (N_18335,N_17323,N_17851);
nor U18336 (N_18336,N_17510,N_17106);
or U18337 (N_18337,N_17529,N_17763);
xor U18338 (N_18338,N_17489,N_17466);
nor U18339 (N_18339,N_17497,N_17035);
or U18340 (N_18340,N_17641,N_17150);
xor U18341 (N_18341,N_17814,N_17326);
or U18342 (N_18342,N_17087,N_17574);
nor U18343 (N_18343,N_17448,N_17204);
and U18344 (N_18344,N_17681,N_17563);
xnor U18345 (N_18345,N_17740,N_17700);
xor U18346 (N_18346,N_17587,N_17101);
nor U18347 (N_18347,N_17813,N_17138);
nor U18348 (N_18348,N_17608,N_17090);
and U18349 (N_18349,N_17393,N_17783);
nor U18350 (N_18350,N_17318,N_17341);
xor U18351 (N_18351,N_17271,N_17290);
nand U18352 (N_18352,N_17838,N_17419);
and U18353 (N_18353,N_17809,N_17818);
nor U18354 (N_18354,N_17373,N_17229);
or U18355 (N_18355,N_17137,N_17409);
nand U18356 (N_18356,N_17172,N_17171);
xor U18357 (N_18357,N_17568,N_17691);
or U18358 (N_18358,N_17821,N_17026);
xnor U18359 (N_18359,N_17153,N_17013);
xor U18360 (N_18360,N_17115,N_17346);
or U18361 (N_18361,N_17121,N_17015);
and U18362 (N_18362,N_17517,N_17908);
nor U18363 (N_18363,N_17648,N_17134);
or U18364 (N_18364,N_17056,N_17930);
or U18365 (N_18365,N_17451,N_17336);
nor U18366 (N_18366,N_17339,N_17482);
and U18367 (N_18367,N_17185,N_17076);
xor U18368 (N_18368,N_17986,N_17519);
or U18369 (N_18369,N_17567,N_17010);
xnor U18370 (N_18370,N_17913,N_17148);
nor U18371 (N_18371,N_17864,N_17956);
and U18372 (N_18372,N_17893,N_17880);
xor U18373 (N_18373,N_17602,N_17849);
nand U18374 (N_18374,N_17680,N_17249);
and U18375 (N_18375,N_17306,N_17504);
xor U18376 (N_18376,N_17820,N_17674);
and U18377 (N_18377,N_17797,N_17561);
nor U18378 (N_18378,N_17462,N_17413);
and U18379 (N_18379,N_17569,N_17627);
and U18380 (N_18380,N_17164,N_17050);
nor U18381 (N_18381,N_17962,N_17606);
nand U18382 (N_18382,N_17578,N_17071);
nand U18383 (N_18383,N_17714,N_17780);
or U18384 (N_18384,N_17457,N_17832);
and U18385 (N_18385,N_17582,N_17360);
xor U18386 (N_18386,N_17828,N_17308);
or U18387 (N_18387,N_17174,N_17916);
nor U18388 (N_18388,N_17027,N_17374);
nand U18389 (N_18389,N_17140,N_17127);
nand U18390 (N_18390,N_17020,N_17196);
or U18391 (N_18391,N_17708,N_17548);
nand U18392 (N_18392,N_17789,N_17827);
or U18393 (N_18393,N_17317,N_17143);
nand U18394 (N_18394,N_17617,N_17982);
or U18395 (N_18395,N_17625,N_17080);
and U18396 (N_18396,N_17710,N_17442);
and U18397 (N_18397,N_17066,N_17546);
nand U18398 (N_18398,N_17992,N_17499);
or U18399 (N_18399,N_17987,N_17146);
nand U18400 (N_18400,N_17758,N_17445);
nor U18401 (N_18401,N_17123,N_17295);
nor U18402 (N_18402,N_17943,N_17767);
nand U18403 (N_18403,N_17559,N_17282);
nor U18404 (N_18404,N_17718,N_17724);
nand U18405 (N_18405,N_17403,N_17261);
or U18406 (N_18406,N_17876,N_17322);
nand U18407 (N_18407,N_17488,N_17687);
nor U18408 (N_18408,N_17274,N_17328);
nor U18409 (N_18409,N_17631,N_17915);
or U18410 (N_18410,N_17557,N_17082);
xnor U18411 (N_18411,N_17273,N_17697);
and U18412 (N_18412,N_17518,N_17386);
nor U18413 (N_18413,N_17542,N_17914);
nand U18414 (N_18414,N_17265,N_17046);
and U18415 (N_18415,N_17464,N_17590);
and U18416 (N_18416,N_17160,N_17435);
nand U18417 (N_18417,N_17808,N_17321);
and U18418 (N_18418,N_17897,N_17803);
nand U18419 (N_18419,N_17296,N_17890);
xnor U18420 (N_18420,N_17636,N_17241);
xor U18421 (N_18421,N_17337,N_17978);
xor U18422 (N_18422,N_17856,N_17949);
and U18423 (N_18423,N_17158,N_17607);
and U18424 (N_18424,N_17385,N_17331);
nand U18425 (N_18425,N_17039,N_17896);
and U18426 (N_18426,N_17284,N_17129);
xnor U18427 (N_18427,N_17664,N_17591);
or U18428 (N_18428,N_17479,N_17948);
or U18429 (N_18429,N_17055,N_17792);
xnor U18430 (N_18430,N_17934,N_17441);
nor U18431 (N_18431,N_17565,N_17554);
nand U18432 (N_18432,N_17778,N_17378);
xor U18433 (N_18433,N_17759,N_17230);
nor U18434 (N_18434,N_17014,N_17354);
nor U18435 (N_18435,N_17157,N_17092);
or U18436 (N_18436,N_17682,N_17340);
or U18437 (N_18437,N_17971,N_17848);
nand U18438 (N_18438,N_17437,N_17376);
nand U18439 (N_18439,N_17686,N_17635);
nand U18440 (N_18440,N_17576,N_17210);
xor U18441 (N_18441,N_17885,N_17988);
nor U18442 (N_18442,N_17945,N_17904);
nor U18443 (N_18443,N_17667,N_17252);
nand U18444 (N_18444,N_17240,N_17872);
nor U18445 (N_18445,N_17214,N_17652);
or U18446 (N_18446,N_17878,N_17260);
and U18447 (N_18447,N_17555,N_17487);
and U18448 (N_18448,N_17500,N_17392);
nand U18449 (N_18449,N_17868,N_17450);
nor U18450 (N_18450,N_17702,N_17281);
nor U18451 (N_18451,N_17043,N_17689);
or U18452 (N_18452,N_17663,N_17162);
nor U18453 (N_18453,N_17940,N_17762);
xor U18454 (N_18454,N_17329,N_17415);
nor U18455 (N_18455,N_17706,N_17757);
or U18456 (N_18456,N_17537,N_17750);
nand U18457 (N_18457,N_17552,N_17879);
xor U18458 (N_18458,N_17147,N_17011);
or U18459 (N_18459,N_17370,N_17966);
xor U18460 (N_18460,N_17391,N_17787);
nor U18461 (N_18461,N_17586,N_17051);
nor U18462 (N_18462,N_17769,N_17734);
nor U18463 (N_18463,N_17455,N_17993);
and U18464 (N_18464,N_17646,N_17377);
or U18465 (N_18465,N_17311,N_17000);
nand U18466 (N_18466,N_17289,N_17266);
nand U18467 (N_18467,N_17325,N_17523);
or U18468 (N_18468,N_17120,N_17438);
xnor U18469 (N_18469,N_17344,N_17283);
xor U18470 (N_18470,N_17739,N_17979);
or U18471 (N_18471,N_17677,N_17021);
xor U18472 (N_18472,N_17072,N_17044);
nor U18473 (N_18473,N_17630,N_17263);
and U18474 (N_18474,N_17061,N_17910);
xnor U18475 (N_18475,N_17959,N_17650);
and U18476 (N_18476,N_17037,N_17721);
and U18477 (N_18477,N_17695,N_17126);
nor U18478 (N_18478,N_17800,N_17881);
or U18479 (N_18479,N_17629,N_17936);
xor U18480 (N_18480,N_17053,N_17884);
nand U18481 (N_18481,N_17513,N_17632);
nor U18482 (N_18482,N_17742,N_17114);
or U18483 (N_18483,N_17776,N_17034);
nor U18484 (N_18484,N_17375,N_17947);
nor U18485 (N_18485,N_17666,N_17744);
or U18486 (N_18486,N_17423,N_17009);
xnor U18487 (N_18487,N_17611,N_17669);
xor U18488 (N_18488,N_17270,N_17980);
xnor U18489 (N_18489,N_17644,N_17428);
and U18490 (N_18490,N_17330,N_17406);
nor U18491 (N_18491,N_17002,N_17859);
or U18492 (N_18492,N_17033,N_17932);
and U18493 (N_18493,N_17760,N_17556);
or U18494 (N_18494,N_17729,N_17422);
and U18495 (N_18495,N_17276,N_17928);
nor U18496 (N_18496,N_17262,N_17125);
nand U18497 (N_18497,N_17278,N_17253);
and U18498 (N_18498,N_17357,N_17343);
nor U18499 (N_18499,N_17177,N_17200);
nand U18500 (N_18500,N_17197,N_17240);
xor U18501 (N_18501,N_17854,N_17391);
or U18502 (N_18502,N_17026,N_17035);
xnor U18503 (N_18503,N_17617,N_17173);
nor U18504 (N_18504,N_17037,N_17931);
xor U18505 (N_18505,N_17596,N_17138);
nor U18506 (N_18506,N_17805,N_17260);
or U18507 (N_18507,N_17885,N_17693);
nor U18508 (N_18508,N_17576,N_17293);
nor U18509 (N_18509,N_17512,N_17710);
xor U18510 (N_18510,N_17284,N_17121);
or U18511 (N_18511,N_17591,N_17244);
nand U18512 (N_18512,N_17992,N_17249);
nor U18513 (N_18513,N_17651,N_17353);
xor U18514 (N_18514,N_17241,N_17522);
xor U18515 (N_18515,N_17396,N_17758);
or U18516 (N_18516,N_17371,N_17968);
xor U18517 (N_18517,N_17384,N_17198);
nor U18518 (N_18518,N_17317,N_17335);
xor U18519 (N_18519,N_17844,N_17581);
and U18520 (N_18520,N_17792,N_17900);
nand U18521 (N_18521,N_17575,N_17112);
nand U18522 (N_18522,N_17513,N_17405);
or U18523 (N_18523,N_17536,N_17828);
xnor U18524 (N_18524,N_17605,N_17985);
nor U18525 (N_18525,N_17599,N_17373);
xnor U18526 (N_18526,N_17819,N_17230);
or U18527 (N_18527,N_17941,N_17991);
and U18528 (N_18528,N_17002,N_17584);
nor U18529 (N_18529,N_17833,N_17003);
or U18530 (N_18530,N_17684,N_17972);
or U18531 (N_18531,N_17734,N_17355);
xnor U18532 (N_18532,N_17674,N_17348);
and U18533 (N_18533,N_17378,N_17652);
or U18534 (N_18534,N_17980,N_17549);
nor U18535 (N_18535,N_17475,N_17894);
and U18536 (N_18536,N_17658,N_17016);
or U18537 (N_18537,N_17359,N_17639);
and U18538 (N_18538,N_17097,N_17326);
and U18539 (N_18539,N_17200,N_17401);
nor U18540 (N_18540,N_17409,N_17302);
xnor U18541 (N_18541,N_17682,N_17229);
nand U18542 (N_18542,N_17671,N_17607);
and U18543 (N_18543,N_17884,N_17844);
xor U18544 (N_18544,N_17470,N_17111);
nor U18545 (N_18545,N_17045,N_17966);
and U18546 (N_18546,N_17735,N_17736);
nor U18547 (N_18547,N_17241,N_17484);
xnor U18548 (N_18548,N_17594,N_17603);
or U18549 (N_18549,N_17557,N_17644);
and U18550 (N_18550,N_17399,N_17701);
or U18551 (N_18551,N_17036,N_17983);
nand U18552 (N_18552,N_17457,N_17155);
and U18553 (N_18553,N_17333,N_17405);
and U18554 (N_18554,N_17050,N_17383);
nand U18555 (N_18555,N_17297,N_17045);
nand U18556 (N_18556,N_17423,N_17395);
nand U18557 (N_18557,N_17177,N_17488);
xor U18558 (N_18558,N_17967,N_17855);
nand U18559 (N_18559,N_17064,N_17649);
nor U18560 (N_18560,N_17174,N_17869);
nand U18561 (N_18561,N_17688,N_17564);
nor U18562 (N_18562,N_17235,N_17444);
and U18563 (N_18563,N_17299,N_17030);
or U18564 (N_18564,N_17952,N_17694);
xnor U18565 (N_18565,N_17608,N_17453);
nand U18566 (N_18566,N_17490,N_17132);
or U18567 (N_18567,N_17379,N_17853);
xnor U18568 (N_18568,N_17170,N_17659);
xor U18569 (N_18569,N_17108,N_17545);
xnor U18570 (N_18570,N_17622,N_17528);
or U18571 (N_18571,N_17671,N_17691);
nor U18572 (N_18572,N_17401,N_17425);
nand U18573 (N_18573,N_17039,N_17396);
or U18574 (N_18574,N_17309,N_17730);
nor U18575 (N_18575,N_17058,N_17353);
and U18576 (N_18576,N_17242,N_17896);
xnor U18577 (N_18577,N_17765,N_17093);
or U18578 (N_18578,N_17469,N_17971);
xor U18579 (N_18579,N_17550,N_17608);
or U18580 (N_18580,N_17795,N_17027);
and U18581 (N_18581,N_17034,N_17313);
nand U18582 (N_18582,N_17216,N_17884);
and U18583 (N_18583,N_17330,N_17942);
nor U18584 (N_18584,N_17470,N_17526);
xor U18585 (N_18585,N_17349,N_17215);
nor U18586 (N_18586,N_17180,N_17333);
nand U18587 (N_18587,N_17408,N_17052);
nor U18588 (N_18588,N_17753,N_17016);
nor U18589 (N_18589,N_17626,N_17380);
nand U18590 (N_18590,N_17624,N_17127);
nor U18591 (N_18591,N_17866,N_17533);
xor U18592 (N_18592,N_17525,N_17712);
xnor U18593 (N_18593,N_17477,N_17936);
and U18594 (N_18594,N_17474,N_17210);
nor U18595 (N_18595,N_17685,N_17919);
nand U18596 (N_18596,N_17010,N_17033);
nor U18597 (N_18597,N_17364,N_17624);
xnor U18598 (N_18598,N_17977,N_17565);
nand U18599 (N_18599,N_17381,N_17010);
or U18600 (N_18600,N_17300,N_17816);
nand U18601 (N_18601,N_17596,N_17617);
nand U18602 (N_18602,N_17436,N_17979);
xnor U18603 (N_18603,N_17463,N_17224);
and U18604 (N_18604,N_17515,N_17231);
or U18605 (N_18605,N_17281,N_17393);
nand U18606 (N_18606,N_17299,N_17788);
nand U18607 (N_18607,N_17439,N_17510);
or U18608 (N_18608,N_17511,N_17576);
xor U18609 (N_18609,N_17641,N_17038);
and U18610 (N_18610,N_17215,N_17776);
nand U18611 (N_18611,N_17028,N_17689);
nand U18612 (N_18612,N_17860,N_17861);
nand U18613 (N_18613,N_17252,N_17764);
or U18614 (N_18614,N_17052,N_17048);
and U18615 (N_18615,N_17002,N_17057);
nor U18616 (N_18616,N_17413,N_17809);
and U18617 (N_18617,N_17593,N_17838);
nor U18618 (N_18618,N_17381,N_17967);
and U18619 (N_18619,N_17308,N_17435);
nor U18620 (N_18620,N_17902,N_17018);
and U18621 (N_18621,N_17506,N_17613);
and U18622 (N_18622,N_17766,N_17985);
nand U18623 (N_18623,N_17100,N_17255);
nor U18624 (N_18624,N_17688,N_17149);
nand U18625 (N_18625,N_17436,N_17628);
or U18626 (N_18626,N_17689,N_17681);
nand U18627 (N_18627,N_17742,N_17582);
nand U18628 (N_18628,N_17759,N_17582);
and U18629 (N_18629,N_17300,N_17607);
nor U18630 (N_18630,N_17805,N_17208);
and U18631 (N_18631,N_17488,N_17137);
nor U18632 (N_18632,N_17804,N_17082);
and U18633 (N_18633,N_17651,N_17772);
and U18634 (N_18634,N_17011,N_17593);
or U18635 (N_18635,N_17216,N_17942);
nand U18636 (N_18636,N_17540,N_17478);
nor U18637 (N_18637,N_17263,N_17256);
nand U18638 (N_18638,N_17917,N_17200);
or U18639 (N_18639,N_17917,N_17759);
nor U18640 (N_18640,N_17241,N_17756);
and U18641 (N_18641,N_17225,N_17006);
or U18642 (N_18642,N_17783,N_17349);
nor U18643 (N_18643,N_17447,N_17163);
and U18644 (N_18644,N_17121,N_17600);
or U18645 (N_18645,N_17068,N_17768);
nand U18646 (N_18646,N_17465,N_17744);
nand U18647 (N_18647,N_17600,N_17235);
nor U18648 (N_18648,N_17208,N_17241);
and U18649 (N_18649,N_17294,N_17585);
and U18650 (N_18650,N_17925,N_17449);
or U18651 (N_18651,N_17256,N_17265);
nand U18652 (N_18652,N_17111,N_17285);
nor U18653 (N_18653,N_17993,N_17429);
and U18654 (N_18654,N_17657,N_17352);
or U18655 (N_18655,N_17962,N_17727);
and U18656 (N_18656,N_17266,N_17325);
or U18657 (N_18657,N_17353,N_17129);
and U18658 (N_18658,N_17154,N_17436);
nor U18659 (N_18659,N_17223,N_17899);
or U18660 (N_18660,N_17909,N_17711);
xor U18661 (N_18661,N_17892,N_17895);
and U18662 (N_18662,N_17293,N_17416);
xor U18663 (N_18663,N_17154,N_17008);
xor U18664 (N_18664,N_17332,N_17571);
or U18665 (N_18665,N_17832,N_17078);
xnor U18666 (N_18666,N_17776,N_17962);
nand U18667 (N_18667,N_17370,N_17267);
and U18668 (N_18668,N_17800,N_17426);
xor U18669 (N_18669,N_17661,N_17438);
nand U18670 (N_18670,N_17637,N_17562);
xnor U18671 (N_18671,N_17624,N_17285);
or U18672 (N_18672,N_17765,N_17569);
nor U18673 (N_18673,N_17114,N_17518);
and U18674 (N_18674,N_17583,N_17046);
nor U18675 (N_18675,N_17913,N_17002);
nand U18676 (N_18676,N_17037,N_17059);
nand U18677 (N_18677,N_17036,N_17547);
xor U18678 (N_18678,N_17963,N_17588);
xnor U18679 (N_18679,N_17955,N_17894);
xnor U18680 (N_18680,N_17390,N_17940);
and U18681 (N_18681,N_17139,N_17168);
xor U18682 (N_18682,N_17152,N_17839);
xor U18683 (N_18683,N_17371,N_17304);
nor U18684 (N_18684,N_17121,N_17384);
or U18685 (N_18685,N_17555,N_17816);
xnor U18686 (N_18686,N_17674,N_17554);
and U18687 (N_18687,N_17429,N_17021);
and U18688 (N_18688,N_17997,N_17952);
nor U18689 (N_18689,N_17219,N_17687);
nand U18690 (N_18690,N_17189,N_17832);
or U18691 (N_18691,N_17097,N_17488);
nor U18692 (N_18692,N_17805,N_17168);
nor U18693 (N_18693,N_17302,N_17163);
nand U18694 (N_18694,N_17448,N_17253);
or U18695 (N_18695,N_17897,N_17725);
or U18696 (N_18696,N_17196,N_17673);
xor U18697 (N_18697,N_17688,N_17023);
xnor U18698 (N_18698,N_17376,N_17836);
nor U18699 (N_18699,N_17901,N_17519);
and U18700 (N_18700,N_17093,N_17457);
xnor U18701 (N_18701,N_17794,N_17025);
or U18702 (N_18702,N_17302,N_17732);
xnor U18703 (N_18703,N_17913,N_17876);
nand U18704 (N_18704,N_17511,N_17677);
or U18705 (N_18705,N_17747,N_17418);
nor U18706 (N_18706,N_17713,N_17584);
nand U18707 (N_18707,N_17807,N_17142);
nand U18708 (N_18708,N_17708,N_17560);
or U18709 (N_18709,N_17753,N_17976);
and U18710 (N_18710,N_17215,N_17682);
and U18711 (N_18711,N_17169,N_17592);
nand U18712 (N_18712,N_17317,N_17084);
nor U18713 (N_18713,N_17680,N_17783);
and U18714 (N_18714,N_17785,N_17126);
or U18715 (N_18715,N_17997,N_17280);
and U18716 (N_18716,N_17205,N_17536);
and U18717 (N_18717,N_17593,N_17572);
nor U18718 (N_18718,N_17352,N_17322);
nand U18719 (N_18719,N_17031,N_17541);
and U18720 (N_18720,N_17860,N_17218);
nand U18721 (N_18721,N_17517,N_17968);
nand U18722 (N_18722,N_17016,N_17407);
and U18723 (N_18723,N_17223,N_17039);
and U18724 (N_18724,N_17462,N_17689);
xor U18725 (N_18725,N_17852,N_17279);
nor U18726 (N_18726,N_17291,N_17527);
nand U18727 (N_18727,N_17820,N_17325);
or U18728 (N_18728,N_17254,N_17837);
and U18729 (N_18729,N_17013,N_17928);
and U18730 (N_18730,N_17672,N_17847);
nand U18731 (N_18731,N_17281,N_17758);
and U18732 (N_18732,N_17548,N_17044);
nand U18733 (N_18733,N_17787,N_17952);
or U18734 (N_18734,N_17742,N_17210);
or U18735 (N_18735,N_17629,N_17565);
or U18736 (N_18736,N_17699,N_17874);
nor U18737 (N_18737,N_17348,N_17751);
nand U18738 (N_18738,N_17861,N_17683);
xor U18739 (N_18739,N_17091,N_17002);
and U18740 (N_18740,N_17295,N_17109);
nor U18741 (N_18741,N_17027,N_17691);
xnor U18742 (N_18742,N_17056,N_17268);
nor U18743 (N_18743,N_17524,N_17988);
and U18744 (N_18744,N_17639,N_17509);
nand U18745 (N_18745,N_17482,N_17271);
xnor U18746 (N_18746,N_17701,N_17940);
or U18747 (N_18747,N_17473,N_17010);
nand U18748 (N_18748,N_17989,N_17652);
and U18749 (N_18749,N_17081,N_17457);
nand U18750 (N_18750,N_17621,N_17794);
nor U18751 (N_18751,N_17872,N_17023);
and U18752 (N_18752,N_17357,N_17344);
or U18753 (N_18753,N_17269,N_17660);
nand U18754 (N_18754,N_17176,N_17353);
nor U18755 (N_18755,N_17220,N_17240);
or U18756 (N_18756,N_17895,N_17801);
or U18757 (N_18757,N_17496,N_17949);
and U18758 (N_18758,N_17865,N_17380);
nand U18759 (N_18759,N_17976,N_17752);
nor U18760 (N_18760,N_17307,N_17254);
and U18761 (N_18761,N_17396,N_17209);
nor U18762 (N_18762,N_17281,N_17089);
and U18763 (N_18763,N_17930,N_17298);
or U18764 (N_18764,N_17815,N_17259);
xor U18765 (N_18765,N_17872,N_17149);
or U18766 (N_18766,N_17982,N_17701);
nor U18767 (N_18767,N_17668,N_17381);
and U18768 (N_18768,N_17610,N_17044);
nor U18769 (N_18769,N_17929,N_17477);
nand U18770 (N_18770,N_17299,N_17944);
nor U18771 (N_18771,N_17700,N_17251);
nand U18772 (N_18772,N_17863,N_17242);
nand U18773 (N_18773,N_17499,N_17554);
and U18774 (N_18774,N_17723,N_17492);
and U18775 (N_18775,N_17779,N_17896);
nor U18776 (N_18776,N_17259,N_17127);
nor U18777 (N_18777,N_17035,N_17168);
and U18778 (N_18778,N_17520,N_17655);
xor U18779 (N_18779,N_17487,N_17394);
nand U18780 (N_18780,N_17805,N_17553);
nand U18781 (N_18781,N_17816,N_17625);
nand U18782 (N_18782,N_17152,N_17583);
or U18783 (N_18783,N_17154,N_17682);
and U18784 (N_18784,N_17274,N_17023);
xnor U18785 (N_18785,N_17497,N_17092);
nand U18786 (N_18786,N_17061,N_17367);
nor U18787 (N_18787,N_17322,N_17533);
and U18788 (N_18788,N_17148,N_17184);
xnor U18789 (N_18789,N_17723,N_17072);
and U18790 (N_18790,N_17790,N_17310);
xor U18791 (N_18791,N_17056,N_17572);
nand U18792 (N_18792,N_17421,N_17487);
xor U18793 (N_18793,N_17566,N_17469);
nand U18794 (N_18794,N_17896,N_17069);
nand U18795 (N_18795,N_17370,N_17226);
nor U18796 (N_18796,N_17213,N_17463);
nor U18797 (N_18797,N_17654,N_17174);
xor U18798 (N_18798,N_17595,N_17317);
xnor U18799 (N_18799,N_17656,N_17902);
xor U18800 (N_18800,N_17094,N_17258);
nor U18801 (N_18801,N_17962,N_17182);
or U18802 (N_18802,N_17123,N_17928);
and U18803 (N_18803,N_17135,N_17247);
nand U18804 (N_18804,N_17416,N_17942);
and U18805 (N_18805,N_17212,N_17201);
xor U18806 (N_18806,N_17122,N_17056);
xor U18807 (N_18807,N_17885,N_17801);
nand U18808 (N_18808,N_17592,N_17792);
xor U18809 (N_18809,N_17192,N_17646);
and U18810 (N_18810,N_17507,N_17096);
or U18811 (N_18811,N_17504,N_17577);
or U18812 (N_18812,N_17398,N_17460);
xor U18813 (N_18813,N_17518,N_17121);
xor U18814 (N_18814,N_17990,N_17806);
xnor U18815 (N_18815,N_17415,N_17241);
nor U18816 (N_18816,N_17592,N_17942);
or U18817 (N_18817,N_17658,N_17140);
xor U18818 (N_18818,N_17707,N_17834);
nand U18819 (N_18819,N_17494,N_17207);
or U18820 (N_18820,N_17803,N_17065);
or U18821 (N_18821,N_17926,N_17487);
nand U18822 (N_18822,N_17760,N_17488);
nand U18823 (N_18823,N_17419,N_17930);
and U18824 (N_18824,N_17684,N_17567);
nor U18825 (N_18825,N_17691,N_17881);
or U18826 (N_18826,N_17562,N_17244);
and U18827 (N_18827,N_17859,N_17029);
nand U18828 (N_18828,N_17822,N_17388);
nor U18829 (N_18829,N_17822,N_17997);
or U18830 (N_18830,N_17566,N_17413);
or U18831 (N_18831,N_17142,N_17383);
nand U18832 (N_18832,N_17794,N_17084);
nor U18833 (N_18833,N_17129,N_17293);
nor U18834 (N_18834,N_17738,N_17161);
or U18835 (N_18835,N_17801,N_17423);
xor U18836 (N_18836,N_17952,N_17626);
nor U18837 (N_18837,N_17740,N_17667);
nand U18838 (N_18838,N_17473,N_17900);
or U18839 (N_18839,N_17053,N_17792);
nor U18840 (N_18840,N_17920,N_17790);
nand U18841 (N_18841,N_17551,N_17159);
or U18842 (N_18842,N_17048,N_17287);
nand U18843 (N_18843,N_17715,N_17761);
nor U18844 (N_18844,N_17853,N_17939);
xor U18845 (N_18845,N_17729,N_17762);
nand U18846 (N_18846,N_17739,N_17675);
and U18847 (N_18847,N_17274,N_17090);
and U18848 (N_18848,N_17793,N_17235);
xnor U18849 (N_18849,N_17070,N_17668);
xnor U18850 (N_18850,N_17685,N_17309);
and U18851 (N_18851,N_17011,N_17251);
nor U18852 (N_18852,N_17074,N_17845);
nor U18853 (N_18853,N_17598,N_17692);
xor U18854 (N_18854,N_17191,N_17993);
nor U18855 (N_18855,N_17031,N_17076);
or U18856 (N_18856,N_17234,N_17345);
nand U18857 (N_18857,N_17536,N_17553);
nand U18858 (N_18858,N_17020,N_17422);
xnor U18859 (N_18859,N_17923,N_17159);
nand U18860 (N_18860,N_17712,N_17138);
nand U18861 (N_18861,N_17777,N_17235);
xor U18862 (N_18862,N_17438,N_17156);
xor U18863 (N_18863,N_17163,N_17487);
or U18864 (N_18864,N_17148,N_17542);
nor U18865 (N_18865,N_17662,N_17003);
and U18866 (N_18866,N_17488,N_17423);
xor U18867 (N_18867,N_17976,N_17211);
or U18868 (N_18868,N_17027,N_17835);
xnor U18869 (N_18869,N_17760,N_17829);
xor U18870 (N_18870,N_17397,N_17348);
nor U18871 (N_18871,N_17640,N_17231);
nand U18872 (N_18872,N_17621,N_17401);
nor U18873 (N_18873,N_17738,N_17158);
xor U18874 (N_18874,N_17927,N_17817);
nor U18875 (N_18875,N_17546,N_17255);
or U18876 (N_18876,N_17082,N_17420);
xor U18877 (N_18877,N_17967,N_17854);
and U18878 (N_18878,N_17329,N_17626);
nand U18879 (N_18879,N_17713,N_17085);
or U18880 (N_18880,N_17423,N_17505);
and U18881 (N_18881,N_17751,N_17704);
xnor U18882 (N_18882,N_17457,N_17792);
and U18883 (N_18883,N_17401,N_17715);
nor U18884 (N_18884,N_17582,N_17397);
xnor U18885 (N_18885,N_17648,N_17659);
or U18886 (N_18886,N_17140,N_17076);
nand U18887 (N_18887,N_17126,N_17170);
and U18888 (N_18888,N_17869,N_17584);
nand U18889 (N_18889,N_17452,N_17332);
nand U18890 (N_18890,N_17757,N_17652);
xor U18891 (N_18891,N_17805,N_17792);
xnor U18892 (N_18892,N_17512,N_17523);
nand U18893 (N_18893,N_17628,N_17168);
nor U18894 (N_18894,N_17394,N_17224);
xnor U18895 (N_18895,N_17002,N_17378);
and U18896 (N_18896,N_17037,N_17936);
nor U18897 (N_18897,N_17796,N_17215);
nor U18898 (N_18898,N_17455,N_17709);
xor U18899 (N_18899,N_17150,N_17286);
xnor U18900 (N_18900,N_17183,N_17381);
or U18901 (N_18901,N_17459,N_17183);
nor U18902 (N_18902,N_17364,N_17208);
nand U18903 (N_18903,N_17630,N_17689);
nand U18904 (N_18904,N_17195,N_17771);
or U18905 (N_18905,N_17736,N_17323);
nand U18906 (N_18906,N_17385,N_17758);
and U18907 (N_18907,N_17435,N_17511);
nand U18908 (N_18908,N_17884,N_17921);
or U18909 (N_18909,N_17488,N_17636);
xnor U18910 (N_18910,N_17077,N_17630);
xor U18911 (N_18911,N_17010,N_17866);
or U18912 (N_18912,N_17319,N_17491);
nand U18913 (N_18913,N_17019,N_17786);
or U18914 (N_18914,N_17915,N_17425);
xnor U18915 (N_18915,N_17093,N_17529);
xor U18916 (N_18916,N_17565,N_17475);
nor U18917 (N_18917,N_17890,N_17321);
xor U18918 (N_18918,N_17239,N_17558);
nor U18919 (N_18919,N_17423,N_17402);
xor U18920 (N_18920,N_17897,N_17628);
and U18921 (N_18921,N_17231,N_17613);
nor U18922 (N_18922,N_17215,N_17848);
nand U18923 (N_18923,N_17289,N_17357);
nor U18924 (N_18924,N_17088,N_17640);
nor U18925 (N_18925,N_17174,N_17148);
xnor U18926 (N_18926,N_17244,N_17681);
or U18927 (N_18927,N_17992,N_17462);
nand U18928 (N_18928,N_17198,N_17972);
nor U18929 (N_18929,N_17193,N_17643);
nand U18930 (N_18930,N_17846,N_17013);
nor U18931 (N_18931,N_17458,N_17115);
or U18932 (N_18932,N_17277,N_17114);
nand U18933 (N_18933,N_17755,N_17640);
nor U18934 (N_18934,N_17572,N_17317);
or U18935 (N_18935,N_17612,N_17654);
xnor U18936 (N_18936,N_17721,N_17966);
nand U18937 (N_18937,N_17913,N_17424);
nand U18938 (N_18938,N_17463,N_17341);
or U18939 (N_18939,N_17119,N_17696);
xnor U18940 (N_18940,N_17709,N_17330);
nand U18941 (N_18941,N_17793,N_17998);
nand U18942 (N_18942,N_17485,N_17942);
nor U18943 (N_18943,N_17068,N_17836);
or U18944 (N_18944,N_17236,N_17726);
and U18945 (N_18945,N_17064,N_17336);
xor U18946 (N_18946,N_17292,N_17630);
and U18947 (N_18947,N_17409,N_17775);
xnor U18948 (N_18948,N_17210,N_17372);
nand U18949 (N_18949,N_17836,N_17958);
xnor U18950 (N_18950,N_17224,N_17885);
nor U18951 (N_18951,N_17479,N_17298);
or U18952 (N_18952,N_17376,N_17960);
or U18953 (N_18953,N_17870,N_17084);
nor U18954 (N_18954,N_17446,N_17980);
xor U18955 (N_18955,N_17687,N_17380);
nand U18956 (N_18956,N_17665,N_17071);
and U18957 (N_18957,N_17796,N_17056);
or U18958 (N_18958,N_17373,N_17401);
nor U18959 (N_18959,N_17695,N_17707);
or U18960 (N_18960,N_17185,N_17510);
or U18961 (N_18961,N_17758,N_17978);
and U18962 (N_18962,N_17172,N_17728);
nand U18963 (N_18963,N_17865,N_17471);
xor U18964 (N_18964,N_17113,N_17855);
or U18965 (N_18965,N_17534,N_17337);
nand U18966 (N_18966,N_17497,N_17110);
xor U18967 (N_18967,N_17203,N_17846);
and U18968 (N_18968,N_17102,N_17644);
nand U18969 (N_18969,N_17666,N_17373);
or U18970 (N_18970,N_17278,N_17551);
and U18971 (N_18971,N_17636,N_17954);
xor U18972 (N_18972,N_17874,N_17486);
xor U18973 (N_18973,N_17489,N_17349);
or U18974 (N_18974,N_17562,N_17682);
or U18975 (N_18975,N_17570,N_17804);
xnor U18976 (N_18976,N_17718,N_17690);
or U18977 (N_18977,N_17914,N_17144);
xor U18978 (N_18978,N_17774,N_17866);
xnor U18979 (N_18979,N_17988,N_17212);
and U18980 (N_18980,N_17898,N_17633);
xor U18981 (N_18981,N_17191,N_17515);
or U18982 (N_18982,N_17819,N_17997);
nor U18983 (N_18983,N_17984,N_17533);
xnor U18984 (N_18984,N_17156,N_17259);
xnor U18985 (N_18985,N_17076,N_17737);
xnor U18986 (N_18986,N_17608,N_17737);
and U18987 (N_18987,N_17094,N_17736);
nand U18988 (N_18988,N_17133,N_17110);
xnor U18989 (N_18989,N_17632,N_17737);
and U18990 (N_18990,N_17510,N_17390);
or U18991 (N_18991,N_17253,N_17045);
or U18992 (N_18992,N_17957,N_17550);
nor U18993 (N_18993,N_17186,N_17568);
and U18994 (N_18994,N_17379,N_17870);
and U18995 (N_18995,N_17487,N_17766);
xnor U18996 (N_18996,N_17528,N_17654);
or U18997 (N_18997,N_17980,N_17258);
nand U18998 (N_18998,N_17892,N_17016);
xnor U18999 (N_18999,N_17128,N_17835);
and U19000 (N_19000,N_18008,N_18874);
and U19001 (N_19001,N_18011,N_18437);
xor U19002 (N_19002,N_18863,N_18359);
nand U19003 (N_19003,N_18763,N_18611);
nand U19004 (N_19004,N_18231,N_18302);
nor U19005 (N_19005,N_18877,N_18978);
nor U19006 (N_19006,N_18868,N_18975);
xnor U19007 (N_19007,N_18639,N_18278);
nand U19008 (N_19008,N_18699,N_18864);
and U19009 (N_19009,N_18123,N_18372);
nor U19010 (N_19010,N_18413,N_18427);
xnor U19011 (N_19011,N_18381,N_18705);
nor U19012 (N_19012,N_18842,N_18766);
or U19013 (N_19013,N_18656,N_18322);
nor U19014 (N_19014,N_18569,N_18325);
xor U19015 (N_19015,N_18233,N_18781);
and U19016 (N_19016,N_18734,N_18308);
nor U19017 (N_19017,N_18519,N_18374);
xor U19018 (N_19018,N_18564,N_18745);
or U19019 (N_19019,N_18720,N_18058);
nand U19020 (N_19020,N_18504,N_18019);
and U19021 (N_19021,N_18502,N_18744);
or U19022 (N_19022,N_18615,N_18009);
nor U19023 (N_19023,N_18222,N_18421);
or U19024 (N_19024,N_18832,N_18886);
or U19025 (N_19025,N_18742,N_18860);
nand U19026 (N_19026,N_18314,N_18809);
and U19027 (N_19027,N_18357,N_18855);
nor U19028 (N_19028,N_18419,N_18884);
xor U19029 (N_19029,N_18342,N_18632);
nand U19030 (N_19030,N_18827,N_18338);
or U19031 (N_19031,N_18549,N_18826);
nand U19032 (N_19032,N_18689,N_18562);
nor U19033 (N_19033,N_18143,N_18708);
and U19034 (N_19034,N_18451,N_18094);
xor U19035 (N_19035,N_18701,N_18186);
xnor U19036 (N_19036,N_18136,N_18944);
or U19037 (N_19037,N_18955,N_18082);
xnor U19038 (N_19038,N_18483,N_18930);
nor U19039 (N_19039,N_18379,N_18003);
and U19040 (N_19040,N_18903,N_18730);
and U19041 (N_19041,N_18212,N_18643);
or U19042 (N_19042,N_18729,N_18459);
or U19043 (N_19043,N_18373,N_18821);
and U19044 (N_19044,N_18259,N_18098);
nand U19045 (N_19045,N_18360,N_18773);
nor U19046 (N_19046,N_18029,N_18382);
nor U19047 (N_19047,N_18588,N_18531);
nand U19048 (N_19048,N_18070,N_18320);
or U19049 (N_19049,N_18608,N_18736);
and U19050 (N_19050,N_18538,N_18468);
nor U19051 (N_19051,N_18568,N_18396);
and U19052 (N_19052,N_18171,N_18797);
nor U19053 (N_19053,N_18445,N_18919);
nor U19054 (N_19054,N_18393,N_18962);
nand U19055 (N_19055,N_18244,N_18316);
or U19056 (N_19056,N_18496,N_18706);
xnor U19057 (N_19057,N_18390,N_18464);
and U19058 (N_19058,N_18587,N_18295);
xor U19059 (N_19059,N_18130,N_18076);
nand U19060 (N_19060,N_18285,N_18274);
and U19061 (N_19061,N_18198,N_18949);
xor U19062 (N_19062,N_18361,N_18916);
and U19063 (N_19063,N_18167,N_18311);
xnor U19064 (N_19064,N_18237,N_18652);
nand U19065 (N_19065,N_18848,N_18328);
and U19066 (N_19066,N_18682,N_18994);
xnor U19067 (N_19067,N_18429,N_18280);
nand U19068 (N_19068,N_18528,N_18087);
and U19069 (N_19069,N_18594,N_18047);
nand U19070 (N_19070,N_18592,N_18432);
xnor U19071 (N_19071,N_18722,N_18931);
xor U19072 (N_19072,N_18966,N_18634);
nand U19073 (N_19073,N_18607,N_18650);
and U19074 (N_19074,N_18854,N_18807);
nand U19075 (N_19075,N_18885,N_18300);
xnor U19076 (N_19076,N_18671,N_18973);
nand U19077 (N_19077,N_18631,N_18152);
nand U19078 (N_19078,N_18619,N_18642);
xnor U19079 (N_19079,N_18754,N_18750);
and U19080 (N_19080,N_18310,N_18490);
nand U19081 (N_19081,N_18190,N_18081);
nand U19082 (N_19082,N_18493,N_18065);
and U19083 (N_19083,N_18574,N_18018);
nand U19084 (N_19084,N_18089,N_18113);
xnor U19085 (N_19085,N_18728,N_18684);
and U19086 (N_19086,N_18911,N_18756);
nor U19087 (N_19087,N_18563,N_18596);
or U19088 (N_19088,N_18108,N_18543);
nand U19089 (N_19089,N_18723,N_18679);
or U19090 (N_19090,N_18238,N_18096);
xor U19091 (N_19091,N_18853,N_18673);
or U19092 (N_19092,N_18120,N_18461);
or U19093 (N_19093,N_18016,N_18272);
xor U19094 (N_19094,N_18192,N_18193);
or U19095 (N_19095,N_18902,N_18028);
nand U19096 (N_19096,N_18250,N_18995);
nor U19097 (N_19097,N_18195,N_18035);
nor U19098 (N_19098,N_18678,N_18450);
nor U19099 (N_19099,N_18454,N_18710);
and U19100 (N_19100,N_18584,N_18824);
nand U19101 (N_19101,N_18103,N_18999);
nor U19102 (N_19102,N_18401,N_18162);
and U19103 (N_19103,N_18297,N_18128);
nand U19104 (N_19104,N_18982,N_18273);
or U19105 (N_19105,N_18808,N_18470);
nor U19106 (N_19106,N_18291,N_18676);
or U19107 (N_19107,N_18001,N_18399);
nand U19108 (N_19108,N_18905,N_18458);
nor U19109 (N_19109,N_18312,N_18606);
or U19110 (N_19110,N_18666,N_18185);
and U19111 (N_19111,N_18668,N_18547);
xor U19112 (N_19112,N_18946,N_18157);
nand U19113 (N_19113,N_18661,N_18332);
or U19114 (N_19114,N_18262,N_18669);
nor U19115 (N_19115,N_18922,N_18918);
nand U19116 (N_19116,N_18474,N_18778);
and U19117 (N_19117,N_18938,N_18201);
or U19118 (N_19118,N_18112,N_18214);
or U19119 (N_19119,N_18500,N_18488);
and U19120 (N_19120,N_18712,N_18789);
nand U19121 (N_19121,N_18782,N_18852);
or U19122 (N_19122,N_18617,N_18337);
and U19123 (N_19123,N_18404,N_18518);
or U19124 (N_19124,N_18200,N_18414);
nor U19125 (N_19125,N_18038,N_18431);
nor U19126 (N_19126,N_18329,N_18635);
nand U19127 (N_19127,N_18106,N_18370);
or U19128 (N_19128,N_18614,N_18585);
xnor U19129 (N_19129,N_18339,N_18024);
nor U19130 (N_19130,N_18784,N_18960);
nand U19131 (N_19131,N_18327,N_18934);
and U19132 (N_19132,N_18392,N_18079);
nor U19133 (N_19133,N_18037,N_18180);
nor U19134 (N_19134,N_18025,N_18846);
nand U19135 (N_19135,N_18915,N_18457);
and U19136 (N_19136,N_18412,N_18448);
or U19137 (N_19137,N_18077,N_18577);
and U19138 (N_19138,N_18558,N_18914);
nor U19139 (N_19139,N_18263,N_18407);
nand U19140 (N_19140,N_18845,N_18276);
or U19141 (N_19141,N_18246,N_18731);
nand U19142 (N_19142,N_18866,N_18565);
and U19143 (N_19143,N_18164,N_18967);
nor U19144 (N_19144,N_18690,N_18172);
nor U19145 (N_19145,N_18403,N_18804);
nor U19146 (N_19146,N_18309,N_18732);
and U19147 (N_19147,N_18232,N_18839);
or U19148 (N_19148,N_18163,N_18674);
xnor U19149 (N_19149,N_18436,N_18012);
nor U19150 (N_19150,N_18304,N_18299);
nor U19151 (N_19151,N_18737,N_18814);
or U19152 (N_19152,N_18741,N_18017);
nor U19153 (N_19153,N_18501,N_18184);
nor U19154 (N_19154,N_18426,N_18770);
xor U19155 (N_19155,N_18665,N_18455);
nor U19156 (N_19156,N_18859,N_18133);
nand U19157 (N_19157,N_18697,N_18121);
nand U19158 (N_19158,N_18397,N_18482);
nor U19159 (N_19159,N_18318,N_18888);
nor U19160 (N_19160,N_18823,N_18229);
nor U19161 (N_19161,N_18509,N_18771);
or U19162 (N_19162,N_18566,N_18385);
and U19163 (N_19163,N_18199,N_18447);
and U19164 (N_19164,N_18050,N_18521);
nand U19165 (N_19165,N_18078,N_18289);
nor U19166 (N_19166,N_18211,N_18939);
and U19167 (N_19167,N_18260,N_18576);
or U19168 (N_19168,N_18896,N_18213);
or U19169 (N_19169,N_18618,N_18168);
nor U19170 (N_19170,N_18027,N_18366);
and U19171 (N_19171,N_18481,N_18176);
nand U19172 (N_19172,N_18672,N_18578);
nor U19173 (N_19173,N_18124,N_18368);
nand U19174 (N_19174,N_18142,N_18159);
nand U19175 (N_19175,N_18970,N_18227);
xnor U19176 (N_19176,N_18725,N_18139);
and U19177 (N_19177,N_18825,N_18872);
nand U19178 (N_19178,N_18529,N_18740);
nor U19179 (N_19179,N_18718,N_18242);
and U19180 (N_19180,N_18252,N_18776);
nand U19181 (N_19181,N_18840,N_18075);
xor U19182 (N_19182,N_18135,N_18284);
or U19183 (N_19183,N_18986,N_18719);
or U19184 (N_19184,N_18616,N_18384);
xnor U19185 (N_19185,N_18867,N_18440);
and U19186 (N_19186,N_18462,N_18803);
and U19187 (N_19187,N_18505,N_18836);
xnor U19188 (N_19188,N_18294,N_18367);
nand U19189 (N_19189,N_18972,N_18216);
nor U19190 (N_19190,N_18834,N_18465);
nor U19191 (N_19191,N_18410,N_18345);
nor U19192 (N_19192,N_18540,N_18453);
and U19193 (N_19193,N_18489,N_18416);
nor U19194 (N_19194,N_18476,N_18156);
or U19195 (N_19195,N_18064,N_18062);
or U19196 (N_19196,N_18129,N_18288);
and U19197 (N_19197,N_18892,N_18704);
or U19198 (N_19198,N_18068,N_18109);
nand U19199 (N_19199,N_18083,N_18411);
or U19200 (N_19200,N_18749,N_18165);
nand U19201 (N_19201,N_18985,N_18015);
nor U19202 (N_19202,N_18871,N_18353);
nand U19203 (N_19203,N_18460,N_18535);
nand U19204 (N_19204,N_18516,N_18929);
nand U19205 (N_19205,N_18685,N_18386);
or U19206 (N_19206,N_18054,N_18467);
and U19207 (N_19207,N_18582,N_18640);
and U19208 (N_19208,N_18444,N_18048);
xnor U19209 (N_19209,N_18768,N_18006);
and U19210 (N_19210,N_18210,N_18542);
or U19211 (N_19211,N_18593,N_18716);
xor U19212 (N_19212,N_18248,N_18556);
xor U19213 (N_19213,N_18228,N_18321);
nor U19214 (N_19214,N_18378,N_18235);
xor U19215 (N_19215,N_18355,N_18182);
nor U19216 (N_19216,N_18988,N_18816);
nand U19217 (N_19217,N_18545,N_18951);
and U19218 (N_19218,N_18950,N_18936);
nor U19219 (N_19219,N_18243,N_18925);
nor U19220 (N_19220,N_18424,N_18567);
and U19221 (N_19221,N_18900,N_18503);
nand U19222 (N_19222,N_18620,N_18645);
or U19223 (N_19223,N_18110,N_18786);
nand U19224 (N_19224,N_18226,N_18980);
or U19225 (N_19225,N_18890,N_18739);
or U19226 (N_19226,N_18755,N_18506);
nor U19227 (N_19227,N_18961,N_18452);
and U19228 (N_19228,N_18230,N_18479);
xor U19229 (N_19229,N_18849,N_18586);
and U19230 (N_19230,N_18344,N_18435);
or U19231 (N_19231,N_18265,N_18319);
nor U19232 (N_19232,N_18658,N_18086);
nor U19233 (N_19233,N_18590,N_18523);
or U19234 (N_19234,N_18910,N_18638);
nand U19235 (N_19235,N_18408,N_18927);
and U19236 (N_19236,N_18194,N_18660);
nand U19237 (N_19237,N_18747,N_18215);
xor U19238 (N_19238,N_18477,N_18948);
nor U19239 (N_19239,N_18933,N_18828);
xnor U19240 (N_19240,N_18598,N_18119);
xnor U19241 (N_19241,N_18107,N_18117);
nor U19242 (N_19242,N_18484,N_18541);
nor U19243 (N_19243,N_18169,N_18356);
and U19244 (N_19244,N_18818,N_18651);
nand U19245 (N_19245,N_18080,N_18630);
or U19246 (N_19246,N_18981,N_18268);
nor U19247 (N_19247,N_18475,N_18769);
xor U19248 (N_19248,N_18063,N_18290);
and U19249 (N_19249,N_18072,N_18223);
nand U19250 (N_19250,N_18251,N_18277);
or U19251 (N_19251,N_18553,N_18882);
xnor U19252 (N_19252,N_18275,N_18515);
and U19253 (N_19253,N_18876,N_18654);
or U19254 (N_19254,N_18264,N_18990);
nand U19255 (N_19255,N_18663,N_18155);
and U19256 (N_19256,N_18205,N_18552);
or U19257 (N_19257,N_18497,N_18149);
nand U19258 (N_19258,N_18066,N_18998);
nor U19259 (N_19259,N_18420,N_18976);
xnor U19260 (N_19260,N_18104,N_18780);
nor U19261 (N_19261,N_18282,N_18625);
nor U19262 (N_19262,N_18217,N_18551);
xor U19263 (N_19263,N_18681,N_18841);
xor U19264 (N_19264,N_18603,N_18622);
nor U19265 (N_19265,N_18659,N_18700);
and U19266 (N_19266,N_18239,N_18560);
xor U19267 (N_19267,N_18443,N_18084);
or U19268 (N_19268,N_18147,N_18984);
and U19269 (N_19269,N_18904,N_18767);
xnor U19270 (N_19270,N_18255,N_18667);
and U19271 (N_19271,N_18683,N_18897);
and U19272 (N_19272,N_18219,N_18137);
nand U19273 (N_19273,N_18032,N_18301);
nand U19274 (N_19274,N_18090,N_18389);
nor U19275 (N_19275,N_18935,N_18533);
xor U19276 (N_19276,N_18711,N_18131);
nand U19277 (N_19277,N_18991,N_18498);
xor U19278 (N_19278,N_18664,N_18945);
and U19279 (N_19279,N_18752,N_18644);
nand U19280 (N_19280,N_18702,N_18323);
xnor U19281 (N_19281,N_18363,N_18177);
nand U19282 (N_19282,N_18626,N_18829);
nand U19283 (N_19283,N_18844,N_18256);
nor U19284 (N_19284,N_18287,N_18597);
xnor U19285 (N_19285,N_18861,N_18920);
xor U19286 (N_19286,N_18485,N_18317);
xor U19287 (N_19287,N_18838,N_18293);
or U19288 (N_19288,N_18810,N_18862);
or U19289 (N_19289,N_18837,N_18398);
and U19290 (N_19290,N_18947,N_18074);
nor U19291 (N_19291,N_18762,N_18023);
and U19292 (N_19292,N_18494,N_18253);
nand U19293 (N_19293,N_18511,N_18899);
nor U19294 (N_19294,N_18013,N_18977);
nand U19295 (N_19295,N_18097,N_18340);
or U19296 (N_19296,N_18191,N_18145);
nand U19297 (N_19297,N_18764,N_18160);
nor U19298 (N_19298,N_18463,N_18456);
xor U19299 (N_19299,N_18613,N_18534);
nand U19300 (N_19300,N_18181,N_18943);
and U19301 (N_19301,N_18480,N_18802);
nor U19302 (N_19302,N_18375,N_18207);
nand U19303 (N_19303,N_18554,N_18572);
or U19304 (N_19304,N_18153,N_18779);
nor U19305 (N_19305,N_18993,N_18092);
nor U19306 (N_19306,N_18873,N_18760);
xor U19307 (N_19307,N_18354,N_18851);
or U19308 (N_19308,N_18983,N_18116);
or U19309 (N_19309,N_18254,N_18111);
nand U19310 (N_19310,N_18279,N_18774);
and U19311 (N_19311,N_18649,N_18724);
and U19312 (N_19312,N_18870,N_18997);
xnor U19313 (N_19313,N_18628,N_18583);
nand U19314 (N_19314,N_18830,N_18388);
or U19315 (N_19315,N_18417,N_18887);
nor U19316 (N_19316,N_18605,N_18772);
xor U19317 (N_19317,N_18031,N_18364);
nand U19318 (N_19318,N_18527,N_18002);
xnor U19319 (N_19319,N_18179,N_18692);
and U19320 (N_19320,N_18472,N_18324);
xor U19321 (N_19321,N_18350,N_18715);
nand U19322 (N_19322,N_18380,N_18795);
or U19323 (N_19323,N_18721,N_18249);
and U19324 (N_19324,N_18695,N_18599);
nor U19325 (N_19325,N_18641,N_18895);
and U19326 (N_19326,N_18801,N_18517);
nand U19327 (N_19327,N_18336,N_18071);
and U19328 (N_19328,N_18788,N_18415);
nand U19329 (N_19329,N_18240,N_18315);
and U19330 (N_19330,N_18775,N_18513);
nor U19331 (N_19331,N_18989,N_18532);
nor U19332 (N_19332,N_18478,N_18258);
or U19333 (N_19333,N_18283,N_18091);
and U19334 (N_19334,N_18428,N_18833);
and U19335 (N_19335,N_18405,N_18921);
and U19336 (N_19336,N_18387,N_18791);
xor U19337 (N_19337,N_18733,N_18600);
xor U19338 (N_19338,N_18236,N_18835);
nand U19339 (N_19339,N_18061,N_18881);
or U19340 (N_19340,N_18765,N_18313);
nand U19341 (N_19341,N_18102,N_18422);
and U19342 (N_19342,N_18843,N_18034);
or U19343 (N_19343,N_18796,N_18224);
and U19344 (N_19344,N_18059,N_18220);
xnor U19345 (N_19345,N_18101,N_18812);
nand U19346 (N_19346,N_18633,N_18161);
nor U19347 (N_19347,N_18857,N_18940);
and U19348 (N_19348,N_18221,N_18100);
and U19349 (N_19349,N_18507,N_18822);
or U19350 (N_19350,N_18968,N_18957);
or U19351 (N_19351,N_18183,N_18783);
and U19352 (N_19352,N_18261,N_18051);
or U19353 (N_19353,N_18657,N_18369);
nor U19354 (N_19354,N_18376,N_18894);
and U19355 (N_19355,N_18811,N_18286);
xor U19356 (N_19356,N_18555,N_18799);
nor U19357 (N_19357,N_18907,N_18798);
and U19358 (N_19358,N_18856,N_18514);
nor U19359 (N_19359,N_18713,N_18306);
xnor U19360 (N_19360,N_18148,N_18806);
xnor U19361 (N_19361,N_18173,N_18141);
nand U19362 (N_19362,N_18418,N_18292);
xnor U19363 (N_19363,N_18007,N_18395);
xor U19364 (N_19364,N_18792,N_18751);
nor U19365 (N_19365,N_18893,N_18790);
nand U19366 (N_19366,N_18127,N_18170);
or U19367 (N_19367,N_18247,N_18166);
nor U19368 (N_19368,N_18073,N_18817);
nand U19369 (N_19369,N_18040,N_18394);
and U19370 (N_19370,N_18202,N_18687);
nor U19371 (N_19371,N_18726,N_18923);
or U19372 (N_19372,N_18492,N_18908);
nor U19373 (N_19373,N_18362,N_18146);
xor U19374 (N_19374,N_18471,N_18438);
nand U19375 (N_19375,N_18913,N_18234);
nor U19376 (N_19376,N_18030,N_18298);
and U19377 (N_19377,N_18307,N_18115);
and U19378 (N_19378,N_18383,N_18020);
xor U19379 (N_19379,N_18043,N_18746);
and U19380 (N_19380,N_18487,N_18869);
nor U19381 (N_19381,N_18805,N_18055);
nor U19382 (N_19382,N_18952,N_18912);
and U19383 (N_19383,N_18257,N_18209);
nor U19384 (N_19384,N_18858,N_18629);
and U19385 (N_19385,N_18813,N_18014);
xnor U19386 (N_19386,N_18486,N_18134);
or U19387 (N_19387,N_18573,N_18901);
nand U19388 (N_19388,N_18875,N_18963);
nor U19389 (N_19389,N_18691,N_18537);
or U19390 (N_19390,N_18204,N_18140);
xnor U19391 (N_19391,N_18266,N_18758);
xor U19392 (N_19392,N_18820,N_18757);
and U19393 (N_19393,N_18536,N_18520);
and U19394 (N_19394,N_18330,N_18510);
nand U19395 (N_19395,N_18847,N_18675);
nor U19396 (N_19396,N_18589,N_18154);
or U19397 (N_19397,N_18879,N_18449);
and U19398 (N_19398,N_18114,N_18093);
and U19399 (N_19399,N_18409,N_18850);
and U19400 (N_19400,N_18609,N_18761);
xor U19401 (N_19401,N_18909,N_18748);
xnor U19402 (N_19402,N_18530,N_18132);
nand U19403 (N_19403,N_18714,N_18522);
or U19404 (N_19404,N_18954,N_18425);
or U19405 (N_19405,N_18270,N_18880);
nor U19406 (N_19406,N_18491,N_18680);
xnor U19407 (N_19407,N_18060,N_18371);
nand U19408 (N_19408,N_18122,N_18971);
xnor U19409 (N_19409,N_18175,N_18296);
and U19410 (N_19410,N_18703,N_18777);
nor U19411 (N_19411,N_18544,N_18348);
and U19412 (N_19412,N_18036,N_18067);
and U19413 (N_19413,N_18677,N_18151);
or U19414 (N_19414,N_18610,N_18591);
or U19415 (N_19415,N_18735,N_18446);
and U19416 (N_19416,N_18000,N_18526);
and U19417 (N_19417,N_18004,N_18267);
or U19418 (N_19418,N_18969,N_18225);
nand U19419 (N_19419,N_18819,N_18891);
xnor U19420 (N_19420,N_18604,N_18430);
and U19421 (N_19421,N_18281,N_18815);
or U19422 (N_19422,N_18546,N_18391);
and U19423 (N_19423,N_18548,N_18878);
or U19424 (N_19424,N_18662,N_18787);
xnor U19425 (N_19425,N_18707,N_18953);
nand U19426 (N_19426,N_18187,N_18346);
nand U19427 (N_19427,N_18964,N_18898);
or U19428 (N_19428,N_18508,N_18580);
nand U19429 (N_19429,N_18144,N_18174);
nand U19430 (N_19430,N_18188,N_18402);
and U19431 (N_19431,N_18974,N_18423);
nand U19432 (N_19432,N_18026,N_18646);
or U19433 (N_19433,N_18305,N_18561);
xor U19434 (N_19434,N_18126,N_18623);
xnor U19435 (N_19435,N_18693,N_18335);
and U19436 (N_19436,N_18406,N_18150);
and U19437 (N_19437,N_18178,N_18334);
or U19438 (N_19438,N_18218,N_18525);
xor U19439 (N_19439,N_18621,N_18512);
nor U19440 (N_19440,N_18624,N_18738);
nand U19441 (N_19441,N_18883,N_18046);
and U19442 (N_19442,N_18579,N_18039);
and U19443 (N_19443,N_18469,N_18595);
and U19444 (N_19444,N_18351,N_18979);
or U19445 (N_19445,N_18612,N_18694);
nor U19446 (N_19446,N_18717,N_18333);
xnor U19447 (N_19447,N_18196,N_18759);
nand U19448 (N_19448,N_18269,N_18800);
nor U19449 (N_19449,N_18889,N_18118);
and U19450 (N_19450,N_18670,N_18377);
xnor U19451 (N_19451,N_18570,N_18696);
or U19452 (N_19452,N_18197,N_18959);
xnor U19453 (N_19453,N_18793,N_18010);
or U19454 (N_19454,N_18203,N_18042);
nand U19455 (N_19455,N_18331,N_18347);
and U19456 (N_19456,N_18571,N_18049);
or U19457 (N_19457,N_18358,N_18158);
xnor U19458 (N_19458,N_18085,N_18785);
nand U19459 (N_19459,N_18996,N_18932);
xnor U19460 (N_19460,N_18326,N_18005);
and U19461 (N_19461,N_18743,N_18653);
xor U19462 (N_19462,N_18352,N_18636);
nand U19463 (N_19463,N_18686,N_18022);
xnor U19464 (N_19464,N_18906,N_18189);
nand U19465 (N_19465,N_18088,N_18956);
nand U19466 (N_19466,N_18753,N_18271);
nor U19467 (N_19467,N_18495,N_18865);
xnor U19468 (N_19468,N_18343,N_18937);
or U19469 (N_19469,N_18138,N_18349);
nand U19470 (N_19470,N_18041,N_18439);
xnor U19471 (N_19471,N_18581,N_18434);
nand U19472 (N_19472,N_18033,N_18575);
and U19473 (N_19473,N_18965,N_18958);
or U19474 (N_19474,N_18052,N_18466);
nor U19475 (N_19475,N_18557,N_18442);
nand U19476 (N_19476,N_18365,N_18473);
and U19477 (N_19477,N_18917,N_18245);
nand U19478 (N_19478,N_18099,N_18831);
nor U19479 (N_19479,N_18559,N_18550);
or U19480 (N_19480,N_18637,N_18794);
xnor U19481 (N_19481,N_18441,N_18105);
and U19482 (N_19482,N_18057,N_18069);
nand U19483 (N_19483,N_18021,N_18206);
xor U19484 (N_19484,N_18539,N_18400);
or U19485 (N_19485,N_18942,N_18688);
nor U19486 (N_19486,N_18992,N_18924);
or U19487 (N_19487,N_18941,N_18727);
nor U19488 (N_19488,N_18709,N_18241);
and U19489 (N_19489,N_18125,N_18655);
nor U19490 (N_19490,N_18095,N_18926);
and U19491 (N_19491,N_18987,N_18044);
xor U19492 (N_19492,N_18045,N_18648);
or U19493 (N_19493,N_18524,N_18056);
nand U19494 (N_19494,N_18698,N_18341);
and U19495 (N_19495,N_18647,N_18602);
nor U19496 (N_19496,N_18499,N_18433);
or U19497 (N_19497,N_18303,N_18601);
nor U19498 (N_19498,N_18208,N_18928);
xnor U19499 (N_19499,N_18627,N_18053);
nor U19500 (N_19500,N_18883,N_18097);
xor U19501 (N_19501,N_18685,N_18359);
xnor U19502 (N_19502,N_18294,N_18434);
nor U19503 (N_19503,N_18311,N_18000);
and U19504 (N_19504,N_18708,N_18539);
or U19505 (N_19505,N_18822,N_18860);
nand U19506 (N_19506,N_18348,N_18901);
nor U19507 (N_19507,N_18828,N_18329);
xor U19508 (N_19508,N_18059,N_18020);
nand U19509 (N_19509,N_18704,N_18604);
nor U19510 (N_19510,N_18204,N_18989);
nand U19511 (N_19511,N_18259,N_18707);
and U19512 (N_19512,N_18569,N_18245);
xnor U19513 (N_19513,N_18806,N_18620);
nand U19514 (N_19514,N_18698,N_18126);
or U19515 (N_19515,N_18319,N_18855);
nor U19516 (N_19516,N_18709,N_18374);
nor U19517 (N_19517,N_18401,N_18603);
and U19518 (N_19518,N_18012,N_18101);
or U19519 (N_19519,N_18737,N_18320);
or U19520 (N_19520,N_18197,N_18259);
and U19521 (N_19521,N_18443,N_18801);
and U19522 (N_19522,N_18754,N_18090);
and U19523 (N_19523,N_18767,N_18119);
nor U19524 (N_19524,N_18770,N_18254);
nor U19525 (N_19525,N_18887,N_18425);
nor U19526 (N_19526,N_18713,N_18299);
nor U19527 (N_19527,N_18950,N_18339);
xor U19528 (N_19528,N_18711,N_18709);
xor U19529 (N_19529,N_18003,N_18832);
or U19530 (N_19530,N_18147,N_18081);
or U19531 (N_19531,N_18060,N_18186);
and U19532 (N_19532,N_18342,N_18735);
xnor U19533 (N_19533,N_18153,N_18240);
nand U19534 (N_19534,N_18826,N_18963);
nor U19535 (N_19535,N_18586,N_18710);
nor U19536 (N_19536,N_18841,N_18217);
xnor U19537 (N_19537,N_18675,N_18707);
or U19538 (N_19538,N_18137,N_18469);
or U19539 (N_19539,N_18443,N_18308);
or U19540 (N_19540,N_18998,N_18575);
nor U19541 (N_19541,N_18703,N_18715);
and U19542 (N_19542,N_18149,N_18034);
nor U19543 (N_19543,N_18366,N_18497);
xnor U19544 (N_19544,N_18366,N_18382);
or U19545 (N_19545,N_18965,N_18226);
nand U19546 (N_19546,N_18583,N_18744);
nor U19547 (N_19547,N_18352,N_18429);
and U19548 (N_19548,N_18735,N_18725);
nand U19549 (N_19549,N_18399,N_18842);
nor U19550 (N_19550,N_18734,N_18897);
nand U19551 (N_19551,N_18793,N_18360);
xnor U19552 (N_19552,N_18497,N_18119);
xnor U19553 (N_19553,N_18301,N_18349);
nor U19554 (N_19554,N_18713,N_18240);
nand U19555 (N_19555,N_18467,N_18968);
nor U19556 (N_19556,N_18939,N_18079);
and U19557 (N_19557,N_18087,N_18104);
xnor U19558 (N_19558,N_18880,N_18207);
or U19559 (N_19559,N_18369,N_18992);
nand U19560 (N_19560,N_18346,N_18199);
and U19561 (N_19561,N_18561,N_18856);
xor U19562 (N_19562,N_18330,N_18393);
and U19563 (N_19563,N_18809,N_18640);
and U19564 (N_19564,N_18343,N_18371);
or U19565 (N_19565,N_18930,N_18861);
xor U19566 (N_19566,N_18321,N_18246);
xor U19567 (N_19567,N_18068,N_18570);
nand U19568 (N_19568,N_18112,N_18650);
nor U19569 (N_19569,N_18586,N_18838);
and U19570 (N_19570,N_18905,N_18377);
nor U19571 (N_19571,N_18816,N_18825);
nand U19572 (N_19572,N_18576,N_18470);
or U19573 (N_19573,N_18129,N_18037);
or U19574 (N_19574,N_18451,N_18247);
or U19575 (N_19575,N_18097,N_18795);
or U19576 (N_19576,N_18886,N_18027);
and U19577 (N_19577,N_18974,N_18498);
xnor U19578 (N_19578,N_18186,N_18199);
nor U19579 (N_19579,N_18813,N_18134);
nand U19580 (N_19580,N_18763,N_18384);
xnor U19581 (N_19581,N_18852,N_18605);
xnor U19582 (N_19582,N_18574,N_18827);
and U19583 (N_19583,N_18077,N_18005);
nor U19584 (N_19584,N_18465,N_18674);
or U19585 (N_19585,N_18676,N_18906);
nor U19586 (N_19586,N_18308,N_18195);
nand U19587 (N_19587,N_18194,N_18391);
xor U19588 (N_19588,N_18821,N_18100);
or U19589 (N_19589,N_18350,N_18874);
nand U19590 (N_19590,N_18367,N_18529);
nor U19591 (N_19591,N_18280,N_18635);
nor U19592 (N_19592,N_18988,N_18424);
nand U19593 (N_19593,N_18186,N_18320);
xor U19594 (N_19594,N_18613,N_18866);
xor U19595 (N_19595,N_18696,N_18714);
nand U19596 (N_19596,N_18183,N_18707);
and U19597 (N_19597,N_18914,N_18105);
nor U19598 (N_19598,N_18533,N_18807);
or U19599 (N_19599,N_18694,N_18723);
and U19600 (N_19600,N_18510,N_18959);
and U19601 (N_19601,N_18709,N_18730);
or U19602 (N_19602,N_18315,N_18060);
nand U19603 (N_19603,N_18571,N_18566);
xor U19604 (N_19604,N_18578,N_18241);
or U19605 (N_19605,N_18982,N_18331);
nor U19606 (N_19606,N_18278,N_18474);
nand U19607 (N_19607,N_18855,N_18139);
and U19608 (N_19608,N_18669,N_18864);
and U19609 (N_19609,N_18313,N_18540);
nor U19610 (N_19610,N_18453,N_18797);
nand U19611 (N_19611,N_18503,N_18244);
and U19612 (N_19612,N_18417,N_18938);
or U19613 (N_19613,N_18830,N_18060);
or U19614 (N_19614,N_18160,N_18351);
xnor U19615 (N_19615,N_18101,N_18202);
or U19616 (N_19616,N_18267,N_18166);
xnor U19617 (N_19617,N_18199,N_18482);
xnor U19618 (N_19618,N_18977,N_18008);
and U19619 (N_19619,N_18137,N_18045);
nand U19620 (N_19620,N_18337,N_18690);
or U19621 (N_19621,N_18728,N_18371);
and U19622 (N_19622,N_18091,N_18030);
or U19623 (N_19623,N_18323,N_18559);
xnor U19624 (N_19624,N_18709,N_18903);
xnor U19625 (N_19625,N_18111,N_18424);
or U19626 (N_19626,N_18149,N_18595);
nor U19627 (N_19627,N_18803,N_18660);
or U19628 (N_19628,N_18466,N_18020);
and U19629 (N_19629,N_18101,N_18330);
or U19630 (N_19630,N_18572,N_18722);
or U19631 (N_19631,N_18306,N_18699);
nand U19632 (N_19632,N_18310,N_18371);
or U19633 (N_19633,N_18149,N_18305);
xnor U19634 (N_19634,N_18783,N_18965);
xnor U19635 (N_19635,N_18329,N_18719);
nor U19636 (N_19636,N_18191,N_18469);
and U19637 (N_19637,N_18648,N_18917);
nor U19638 (N_19638,N_18691,N_18203);
nor U19639 (N_19639,N_18789,N_18026);
nand U19640 (N_19640,N_18795,N_18204);
xnor U19641 (N_19641,N_18577,N_18051);
or U19642 (N_19642,N_18498,N_18307);
and U19643 (N_19643,N_18251,N_18362);
nand U19644 (N_19644,N_18973,N_18799);
and U19645 (N_19645,N_18195,N_18068);
xnor U19646 (N_19646,N_18949,N_18002);
nand U19647 (N_19647,N_18238,N_18899);
nor U19648 (N_19648,N_18046,N_18685);
xor U19649 (N_19649,N_18202,N_18236);
nor U19650 (N_19650,N_18681,N_18307);
nor U19651 (N_19651,N_18709,N_18161);
nor U19652 (N_19652,N_18220,N_18819);
and U19653 (N_19653,N_18080,N_18013);
xor U19654 (N_19654,N_18150,N_18333);
or U19655 (N_19655,N_18981,N_18466);
xor U19656 (N_19656,N_18454,N_18921);
nor U19657 (N_19657,N_18092,N_18001);
nand U19658 (N_19658,N_18731,N_18307);
or U19659 (N_19659,N_18489,N_18850);
and U19660 (N_19660,N_18676,N_18562);
xnor U19661 (N_19661,N_18274,N_18890);
nand U19662 (N_19662,N_18914,N_18278);
and U19663 (N_19663,N_18898,N_18698);
and U19664 (N_19664,N_18397,N_18915);
or U19665 (N_19665,N_18921,N_18052);
nand U19666 (N_19666,N_18927,N_18097);
xnor U19667 (N_19667,N_18577,N_18015);
nor U19668 (N_19668,N_18774,N_18708);
nor U19669 (N_19669,N_18265,N_18190);
and U19670 (N_19670,N_18746,N_18412);
and U19671 (N_19671,N_18043,N_18342);
nor U19672 (N_19672,N_18296,N_18945);
or U19673 (N_19673,N_18613,N_18090);
or U19674 (N_19674,N_18037,N_18293);
nor U19675 (N_19675,N_18503,N_18970);
nand U19676 (N_19676,N_18585,N_18530);
and U19677 (N_19677,N_18504,N_18522);
nor U19678 (N_19678,N_18298,N_18144);
or U19679 (N_19679,N_18835,N_18851);
nand U19680 (N_19680,N_18139,N_18118);
nand U19681 (N_19681,N_18392,N_18529);
and U19682 (N_19682,N_18327,N_18556);
xor U19683 (N_19683,N_18849,N_18653);
and U19684 (N_19684,N_18804,N_18910);
and U19685 (N_19685,N_18832,N_18974);
and U19686 (N_19686,N_18580,N_18063);
and U19687 (N_19687,N_18405,N_18815);
and U19688 (N_19688,N_18368,N_18361);
nor U19689 (N_19689,N_18357,N_18721);
or U19690 (N_19690,N_18219,N_18979);
and U19691 (N_19691,N_18673,N_18134);
and U19692 (N_19692,N_18058,N_18624);
nand U19693 (N_19693,N_18693,N_18684);
nand U19694 (N_19694,N_18260,N_18467);
nand U19695 (N_19695,N_18435,N_18429);
and U19696 (N_19696,N_18594,N_18586);
or U19697 (N_19697,N_18025,N_18824);
nor U19698 (N_19698,N_18166,N_18522);
or U19699 (N_19699,N_18815,N_18414);
and U19700 (N_19700,N_18341,N_18464);
and U19701 (N_19701,N_18758,N_18631);
xnor U19702 (N_19702,N_18827,N_18264);
and U19703 (N_19703,N_18620,N_18443);
and U19704 (N_19704,N_18020,N_18019);
or U19705 (N_19705,N_18390,N_18035);
or U19706 (N_19706,N_18038,N_18482);
nand U19707 (N_19707,N_18787,N_18163);
nor U19708 (N_19708,N_18214,N_18808);
nand U19709 (N_19709,N_18709,N_18590);
xor U19710 (N_19710,N_18014,N_18798);
and U19711 (N_19711,N_18155,N_18008);
or U19712 (N_19712,N_18061,N_18829);
or U19713 (N_19713,N_18079,N_18993);
nand U19714 (N_19714,N_18384,N_18785);
nand U19715 (N_19715,N_18533,N_18230);
nand U19716 (N_19716,N_18385,N_18265);
and U19717 (N_19717,N_18439,N_18846);
and U19718 (N_19718,N_18293,N_18786);
or U19719 (N_19719,N_18254,N_18496);
and U19720 (N_19720,N_18842,N_18088);
xor U19721 (N_19721,N_18496,N_18187);
xor U19722 (N_19722,N_18031,N_18567);
or U19723 (N_19723,N_18475,N_18879);
nand U19724 (N_19724,N_18376,N_18074);
nand U19725 (N_19725,N_18054,N_18704);
and U19726 (N_19726,N_18748,N_18794);
nor U19727 (N_19727,N_18484,N_18480);
or U19728 (N_19728,N_18516,N_18428);
xor U19729 (N_19729,N_18268,N_18104);
nand U19730 (N_19730,N_18922,N_18011);
nor U19731 (N_19731,N_18548,N_18297);
xnor U19732 (N_19732,N_18224,N_18254);
nor U19733 (N_19733,N_18363,N_18069);
and U19734 (N_19734,N_18543,N_18013);
xnor U19735 (N_19735,N_18198,N_18686);
xor U19736 (N_19736,N_18364,N_18700);
xnor U19737 (N_19737,N_18222,N_18870);
nand U19738 (N_19738,N_18747,N_18837);
and U19739 (N_19739,N_18190,N_18322);
nand U19740 (N_19740,N_18718,N_18356);
xnor U19741 (N_19741,N_18974,N_18375);
xnor U19742 (N_19742,N_18294,N_18573);
and U19743 (N_19743,N_18197,N_18807);
nand U19744 (N_19744,N_18713,N_18801);
or U19745 (N_19745,N_18802,N_18934);
nor U19746 (N_19746,N_18609,N_18760);
or U19747 (N_19747,N_18823,N_18254);
and U19748 (N_19748,N_18434,N_18598);
nor U19749 (N_19749,N_18265,N_18484);
or U19750 (N_19750,N_18027,N_18763);
nor U19751 (N_19751,N_18096,N_18836);
or U19752 (N_19752,N_18954,N_18953);
xnor U19753 (N_19753,N_18167,N_18949);
nor U19754 (N_19754,N_18571,N_18300);
xnor U19755 (N_19755,N_18753,N_18298);
xnor U19756 (N_19756,N_18303,N_18084);
nand U19757 (N_19757,N_18960,N_18780);
nand U19758 (N_19758,N_18480,N_18495);
nor U19759 (N_19759,N_18957,N_18858);
or U19760 (N_19760,N_18569,N_18747);
nand U19761 (N_19761,N_18602,N_18233);
nor U19762 (N_19762,N_18933,N_18636);
xor U19763 (N_19763,N_18209,N_18206);
nand U19764 (N_19764,N_18557,N_18156);
or U19765 (N_19765,N_18524,N_18895);
or U19766 (N_19766,N_18921,N_18097);
xnor U19767 (N_19767,N_18893,N_18788);
nor U19768 (N_19768,N_18996,N_18257);
xnor U19769 (N_19769,N_18269,N_18198);
and U19770 (N_19770,N_18767,N_18303);
nor U19771 (N_19771,N_18422,N_18515);
or U19772 (N_19772,N_18343,N_18672);
xnor U19773 (N_19773,N_18522,N_18913);
xnor U19774 (N_19774,N_18332,N_18497);
or U19775 (N_19775,N_18133,N_18780);
xor U19776 (N_19776,N_18173,N_18431);
nor U19777 (N_19777,N_18895,N_18441);
nand U19778 (N_19778,N_18874,N_18876);
and U19779 (N_19779,N_18001,N_18808);
and U19780 (N_19780,N_18848,N_18420);
or U19781 (N_19781,N_18825,N_18812);
nand U19782 (N_19782,N_18833,N_18781);
nand U19783 (N_19783,N_18195,N_18950);
xor U19784 (N_19784,N_18465,N_18534);
or U19785 (N_19785,N_18927,N_18489);
nor U19786 (N_19786,N_18528,N_18055);
nand U19787 (N_19787,N_18705,N_18671);
nand U19788 (N_19788,N_18261,N_18792);
nor U19789 (N_19789,N_18710,N_18792);
nor U19790 (N_19790,N_18273,N_18970);
nor U19791 (N_19791,N_18670,N_18767);
or U19792 (N_19792,N_18171,N_18879);
xor U19793 (N_19793,N_18999,N_18127);
or U19794 (N_19794,N_18968,N_18186);
and U19795 (N_19795,N_18576,N_18585);
nor U19796 (N_19796,N_18942,N_18176);
and U19797 (N_19797,N_18301,N_18225);
nor U19798 (N_19798,N_18512,N_18904);
or U19799 (N_19799,N_18617,N_18657);
xor U19800 (N_19800,N_18095,N_18709);
or U19801 (N_19801,N_18864,N_18578);
nor U19802 (N_19802,N_18724,N_18743);
or U19803 (N_19803,N_18784,N_18276);
xnor U19804 (N_19804,N_18580,N_18072);
nand U19805 (N_19805,N_18773,N_18554);
or U19806 (N_19806,N_18932,N_18921);
and U19807 (N_19807,N_18105,N_18134);
nand U19808 (N_19808,N_18602,N_18464);
nor U19809 (N_19809,N_18661,N_18969);
nand U19810 (N_19810,N_18275,N_18046);
xnor U19811 (N_19811,N_18264,N_18768);
nand U19812 (N_19812,N_18288,N_18336);
and U19813 (N_19813,N_18024,N_18136);
xnor U19814 (N_19814,N_18812,N_18770);
or U19815 (N_19815,N_18227,N_18220);
xnor U19816 (N_19816,N_18478,N_18293);
xor U19817 (N_19817,N_18889,N_18978);
xor U19818 (N_19818,N_18620,N_18204);
and U19819 (N_19819,N_18960,N_18653);
xnor U19820 (N_19820,N_18824,N_18918);
nand U19821 (N_19821,N_18296,N_18696);
xnor U19822 (N_19822,N_18911,N_18056);
and U19823 (N_19823,N_18240,N_18526);
or U19824 (N_19824,N_18187,N_18819);
xor U19825 (N_19825,N_18096,N_18751);
nand U19826 (N_19826,N_18888,N_18999);
xor U19827 (N_19827,N_18337,N_18208);
xnor U19828 (N_19828,N_18829,N_18955);
xnor U19829 (N_19829,N_18065,N_18466);
xor U19830 (N_19830,N_18879,N_18443);
nand U19831 (N_19831,N_18277,N_18441);
and U19832 (N_19832,N_18104,N_18570);
or U19833 (N_19833,N_18872,N_18108);
nor U19834 (N_19834,N_18550,N_18119);
nand U19835 (N_19835,N_18199,N_18103);
and U19836 (N_19836,N_18396,N_18202);
xor U19837 (N_19837,N_18385,N_18143);
xnor U19838 (N_19838,N_18987,N_18817);
and U19839 (N_19839,N_18355,N_18870);
or U19840 (N_19840,N_18466,N_18298);
or U19841 (N_19841,N_18495,N_18121);
or U19842 (N_19842,N_18042,N_18529);
or U19843 (N_19843,N_18849,N_18830);
xor U19844 (N_19844,N_18013,N_18955);
xnor U19845 (N_19845,N_18998,N_18356);
nand U19846 (N_19846,N_18613,N_18569);
nand U19847 (N_19847,N_18946,N_18700);
nor U19848 (N_19848,N_18048,N_18935);
xor U19849 (N_19849,N_18836,N_18141);
xnor U19850 (N_19850,N_18379,N_18857);
xor U19851 (N_19851,N_18834,N_18114);
and U19852 (N_19852,N_18610,N_18249);
nor U19853 (N_19853,N_18727,N_18301);
or U19854 (N_19854,N_18665,N_18541);
nand U19855 (N_19855,N_18617,N_18317);
and U19856 (N_19856,N_18643,N_18959);
or U19857 (N_19857,N_18096,N_18589);
or U19858 (N_19858,N_18459,N_18200);
nor U19859 (N_19859,N_18778,N_18986);
or U19860 (N_19860,N_18456,N_18621);
nor U19861 (N_19861,N_18791,N_18026);
nor U19862 (N_19862,N_18467,N_18392);
nand U19863 (N_19863,N_18271,N_18907);
nand U19864 (N_19864,N_18714,N_18290);
and U19865 (N_19865,N_18067,N_18033);
and U19866 (N_19866,N_18334,N_18357);
nor U19867 (N_19867,N_18136,N_18924);
nand U19868 (N_19868,N_18894,N_18230);
or U19869 (N_19869,N_18230,N_18981);
nor U19870 (N_19870,N_18169,N_18272);
nor U19871 (N_19871,N_18241,N_18633);
nor U19872 (N_19872,N_18184,N_18101);
nor U19873 (N_19873,N_18844,N_18705);
nand U19874 (N_19874,N_18369,N_18913);
nand U19875 (N_19875,N_18226,N_18791);
or U19876 (N_19876,N_18259,N_18455);
and U19877 (N_19877,N_18672,N_18328);
xnor U19878 (N_19878,N_18891,N_18282);
xnor U19879 (N_19879,N_18666,N_18677);
nand U19880 (N_19880,N_18589,N_18360);
nor U19881 (N_19881,N_18255,N_18946);
and U19882 (N_19882,N_18355,N_18038);
nand U19883 (N_19883,N_18637,N_18734);
nand U19884 (N_19884,N_18668,N_18563);
or U19885 (N_19885,N_18258,N_18244);
nor U19886 (N_19886,N_18760,N_18571);
and U19887 (N_19887,N_18824,N_18542);
and U19888 (N_19888,N_18886,N_18518);
nor U19889 (N_19889,N_18044,N_18654);
nand U19890 (N_19890,N_18974,N_18092);
nor U19891 (N_19891,N_18537,N_18149);
xor U19892 (N_19892,N_18942,N_18597);
xnor U19893 (N_19893,N_18867,N_18828);
or U19894 (N_19894,N_18615,N_18305);
and U19895 (N_19895,N_18064,N_18402);
xor U19896 (N_19896,N_18151,N_18737);
nor U19897 (N_19897,N_18224,N_18492);
or U19898 (N_19898,N_18153,N_18262);
xnor U19899 (N_19899,N_18118,N_18125);
nor U19900 (N_19900,N_18941,N_18758);
or U19901 (N_19901,N_18299,N_18282);
xnor U19902 (N_19902,N_18925,N_18175);
or U19903 (N_19903,N_18017,N_18128);
nor U19904 (N_19904,N_18228,N_18764);
xnor U19905 (N_19905,N_18110,N_18448);
or U19906 (N_19906,N_18683,N_18428);
xnor U19907 (N_19907,N_18700,N_18497);
and U19908 (N_19908,N_18767,N_18745);
or U19909 (N_19909,N_18504,N_18059);
xnor U19910 (N_19910,N_18284,N_18683);
xor U19911 (N_19911,N_18310,N_18479);
nand U19912 (N_19912,N_18013,N_18390);
or U19913 (N_19913,N_18667,N_18908);
or U19914 (N_19914,N_18887,N_18227);
and U19915 (N_19915,N_18797,N_18026);
xnor U19916 (N_19916,N_18285,N_18162);
and U19917 (N_19917,N_18446,N_18522);
and U19918 (N_19918,N_18339,N_18661);
xnor U19919 (N_19919,N_18166,N_18490);
nand U19920 (N_19920,N_18688,N_18608);
nand U19921 (N_19921,N_18098,N_18230);
xnor U19922 (N_19922,N_18911,N_18110);
or U19923 (N_19923,N_18143,N_18214);
nand U19924 (N_19924,N_18500,N_18781);
and U19925 (N_19925,N_18398,N_18073);
and U19926 (N_19926,N_18815,N_18698);
nor U19927 (N_19927,N_18592,N_18525);
nand U19928 (N_19928,N_18048,N_18186);
and U19929 (N_19929,N_18906,N_18528);
nand U19930 (N_19930,N_18681,N_18569);
and U19931 (N_19931,N_18434,N_18105);
nand U19932 (N_19932,N_18222,N_18286);
or U19933 (N_19933,N_18366,N_18249);
or U19934 (N_19934,N_18899,N_18482);
and U19935 (N_19935,N_18284,N_18280);
or U19936 (N_19936,N_18955,N_18681);
or U19937 (N_19937,N_18349,N_18303);
nor U19938 (N_19938,N_18491,N_18060);
xnor U19939 (N_19939,N_18776,N_18710);
xor U19940 (N_19940,N_18050,N_18789);
nand U19941 (N_19941,N_18938,N_18249);
nand U19942 (N_19942,N_18489,N_18727);
nor U19943 (N_19943,N_18567,N_18456);
nand U19944 (N_19944,N_18088,N_18324);
nor U19945 (N_19945,N_18675,N_18225);
nor U19946 (N_19946,N_18865,N_18332);
nand U19947 (N_19947,N_18784,N_18586);
and U19948 (N_19948,N_18493,N_18172);
nand U19949 (N_19949,N_18397,N_18603);
and U19950 (N_19950,N_18866,N_18633);
nand U19951 (N_19951,N_18680,N_18451);
and U19952 (N_19952,N_18995,N_18526);
nand U19953 (N_19953,N_18028,N_18278);
xor U19954 (N_19954,N_18797,N_18521);
or U19955 (N_19955,N_18948,N_18509);
xor U19956 (N_19956,N_18048,N_18191);
or U19957 (N_19957,N_18526,N_18673);
nor U19958 (N_19958,N_18340,N_18124);
or U19959 (N_19959,N_18667,N_18453);
xnor U19960 (N_19960,N_18031,N_18113);
nand U19961 (N_19961,N_18899,N_18981);
xor U19962 (N_19962,N_18669,N_18356);
or U19963 (N_19963,N_18304,N_18661);
or U19964 (N_19964,N_18670,N_18333);
xnor U19965 (N_19965,N_18667,N_18503);
nand U19966 (N_19966,N_18296,N_18022);
and U19967 (N_19967,N_18113,N_18894);
nor U19968 (N_19968,N_18011,N_18970);
and U19969 (N_19969,N_18489,N_18550);
nor U19970 (N_19970,N_18314,N_18443);
and U19971 (N_19971,N_18003,N_18260);
xor U19972 (N_19972,N_18313,N_18243);
or U19973 (N_19973,N_18029,N_18130);
and U19974 (N_19974,N_18370,N_18768);
and U19975 (N_19975,N_18036,N_18693);
and U19976 (N_19976,N_18600,N_18952);
or U19977 (N_19977,N_18016,N_18398);
and U19978 (N_19978,N_18834,N_18488);
or U19979 (N_19979,N_18551,N_18956);
or U19980 (N_19980,N_18167,N_18804);
or U19981 (N_19981,N_18015,N_18393);
nor U19982 (N_19982,N_18586,N_18139);
xnor U19983 (N_19983,N_18240,N_18084);
xor U19984 (N_19984,N_18767,N_18302);
or U19985 (N_19985,N_18062,N_18238);
nor U19986 (N_19986,N_18978,N_18977);
nand U19987 (N_19987,N_18578,N_18555);
nand U19988 (N_19988,N_18486,N_18015);
and U19989 (N_19989,N_18706,N_18310);
nand U19990 (N_19990,N_18516,N_18180);
nor U19991 (N_19991,N_18800,N_18907);
and U19992 (N_19992,N_18727,N_18908);
and U19993 (N_19993,N_18294,N_18307);
nor U19994 (N_19994,N_18130,N_18495);
nor U19995 (N_19995,N_18016,N_18365);
or U19996 (N_19996,N_18289,N_18698);
and U19997 (N_19997,N_18322,N_18111);
or U19998 (N_19998,N_18177,N_18843);
nand U19999 (N_19999,N_18423,N_18522);
xnor U20000 (N_20000,N_19562,N_19108);
xnor U20001 (N_20001,N_19567,N_19252);
and U20002 (N_20002,N_19584,N_19370);
nand U20003 (N_20003,N_19468,N_19564);
or U20004 (N_20004,N_19844,N_19967);
and U20005 (N_20005,N_19217,N_19080);
and U20006 (N_20006,N_19923,N_19426);
and U20007 (N_20007,N_19524,N_19183);
or U20008 (N_20008,N_19433,N_19409);
xnor U20009 (N_20009,N_19750,N_19385);
or U20010 (N_20010,N_19261,N_19737);
and U20011 (N_20011,N_19942,N_19281);
xor U20012 (N_20012,N_19479,N_19194);
and U20013 (N_20013,N_19911,N_19098);
nor U20014 (N_20014,N_19420,N_19044);
or U20015 (N_20015,N_19221,N_19554);
xor U20016 (N_20016,N_19587,N_19401);
or U20017 (N_20017,N_19561,N_19984);
nand U20018 (N_20018,N_19971,N_19542);
nand U20019 (N_20019,N_19403,N_19817);
or U20020 (N_20020,N_19376,N_19444);
and U20021 (N_20021,N_19248,N_19665);
nand U20022 (N_20022,N_19886,N_19210);
and U20023 (N_20023,N_19769,N_19768);
nor U20024 (N_20024,N_19241,N_19075);
and U20025 (N_20025,N_19621,N_19849);
or U20026 (N_20026,N_19135,N_19094);
and U20027 (N_20027,N_19440,N_19400);
nor U20028 (N_20028,N_19880,N_19710);
nor U20029 (N_20029,N_19583,N_19349);
nand U20030 (N_20030,N_19458,N_19371);
nand U20031 (N_20031,N_19498,N_19841);
and U20032 (N_20032,N_19311,N_19117);
and U20033 (N_20033,N_19560,N_19472);
nand U20034 (N_20034,N_19027,N_19720);
xor U20035 (N_20035,N_19136,N_19480);
or U20036 (N_20036,N_19619,N_19388);
xnor U20037 (N_20037,N_19436,N_19973);
or U20038 (N_20038,N_19744,N_19302);
xnor U20039 (N_20039,N_19758,N_19794);
and U20040 (N_20040,N_19310,N_19660);
and U20041 (N_20041,N_19211,N_19839);
and U20042 (N_20042,N_19188,N_19414);
xor U20043 (N_20043,N_19539,N_19432);
or U20044 (N_20044,N_19642,N_19446);
nand U20045 (N_20045,N_19452,N_19378);
or U20046 (N_20046,N_19674,N_19305);
xnor U20047 (N_20047,N_19990,N_19928);
nor U20048 (N_20048,N_19068,N_19050);
nor U20049 (N_20049,N_19791,N_19303);
or U20050 (N_20050,N_19258,N_19919);
nor U20051 (N_20051,N_19995,N_19058);
nor U20052 (N_20052,N_19566,N_19986);
or U20053 (N_20053,N_19657,N_19792);
or U20054 (N_20054,N_19755,N_19507);
nor U20055 (N_20055,N_19353,N_19778);
or U20056 (N_20056,N_19515,N_19502);
nand U20057 (N_20057,N_19228,N_19447);
or U20058 (N_20058,N_19394,N_19474);
xnor U20059 (N_20059,N_19666,N_19010);
or U20060 (N_20060,N_19042,N_19985);
nor U20061 (N_20061,N_19589,N_19127);
or U20062 (N_20062,N_19115,N_19121);
and U20063 (N_20063,N_19675,N_19932);
and U20064 (N_20064,N_19918,N_19785);
xor U20065 (N_20065,N_19910,N_19213);
and U20066 (N_20066,N_19784,N_19585);
and U20067 (N_20067,N_19826,N_19280);
nand U20068 (N_20068,N_19747,N_19611);
or U20069 (N_20069,N_19150,N_19586);
nor U20070 (N_20070,N_19391,N_19820);
nand U20071 (N_20071,N_19837,N_19952);
or U20072 (N_20072,N_19927,N_19380);
nand U20073 (N_20073,N_19187,N_19416);
or U20074 (N_20074,N_19428,N_19065);
or U20075 (N_20075,N_19312,N_19531);
and U20076 (N_20076,N_19590,N_19399);
and U20077 (N_20077,N_19043,N_19714);
or U20078 (N_20078,N_19193,N_19842);
or U20079 (N_20079,N_19291,N_19204);
nor U20080 (N_20080,N_19934,N_19680);
or U20081 (N_20081,N_19015,N_19701);
nor U20082 (N_20082,N_19969,N_19717);
or U20083 (N_20083,N_19612,N_19095);
xor U20084 (N_20084,N_19572,N_19945);
or U20085 (N_20085,N_19079,N_19462);
xor U20086 (N_20086,N_19026,N_19090);
and U20087 (N_20087,N_19746,N_19898);
nor U20088 (N_20088,N_19286,N_19111);
and U20089 (N_20089,N_19815,N_19088);
and U20090 (N_20090,N_19489,N_19743);
or U20091 (N_20091,N_19519,N_19738);
and U20092 (N_20092,N_19574,N_19639);
and U20093 (N_20093,N_19569,N_19877);
and U20094 (N_20094,N_19682,N_19845);
xor U20095 (N_20095,N_19308,N_19555);
nor U20096 (N_20096,N_19259,N_19355);
and U20097 (N_20097,N_19897,N_19697);
nor U20098 (N_20098,N_19646,N_19907);
nand U20099 (N_20099,N_19406,N_19254);
nand U20100 (N_20100,N_19848,N_19534);
and U20101 (N_20101,N_19182,N_19290);
nand U20102 (N_20102,N_19441,N_19632);
or U20103 (N_20103,N_19236,N_19604);
nor U20104 (N_20104,N_19072,N_19756);
and U20105 (N_20105,N_19445,N_19008);
nor U20106 (N_20106,N_19151,N_19689);
and U20107 (N_20107,N_19958,N_19266);
and U20108 (N_20108,N_19484,N_19481);
or U20109 (N_20109,N_19262,N_19061);
or U20110 (N_20110,N_19402,N_19723);
and U20111 (N_20111,N_19243,N_19997);
and U20112 (N_20112,N_19673,N_19702);
and U20113 (N_20113,N_19272,N_19014);
or U20114 (N_20114,N_19025,N_19802);
and U20115 (N_20115,N_19944,N_19074);
nor U20116 (N_20116,N_19361,N_19664);
nor U20117 (N_20117,N_19488,N_19225);
nand U20118 (N_20118,N_19729,N_19506);
xnor U20119 (N_20119,N_19640,N_19206);
or U20120 (N_20120,N_19753,N_19885);
and U20121 (N_20121,N_19754,N_19018);
nor U20122 (N_20122,N_19974,N_19705);
and U20123 (N_20123,N_19625,N_19497);
or U20124 (N_20124,N_19707,N_19889);
xor U20125 (N_20125,N_19320,N_19887);
nand U20126 (N_20126,N_19890,N_19981);
or U20127 (N_20127,N_19033,N_19197);
nand U20128 (N_20128,N_19571,N_19238);
xor U20129 (N_20129,N_19933,N_19662);
nor U20130 (N_20130,N_19641,N_19669);
and U20131 (N_20131,N_19977,N_19681);
or U20132 (N_20132,N_19263,N_19017);
nand U20133 (N_20133,N_19102,N_19327);
nor U20134 (N_20134,N_19732,N_19854);
or U20135 (N_20135,N_19396,N_19718);
xor U20136 (N_20136,N_19089,N_19964);
xor U20137 (N_20137,N_19030,N_19623);
or U20138 (N_20138,N_19580,N_19633);
or U20139 (N_20139,N_19850,N_19215);
xnor U20140 (N_20140,N_19980,N_19093);
nor U20141 (N_20141,N_19801,N_19028);
nand U20142 (N_20142,N_19455,N_19359);
and U20143 (N_20143,N_19199,N_19888);
xnor U20144 (N_20144,N_19374,N_19896);
and U20145 (N_20145,N_19871,N_19443);
nand U20146 (N_20146,N_19721,N_19367);
or U20147 (N_20147,N_19282,N_19096);
nor U20148 (N_20148,N_19740,N_19292);
nand U20149 (N_20149,N_19141,N_19722);
xnor U20150 (N_20150,N_19894,N_19078);
xnor U20151 (N_20151,N_19267,N_19270);
or U20152 (N_20152,N_19698,N_19514);
and U20153 (N_20153,N_19786,N_19430);
or U20154 (N_20154,N_19996,N_19712);
nor U20155 (N_20155,N_19955,N_19553);
nor U20156 (N_20156,N_19289,N_19766);
nand U20157 (N_20157,N_19734,N_19203);
or U20158 (N_20158,N_19570,N_19427);
and U20159 (N_20159,N_19763,N_19004);
or U20160 (N_20160,N_19608,N_19276);
nor U20161 (N_20161,N_19132,N_19176);
nand U20162 (N_20162,N_19836,N_19548);
xor U20163 (N_20163,N_19774,N_19867);
or U20164 (N_20164,N_19139,N_19363);
or U20165 (N_20165,N_19654,N_19856);
nor U20166 (N_20166,N_19450,N_19034);
or U20167 (N_20167,N_19522,N_19954);
nand U20168 (N_20168,N_19685,N_19179);
nand U20169 (N_20169,N_19109,N_19777);
nor U20170 (N_20170,N_19067,N_19816);
nand U20171 (N_20171,N_19776,N_19160);
xor U20172 (N_20172,N_19157,N_19828);
or U20173 (N_20173,N_19318,N_19071);
and U20174 (N_20174,N_19227,N_19807);
and U20175 (N_20175,N_19260,N_19987);
xnor U20176 (N_20176,N_19235,N_19195);
nand U20177 (N_20177,N_19032,N_19645);
and U20178 (N_20178,N_19949,N_19822);
nand U20179 (N_20179,N_19216,N_19706);
xnor U20180 (N_20180,N_19843,N_19331);
nand U20181 (N_20181,N_19775,N_19338);
or U20182 (N_20182,N_19667,N_19048);
nor U20183 (N_20183,N_19366,N_19404);
or U20184 (N_20184,N_19460,N_19512);
xnor U20185 (N_20185,N_19762,N_19827);
or U20186 (N_20186,N_19222,N_19797);
nor U20187 (N_20187,N_19883,N_19556);
xnor U20188 (N_20188,N_19806,N_19953);
nor U20189 (N_20189,N_19838,N_19693);
nor U20190 (N_20190,N_19761,N_19869);
nor U20191 (N_20191,N_19509,N_19520);
xnor U20192 (N_20192,N_19476,N_19429);
xor U20193 (N_20193,N_19156,N_19704);
or U20194 (N_20194,N_19020,N_19676);
and U20195 (N_20195,N_19741,N_19821);
nor U20196 (N_20196,N_19314,N_19390);
xor U20197 (N_20197,N_19405,N_19630);
xnor U20198 (N_20198,N_19129,N_19961);
and U20199 (N_20199,N_19185,N_19456);
nor U20200 (N_20200,N_19609,N_19749);
and U20201 (N_20201,N_19679,N_19490);
nor U20202 (N_20202,N_19459,N_19013);
nand U20203 (N_20203,N_19552,N_19862);
nor U20204 (N_20204,N_19434,N_19528);
xor U20205 (N_20205,N_19105,N_19035);
nor U20206 (N_20206,N_19190,N_19508);
nand U20207 (N_20207,N_19870,N_19299);
nand U20208 (N_20208,N_19631,N_19736);
and U20209 (N_20209,N_19988,N_19334);
and U20210 (N_20210,N_19541,N_19943);
nor U20211 (N_20211,N_19148,N_19809);
nand U20212 (N_20212,N_19811,N_19167);
or U20213 (N_20213,N_19752,N_19052);
and U20214 (N_20214,N_19411,N_19819);
or U20215 (N_20215,N_19155,N_19172);
and U20216 (N_20216,N_19573,N_19650);
or U20217 (N_20217,N_19626,N_19125);
and U20218 (N_20218,N_19073,N_19576);
xor U20219 (N_20219,N_19965,N_19638);
and U20220 (N_20220,N_19847,N_19438);
nand U20221 (N_20221,N_19373,N_19083);
nor U20222 (N_20222,N_19543,N_19000);
or U20223 (N_20223,N_19200,N_19607);
or U20224 (N_20224,N_19239,N_19782);
nor U20225 (N_20225,N_19285,N_19739);
nand U20226 (N_20226,N_19087,N_19387);
or U20227 (N_20227,N_19670,N_19473);
and U20228 (N_20228,N_19959,N_19579);
nand U20229 (N_20229,N_19091,N_19039);
or U20230 (N_20230,N_19466,N_19419);
nor U20231 (N_20231,N_19144,N_19901);
nand U20232 (N_20232,N_19873,N_19233);
or U20233 (N_20233,N_19525,N_19180);
nor U20234 (N_20234,N_19582,N_19711);
nor U20235 (N_20235,N_19174,N_19866);
or U20236 (N_20236,N_19780,N_19687);
nand U20237 (N_20237,N_19315,N_19076);
xor U20238 (N_20238,N_19306,N_19523);
nand U20239 (N_20239,N_19325,N_19283);
nor U20240 (N_20240,N_19596,N_19728);
xor U20241 (N_20241,N_19765,N_19513);
or U20242 (N_20242,N_19166,N_19137);
nor U20243 (N_20243,N_19731,N_19602);
or U20244 (N_20244,N_19909,N_19535);
nor U20245 (N_20245,N_19656,N_19904);
nand U20246 (N_20246,N_19342,N_19330);
or U20247 (N_20247,N_19859,N_19124);
xor U20248 (N_20248,N_19659,N_19477);
nand U20249 (N_20249,N_19863,N_19277);
and U20250 (N_20250,N_19500,N_19536);
xnor U20251 (N_20251,N_19407,N_19163);
or U20252 (N_20252,N_19647,N_19966);
and U20253 (N_20253,N_19540,N_19063);
and U20254 (N_20254,N_19692,N_19627);
nor U20255 (N_20255,N_19830,N_19397);
xnor U20256 (N_20256,N_19603,N_19501);
xor U20257 (N_20257,N_19365,N_19767);
xor U20258 (N_20258,N_19624,N_19360);
nand U20259 (N_20259,N_19250,N_19049);
or U20260 (N_20260,N_19364,N_19437);
or U20261 (N_20261,N_19865,N_19324);
or U20262 (N_20262,N_19099,N_19972);
xnor U20263 (N_20263,N_19588,N_19170);
and U20264 (N_20264,N_19439,N_19134);
nand U20265 (N_20265,N_19558,N_19983);
nand U20266 (N_20266,N_19637,N_19143);
xnor U20267 (N_20267,N_19695,N_19852);
nor U20268 (N_20268,N_19831,N_19518);
nor U20269 (N_20269,N_19715,N_19293);
nand U20270 (N_20270,N_19655,N_19796);
xor U20271 (N_20271,N_19005,N_19678);
nor U20272 (N_20272,N_19348,N_19884);
nand U20273 (N_20273,N_19920,N_19086);
and U20274 (N_20274,N_19247,N_19386);
and U20275 (N_20275,N_19142,N_19823);
xor U20276 (N_20276,N_19202,N_19045);
nor U20277 (N_20277,N_19181,N_19748);
and U20278 (N_20278,N_19581,N_19635);
xnor U20279 (N_20279,N_19878,N_19726);
nor U20280 (N_20280,N_19788,N_19410);
nand U20281 (N_20281,N_19264,N_19357);
nand U20282 (N_20282,N_19321,N_19773);
nand U20283 (N_20283,N_19224,N_19597);
and U20284 (N_20284,N_19812,N_19092);
xnor U20285 (N_20285,N_19064,N_19173);
nor U20286 (N_20286,N_19496,N_19464);
and U20287 (N_20287,N_19384,N_19708);
or U20288 (N_20288,N_19658,N_19278);
nand U20289 (N_20289,N_19691,N_19421);
nand U20290 (N_20290,N_19529,N_19527);
or U20291 (N_20291,N_19993,N_19700);
and U20292 (N_20292,N_19652,N_19803);
or U20293 (N_20293,N_19677,N_19425);
nor U20294 (N_20294,N_19212,N_19230);
xor U20295 (N_20295,N_19516,N_19177);
and U20296 (N_20296,N_19493,N_19486);
xnor U20297 (N_20297,N_19661,N_19002);
xnor U20298 (N_20298,N_19454,N_19629);
xor U20299 (N_20299,N_19234,N_19417);
nor U20300 (N_20300,N_19799,N_19947);
xnor U20301 (N_20301,N_19671,N_19913);
nor U20302 (N_20302,N_19381,N_19912);
xor U20303 (N_20303,N_19694,N_19846);
nor U20304 (N_20304,N_19495,N_19304);
or U20305 (N_20305,N_19169,N_19333);
xor U20306 (N_20306,N_19779,N_19295);
and U20307 (N_20307,N_19899,N_19851);
or U20308 (N_20308,N_19379,N_19551);
nand U20309 (N_20309,N_19683,N_19245);
and U20310 (N_20310,N_19924,N_19081);
nand U20311 (N_20311,N_19059,N_19499);
and U20312 (N_20312,N_19413,N_19352);
nand U20313 (N_20313,N_19902,N_19418);
and U20314 (N_20314,N_19544,N_19307);
nand U20315 (N_20315,N_19592,N_19377);
or U20316 (N_20316,N_19253,N_19001);
nor U20317 (N_20317,N_19103,N_19244);
xor U20318 (N_20318,N_19246,N_19601);
and U20319 (N_20319,N_19644,N_19146);
and U20320 (N_20320,N_19937,N_19908);
nand U20321 (N_20321,N_19892,N_19175);
nor U20322 (N_20322,N_19643,N_19875);
or U20323 (N_20323,N_19356,N_19936);
nor U20324 (N_20324,N_19284,N_19724);
or U20325 (N_20325,N_19686,N_19240);
and U20326 (N_20326,N_19941,N_19184);
or U20327 (N_20327,N_19408,N_19946);
nor U20328 (N_20328,N_19024,N_19636);
and U20329 (N_20329,N_19300,N_19168);
and U20330 (N_20330,N_19249,N_19857);
nand U20331 (N_20331,N_19189,N_19341);
xor U20332 (N_20332,N_19696,N_19467);
nand U20333 (N_20333,N_19975,N_19346);
or U20334 (N_20334,N_19389,N_19921);
or U20335 (N_20335,N_19273,N_19808);
nand U20336 (N_20336,N_19804,N_19201);
or U20337 (N_20337,N_19978,N_19790);
nand U20338 (N_20338,N_19021,N_19872);
or U20339 (N_20339,N_19457,N_19825);
nor U20340 (N_20340,N_19463,N_19511);
xnor U20341 (N_20341,N_19060,N_19550);
xnor U20342 (N_20342,N_19223,N_19577);
and U20343 (N_20343,N_19532,N_19960);
xnor U20344 (N_20344,N_19053,N_19818);
and U20345 (N_20345,N_19424,N_19147);
and U20346 (N_20346,N_19023,N_19521);
xnor U20347 (N_20347,N_19565,N_19232);
or U20348 (N_20348,N_19153,N_19620);
and U20349 (N_20349,N_19326,N_19595);
nor U20350 (N_20350,N_19084,N_19547);
or U20351 (N_20351,N_19733,N_19145);
and U20352 (N_20352,N_19412,N_19340);
and U20353 (N_20353,N_19713,N_19296);
xnor U20354 (N_20354,N_19614,N_19989);
nand U20355 (N_20355,N_19178,N_19047);
or U20356 (N_20356,N_19198,N_19041);
or U20357 (N_20357,N_19011,N_19688);
nor U20358 (N_20358,N_19337,N_19110);
and U20359 (N_20359,N_19475,N_19874);
nor U20360 (N_20360,N_19165,N_19929);
xor U20361 (N_20361,N_19133,N_19375);
and U20362 (N_20362,N_19478,N_19107);
xnor U20363 (N_20363,N_19760,N_19393);
nand U20364 (N_20364,N_19158,N_19470);
xor U20365 (N_20365,N_19668,N_19787);
and U20366 (N_20366,N_19526,N_19171);
and U20367 (N_20367,N_19893,N_19951);
or U20368 (N_20368,N_19016,N_19226);
xor U20369 (N_20369,N_19970,N_19274);
xnor U20370 (N_20370,N_19112,N_19745);
xnor U20371 (N_20371,N_19069,N_19616);
or U20372 (N_20372,N_19855,N_19591);
xnor U20373 (N_20373,N_19159,N_19622);
and U20374 (N_20374,N_19383,N_19840);
or U20375 (N_20375,N_19976,N_19162);
nand U20376 (N_20376,N_19999,N_19824);
or U20377 (N_20377,N_19448,N_19881);
or U20378 (N_20378,N_19265,N_19789);
nor U20379 (N_20379,N_19895,N_19126);
nand U20380 (N_20380,N_19022,N_19926);
and U20381 (N_20381,N_19759,N_19012);
nor U20382 (N_20382,N_19122,N_19557);
or U20383 (N_20383,N_19268,N_19279);
nand U20384 (N_20384,N_19810,N_19336);
or U20385 (N_20385,N_19492,N_19219);
xor U20386 (N_20386,N_19530,N_19751);
nand U20387 (N_20387,N_19350,N_19628);
nand U20388 (N_20388,N_19335,N_19319);
or U20389 (N_20389,N_19347,N_19196);
nand U20390 (N_20390,N_19930,N_19716);
and U20391 (N_20391,N_19963,N_19709);
nand U20392 (N_20392,N_19056,N_19510);
xnor U20393 (N_20393,N_19593,N_19007);
nor U20394 (N_20394,N_19343,N_19925);
or U20395 (N_20395,N_19271,N_19793);
xnor U20396 (N_20396,N_19992,N_19517);
and U20397 (N_20397,N_19164,N_19298);
nand U20398 (N_20398,N_19309,N_19422);
nand U20399 (N_20399,N_19036,N_19207);
nand U20400 (N_20400,N_19152,N_19882);
and U20401 (N_20401,N_19040,N_19699);
nor U20402 (N_20402,N_19392,N_19615);
nand U20403 (N_20403,N_19719,N_19003);
nand U20404 (N_20404,N_19113,N_19275);
nand U20405 (N_20405,N_19914,N_19322);
and U20406 (N_20406,N_19915,N_19482);
and U20407 (N_20407,N_19301,N_19297);
nor U20408 (N_20408,N_19231,N_19800);
or U20409 (N_20409,N_19939,N_19648);
xor U20410 (N_20410,N_19684,N_19771);
nor U20411 (N_20411,N_19533,N_19653);
nor U20412 (N_20412,N_19982,N_19237);
or U20413 (N_20413,N_19354,N_19876);
or U20414 (N_20414,N_19503,N_19186);
nor U20415 (N_20415,N_19019,N_19332);
nand U20416 (N_20416,N_19725,N_19205);
nor U20417 (N_20417,N_19764,N_19128);
and U20418 (N_20418,N_19192,N_19051);
xor U20419 (N_20419,N_19077,N_19031);
nand U20420 (N_20420,N_19940,N_19832);
nand U20421 (N_20421,N_19287,N_19372);
nand U20422 (N_20422,N_19453,N_19317);
or U20423 (N_20423,N_19491,N_19351);
or U20424 (N_20424,N_19323,N_19485);
nor U20425 (N_20425,N_19879,N_19362);
nor U20426 (N_20426,N_19242,N_19922);
xnor U20427 (N_20427,N_19559,N_19316);
or U20428 (N_20428,N_19269,N_19009);
or U20429 (N_20429,N_19598,N_19605);
nand U20430 (N_20430,N_19672,N_19038);
or U20431 (N_20431,N_19329,N_19255);
nor U20432 (N_20432,N_19549,N_19906);
nand U20433 (N_20433,N_19055,N_19957);
or U20434 (N_20434,N_19853,N_19130);
nor U20435 (N_20435,N_19123,N_19735);
xor U20436 (N_20436,N_19229,N_19613);
and U20437 (N_20437,N_19191,N_19037);
xnor U20438 (N_20438,N_19119,N_19114);
xnor U20439 (N_20439,N_19568,N_19461);
nand U20440 (N_20440,N_19442,N_19594);
and U20441 (N_20441,N_19085,N_19814);
or U20442 (N_20442,N_19465,N_19916);
or U20443 (N_20443,N_19575,N_19546);
or U20444 (N_20444,N_19288,N_19220);
xor U20445 (N_20445,N_19339,N_19829);
or U20446 (N_20446,N_19617,N_19903);
nand U20447 (N_20447,N_19294,N_19860);
xor U20448 (N_20448,N_19795,N_19066);
or U20449 (N_20449,N_19368,N_19423);
nor U20450 (N_20450,N_19833,N_19649);
and U20451 (N_20451,N_19057,N_19868);
and U20452 (N_20452,N_19861,N_19663);
nor U20453 (N_20453,N_19962,N_19161);
and U20454 (N_20454,N_19835,N_19106);
and U20455 (N_20455,N_19798,N_19118);
nand U20456 (N_20456,N_19690,N_19805);
xor U20457 (N_20457,N_19979,N_19991);
and U20458 (N_20458,N_19994,N_19950);
nand U20459 (N_20459,N_19029,N_19651);
and U20460 (N_20460,N_19449,N_19606);
nand U20461 (N_20461,N_19415,N_19257);
and U20462 (N_20462,N_19131,N_19154);
or U20463 (N_20463,N_19070,N_19435);
nor U20464 (N_20464,N_19834,N_19344);
nand U20465 (N_20465,N_19218,N_19256);
and U20466 (N_20466,N_19062,N_19345);
nor U20467 (N_20467,N_19382,N_19369);
nor U20468 (N_20468,N_19398,N_19634);
nor U20469 (N_20469,N_19858,N_19956);
or U20470 (N_20470,N_19313,N_19727);
and U20471 (N_20471,N_19214,N_19504);
xnor U20472 (N_20472,N_19140,N_19563);
nand U20473 (N_20473,N_19599,N_19781);
and U20474 (N_20474,N_19104,N_19968);
or U20475 (N_20475,N_19395,N_19703);
or U20476 (N_20476,N_19054,N_19757);
xor U20477 (N_20477,N_19864,N_19469);
nor U20478 (N_20478,N_19100,N_19600);
and U20479 (N_20479,N_19998,N_19251);
nor U20480 (N_20480,N_19538,N_19358);
and U20481 (N_20481,N_19116,N_19046);
or U20482 (N_20482,N_19545,N_19931);
nor U20483 (N_20483,N_19537,N_19006);
and U20484 (N_20484,N_19082,N_19618);
or U20485 (N_20485,N_19494,N_19783);
and U20486 (N_20486,N_19948,N_19917);
nor U20487 (N_20487,N_19483,N_19149);
or U20488 (N_20488,N_19610,N_19935);
xnor U20489 (N_20489,N_19208,N_19905);
xor U20490 (N_20490,N_19097,N_19101);
xnor U20491 (N_20491,N_19770,N_19772);
xnor U20492 (N_20492,N_19891,N_19505);
nand U20493 (N_20493,N_19328,N_19938);
or U20494 (N_20494,N_19138,N_19730);
or U20495 (N_20495,N_19431,N_19471);
nand U20496 (N_20496,N_19120,N_19209);
nor U20497 (N_20497,N_19813,N_19451);
or U20498 (N_20498,N_19578,N_19742);
nor U20499 (N_20499,N_19900,N_19487);
or U20500 (N_20500,N_19543,N_19106);
nand U20501 (N_20501,N_19777,N_19103);
nor U20502 (N_20502,N_19190,N_19236);
nand U20503 (N_20503,N_19912,N_19110);
nor U20504 (N_20504,N_19603,N_19956);
or U20505 (N_20505,N_19533,N_19568);
or U20506 (N_20506,N_19646,N_19397);
nand U20507 (N_20507,N_19481,N_19210);
xor U20508 (N_20508,N_19990,N_19554);
nand U20509 (N_20509,N_19848,N_19868);
nand U20510 (N_20510,N_19712,N_19501);
or U20511 (N_20511,N_19695,N_19438);
nand U20512 (N_20512,N_19834,N_19779);
nand U20513 (N_20513,N_19661,N_19807);
nor U20514 (N_20514,N_19063,N_19663);
or U20515 (N_20515,N_19263,N_19933);
nor U20516 (N_20516,N_19448,N_19830);
nor U20517 (N_20517,N_19923,N_19860);
nor U20518 (N_20518,N_19550,N_19519);
and U20519 (N_20519,N_19585,N_19797);
xor U20520 (N_20520,N_19497,N_19492);
xnor U20521 (N_20521,N_19852,N_19210);
or U20522 (N_20522,N_19752,N_19994);
and U20523 (N_20523,N_19580,N_19448);
and U20524 (N_20524,N_19779,N_19959);
or U20525 (N_20525,N_19167,N_19726);
nor U20526 (N_20526,N_19611,N_19162);
and U20527 (N_20527,N_19304,N_19233);
nand U20528 (N_20528,N_19924,N_19125);
and U20529 (N_20529,N_19097,N_19995);
or U20530 (N_20530,N_19391,N_19180);
or U20531 (N_20531,N_19275,N_19967);
or U20532 (N_20532,N_19653,N_19987);
nand U20533 (N_20533,N_19095,N_19705);
xnor U20534 (N_20534,N_19374,N_19310);
nand U20535 (N_20535,N_19876,N_19707);
nor U20536 (N_20536,N_19074,N_19616);
or U20537 (N_20537,N_19225,N_19828);
nor U20538 (N_20538,N_19258,N_19163);
or U20539 (N_20539,N_19889,N_19178);
nor U20540 (N_20540,N_19512,N_19935);
or U20541 (N_20541,N_19876,N_19975);
nor U20542 (N_20542,N_19260,N_19644);
xnor U20543 (N_20543,N_19081,N_19545);
nand U20544 (N_20544,N_19249,N_19648);
nand U20545 (N_20545,N_19985,N_19083);
or U20546 (N_20546,N_19810,N_19856);
xnor U20547 (N_20547,N_19822,N_19843);
nand U20548 (N_20548,N_19044,N_19993);
nand U20549 (N_20549,N_19343,N_19142);
or U20550 (N_20550,N_19728,N_19607);
and U20551 (N_20551,N_19119,N_19201);
and U20552 (N_20552,N_19842,N_19138);
nand U20553 (N_20553,N_19919,N_19294);
and U20554 (N_20554,N_19719,N_19824);
nand U20555 (N_20555,N_19856,N_19737);
or U20556 (N_20556,N_19113,N_19184);
xor U20557 (N_20557,N_19730,N_19654);
or U20558 (N_20558,N_19606,N_19387);
or U20559 (N_20559,N_19316,N_19639);
and U20560 (N_20560,N_19199,N_19669);
xor U20561 (N_20561,N_19156,N_19504);
nand U20562 (N_20562,N_19425,N_19376);
nand U20563 (N_20563,N_19625,N_19225);
nor U20564 (N_20564,N_19512,N_19926);
xor U20565 (N_20565,N_19719,N_19407);
nor U20566 (N_20566,N_19249,N_19437);
and U20567 (N_20567,N_19495,N_19039);
and U20568 (N_20568,N_19430,N_19911);
and U20569 (N_20569,N_19098,N_19449);
or U20570 (N_20570,N_19969,N_19191);
xor U20571 (N_20571,N_19492,N_19298);
nand U20572 (N_20572,N_19780,N_19312);
nand U20573 (N_20573,N_19096,N_19830);
xor U20574 (N_20574,N_19639,N_19543);
nor U20575 (N_20575,N_19517,N_19186);
nand U20576 (N_20576,N_19869,N_19712);
nor U20577 (N_20577,N_19106,N_19602);
nor U20578 (N_20578,N_19394,N_19986);
nor U20579 (N_20579,N_19766,N_19568);
xnor U20580 (N_20580,N_19324,N_19352);
nand U20581 (N_20581,N_19683,N_19933);
nor U20582 (N_20582,N_19010,N_19524);
xnor U20583 (N_20583,N_19504,N_19998);
and U20584 (N_20584,N_19958,N_19635);
nand U20585 (N_20585,N_19236,N_19325);
xnor U20586 (N_20586,N_19978,N_19720);
nor U20587 (N_20587,N_19936,N_19933);
xnor U20588 (N_20588,N_19226,N_19521);
nand U20589 (N_20589,N_19029,N_19519);
nand U20590 (N_20590,N_19373,N_19473);
nor U20591 (N_20591,N_19200,N_19799);
or U20592 (N_20592,N_19654,N_19846);
nor U20593 (N_20593,N_19969,N_19744);
and U20594 (N_20594,N_19503,N_19435);
xor U20595 (N_20595,N_19758,N_19421);
or U20596 (N_20596,N_19437,N_19218);
xnor U20597 (N_20597,N_19974,N_19201);
and U20598 (N_20598,N_19290,N_19163);
or U20599 (N_20599,N_19075,N_19200);
and U20600 (N_20600,N_19853,N_19565);
and U20601 (N_20601,N_19308,N_19062);
or U20602 (N_20602,N_19363,N_19849);
nand U20603 (N_20603,N_19171,N_19808);
nor U20604 (N_20604,N_19017,N_19014);
xnor U20605 (N_20605,N_19398,N_19174);
nor U20606 (N_20606,N_19686,N_19576);
xnor U20607 (N_20607,N_19419,N_19839);
or U20608 (N_20608,N_19082,N_19339);
nor U20609 (N_20609,N_19291,N_19333);
nor U20610 (N_20610,N_19712,N_19175);
or U20611 (N_20611,N_19759,N_19446);
xor U20612 (N_20612,N_19367,N_19511);
nor U20613 (N_20613,N_19728,N_19857);
or U20614 (N_20614,N_19023,N_19965);
nor U20615 (N_20615,N_19408,N_19593);
xnor U20616 (N_20616,N_19025,N_19847);
xnor U20617 (N_20617,N_19219,N_19230);
nor U20618 (N_20618,N_19863,N_19979);
nand U20619 (N_20619,N_19069,N_19383);
or U20620 (N_20620,N_19540,N_19830);
xor U20621 (N_20621,N_19338,N_19779);
or U20622 (N_20622,N_19524,N_19843);
and U20623 (N_20623,N_19247,N_19394);
and U20624 (N_20624,N_19491,N_19367);
nor U20625 (N_20625,N_19022,N_19251);
nand U20626 (N_20626,N_19544,N_19717);
and U20627 (N_20627,N_19519,N_19894);
nand U20628 (N_20628,N_19492,N_19290);
or U20629 (N_20629,N_19022,N_19782);
nor U20630 (N_20630,N_19684,N_19030);
or U20631 (N_20631,N_19877,N_19995);
xor U20632 (N_20632,N_19766,N_19060);
and U20633 (N_20633,N_19714,N_19287);
or U20634 (N_20634,N_19904,N_19890);
nand U20635 (N_20635,N_19950,N_19055);
nand U20636 (N_20636,N_19366,N_19544);
or U20637 (N_20637,N_19388,N_19080);
nand U20638 (N_20638,N_19063,N_19505);
and U20639 (N_20639,N_19133,N_19916);
or U20640 (N_20640,N_19998,N_19709);
nand U20641 (N_20641,N_19514,N_19441);
nor U20642 (N_20642,N_19438,N_19340);
nand U20643 (N_20643,N_19547,N_19826);
or U20644 (N_20644,N_19617,N_19017);
or U20645 (N_20645,N_19854,N_19717);
nor U20646 (N_20646,N_19311,N_19516);
and U20647 (N_20647,N_19862,N_19428);
nor U20648 (N_20648,N_19001,N_19414);
xor U20649 (N_20649,N_19608,N_19461);
nand U20650 (N_20650,N_19793,N_19325);
or U20651 (N_20651,N_19113,N_19242);
or U20652 (N_20652,N_19716,N_19587);
nor U20653 (N_20653,N_19034,N_19700);
xnor U20654 (N_20654,N_19446,N_19903);
xnor U20655 (N_20655,N_19261,N_19211);
nor U20656 (N_20656,N_19776,N_19669);
nand U20657 (N_20657,N_19409,N_19548);
nor U20658 (N_20658,N_19016,N_19162);
and U20659 (N_20659,N_19402,N_19571);
and U20660 (N_20660,N_19594,N_19749);
xnor U20661 (N_20661,N_19678,N_19928);
nand U20662 (N_20662,N_19039,N_19832);
or U20663 (N_20663,N_19136,N_19779);
nor U20664 (N_20664,N_19464,N_19772);
or U20665 (N_20665,N_19984,N_19721);
nand U20666 (N_20666,N_19012,N_19965);
nor U20667 (N_20667,N_19265,N_19417);
and U20668 (N_20668,N_19270,N_19318);
or U20669 (N_20669,N_19760,N_19019);
xor U20670 (N_20670,N_19463,N_19371);
or U20671 (N_20671,N_19196,N_19327);
nand U20672 (N_20672,N_19031,N_19668);
nor U20673 (N_20673,N_19290,N_19516);
nor U20674 (N_20674,N_19314,N_19490);
or U20675 (N_20675,N_19663,N_19355);
xor U20676 (N_20676,N_19565,N_19407);
nand U20677 (N_20677,N_19100,N_19730);
nand U20678 (N_20678,N_19781,N_19856);
xor U20679 (N_20679,N_19289,N_19911);
xnor U20680 (N_20680,N_19228,N_19151);
and U20681 (N_20681,N_19458,N_19910);
and U20682 (N_20682,N_19280,N_19167);
or U20683 (N_20683,N_19344,N_19385);
xnor U20684 (N_20684,N_19264,N_19997);
and U20685 (N_20685,N_19359,N_19130);
or U20686 (N_20686,N_19827,N_19021);
or U20687 (N_20687,N_19982,N_19530);
xor U20688 (N_20688,N_19444,N_19723);
xor U20689 (N_20689,N_19159,N_19811);
xnor U20690 (N_20690,N_19559,N_19233);
nand U20691 (N_20691,N_19778,N_19581);
xnor U20692 (N_20692,N_19481,N_19446);
nand U20693 (N_20693,N_19543,N_19349);
nand U20694 (N_20694,N_19728,N_19964);
xor U20695 (N_20695,N_19037,N_19507);
xor U20696 (N_20696,N_19715,N_19129);
or U20697 (N_20697,N_19742,N_19790);
and U20698 (N_20698,N_19400,N_19781);
nor U20699 (N_20699,N_19797,N_19102);
and U20700 (N_20700,N_19867,N_19788);
nor U20701 (N_20701,N_19860,N_19410);
and U20702 (N_20702,N_19748,N_19872);
and U20703 (N_20703,N_19724,N_19091);
and U20704 (N_20704,N_19707,N_19073);
and U20705 (N_20705,N_19561,N_19742);
xnor U20706 (N_20706,N_19233,N_19793);
and U20707 (N_20707,N_19585,N_19234);
xnor U20708 (N_20708,N_19821,N_19396);
and U20709 (N_20709,N_19841,N_19113);
or U20710 (N_20710,N_19982,N_19798);
nor U20711 (N_20711,N_19830,N_19592);
or U20712 (N_20712,N_19371,N_19041);
or U20713 (N_20713,N_19751,N_19237);
nand U20714 (N_20714,N_19890,N_19919);
nand U20715 (N_20715,N_19688,N_19997);
xor U20716 (N_20716,N_19076,N_19765);
xor U20717 (N_20717,N_19891,N_19376);
xnor U20718 (N_20718,N_19488,N_19475);
xnor U20719 (N_20719,N_19310,N_19506);
and U20720 (N_20720,N_19167,N_19666);
xor U20721 (N_20721,N_19731,N_19557);
or U20722 (N_20722,N_19282,N_19750);
nand U20723 (N_20723,N_19695,N_19175);
nand U20724 (N_20724,N_19519,N_19491);
xnor U20725 (N_20725,N_19536,N_19540);
xor U20726 (N_20726,N_19217,N_19048);
and U20727 (N_20727,N_19086,N_19163);
nor U20728 (N_20728,N_19541,N_19029);
nand U20729 (N_20729,N_19303,N_19599);
nor U20730 (N_20730,N_19441,N_19123);
or U20731 (N_20731,N_19050,N_19098);
and U20732 (N_20732,N_19386,N_19293);
xor U20733 (N_20733,N_19121,N_19592);
xnor U20734 (N_20734,N_19101,N_19851);
nand U20735 (N_20735,N_19508,N_19578);
xor U20736 (N_20736,N_19653,N_19888);
nand U20737 (N_20737,N_19080,N_19667);
or U20738 (N_20738,N_19477,N_19893);
and U20739 (N_20739,N_19284,N_19048);
and U20740 (N_20740,N_19976,N_19430);
and U20741 (N_20741,N_19091,N_19404);
nand U20742 (N_20742,N_19998,N_19915);
nor U20743 (N_20743,N_19844,N_19803);
and U20744 (N_20744,N_19569,N_19374);
nor U20745 (N_20745,N_19799,N_19824);
nand U20746 (N_20746,N_19370,N_19074);
nand U20747 (N_20747,N_19771,N_19515);
or U20748 (N_20748,N_19128,N_19186);
xnor U20749 (N_20749,N_19151,N_19608);
or U20750 (N_20750,N_19955,N_19601);
nand U20751 (N_20751,N_19815,N_19149);
xor U20752 (N_20752,N_19604,N_19788);
nor U20753 (N_20753,N_19466,N_19217);
nor U20754 (N_20754,N_19597,N_19027);
nand U20755 (N_20755,N_19762,N_19749);
xor U20756 (N_20756,N_19060,N_19992);
or U20757 (N_20757,N_19384,N_19924);
xnor U20758 (N_20758,N_19627,N_19972);
or U20759 (N_20759,N_19444,N_19305);
nor U20760 (N_20760,N_19894,N_19946);
and U20761 (N_20761,N_19995,N_19665);
or U20762 (N_20762,N_19264,N_19648);
or U20763 (N_20763,N_19255,N_19775);
nand U20764 (N_20764,N_19392,N_19304);
nand U20765 (N_20765,N_19217,N_19497);
nand U20766 (N_20766,N_19425,N_19195);
nand U20767 (N_20767,N_19472,N_19699);
xor U20768 (N_20768,N_19597,N_19207);
and U20769 (N_20769,N_19575,N_19820);
or U20770 (N_20770,N_19189,N_19560);
nor U20771 (N_20771,N_19319,N_19188);
nand U20772 (N_20772,N_19430,N_19064);
xnor U20773 (N_20773,N_19770,N_19803);
nor U20774 (N_20774,N_19234,N_19568);
xnor U20775 (N_20775,N_19672,N_19140);
nand U20776 (N_20776,N_19951,N_19949);
xor U20777 (N_20777,N_19437,N_19828);
nor U20778 (N_20778,N_19365,N_19594);
or U20779 (N_20779,N_19077,N_19279);
nor U20780 (N_20780,N_19920,N_19237);
and U20781 (N_20781,N_19499,N_19583);
and U20782 (N_20782,N_19802,N_19339);
nor U20783 (N_20783,N_19846,N_19516);
nand U20784 (N_20784,N_19302,N_19787);
and U20785 (N_20785,N_19000,N_19497);
xor U20786 (N_20786,N_19265,N_19012);
or U20787 (N_20787,N_19745,N_19553);
or U20788 (N_20788,N_19317,N_19842);
or U20789 (N_20789,N_19779,N_19322);
xnor U20790 (N_20790,N_19896,N_19661);
nor U20791 (N_20791,N_19563,N_19951);
nor U20792 (N_20792,N_19410,N_19082);
nor U20793 (N_20793,N_19299,N_19218);
xnor U20794 (N_20794,N_19122,N_19034);
or U20795 (N_20795,N_19421,N_19035);
or U20796 (N_20796,N_19284,N_19938);
nor U20797 (N_20797,N_19747,N_19444);
nand U20798 (N_20798,N_19222,N_19291);
nor U20799 (N_20799,N_19056,N_19066);
or U20800 (N_20800,N_19949,N_19049);
nor U20801 (N_20801,N_19600,N_19295);
xor U20802 (N_20802,N_19389,N_19616);
nor U20803 (N_20803,N_19609,N_19660);
xnor U20804 (N_20804,N_19038,N_19647);
nand U20805 (N_20805,N_19807,N_19415);
nand U20806 (N_20806,N_19593,N_19263);
nor U20807 (N_20807,N_19806,N_19031);
nor U20808 (N_20808,N_19688,N_19260);
nor U20809 (N_20809,N_19454,N_19932);
nor U20810 (N_20810,N_19117,N_19027);
and U20811 (N_20811,N_19943,N_19004);
nand U20812 (N_20812,N_19788,N_19752);
or U20813 (N_20813,N_19079,N_19622);
xor U20814 (N_20814,N_19596,N_19164);
xnor U20815 (N_20815,N_19089,N_19936);
and U20816 (N_20816,N_19545,N_19226);
and U20817 (N_20817,N_19240,N_19849);
or U20818 (N_20818,N_19446,N_19823);
and U20819 (N_20819,N_19534,N_19834);
nand U20820 (N_20820,N_19791,N_19806);
nand U20821 (N_20821,N_19031,N_19012);
or U20822 (N_20822,N_19977,N_19335);
nor U20823 (N_20823,N_19858,N_19372);
nand U20824 (N_20824,N_19833,N_19320);
or U20825 (N_20825,N_19952,N_19464);
and U20826 (N_20826,N_19183,N_19336);
nor U20827 (N_20827,N_19386,N_19588);
and U20828 (N_20828,N_19662,N_19820);
nor U20829 (N_20829,N_19573,N_19481);
xor U20830 (N_20830,N_19870,N_19187);
nor U20831 (N_20831,N_19474,N_19154);
or U20832 (N_20832,N_19546,N_19865);
xor U20833 (N_20833,N_19032,N_19168);
xnor U20834 (N_20834,N_19935,N_19548);
nor U20835 (N_20835,N_19218,N_19386);
and U20836 (N_20836,N_19552,N_19535);
nand U20837 (N_20837,N_19248,N_19427);
and U20838 (N_20838,N_19148,N_19108);
xnor U20839 (N_20839,N_19413,N_19268);
or U20840 (N_20840,N_19678,N_19827);
xor U20841 (N_20841,N_19228,N_19659);
xnor U20842 (N_20842,N_19811,N_19737);
nor U20843 (N_20843,N_19567,N_19657);
nor U20844 (N_20844,N_19499,N_19846);
nor U20845 (N_20845,N_19012,N_19584);
and U20846 (N_20846,N_19334,N_19980);
xor U20847 (N_20847,N_19098,N_19233);
nand U20848 (N_20848,N_19987,N_19852);
nor U20849 (N_20849,N_19491,N_19295);
xor U20850 (N_20850,N_19610,N_19286);
and U20851 (N_20851,N_19439,N_19456);
nand U20852 (N_20852,N_19397,N_19105);
and U20853 (N_20853,N_19907,N_19957);
xnor U20854 (N_20854,N_19457,N_19117);
or U20855 (N_20855,N_19364,N_19687);
or U20856 (N_20856,N_19879,N_19889);
and U20857 (N_20857,N_19214,N_19397);
or U20858 (N_20858,N_19346,N_19183);
xnor U20859 (N_20859,N_19654,N_19457);
nand U20860 (N_20860,N_19601,N_19293);
xnor U20861 (N_20861,N_19635,N_19038);
and U20862 (N_20862,N_19267,N_19766);
xor U20863 (N_20863,N_19808,N_19125);
nor U20864 (N_20864,N_19945,N_19148);
nor U20865 (N_20865,N_19096,N_19112);
nor U20866 (N_20866,N_19606,N_19907);
and U20867 (N_20867,N_19905,N_19079);
nor U20868 (N_20868,N_19131,N_19034);
or U20869 (N_20869,N_19646,N_19772);
nor U20870 (N_20870,N_19434,N_19180);
nor U20871 (N_20871,N_19466,N_19117);
xnor U20872 (N_20872,N_19203,N_19497);
nor U20873 (N_20873,N_19611,N_19172);
nand U20874 (N_20874,N_19439,N_19856);
nand U20875 (N_20875,N_19476,N_19194);
and U20876 (N_20876,N_19252,N_19057);
and U20877 (N_20877,N_19537,N_19496);
and U20878 (N_20878,N_19109,N_19089);
and U20879 (N_20879,N_19714,N_19491);
or U20880 (N_20880,N_19556,N_19630);
and U20881 (N_20881,N_19024,N_19377);
nor U20882 (N_20882,N_19619,N_19086);
nand U20883 (N_20883,N_19550,N_19278);
nand U20884 (N_20884,N_19839,N_19084);
xor U20885 (N_20885,N_19775,N_19066);
xnor U20886 (N_20886,N_19273,N_19643);
xnor U20887 (N_20887,N_19688,N_19374);
xor U20888 (N_20888,N_19118,N_19747);
or U20889 (N_20889,N_19202,N_19125);
xor U20890 (N_20890,N_19805,N_19174);
and U20891 (N_20891,N_19772,N_19775);
or U20892 (N_20892,N_19731,N_19492);
xor U20893 (N_20893,N_19464,N_19906);
xor U20894 (N_20894,N_19178,N_19154);
nand U20895 (N_20895,N_19422,N_19121);
and U20896 (N_20896,N_19728,N_19552);
and U20897 (N_20897,N_19754,N_19961);
and U20898 (N_20898,N_19986,N_19987);
nor U20899 (N_20899,N_19483,N_19415);
and U20900 (N_20900,N_19585,N_19272);
nand U20901 (N_20901,N_19624,N_19548);
and U20902 (N_20902,N_19430,N_19572);
nor U20903 (N_20903,N_19026,N_19489);
and U20904 (N_20904,N_19030,N_19927);
and U20905 (N_20905,N_19819,N_19130);
or U20906 (N_20906,N_19401,N_19334);
nand U20907 (N_20907,N_19549,N_19079);
or U20908 (N_20908,N_19354,N_19673);
and U20909 (N_20909,N_19701,N_19666);
or U20910 (N_20910,N_19096,N_19577);
and U20911 (N_20911,N_19063,N_19846);
xor U20912 (N_20912,N_19043,N_19216);
and U20913 (N_20913,N_19389,N_19296);
and U20914 (N_20914,N_19934,N_19415);
nand U20915 (N_20915,N_19699,N_19546);
nor U20916 (N_20916,N_19813,N_19025);
nand U20917 (N_20917,N_19815,N_19765);
xor U20918 (N_20918,N_19311,N_19224);
and U20919 (N_20919,N_19137,N_19621);
xnor U20920 (N_20920,N_19702,N_19762);
nand U20921 (N_20921,N_19416,N_19433);
and U20922 (N_20922,N_19890,N_19908);
nor U20923 (N_20923,N_19966,N_19980);
and U20924 (N_20924,N_19642,N_19541);
nor U20925 (N_20925,N_19856,N_19454);
nor U20926 (N_20926,N_19003,N_19347);
xor U20927 (N_20927,N_19213,N_19639);
nor U20928 (N_20928,N_19236,N_19822);
nand U20929 (N_20929,N_19870,N_19935);
and U20930 (N_20930,N_19592,N_19251);
and U20931 (N_20931,N_19652,N_19920);
and U20932 (N_20932,N_19549,N_19183);
nor U20933 (N_20933,N_19107,N_19764);
nand U20934 (N_20934,N_19519,N_19562);
or U20935 (N_20935,N_19977,N_19345);
nand U20936 (N_20936,N_19916,N_19319);
nor U20937 (N_20937,N_19027,N_19465);
nand U20938 (N_20938,N_19994,N_19203);
and U20939 (N_20939,N_19204,N_19416);
xnor U20940 (N_20940,N_19553,N_19822);
nor U20941 (N_20941,N_19397,N_19244);
and U20942 (N_20942,N_19293,N_19156);
nand U20943 (N_20943,N_19512,N_19704);
and U20944 (N_20944,N_19347,N_19671);
nor U20945 (N_20945,N_19977,N_19329);
nand U20946 (N_20946,N_19416,N_19023);
and U20947 (N_20947,N_19126,N_19619);
nand U20948 (N_20948,N_19469,N_19647);
xor U20949 (N_20949,N_19521,N_19692);
or U20950 (N_20950,N_19989,N_19129);
xnor U20951 (N_20951,N_19931,N_19478);
nand U20952 (N_20952,N_19676,N_19850);
nand U20953 (N_20953,N_19097,N_19618);
nor U20954 (N_20954,N_19416,N_19788);
and U20955 (N_20955,N_19288,N_19198);
nand U20956 (N_20956,N_19461,N_19682);
or U20957 (N_20957,N_19486,N_19888);
xor U20958 (N_20958,N_19841,N_19280);
nand U20959 (N_20959,N_19270,N_19707);
nor U20960 (N_20960,N_19444,N_19346);
or U20961 (N_20961,N_19846,N_19402);
and U20962 (N_20962,N_19460,N_19366);
nand U20963 (N_20963,N_19713,N_19432);
or U20964 (N_20964,N_19818,N_19059);
xnor U20965 (N_20965,N_19648,N_19365);
and U20966 (N_20966,N_19848,N_19485);
nand U20967 (N_20967,N_19634,N_19264);
xor U20968 (N_20968,N_19357,N_19025);
xnor U20969 (N_20969,N_19387,N_19737);
nand U20970 (N_20970,N_19613,N_19459);
and U20971 (N_20971,N_19235,N_19186);
and U20972 (N_20972,N_19230,N_19528);
nor U20973 (N_20973,N_19380,N_19026);
xnor U20974 (N_20974,N_19589,N_19734);
and U20975 (N_20975,N_19592,N_19067);
xnor U20976 (N_20976,N_19560,N_19738);
nor U20977 (N_20977,N_19868,N_19730);
or U20978 (N_20978,N_19616,N_19737);
nor U20979 (N_20979,N_19567,N_19766);
xnor U20980 (N_20980,N_19587,N_19421);
xnor U20981 (N_20981,N_19798,N_19940);
or U20982 (N_20982,N_19088,N_19037);
and U20983 (N_20983,N_19414,N_19128);
nand U20984 (N_20984,N_19991,N_19911);
xor U20985 (N_20985,N_19359,N_19774);
or U20986 (N_20986,N_19409,N_19325);
and U20987 (N_20987,N_19702,N_19356);
nor U20988 (N_20988,N_19708,N_19450);
nor U20989 (N_20989,N_19257,N_19679);
nand U20990 (N_20990,N_19999,N_19023);
nand U20991 (N_20991,N_19545,N_19827);
or U20992 (N_20992,N_19672,N_19918);
nand U20993 (N_20993,N_19105,N_19861);
or U20994 (N_20994,N_19897,N_19104);
and U20995 (N_20995,N_19434,N_19816);
or U20996 (N_20996,N_19589,N_19283);
xnor U20997 (N_20997,N_19342,N_19154);
or U20998 (N_20998,N_19058,N_19563);
xor U20999 (N_20999,N_19666,N_19904);
xor U21000 (N_21000,N_20593,N_20959);
nand U21001 (N_21001,N_20394,N_20791);
xor U21002 (N_21002,N_20958,N_20182);
nor U21003 (N_21003,N_20592,N_20134);
nand U21004 (N_21004,N_20420,N_20555);
nor U21005 (N_21005,N_20240,N_20190);
and U21006 (N_21006,N_20434,N_20156);
nor U21007 (N_21007,N_20838,N_20108);
xnor U21008 (N_21008,N_20849,N_20680);
nand U21009 (N_21009,N_20109,N_20554);
nand U21010 (N_21010,N_20743,N_20327);
xor U21011 (N_21011,N_20759,N_20616);
nor U21012 (N_21012,N_20633,N_20149);
and U21013 (N_21013,N_20168,N_20550);
nor U21014 (N_21014,N_20102,N_20748);
or U21015 (N_21015,N_20423,N_20448);
nand U21016 (N_21016,N_20067,N_20021);
or U21017 (N_21017,N_20500,N_20981);
and U21018 (N_21018,N_20882,N_20489);
nor U21019 (N_21019,N_20010,N_20378);
xnor U21020 (N_21020,N_20294,N_20412);
nor U21021 (N_21021,N_20545,N_20407);
and U21022 (N_21022,N_20399,N_20160);
and U21023 (N_21023,N_20975,N_20558);
nand U21024 (N_21024,N_20047,N_20103);
nor U21025 (N_21025,N_20366,N_20185);
or U21026 (N_21026,N_20512,N_20145);
nand U21027 (N_21027,N_20004,N_20364);
xor U21028 (N_21028,N_20717,N_20721);
nand U21029 (N_21029,N_20792,N_20402);
nand U21030 (N_21030,N_20979,N_20330);
nor U21031 (N_21031,N_20628,N_20234);
nand U21032 (N_21032,N_20306,N_20629);
nand U21033 (N_21033,N_20175,N_20869);
nand U21034 (N_21034,N_20323,N_20169);
and U21035 (N_21035,N_20363,N_20510);
or U21036 (N_21036,N_20013,N_20615);
nor U21037 (N_21037,N_20850,N_20915);
xnor U21038 (N_21038,N_20964,N_20614);
or U21039 (N_21039,N_20579,N_20734);
or U21040 (N_21040,N_20447,N_20695);
or U21041 (N_21041,N_20204,N_20215);
nand U21042 (N_21042,N_20408,N_20427);
or U21043 (N_21043,N_20926,N_20119);
xnor U21044 (N_21044,N_20783,N_20426);
and U21045 (N_21045,N_20284,N_20546);
nor U21046 (N_21046,N_20884,N_20501);
xnor U21047 (N_21047,N_20523,N_20467);
nor U21048 (N_21048,N_20745,N_20502);
or U21049 (N_21049,N_20454,N_20425);
nand U21050 (N_21050,N_20329,N_20357);
xnor U21051 (N_21051,N_20821,N_20674);
xor U21052 (N_21052,N_20940,N_20410);
xnor U21053 (N_21053,N_20049,N_20273);
nor U21054 (N_21054,N_20075,N_20752);
or U21055 (N_21055,N_20538,N_20058);
and U21056 (N_21056,N_20729,N_20456);
nor U21057 (N_21057,N_20601,N_20564);
nand U21058 (N_21058,N_20604,N_20705);
and U21059 (N_21059,N_20391,N_20999);
nor U21060 (N_21060,N_20813,N_20380);
nand U21061 (N_21061,N_20794,N_20386);
xnor U21062 (N_21062,N_20480,N_20007);
or U21063 (N_21063,N_20080,N_20862);
xor U21064 (N_21064,N_20161,N_20889);
nor U21065 (N_21065,N_20507,N_20811);
nor U21066 (N_21066,N_20655,N_20074);
nor U21067 (N_21067,N_20126,N_20097);
nor U21068 (N_21068,N_20296,N_20218);
xor U21069 (N_21069,N_20219,N_20909);
or U21070 (N_21070,N_20223,N_20430);
and U21071 (N_21071,N_20228,N_20322);
nor U21072 (N_21072,N_20347,N_20871);
nor U21073 (N_21073,N_20266,N_20247);
or U21074 (N_21074,N_20693,N_20084);
or U21075 (N_21075,N_20667,N_20584);
or U21076 (N_21076,N_20398,N_20776);
xnor U21077 (N_21077,N_20362,N_20626);
and U21078 (N_21078,N_20388,N_20934);
xor U21079 (N_21079,N_20673,N_20005);
xnor U21080 (N_21080,N_20509,N_20451);
and U21081 (N_21081,N_20908,N_20775);
nor U21082 (N_21082,N_20553,N_20636);
nor U21083 (N_21083,N_20913,N_20848);
nand U21084 (N_21084,N_20853,N_20320);
nor U21085 (N_21085,N_20262,N_20582);
or U21086 (N_21086,N_20381,N_20290);
and U21087 (N_21087,N_20462,N_20722);
nand U21088 (N_21088,N_20551,N_20701);
nand U21089 (N_21089,N_20060,N_20491);
xor U21090 (N_21090,N_20498,N_20880);
and U21091 (N_21091,N_20755,N_20164);
or U21092 (N_21092,N_20267,N_20231);
or U21093 (N_21093,N_20805,N_20086);
xor U21094 (N_21094,N_20295,N_20860);
nor U21095 (N_21095,N_20872,N_20460);
nand U21096 (N_21096,N_20377,N_20640);
and U21097 (N_21097,N_20540,N_20968);
nor U21098 (N_21098,N_20736,N_20374);
and U21099 (N_21099,N_20799,N_20985);
nand U21100 (N_21100,N_20116,N_20072);
xnor U21101 (N_21101,N_20866,N_20779);
or U21102 (N_21102,N_20963,N_20369);
or U21103 (N_21103,N_20360,N_20300);
and U21104 (N_21104,N_20657,N_20099);
nand U21105 (N_21105,N_20230,N_20568);
and U21106 (N_21106,N_20557,N_20292);
nand U21107 (N_21107,N_20609,N_20733);
xnor U21108 (N_21108,N_20382,N_20669);
nand U21109 (N_21109,N_20651,N_20332);
nand U21110 (N_21110,N_20036,N_20587);
nand U21111 (N_21111,N_20948,N_20839);
xnor U21112 (N_21112,N_20343,N_20521);
nand U21113 (N_21113,N_20022,N_20982);
xnor U21114 (N_21114,N_20666,N_20191);
and U21115 (N_21115,N_20144,N_20907);
nand U21116 (N_21116,N_20571,N_20875);
nand U21117 (N_21117,N_20678,N_20668);
nand U21118 (N_21118,N_20508,N_20368);
or U21119 (N_21119,N_20073,N_20588);
and U21120 (N_21120,N_20814,N_20504);
or U21121 (N_21121,N_20416,N_20229);
nor U21122 (N_21122,N_20539,N_20112);
or U21123 (N_21123,N_20534,N_20921);
xnor U21124 (N_21124,N_20682,N_20123);
nor U21125 (N_21125,N_20561,N_20459);
and U21126 (N_21126,N_20146,N_20195);
or U21127 (N_21127,N_20000,N_20549);
nor U21128 (N_21128,N_20795,N_20727);
xnor U21129 (N_21129,N_20346,N_20591);
or U21130 (N_21130,N_20232,N_20034);
nand U21131 (N_21131,N_20663,N_20261);
xnor U21132 (N_21132,N_20253,N_20784);
nor U21133 (N_21133,N_20044,N_20291);
or U21134 (N_21134,N_20793,N_20763);
nand U21135 (N_21135,N_20068,N_20283);
and U21136 (N_21136,N_20024,N_20418);
xor U21137 (N_21137,N_20586,N_20048);
nand U21138 (N_21138,N_20248,N_20954);
xnor U21139 (N_21139,N_20438,N_20038);
nor U21140 (N_21140,N_20768,N_20379);
xor U21141 (N_21141,N_20245,N_20409);
nor U21142 (N_21142,N_20387,N_20861);
xnor U21143 (N_21143,N_20444,N_20192);
or U21144 (N_21144,N_20331,N_20809);
nor U21145 (N_21145,N_20688,N_20354);
xor U21146 (N_21146,N_20762,N_20313);
or U21147 (N_21147,N_20656,N_20879);
xnor U21148 (N_21148,N_20455,N_20213);
nor U21149 (N_21149,N_20702,N_20281);
nand U21150 (N_21150,N_20772,N_20578);
xnor U21151 (N_21151,N_20524,N_20599);
xnor U21152 (N_21152,N_20170,N_20713);
or U21153 (N_21153,N_20902,N_20453);
nand U21154 (N_21154,N_20585,N_20239);
xnor U21155 (N_21155,N_20339,N_20897);
nand U21156 (N_21156,N_20819,N_20874);
and U21157 (N_21157,N_20043,N_20096);
nor U21158 (N_21158,N_20457,N_20474);
nand U21159 (N_21159,N_20978,N_20530);
nor U21160 (N_21160,N_20856,N_20841);
and U21161 (N_21161,N_20827,N_20351);
nand U21162 (N_21162,N_20147,N_20644);
and U21163 (N_21163,N_20167,N_20596);
and U21164 (N_21164,N_20817,N_20015);
nor U21165 (N_21165,N_20417,N_20518);
nand U21166 (N_21166,N_20634,N_20194);
nand U21167 (N_21167,N_20531,N_20199);
nand U21168 (N_21168,N_20319,N_20970);
or U21169 (N_21169,N_20552,N_20843);
and U21170 (N_21170,N_20929,N_20259);
xor U21171 (N_21171,N_20962,N_20773);
xnor U21172 (N_21172,N_20172,N_20479);
and U21173 (N_21173,N_20488,N_20321);
nand U21174 (N_21174,N_20181,N_20898);
xnor U21175 (N_21175,N_20336,N_20730);
and U21176 (N_21176,N_20210,N_20804);
or U21177 (N_21177,N_20053,N_20490);
and U21178 (N_21178,N_20506,N_20282);
nor U21179 (N_21179,N_20355,N_20085);
nor U21180 (N_21180,N_20285,N_20404);
xor U21181 (N_21181,N_20422,N_20411);
nor U21182 (N_21182,N_20961,N_20868);
xor U21183 (N_21183,N_20774,N_20125);
nor U21184 (N_21184,N_20098,N_20661);
xor U21185 (N_21185,N_20101,N_20766);
nand U21186 (N_21186,N_20780,N_20260);
xnor U21187 (N_21187,N_20335,N_20625);
and U21188 (N_21188,N_20767,N_20939);
nor U21189 (N_21189,N_20649,N_20106);
nand U21190 (N_21190,N_20340,N_20415);
nor U21191 (N_21191,N_20243,N_20960);
or U21192 (N_21192,N_20050,N_20638);
or U21193 (N_21193,N_20001,N_20672);
nor U21194 (N_21194,N_20997,N_20069);
nor U21195 (N_21195,N_20188,N_20900);
nand U21196 (N_21196,N_20173,N_20694);
nand U21197 (N_21197,N_20706,N_20392);
or U21198 (N_21198,N_20764,N_20468);
and U21199 (N_21199,N_20641,N_20989);
nand U21200 (N_21200,N_20435,N_20837);
and U21201 (N_21201,N_20977,N_20692);
and U21202 (N_21202,N_20028,N_20439);
nand U21203 (N_21203,N_20133,N_20361);
nand U21204 (N_21204,N_20936,N_20761);
and U21205 (N_21205,N_20120,N_20304);
nor U21206 (N_21206,N_20946,N_20619);
nand U21207 (N_21207,N_20481,N_20603);
nand U21208 (N_21208,N_20252,N_20876);
nand U21209 (N_21209,N_20815,N_20345);
nand U21210 (N_21210,N_20808,N_20786);
and U21211 (N_21211,N_20225,N_20485);
and U21212 (N_21212,N_20716,N_20824);
and U21213 (N_21213,N_20520,N_20442);
nand U21214 (N_21214,N_20613,N_20428);
nand U21215 (N_21215,N_20174,N_20751);
xnor U21216 (N_21216,N_20831,N_20949);
and U21217 (N_21217,N_20041,N_20371);
and U21218 (N_21218,N_20206,N_20951);
or U21219 (N_21219,N_20810,N_20781);
or U21220 (N_21220,N_20567,N_20037);
or U21221 (N_21221,N_20476,N_20401);
nor U21222 (N_21222,N_20186,N_20054);
and U21223 (N_21223,N_20155,N_20574);
nand U21224 (N_21224,N_20264,N_20200);
nor U21225 (N_21225,N_20844,N_20527);
or U21226 (N_21226,N_20316,N_20857);
xnor U21227 (N_21227,N_20452,N_20042);
and U21228 (N_21228,N_20393,N_20424);
and U21229 (N_21229,N_20405,N_20492);
and U21230 (N_21230,N_20431,N_20464);
or U21231 (N_21231,N_20026,N_20986);
or U21232 (N_21232,N_20222,N_20632);
nor U21233 (N_21233,N_20516,N_20178);
nand U21234 (N_21234,N_20803,N_20272);
xnor U21235 (N_21235,N_20317,N_20542);
or U21236 (N_21236,N_20933,N_20529);
or U21237 (N_21237,N_20923,N_20893);
nor U21238 (N_21238,N_20870,N_20138);
nor U21239 (N_21239,N_20177,N_20016);
or U21240 (N_21240,N_20966,N_20890);
nand U21241 (N_21241,N_20910,N_20356);
nor U21242 (N_21242,N_20770,N_20494);
or U21243 (N_21243,N_20312,N_20255);
nor U21244 (N_21244,N_20718,N_20864);
or U21245 (N_21245,N_20639,N_20901);
or U21246 (N_21246,N_20279,N_20525);
and U21247 (N_21247,N_20214,N_20836);
nor U21248 (N_21248,N_20757,N_20895);
and U21249 (N_21249,N_20483,N_20136);
xnor U21250 (N_21250,N_20541,N_20569);
nand U21251 (N_21251,N_20517,N_20166);
or U21252 (N_21252,N_20113,N_20244);
nor U21253 (N_21253,N_20246,N_20238);
xor U21254 (N_21254,N_20974,N_20220);
xnor U21255 (N_21255,N_20432,N_20943);
nor U21256 (N_21256,N_20710,N_20737);
or U21257 (N_21257,N_20076,N_20056);
and U21258 (N_21258,N_20018,N_20196);
xor U21259 (N_21259,N_20227,N_20698);
nand U21260 (N_21260,N_20715,N_20265);
and U21261 (N_21261,N_20079,N_20445);
or U21262 (N_21262,N_20493,N_20338);
and U21263 (N_21263,N_20251,N_20973);
xor U21264 (N_21264,N_20159,N_20217);
nor U21265 (N_21265,N_20201,N_20699);
and U21266 (N_21266,N_20270,N_20132);
xnor U21267 (N_21267,N_20203,N_20040);
and U21268 (N_21268,N_20570,N_20091);
nor U21269 (N_21269,N_20746,N_20437);
and U21270 (N_21270,N_20122,N_20611);
xor U21271 (N_21271,N_20463,N_20288);
xor U21272 (N_21272,N_20709,N_20208);
nand U21273 (N_21273,N_20165,N_20528);
xor U21274 (N_21274,N_20675,N_20535);
xor U21275 (N_21275,N_20446,N_20664);
or U21276 (N_21276,N_20376,N_20139);
nand U21277 (N_21277,N_20278,N_20679);
or U21278 (N_21278,N_20903,N_20988);
nor U21279 (N_21279,N_20150,N_20148);
nor U21280 (N_21280,N_20691,N_20031);
xnor U21281 (N_21281,N_20575,N_20419);
and U21282 (N_21282,N_20092,N_20082);
or U21283 (N_21283,N_20724,N_20469);
or U21284 (N_21284,N_20620,N_20372);
nor U21285 (N_21285,N_20996,N_20179);
or U21286 (N_21286,N_20237,N_20742);
or U21287 (N_21287,N_20747,N_20344);
and U21288 (N_21288,N_20211,N_20153);
xor U21289 (N_21289,N_20956,N_20732);
or U21290 (N_21290,N_20057,N_20003);
nor U21291 (N_21291,N_20918,N_20497);
xor U21292 (N_21292,N_20832,N_20128);
or U21293 (N_21293,N_20070,N_20957);
nand U21294 (N_21294,N_20183,N_20565);
or U21295 (N_21295,N_20383,N_20482);
and U21296 (N_21296,N_20665,N_20274);
nand U21297 (N_21297,N_20928,N_20605);
or U21298 (N_21298,N_20293,N_20833);
nor U21299 (N_21299,N_20342,N_20127);
xnor U21300 (N_21300,N_20030,N_20250);
and U21301 (N_21301,N_20373,N_20580);
nand U21302 (N_21302,N_20140,N_20697);
and U21303 (N_21303,N_20515,N_20576);
xnor U21304 (N_21304,N_20847,N_20124);
nand U21305 (N_21305,N_20055,N_20078);
nor U21306 (N_21306,N_20107,N_20807);
xor U21307 (N_21307,N_20352,N_20820);
or U21308 (N_21308,N_20532,N_20257);
nor U21309 (N_21309,N_20443,N_20006);
nand U21310 (N_21310,N_20522,N_20413);
or U21311 (N_21311,N_20711,N_20750);
or U21312 (N_21312,N_20927,N_20287);
xor U21313 (N_21313,N_20104,N_20859);
or U21314 (N_21314,N_20242,N_20105);
and U21315 (N_21315,N_20806,N_20256);
xor U21316 (N_21316,N_20315,N_20471);
or U21317 (N_21317,N_20023,N_20142);
nand U21318 (N_21318,N_20461,N_20544);
or U21319 (N_21319,N_20931,N_20993);
nor U21320 (N_21320,N_20938,N_20618);
nand U21321 (N_21321,N_20135,N_20941);
or U21322 (N_21322,N_20712,N_20987);
or U21323 (N_21323,N_20881,N_20822);
and U21324 (N_21324,N_20912,N_20011);
xnor U21325 (N_21325,N_20624,N_20930);
and U21326 (N_21326,N_20790,N_20158);
and U21327 (N_21327,N_20189,N_20472);
nor U21328 (N_21328,N_20719,N_20513);
or U21329 (N_21329,N_20749,N_20466);
or U21330 (N_21330,N_20499,N_20458);
and U21331 (N_21331,N_20298,N_20090);
nor U21332 (N_21332,N_20741,N_20514);
xnor U21333 (N_21333,N_20235,N_20677);
or U21334 (N_21334,N_20914,N_20944);
nor U21335 (N_21335,N_20397,N_20162);
or U21336 (N_21336,N_20062,N_20690);
xnor U21337 (N_21337,N_20562,N_20911);
nor U21338 (N_21338,N_20789,N_20560);
and U21339 (N_21339,N_20268,N_20137);
nand U21340 (N_21340,N_20816,N_20899);
and U21341 (N_21341,N_20777,N_20171);
xnor U21342 (N_21342,N_20648,N_20904);
and U21343 (N_21343,N_20400,N_20314);
nand U21344 (N_21344,N_20796,N_20583);
nand U21345 (N_21345,N_20311,N_20846);
and U21346 (N_21346,N_20888,N_20801);
and U21347 (N_21347,N_20708,N_20349);
nor U21348 (N_21348,N_20297,N_20367);
nor U21349 (N_21349,N_20896,N_20704);
xor U21350 (N_21350,N_20917,N_20654);
xor U21351 (N_21351,N_20754,N_20365);
xnor U21352 (N_21352,N_20117,N_20787);
nor U21353 (N_21353,N_20765,N_20406);
xor U21354 (N_21354,N_20725,N_20925);
nor U21355 (N_21355,N_20051,N_20328);
and U21356 (N_21356,N_20830,N_20598);
or U21357 (N_21357,N_20867,N_20033);
or U21358 (N_21358,N_20589,N_20818);
and U21359 (N_21359,N_20543,N_20852);
xnor U21360 (N_21360,N_20646,N_20019);
nand U21361 (N_21361,N_20429,N_20151);
and U21362 (N_21362,N_20563,N_20025);
or U21363 (N_21363,N_20353,N_20647);
and U21364 (N_21364,N_20995,N_20505);
nor U21365 (N_21365,N_20039,N_20375);
nor U21366 (N_21366,N_20828,N_20612);
nor U21367 (N_21367,N_20045,N_20121);
xnor U21368 (N_21368,N_20280,N_20707);
or U21369 (N_21369,N_20660,N_20891);
nand U21370 (N_21370,N_20671,N_20029);
nor U21371 (N_21371,N_20157,N_20236);
xnor U21372 (N_21372,N_20334,N_20308);
and U21373 (N_21373,N_20083,N_20782);
nor U21374 (N_21374,N_20658,N_20731);
nand U21375 (N_21375,N_20622,N_20289);
xnor U21376 (N_21376,N_20953,N_20630);
or U21377 (N_21377,N_20797,N_20976);
xor U21378 (N_21378,N_20887,N_20299);
or U21379 (N_21379,N_20798,N_20046);
xor U21380 (N_21380,N_20714,N_20100);
xor U21381 (N_21381,N_20014,N_20617);
xnor U21382 (N_21382,N_20610,N_20920);
xnor U21383 (N_21383,N_20990,N_20325);
nand U21384 (N_21384,N_20686,N_20027);
and U21385 (N_21385,N_20275,N_20307);
and U21386 (N_21386,N_20855,N_20627);
nor U21387 (N_21387,N_20744,N_20081);
or U21388 (N_21388,N_20607,N_20684);
nor U21389 (N_21389,N_20301,N_20495);
or U21390 (N_21390,N_20998,N_20720);
or U21391 (N_21391,N_20597,N_20348);
xnor U21392 (N_21392,N_20905,N_20152);
nor U21393 (N_21393,N_20892,N_20785);
and U21394 (N_21394,N_20197,N_20723);
and U21395 (N_21395,N_20198,N_20703);
xnor U21396 (N_21396,N_20886,N_20536);
or U21397 (N_21397,N_20254,N_20935);
nor U21398 (N_21398,N_20478,N_20919);
or U21399 (N_21399,N_20676,N_20788);
nand U21400 (N_21400,N_20473,N_20114);
or U21401 (N_21401,N_20176,N_20756);
and U21402 (N_21402,N_20477,N_20577);
and U21403 (N_21403,N_20700,N_20358);
nor U21404 (N_21404,N_20623,N_20110);
nand U21405 (N_21405,N_20035,N_20590);
xor U21406 (N_21406,N_20318,N_20008);
or U21407 (N_21407,N_20854,N_20111);
and U21408 (N_21408,N_20350,N_20224);
nor U21409 (N_21409,N_20421,N_20249);
and U21410 (N_21410,N_20143,N_20594);
or U21411 (N_21411,N_20475,N_20258);
xnor U21412 (N_21412,N_20017,N_20631);
nand U21413 (N_21413,N_20696,N_20233);
nand U21414 (N_21414,N_20303,N_20450);
and U21415 (N_21415,N_20556,N_20606);
xnor U21416 (N_21416,N_20305,N_20118);
or U21417 (N_21417,N_20163,N_20269);
or U21418 (N_21418,N_20608,N_20826);
nand U21419 (N_21419,N_20942,N_20310);
nor U21420 (N_21420,N_20842,N_20865);
and U21421 (N_21421,N_20595,N_20263);
xor U21422 (N_21422,N_20771,N_20878);
and U21423 (N_21423,N_20971,N_20834);
nor U21424 (N_21424,N_20937,N_20945);
nand U21425 (N_21425,N_20685,N_20922);
or U21426 (N_21426,N_20071,N_20087);
xor U21427 (N_21427,N_20212,N_20093);
xor U21428 (N_21428,N_20753,N_20337);
nor U21429 (N_21429,N_20802,N_20980);
and U21430 (N_21430,N_20077,N_20645);
nand U21431 (N_21431,N_20012,N_20395);
nand U21432 (N_21432,N_20440,N_20950);
or U21433 (N_21433,N_20484,N_20825);
xor U21434 (N_21434,N_20065,N_20969);
nor U21435 (N_21435,N_20063,N_20687);
nor U21436 (N_21436,N_20728,N_20533);
nor U21437 (N_21437,N_20389,N_20449);
nor U21438 (N_21438,N_20370,N_20760);
nand U21439 (N_21439,N_20600,N_20681);
and U21440 (N_21440,N_20020,N_20095);
nand U21441 (N_21441,N_20835,N_20436);
or U21442 (N_21442,N_20559,N_20906);
or U21443 (N_21443,N_20286,N_20840);
nor U21444 (N_21444,N_20441,N_20851);
and U21445 (N_21445,N_20309,N_20984);
nand U21446 (N_21446,N_20863,N_20180);
nand U21447 (N_21447,N_20276,N_20566);
nor U21448 (N_21448,N_20226,N_20032);
nor U21449 (N_21449,N_20059,N_20581);
xor U21450 (N_21450,N_20187,N_20967);
nand U21451 (N_21451,N_20735,N_20873);
nor U21452 (N_21452,N_20740,N_20650);
xnor U21453 (N_21453,N_20129,N_20486);
nand U21454 (N_21454,N_20193,N_20652);
or U21455 (N_21455,N_20241,N_20052);
or U21456 (N_21456,N_20947,N_20829);
nor U21457 (N_21457,N_20738,N_20548);
nor U21458 (N_21458,N_20845,N_20972);
nand U21459 (N_21459,N_20202,N_20769);
nand U21460 (N_21460,N_20924,N_20916);
nor U21461 (N_21461,N_20009,N_20433);
xor U21462 (N_21462,N_20983,N_20184);
nor U21463 (N_21463,N_20643,N_20496);
or U21464 (N_21464,N_20130,N_20396);
nor U21465 (N_21465,N_20341,N_20662);
nor U21466 (N_21466,N_20894,N_20324);
and U21467 (N_21467,N_20390,N_20216);
or U21468 (N_21468,N_20739,N_20115);
and U21469 (N_21469,N_20885,N_20932);
or U21470 (N_21470,N_20670,N_20858);
xor U21471 (N_21471,N_20991,N_20088);
nor U21472 (N_21472,N_20511,N_20385);
nand U21473 (N_21473,N_20487,N_20205);
and U21474 (N_21474,N_20547,N_20519);
nor U21475 (N_21475,N_20465,N_20154);
or U21476 (N_21476,N_20002,N_20333);
and U21477 (N_21477,N_20621,N_20812);
and U21478 (N_21478,N_20326,N_20572);
and U21479 (N_21479,N_20141,N_20952);
or U21480 (N_21480,N_20221,N_20066);
nor U21481 (N_21481,N_20277,N_20089);
xnor U21482 (N_21482,N_20758,N_20537);
xnor U21483 (N_21483,N_20635,N_20094);
xnor U21484 (N_21484,N_20883,N_20994);
xnor U21485 (N_21485,N_20503,N_20414);
nor U21486 (N_21486,N_20726,N_20778);
and U21487 (N_21487,N_20131,N_20384);
nor U21488 (N_21488,N_20689,N_20637);
or U21489 (N_21489,N_20209,N_20877);
or U21490 (N_21490,N_20573,N_20965);
nand U21491 (N_21491,N_20271,N_20653);
xnor U21492 (N_21492,N_20470,N_20526);
or U21493 (N_21493,N_20659,N_20642);
or U21494 (N_21494,N_20823,N_20800);
or U21495 (N_21495,N_20683,N_20403);
or U21496 (N_21496,N_20061,N_20302);
nand U21497 (N_21497,N_20992,N_20207);
nor U21498 (N_21498,N_20359,N_20955);
nor U21499 (N_21499,N_20064,N_20602);
xor U21500 (N_21500,N_20258,N_20964);
xnor U21501 (N_21501,N_20943,N_20127);
xnor U21502 (N_21502,N_20117,N_20373);
and U21503 (N_21503,N_20277,N_20459);
nand U21504 (N_21504,N_20282,N_20476);
nand U21505 (N_21505,N_20218,N_20881);
xnor U21506 (N_21506,N_20666,N_20761);
and U21507 (N_21507,N_20059,N_20050);
and U21508 (N_21508,N_20223,N_20651);
or U21509 (N_21509,N_20108,N_20101);
nand U21510 (N_21510,N_20281,N_20046);
xnor U21511 (N_21511,N_20651,N_20356);
or U21512 (N_21512,N_20546,N_20847);
nand U21513 (N_21513,N_20831,N_20487);
nand U21514 (N_21514,N_20171,N_20302);
and U21515 (N_21515,N_20137,N_20869);
and U21516 (N_21516,N_20800,N_20825);
xor U21517 (N_21517,N_20848,N_20898);
nand U21518 (N_21518,N_20863,N_20507);
and U21519 (N_21519,N_20416,N_20748);
xor U21520 (N_21520,N_20210,N_20278);
or U21521 (N_21521,N_20784,N_20041);
nand U21522 (N_21522,N_20484,N_20236);
or U21523 (N_21523,N_20368,N_20250);
nand U21524 (N_21524,N_20026,N_20558);
nor U21525 (N_21525,N_20213,N_20952);
or U21526 (N_21526,N_20165,N_20413);
nand U21527 (N_21527,N_20423,N_20828);
and U21528 (N_21528,N_20555,N_20238);
nor U21529 (N_21529,N_20530,N_20692);
or U21530 (N_21530,N_20637,N_20937);
nor U21531 (N_21531,N_20212,N_20958);
nand U21532 (N_21532,N_20606,N_20795);
and U21533 (N_21533,N_20047,N_20774);
nand U21534 (N_21534,N_20290,N_20564);
nand U21535 (N_21535,N_20838,N_20685);
nor U21536 (N_21536,N_20770,N_20306);
xor U21537 (N_21537,N_20905,N_20744);
nor U21538 (N_21538,N_20002,N_20361);
xnor U21539 (N_21539,N_20582,N_20784);
or U21540 (N_21540,N_20951,N_20853);
and U21541 (N_21541,N_20720,N_20556);
nand U21542 (N_21542,N_20826,N_20596);
xnor U21543 (N_21543,N_20043,N_20809);
nand U21544 (N_21544,N_20677,N_20755);
nand U21545 (N_21545,N_20528,N_20548);
nand U21546 (N_21546,N_20055,N_20359);
nand U21547 (N_21547,N_20464,N_20594);
nor U21548 (N_21548,N_20791,N_20205);
and U21549 (N_21549,N_20022,N_20673);
nand U21550 (N_21550,N_20970,N_20785);
or U21551 (N_21551,N_20962,N_20820);
xnor U21552 (N_21552,N_20101,N_20958);
xor U21553 (N_21553,N_20399,N_20135);
and U21554 (N_21554,N_20735,N_20450);
or U21555 (N_21555,N_20823,N_20933);
or U21556 (N_21556,N_20076,N_20289);
nor U21557 (N_21557,N_20093,N_20708);
nor U21558 (N_21558,N_20096,N_20036);
or U21559 (N_21559,N_20977,N_20237);
nor U21560 (N_21560,N_20250,N_20588);
nand U21561 (N_21561,N_20638,N_20433);
and U21562 (N_21562,N_20563,N_20710);
or U21563 (N_21563,N_20251,N_20913);
nand U21564 (N_21564,N_20220,N_20751);
xor U21565 (N_21565,N_20112,N_20598);
nor U21566 (N_21566,N_20284,N_20020);
nor U21567 (N_21567,N_20466,N_20576);
or U21568 (N_21568,N_20342,N_20661);
and U21569 (N_21569,N_20419,N_20311);
or U21570 (N_21570,N_20296,N_20416);
and U21571 (N_21571,N_20647,N_20763);
and U21572 (N_21572,N_20957,N_20689);
or U21573 (N_21573,N_20402,N_20767);
nand U21574 (N_21574,N_20190,N_20160);
or U21575 (N_21575,N_20707,N_20658);
nand U21576 (N_21576,N_20471,N_20573);
xnor U21577 (N_21577,N_20766,N_20210);
nor U21578 (N_21578,N_20158,N_20344);
or U21579 (N_21579,N_20532,N_20583);
nor U21580 (N_21580,N_20152,N_20373);
and U21581 (N_21581,N_20178,N_20601);
nor U21582 (N_21582,N_20902,N_20511);
nor U21583 (N_21583,N_20224,N_20868);
and U21584 (N_21584,N_20836,N_20464);
or U21585 (N_21585,N_20793,N_20572);
and U21586 (N_21586,N_20841,N_20313);
and U21587 (N_21587,N_20733,N_20155);
nor U21588 (N_21588,N_20231,N_20848);
xnor U21589 (N_21589,N_20972,N_20507);
nor U21590 (N_21590,N_20668,N_20069);
xnor U21591 (N_21591,N_20557,N_20372);
nand U21592 (N_21592,N_20398,N_20028);
nand U21593 (N_21593,N_20751,N_20135);
nand U21594 (N_21594,N_20726,N_20458);
or U21595 (N_21595,N_20935,N_20588);
xor U21596 (N_21596,N_20094,N_20937);
or U21597 (N_21597,N_20245,N_20196);
and U21598 (N_21598,N_20492,N_20863);
nor U21599 (N_21599,N_20467,N_20521);
nand U21600 (N_21600,N_20933,N_20938);
and U21601 (N_21601,N_20892,N_20982);
or U21602 (N_21602,N_20246,N_20637);
and U21603 (N_21603,N_20207,N_20957);
nand U21604 (N_21604,N_20124,N_20946);
and U21605 (N_21605,N_20954,N_20112);
or U21606 (N_21606,N_20571,N_20770);
and U21607 (N_21607,N_20022,N_20893);
or U21608 (N_21608,N_20343,N_20026);
nor U21609 (N_21609,N_20524,N_20159);
or U21610 (N_21610,N_20335,N_20175);
xnor U21611 (N_21611,N_20146,N_20404);
and U21612 (N_21612,N_20748,N_20055);
nor U21613 (N_21613,N_20211,N_20315);
or U21614 (N_21614,N_20743,N_20408);
xor U21615 (N_21615,N_20121,N_20364);
or U21616 (N_21616,N_20911,N_20407);
or U21617 (N_21617,N_20283,N_20812);
nand U21618 (N_21618,N_20445,N_20287);
xnor U21619 (N_21619,N_20833,N_20635);
nor U21620 (N_21620,N_20806,N_20018);
nor U21621 (N_21621,N_20287,N_20749);
or U21622 (N_21622,N_20429,N_20013);
nand U21623 (N_21623,N_20894,N_20167);
and U21624 (N_21624,N_20510,N_20880);
nand U21625 (N_21625,N_20340,N_20083);
nor U21626 (N_21626,N_20416,N_20152);
nand U21627 (N_21627,N_20890,N_20532);
nor U21628 (N_21628,N_20940,N_20203);
nor U21629 (N_21629,N_20360,N_20047);
or U21630 (N_21630,N_20254,N_20165);
xor U21631 (N_21631,N_20950,N_20138);
xnor U21632 (N_21632,N_20852,N_20275);
nor U21633 (N_21633,N_20048,N_20986);
nor U21634 (N_21634,N_20801,N_20573);
nand U21635 (N_21635,N_20465,N_20998);
nand U21636 (N_21636,N_20588,N_20799);
nor U21637 (N_21637,N_20759,N_20036);
and U21638 (N_21638,N_20182,N_20909);
xnor U21639 (N_21639,N_20979,N_20795);
nand U21640 (N_21640,N_20954,N_20450);
nor U21641 (N_21641,N_20626,N_20434);
and U21642 (N_21642,N_20894,N_20011);
nand U21643 (N_21643,N_20727,N_20510);
nor U21644 (N_21644,N_20475,N_20093);
nand U21645 (N_21645,N_20232,N_20809);
and U21646 (N_21646,N_20334,N_20667);
nor U21647 (N_21647,N_20794,N_20561);
nor U21648 (N_21648,N_20003,N_20571);
nor U21649 (N_21649,N_20262,N_20471);
and U21650 (N_21650,N_20970,N_20365);
xor U21651 (N_21651,N_20991,N_20357);
nor U21652 (N_21652,N_20452,N_20847);
and U21653 (N_21653,N_20616,N_20894);
nand U21654 (N_21654,N_20510,N_20171);
nor U21655 (N_21655,N_20716,N_20912);
xor U21656 (N_21656,N_20747,N_20923);
nand U21657 (N_21657,N_20502,N_20317);
or U21658 (N_21658,N_20528,N_20449);
or U21659 (N_21659,N_20945,N_20164);
or U21660 (N_21660,N_20726,N_20733);
nand U21661 (N_21661,N_20544,N_20429);
or U21662 (N_21662,N_20263,N_20293);
and U21663 (N_21663,N_20342,N_20509);
or U21664 (N_21664,N_20479,N_20240);
nand U21665 (N_21665,N_20644,N_20990);
xor U21666 (N_21666,N_20490,N_20800);
and U21667 (N_21667,N_20357,N_20021);
nor U21668 (N_21668,N_20140,N_20292);
nand U21669 (N_21669,N_20717,N_20067);
xor U21670 (N_21670,N_20496,N_20806);
and U21671 (N_21671,N_20741,N_20604);
nand U21672 (N_21672,N_20120,N_20380);
nor U21673 (N_21673,N_20433,N_20806);
nor U21674 (N_21674,N_20187,N_20697);
and U21675 (N_21675,N_20644,N_20317);
or U21676 (N_21676,N_20350,N_20489);
nand U21677 (N_21677,N_20985,N_20902);
nand U21678 (N_21678,N_20130,N_20113);
nand U21679 (N_21679,N_20249,N_20172);
nand U21680 (N_21680,N_20686,N_20926);
or U21681 (N_21681,N_20579,N_20129);
nor U21682 (N_21682,N_20874,N_20164);
and U21683 (N_21683,N_20162,N_20944);
nand U21684 (N_21684,N_20677,N_20282);
nor U21685 (N_21685,N_20047,N_20602);
xnor U21686 (N_21686,N_20265,N_20951);
xor U21687 (N_21687,N_20618,N_20082);
or U21688 (N_21688,N_20055,N_20637);
nand U21689 (N_21689,N_20020,N_20826);
nor U21690 (N_21690,N_20848,N_20579);
nand U21691 (N_21691,N_20369,N_20742);
nor U21692 (N_21692,N_20556,N_20021);
nand U21693 (N_21693,N_20411,N_20398);
xor U21694 (N_21694,N_20243,N_20904);
xnor U21695 (N_21695,N_20496,N_20770);
xor U21696 (N_21696,N_20531,N_20745);
and U21697 (N_21697,N_20427,N_20690);
xnor U21698 (N_21698,N_20914,N_20922);
or U21699 (N_21699,N_20983,N_20762);
or U21700 (N_21700,N_20556,N_20000);
nor U21701 (N_21701,N_20492,N_20476);
nand U21702 (N_21702,N_20424,N_20963);
nor U21703 (N_21703,N_20232,N_20627);
or U21704 (N_21704,N_20855,N_20351);
or U21705 (N_21705,N_20415,N_20427);
or U21706 (N_21706,N_20731,N_20886);
and U21707 (N_21707,N_20090,N_20699);
or U21708 (N_21708,N_20923,N_20287);
nor U21709 (N_21709,N_20091,N_20527);
nor U21710 (N_21710,N_20413,N_20468);
nand U21711 (N_21711,N_20801,N_20493);
xor U21712 (N_21712,N_20274,N_20976);
or U21713 (N_21713,N_20683,N_20301);
and U21714 (N_21714,N_20759,N_20199);
or U21715 (N_21715,N_20741,N_20504);
and U21716 (N_21716,N_20847,N_20571);
or U21717 (N_21717,N_20458,N_20913);
and U21718 (N_21718,N_20103,N_20124);
nand U21719 (N_21719,N_20134,N_20878);
or U21720 (N_21720,N_20833,N_20830);
xnor U21721 (N_21721,N_20366,N_20056);
nand U21722 (N_21722,N_20025,N_20775);
and U21723 (N_21723,N_20997,N_20279);
nor U21724 (N_21724,N_20150,N_20513);
nor U21725 (N_21725,N_20648,N_20256);
or U21726 (N_21726,N_20873,N_20887);
or U21727 (N_21727,N_20454,N_20346);
and U21728 (N_21728,N_20573,N_20781);
or U21729 (N_21729,N_20205,N_20556);
xnor U21730 (N_21730,N_20288,N_20224);
nand U21731 (N_21731,N_20314,N_20479);
xnor U21732 (N_21732,N_20419,N_20993);
or U21733 (N_21733,N_20871,N_20191);
nor U21734 (N_21734,N_20959,N_20042);
or U21735 (N_21735,N_20856,N_20889);
nand U21736 (N_21736,N_20280,N_20316);
xor U21737 (N_21737,N_20453,N_20917);
xnor U21738 (N_21738,N_20519,N_20846);
and U21739 (N_21739,N_20015,N_20581);
or U21740 (N_21740,N_20112,N_20335);
xnor U21741 (N_21741,N_20881,N_20223);
xnor U21742 (N_21742,N_20538,N_20150);
and U21743 (N_21743,N_20303,N_20127);
xor U21744 (N_21744,N_20659,N_20459);
xor U21745 (N_21745,N_20868,N_20965);
nand U21746 (N_21746,N_20411,N_20878);
or U21747 (N_21747,N_20865,N_20185);
or U21748 (N_21748,N_20438,N_20138);
and U21749 (N_21749,N_20183,N_20538);
nand U21750 (N_21750,N_20090,N_20446);
nor U21751 (N_21751,N_20299,N_20945);
or U21752 (N_21752,N_20972,N_20796);
nor U21753 (N_21753,N_20945,N_20614);
nand U21754 (N_21754,N_20842,N_20881);
or U21755 (N_21755,N_20517,N_20142);
nand U21756 (N_21756,N_20770,N_20329);
xnor U21757 (N_21757,N_20742,N_20323);
nand U21758 (N_21758,N_20410,N_20515);
nand U21759 (N_21759,N_20427,N_20046);
and U21760 (N_21760,N_20883,N_20348);
nand U21761 (N_21761,N_20612,N_20244);
and U21762 (N_21762,N_20005,N_20513);
or U21763 (N_21763,N_20865,N_20059);
nor U21764 (N_21764,N_20168,N_20484);
or U21765 (N_21765,N_20715,N_20778);
xnor U21766 (N_21766,N_20698,N_20479);
and U21767 (N_21767,N_20018,N_20936);
nand U21768 (N_21768,N_20529,N_20394);
and U21769 (N_21769,N_20998,N_20718);
nand U21770 (N_21770,N_20702,N_20219);
nand U21771 (N_21771,N_20443,N_20198);
xor U21772 (N_21772,N_20836,N_20388);
nand U21773 (N_21773,N_20759,N_20462);
xor U21774 (N_21774,N_20150,N_20152);
xnor U21775 (N_21775,N_20584,N_20638);
and U21776 (N_21776,N_20660,N_20635);
or U21777 (N_21777,N_20834,N_20492);
nor U21778 (N_21778,N_20223,N_20557);
nand U21779 (N_21779,N_20439,N_20431);
or U21780 (N_21780,N_20284,N_20630);
or U21781 (N_21781,N_20727,N_20541);
nand U21782 (N_21782,N_20518,N_20547);
and U21783 (N_21783,N_20549,N_20302);
or U21784 (N_21784,N_20937,N_20309);
nor U21785 (N_21785,N_20922,N_20991);
and U21786 (N_21786,N_20037,N_20798);
and U21787 (N_21787,N_20486,N_20531);
or U21788 (N_21788,N_20709,N_20339);
and U21789 (N_21789,N_20772,N_20646);
nor U21790 (N_21790,N_20469,N_20340);
or U21791 (N_21791,N_20018,N_20894);
xor U21792 (N_21792,N_20768,N_20216);
xnor U21793 (N_21793,N_20719,N_20291);
xor U21794 (N_21794,N_20909,N_20941);
nand U21795 (N_21795,N_20462,N_20141);
or U21796 (N_21796,N_20653,N_20397);
xor U21797 (N_21797,N_20406,N_20600);
nand U21798 (N_21798,N_20277,N_20848);
xor U21799 (N_21799,N_20245,N_20671);
or U21800 (N_21800,N_20034,N_20270);
nand U21801 (N_21801,N_20031,N_20415);
and U21802 (N_21802,N_20798,N_20060);
nor U21803 (N_21803,N_20637,N_20628);
or U21804 (N_21804,N_20320,N_20759);
or U21805 (N_21805,N_20674,N_20538);
and U21806 (N_21806,N_20322,N_20737);
and U21807 (N_21807,N_20711,N_20046);
or U21808 (N_21808,N_20075,N_20640);
nor U21809 (N_21809,N_20257,N_20202);
or U21810 (N_21810,N_20507,N_20142);
nor U21811 (N_21811,N_20350,N_20857);
nand U21812 (N_21812,N_20617,N_20493);
xnor U21813 (N_21813,N_20187,N_20633);
nor U21814 (N_21814,N_20992,N_20476);
nand U21815 (N_21815,N_20445,N_20005);
and U21816 (N_21816,N_20186,N_20842);
nor U21817 (N_21817,N_20069,N_20869);
or U21818 (N_21818,N_20335,N_20763);
and U21819 (N_21819,N_20406,N_20588);
xnor U21820 (N_21820,N_20827,N_20223);
and U21821 (N_21821,N_20367,N_20764);
nand U21822 (N_21822,N_20650,N_20306);
nand U21823 (N_21823,N_20780,N_20831);
nor U21824 (N_21824,N_20057,N_20327);
and U21825 (N_21825,N_20743,N_20934);
and U21826 (N_21826,N_20708,N_20255);
xnor U21827 (N_21827,N_20230,N_20776);
or U21828 (N_21828,N_20453,N_20966);
nand U21829 (N_21829,N_20711,N_20247);
nor U21830 (N_21830,N_20310,N_20921);
nor U21831 (N_21831,N_20728,N_20606);
nand U21832 (N_21832,N_20086,N_20401);
and U21833 (N_21833,N_20483,N_20564);
nand U21834 (N_21834,N_20984,N_20303);
nor U21835 (N_21835,N_20085,N_20346);
nor U21836 (N_21836,N_20500,N_20686);
and U21837 (N_21837,N_20364,N_20655);
nor U21838 (N_21838,N_20151,N_20761);
or U21839 (N_21839,N_20143,N_20103);
and U21840 (N_21840,N_20257,N_20237);
nand U21841 (N_21841,N_20282,N_20733);
xnor U21842 (N_21842,N_20337,N_20338);
and U21843 (N_21843,N_20834,N_20262);
nor U21844 (N_21844,N_20805,N_20716);
or U21845 (N_21845,N_20730,N_20950);
nand U21846 (N_21846,N_20070,N_20045);
or U21847 (N_21847,N_20515,N_20814);
nand U21848 (N_21848,N_20949,N_20733);
nor U21849 (N_21849,N_20848,N_20884);
or U21850 (N_21850,N_20516,N_20673);
nor U21851 (N_21851,N_20444,N_20847);
nor U21852 (N_21852,N_20190,N_20591);
or U21853 (N_21853,N_20994,N_20356);
nand U21854 (N_21854,N_20497,N_20992);
or U21855 (N_21855,N_20918,N_20289);
or U21856 (N_21856,N_20834,N_20610);
and U21857 (N_21857,N_20385,N_20865);
xnor U21858 (N_21858,N_20033,N_20716);
xnor U21859 (N_21859,N_20984,N_20897);
and U21860 (N_21860,N_20405,N_20361);
and U21861 (N_21861,N_20069,N_20237);
and U21862 (N_21862,N_20048,N_20100);
nor U21863 (N_21863,N_20504,N_20277);
nand U21864 (N_21864,N_20629,N_20593);
nand U21865 (N_21865,N_20540,N_20440);
nand U21866 (N_21866,N_20303,N_20888);
nor U21867 (N_21867,N_20371,N_20241);
nor U21868 (N_21868,N_20812,N_20265);
or U21869 (N_21869,N_20026,N_20165);
and U21870 (N_21870,N_20047,N_20655);
and U21871 (N_21871,N_20014,N_20307);
nor U21872 (N_21872,N_20288,N_20069);
and U21873 (N_21873,N_20976,N_20784);
xnor U21874 (N_21874,N_20271,N_20900);
nand U21875 (N_21875,N_20553,N_20085);
xnor U21876 (N_21876,N_20928,N_20260);
and U21877 (N_21877,N_20242,N_20351);
xnor U21878 (N_21878,N_20335,N_20780);
nand U21879 (N_21879,N_20724,N_20294);
nand U21880 (N_21880,N_20401,N_20856);
nor U21881 (N_21881,N_20406,N_20499);
nor U21882 (N_21882,N_20381,N_20576);
or U21883 (N_21883,N_20062,N_20857);
xnor U21884 (N_21884,N_20566,N_20248);
xor U21885 (N_21885,N_20214,N_20826);
or U21886 (N_21886,N_20332,N_20767);
nor U21887 (N_21887,N_20811,N_20735);
nand U21888 (N_21888,N_20355,N_20956);
xnor U21889 (N_21889,N_20246,N_20282);
xor U21890 (N_21890,N_20624,N_20905);
nand U21891 (N_21891,N_20986,N_20145);
nand U21892 (N_21892,N_20897,N_20167);
or U21893 (N_21893,N_20405,N_20927);
xor U21894 (N_21894,N_20280,N_20071);
nor U21895 (N_21895,N_20770,N_20553);
nor U21896 (N_21896,N_20320,N_20180);
nand U21897 (N_21897,N_20334,N_20754);
and U21898 (N_21898,N_20567,N_20484);
nand U21899 (N_21899,N_20363,N_20724);
or U21900 (N_21900,N_20718,N_20189);
and U21901 (N_21901,N_20262,N_20607);
and U21902 (N_21902,N_20528,N_20969);
and U21903 (N_21903,N_20213,N_20780);
xor U21904 (N_21904,N_20884,N_20508);
and U21905 (N_21905,N_20284,N_20155);
xnor U21906 (N_21906,N_20830,N_20462);
nand U21907 (N_21907,N_20053,N_20876);
nor U21908 (N_21908,N_20778,N_20326);
or U21909 (N_21909,N_20263,N_20650);
nor U21910 (N_21910,N_20134,N_20716);
xnor U21911 (N_21911,N_20052,N_20228);
nand U21912 (N_21912,N_20414,N_20444);
nand U21913 (N_21913,N_20509,N_20911);
xnor U21914 (N_21914,N_20048,N_20993);
and U21915 (N_21915,N_20170,N_20743);
and U21916 (N_21916,N_20296,N_20866);
or U21917 (N_21917,N_20850,N_20856);
or U21918 (N_21918,N_20638,N_20494);
nand U21919 (N_21919,N_20067,N_20790);
nand U21920 (N_21920,N_20908,N_20647);
or U21921 (N_21921,N_20816,N_20608);
or U21922 (N_21922,N_20307,N_20407);
or U21923 (N_21923,N_20066,N_20012);
nand U21924 (N_21924,N_20309,N_20690);
nand U21925 (N_21925,N_20187,N_20374);
xor U21926 (N_21926,N_20154,N_20048);
and U21927 (N_21927,N_20553,N_20587);
or U21928 (N_21928,N_20497,N_20287);
nand U21929 (N_21929,N_20835,N_20676);
nand U21930 (N_21930,N_20204,N_20485);
and U21931 (N_21931,N_20591,N_20595);
nor U21932 (N_21932,N_20479,N_20332);
and U21933 (N_21933,N_20267,N_20295);
nor U21934 (N_21934,N_20779,N_20765);
nor U21935 (N_21935,N_20459,N_20341);
nand U21936 (N_21936,N_20482,N_20266);
or U21937 (N_21937,N_20441,N_20673);
and U21938 (N_21938,N_20727,N_20357);
nor U21939 (N_21939,N_20869,N_20768);
nand U21940 (N_21940,N_20542,N_20336);
xor U21941 (N_21941,N_20112,N_20017);
xor U21942 (N_21942,N_20400,N_20473);
and U21943 (N_21943,N_20469,N_20428);
xnor U21944 (N_21944,N_20529,N_20686);
nand U21945 (N_21945,N_20080,N_20775);
and U21946 (N_21946,N_20414,N_20746);
or U21947 (N_21947,N_20120,N_20657);
nand U21948 (N_21948,N_20086,N_20566);
and U21949 (N_21949,N_20572,N_20993);
and U21950 (N_21950,N_20646,N_20784);
nand U21951 (N_21951,N_20651,N_20978);
nor U21952 (N_21952,N_20781,N_20491);
nand U21953 (N_21953,N_20874,N_20791);
nand U21954 (N_21954,N_20890,N_20001);
or U21955 (N_21955,N_20306,N_20733);
or U21956 (N_21956,N_20490,N_20643);
and U21957 (N_21957,N_20032,N_20114);
xnor U21958 (N_21958,N_20889,N_20787);
xor U21959 (N_21959,N_20102,N_20201);
nand U21960 (N_21960,N_20584,N_20698);
and U21961 (N_21961,N_20683,N_20276);
and U21962 (N_21962,N_20857,N_20842);
and U21963 (N_21963,N_20977,N_20776);
or U21964 (N_21964,N_20040,N_20822);
and U21965 (N_21965,N_20275,N_20438);
nor U21966 (N_21966,N_20915,N_20111);
xnor U21967 (N_21967,N_20967,N_20759);
nor U21968 (N_21968,N_20642,N_20311);
nand U21969 (N_21969,N_20637,N_20949);
nand U21970 (N_21970,N_20621,N_20589);
nor U21971 (N_21971,N_20471,N_20697);
nor U21972 (N_21972,N_20944,N_20533);
or U21973 (N_21973,N_20697,N_20080);
nor U21974 (N_21974,N_20152,N_20102);
nor U21975 (N_21975,N_20549,N_20797);
xnor U21976 (N_21976,N_20868,N_20880);
and U21977 (N_21977,N_20886,N_20814);
nor U21978 (N_21978,N_20832,N_20891);
xnor U21979 (N_21979,N_20800,N_20041);
xnor U21980 (N_21980,N_20853,N_20945);
nand U21981 (N_21981,N_20793,N_20711);
or U21982 (N_21982,N_20322,N_20093);
nor U21983 (N_21983,N_20150,N_20683);
xor U21984 (N_21984,N_20613,N_20220);
or U21985 (N_21985,N_20620,N_20762);
nand U21986 (N_21986,N_20207,N_20055);
nand U21987 (N_21987,N_20678,N_20733);
nand U21988 (N_21988,N_20830,N_20677);
and U21989 (N_21989,N_20702,N_20107);
nand U21990 (N_21990,N_20974,N_20711);
or U21991 (N_21991,N_20314,N_20631);
xor U21992 (N_21992,N_20878,N_20856);
nor U21993 (N_21993,N_20609,N_20970);
and U21994 (N_21994,N_20009,N_20754);
xor U21995 (N_21995,N_20692,N_20208);
xnor U21996 (N_21996,N_20018,N_20586);
or U21997 (N_21997,N_20522,N_20333);
nor U21998 (N_21998,N_20568,N_20059);
nor U21999 (N_21999,N_20729,N_20664);
nand U22000 (N_22000,N_21556,N_21999);
nor U22001 (N_22001,N_21872,N_21978);
or U22002 (N_22002,N_21738,N_21963);
and U22003 (N_22003,N_21064,N_21759);
xnor U22004 (N_22004,N_21722,N_21029);
nand U22005 (N_22005,N_21338,N_21093);
or U22006 (N_22006,N_21377,N_21318);
xnor U22007 (N_22007,N_21502,N_21256);
nand U22008 (N_22008,N_21662,N_21208);
or U22009 (N_22009,N_21292,N_21816);
nor U22010 (N_22010,N_21238,N_21656);
nand U22011 (N_22011,N_21883,N_21640);
nor U22012 (N_22012,N_21427,N_21515);
xor U22013 (N_22013,N_21776,N_21688);
nand U22014 (N_22014,N_21651,N_21448);
nor U22015 (N_22015,N_21658,N_21231);
nand U22016 (N_22016,N_21060,N_21406);
or U22017 (N_22017,N_21701,N_21416);
xnor U22018 (N_22018,N_21123,N_21160);
or U22019 (N_22019,N_21714,N_21798);
xor U22020 (N_22020,N_21127,N_21147);
nand U22021 (N_22021,N_21576,N_21201);
xnor U22022 (N_22022,N_21339,N_21789);
xor U22023 (N_22023,N_21811,N_21285);
nand U22024 (N_22024,N_21196,N_21943);
or U22025 (N_22025,N_21321,N_21846);
xor U22026 (N_22026,N_21859,N_21895);
nor U22027 (N_22027,N_21408,N_21158);
and U22028 (N_22028,N_21031,N_21597);
xnor U22029 (N_22029,N_21362,N_21004);
and U22030 (N_22030,N_21552,N_21211);
xor U22031 (N_22031,N_21352,N_21777);
xnor U22032 (N_22032,N_21126,N_21180);
or U22033 (N_22033,N_21849,N_21232);
nor U22034 (N_22034,N_21258,N_21106);
nand U22035 (N_22035,N_21069,N_21546);
or U22036 (N_22036,N_21359,N_21372);
or U22037 (N_22037,N_21964,N_21644);
nand U22038 (N_22038,N_21979,N_21760);
or U22039 (N_22039,N_21888,N_21508);
xor U22040 (N_22040,N_21272,N_21025);
or U22041 (N_22041,N_21466,N_21353);
nand U22042 (N_22042,N_21451,N_21298);
xor U22043 (N_22043,N_21428,N_21340);
and U22044 (N_22044,N_21347,N_21643);
nand U22045 (N_22045,N_21542,N_21354);
xor U22046 (N_22046,N_21941,N_21570);
xor U22047 (N_22047,N_21740,N_21728);
or U22048 (N_22048,N_21115,N_21003);
or U22049 (N_22049,N_21048,N_21241);
nor U22050 (N_22050,N_21631,N_21244);
xnor U22051 (N_22051,N_21344,N_21161);
or U22052 (N_22052,N_21938,N_21381);
or U22053 (N_22053,N_21269,N_21898);
or U22054 (N_22054,N_21976,N_21178);
nor U22055 (N_22055,N_21392,N_21483);
nor U22056 (N_22056,N_21578,N_21215);
nor U22057 (N_22057,N_21450,N_21748);
nand U22058 (N_22058,N_21476,N_21646);
nor U22059 (N_22059,N_21179,N_21489);
xor U22060 (N_22060,N_21854,N_21249);
nor U22061 (N_22061,N_21595,N_21418);
nand U22062 (N_22062,N_21128,N_21493);
nor U22063 (N_22063,N_21246,N_21663);
or U22064 (N_22064,N_21781,N_21757);
nand U22065 (N_22065,N_21844,N_21625);
or U22066 (N_22066,N_21474,N_21412);
xnor U22067 (N_22067,N_21561,N_21050);
nand U22068 (N_22068,N_21763,N_21495);
xor U22069 (N_22069,N_21810,N_21548);
nand U22070 (N_22070,N_21108,N_21700);
and U22071 (N_22071,N_21582,N_21946);
xor U22072 (N_22072,N_21016,N_21132);
and U22073 (N_22073,N_21614,N_21709);
nor U22074 (N_22074,N_21809,N_21299);
nand U22075 (N_22075,N_21655,N_21873);
xor U22076 (N_22076,N_21550,N_21762);
nand U22077 (N_22077,N_21681,N_21358);
nand U22078 (N_22078,N_21420,N_21991);
xnor U22079 (N_22079,N_21937,N_21779);
nand U22080 (N_22080,N_21112,N_21404);
nor U22081 (N_22081,N_21829,N_21784);
nor U22082 (N_22082,N_21150,N_21113);
xor U22083 (N_22083,N_21671,N_21910);
and U22084 (N_22084,N_21635,N_21346);
or U22085 (N_22085,N_21472,N_21511);
nor U22086 (N_22086,N_21972,N_21695);
and U22087 (N_22087,N_21350,N_21257);
xnor U22088 (N_22088,N_21438,N_21773);
or U22089 (N_22089,N_21812,N_21345);
or U22090 (N_22090,N_21043,N_21044);
or U22091 (N_22091,N_21806,N_21574);
nor U22092 (N_22092,N_21716,N_21379);
nor U22093 (N_22093,N_21666,N_21205);
nor U22094 (N_22094,N_21554,N_21698);
or U22095 (N_22095,N_21683,N_21731);
and U22096 (N_22096,N_21385,N_21324);
nand U22097 (N_22097,N_21817,N_21772);
nor U22098 (N_22098,N_21674,N_21694);
nor U22099 (N_22099,N_21620,N_21530);
and U22100 (N_22100,N_21442,N_21302);
nor U22101 (N_22101,N_21818,N_21587);
or U22102 (N_22102,N_21068,N_21726);
and U22103 (N_22103,N_21154,N_21797);
nor U22104 (N_22104,N_21930,N_21611);
nor U22105 (N_22105,N_21920,N_21725);
nand U22106 (N_22106,N_21390,N_21973);
or U22107 (N_22107,N_21330,N_21949);
xor U22108 (N_22108,N_21743,N_21053);
and U22109 (N_22109,N_21838,N_21107);
nor U22110 (N_22110,N_21761,N_21851);
nand U22111 (N_22111,N_21423,N_21672);
nor U22112 (N_22112,N_21081,N_21553);
and U22113 (N_22113,N_21363,N_21922);
or U22114 (N_22114,N_21366,N_21952);
nand U22115 (N_22115,N_21045,N_21936);
and U22116 (N_22116,N_21724,N_21300);
xnor U22117 (N_22117,N_21456,N_21690);
nor U22118 (N_22118,N_21075,N_21268);
nor U22119 (N_22119,N_21932,N_21230);
xor U22120 (N_22120,N_21320,N_21543);
and U22121 (N_22121,N_21845,N_21368);
and U22122 (N_22122,N_21110,N_21109);
or U22123 (N_22123,N_21415,N_21296);
and U22124 (N_22124,N_21317,N_21692);
nand U22125 (N_22125,N_21233,N_21284);
xor U22126 (N_22126,N_21008,N_21856);
and U22127 (N_22127,N_21609,N_21225);
nor U22128 (N_22128,N_21216,N_21875);
and U22129 (N_22129,N_21305,N_21136);
or U22130 (N_22130,N_21638,N_21329);
or U22131 (N_22131,N_21468,N_21892);
or U22132 (N_22132,N_21783,N_21867);
or U22133 (N_22133,N_21794,N_21307);
and U22134 (N_22134,N_21598,N_21617);
and U22135 (N_22135,N_21580,N_21471);
or U22136 (N_22136,N_21301,N_21182);
nor U22137 (N_22137,N_21015,N_21325);
nand U22138 (N_22138,N_21156,N_21222);
nand U22139 (N_22139,N_21054,N_21122);
xor U22140 (N_22140,N_21842,N_21860);
nand U22141 (N_22141,N_21984,N_21135);
xnor U22142 (N_22142,N_21193,N_21955);
nor U22143 (N_22143,N_21207,N_21030);
nor U22144 (N_22144,N_21168,N_21038);
xor U22145 (N_22145,N_21174,N_21090);
and U22146 (N_22146,N_21914,N_21988);
nand U22147 (N_22147,N_21061,N_21583);
or U22148 (N_22148,N_21791,N_21278);
nor U22149 (N_22149,N_21808,N_21371);
or U22150 (N_22150,N_21417,N_21447);
nor U22151 (N_22151,N_21435,N_21440);
nor U22152 (N_22152,N_21009,N_21924);
or U22153 (N_22153,N_21388,N_21697);
nor U22154 (N_22154,N_21685,N_21478);
nor U22155 (N_22155,N_21020,N_21261);
nand U22156 (N_22156,N_21190,N_21537);
nor U22157 (N_22157,N_21629,N_21501);
and U22158 (N_22158,N_21169,N_21933);
or U22159 (N_22159,N_21968,N_21032);
nand U22160 (N_22160,N_21006,N_21585);
or U22161 (N_22161,N_21336,N_21188);
nand U22162 (N_22162,N_21071,N_21981);
xor U22163 (N_22163,N_21705,N_21486);
nand U22164 (N_22164,N_21903,N_21349);
xnor U22165 (N_22165,N_21526,N_21260);
nor U22166 (N_22166,N_21962,N_21036);
and U22167 (N_22167,N_21274,N_21891);
nand U22168 (N_22168,N_21669,N_21144);
nand U22169 (N_22169,N_21198,N_21567);
and U22170 (N_22170,N_21923,N_21391);
nand U22171 (N_22171,N_21459,N_21619);
nand U22172 (N_22172,N_21488,N_21209);
and U22173 (N_22173,N_21591,N_21840);
xor U22174 (N_22174,N_21102,N_21096);
xnor U22175 (N_22175,N_21535,N_21490);
or U22176 (N_22176,N_21103,N_21091);
and U22177 (N_22177,N_21841,N_21376);
xnor U22178 (N_22178,N_21473,N_21204);
nand U22179 (N_22179,N_21058,N_21608);
nand U22180 (N_22180,N_21869,N_21790);
or U22181 (N_22181,N_21622,N_21639);
nor U22182 (N_22182,N_21239,N_21152);
xor U22183 (N_22183,N_21675,N_21547);
or U22184 (N_22184,N_21876,N_21327);
xnor U22185 (N_22185,N_21835,N_21744);
or U22186 (N_22186,N_21453,N_21531);
nand U22187 (N_22187,N_21315,N_21277);
or U22188 (N_22188,N_21282,N_21125);
xnor U22189 (N_22189,N_21148,N_21199);
nand U22190 (N_22190,N_21017,N_21293);
nand U22191 (N_22191,N_21727,N_21802);
nand U22192 (N_22192,N_21568,N_21186);
xor U22193 (N_22193,N_21076,N_21119);
nor U22194 (N_22194,N_21118,N_21078);
xnor U22195 (N_22195,N_21626,N_21995);
and U22196 (N_22196,N_21026,N_21729);
and U22197 (N_22197,N_21281,N_21831);
and U22198 (N_22198,N_21953,N_21263);
nor U22199 (N_22199,N_21704,N_21960);
nor U22200 (N_22200,N_21303,N_21437);
or U22201 (N_22201,N_21411,N_21954);
nand U22202 (N_22202,N_21885,N_21458);
or U22203 (N_22203,N_21312,N_21807);
and U22204 (N_22204,N_21540,N_21539);
or U22205 (N_22205,N_21771,N_21730);
or U22206 (N_22206,N_21921,N_21331);
and U22207 (N_22207,N_21558,N_21848);
or U22208 (N_22208,N_21997,N_21191);
nor U22209 (N_22209,N_21879,N_21266);
xor U22210 (N_22210,N_21077,N_21504);
or U22211 (N_22211,N_21993,N_21819);
nor U22212 (N_22212,N_21880,N_21627);
nand U22213 (N_22213,N_21273,N_21323);
or U22214 (N_22214,N_21652,N_21151);
nor U22215 (N_22215,N_21507,N_21686);
nor U22216 (N_22216,N_21469,N_21477);
and U22217 (N_22217,N_21089,N_21073);
nand U22218 (N_22218,N_21706,N_21657);
and U22219 (N_22219,N_21005,N_21827);
nand U22220 (N_22220,N_21514,N_21801);
or U22221 (N_22221,N_21202,N_21481);
nand U22222 (N_22222,N_21037,N_21940);
nand U22223 (N_22223,N_21862,N_21906);
and U22224 (N_22224,N_21236,N_21001);
xnor U22225 (N_22225,N_21059,N_21575);
and U22226 (N_22226,N_21010,N_21171);
nor U22227 (N_22227,N_21375,N_21642);
nor U22228 (N_22228,N_21304,N_21162);
nor U22229 (N_22229,N_21176,N_21874);
xor U22230 (N_22230,N_21289,N_21117);
nor U22231 (N_22231,N_21648,N_21533);
nand U22232 (N_22232,N_21498,N_21902);
or U22233 (N_22233,N_21755,N_21389);
or U22234 (N_22234,N_21825,N_21141);
or U22235 (N_22235,N_21918,N_21314);
and U22236 (N_22236,N_21881,N_21400);
or U22237 (N_22237,N_21099,N_21971);
nor U22238 (N_22238,N_21181,N_21749);
and U22239 (N_22239,N_21383,N_21213);
and U22240 (N_22240,N_21401,N_21452);
nor U22241 (N_22241,N_21894,N_21661);
nor U22242 (N_22242,N_21034,N_21623);
xnor U22243 (N_22243,N_21255,N_21097);
or U22244 (N_22244,N_21708,N_21227);
or U22245 (N_22245,N_21434,N_21436);
or U22246 (N_22246,N_21287,N_21649);
or U22247 (N_22247,N_21133,N_21240);
nand U22248 (N_22248,N_21929,N_21769);
nand U22249 (N_22249,N_21254,N_21157);
nor U22250 (N_22250,N_21633,N_21928);
or U22251 (N_22251,N_21279,N_21494);
or U22252 (N_22252,N_21087,N_21521);
nand U22253 (N_22253,N_21586,N_21986);
and U22254 (N_22254,N_21429,N_21822);
nand U22255 (N_22255,N_21828,N_21713);
nand U22256 (N_22256,N_21710,N_21907);
or U22257 (N_22257,N_21092,N_21288);
nor U22258 (N_22258,N_21394,N_21788);
nor U22259 (N_22259,N_21560,N_21335);
nand U22260 (N_22260,N_21956,N_21998);
nand U22261 (N_22261,N_21114,N_21736);
xnor U22262 (N_22262,N_21847,N_21041);
nor U22263 (N_22263,N_21950,N_21100);
xor U22264 (N_22264,N_21513,N_21002);
and U22265 (N_22265,N_21341,N_21397);
or U22266 (N_22266,N_21121,N_21267);
and U22267 (N_22267,N_21621,N_21264);
nor U22268 (N_22268,N_21173,N_21313);
xnor U22269 (N_22269,N_21140,N_21419);
nand U22270 (N_22270,N_21441,N_21563);
and U22271 (N_22271,N_21055,N_21764);
xor U22272 (N_22272,N_21718,N_21393);
nor U22273 (N_22273,N_21541,N_21958);
xor U22274 (N_22274,N_21589,N_21022);
or U22275 (N_22275,N_21185,N_21479);
nor U22276 (N_22276,N_21219,N_21572);
or U22277 (N_22277,N_21605,N_21983);
nor U22278 (N_22278,N_21356,N_21593);
or U22279 (N_22279,N_21163,N_21813);
nand U22280 (N_22280,N_21590,N_21987);
or U22281 (N_22281,N_21630,N_21088);
xor U22282 (N_22282,N_21210,N_21673);
nand U22283 (N_22283,N_21850,N_21384);
nor U22284 (N_22284,N_21606,N_21243);
xnor U22285 (N_22285,N_21720,N_21310);
nand U22286 (N_22286,N_21534,N_21711);
nand U22287 (N_22287,N_21214,N_21821);
and U22288 (N_22288,N_21374,N_21868);
nor U22289 (N_22289,N_21691,N_21187);
or U22290 (N_22290,N_21155,N_21294);
nor U22291 (N_22291,N_21858,N_21670);
xnor U22292 (N_22292,N_21386,N_21382);
nand U22293 (N_22293,N_21654,N_21607);
or U22294 (N_22294,N_21270,N_21564);
and U22295 (N_22295,N_21782,N_21322);
xor U22296 (N_22296,N_21405,N_21484);
xor U22297 (N_22297,N_21739,N_21717);
xnor U22298 (N_22298,N_21834,N_21316);
and U22299 (N_22299,N_21610,N_21990);
nor U22300 (N_22300,N_21079,N_21889);
or U22301 (N_22301,N_21021,N_21820);
or U22302 (N_22302,N_21070,N_21684);
or U22303 (N_22303,N_21457,N_21805);
and U22304 (N_22304,N_21104,N_21925);
and U22305 (N_22305,N_21407,N_21992);
or U22306 (N_22306,N_21696,N_21311);
and U22307 (N_22307,N_21573,N_21975);
and U22308 (N_22308,N_21083,N_21687);
or U22309 (N_22309,N_21853,N_21035);
and U22310 (N_22310,N_21723,N_21896);
or U22311 (N_22311,N_21482,N_21057);
xor U22312 (N_22312,N_21569,N_21337);
or U22313 (N_22313,N_21766,N_21616);
nand U22314 (N_22314,N_21403,N_21226);
nor U22315 (N_22315,N_21887,N_21252);
and U22316 (N_22316,N_21839,N_21056);
nand U22317 (N_22317,N_21082,N_21503);
and U22318 (N_22318,N_21814,N_21786);
xnor U22319 (N_22319,N_21033,N_21497);
or U22320 (N_22320,N_21832,N_21577);
nand U22321 (N_22321,N_21945,N_21985);
nand U22322 (N_22322,N_21410,N_21013);
or U22323 (N_22323,N_21980,N_21909);
and U22324 (N_22324,N_21712,N_21245);
or U22325 (N_22325,N_21912,N_21012);
or U22326 (N_22326,N_21523,N_21520);
nand U22327 (N_22327,N_21636,N_21228);
nor U22328 (N_22328,N_21977,N_21116);
or U22329 (N_22329,N_21139,N_21192);
or U22330 (N_22330,N_21966,N_21265);
or U22331 (N_22331,N_21027,N_21051);
or U22332 (N_22332,N_21409,N_21742);
xnor U22333 (N_22333,N_21913,N_21908);
nor U22334 (N_22334,N_21917,N_21348);
or U22335 (N_22335,N_21942,N_21934);
and U22336 (N_22336,N_21948,N_21512);
nand U22337 (N_22337,N_21224,N_21679);
and U22338 (N_22338,N_21175,N_21200);
and U22339 (N_22339,N_21768,N_21664);
xnor U22340 (N_22340,N_21167,N_21120);
nor U22341 (N_22341,N_21291,N_21250);
nor U22342 (N_22342,N_21221,N_21852);
nor U22343 (N_22343,N_21525,N_21007);
or U22344 (N_22344,N_21588,N_21276);
or U22345 (N_22345,N_21733,N_21464);
nor U22346 (N_22346,N_21319,N_21164);
or U22347 (N_22347,N_21601,N_21746);
xor U22348 (N_22348,N_21461,N_21105);
or U22349 (N_22349,N_21599,N_21170);
and U22350 (N_22350,N_21800,N_21653);
nor U22351 (N_22351,N_21780,N_21677);
and U22352 (N_22352,N_21785,N_21778);
and U22353 (N_22353,N_21596,N_21565);
nor U22354 (N_22354,N_21624,N_21446);
or U22355 (N_22355,N_21861,N_21124);
and U22356 (N_22356,N_21680,N_21866);
and U22357 (N_22357,N_21046,N_21815);
xor U22358 (N_22358,N_21538,N_21387);
and U22359 (N_22359,N_21023,N_21877);
nor U22360 (N_22360,N_21138,N_21947);
nand U22361 (N_22361,N_21864,N_21905);
nor U22362 (N_22362,N_21901,N_21965);
and U22363 (N_22363,N_21893,N_21449);
nor U22364 (N_22364,N_21470,N_21234);
or U22365 (N_22365,N_21129,N_21066);
nor U22366 (N_22366,N_21342,N_21177);
or U22367 (N_22367,N_21430,N_21989);
xor U22368 (N_22368,N_21475,N_21422);
xor U22369 (N_22369,N_21796,N_21364);
nor U22370 (N_22370,N_21668,N_21247);
xor U22371 (N_22371,N_21959,N_21189);
nor U22372 (N_22372,N_21424,N_21799);
xor U22373 (N_22373,N_21689,N_21927);
and U22374 (N_22374,N_21758,N_21765);
nand U22375 (N_22375,N_21235,N_21824);
nor U22376 (N_22376,N_21833,N_21702);
nand U22377 (N_22377,N_21641,N_21480);
nor U22378 (N_22378,N_21396,N_21613);
nand U22379 (N_22379,N_21719,N_21734);
xnor U22380 (N_22380,N_21443,N_21491);
or U22381 (N_22381,N_21000,N_21165);
nor U22382 (N_22382,N_21220,N_21793);
and U22383 (N_22383,N_21134,N_21737);
and U22384 (N_22384,N_21579,N_21149);
nor U22385 (N_22385,N_21496,N_21571);
or U22386 (N_22386,N_21398,N_21982);
or U22387 (N_22387,N_21890,N_21628);
xnor U22388 (N_22388,N_21280,N_21425);
nor U22389 (N_22389,N_21380,N_21732);
xor U22390 (N_22390,N_21248,N_21615);
or U22391 (N_22391,N_21067,N_21604);
nor U22392 (N_22392,N_21295,N_21455);
nor U22393 (N_22393,N_21774,N_21262);
xnor U22394 (N_22394,N_21444,N_21944);
xor U22395 (N_22395,N_21334,N_21145);
and U22396 (N_22396,N_21855,N_21970);
nand U22397 (N_22397,N_21754,N_21603);
nor U22398 (N_22398,N_21926,N_21871);
or U22399 (N_22399,N_21098,N_21259);
nand U22400 (N_22400,N_21522,N_21996);
nand U22401 (N_22401,N_21826,N_21142);
nor U22402 (N_22402,N_21130,N_21166);
and U22403 (N_22403,N_21492,N_21378);
or U22404 (N_22404,N_21823,N_21865);
xor U22405 (N_22405,N_21527,N_21351);
or U22406 (N_22406,N_21667,N_21974);
or U22407 (N_22407,N_21857,N_21367);
or U22408 (N_22408,N_21555,N_21645);
and U22409 (N_22409,N_21594,N_21557);
nor U22410 (N_22410,N_21217,N_21516);
nand U22411 (N_22411,N_21326,N_21904);
and U22412 (N_22412,N_21195,N_21499);
nor U22413 (N_22413,N_21602,N_21682);
nand U22414 (N_22414,N_21131,N_21545);
xor U22415 (N_22415,N_21343,N_21767);
and U22416 (N_22416,N_21237,N_21703);
nor U22417 (N_22417,N_21357,N_21137);
or U22418 (N_22418,N_21086,N_21549);
nor U22419 (N_22419,N_21018,N_21332);
and U22420 (N_22420,N_21693,N_21506);
and U22421 (N_22421,N_21275,N_21111);
and U22422 (N_22422,N_21040,N_21707);
and U22423 (N_22423,N_21961,N_21884);
nor U22424 (N_22424,N_21735,N_21445);
nor U22425 (N_22425,N_21863,N_21333);
nand U22426 (N_22426,N_21741,N_21939);
xnor U22427 (N_22427,N_21510,N_21467);
nand U22428 (N_22428,N_21886,N_21146);
xor U22429 (N_22429,N_21792,N_21536);
nor U22430 (N_22430,N_21969,N_21753);
nor U22431 (N_22431,N_21637,N_21935);
nor U22432 (N_22432,N_21223,N_21084);
xnor U22433 (N_22433,N_21634,N_21836);
nor U22434 (N_22434,N_21612,N_21803);
or U22435 (N_22435,N_21751,N_21308);
xnor U22436 (N_22436,N_21957,N_21360);
nor U22437 (N_22437,N_21253,N_21062);
xnor U22438 (N_22438,N_21439,N_21206);
or U22439 (N_22439,N_21951,N_21900);
nor U22440 (N_22440,N_21361,N_21203);
nor U22441 (N_22441,N_21218,N_21665);
and U22442 (N_22442,N_21916,N_21251);
xor U22443 (N_22443,N_21432,N_21011);
and U22444 (N_22444,N_21460,N_21433);
or U22445 (N_22445,N_21395,N_21529);
nor U22446 (N_22446,N_21650,N_21660);
xor U22447 (N_22447,N_21678,N_21229);
or U22448 (N_22448,N_21063,N_21804);
nor U22449 (N_22449,N_21787,N_21967);
nor U22450 (N_22450,N_21899,N_21775);
nor U22451 (N_22451,N_21463,N_21286);
nand U22452 (N_22452,N_21355,N_21283);
nor U22453 (N_22453,N_21212,N_21414);
or U22454 (N_22454,N_21747,N_21830);
xnor U22455 (N_22455,N_21870,N_21197);
xnor U22456 (N_22456,N_21194,N_21878);
nor U22457 (N_22457,N_21919,N_21028);
xnor U22458 (N_22458,N_21052,N_21024);
and U22459 (N_22459,N_21413,N_21306);
nand U22460 (N_22460,N_21042,N_21882);
or U22461 (N_22461,N_21328,N_21752);
and U22462 (N_22462,N_21632,N_21994);
nand U22463 (N_22463,N_21465,N_21290);
or U22464 (N_22464,N_21369,N_21911);
nor U22465 (N_22465,N_21039,N_21019);
xor U22466 (N_22466,N_21544,N_21421);
nor U22467 (N_22467,N_21750,N_21519);
or U22468 (N_22468,N_21715,N_21184);
and U22469 (N_22469,N_21562,N_21795);
nand U22470 (N_22470,N_21159,N_21592);
xor U22471 (N_22471,N_21454,N_21699);
nor U22472 (N_22472,N_21095,N_21143);
nor U22473 (N_22473,N_21745,N_21370);
nor U22474 (N_22474,N_21485,N_21528);
nand U22475 (N_22475,N_21915,N_21837);
nand U22476 (N_22476,N_21566,N_21532);
xnor U22477 (N_22477,N_21647,N_21074);
nor U22478 (N_22478,N_21049,N_21172);
and U22479 (N_22479,N_21721,N_21431);
or U22480 (N_22480,N_21659,N_21509);
nand U22481 (N_22481,N_21505,N_21843);
and U22482 (N_22482,N_21487,N_21756);
xor U22483 (N_22483,N_21402,N_21897);
or U22484 (N_22484,N_21584,N_21618);
or U22485 (N_22485,N_21524,N_21047);
or U22486 (N_22486,N_21072,N_21085);
or U22487 (N_22487,N_21517,N_21365);
nor U22488 (N_22488,N_21600,N_21518);
nor U22489 (N_22489,N_21242,N_21094);
nor U22490 (N_22490,N_21014,N_21183);
and U22491 (N_22491,N_21309,N_21581);
nand U22492 (N_22492,N_21297,N_21551);
or U22493 (N_22493,N_21426,N_21153);
or U22494 (N_22494,N_21271,N_21065);
or U22495 (N_22495,N_21931,N_21676);
nand U22496 (N_22496,N_21559,N_21101);
nor U22497 (N_22497,N_21500,N_21770);
and U22498 (N_22498,N_21462,N_21399);
nor U22499 (N_22499,N_21373,N_21080);
and U22500 (N_22500,N_21361,N_21130);
xnor U22501 (N_22501,N_21828,N_21475);
xnor U22502 (N_22502,N_21342,N_21960);
nand U22503 (N_22503,N_21092,N_21712);
or U22504 (N_22504,N_21664,N_21472);
xor U22505 (N_22505,N_21880,N_21228);
xor U22506 (N_22506,N_21685,N_21290);
nand U22507 (N_22507,N_21387,N_21080);
nand U22508 (N_22508,N_21910,N_21942);
xor U22509 (N_22509,N_21374,N_21580);
xnor U22510 (N_22510,N_21050,N_21841);
xnor U22511 (N_22511,N_21282,N_21695);
nand U22512 (N_22512,N_21112,N_21633);
and U22513 (N_22513,N_21631,N_21174);
and U22514 (N_22514,N_21014,N_21919);
nor U22515 (N_22515,N_21038,N_21539);
and U22516 (N_22516,N_21529,N_21849);
xor U22517 (N_22517,N_21988,N_21465);
xnor U22518 (N_22518,N_21504,N_21303);
nor U22519 (N_22519,N_21065,N_21711);
nor U22520 (N_22520,N_21871,N_21855);
nand U22521 (N_22521,N_21189,N_21777);
nand U22522 (N_22522,N_21604,N_21193);
nor U22523 (N_22523,N_21800,N_21400);
or U22524 (N_22524,N_21494,N_21342);
nor U22525 (N_22525,N_21177,N_21769);
nor U22526 (N_22526,N_21802,N_21632);
xor U22527 (N_22527,N_21733,N_21340);
xor U22528 (N_22528,N_21204,N_21620);
nand U22529 (N_22529,N_21629,N_21985);
nor U22530 (N_22530,N_21184,N_21013);
and U22531 (N_22531,N_21289,N_21338);
or U22532 (N_22532,N_21041,N_21868);
nand U22533 (N_22533,N_21763,N_21807);
and U22534 (N_22534,N_21695,N_21504);
nand U22535 (N_22535,N_21136,N_21359);
nor U22536 (N_22536,N_21427,N_21651);
or U22537 (N_22537,N_21211,N_21274);
nor U22538 (N_22538,N_21937,N_21044);
or U22539 (N_22539,N_21842,N_21988);
and U22540 (N_22540,N_21068,N_21691);
nand U22541 (N_22541,N_21051,N_21769);
and U22542 (N_22542,N_21411,N_21273);
xnor U22543 (N_22543,N_21186,N_21173);
xor U22544 (N_22544,N_21732,N_21185);
nor U22545 (N_22545,N_21725,N_21313);
nor U22546 (N_22546,N_21834,N_21685);
or U22547 (N_22547,N_21235,N_21725);
nand U22548 (N_22548,N_21543,N_21861);
and U22549 (N_22549,N_21001,N_21098);
and U22550 (N_22550,N_21264,N_21295);
and U22551 (N_22551,N_21402,N_21566);
and U22552 (N_22552,N_21696,N_21423);
nand U22553 (N_22553,N_21533,N_21673);
nor U22554 (N_22554,N_21101,N_21779);
xor U22555 (N_22555,N_21323,N_21887);
nor U22556 (N_22556,N_21489,N_21128);
nand U22557 (N_22557,N_21307,N_21535);
nor U22558 (N_22558,N_21938,N_21842);
and U22559 (N_22559,N_21518,N_21074);
or U22560 (N_22560,N_21869,N_21099);
nor U22561 (N_22561,N_21504,N_21213);
nand U22562 (N_22562,N_21034,N_21795);
nand U22563 (N_22563,N_21671,N_21554);
and U22564 (N_22564,N_21862,N_21602);
nand U22565 (N_22565,N_21060,N_21713);
or U22566 (N_22566,N_21954,N_21027);
or U22567 (N_22567,N_21717,N_21915);
or U22568 (N_22568,N_21592,N_21662);
nand U22569 (N_22569,N_21719,N_21685);
or U22570 (N_22570,N_21595,N_21492);
nand U22571 (N_22571,N_21722,N_21301);
nand U22572 (N_22572,N_21962,N_21281);
or U22573 (N_22573,N_21784,N_21697);
nor U22574 (N_22574,N_21653,N_21968);
and U22575 (N_22575,N_21612,N_21319);
and U22576 (N_22576,N_21330,N_21361);
xnor U22577 (N_22577,N_21404,N_21150);
nand U22578 (N_22578,N_21600,N_21150);
nand U22579 (N_22579,N_21262,N_21216);
nor U22580 (N_22580,N_21992,N_21408);
nand U22581 (N_22581,N_21676,N_21659);
nor U22582 (N_22582,N_21838,N_21473);
or U22583 (N_22583,N_21638,N_21021);
xnor U22584 (N_22584,N_21359,N_21922);
xor U22585 (N_22585,N_21989,N_21804);
nand U22586 (N_22586,N_21559,N_21995);
or U22587 (N_22587,N_21542,N_21409);
nand U22588 (N_22588,N_21649,N_21620);
or U22589 (N_22589,N_21569,N_21235);
or U22590 (N_22590,N_21632,N_21571);
nor U22591 (N_22591,N_21155,N_21045);
nand U22592 (N_22592,N_21392,N_21905);
and U22593 (N_22593,N_21997,N_21180);
xor U22594 (N_22594,N_21202,N_21156);
or U22595 (N_22595,N_21660,N_21119);
or U22596 (N_22596,N_21269,N_21143);
or U22597 (N_22597,N_21889,N_21189);
nor U22598 (N_22598,N_21460,N_21970);
or U22599 (N_22599,N_21234,N_21318);
nand U22600 (N_22600,N_21304,N_21327);
xor U22601 (N_22601,N_21270,N_21391);
and U22602 (N_22602,N_21459,N_21610);
or U22603 (N_22603,N_21845,N_21707);
or U22604 (N_22604,N_21626,N_21001);
and U22605 (N_22605,N_21925,N_21340);
or U22606 (N_22606,N_21172,N_21849);
nor U22607 (N_22607,N_21399,N_21116);
nand U22608 (N_22608,N_21883,N_21258);
nand U22609 (N_22609,N_21984,N_21569);
and U22610 (N_22610,N_21433,N_21104);
xor U22611 (N_22611,N_21697,N_21186);
or U22612 (N_22612,N_21096,N_21644);
or U22613 (N_22613,N_21153,N_21030);
or U22614 (N_22614,N_21325,N_21757);
or U22615 (N_22615,N_21991,N_21935);
nand U22616 (N_22616,N_21971,N_21675);
xor U22617 (N_22617,N_21889,N_21405);
nand U22618 (N_22618,N_21143,N_21593);
or U22619 (N_22619,N_21904,N_21266);
nor U22620 (N_22620,N_21939,N_21792);
and U22621 (N_22621,N_21254,N_21219);
or U22622 (N_22622,N_21064,N_21494);
xor U22623 (N_22623,N_21242,N_21895);
nor U22624 (N_22624,N_21379,N_21707);
and U22625 (N_22625,N_21523,N_21171);
xnor U22626 (N_22626,N_21923,N_21392);
or U22627 (N_22627,N_21300,N_21335);
or U22628 (N_22628,N_21316,N_21102);
nand U22629 (N_22629,N_21338,N_21748);
nor U22630 (N_22630,N_21867,N_21659);
nand U22631 (N_22631,N_21842,N_21607);
xor U22632 (N_22632,N_21461,N_21198);
xor U22633 (N_22633,N_21061,N_21389);
nor U22634 (N_22634,N_21703,N_21680);
xnor U22635 (N_22635,N_21869,N_21494);
nand U22636 (N_22636,N_21792,N_21039);
or U22637 (N_22637,N_21512,N_21724);
or U22638 (N_22638,N_21456,N_21336);
xnor U22639 (N_22639,N_21480,N_21611);
xor U22640 (N_22640,N_21343,N_21314);
nand U22641 (N_22641,N_21568,N_21087);
or U22642 (N_22642,N_21477,N_21875);
and U22643 (N_22643,N_21211,N_21043);
xnor U22644 (N_22644,N_21454,N_21089);
or U22645 (N_22645,N_21958,N_21948);
xor U22646 (N_22646,N_21624,N_21973);
and U22647 (N_22647,N_21460,N_21391);
or U22648 (N_22648,N_21348,N_21339);
xnor U22649 (N_22649,N_21680,N_21779);
or U22650 (N_22650,N_21624,N_21462);
nor U22651 (N_22651,N_21192,N_21102);
and U22652 (N_22652,N_21580,N_21166);
and U22653 (N_22653,N_21222,N_21311);
xor U22654 (N_22654,N_21623,N_21545);
and U22655 (N_22655,N_21237,N_21611);
or U22656 (N_22656,N_21636,N_21748);
or U22657 (N_22657,N_21895,N_21875);
nor U22658 (N_22658,N_21992,N_21593);
or U22659 (N_22659,N_21863,N_21400);
nand U22660 (N_22660,N_21213,N_21996);
or U22661 (N_22661,N_21096,N_21145);
xor U22662 (N_22662,N_21257,N_21874);
and U22663 (N_22663,N_21357,N_21280);
or U22664 (N_22664,N_21540,N_21914);
or U22665 (N_22665,N_21804,N_21641);
nor U22666 (N_22666,N_21666,N_21694);
and U22667 (N_22667,N_21534,N_21855);
xor U22668 (N_22668,N_21100,N_21459);
and U22669 (N_22669,N_21242,N_21536);
nand U22670 (N_22670,N_21049,N_21991);
or U22671 (N_22671,N_21228,N_21954);
or U22672 (N_22672,N_21902,N_21866);
and U22673 (N_22673,N_21486,N_21801);
nor U22674 (N_22674,N_21173,N_21629);
nor U22675 (N_22675,N_21848,N_21426);
nor U22676 (N_22676,N_21142,N_21225);
nor U22677 (N_22677,N_21384,N_21119);
nand U22678 (N_22678,N_21708,N_21765);
nand U22679 (N_22679,N_21825,N_21305);
nand U22680 (N_22680,N_21914,N_21548);
xor U22681 (N_22681,N_21554,N_21829);
or U22682 (N_22682,N_21271,N_21078);
and U22683 (N_22683,N_21993,N_21558);
nor U22684 (N_22684,N_21528,N_21486);
xnor U22685 (N_22685,N_21118,N_21050);
nor U22686 (N_22686,N_21145,N_21163);
and U22687 (N_22687,N_21591,N_21386);
and U22688 (N_22688,N_21134,N_21252);
nand U22689 (N_22689,N_21719,N_21736);
or U22690 (N_22690,N_21817,N_21407);
nand U22691 (N_22691,N_21769,N_21747);
nor U22692 (N_22692,N_21786,N_21104);
and U22693 (N_22693,N_21547,N_21683);
nor U22694 (N_22694,N_21169,N_21926);
nand U22695 (N_22695,N_21571,N_21901);
xnor U22696 (N_22696,N_21164,N_21038);
or U22697 (N_22697,N_21419,N_21884);
nand U22698 (N_22698,N_21649,N_21480);
nor U22699 (N_22699,N_21017,N_21933);
xnor U22700 (N_22700,N_21045,N_21739);
or U22701 (N_22701,N_21930,N_21712);
xnor U22702 (N_22702,N_21807,N_21682);
nand U22703 (N_22703,N_21543,N_21044);
or U22704 (N_22704,N_21637,N_21366);
and U22705 (N_22705,N_21385,N_21510);
xor U22706 (N_22706,N_21340,N_21508);
nand U22707 (N_22707,N_21320,N_21234);
nand U22708 (N_22708,N_21241,N_21761);
or U22709 (N_22709,N_21193,N_21300);
and U22710 (N_22710,N_21339,N_21788);
nand U22711 (N_22711,N_21604,N_21553);
and U22712 (N_22712,N_21823,N_21190);
nand U22713 (N_22713,N_21201,N_21093);
and U22714 (N_22714,N_21049,N_21744);
nand U22715 (N_22715,N_21480,N_21708);
nor U22716 (N_22716,N_21335,N_21575);
nand U22717 (N_22717,N_21918,N_21406);
nor U22718 (N_22718,N_21546,N_21904);
nor U22719 (N_22719,N_21836,N_21262);
nand U22720 (N_22720,N_21040,N_21259);
xor U22721 (N_22721,N_21090,N_21558);
and U22722 (N_22722,N_21588,N_21714);
and U22723 (N_22723,N_21114,N_21872);
xor U22724 (N_22724,N_21329,N_21478);
xnor U22725 (N_22725,N_21384,N_21527);
nand U22726 (N_22726,N_21999,N_21500);
nor U22727 (N_22727,N_21221,N_21802);
nor U22728 (N_22728,N_21358,N_21729);
xnor U22729 (N_22729,N_21752,N_21576);
or U22730 (N_22730,N_21925,N_21692);
or U22731 (N_22731,N_21768,N_21268);
and U22732 (N_22732,N_21265,N_21489);
or U22733 (N_22733,N_21380,N_21237);
nand U22734 (N_22734,N_21250,N_21221);
nand U22735 (N_22735,N_21298,N_21048);
nor U22736 (N_22736,N_21056,N_21588);
nor U22737 (N_22737,N_21477,N_21395);
nor U22738 (N_22738,N_21684,N_21763);
or U22739 (N_22739,N_21626,N_21753);
xor U22740 (N_22740,N_21951,N_21850);
nor U22741 (N_22741,N_21902,N_21820);
nor U22742 (N_22742,N_21939,N_21173);
or U22743 (N_22743,N_21618,N_21736);
nor U22744 (N_22744,N_21515,N_21744);
nor U22745 (N_22745,N_21030,N_21681);
xnor U22746 (N_22746,N_21810,N_21199);
xnor U22747 (N_22747,N_21465,N_21959);
nor U22748 (N_22748,N_21133,N_21334);
nor U22749 (N_22749,N_21486,N_21011);
or U22750 (N_22750,N_21830,N_21609);
xnor U22751 (N_22751,N_21999,N_21863);
or U22752 (N_22752,N_21560,N_21710);
or U22753 (N_22753,N_21922,N_21565);
and U22754 (N_22754,N_21363,N_21516);
and U22755 (N_22755,N_21745,N_21754);
xnor U22756 (N_22756,N_21578,N_21167);
or U22757 (N_22757,N_21415,N_21995);
xor U22758 (N_22758,N_21851,N_21628);
nor U22759 (N_22759,N_21732,N_21650);
and U22760 (N_22760,N_21688,N_21080);
nor U22761 (N_22761,N_21709,N_21364);
xnor U22762 (N_22762,N_21700,N_21203);
nand U22763 (N_22763,N_21697,N_21456);
and U22764 (N_22764,N_21609,N_21059);
and U22765 (N_22765,N_21646,N_21883);
nand U22766 (N_22766,N_21147,N_21891);
or U22767 (N_22767,N_21636,N_21981);
nor U22768 (N_22768,N_21429,N_21684);
xor U22769 (N_22769,N_21134,N_21705);
or U22770 (N_22770,N_21629,N_21735);
nor U22771 (N_22771,N_21670,N_21969);
nand U22772 (N_22772,N_21426,N_21534);
nor U22773 (N_22773,N_21211,N_21570);
nor U22774 (N_22774,N_21374,N_21217);
nand U22775 (N_22775,N_21801,N_21331);
and U22776 (N_22776,N_21829,N_21761);
nor U22777 (N_22777,N_21679,N_21947);
nor U22778 (N_22778,N_21331,N_21884);
nor U22779 (N_22779,N_21897,N_21115);
nor U22780 (N_22780,N_21211,N_21565);
nor U22781 (N_22781,N_21037,N_21382);
and U22782 (N_22782,N_21651,N_21737);
nor U22783 (N_22783,N_21363,N_21619);
xnor U22784 (N_22784,N_21782,N_21546);
xnor U22785 (N_22785,N_21056,N_21806);
or U22786 (N_22786,N_21027,N_21439);
or U22787 (N_22787,N_21520,N_21018);
and U22788 (N_22788,N_21437,N_21997);
xor U22789 (N_22789,N_21639,N_21584);
xor U22790 (N_22790,N_21343,N_21282);
nor U22791 (N_22791,N_21359,N_21076);
xnor U22792 (N_22792,N_21781,N_21592);
xnor U22793 (N_22793,N_21210,N_21871);
xnor U22794 (N_22794,N_21160,N_21108);
or U22795 (N_22795,N_21545,N_21584);
nand U22796 (N_22796,N_21652,N_21786);
and U22797 (N_22797,N_21780,N_21435);
nor U22798 (N_22798,N_21368,N_21944);
nor U22799 (N_22799,N_21106,N_21552);
xnor U22800 (N_22800,N_21956,N_21707);
and U22801 (N_22801,N_21088,N_21592);
nor U22802 (N_22802,N_21464,N_21682);
nor U22803 (N_22803,N_21319,N_21128);
xor U22804 (N_22804,N_21704,N_21025);
nor U22805 (N_22805,N_21098,N_21135);
nor U22806 (N_22806,N_21035,N_21733);
or U22807 (N_22807,N_21891,N_21756);
xnor U22808 (N_22808,N_21685,N_21560);
or U22809 (N_22809,N_21665,N_21650);
and U22810 (N_22810,N_21164,N_21072);
xor U22811 (N_22811,N_21294,N_21998);
or U22812 (N_22812,N_21623,N_21206);
or U22813 (N_22813,N_21236,N_21160);
nand U22814 (N_22814,N_21174,N_21817);
xor U22815 (N_22815,N_21091,N_21973);
nand U22816 (N_22816,N_21715,N_21000);
or U22817 (N_22817,N_21358,N_21857);
nand U22818 (N_22818,N_21075,N_21713);
and U22819 (N_22819,N_21679,N_21816);
xor U22820 (N_22820,N_21713,N_21134);
nand U22821 (N_22821,N_21102,N_21348);
or U22822 (N_22822,N_21084,N_21237);
and U22823 (N_22823,N_21302,N_21333);
or U22824 (N_22824,N_21501,N_21162);
nand U22825 (N_22825,N_21250,N_21485);
nor U22826 (N_22826,N_21223,N_21380);
and U22827 (N_22827,N_21826,N_21288);
and U22828 (N_22828,N_21178,N_21549);
nor U22829 (N_22829,N_21184,N_21566);
or U22830 (N_22830,N_21546,N_21409);
and U22831 (N_22831,N_21471,N_21131);
and U22832 (N_22832,N_21992,N_21781);
nand U22833 (N_22833,N_21599,N_21085);
or U22834 (N_22834,N_21289,N_21540);
xnor U22835 (N_22835,N_21937,N_21984);
nand U22836 (N_22836,N_21889,N_21627);
xnor U22837 (N_22837,N_21980,N_21461);
and U22838 (N_22838,N_21705,N_21816);
nand U22839 (N_22839,N_21927,N_21614);
nor U22840 (N_22840,N_21174,N_21689);
nand U22841 (N_22841,N_21082,N_21908);
or U22842 (N_22842,N_21909,N_21803);
nor U22843 (N_22843,N_21445,N_21216);
nand U22844 (N_22844,N_21570,N_21487);
or U22845 (N_22845,N_21776,N_21528);
or U22846 (N_22846,N_21915,N_21473);
xnor U22847 (N_22847,N_21100,N_21015);
and U22848 (N_22848,N_21572,N_21602);
and U22849 (N_22849,N_21305,N_21820);
or U22850 (N_22850,N_21710,N_21100);
xor U22851 (N_22851,N_21051,N_21750);
and U22852 (N_22852,N_21445,N_21141);
xor U22853 (N_22853,N_21716,N_21856);
nor U22854 (N_22854,N_21281,N_21459);
nand U22855 (N_22855,N_21102,N_21727);
nand U22856 (N_22856,N_21791,N_21554);
or U22857 (N_22857,N_21728,N_21068);
or U22858 (N_22858,N_21467,N_21213);
nand U22859 (N_22859,N_21975,N_21244);
nor U22860 (N_22860,N_21372,N_21955);
nand U22861 (N_22861,N_21997,N_21891);
nor U22862 (N_22862,N_21181,N_21214);
nor U22863 (N_22863,N_21438,N_21397);
nor U22864 (N_22864,N_21747,N_21374);
xor U22865 (N_22865,N_21991,N_21227);
nor U22866 (N_22866,N_21657,N_21601);
nor U22867 (N_22867,N_21933,N_21222);
xnor U22868 (N_22868,N_21514,N_21231);
and U22869 (N_22869,N_21312,N_21705);
or U22870 (N_22870,N_21157,N_21129);
nand U22871 (N_22871,N_21618,N_21935);
and U22872 (N_22872,N_21464,N_21546);
xnor U22873 (N_22873,N_21690,N_21654);
and U22874 (N_22874,N_21162,N_21724);
nor U22875 (N_22875,N_21958,N_21660);
nor U22876 (N_22876,N_21312,N_21441);
xor U22877 (N_22877,N_21663,N_21101);
xnor U22878 (N_22878,N_21457,N_21525);
nand U22879 (N_22879,N_21217,N_21958);
or U22880 (N_22880,N_21934,N_21174);
xnor U22881 (N_22881,N_21988,N_21027);
or U22882 (N_22882,N_21395,N_21095);
or U22883 (N_22883,N_21174,N_21865);
and U22884 (N_22884,N_21039,N_21157);
nor U22885 (N_22885,N_21131,N_21003);
and U22886 (N_22886,N_21211,N_21883);
nor U22887 (N_22887,N_21470,N_21871);
or U22888 (N_22888,N_21100,N_21609);
nor U22889 (N_22889,N_21529,N_21881);
nor U22890 (N_22890,N_21812,N_21876);
nor U22891 (N_22891,N_21621,N_21259);
and U22892 (N_22892,N_21781,N_21418);
nor U22893 (N_22893,N_21876,N_21324);
nand U22894 (N_22894,N_21117,N_21677);
xnor U22895 (N_22895,N_21217,N_21268);
nand U22896 (N_22896,N_21866,N_21808);
nor U22897 (N_22897,N_21755,N_21380);
or U22898 (N_22898,N_21660,N_21818);
xnor U22899 (N_22899,N_21271,N_21653);
nand U22900 (N_22900,N_21006,N_21625);
nand U22901 (N_22901,N_21814,N_21430);
and U22902 (N_22902,N_21964,N_21000);
and U22903 (N_22903,N_21519,N_21216);
or U22904 (N_22904,N_21604,N_21549);
nor U22905 (N_22905,N_21205,N_21957);
nor U22906 (N_22906,N_21302,N_21261);
nor U22907 (N_22907,N_21468,N_21990);
xor U22908 (N_22908,N_21405,N_21458);
and U22909 (N_22909,N_21751,N_21519);
and U22910 (N_22910,N_21808,N_21548);
nand U22911 (N_22911,N_21550,N_21102);
xor U22912 (N_22912,N_21853,N_21449);
or U22913 (N_22913,N_21961,N_21707);
xor U22914 (N_22914,N_21889,N_21863);
and U22915 (N_22915,N_21083,N_21015);
or U22916 (N_22916,N_21768,N_21749);
nand U22917 (N_22917,N_21162,N_21218);
nand U22918 (N_22918,N_21811,N_21300);
or U22919 (N_22919,N_21611,N_21575);
and U22920 (N_22920,N_21121,N_21511);
nand U22921 (N_22921,N_21642,N_21111);
nand U22922 (N_22922,N_21814,N_21914);
or U22923 (N_22923,N_21271,N_21534);
or U22924 (N_22924,N_21952,N_21393);
nor U22925 (N_22925,N_21993,N_21655);
nand U22926 (N_22926,N_21475,N_21356);
xor U22927 (N_22927,N_21900,N_21262);
nor U22928 (N_22928,N_21286,N_21379);
nand U22929 (N_22929,N_21537,N_21378);
nand U22930 (N_22930,N_21999,N_21403);
xnor U22931 (N_22931,N_21210,N_21330);
or U22932 (N_22932,N_21735,N_21767);
nor U22933 (N_22933,N_21908,N_21251);
nand U22934 (N_22934,N_21696,N_21085);
nand U22935 (N_22935,N_21169,N_21472);
and U22936 (N_22936,N_21087,N_21750);
or U22937 (N_22937,N_21535,N_21003);
nand U22938 (N_22938,N_21426,N_21420);
nand U22939 (N_22939,N_21630,N_21843);
and U22940 (N_22940,N_21345,N_21421);
nand U22941 (N_22941,N_21663,N_21120);
and U22942 (N_22942,N_21911,N_21671);
nor U22943 (N_22943,N_21632,N_21655);
nand U22944 (N_22944,N_21115,N_21559);
or U22945 (N_22945,N_21157,N_21835);
nor U22946 (N_22946,N_21961,N_21185);
or U22947 (N_22947,N_21074,N_21273);
and U22948 (N_22948,N_21874,N_21913);
nand U22949 (N_22949,N_21786,N_21060);
xor U22950 (N_22950,N_21953,N_21029);
and U22951 (N_22951,N_21912,N_21727);
xnor U22952 (N_22952,N_21284,N_21501);
or U22953 (N_22953,N_21251,N_21803);
nor U22954 (N_22954,N_21416,N_21401);
nor U22955 (N_22955,N_21468,N_21531);
nor U22956 (N_22956,N_21909,N_21982);
nor U22957 (N_22957,N_21504,N_21125);
nand U22958 (N_22958,N_21738,N_21413);
nor U22959 (N_22959,N_21319,N_21512);
or U22960 (N_22960,N_21001,N_21042);
nor U22961 (N_22961,N_21350,N_21273);
and U22962 (N_22962,N_21610,N_21880);
or U22963 (N_22963,N_21097,N_21446);
nand U22964 (N_22964,N_21259,N_21402);
xnor U22965 (N_22965,N_21828,N_21014);
xor U22966 (N_22966,N_21993,N_21246);
xor U22967 (N_22967,N_21111,N_21607);
xnor U22968 (N_22968,N_21658,N_21095);
or U22969 (N_22969,N_21552,N_21715);
xor U22970 (N_22970,N_21720,N_21789);
and U22971 (N_22971,N_21186,N_21625);
or U22972 (N_22972,N_21537,N_21545);
nor U22973 (N_22973,N_21684,N_21608);
and U22974 (N_22974,N_21821,N_21331);
nand U22975 (N_22975,N_21728,N_21072);
nand U22976 (N_22976,N_21150,N_21987);
nand U22977 (N_22977,N_21102,N_21655);
and U22978 (N_22978,N_21002,N_21639);
and U22979 (N_22979,N_21749,N_21366);
nand U22980 (N_22980,N_21777,N_21021);
nor U22981 (N_22981,N_21721,N_21534);
nand U22982 (N_22982,N_21173,N_21681);
and U22983 (N_22983,N_21834,N_21456);
nor U22984 (N_22984,N_21865,N_21616);
nand U22985 (N_22985,N_21127,N_21949);
nor U22986 (N_22986,N_21879,N_21388);
nor U22987 (N_22987,N_21158,N_21428);
nand U22988 (N_22988,N_21613,N_21261);
xnor U22989 (N_22989,N_21150,N_21800);
and U22990 (N_22990,N_21970,N_21314);
nand U22991 (N_22991,N_21270,N_21550);
nand U22992 (N_22992,N_21316,N_21621);
xor U22993 (N_22993,N_21149,N_21715);
xor U22994 (N_22994,N_21070,N_21407);
nor U22995 (N_22995,N_21949,N_21887);
nor U22996 (N_22996,N_21670,N_21198);
and U22997 (N_22997,N_21783,N_21870);
or U22998 (N_22998,N_21153,N_21330);
or U22999 (N_22999,N_21994,N_21241);
nand U23000 (N_23000,N_22659,N_22756);
and U23001 (N_23001,N_22210,N_22066);
or U23002 (N_23002,N_22579,N_22840);
xnor U23003 (N_23003,N_22107,N_22959);
and U23004 (N_23004,N_22972,N_22029);
or U23005 (N_23005,N_22228,N_22895);
xor U23006 (N_23006,N_22908,N_22333);
xnor U23007 (N_23007,N_22578,N_22682);
xor U23008 (N_23008,N_22047,N_22850);
or U23009 (N_23009,N_22156,N_22829);
nand U23010 (N_23010,N_22511,N_22008);
and U23011 (N_23011,N_22764,N_22742);
nor U23012 (N_23012,N_22015,N_22572);
and U23013 (N_23013,N_22658,N_22433);
xor U23014 (N_23014,N_22813,N_22241);
and U23015 (N_23015,N_22023,N_22062);
nand U23016 (N_23016,N_22105,N_22584);
xnor U23017 (N_23017,N_22527,N_22833);
nor U23018 (N_23018,N_22541,N_22346);
nor U23019 (N_23019,N_22197,N_22858);
and U23020 (N_23020,N_22627,N_22362);
or U23021 (N_23021,N_22053,N_22547);
xor U23022 (N_23022,N_22724,N_22688);
and U23023 (N_23023,N_22063,N_22891);
nor U23024 (N_23024,N_22815,N_22302);
nand U23025 (N_23025,N_22316,N_22038);
xor U23026 (N_23026,N_22291,N_22538);
xor U23027 (N_23027,N_22426,N_22336);
and U23028 (N_23028,N_22952,N_22759);
nor U23029 (N_23029,N_22088,N_22723);
and U23030 (N_23030,N_22184,N_22936);
and U23031 (N_23031,N_22423,N_22803);
nand U23032 (N_23032,N_22513,N_22109);
xor U23033 (N_23033,N_22490,N_22190);
and U23034 (N_23034,N_22535,N_22473);
nand U23035 (N_23035,N_22215,N_22152);
or U23036 (N_23036,N_22252,N_22312);
nor U23037 (N_23037,N_22639,N_22404);
or U23038 (N_23038,N_22624,N_22502);
or U23039 (N_23039,N_22112,N_22505);
and U23040 (N_23040,N_22776,N_22982);
nor U23041 (N_23041,N_22748,N_22516);
xnor U23042 (N_23042,N_22458,N_22129);
and U23043 (N_23043,N_22454,N_22626);
and U23044 (N_23044,N_22366,N_22674);
xor U23045 (N_23045,N_22159,N_22397);
xor U23046 (N_23046,N_22836,N_22180);
or U23047 (N_23047,N_22232,N_22126);
and U23048 (N_23048,N_22263,N_22844);
and U23049 (N_23049,N_22668,N_22260);
nor U23050 (N_23050,N_22977,N_22418);
or U23051 (N_23051,N_22492,N_22323);
or U23052 (N_23052,N_22712,N_22777);
xor U23053 (N_23053,N_22650,N_22837);
nand U23054 (N_23054,N_22567,N_22163);
nor U23055 (N_23055,N_22189,N_22436);
or U23056 (N_23056,N_22407,N_22235);
nor U23057 (N_23057,N_22760,N_22622);
and U23058 (N_23058,N_22005,N_22380);
xor U23059 (N_23059,N_22595,N_22512);
nand U23060 (N_23060,N_22093,N_22570);
or U23061 (N_23061,N_22245,N_22564);
nor U23062 (N_23062,N_22052,N_22830);
and U23063 (N_23063,N_22827,N_22918);
xor U23064 (N_23064,N_22374,N_22821);
nand U23065 (N_23065,N_22213,N_22306);
nand U23066 (N_23066,N_22892,N_22343);
nand U23067 (N_23067,N_22354,N_22986);
nor U23068 (N_23068,N_22611,N_22589);
nor U23069 (N_23069,N_22873,N_22887);
nor U23070 (N_23070,N_22035,N_22137);
xor U23071 (N_23071,N_22084,N_22270);
xor U23072 (N_23072,N_22934,N_22305);
and U23073 (N_23073,N_22657,N_22161);
and U23074 (N_23074,N_22583,N_22471);
nand U23075 (N_23075,N_22722,N_22335);
nor U23076 (N_23076,N_22314,N_22510);
xnor U23077 (N_23077,N_22025,N_22546);
nand U23078 (N_23078,N_22728,N_22714);
nor U23079 (N_23079,N_22277,N_22104);
nand U23080 (N_23080,N_22898,N_22179);
xnor U23081 (N_23081,N_22809,N_22805);
or U23082 (N_23082,N_22962,N_22793);
and U23083 (N_23083,N_22010,N_22654);
and U23084 (N_23084,N_22922,N_22839);
and U23085 (N_23085,N_22816,N_22287);
xor U23086 (N_23086,N_22139,N_22021);
or U23087 (N_23087,N_22296,N_22676);
nand U23088 (N_23088,N_22504,N_22440);
and U23089 (N_23089,N_22229,N_22610);
or U23090 (N_23090,N_22470,N_22644);
nand U23091 (N_23091,N_22966,N_22355);
or U23092 (N_23092,N_22715,N_22530);
nor U23093 (N_23093,N_22710,N_22975);
nand U23094 (N_23094,N_22158,N_22620);
nor U23095 (N_23095,N_22603,N_22846);
nor U23096 (N_23096,N_22613,N_22540);
or U23097 (N_23097,N_22716,N_22906);
or U23098 (N_23098,N_22274,N_22810);
nor U23099 (N_23099,N_22162,N_22135);
or U23100 (N_23100,N_22834,N_22963);
and U23101 (N_23101,N_22704,N_22032);
xor U23102 (N_23102,N_22787,N_22880);
nor U23103 (N_23103,N_22170,N_22662);
or U23104 (N_23104,N_22209,N_22557);
nor U23105 (N_23105,N_22957,N_22794);
nand U23106 (N_23106,N_22762,N_22482);
xnor U23107 (N_23107,N_22831,N_22993);
nand U23108 (N_23108,N_22623,N_22905);
or U23109 (N_23109,N_22698,N_22771);
and U23110 (N_23110,N_22544,N_22186);
nor U23111 (N_23111,N_22690,N_22985);
xor U23112 (N_23112,N_22528,N_22325);
and U23113 (N_23113,N_22636,N_22082);
nand U23114 (N_23114,N_22980,N_22476);
nand U23115 (N_23115,N_22819,N_22466);
nor U23116 (N_23116,N_22609,N_22070);
xnor U23117 (N_23117,N_22331,N_22749);
or U23118 (N_23118,N_22717,N_22818);
and U23119 (N_23119,N_22119,N_22264);
nand U23120 (N_23120,N_22747,N_22751);
xor U23121 (N_23121,N_22883,N_22097);
or U23122 (N_23122,N_22389,N_22849);
xnor U23123 (N_23123,N_22702,N_22689);
xnor U23124 (N_23124,N_22775,N_22143);
nand U23125 (N_23125,N_22381,N_22003);
and U23126 (N_23126,N_22856,N_22876);
nand U23127 (N_23127,N_22780,N_22140);
nand U23128 (N_23128,N_22591,N_22920);
nand U23129 (N_23129,N_22428,N_22236);
or U23130 (N_23130,N_22442,N_22487);
and U23131 (N_23131,N_22561,N_22048);
xnor U23132 (N_23132,N_22011,N_22318);
or U23133 (N_23133,N_22700,N_22479);
or U23134 (N_23134,N_22000,N_22969);
or U23135 (N_23135,N_22281,N_22046);
xor U23136 (N_23136,N_22503,N_22413);
nand U23137 (N_23137,N_22339,N_22594);
nand U23138 (N_23138,N_22902,N_22110);
and U23139 (N_23139,N_22649,N_22631);
or U23140 (N_23140,N_22637,N_22548);
xor U23141 (N_23141,N_22736,N_22480);
nor U23142 (N_23142,N_22246,N_22640);
nand U23143 (N_23143,N_22022,N_22795);
nand U23144 (N_23144,N_22164,N_22486);
and U23145 (N_23145,N_22151,N_22211);
and U23146 (N_23146,N_22387,N_22198);
nand U23147 (N_23147,N_22709,N_22746);
nand U23148 (N_23148,N_22953,N_22995);
xor U23149 (N_23149,N_22201,N_22896);
or U23150 (N_23150,N_22327,N_22185);
nand U23151 (N_23151,N_22410,N_22243);
nor U23152 (N_23152,N_22990,N_22757);
and U23153 (N_23153,N_22981,N_22814);
or U23154 (N_23154,N_22525,N_22117);
or U23155 (N_23155,N_22067,N_22449);
or U23156 (N_23156,N_22761,N_22064);
nand U23157 (N_23157,N_22019,N_22884);
nand U23158 (N_23158,N_22313,N_22563);
nand U23159 (N_23159,N_22108,N_22812);
or U23160 (N_23160,N_22373,N_22597);
nand U23161 (N_23161,N_22265,N_22932);
or U23162 (N_23162,N_22566,N_22099);
or U23163 (N_23163,N_22645,N_22462);
nand U23164 (N_23164,N_22721,N_22853);
or U23165 (N_23165,N_22169,N_22670);
nor U23166 (N_23166,N_22732,N_22020);
nand U23167 (N_23167,N_22695,N_22092);
nor U23168 (N_23168,N_22868,N_22259);
xor U23169 (N_23169,N_22452,N_22116);
nor U23170 (N_23170,N_22073,N_22669);
nor U23171 (N_23171,N_22177,N_22802);
xor U23172 (N_23172,N_22974,N_22133);
and U23173 (N_23173,N_22964,N_22155);
and U23174 (N_23174,N_22823,N_22522);
and U23175 (N_23175,N_22317,N_22435);
or U23176 (N_23176,N_22944,N_22489);
and U23177 (N_23177,N_22171,N_22808);
nand U23178 (N_23178,N_22562,N_22128);
nand U23179 (N_23179,N_22027,N_22172);
and U23180 (N_23180,N_22324,N_22847);
nor U23181 (N_23181,N_22592,N_22446);
xnor U23182 (N_23182,N_22390,N_22766);
xor U23183 (N_23183,N_22792,N_22531);
and U23184 (N_23184,N_22743,N_22465);
nor U23185 (N_23185,N_22148,N_22641);
nor U23186 (N_23186,N_22311,N_22890);
xnor U23187 (N_23187,N_22731,N_22474);
nand U23188 (N_23188,N_22739,N_22612);
nand U23189 (N_23189,N_22988,N_22520);
nor U23190 (N_23190,N_22300,N_22590);
and U23191 (N_23191,N_22874,N_22055);
and U23192 (N_23192,N_22036,N_22045);
nor U23193 (N_23193,N_22927,N_22191);
and U23194 (N_23194,N_22131,N_22615);
nand U23195 (N_23195,N_22677,N_22016);
nand U23196 (N_23196,N_22176,N_22534);
and U23197 (N_23197,N_22586,N_22004);
and U23198 (N_23198,N_22899,N_22838);
xor U23199 (N_23199,N_22483,N_22220);
or U23200 (N_23200,N_22194,N_22582);
and U23201 (N_23201,N_22678,N_22338);
and U23202 (N_23202,N_22574,N_22276);
nor U23203 (N_23203,N_22142,N_22102);
nand U23204 (N_23204,N_22219,N_22629);
xor U23205 (N_23205,N_22864,N_22351);
nor U23206 (N_23206,N_22877,N_22309);
xnor U23207 (N_23207,N_22225,N_22608);
nor U23208 (N_23208,N_22076,N_22683);
xor U23209 (N_23209,N_22687,N_22931);
nor U23210 (N_23210,N_22568,N_22051);
nor U23211 (N_23211,N_22271,N_22845);
and U23212 (N_23212,N_22577,N_22205);
or U23213 (N_23213,N_22227,N_22488);
or U23214 (N_23214,N_22854,N_22679);
nand U23215 (N_23215,N_22217,N_22691);
nor U23216 (N_23216,N_22681,N_22365);
nor U23217 (N_23217,N_22956,N_22915);
and U23218 (N_23218,N_22571,N_22240);
nor U23219 (N_23219,N_22187,N_22059);
or U23220 (N_23220,N_22353,N_22917);
nand U23221 (N_23221,N_22885,N_22031);
nor U23222 (N_23222,N_22098,N_22765);
nand U23223 (N_23223,N_22258,N_22869);
xor U23224 (N_23224,N_22167,N_22028);
or U23225 (N_23225,N_22587,N_22299);
nand U23226 (N_23226,N_22293,N_22282);
nor U23227 (N_23227,N_22014,N_22118);
nand U23228 (N_23228,N_22332,N_22524);
xor U23229 (N_23229,N_22904,N_22507);
xor U23230 (N_23230,N_22310,N_22234);
or U23231 (N_23231,N_22686,N_22954);
nand U23232 (N_23232,N_22653,N_22481);
nand U23233 (N_23233,N_22782,N_22477);
nor U23234 (N_23234,N_22938,N_22315);
nand U23235 (N_23235,N_22249,N_22393);
nor U23236 (N_23236,N_22464,N_22519);
xnor U23237 (N_23237,N_22086,N_22146);
nor U23238 (N_23238,N_22879,N_22556);
nor U23239 (N_23239,N_22718,N_22784);
nand U23240 (N_23240,N_22559,N_22439);
nor U23241 (N_23241,N_22634,N_22242);
xor U23242 (N_23242,N_22072,N_22857);
nand U23243 (N_23243,N_22937,N_22999);
or U23244 (N_23244,N_22041,N_22797);
or U23245 (N_23245,N_22412,N_22575);
and U23246 (N_23246,N_22337,N_22149);
xor U23247 (N_23247,N_22788,N_22350);
and U23248 (N_23248,N_22278,N_22729);
nor U23249 (N_23249,N_22870,N_22196);
and U23250 (N_23250,N_22453,N_22842);
nand U23251 (N_23251,N_22506,N_22208);
and U23252 (N_23252,N_22537,N_22606);
and U23253 (N_23253,N_22496,N_22786);
xor U23254 (N_23254,N_22168,N_22817);
xor U23255 (N_23255,N_22065,N_22266);
or U23256 (N_23256,N_22866,N_22713);
and U23257 (N_23257,N_22083,N_22372);
or U23258 (N_23258,N_22984,N_22971);
nor U23259 (N_23259,N_22319,N_22888);
nor U23260 (N_23260,N_22848,N_22256);
or U23261 (N_23261,N_22536,N_22445);
nand U23262 (N_23262,N_22212,N_22370);
nor U23263 (N_23263,N_22773,N_22860);
nand U23264 (N_23264,N_22068,N_22382);
xor U23265 (N_23265,N_22960,N_22214);
and U23266 (N_23266,N_22304,N_22642);
or U23267 (N_23267,N_22095,N_22111);
nor U23268 (N_23268,N_22414,N_22203);
nand U23269 (N_23269,N_22855,N_22921);
nand U23270 (N_23270,N_22223,N_22386);
xnor U23271 (N_23271,N_22497,N_22741);
nor U23272 (N_23272,N_22006,N_22257);
and U23273 (N_23273,N_22134,N_22114);
nand U23274 (N_23274,N_22206,N_22132);
or U23275 (N_23275,N_22268,N_22284);
or U23276 (N_23276,N_22017,N_22286);
or U23277 (N_23277,N_22123,N_22970);
and U23278 (N_23278,N_22181,N_22752);
nand U23279 (N_23279,N_22138,N_22926);
xor U23280 (N_23280,N_22307,N_22878);
or U23281 (N_23281,N_22468,N_22588);
nand U23282 (N_23282,N_22843,N_22456);
xnor U23283 (N_23283,N_22434,N_22925);
nand U23284 (N_23284,N_22665,N_22165);
or U23285 (N_23285,N_22983,N_22460);
xor U23286 (N_23286,N_22554,N_22648);
xor U23287 (N_23287,N_22744,N_22673);
or U23288 (N_23288,N_22916,N_22628);
nand U23289 (N_23289,N_22253,N_22224);
or U23290 (N_23290,N_22545,N_22529);
xnor U23291 (N_23291,N_22417,N_22419);
xor U23292 (N_23292,N_22935,N_22207);
nand U23293 (N_23293,N_22406,N_22075);
and U23294 (N_23294,N_22621,N_22774);
and U23295 (N_23295,N_22395,N_22851);
and U23296 (N_23296,N_22369,N_22030);
nor U23297 (N_23297,N_22283,N_22705);
and U23298 (N_23298,N_22120,N_22074);
nand U23299 (N_23299,N_22290,N_22987);
and U23300 (N_23300,N_22785,N_22614);
xor U23301 (N_23301,N_22396,N_22919);
and U23302 (N_23302,N_22897,N_22034);
nor U23303 (N_23303,N_22320,N_22499);
and U23304 (N_23304,N_22192,N_22825);
nor U23305 (N_23305,N_22244,N_22948);
nand U23306 (N_23306,N_22272,N_22523);
nor U23307 (N_23307,N_22427,N_22552);
and U23308 (N_23308,N_22438,N_22361);
or U23309 (N_23309,N_22100,N_22989);
and U23310 (N_23310,N_22360,N_22852);
nand U23311 (N_23311,N_22632,N_22448);
xnor U23312 (N_23312,N_22367,N_22493);
nand U23313 (N_23313,N_22607,N_22889);
or U23314 (N_23314,N_22383,N_22175);
nand U23315 (N_23315,N_22933,N_22719);
nand U23316 (N_23316,N_22781,N_22371);
and U23317 (N_23317,N_22924,N_22501);
nand U23318 (N_23318,N_22357,N_22949);
nor U23319 (N_23319,N_22798,N_22633);
and U23320 (N_23320,N_22997,N_22872);
and U23321 (N_23321,N_22711,N_22432);
and U23322 (N_23322,N_22239,N_22391);
or U23323 (N_23323,N_22292,N_22248);
or U23324 (N_23324,N_22976,N_22080);
and U23325 (N_23325,N_22349,N_22461);
nor U23326 (N_23326,N_22498,N_22392);
or U23327 (N_23327,N_22024,N_22772);
or U23328 (N_23328,N_22940,N_22136);
nand U23329 (N_23329,N_22422,N_22231);
xor U23330 (N_23330,N_22160,N_22707);
or U23331 (N_23331,N_22044,N_22576);
and U23332 (N_23332,N_22409,N_22911);
and U23333 (N_23333,N_22437,N_22593);
xnor U23334 (N_23334,N_22734,N_22804);
nor U23335 (N_23335,N_22929,N_22195);
nor U23336 (N_23336,N_22221,N_22778);
nand U23337 (N_23337,N_22725,N_22923);
nor U23338 (N_23338,N_22193,N_22913);
nand U23339 (N_23339,N_22754,N_22012);
or U23340 (N_23340,N_22280,N_22951);
nand U23341 (N_23341,N_22824,N_22182);
xor U23342 (N_23342,N_22183,N_22753);
xnor U23343 (N_23343,N_22735,N_22551);
xor U23344 (N_23344,N_22144,N_22871);
nand U23345 (N_23345,N_22153,N_22101);
xor U23346 (N_23346,N_22125,N_22881);
nand U23347 (N_23347,N_22421,N_22580);
xnor U23348 (N_23348,N_22893,N_22533);
xnor U23349 (N_23349,N_22672,N_22894);
and U23350 (N_23350,N_22222,N_22115);
xnor U23351 (N_23351,N_22174,N_22178);
or U23352 (N_23352,N_22758,N_22667);
xor U23353 (N_23353,N_22618,N_22832);
nand U23354 (N_23354,N_22909,N_22420);
nor U23355 (N_23355,N_22684,N_22820);
and U23356 (N_23356,N_22945,N_22532);
xor U23357 (N_23357,N_22424,N_22549);
nor U23358 (N_23358,N_22900,N_22250);
xor U23359 (N_23359,N_22750,N_22903);
and U23360 (N_23360,N_22301,N_22991);
and U23361 (N_23361,N_22475,N_22965);
nand U23362 (N_23362,N_22238,N_22455);
xnor U23363 (N_23363,N_22643,N_22364);
and U23364 (N_23364,N_22375,N_22769);
or U23365 (N_23365,N_22385,N_22500);
or U23366 (N_23366,N_22121,N_22297);
and U23367 (N_23367,N_22550,N_22675);
or U23368 (N_23368,N_22457,N_22326);
nor U23369 (N_23369,N_22585,N_22968);
and U23370 (N_23370,N_22275,N_22443);
and U23371 (N_23371,N_22049,N_22009);
xnor U23372 (N_23372,N_22321,N_22518);
nor U23373 (N_23373,N_22617,N_22912);
xnor U23374 (N_23374,N_22727,N_22596);
nor U23375 (N_23375,N_22166,N_22103);
nand U23376 (N_23376,N_22237,N_22463);
nand U23377 (N_23377,N_22368,N_22660);
nor U23378 (N_23378,N_22451,N_22791);
xnor U23379 (N_23379,N_22042,N_22763);
or U23380 (N_23380,N_22033,N_22616);
nand U23381 (N_23381,N_22699,N_22602);
or U23382 (N_23382,N_22807,N_22060);
and U23383 (N_23383,N_22875,N_22061);
nand U23384 (N_23384,N_22539,N_22910);
nor U23385 (N_23385,N_22069,N_22394);
nand U23386 (N_23386,N_22150,N_22811);
nor U23387 (N_23387,N_22967,N_22569);
xnor U23388 (N_23388,N_22154,N_22619);
or U23389 (N_23389,N_22755,N_22001);
or U23390 (N_23390,N_22429,N_22113);
and U23391 (N_23391,N_22405,N_22992);
and U23392 (N_23392,N_22979,N_22130);
or U23393 (N_23393,N_22862,N_22950);
nor U23394 (N_23394,N_22106,N_22835);
and U23395 (N_23395,N_22285,N_22216);
or U23396 (N_23396,N_22646,N_22961);
and U23397 (N_23397,N_22859,N_22491);
and U23398 (N_23398,N_22091,N_22581);
and U23399 (N_23399,N_22441,N_22018);
xnor U23400 (N_23400,N_22796,N_22730);
or U23401 (N_23401,N_22400,N_22604);
or U23402 (N_23402,N_22226,N_22661);
and U23403 (N_23403,N_22696,N_22694);
nor U23404 (N_23404,N_22701,N_22789);
nand U23405 (N_23405,N_22200,N_22273);
xnor U23406 (N_23406,N_22342,N_22334);
or U23407 (N_23407,N_22543,N_22901);
or U23408 (N_23408,N_22647,N_22251);
nand U23409 (N_23409,N_22288,N_22625);
xnor U23410 (N_23410,N_22998,N_22955);
nor U23411 (N_23411,N_22233,N_22826);
or U23412 (N_23412,N_22403,N_22348);
or U23413 (N_23413,N_22865,N_22444);
and U23414 (N_23414,N_22345,N_22359);
and U23415 (N_23415,N_22630,N_22040);
xor U23416 (N_23416,N_22720,N_22599);
and U23417 (N_23417,N_22726,N_22402);
nand U23418 (N_23418,N_22996,N_22939);
nor U23419 (N_23419,N_22322,N_22664);
and U23420 (N_23420,N_22379,N_22886);
nand U23421 (N_23421,N_22666,N_22090);
or U23422 (N_23422,N_22656,N_22745);
nor U23423 (N_23423,N_22430,N_22882);
xnor U23424 (N_23424,N_22655,N_22768);
xnor U23425 (N_23425,N_22494,N_22261);
and U23426 (N_23426,N_22199,N_22340);
xor U23427 (N_23427,N_22994,N_22295);
xnor U23428 (N_23428,N_22425,N_22692);
nor U23429 (N_23429,N_22509,N_22973);
nor U23430 (N_23430,N_22560,N_22328);
nor U23431 (N_23431,N_22363,N_22378);
xnor U23432 (N_23432,N_22605,N_22401);
and U23433 (N_23433,N_22914,N_22037);
and U23434 (N_23434,N_22352,N_22467);
nand U23435 (N_23435,N_22254,N_22247);
nand U23436 (N_23436,N_22077,N_22638);
or U23437 (N_23437,N_22377,N_22930);
nand U23438 (N_23438,N_22415,N_22685);
or U23439 (N_23439,N_22002,N_22267);
xnor U23440 (N_23440,N_22384,N_22517);
xnor U23441 (N_23441,N_22303,N_22867);
nand U23442 (N_23442,N_22478,N_22783);
and U23443 (N_23443,N_22054,N_22558);
and U23444 (N_23444,N_22738,N_22122);
nand U23445 (N_23445,N_22770,N_22508);
or U23446 (N_23446,N_22089,N_22861);
nand U23447 (N_23447,N_22141,N_22469);
nand U23448 (N_23448,N_22431,N_22459);
nand U23449 (N_23449,N_22841,N_22147);
and U23450 (N_23450,N_22050,N_22416);
and U23451 (N_23451,N_22329,N_22085);
nand U23452 (N_23452,N_22800,N_22096);
or U23453 (N_23453,N_22693,N_22799);
nand U23454 (N_23454,N_22078,N_22706);
nor U23455 (N_23455,N_22145,N_22946);
xnor U23456 (N_23456,N_22087,N_22740);
xor U23457 (N_23457,N_22801,N_22341);
nor U23458 (N_23458,N_22039,N_22863);
or U23459 (N_23459,N_22124,N_22978);
nor U23460 (N_23460,N_22928,N_22269);
and U23461 (N_23461,N_22472,N_22941);
nor U23462 (N_23462,N_22157,N_22255);
and U23463 (N_23463,N_22958,N_22347);
nand U23464 (N_23464,N_22330,N_22279);
xnor U23465 (N_23465,N_22943,N_22399);
nor U23466 (N_23466,N_22542,N_22202);
xor U23467 (N_23467,N_22651,N_22043);
and U23468 (N_23468,N_22388,N_22204);
and U23469 (N_23469,N_22127,N_22555);
and U23470 (N_23470,N_22733,N_22942);
xor U23471 (N_23471,N_22358,N_22779);
nand U23472 (N_23472,N_22218,N_22553);
and U23473 (N_23473,N_22485,N_22308);
or U23474 (N_23474,N_22013,N_22598);
and U23475 (N_23475,N_22680,N_22907);
xor U23476 (N_23476,N_22447,N_22071);
and U23477 (N_23477,N_22294,N_22565);
nor U23478 (N_23478,N_22828,N_22411);
and U23479 (N_23479,N_22600,N_22495);
xnor U23480 (N_23480,N_22173,N_22056);
xor U23481 (N_23481,N_22408,N_22514);
or U23482 (N_23482,N_22094,N_22079);
xor U23483 (N_23483,N_22450,N_22188);
xnor U23484 (N_23484,N_22262,N_22703);
nand U23485 (N_23485,N_22344,N_22635);
xnor U23486 (N_23486,N_22298,N_22484);
or U23487 (N_23487,N_22790,N_22376);
and U23488 (N_23488,N_22947,N_22806);
nor U23489 (N_23489,N_22767,N_22007);
or U23490 (N_23490,N_22822,N_22737);
nor U23491 (N_23491,N_22289,N_22526);
nor U23492 (N_23492,N_22573,N_22697);
or U23493 (N_23493,N_22398,N_22521);
or U23494 (N_23494,N_22708,N_22671);
xnor U23495 (N_23495,N_22663,N_22081);
and U23496 (N_23496,N_22356,N_22230);
nor U23497 (N_23497,N_22058,N_22057);
and U23498 (N_23498,N_22652,N_22026);
nand U23499 (N_23499,N_22601,N_22515);
nor U23500 (N_23500,N_22378,N_22337);
nor U23501 (N_23501,N_22455,N_22594);
or U23502 (N_23502,N_22887,N_22453);
and U23503 (N_23503,N_22804,N_22942);
nor U23504 (N_23504,N_22219,N_22331);
and U23505 (N_23505,N_22536,N_22045);
xor U23506 (N_23506,N_22565,N_22682);
xor U23507 (N_23507,N_22544,N_22308);
or U23508 (N_23508,N_22808,N_22862);
and U23509 (N_23509,N_22307,N_22371);
or U23510 (N_23510,N_22958,N_22613);
and U23511 (N_23511,N_22634,N_22023);
xor U23512 (N_23512,N_22840,N_22860);
nand U23513 (N_23513,N_22454,N_22244);
nand U23514 (N_23514,N_22640,N_22727);
nor U23515 (N_23515,N_22439,N_22720);
xnor U23516 (N_23516,N_22401,N_22771);
or U23517 (N_23517,N_22658,N_22597);
nor U23518 (N_23518,N_22245,N_22613);
or U23519 (N_23519,N_22727,N_22890);
or U23520 (N_23520,N_22004,N_22533);
xor U23521 (N_23521,N_22381,N_22146);
xnor U23522 (N_23522,N_22979,N_22797);
nand U23523 (N_23523,N_22914,N_22680);
and U23524 (N_23524,N_22835,N_22574);
xor U23525 (N_23525,N_22877,N_22899);
nor U23526 (N_23526,N_22586,N_22220);
and U23527 (N_23527,N_22543,N_22244);
nand U23528 (N_23528,N_22677,N_22797);
nor U23529 (N_23529,N_22863,N_22676);
or U23530 (N_23530,N_22263,N_22559);
nand U23531 (N_23531,N_22600,N_22462);
or U23532 (N_23532,N_22651,N_22277);
nor U23533 (N_23533,N_22841,N_22877);
or U23534 (N_23534,N_22790,N_22064);
and U23535 (N_23535,N_22533,N_22770);
nor U23536 (N_23536,N_22689,N_22501);
or U23537 (N_23537,N_22041,N_22569);
or U23538 (N_23538,N_22050,N_22113);
nand U23539 (N_23539,N_22199,N_22141);
or U23540 (N_23540,N_22917,N_22091);
nor U23541 (N_23541,N_22486,N_22153);
or U23542 (N_23542,N_22252,N_22594);
xor U23543 (N_23543,N_22850,N_22510);
nand U23544 (N_23544,N_22290,N_22441);
or U23545 (N_23545,N_22087,N_22916);
nor U23546 (N_23546,N_22478,N_22650);
nand U23547 (N_23547,N_22214,N_22891);
xor U23548 (N_23548,N_22193,N_22818);
or U23549 (N_23549,N_22982,N_22599);
nor U23550 (N_23550,N_22563,N_22428);
nand U23551 (N_23551,N_22897,N_22112);
and U23552 (N_23552,N_22307,N_22659);
or U23553 (N_23553,N_22912,N_22904);
xnor U23554 (N_23554,N_22980,N_22364);
or U23555 (N_23555,N_22218,N_22636);
nand U23556 (N_23556,N_22548,N_22090);
and U23557 (N_23557,N_22025,N_22189);
or U23558 (N_23558,N_22016,N_22979);
xnor U23559 (N_23559,N_22952,N_22716);
nand U23560 (N_23560,N_22360,N_22420);
and U23561 (N_23561,N_22943,N_22095);
nor U23562 (N_23562,N_22132,N_22381);
nor U23563 (N_23563,N_22771,N_22831);
and U23564 (N_23564,N_22825,N_22686);
and U23565 (N_23565,N_22742,N_22505);
xor U23566 (N_23566,N_22370,N_22696);
nor U23567 (N_23567,N_22562,N_22304);
or U23568 (N_23568,N_22179,N_22610);
xor U23569 (N_23569,N_22042,N_22509);
and U23570 (N_23570,N_22548,N_22885);
and U23571 (N_23571,N_22859,N_22950);
and U23572 (N_23572,N_22242,N_22100);
xor U23573 (N_23573,N_22884,N_22835);
xnor U23574 (N_23574,N_22740,N_22636);
xor U23575 (N_23575,N_22112,N_22499);
and U23576 (N_23576,N_22447,N_22048);
or U23577 (N_23577,N_22337,N_22928);
and U23578 (N_23578,N_22003,N_22365);
nand U23579 (N_23579,N_22676,N_22062);
and U23580 (N_23580,N_22527,N_22116);
nor U23581 (N_23581,N_22249,N_22460);
nand U23582 (N_23582,N_22543,N_22583);
or U23583 (N_23583,N_22594,N_22526);
or U23584 (N_23584,N_22135,N_22506);
xnor U23585 (N_23585,N_22240,N_22307);
nand U23586 (N_23586,N_22188,N_22030);
or U23587 (N_23587,N_22159,N_22036);
nand U23588 (N_23588,N_22155,N_22003);
and U23589 (N_23589,N_22073,N_22447);
and U23590 (N_23590,N_22317,N_22645);
or U23591 (N_23591,N_22362,N_22612);
xor U23592 (N_23592,N_22127,N_22103);
or U23593 (N_23593,N_22039,N_22970);
nand U23594 (N_23594,N_22069,N_22788);
nor U23595 (N_23595,N_22235,N_22818);
or U23596 (N_23596,N_22727,N_22526);
or U23597 (N_23597,N_22204,N_22776);
xnor U23598 (N_23598,N_22627,N_22178);
xnor U23599 (N_23599,N_22846,N_22809);
and U23600 (N_23600,N_22428,N_22188);
nor U23601 (N_23601,N_22470,N_22044);
or U23602 (N_23602,N_22750,N_22954);
nor U23603 (N_23603,N_22240,N_22382);
or U23604 (N_23604,N_22323,N_22851);
nand U23605 (N_23605,N_22579,N_22909);
and U23606 (N_23606,N_22154,N_22256);
xor U23607 (N_23607,N_22795,N_22206);
nand U23608 (N_23608,N_22213,N_22411);
nand U23609 (N_23609,N_22666,N_22087);
and U23610 (N_23610,N_22807,N_22984);
or U23611 (N_23611,N_22666,N_22553);
nor U23612 (N_23612,N_22022,N_22633);
xnor U23613 (N_23613,N_22604,N_22732);
xor U23614 (N_23614,N_22182,N_22951);
nor U23615 (N_23615,N_22935,N_22452);
nand U23616 (N_23616,N_22169,N_22902);
xnor U23617 (N_23617,N_22191,N_22356);
xnor U23618 (N_23618,N_22184,N_22750);
nand U23619 (N_23619,N_22565,N_22419);
or U23620 (N_23620,N_22371,N_22129);
and U23621 (N_23621,N_22149,N_22787);
and U23622 (N_23622,N_22374,N_22166);
and U23623 (N_23623,N_22840,N_22948);
nor U23624 (N_23624,N_22980,N_22467);
or U23625 (N_23625,N_22515,N_22441);
or U23626 (N_23626,N_22687,N_22257);
nor U23627 (N_23627,N_22175,N_22464);
nand U23628 (N_23628,N_22201,N_22065);
or U23629 (N_23629,N_22863,N_22885);
nor U23630 (N_23630,N_22417,N_22054);
nor U23631 (N_23631,N_22642,N_22292);
or U23632 (N_23632,N_22637,N_22612);
and U23633 (N_23633,N_22690,N_22027);
nor U23634 (N_23634,N_22637,N_22215);
or U23635 (N_23635,N_22825,N_22460);
nor U23636 (N_23636,N_22172,N_22184);
xnor U23637 (N_23637,N_22697,N_22061);
or U23638 (N_23638,N_22359,N_22994);
and U23639 (N_23639,N_22929,N_22199);
xor U23640 (N_23640,N_22923,N_22336);
xor U23641 (N_23641,N_22698,N_22776);
or U23642 (N_23642,N_22685,N_22589);
xnor U23643 (N_23643,N_22444,N_22605);
nand U23644 (N_23644,N_22890,N_22035);
and U23645 (N_23645,N_22667,N_22978);
xor U23646 (N_23646,N_22378,N_22037);
nor U23647 (N_23647,N_22402,N_22155);
and U23648 (N_23648,N_22082,N_22813);
nor U23649 (N_23649,N_22191,N_22225);
or U23650 (N_23650,N_22897,N_22560);
or U23651 (N_23651,N_22774,N_22158);
and U23652 (N_23652,N_22794,N_22931);
nor U23653 (N_23653,N_22100,N_22068);
nor U23654 (N_23654,N_22863,N_22343);
nor U23655 (N_23655,N_22294,N_22720);
xor U23656 (N_23656,N_22784,N_22521);
nand U23657 (N_23657,N_22555,N_22303);
nor U23658 (N_23658,N_22288,N_22898);
or U23659 (N_23659,N_22918,N_22529);
or U23660 (N_23660,N_22737,N_22651);
or U23661 (N_23661,N_22402,N_22903);
xnor U23662 (N_23662,N_22836,N_22484);
nor U23663 (N_23663,N_22616,N_22287);
or U23664 (N_23664,N_22449,N_22633);
and U23665 (N_23665,N_22012,N_22340);
xnor U23666 (N_23666,N_22869,N_22892);
or U23667 (N_23667,N_22660,N_22294);
nor U23668 (N_23668,N_22297,N_22556);
nor U23669 (N_23669,N_22571,N_22245);
and U23670 (N_23670,N_22782,N_22778);
nor U23671 (N_23671,N_22411,N_22512);
nand U23672 (N_23672,N_22160,N_22994);
xor U23673 (N_23673,N_22035,N_22132);
or U23674 (N_23674,N_22646,N_22998);
nor U23675 (N_23675,N_22331,N_22523);
nand U23676 (N_23676,N_22869,N_22889);
xnor U23677 (N_23677,N_22338,N_22517);
nor U23678 (N_23678,N_22854,N_22622);
xor U23679 (N_23679,N_22895,N_22321);
or U23680 (N_23680,N_22426,N_22974);
or U23681 (N_23681,N_22353,N_22728);
or U23682 (N_23682,N_22506,N_22802);
xnor U23683 (N_23683,N_22342,N_22663);
nor U23684 (N_23684,N_22396,N_22253);
or U23685 (N_23685,N_22057,N_22569);
nor U23686 (N_23686,N_22566,N_22572);
or U23687 (N_23687,N_22757,N_22015);
nor U23688 (N_23688,N_22781,N_22396);
nor U23689 (N_23689,N_22553,N_22568);
xnor U23690 (N_23690,N_22039,N_22708);
nor U23691 (N_23691,N_22963,N_22698);
xnor U23692 (N_23692,N_22419,N_22199);
xor U23693 (N_23693,N_22113,N_22145);
or U23694 (N_23694,N_22423,N_22782);
nand U23695 (N_23695,N_22859,N_22968);
nand U23696 (N_23696,N_22270,N_22370);
xnor U23697 (N_23697,N_22429,N_22623);
and U23698 (N_23698,N_22980,N_22115);
xor U23699 (N_23699,N_22036,N_22263);
xor U23700 (N_23700,N_22691,N_22492);
xnor U23701 (N_23701,N_22311,N_22697);
and U23702 (N_23702,N_22333,N_22893);
xor U23703 (N_23703,N_22572,N_22149);
nand U23704 (N_23704,N_22265,N_22259);
nand U23705 (N_23705,N_22843,N_22601);
nand U23706 (N_23706,N_22165,N_22208);
nor U23707 (N_23707,N_22773,N_22688);
nor U23708 (N_23708,N_22022,N_22762);
nor U23709 (N_23709,N_22299,N_22062);
nor U23710 (N_23710,N_22633,N_22741);
nand U23711 (N_23711,N_22637,N_22162);
xnor U23712 (N_23712,N_22534,N_22636);
nand U23713 (N_23713,N_22237,N_22467);
or U23714 (N_23714,N_22222,N_22330);
and U23715 (N_23715,N_22163,N_22964);
xnor U23716 (N_23716,N_22688,N_22845);
nand U23717 (N_23717,N_22560,N_22388);
nor U23718 (N_23718,N_22534,N_22585);
and U23719 (N_23719,N_22436,N_22272);
xnor U23720 (N_23720,N_22148,N_22797);
and U23721 (N_23721,N_22563,N_22279);
and U23722 (N_23722,N_22589,N_22585);
xor U23723 (N_23723,N_22766,N_22183);
nand U23724 (N_23724,N_22018,N_22292);
and U23725 (N_23725,N_22949,N_22908);
and U23726 (N_23726,N_22461,N_22547);
and U23727 (N_23727,N_22365,N_22114);
or U23728 (N_23728,N_22210,N_22017);
and U23729 (N_23729,N_22117,N_22813);
xnor U23730 (N_23730,N_22851,N_22358);
and U23731 (N_23731,N_22535,N_22866);
xor U23732 (N_23732,N_22027,N_22827);
nor U23733 (N_23733,N_22863,N_22848);
or U23734 (N_23734,N_22861,N_22647);
and U23735 (N_23735,N_22917,N_22815);
or U23736 (N_23736,N_22265,N_22390);
nand U23737 (N_23737,N_22982,N_22299);
and U23738 (N_23738,N_22469,N_22054);
or U23739 (N_23739,N_22752,N_22520);
or U23740 (N_23740,N_22940,N_22204);
or U23741 (N_23741,N_22038,N_22794);
and U23742 (N_23742,N_22104,N_22643);
or U23743 (N_23743,N_22885,N_22918);
and U23744 (N_23744,N_22145,N_22134);
and U23745 (N_23745,N_22719,N_22760);
xnor U23746 (N_23746,N_22636,N_22994);
nand U23747 (N_23747,N_22846,N_22445);
or U23748 (N_23748,N_22982,N_22351);
xnor U23749 (N_23749,N_22840,N_22256);
and U23750 (N_23750,N_22828,N_22388);
xnor U23751 (N_23751,N_22737,N_22870);
and U23752 (N_23752,N_22926,N_22204);
nor U23753 (N_23753,N_22988,N_22961);
or U23754 (N_23754,N_22683,N_22271);
nor U23755 (N_23755,N_22171,N_22416);
xor U23756 (N_23756,N_22708,N_22093);
or U23757 (N_23757,N_22072,N_22057);
or U23758 (N_23758,N_22554,N_22711);
nor U23759 (N_23759,N_22923,N_22169);
nand U23760 (N_23760,N_22619,N_22218);
and U23761 (N_23761,N_22360,N_22462);
nor U23762 (N_23762,N_22391,N_22998);
nand U23763 (N_23763,N_22509,N_22945);
nor U23764 (N_23764,N_22036,N_22910);
xnor U23765 (N_23765,N_22880,N_22171);
nor U23766 (N_23766,N_22568,N_22734);
and U23767 (N_23767,N_22843,N_22837);
nand U23768 (N_23768,N_22518,N_22920);
nand U23769 (N_23769,N_22843,N_22881);
nor U23770 (N_23770,N_22101,N_22205);
or U23771 (N_23771,N_22337,N_22042);
and U23772 (N_23772,N_22045,N_22002);
xnor U23773 (N_23773,N_22916,N_22394);
and U23774 (N_23774,N_22278,N_22345);
and U23775 (N_23775,N_22773,N_22057);
nand U23776 (N_23776,N_22790,N_22189);
or U23777 (N_23777,N_22292,N_22965);
and U23778 (N_23778,N_22829,N_22682);
xor U23779 (N_23779,N_22457,N_22214);
and U23780 (N_23780,N_22329,N_22218);
and U23781 (N_23781,N_22217,N_22470);
or U23782 (N_23782,N_22021,N_22448);
nand U23783 (N_23783,N_22893,N_22306);
nor U23784 (N_23784,N_22405,N_22191);
xnor U23785 (N_23785,N_22032,N_22208);
nand U23786 (N_23786,N_22404,N_22231);
or U23787 (N_23787,N_22092,N_22394);
xnor U23788 (N_23788,N_22405,N_22697);
xor U23789 (N_23789,N_22816,N_22679);
xnor U23790 (N_23790,N_22569,N_22666);
nand U23791 (N_23791,N_22373,N_22108);
and U23792 (N_23792,N_22964,N_22708);
and U23793 (N_23793,N_22337,N_22836);
or U23794 (N_23794,N_22683,N_22285);
nor U23795 (N_23795,N_22864,N_22936);
xor U23796 (N_23796,N_22545,N_22118);
nand U23797 (N_23797,N_22736,N_22455);
and U23798 (N_23798,N_22484,N_22007);
nor U23799 (N_23799,N_22038,N_22918);
and U23800 (N_23800,N_22281,N_22897);
nand U23801 (N_23801,N_22267,N_22574);
xnor U23802 (N_23802,N_22558,N_22220);
or U23803 (N_23803,N_22654,N_22669);
nand U23804 (N_23804,N_22136,N_22694);
xnor U23805 (N_23805,N_22730,N_22749);
xnor U23806 (N_23806,N_22162,N_22420);
xnor U23807 (N_23807,N_22029,N_22794);
xnor U23808 (N_23808,N_22682,N_22656);
or U23809 (N_23809,N_22995,N_22229);
nand U23810 (N_23810,N_22619,N_22616);
xor U23811 (N_23811,N_22857,N_22407);
xnor U23812 (N_23812,N_22599,N_22692);
xnor U23813 (N_23813,N_22938,N_22544);
nand U23814 (N_23814,N_22330,N_22119);
nand U23815 (N_23815,N_22579,N_22294);
nor U23816 (N_23816,N_22532,N_22198);
and U23817 (N_23817,N_22810,N_22129);
nor U23818 (N_23818,N_22569,N_22468);
nor U23819 (N_23819,N_22119,N_22702);
and U23820 (N_23820,N_22062,N_22823);
nand U23821 (N_23821,N_22285,N_22782);
or U23822 (N_23822,N_22651,N_22834);
and U23823 (N_23823,N_22519,N_22941);
xor U23824 (N_23824,N_22784,N_22329);
xor U23825 (N_23825,N_22182,N_22581);
xor U23826 (N_23826,N_22120,N_22535);
nor U23827 (N_23827,N_22037,N_22247);
or U23828 (N_23828,N_22417,N_22050);
or U23829 (N_23829,N_22409,N_22491);
nor U23830 (N_23830,N_22151,N_22316);
nor U23831 (N_23831,N_22592,N_22295);
nor U23832 (N_23832,N_22759,N_22253);
and U23833 (N_23833,N_22743,N_22641);
nor U23834 (N_23834,N_22877,N_22703);
xor U23835 (N_23835,N_22997,N_22126);
nor U23836 (N_23836,N_22380,N_22479);
nor U23837 (N_23837,N_22857,N_22642);
nor U23838 (N_23838,N_22428,N_22906);
xnor U23839 (N_23839,N_22393,N_22862);
or U23840 (N_23840,N_22083,N_22584);
and U23841 (N_23841,N_22986,N_22754);
or U23842 (N_23842,N_22672,N_22093);
nand U23843 (N_23843,N_22794,N_22792);
or U23844 (N_23844,N_22353,N_22661);
nand U23845 (N_23845,N_22919,N_22466);
or U23846 (N_23846,N_22749,N_22426);
and U23847 (N_23847,N_22232,N_22346);
nand U23848 (N_23848,N_22431,N_22082);
or U23849 (N_23849,N_22657,N_22033);
xor U23850 (N_23850,N_22799,N_22964);
or U23851 (N_23851,N_22060,N_22500);
and U23852 (N_23852,N_22255,N_22655);
nor U23853 (N_23853,N_22007,N_22989);
or U23854 (N_23854,N_22930,N_22136);
xor U23855 (N_23855,N_22090,N_22503);
nor U23856 (N_23856,N_22900,N_22127);
and U23857 (N_23857,N_22763,N_22987);
or U23858 (N_23858,N_22396,N_22388);
xor U23859 (N_23859,N_22160,N_22865);
xor U23860 (N_23860,N_22551,N_22245);
xnor U23861 (N_23861,N_22415,N_22173);
and U23862 (N_23862,N_22791,N_22330);
and U23863 (N_23863,N_22035,N_22821);
or U23864 (N_23864,N_22825,N_22858);
or U23865 (N_23865,N_22753,N_22745);
or U23866 (N_23866,N_22879,N_22108);
or U23867 (N_23867,N_22563,N_22846);
nand U23868 (N_23868,N_22352,N_22224);
nor U23869 (N_23869,N_22975,N_22213);
and U23870 (N_23870,N_22808,N_22262);
nor U23871 (N_23871,N_22776,N_22011);
and U23872 (N_23872,N_22134,N_22498);
nand U23873 (N_23873,N_22256,N_22505);
xor U23874 (N_23874,N_22543,N_22300);
nand U23875 (N_23875,N_22536,N_22280);
or U23876 (N_23876,N_22755,N_22686);
and U23877 (N_23877,N_22470,N_22687);
xor U23878 (N_23878,N_22819,N_22467);
nor U23879 (N_23879,N_22180,N_22062);
or U23880 (N_23880,N_22079,N_22820);
xor U23881 (N_23881,N_22488,N_22553);
nand U23882 (N_23882,N_22186,N_22244);
xor U23883 (N_23883,N_22812,N_22017);
and U23884 (N_23884,N_22865,N_22854);
nand U23885 (N_23885,N_22498,N_22489);
nor U23886 (N_23886,N_22025,N_22430);
nand U23887 (N_23887,N_22560,N_22093);
nand U23888 (N_23888,N_22193,N_22503);
nor U23889 (N_23889,N_22143,N_22811);
nor U23890 (N_23890,N_22269,N_22312);
nand U23891 (N_23891,N_22331,N_22302);
nor U23892 (N_23892,N_22688,N_22698);
nor U23893 (N_23893,N_22938,N_22878);
or U23894 (N_23894,N_22881,N_22257);
nor U23895 (N_23895,N_22118,N_22679);
xor U23896 (N_23896,N_22745,N_22351);
nor U23897 (N_23897,N_22087,N_22622);
and U23898 (N_23898,N_22773,N_22610);
nor U23899 (N_23899,N_22050,N_22060);
nand U23900 (N_23900,N_22139,N_22272);
nand U23901 (N_23901,N_22537,N_22490);
nand U23902 (N_23902,N_22563,N_22123);
or U23903 (N_23903,N_22946,N_22672);
nor U23904 (N_23904,N_22439,N_22357);
xor U23905 (N_23905,N_22654,N_22559);
nor U23906 (N_23906,N_22956,N_22600);
and U23907 (N_23907,N_22439,N_22938);
nand U23908 (N_23908,N_22955,N_22305);
or U23909 (N_23909,N_22381,N_22375);
or U23910 (N_23910,N_22263,N_22513);
nand U23911 (N_23911,N_22629,N_22196);
or U23912 (N_23912,N_22452,N_22724);
nand U23913 (N_23913,N_22710,N_22747);
and U23914 (N_23914,N_22063,N_22283);
xor U23915 (N_23915,N_22297,N_22748);
and U23916 (N_23916,N_22081,N_22266);
nor U23917 (N_23917,N_22577,N_22447);
xnor U23918 (N_23918,N_22624,N_22357);
or U23919 (N_23919,N_22418,N_22815);
or U23920 (N_23920,N_22719,N_22021);
and U23921 (N_23921,N_22524,N_22364);
xor U23922 (N_23922,N_22101,N_22368);
xor U23923 (N_23923,N_22094,N_22217);
or U23924 (N_23924,N_22226,N_22284);
and U23925 (N_23925,N_22889,N_22387);
and U23926 (N_23926,N_22134,N_22004);
nand U23927 (N_23927,N_22197,N_22580);
or U23928 (N_23928,N_22308,N_22602);
nor U23929 (N_23929,N_22219,N_22486);
nor U23930 (N_23930,N_22216,N_22646);
and U23931 (N_23931,N_22462,N_22653);
nor U23932 (N_23932,N_22271,N_22350);
or U23933 (N_23933,N_22682,N_22709);
and U23934 (N_23934,N_22005,N_22315);
or U23935 (N_23935,N_22587,N_22026);
xor U23936 (N_23936,N_22338,N_22320);
nor U23937 (N_23937,N_22216,N_22912);
xor U23938 (N_23938,N_22409,N_22122);
nor U23939 (N_23939,N_22620,N_22236);
xor U23940 (N_23940,N_22400,N_22582);
nor U23941 (N_23941,N_22984,N_22558);
or U23942 (N_23942,N_22745,N_22011);
and U23943 (N_23943,N_22792,N_22600);
and U23944 (N_23944,N_22707,N_22829);
nor U23945 (N_23945,N_22263,N_22407);
and U23946 (N_23946,N_22515,N_22333);
nand U23947 (N_23947,N_22091,N_22403);
xnor U23948 (N_23948,N_22309,N_22573);
and U23949 (N_23949,N_22978,N_22691);
or U23950 (N_23950,N_22176,N_22991);
nand U23951 (N_23951,N_22401,N_22402);
nand U23952 (N_23952,N_22544,N_22192);
xor U23953 (N_23953,N_22656,N_22128);
xnor U23954 (N_23954,N_22507,N_22426);
xnor U23955 (N_23955,N_22231,N_22639);
xor U23956 (N_23956,N_22585,N_22780);
or U23957 (N_23957,N_22855,N_22729);
nor U23958 (N_23958,N_22254,N_22436);
and U23959 (N_23959,N_22815,N_22704);
nand U23960 (N_23960,N_22645,N_22780);
or U23961 (N_23961,N_22575,N_22343);
and U23962 (N_23962,N_22664,N_22224);
nand U23963 (N_23963,N_22703,N_22656);
nand U23964 (N_23964,N_22957,N_22047);
or U23965 (N_23965,N_22875,N_22507);
and U23966 (N_23966,N_22164,N_22311);
nor U23967 (N_23967,N_22225,N_22340);
and U23968 (N_23968,N_22297,N_22831);
or U23969 (N_23969,N_22567,N_22676);
or U23970 (N_23970,N_22960,N_22821);
or U23971 (N_23971,N_22991,N_22184);
nor U23972 (N_23972,N_22483,N_22965);
and U23973 (N_23973,N_22185,N_22514);
or U23974 (N_23974,N_22099,N_22478);
xnor U23975 (N_23975,N_22594,N_22571);
or U23976 (N_23976,N_22693,N_22418);
and U23977 (N_23977,N_22898,N_22492);
xnor U23978 (N_23978,N_22512,N_22581);
and U23979 (N_23979,N_22129,N_22838);
or U23980 (N_23980,N_22376,N_22611);
xor U23981 (N_23981,N_22264,N_22226);
or U23982 (N_23982,N_22767,N_22765);
and U23983 (N_23983,N_22686,N_22160);
nand U23984 (N_23984,N_22485,N_22422);
and U23985 (N_23985,N_22866,N_22679);
xnor U23986 (N_23986,N_22354,N_22938);
and U23987 (N_23987,N_22155,N_22683);
xor U23988 (N_23988,N_22848,N_22696);
and U23989 (N_23989,N_22250,N_22981);
nand U23990 (N_23990,N_22097,N_22184);
xnor U23991 (N_23991,N_22839,N_22003);
and U23992 (N_23992,N_22774,N_22237);
nand U23993 (N_23993,N_22000,N_22047);
or U23994 (N_23994,N_22505,N_22671);
nor U23995 (N_23995,N_22397,N_22078);
xnor U23996 (N_23996,N_22395,N_22811);
and U23997 (N_23997,N_22164,N_22769);
nand U23998 (N_23998,N_22774,N_22752);
and U23999 (N_23999,N_22758,N_22614);
or U24000 (N_24000,N_23720,N_23646);
or U24001 (N_24001,N_23181,N_23619);
and U24002 (N_24002,N_23626,N_23403);
xor U24003 (N_24003,N_23744,N_23902);
nor U24004 (N_24004,N_23194,N_23889);
and U24005 (N_24005,N_23481,N_23593);
nand U24006 (N_24006,N_23662,N_23800);
and U24007 (N_24007,N_23964,N_23219);
and U24008 (N_24008,N_23732,N_23923);
xor U24009 (N_24009,N_23003,N_23274);
and U24010 (N_24010,N_23470,N_23095);
nor U24011 (N_24011,N_23221,N_23484);
nor U24012 (N_24012,N_23308,N_23913);
nor U24013 (N_24013,N_23021,N_23955);
or U24014 (N_24014,N_23010,N_23891);
and U24015 (N_24015,N_23556,N_23629);
xor U24016 (N_24016,N_23085,N_23642);
nor U24017 (N_24017,N_23271,N_23984);
nor U24018 (N_24018,N_23270,N_23353);
or U24019 (N_24019,N_23237,N_23075);
and U24020 (N_24020,N_23313,N_23376);
or U24021 (N_24021,N_23538,N_23536);
or U24022 (N_24022,N_23125,N_23974);
and U24023 (N_24023,N_23367,N_23290);
and U24024 (N_24024,N_23385,N_23548);
nor U24025 (N_24025,N_23321,N_23763);
or U24026 (N_24026,N_23760,N_23609);
nand U24027 (N_24027,N_23232,N_23083);
nand U24028 (N_24028,N_23413,N_23968);
nor U24029 (N_24029,N_23396,N_23129);
or U24030 (N_24030,N_23144,N_23530);
nor U24031 (N_24031,N_23192,N_23648);
nand U24032 (N_24032,N_23013,N_23643);
nand U24033 (N_24033,N_23424,N_23846);
and U24034 (N_24034,N_23722,N_23737);
xor U24035 (N_24035,N_23865,N_23289);
xnor U24036 (N_24036,N_23569,N_23005);
nand U24037 (N_24037,N_23517,N_23611);
nand U24038 (N_24038,N_23292,N_23751);
xor U24039 (N_24039,N_23475,N_23001);
or U24040 (N_24040,N_23717,N_23450);
xnor U24041 (N_24041,N_23836,N_23983);
or U24042 (N_24042,N_23068,N_23153);
and U24043 (N_24043,N_23358,N_23486);
and U24044 (N_24044,N_23528,N_23374);
xor U24045 (N_24045,N_23327,N_23146);
or U24046 (N_24046,N_23541,N_23465);
xnor U24047 (N_24047,N_23670,N_23186);
nor U24048 (N_24048,N_23698,N_23912);
and U24049 (N_24049,N_23254,N_23857);
and U24050 (N_24050,N_23847,N_23049);
or U24051 (N_24051,N_23755,N_23971);
nand U24052 (N_24052,N_23810,N_23595);
and U24053 (N_24053,N_23037,N_23754);
or U24054 (N_24054,N_23540,N_23750);
nor U24055 (N_24055,N_23918,N_23170);
and U24056 (N_24056,N_23561,N_23654);
and U24057 (N_24057,N_23208,N_23636);
nor U24058 (N_24058,N_23697,N_23317);
or U24059 (N_24059,N_23659,N_23600);
nand U24060 (N_24060,N_23565,N_23672);
and U24061 (N_24061,N_23684,N_23128);
and U24062 (N_24062,N_23514,N_23050);
and U24063 (N_24063,N_23917,N_23956);
xor U24064 (N_24064,N_23236,N_23265);
and U24065 (N_24065,N_23038,N_23507);
nand U24066 (N_24066,N_23625,N_23425);
nor U24067 (N_24067,N_23195,N_23411);
nand U24068 (N_24068,N_23390,N_23703);
and U24069 (N_24069,N_23036,N_23603);
nor U24070 (N_24070,N_23859,N_23069);
and U24071 (N_24071,N_23803,N_23577);
or U24072 (N_24072,N_23812,N_23771);
and U24073 (N_24073,N_23238,N_23903);
nor U24074 (N_24074,N_23849,N_23117);
or U24075 (N_24075,N_23513,N_23077);
nor U24076 (N_24076,N_23777,N_23942);
or U24077 (N_24077,N_23071,N_23597);
nand U24078 (N_24078,N_23025,N_23349);
or U24079 (N_24079,N_23925,N_23973);
nand U24080 (N_24080,N_23252,N_23305);
nand U24081 (N_24081,N_23651,N_23065);
nor U24082 (N_24082,N_23328,N_23985);
nor U24083 (N_24083,N_23915,N_23341);
nand U24084 (N_24084,N_23681,N_23734);
nor U24085 (N_24085,N_23899,N_23892);
or U24086 (N_24086,N_23993,N_23553);
or U24087 (N_24087,N_23512,N_23430);
or U24088 (N_24088,N_23306,N_23753);
or U24089 (N_24089,N_23897,N_23419);
nor U24090 (N_24090,N_23980,N_23620);
nor U24091 (N_24091,N_23216,N_23241);
xor U24092 (N_24092,N_23665,N_23420);
nor U24093 (N_24093,N_23024,N_23004);
nand U24094 (N_24094,N_23559,N_23570);
nor U24095 (N_24095,N_23933,N_23088);
and U24096 (N_24096,N_23579,N_23711);
nor U24097 (N_24097,N_23791,N_23310);
and U24098 (N_24098,N_23360,N_23158);
nand U24099 (N_24099,N_23335,N_23124);
or U24100 (N_24100,N_23275,N_23808);
nor U24101 (N_24101,N_23695,N_23299);
nand U24102 (N_24102,N_23961,N_23965);
or U24103 (N_24103,N_23231,N_23078);
and U24104 (N_24104,N_23279,N_23246);
or U24105 (N_24105,N_23458,N_23023);
nand U24106 (N_24106,N_23293,N_23802);
and U24107 (N_24107,N_23825,N_23444);
nor U24108 (N_24108,N_23463,N_23140);
or U24109 (N_24109,N_23161,N_23886);
xor U24110 (N_24110,N_23788,N_23362);
or U24111 (N_24111,N_23832,N_23082);
or U24112 (N_24112,N_23101,N_23446);
and U24113 (N_24113,N_23845,N_23368);
xor U24114 (N_24114,N_23340,N_23946);
and U24115 (N_24115,N_23172,N_23426);
and U24116 (N_24116,N_23028,N_23987);
nor U24117 (N_24117,N_23156,N_23029);
and U24118 (N_24118,N_23397,N_23945);
nand U24119 (N_24119,N_23989,N_23671);
xor U24120 (N_24120,N_23908,N_23322);
and U24121 (N_24121,N_23401,N_23584);
xnor U24122 (N_24122,N_23778,N_23007);
nand U24123 (N_24123,N_23949,N_23015);
or U24124 (N_24124,N_23572,N_23494);
and U24125 (N_24125,N_23690,N_23201);
or U24126 (N_24126,N_23014,N_23460);
or U24127 (N_24127,N_23476,N_23346);
xor U24128 (N_24128,N_23727,N_23418);
or U24129 (N_24129,N_23852,N_23647);
and U24130 (N_24130,N_23053,N_23392);
nand U24131 (N_24131,N_23728,N_23854);
nand U24132 (N_24132,N_23423,N_23157);
nand U24133 (N_24133,N_23377,N_23228);
and U24134 (N_24134,N_23045,N_23459);
nand U24135 (N_24135,N_23116,N_23137);
nand U24136 (N_24136,N_23519,N_23986);
xor U24137 (N_24137,N_23818,N_23482);
or U24138 (N_24138,N_23640,N_23834);
xor U24139 (N_24139,N_23704,N_23819);
and U24140 (N_24140,N_23009,N_23109);
nor U24141 (N_24141,N_23888,N_23355);
and U24142 (N_24142,N_23652,N_23780);
and U24143 (N_24143,N_23999,N_23248);
or U24144 (N_24144,N_23785,N_23474);
xor U24145 (N_24145,N_23537,N_23111);
or U24146 (N_24146,N_23667,N_23885);
nand U24147 (N_24147,N_23894,N_23781);
or U24148 (N_24148,N_23006,N_23615);
and U24149 (N_24149,N_23926,N_23747);
nand U24150 (N_24150,N_23757,N_23469);
nor U24151 (N_24151,N_23199,N_23693);
and U24152 (N_24152,N_23872,N_23590);
nor U24153 (N_24153,N_23239,N_23884);
xnor U24154 (N_24154,N_23844,N_23505);
or U24155 (N_24155,N_23381,N_23227);
nand U24156 (N_24156,N_23303,N_23539);
nand U24157 (N_24157,N_23914,N_23408);
or U24158 (N_24158,N_23841,N_23831);
and U24159 (N_24159,N_23745,N_23414);
xnor U24160 (N_24160,N_23765,N_23998);
nor U24161 (N_24161,N_23243,N_23784);
and U24162 (N_24162,N_23749,N_23415);
and U24163 (N_24163,N_23268,N_23256);
and U24164 (N_24164,N_23323,N_23574);
nand U24165 (N_24165,N_23938,N_23516);
and U24166 (N_24166,N_23566,N_23527);
xnor U24167 (N_24167,N_23633,N_23017);
and U24168 (N_24168,N_23213,N_23115);
nand U24169 (N_24169,N_23466,N_23969);
or U24170 (N_24170,N_23438,N_23104);
nand U24171 (N_24171,N_23188,N_23978);
xnor U24172 (N_24172,N_23668,N_23073);
nand U24173 (N_24173,N_23225,N_23016);
and U24174 (N_24174,N_23543,N_23108);
or U24175 (N_24175,N_23931,N_23046);
and U24176 (N_24176,N_23582,N_23361);
xor U24177 (N_24177,N_23097,N_23692);
nor U24178 (N_24178,N_23976,N_23112);
nand U24179 (N_24179,N_23247,N_23002);
nand U24180 (N_24180,N_23373,N_23165);
xor U24181 (N_24181,N_23162,N_23389);
or U24182 (N_24182,N_23276,N_23394);
and U24183 (N_24183,N_23176,N_23296);
nor U24184 (N_24184,N_23131,N_23730);
nand U24185 (N_24185,N_23487,N_23916);
xor U24186 (N_24186,N_23257,N_23554);
and U24187 (N_24187,N_23145,N_23316);
or U24188 (N_24188,N_23877,N_23179);
and U24189 (N_24189,N_23649,N_23178);
xor U24190 (N_24190,N_23525,N_23526);
nand U24191 (N_24191,N_23019,N_23545);
nand U24192 (N_24192,N_23655,N_23712);
and U24193 (N_24193,N_23027,N_23233);
nand U24194 (N_24194,N_23200,N_23359);
and U24195 (N_24195,N_23325,N_23052);
and U24196 (N_24196,N_23988,N_23963);
xor U24197 (N_24197,N_23868,N_23714);
xor U24198 (N_24198,N_23850,N_23990);
nor U24199 (N_24199,N_23521,N_23645);
nor U24200 (N_24200,N_23550,N_23092);
xor U24201 (N_24201,N_23434,N_23848);
and U24202 (N_24202,N_23365,N_23467);
nand U24203 (N_24203,N_23705,N_23713);
nor U24204 (N_24204,N_23863,N_23607);
or U24205 (N_24205,N_23473,N_23464);
and U24206 (N_24206,N_23827,N_23683);
nand U24207 (N_24207,N_23842,N_23503);
nor U24208 (N_24208,N_23206,N_23410);
xnor U24209 (N_24209,N_23534,N_23860);
nand U24210 (N_24210,N_23601,N_23947);
and U24211 (N_24211,N_23710,N_23409);
nor U24212 (N_24212,N_23008,N_23960);
and U24213 (N_24213,N_23442,N_23743);
nor U24214 (N_24214,N_23682,N_23518);
nor U24215 (N_24215,N_23687,N_23339);
nand U24216 (N_24216,N_23996,N_23840);
xor U24217 (N_24217,N_23816,N_23883);
xnor U24218 (N_24218,N_23972,N_23921);
nand U24219 (N_24219,N_23059,N_23149);
xnor U24220 (N_24220,N_23447,N_23063);
or U24221 (N_24221,N_23515,N_23813);
and U24222 (N_24222,N_23291,N_23240);
or U24223 (N_24223,N_23634,N_23608);
nand U24224 (N_24224,N_23853,N_23679);
nand U24225 (N_24225,N_23560,N_23220);
and U24226 (N_24226,N_23106,N_23074);
xnor U24227 (N_24227,N_23624,N_23524);
xor U24228 (N_24228,N_23187,N_23948);
and U24229 (N_24229,N_23522,N_23372);
or U24230 (N_24230,N_23344,N_23269);
xnor U24231 (N_24231,N_23040,N_23455);
or U24232 (N_24232,N_23631,N_23263);
or U24233 (N_24233,N_23838,N_23740);
nor U24234 (N_24234,N_23490,N_23927);
xnor U24235 (N_24235,N_23141,N_23782);
xor U24236 (N_24236,N_23301,N_23384);
nor U24237 (N_24237,N_23242,N_23953);
nand U24238 (N_24238,N_23431,N_23719);
xor U24239 (N_24239,N_23520,N_23315);
xor U24240 (N_24240,N_23930,N_23641);
nor U24241 (N_24241,N_23991,N_23909);
xnor U24242 (N_24242,N_23779,N_23664);
and U24243 (N_24243,N_23542,N_23614);
nor U24244 (N_24244,N_23571,N_23084);
and U24245 (N_24245,N_23443,N_23087);
nor U24246 (N_24246,N_23311,N_23471);
nand U24247 (N_24247,N_23992,N_23715);
nand U24248 (N_24248,N_23689,N_23066);
xor U24249 (N_24249,N_23851,N_23307);
xor U24250 (N_24250,N_23770,N_23793);
and U24251 (N_24251,N_23900,N_23148);
and U24252 (N_24252,N_23298,N_23499);
or U24253 (N_24253,N_23427,N_23523);
and U24254 (N_24254,N_23576,N_23058);
and U24255 (N_24255,N_23922,N_23214);
nor U24256 (N_24256,N_23907,N_23875);
and U24257 (N_24257,N_23962,N_23606);
or U24258 (N_24258,N_23429,N_23485);
nand U24259 (N_24259,N_23034,N_23511);
nor U24260 (N_24260,N_23555,N_23653);
or U24261 (N_24261,N_23970,N_23501);
nand U24262 (N_24262,N_23267,N_23762);
nor U24263 (N_24263,N_23508,N_23591);
xor U24264 (N_24264,N_23336,N_23107);
nor U24265 (N_24265,N_23628,N_23099);
nand U24266 (N_24266,N_23635,N_23975);
nand U24267 (N_24267,N_23399,N_23959);
or U24268 (N_24268,N_23578,N_23596);
nor U24269 (N_24269,N_23580,N_23472);
and U24270 (N_24270,N_23212,N_23086);
nor U24271 (N_24271,N_23563,N_23613);
nand U24272 (N_24272,N_23379,N_23795);
and U24273 (N_24273,N_23935,N_23363);
xor U24274 (N_24274,N_23799,N_23205);
nand U24275 (N_24275,N_23309,N_23378);
nand U24276 (N_24276,N_23433,N_23869);
nor U24277 (N_24277,N_23076,N_23929);
xnor U24278 (N_24278,N_23169,N_23792);
nor U24279 (N_24279,N_23143,N_23588);
xor U24280 (N_24280,N_23405,N_23500);
and U24281 (N_24281,N_23958,N_23185);
or U24282 (N_24282,N_23746,N_23604);
nor U24283 (N_24283,N_23796,N_23742);
nor U24284 (N_24284,N_23650,N_23417);
or U24285 (N_24285,N_23531,N_23943);
nand U24286 (N_24286,N_23167,N_23822);
and U24287 (N_24287,N_23637,N_23491);
nand U24288 (N_24288,N_23839,N_23197);
nand U24289 (N_24289,N_23318,N_23766);
nand U24290 (N_24290,N_23830,N_23151);
and U24291 (N_24291,N_23977,N_23294);
nor U24292 (N_24292,N_23051,N_23870);
nand U24293 (N_24293,N_23127,N_23686);
xnor U24294 (N_24294,N_23400,N_23030);
or U24295 (N_24295,N_23627,N_23056);
nand U24296 (N_24296,N_23067,N_23954);
or U24297 (N_24297,N_23031,N_23495);
nand U24298 (N_24298,N_23333,N_23529);
nand U24299 (N_24299,N_23393,N_23215);
and U24300 (N_24300,N_23618,N_23044);
nor U24301 (N_24301,N_23549,N_23057);
xnor U24302 (N_24302,N_23168,N_23700);
xor U24303 (N_24303,N_23807,N_23906);
nand U24304 (N_24304,N_23787,N_23436);
nor U24305 (N_24305,N_23552,N_23982);
nand U24306 (N_24306,N_23422,N_23739);
nor U24307 (N_24307,N_23901,N_23300);
nor U24308 (N_24308,N_23312,N_23375);
nor U24309 (N_24309,N_23055,N_23801);
xnor U24310 (N_24310,N_23264,N_23941);
xnor U24311 (N_24311,N_23814,N_23272);
nor U24312 (N_24312,N_23966,N_23121);
or U24313 (N_24313,N_23786,N_23895);
xnor U24314 (N_24314,N_23504,N_23533);
nor U24315 (N_24315,N_23391,N_23478);
nor U24316 (N_24316,N_23454,N_23725);
or U24317 (N_24317,N_23000,N_23716);
nor U24318 (N_24318,N_23890,N_23110);
nand U24319 (N_24319,N_23022,N_23026);
xnor U24320 (N_24320,N_23183,N_23229);
nand U24321 (N_24321,N_23196,N_23326);
xnor U24322 (N_24322,N_23871,N_23171);
and U24323 (N_24323,N_23691,N_23159);
or U24324 (N_24324,N_23398,N_23492);
nor U24325 (N_24325,N_23677,N_23674);
nand U24326 (N_24326,N_23882,N_23821);
nand U24327 (N_24327,N_23147,N_23567);
xor U24328 (N_24328,N_23283,N_23581);
or U24329 (N_24329,N_23448,N_23119);
nand U24330 (N_24330,N_23610,N_23456);
or U24331 (N_24331,N_23366,N_23062);
and U24332 (N_24332,N_23284,N_23054);
nor U24333 (N_24333,N_23558,N_23380);
and U24334 (N_24334,N_23630,N_23598);
nand U24335 (N_24335,N_23773,N_23338);
and U24336 (N_24336,N_23421,N_23139);
xor U24337 (N_24337,N_23605,N_23287);
nand U24338 (N_24338,N_23136,N_23286);
or U24339 (N_24339,N_23035,N_23250);
xor U24340 (N_24340,N_23295,N_23061);
xnor U24341 (N_24341,N_23297,N_23936);
nor U24342 (N_24342,N_23060,N_23709);
nor U24343 (N_24343,N_23018,N_23130);
nand U24344 (N_24344,N_23189,N_23707);
or U24345 (N_24345,N_23488,N_23102);
nor U24346 (N_24346,N_23497,N_23881);
nand U24347 (N_24347,N_23680,N_23950);
xor U24348 (N_24348,N_23879,N_23209);
xor U24349 (N_24349,N_23480,N_23723);
nor U24350 (N_24350,N_23395,N_23873);
or U24351 (N_24351,N_23612,N_23688);
or U24352 (N_24352,N_23160,N_23856);
xor U24353 (N_24353,N_23190,N_23126);
or U24354 (N_24354,N_23132,N_23449);
or U24355 (N_24355,N_23828,N_23661);
xor U24356 (N_24356,N_23741,N_23352);
or U24357 (N_24357,N_23940,N_23226);
and U24358 (N_24358,N_23660,N_23564);
xnor U24359 (N_24359,N_23211,N_23676);
xor U24360 (N_24360,N_23253,N_23783);
nor U24361 (N_24361,N_23461,N_23331);
xnor U24362 (N_24362,N_23357,N_23218);
or U24363 (N_24363,N_23994,N_23404);
nand U24364 (N_24364,N_23833,N_23920);
and U24365 (N_24365,N_23244,N_23383);
xor U24366 (N_24366,N_23382,N_23817);
or U24367 (N_24367,N_23462,N_23748);
or U24368 (N_24368,N_23724,N_23798);
nand U24369 (N_24369,N_23428,N_23319);
nand U24370 (N_24370,N_23509,N_23020);
and U24371 (N_24371,N_23314,N_23334);
or U24372 (N_24372,N_23789,N_23324);
nand U24373 (N_24373,N_23806,N_23193);
and U24374 (N_24374,N_23911,N_23811);
or U24375 (N_24375,N_23867,N_23251);
nor U24376 (N_24376,N_23592,N_23175);
xor U24377 (N_24377,N_23893,N_23412);
nand U24378 (N_24378,N_23120,N_23735);
nor U24379 (N_24379,N_23502,N_23769);
xor U24380 (N_24380,N_23098,N_23752);
and U24381 (N_24381,N_23135,N_23804);
nor U24382 (N_24382,N_23342,N_23685);
nand U24383 (N_24383,N_23445,N_23721);
or U24384 (N_24384,N_23862,N_23280);
or U24385 (N_24385,N_23876,N_23387);
xor U24386 (N_24386,N_23775,N_23261);
nand U24387 (N_24387,N_23207,N_23731);
and U24388 (N_24388,N_23198,N_23100);
nand U24389 (N_24389,N_23369,N_23350);
nor U24390 (N_24390,N_23090,N_23043);
and U24391 (N_24391,N_23623,N_23656);
nand U24392 (N_24392,N_23809,N_23154);
nand U24393 (N_24393,N_23837,N_23259);
xor U24394 (N_24394,N_23493,N_23774);
and U24395 (N_24395,N_23439,N_23096);
nand U24396 (N_24396,N_23032,N_23701);
nand U24397 (N_24397,N_23416,N_23794);
nor U24398 (N_24398,N_23105,N_23451);
xnor U24399 (N_24399,N_23639,N_23235);
xnor U24400 (N_24400,N_23118,N_23937);
xnor U24401 (N_24401,N_23388,N_23138);
nand U24402 (N_24402,N_23222,N_23278);
and U24403 (N_24403,N_23266,N_23166);
and U24404 (N_24404,N_23164,N_23210);
xnor U24405 (N_24405,N_23573,N_23173);
xor U24406 (N_24406,N_23657,N_23288);
and U24407 (N_24407,N_23356,N_23616);
nor U24408 (N_24408,N_23928,N_23047);
xnor U24409 (N_24409,N_23048,N_23562);
nor U24410 (N_24410,N_23858,N_23260);
nand U24411 (N_24411,N_23934,N_23557);
or U24412 (N_24412,N_23878,N_23738);
xor U24413 (N_24413,N_23669,N_23820);
or U24414 (N_24414,N_23012,N_23432);
or U24415 (N_24415,N_23435,N_23155);
xor U24416 (N_24416,N_23262,N_23726);
xnor U24417 (N_24417,N_23594,N_23437);
xor U24418 (N_24418,N_23457,N_23079);
nand U24419 (N_24419,N_23924,N_23997);
or U24420 (N_24420,N_23952,N_23330);
and U24421 (N_24421,N_23406,N_23632);
and U24422 (N_24422,N_23245,N_23758);
nand U24423 (N_24423,N_23042,N_23150);
nand U24424 (N_24424,N_23733,N_23932);
xnor U24425 (N_24425,N_23658,N_23904);
nor U24426 (N_24426,N_23407,N_23638);
nor U24427 (N_24427,N_23905,N_23202);
nand U24428 (N_24428,N_23332,N_23113);
and U24429 (N_24429,N_23772,N_23386);
nor U24430 (N_24430,N_23824,N_23535);
nor U24431 (N_24431,N_23910,N_23320);
xor U24432 (N_24432,N_23134,N_23644);
nand U24433 (N_24433,N_23094,N_23223);
and U24434 (N_24434,N_23547,N_23343);
and U24435 (N_24435,N_23203,N_23544);
and U24436 (N_24436,N_23694,N_23699);
or U24437 (N_24437,N_23621,N_23347);
nor U24438 (N_24438,N_23285,N_23337);
xor U24439 (N_24439,N_23599,N_23696);
and U24440 (N_24440,N_23957,N_23761);
or U24441 (N_24441,N_23759,N_23896);
nor U24442 (N_24442,N_23093,N_23981);
or U24443 (N_24443,N_23589,N_23979);
nand U24444 (N_24444,N_23453,N_23675);
nand U24445 (N_24445,N_23234,N_23114);
nor U24446 (N_24446,N_23510,N_23826);
and U24447 (N_24447,N_23282,N_23708);
nand U24448 (N_24448,N_23866,N_23551);
nor U24449 (N_24449,N_23776,N_23370);
and U24450 (N_24450,N_23177,N_23678);
xor U24451 (N_24451,N_23152,N_23142);
or U24452 (N_24452,N_23874,N_23829);
and U24453 (N_24453,N_23354,N_23919);
nand U24454 (N_24454,N_23255,N_23835);
and U24455 (N_24455,N_23258,N_23191);
nand U24456 (N_24456,N_23702,N_23756);
nor U24457 (N_24457,N_23163,N_23249);
xnor U24458 (N_24458,N_23224,N_23805);
xnor U24459 (N_24459,N_23568,N_23583);
xnor U24460 (N_24460,N_23184,N_23204);
and U24461 (N_24461,N_23887,N_23033);
and U24462 (N_24462,N_23182,N_23452);
and U24463 (N_24463,N_23304,N_23217);
or U24464 (N_24464,N_23483,N_23764);
xnor U24465 (N_24465,N_23351,N_23864);
nand U24466 (N_24466,N_23587,N_23174);
nand U24467 (N_24467,N_23348,N_23586);
xnor U24468 (N_24468,N_23180,N_23673);
or U24469 (N_24469,N_23736,N_23546);
xor U24470 (N_24470,N_23855,N_23080);
or U24471 (N_24471,N_23277,N_23441);
nor U24472 (N_24472,N_23402,N_23281);
nand U24473 (N_24473,N_23122,N_23371);
nor U24474 (N_24474,N_23081,N_23498);
or U24475 (N_24475,N_23880,N_23496);
nand U24476 (N_24476,N_23995,N_23345);
and U24477 (N_24477,N_23666,N_23364);
nor U24478 (N_24478,N_23039,N_23230);
nor U24479 (N_24479,N_23329,N_23532);
and U24480 (N_24480,N_23622,N_23091);
nand U24481 (N_24481,N_23011,N_23072);
or U24482 (N_24482,N_23706,N_23602);
and U24483 (N_24483,N_23898,N_23575);
xnor U24484 (N_24484,N_23861,N_23440);
xnor U24485 (N_24485,N_23790,N_23489);
nand U24486 (N_24486,N_23479,N_23729);
xor U24487 (N_24487,N_23815,N_23939);
or U24488 (N_24488,N_23843,N_23951);
or U24489 (N_24489,N_23617,N_23273);
xnor U24490 (N_24490,N_23768,N_23967);
and U24491 (N_24491,N_23585,N_23797);
or U24492 (N_24492,N_23767,N_23133);
xnor U24493 (N_24493,N_23302,N_23944);
nor U24494 (N_24494,N_23506,N_23103);
xnor U24495 (N_24495,N_23123,N_23089);
xnor U24496 (N_24496,N_23477,N_23663);
or U24497 (N_24497,N_23468,N_23823);
xor U24498 (N_24498,N_23070,N_23718);
nand U24499 (N_24499,N_23041,N_23064);
nor U24500 (N_24500,N_23233,N_23250);
xor U24501 (N_24501,N_23721,N_23701);
and U24502 (N_24502,N_23147,N_23204);
and U24503 (N_24503,N_23958,N_23249);
or U24504 (N_24504,N_23562,N_23490);
nor U24505 (N_24505,N_23705,N_23581);
nor U24506 (N_24506,N_23395,N_23489);
or U24507 (N_24507,N_23734,N_23750);
or U24508 (N_24508,N_23728,N_23410);
or U24509 (N_24509,N_23772,N_23140);
or U24510 (N_24510,N_23191,N_23814);
or U24511 (N_24511,N_23610,N_23271);
nand U24512 (N_24512,N_23832,N_23598);
xor U24513 (N_24513,N_23957,N_23010);
nor U24514 (N_24514,N_23604,N_23703);
nand U24515 (N_24515,N_23736,N_23354);
nor U24516 (N_24516,N_23151,N_23120);
nand U24517 (N_24517,N_23214,N_23655);
xnor U24518 (N_24518,N_23687,N_23863);
nor U24519 (N_24519,N_23485,N_23137);
xnor U24520 (N_24520,N_23327,N_23650);
nor U24521 (N_24521,N_23502,N_23938);
xnor U24522 (N_24522,N_23701,N_23461);
nand U24523 (N_24523,N_23648,N_23834);
and U24524 (N_24524,N_23525,N_23861);
and U24525 (N_24525,N_23960,N_23763);
nor U24526 (N_24526,N_23568,N_23220);
xor U24527 (N_24527,N_23378,N_23026);
nor U24528 (N_24528,N_23959,N_23966);
xor U24529 (N_24529,N_23471,N_23602);
nor U24530 (N_24530,N_23460,N_23599);
nor U24531 (N_24531,N_23917,N_23003);
or U24532 (N_24532,N_23479,N_23970);
and U24533 (N_24533,N_23975,N_23386);
and U24534 (N_24534,N_23677,N_23778);
or U24535 (N_24535,N_23677,N_23381);
and U24536 (N_24536,N_23895,N_23371);
and U24537 (N_24537,N_23348,N_23373);
or U24538 (N_24538,N_23247,N_23113);
nor U24539 (N_24539,N_23094,N_23104);
or U24540 (N_24540,N_23022,N_23391);
or U24541 (N_24541,N_23044,N_23637);
nor U24542 (N_24542,N_23290,N_23236);
xnor U24543 (N_24543,N_23817,N_23332);
or U24544 (N_24544,N_23362,N_23346);
nand U24545 (N_24545,N_23345,N_23401);
xnor U24546 (N_24546,N_23926,N_23464);
xor U24547 (N_24547,N_23215,N_23989);
nor U24548 (N_24548,N_23782,N_23472);
nand U24549 (N_24549,N_23431,N_23352);
xor U24550 (N_24550,N_23247,N_23107);
nand U24551 (N_24551,N_23243,N_23218);
or U24552 (N_24552,N_23392,N_23442);
and U24553 (N_24553,N_23037,N_23926);
and U24554 (N_24554,N_23064,N_23328);
nand U24555 (N_24555,N_23087,N_23469);
xnor U24556 (N_24556,N_23004,N_23960);
nand U24557 (N_24557,N_23452,N_23722);
or U24558 (N_24558,N_23172,N_23372);
nand U24559 (N_24559,N_23177,N_23072);
nor U24560 (N_24560,N_23894,N_23763);
nand U24561 (N_24561,N_23820,N_23589);
and U24562 (N_24562,N_23948,N_23132);
or U24563 (N_24563,N_23638,N_23525);
and U24564 (N_24564,N_23377,N_23583);
nand U24565 (N_24565,N_23403,N_23670);
and U24566 (N_24566,N_23686,N_23353);
nand U24567 (N_24567,N_23488,N_23351);
xor U24568 (N_24568,N_23572,N_23074);
xor U24569 (N_24569,N_23226,N_23044);
xnor U24570 (N_24570,N_23956,N_23121);
or U24571 (N_24571,N_23134,N_23570);
nor U24572 (N_24572,N_23446,N_23194);
or U24573 (N_24573,N_23618,N_23553);
or U24574 (N_24574,N_23564,N_23844);
and U24575 (N_24575,N_23702,N_23434);
and U24576 (N_24576,N_23173,N_23141);
and U24577 (N_24577,N_23904,N_23074);
xor U24578 (N_24578,N_23321,N_23898);
nand U24579 (N_24579,N_23431,N_23577);
nand U24580 (N_24580,N_23265,N_23218);
xor U24581 (N_24581,N_23661,N_23612);
nor U24582 (N_24582,N_23884,N_23597);
and U24583 (N_24583,N_23888,N_23220);
xnor U24584 (N_24584,N_23895,N_23555);
nand U24585 (N_24585,N_23610,N_23651);
nor U24586 (N_24586,N_23287,N_23368);
or U24587 (N_24587,N_23371,N_23834);
or U24588 (N_24588,N_23208,N_23213);
nor U24589 (N_24589,N_23106,N_23075);
nand U24590 (N_24590,N_23238,N_23446);
and U24591 (N_24591,N_23509,N_23309);
xor U24592 (N_24592,N_23679,N_23660);
or U24593 (N_24593,N_23108,N_23604);
nor U24594 (N_24594,N_23097,N_23648);
xor U24595 (N_24595,N_23609,N_23325);
or U24596 (N_24596,N_23978,N_23397);
or U24597 (N_24597,N_23498,N_23316);
and U24598 (N_24598,N_23069,N_23180);
nand U24599 (N_24599,N_23942,N_23444);
xor U24600 (N_24600,N_23780,N_23800);
and U24601 (N_24601,N_23021,N_23418);
and U24602 (N_24602,N_23996,N_23977);
or U24603 (N_24603,N_23433,N_23387);
and U24604 (N_24604,N_23759,N_23505);
xor U24605 (N_24605,N_23448,N_23744);
xor U24606 (N_24606,N_23333,N_23898);
nor U24607 (N_24607,N_23194,N_23006);
xor U24608 (N_24608,N_23743,N_23911);
and U24609 (N_24609,N_23551,N_23397);
nor U24610 (N_24610,N_23120,N_23032);
nand U24611 (N_24611,N_23511,N_23987);
xor U24612 (N_24612,N_23763,N_23783);
and U24613 (N_24613,N_23622,N_23600);
xnor U24614 (N_24614,N_23349,N_23487);
nor U24615 (N_24615,N_23849,N_23225);
nand U24616 (N_24616,N_23002,N_23960);
nor U24617 (N_24617,N_23301,N_23987);
nor U24618 (N_24618,N_23273,N_23934);
and U24619 (N_24619,N_23579,N_23580);
or U24620 (N_24620,N_23254,N_23718);
and U24621 (N_24621,N_23539,N_23448);
or U24622 (N_24622,N_23954,N_23009);
xnor U24623 (N_24623,N_23413,N_23525);
or U24624 (N_24624,N_23282,N_23679);
nand U24625 (N_24625,N_23690,N_23967);
nand U24626 (N_24626,N_23428,N_23194);
xor U24627 (N_24627,N_23262,N_23427);
and U24628 (N_24628,N_23909,N_23823);
and U24629 (N_24629,N_23612,N_23408);
nand U24630 (N_24630,N_23212,N_23272);
and U24631 (N_24631,N_23813,N_23236);
nand U24632 (N_24632,N_23673,N_23277);
nor U24633 (N_24633,N_23351,N_23411);
or U24634 (N_24634,N_23809,N_23182);
or U24635 (N_24635,N_23732,N_23012);
and U24636 (N_24636,N_23969,N_23427);
nand U24637 (N_24637,N_23026,N_23994);
or U24638 (N_24638,N_23191,N_23782);
xor U24639 (N_24639,N_23629,N_23097);
and U24640 (N_24640,N_23336,N_23799);
nor U24641 (N_24641,N_23995,N_23964);
nor U24642 (N_24642,N_23065,N_23376);
or U24643 (N_24643,N_23370,N_23028);
nor U24644 (N_24644,N_23759,N_23466);
or U24645 (N_24645,N_23008,N_23727);
nand U24646 (N_24646,N_23613,N_23459);
or U24647 (N_24647,N_23861,N_23445);
and U24648 (N_24648,N_23559,N_23633);
nand U24649 (N_24649,N_23945,N_23959);
and U24650 (N_24650,N_23666,N_23757);
and U24651 (N_24651,N_23892,N_23443);
nor U24652 (N_24652,N_23668,N_23378);
nand U24653 (N_24653,N_23075,N_23495);
xnor U24654 (N_24654,N_23366,N_23386);
or U24655 (N_24655,N_23556,N_23246);
nor U24656 (N_24656,N_23500,N_23476);
and U24657 (N_24657,N_23116,N_23901);
nor U24658 (N_24658,N_23399,N_23679);
xor U24659 (N_24659,N_23286,N_23934);
nand U24660 (N_24660,N_23055,N_23423);
xor U24661 (N_24661,N_23596,N_23355);
nand U24662 (N_24662,N_23383,N_23864);
nor U24663 (N_24663,N_23600,N_23349);
nand U24664 (N_24664,N_23953,N_23189);
xnor U24665 (N_24665,N_23098,N_23649);
or U24666 (N_24666,N_23249,N_23101);
nand U24667 (N_24667,N_23347,N_23350);
xor U24668 (N_24668,N_23353,N_23688);
xor U24669 (N_24669,N_23005,N_23824);
nand U24670 (N_24670,N_23626,N_23558);
and U24671 (N_24671,N_23093,N_23102);
or U24672 (N_24672,N_23666,N_23570);
and U24673 (N_24673,N_23001,N_23212);
or U24674 (N_24674,N_23225,N_23820);
or U24675 (N_24675,N_23590,N_23294);
nor U24676 (N_24676,N_23971,N_23741);
xor U24677 (N_24677,N_23062,N_23369);
or U24678 (N_24678,N_23277,N_23256);
xor U24679 (N_24679,N_23529,N_23763);
and U24680 (N_24680,N_23870,N_23168);
and U24681 (N_24681,N_23614,N_23705);
or U24682 (N_24682,N_23116,N_23919);
xor U24683 (N_24683,N_23424,N_23062);
or U24684 (N_24684,N_23141,N_23435);
and U24685 (N_24685,N_23278,N_23695);
and U24686 (N_24686,N_23896,N_23304);
nand U24687 (N_24687,N_23607,N_23762);
nand U24688 (N_24688,N_23201,N_23841);
nor U24689 (N_24689,N_23851,N_23775);
or U24690 (N_24690,N_23111,N_23008);
or U24691 (N_24691,N_23533,N_23765);
xnor U24692 (N_24692,N_23793,N_23378);
nand U24693 (N_24693,N_23127,N_23007);
xnor U24694 (N_24694,N_23289,N_23702);
xor U24695 (N_24695,N_23971,N_23802);
or U24696 (N_24696,N_23121,N_23475);
nor U24697 (N_24697,N_23996,N_23871);
nor U24698 (N_24698,N_23790,N_23969);
xor U24699 (N_24699,N_23937,N_23710);
or U24700 (N_24700,N_23686,N_23890);
xor U24701 (N_24701,N_23184,N_23725);
or U24702 (N_24702,N_23221,N_23429);
nor U24703 (N_24703,N_23879,N_23246);
and U24704 (N_24704,N_23051,N_23936);
nand U24705 (N_24705,N_23929,N_23552);
or U24706 (N_24706,N_23534,N_23712);
and U24707 (N_24707,N_23728,N_23165);
nor U24708 (N_24708,N_23869,N_23714);
and U24709 (N_24709,N_23441,N_23115);
and U24710 (N_24710,N_23965,N_23329);
nor U24711 (N_24711,N_23799,N_23404);
and U24712 (N_24712,N_23235,N_23565);
and U24713 (N_24713,N_23379,N_23757);
xor U24714 (N_24714,N_23423,N_23675);
nor U24715 (N_24715,N_23010,N_23988);
nor U24716 (N_24716,N_23620,N_23330);
xor U24717 (N_24717,N_23770,N_23150);
or U24718 (N_24718,N_23851,N_23610);
nor U24719 (N_24719,N_23879,N_23420);
nand U24720 (N_24720,N_23717,N_23915);
nand U24721 (N_24721,N_23447,N_23829);
or U24722 (N_24722,N_23053,N_23746);
xor U24723 (N_24723,N_23961,N_23432);
or U24724 (N_24724,N_23265,N_23580);
nor U24725 (N_24725,N_23684,N_23544);
and U24726 (N_24726,N_23443,N_23042);
nor U24727 (N_24727,N_23207,N_23384);
and U24728 (N_24728,N_23975,N_23877);
or U24729 (N_24729,N_23298,N_23780);
xor U24730 (N_24730,N_23103,N_23689);
nor U24731 (N_24731,N_23549,N_23075);
or U24732 (N_24732,N_23480,N_23638);
nand U24733 (N_24733,N_23421,N_23591);
and U24734 (N_24734,N_23580,N_23805);
and U24735 (N_24735,N_23437,N_23468);
nand U24736 (N_24736,N_23090,N_23514);
and U24737 (N_24737,N_23966,N_23829);
nor U24738 (N_24738,N_23801,N_23383);
and U24739 (N_24739,N_23719,N_23419);
or U24740 (N_24740,N_23908,N_23691);
or U24741 (N_24741,N_23522,N_23445);
and U24742 (N_24742,N_23470,N_23761);
xor U24743 (N_24743,N_23064,N_23312);
and U24744 (N_24744,N_23664,N_23743);
xnor U24745 (N_24745,N_23406,N_23150);
and U24746 (N_24746,N_23264,N_23488);
or U24747 (N_24747,N_23882,N_23873);
nand U24748 (N_24748,N_23505,N_23068);
xor U24749 (N_24749,N_23209,N_23251);
nor U24750 (N_24750,N_23239,N_23332);
xor U24751 (N_24751,N_23205,N_23095);
nor U24752 (N_24752,N_23917,N_23277);
or U24753 (N_24753,N_23971,N_23351);
nand U24754 (N_24754,N_23279,N_23425);
xor U24755 (N_24755,N_23556,N_23325);
and U24756 (N_24756,N_23313,N_23734);
nand U24757 (N_24757,N_23844,N_23545);
nand U24758 (N_24758,N_23528,N_23632);
or U24759 (N_24759,N_23771,N_23986);
nor U24760 (N_24760,N_23386,N_23294);
or U24761 (N_24761,N_23684,N_23541);
nor U24762 (N_24762,N_23856,N_23385);
nor U24763 (N_24763,N_23191,N_23035);
nand U24764 (N_24764,N_23310,N_23368);
nand U24765 (N_24765,N_23957,N_23926);
nor U24766 (N_24766,N_23806,N_23259);
or U24767 (N_24767,N_23205,N_23971);
nand U24768 (N_24768,N_23992,N_23758);
and U24769 (N_24769,N_23370,N_23892);
and U24770 (N_24770,N_23455,N_23338);
nor U24771 (N_24771,N_23517,N_23652);
nand U24772 (N_24772,N_23436,N_23113);
xor U24773 (N_24773,N_23655,N_23348);
nand U24774 (N_24774,N_23084,N_23809);
and U24775 (N_24775,N_23028,N_23289);
xnor U24776 (N_24776,N_23552,N_23082);
nand U24777 (N_24777,N_23952,N_23740);
and U24778 (N_24778,N_23925,N_23321);
nand U24779 (N_24779,N_23287,N_23608);
nor U24780 (N_24780,N_23842,N_23908);
nor U24781 (N_24781,N_23660,N_23293);
nand U24782 (N_24782,N_23344,N_23056);
xnor U24783 (N_24783,N_23329,N_23401);
nand U24784 (N_24784,N_23523,N_23484);
nor U24785 (N_24785,N_23939,N_23916);
or U24786 (N_24786,N_23025,N_23960);
xnor U24787 (N_24787,N_23702,N_23778);
xnor U24788 (N_24788,N_23018,N_23864);
nor U24789 (N_24789,N_23768,N_23939);
and U24790 (N_24790,N_23950,N_23566);
or U24791 (N_24791,N_23032,N_23704);
nor U24792 (N_24792,N_23109,N_23943);
xor U24793 (N_24793,N_23923,N_23801);
nor U24794 (N_24794,N_23635,N_23285);
nor U24795 (N_24795,N_23686,N_23794);
xor U24796 (N_24796,N_23623,N_23213);
or U24797 (N_24797,N_23389,N_23219);
nand U24798 (N_24798,N_23723,N_23376);
nor U24799 (N_24799,N_23301,N_23426);
nor U24800 (N_24800,N_23105,N_23181);
and U24801 (N_24801,N_23454,N_23442);
nand U24802 (N_24802,N_23976,N_23783);
nand U24803 (N_24803,N_23002,N_23566);
nand U24804 (N_24804,N_23903,N_23093);
nor U24805 (N_24805,N_23329,N_23302);
nand U24806 (N_24806,N_23795,N_23839);
or U24807 (N_24807,N_23010,N_23980);
nand U24808 (N_24808,N_23467,N_23331);
xor U24809 (N_24809,N_23289,N_23589);
nand U24810 (N_24810,N_23554,N_23479);
nand U24811 (N_24811,N_23773,N_23163);
xnor U24812 (N_24812,N_23446,N_23222);
nand U24813 (N_24813,N_23552,N_23048);
or U24814 (N_24814,N_23793,N_23209);
or U24815 (N_24815,N_23786,N_23361);
or U24816 (N_24816,N_23511,N_23082);
xor U24817 (N_24817,N_23648,N_23738);
nand U24818 (N_24818,N_23155,N_23227);
xnor U24819 (N_24819,N_23827,N_23137);
and U24820 (N_24820,N_23612,N_23958);
xor U24821 (N_24821,N_23027,N_23292);
nand U24822 (N_24822,N_23944,N_23278);
or U24823 (N_24823,N_23334,N_23414);
nand U24824 (N_24824,N_23060,N_23282);
or U24825 (N_24825,N_23436,N_23936);
or U24826 (N_24826,N_23084,N_23209);
or U24827 (N_24827,N_23348,N_23763);
and U24828 (N_24828,N_23572,N_23557);
xor U24829 (N_24829,N_23055,N_23941);
xnor U24830 (N_24830,N_23298,N_23304);
and U24831 (N_24831,N_23080,N_23426);
and U24832 (N_24832,N_23846,N_23482);
xnor U24833 (N_24833,N_23177,N_23983);
xor U24834 (N_24834,N_23686,N_23843);
nor U24835 (N_24835,N_23167,N_23229);
and U24836 (N_24836,N_23224,N_23533);
or U24837 (N_24837,N_23433,N_23952);
and U24838 (N_24838,N_23040,N_23090);
or U24839 (N_24839,N_23398,N_23235);
or U24840 (N_24840,N_23920,N_23762);
or U24841 (N_24841,N_23418,N_23479);
and U24842 (N_24842,N_23095,N_23801);
and U24843 (N_24843,N_23183,N_23659);
nor U24844 (N_24844,N_23054,N_23939);
nor U24845 (N_24845,N_23083,N_23536);
xnor U24846 (N_24846,N_23581,N_23376);
nor U24847 (N_24847,N_23213,N_23587);
or U24848 (N_24848,N_23390,N_23700);
or U24849 (N_24849,N_23793,N_23009);
or U24850 (N_24850,N_23061,N_23985);
nor U24851 (N_24851,N_23053,N_23282);
and U24852 (N_24852,N_23240,N_23162);
nor U24853 (N_24853,N_23040,N_23451);
xor U24854 (N_24854,N_23707,N_23049);
nor U24855 (N_24855,N_23018,N_23771);
nand U24856 (N_24856,N_23778,N_23372);
or U24857 (N_24857,N_23327,N_23618);
nand U24858 (N_24858,N_23220,N_23537);
nand U24859 (N_24859,N_23768,N_23799);
xnor U24860 (N_24860,N_23359,N_23841);
xor U24861 (N_24861,N_23165,N_23619);
or U24862 (N_24862,N_23313,N_23608);
nand U24863 (N_24863,N_23825,N_23582);
and U24864 (N_24864,N_23980,N_23699);
or U24865 (N_24865,N_23654,N_23980);
or U24866 (N_24866,N_23679,N_23662);
nand U24867 (N_24867,N_23089,N_23484);
nand U24868 (N_24868,N_23899,N_23777);
and U24869 (N_24869,N_23568,N_23862);
or U24870 (N_24870,N_23470,N_23777);
or U24871 (N_24871,N_23377,N_23806);
nor U24872 (N_24872,N_23978,N_23586);
nand U24873 (N_24873,N_23397,N_23652);
xnor U24874 (N_24874,N_23852,N_23319);
nor U24875 (N_24875,N_23600,N_23406);
xnor U24876 (N_24876,N_23790,N_23922);
or U24877 (N_24877,N_23757,N_23740);
nand U24878 (N_24878,N_23672,N_23831);
or U24879 (N_24879,N_23273,N_23088);
or U24880 (N_24880,N_23117,N_23564);
nor U24881 (N_24881,N_23244,N_23941);
nor U24882 (N_24882,N_23794,N_23850);
and U24883 (N_24883,N_23076,N_23268);
and U24884 (N_24884,N_23976,N_23498);
and U24885 (N_24885,N_23660,N_23199);
and U24886 (N_24886,N_23428,N_23950);
nor U24887 (N_24887,N_23132,N_23963);
nand U24888 (N_24888,N_23815,N_23129);
or U24889 (N_24889,N_23481,N_23641);
nand U24890 (N_24890,N_23902,N_23723);
xor U24891 (N_24891,N_23846,N_23004);
nor U24892 (N_24892,N_23772,N_23715);
or U24893 (N_24893,N_23315,N_23060);
nor U24894 (N_24894,N_23393,N_23067);
xnor U24895 (N_24895,N_23907,N_23952);
and U24896 (N_24896,N_23600,N_23754);
and U24897 (N_24897,N_23207,N_23727);
nand U24898 (N_24898,N_23468,N_23130);
nor U24899 (N_24899,N_23099,N_23025);
nand U24900 (N_24900,N_23258,N_23123);
nand U24901 (N_24901,N_23038,N_23969);
nand U24902 (N_24902,N_23110,N_23052);
or U24903 (N_24903,N_23039,N_23446);
nor U24904 (N_24904,N_23947,N_23360);
or U24905 (N_24905,N_23028,N_23136);
xor U24906 (N_24906,N_23720,N_23317);
nand U24907 (N_24907,N_23232,N_23367);
nand U24908 (N_24908,N_23784,N_23497);
nor U24909 (N_24909,N_23865,N_23417);
xnor U24910 (N_24910,N_23839,N_23842);
xnor U24911 (N_24911,N_23939,N_23911);
nand U24912 (N_24912,N_23684,N_23346);
xnor U24913 (N_24913,N_23700,N_23189);
nand U24914 (N_24914,N_23915,N_23730);
or U24915 (N_24915,N_23069,N_23372);
nor U24916 (N_24916,N_23478,N_23217);
nand U24917 (N_24917,N_23701,N_23335);
or U24918 (N_24918,N_23886,N_23136);
and U24919 (N_24919,N_23883,N_23460);
or U24920 (N_24920,N_23755,N_23769);
and U24921 (N_24921,N_23386,N_23304);
or U24922 (N_24922,N_23422,N_23387);
xnor U24923 (N_24923,N_23407,N_23334);
nor U24924 (N_24924,N_23162,N_23219);
and U24925 (N_24925,N_23354,N_23245);
and U24926 (N_24926,N_23395,N_23839);
nor U24927 (N_24927,N_23104,N_23830);
or U24928 (N_24928,N_23702,N_23498);
and U24929 (N_24929,N_23135,N_23060);
or U24930 (N_24930,N_23855,N_23901);
and U24931 (N_24931,N_23599,N_23313);
and U24932 (N_24932,N_23454,N_23131);
or U24933 (N_24933,N_23910,N_23338);
xnor U24934 (N_24934,N_23183,N_23367);
nor U24935 (N_24935,N_23111,N_23753);
nor U24936 (N_24936,N_23732,N_23323);
xor U24937 (N_24937,N_23486,N_23494);
and U24938 (N_24938,N_23332,N_23749);
xnor U24939 (N_24939,N_23454,N_23827);
xnor U24940 (N_24940,N_23181,N_23980);
and U24941 (N_24941,N_23782,N_23598);
or U24942 (N_24942,N_23949,N_23542);
nand U24943 (N_24943,N_23122,N_23194);
nor U24944 (N_24944,N_23677,N_23962);
and U24945 (N_24945,N_23110,N_23286);
and U24946 (N_24946,N_23383,N_23638);
xnor U24947 (N_24947,N_23211,N_23417);
or U24948 (N_24948,N_23979,N_23847);
nor U24949 (N_24949,N_23136,N_23446);
or U24950 (N_24950,N_23501,N_23597);
nor U24951 (N_24951,N_23897,N_23049);
nand U24952 (N_24952,N_23081,N_23954);
nor U24953 (N_24953,N_23906,N_23517);
nor U24954 (N_24954,N_23750,N_23239);
xnor U24955 (N_24955,N_23087,N_23526);
xnor U24956 (N_24956,N_23103,N_23718);
or U24957 (N_24957,N_23210,N_23819);
nand U24958 (N_24958,N_23459,N_23475);
nand U24959 (N_24959,N_23237,N_23285);
nor U24960 (N_24960,N_23338,N_23190);
or U24961 (N_24961,N_23647,N_23849);
xor U24962 (N_24962,N_23706,N_23827);
nand U24963 (N_24963,N_23166,N_23133);
or U24964 (N_24964,N_23947,N_23385);
or U24965 (N_24965,N_23556,N_23627);
and U24966 (N_24966,N_23332,N_23790);
nor U24967 (N_24967,N_23806,N_23709);
and U24968 (N_24968,N_23992,N_23446);
or U24969 (N_24969,N_23627,N_23787);
or U24970 (N_24970,N_23963,N_23759);
nand U24971 (N_24971,N_23636,N_23207);
nand U24972 (N_24972,N_23529,N_23100);
nor U24973 (N_24973,N_23101,N_23608);
nor U24974 (N_24974,N_23703,N_23125);
or U24975 (N_24975,N_23239,N_23131);
nor U24976 (N_24976,N_23557,N_23712);
nand U24977 (N_24977,N_23252,N_23955);
xnor U24978 (N_24978,N_23638,N_23832);
xnor U24979 (N_24979,N_23049,N_23805);
nor U24980 (N_24980,N_23771,N_23120);
and U24981 (N_24981,N_23387,N_23456);
nand U24982 (N_24982,N_23016,N_23347);
nand U24983 (N_24983,N_23501,N_23897);
nand U24984 (N_24984,N_23542,N_23852);
or U24985 (N_24985,N_23902,N_23879);
xnor U24986 (N_24986,N_23625,N_23472);
and U24987 (N_24987,N_23887,N_23923);
and U24988 (N_24988,N_23876,N_23652);
xnor U24989 (N_24989,N_23591,N_23673);
or U24990 (N_24990,N_23724,N_23019);
or U24991 (N_24991,N_23369,N_23154);
nor U24992 (N_24992,N_23055,N_23823);
nor U24993 (N_24993,N_23459,N_23431);
xor U24994 (N_24994,N_23126,N_23540);
or U24995 (N_24995,N_23413,N_23848);
nand U24996 (N_24996,N_23476,N_23409);
or U24997 (N_24997,N_23941,N_23534);
and U24998 (N_24998,N_23742,N_23960);
xnor U24999 (N_24999,N_23355,N_23515);
and U25000 (N_25000,N_24927,N_24064);
nor U25001 (N_25001,N_24906,N_24628);
xnor U25002 (N_25002,N_24698,N_24543);
and U25003 (N_25003,N_24940,N_24181);
and U25004 (N_25004,N_24569,N_24886);
nor U25005 (N_25005,N_24245,N_24887);
nor U25006 (N_25006,N_24148,N_24345);
or U25007 (N_25007,N_24807,N_24743);
and U25008 (N_25008,N_24229,N_24176);
or U25009 (N_25009,N_24973,N_24028);
nor U25010 (N_25010,N_24739,N_24109);
nor U25011 (N_25011,N_24343,N_24526);
or U25012 (N_25012,N_24684,N_24240);
or U25013 (N_25013,N_24700,N_24276);
or U25014 (N_25014,N_24018,N_24542);
nor U25015 (N_25015,N_24790,N_24958);
nand U25016 (N_25016,N_24004,N_24061);
or U25017 (N_25017,N_24034,N_24848);
and U25018 (N_25018,N_24406,N_24688);
nor U25019 (N_25019,N_24072,N_24612);
nand U25020 (N_25020,N_24454,N_24771);
or U25021 (N_25021,N_24507,N_24947);
nand U25022 (N_25022,N_24270,N_24726);
xor U25023 (N_25023,N_24400,N_24774);
nor U25024 (N_25024,N_24680,N_24335);
nand U25025 (N_25025,N_24627,N_24528);
and U25026 (N_25026,N_24172,N_24673);
and U25027 (N_25027,N_24556,N_24896);
and U25028 (N_25028,N_24654,N_24185);
nand U25029 (N_25029,N_24697,N_24530);
nand U25030 (N_25030,N_24911,N_24226);
nor U25031 (N_25031,N_24557,N_24024);
and U25032 (N_25032,N_24433,N_24816);
and U25033 (N_25033,N_24337,N_24964);
and U25034 (N_25034,N_24128,N_24385);
xor U25035 (N_25035,N_24859,N_24141);
nand U25036 (N_25036,N_24699,N_24903);
and U25037 (N_25037,N_24564,N_24768);
or U25038 (N_25038,N_24231,N_24279);
and U25039 (N_25039,N_24863,N_24587);
or U25040 (N_25040,N_24716,N_24455);
xnor U25041 (N_25041,N_24983,N_24264);
or U25042 (N_25042,N_24052,N_24630);
xnor U25043 (N_25043,N_24670,N_24463);
nor U25044 (N_25044,N_24363,N_24675);
and U25045 (N_25045,N_24418,N_24972);
xnor U25046 (N_25046,N_24219,N_24519);
xnor U25047 (N_25047,N_24862,N_24312);
nand U25048 (N_25048,N_24732,N_24423);
xor U25049 (N_25049,N_24509,N_24429);
nand U25050 (N_25050,N_24459,N_24549);
nand U25051 (N_25051,N_24631,N_24171);
and U25052 (N_25052,N_24250,N_24856);
nor U25053 (N_25053,N_24646,N_24763);
nand U25054 (N_25054,N_24137,N_24939);
nand U25055 (N_25055,N_24027,N_24336);
nand U25056 (N_25056,N_24709,N_24382);
and U25057 (N_25057,N_24754,N_24537);
nand U25058 (N_25058,N_24127,N_24092);
and U25059 (N_25059,N_24523,N_24489);
or U25060 (N_25060,N_24998,N_24495);
nor U25061 (N_25061,N_24042,N_24291);
or U25062 (N_25062,N_24843,N_24297);
and U25063 (N_25063,N_24305,N_24430);
nand U25064 (N_25064,N_24550,N_24540);
or U25065 (N_25065,N_24908,N_24545);
xor U25066 (N_25066,N_24987,N_24614);
nand U25067 (N_25067,N_24687,N_24205);
nor U25068 (N_25068,N_24031,N_24686);
nor U25069 (N_25069,N_24645,N_24674);
or U25070 (N_25070,N_24585,N_24167);
nand U25071 (N_25071,N_24261,N_24837);
nand U25072 (N_25072,N_24131,N_24573);
nor U25073 (N_25073,N_24602,N_24372);
or U25074 (N_25074,N_24232,N_24010);
or U25075 (N_25075,N_24875,N_24020);
nand U25076 (N_25076,N_24281,N_24230);
nand U25077 (N_25077,N_24233,N_24002);
nor U25078 (N_25078,N_24574,N_24635);
nor U25079 (N_25079,N_24085,N_24050);
xnor U25080 (N_25080,N_24091,N_24346);
and U25081 (N_25081,N_24681,N_24948);
xor U25082 (N_25082,N_24154,N_24701);
and U25083 (N_25083,N_24431,N_24100);
nand U25084 (N_25084,N_24373,N_24228);
xnor U25085 (N_25085,N_24473,N_24084);
or U25086 (N_25086,N_24753,N_24620);
nand U25087 (N_25087,N_24932,N_24718);
xor U25088 (N_25088,N_24395,N_24211);
and U25089 (N_25089,N_24394,N_24735);
and U25090 (N_25090,N_24969,N_24356);
and U25091 (N_25091,N_24090,N_24477);
nand U25092 (N_25092,N_24355,N_24583);
or U25093 (N_25093,N_24491,N_24227);
xor U25094 (N_25094,N_24640,N_24685);
and U25095 (N_25095,N_24444,N_24009);
nand U25096 (N_25096,N_24835,N_24182);
nor U25097 (N_25097,N_24340,N_24876);
xnor U25098 (N_25098,N_24690,N_24821);
nor U25099 (N_25099,N_24599,N_24584);
nand U25100 (N_25100,N_24575,N_24005);
xnor U25101 (N_25101,N_24970,N_24360);
nor U25102 (N_25102,N_24689,N_24854);
xnor U25103 (N_25103,N_24191,N_24610);
or U25104 (N_25104,N_24524,N_24235);
nand U25105 (N_25105,N_24300,N_24525);
nand U25106 (N_25106,N_24707,N_24963);
nor U25107 (N_25107,N_24462,N_24880);
nand U25108 (N_25108,N_24581,N_24480);
and U25109 (N_25109,N_24249,N_24458);
and U25110 (N_25110,N_24098,N_24273);
xnor U25111 (N_25111,N_24658,N_24762);
nand U25112 (N_25112,N_24781,N_24015);
nand U25113 (N_25113,N_24499,N_24286);
and U25114 (N_25114,N_24888,N_24786);
and U25115 (N_25115,N_24012,N_24590);
or U25116 (N_25116,N_24745,N_24303);
or U25117 (N_25117,N_24190,N_24905);
xnor U25118 (N_25118,N_24955,N_24892);
nor U25119 (N_25119,N_24466,N_24660);
nor U25120 (N_25120,N_24889,N_24330);
or U25121 (N_25121,N_24915,N_24661);
or U25122 (N_25122,N_24870,N_24693);
nand U25123 (N_25123,N_24323,N_24411);
xor U25124 (N_25124,N_24795,N_24421);
nor U25125 (N_25125,N_24502,N_24089);
and U25126 (N_25126,N_24634,N_24551);
nand U25127 (N_25127,N_24819,N_24078);
nor U25128 (N_25128,N_24313,N_24285);
and U25129 (N_25129,N_24357,N_24508);
nor U25130 (N_25130,N_24811,N_24597);
or U25131 (N_25131,N_24598,N_24571);
xor U25132 (N_25132,N_24033,N_24731);
nand U25133 (N_25133,N_24222,N_24368);
or U25134 (N_25134,N_24582,N_24445);
nand U25135 (N_25135,N_24505,N_24215);
nand U25136 (N_25136,N_24725,N_24319);
and U25137 (N_25137,N_24621,N_24941);
xnor U25138 (N_25138,N_24653,N_24991);
and U25139 (N_25139,N_24138,N_24760);
xnor U25140 (N_25140,N_24331,N_24021);
xor U25141 (N_25141,N_24103,N_24516);
xor U25142 (N_25142,N_24568,N_24006);
nand U25143 (N_25143,N_24825,N_24828);
nand U25144 (N_25144,N_24500,N_24649);
xnor U25145 (N_25145,N_24920,N_24623);
xnor U25146 (N_25146,N_24405,N_24789);
nor U25147 (N_25147,N_24785,N_24521);
and U25148 (N_25148,N_24759,N_24490);
and U25149 (N_25149,N_24456,N_24591);
or U25150 (N_25150,N_24334,N_24643);
or U25151 (N_25151,N_24362,N_24189);
and U25152 (N_25152,N_24810,N_24910);
nand U25153 (N_25153,N_24208,N_24570);
nand U25154 (N_25154,N_24923,N_24580);
nor U25155 (N_25155,N_24861,N_24217);
nor U25156 (N_25156,N_24596,N_24600);
or U25157 (N_25157,N_24472,N_24413);
nand U25158 (N_25158,N_24225,N_24277);
xnor U25159 (N_25159,N_24199,N_24997);
nand U25160 (N_25160,N_24943,N_24547);
and U25161 (N_25161,N_24946,N_24953);
xor U25162 (N_25162,N_24691,N_24160);
xnor U25163 (N_25163,N_24197,N_24769);
or U25164 (N_25164,N_24173,N_24982);
and U25165 (N_25165,N_24717,N_24517);
and U25166 (N_25166,N_24038,N_24234);
or U25167 (N_25167,N_24711,N_24874);
xnor U25168 (N_25168,N_24265,N_24989);
nand U25169 (N_25169,N_24986,N_24164);
nand U25170 (N_25170,N_24655,N_24678);
xor U25171 (N_25171,N_24579,N_24961);
xnor U25172 (N_25172,N_24377,N_24813);
and U25173 (N_25173,N_24398,N_24605);
xnor U25174 (N_25174,N_24301,N_24284);
and U25175 (N_25175,N_24352,N_24316);
and U25176 (N_25176,N_24387,N_24648);
nand U25177 (N_25177,N_24026,N_24820);
nand U25178 (N_25178,N_24396,N_24783);
xnor U25179 (N_25179,N_24824,N_24901);
or U25180 (N_25180,N_24529,N_24822);
or U25181 (N_25181,N_24102,N_24375);
and U25182 (N_25182,N_24294,N_24259);
and U25183 (N_25183,N_24081,N_24916);
or U25184 (N_25184,N_24310,N_24485);
xor U25185 (N_25185,N_24317,N_24761);
or U25186 (N_25186,N_24036,N_24562);
and U25187 (N_25187,N_24194,N_24683);
and U25188 (N_25188,N_24840,N_24775);
or U25189 (N_25189,N_24358,N_24133);
and U25190 (N_25190,N_24115,N_24032);
nand U25191 (N_25191,N_24384,N_24978);
xor U25192 (N_25192,N_24696,N_24296);
and U25193 (N_25193,N_24980,N_24512);
and U25194 (N_25194,N_24535,N_24757);
or U25195 (N_25195,N_24515,N_24561);
nor U25196 (N_25196,N_24846,N_24283);
and U25197 (N_25197,N_24143,N_24448);
nand U25198 (N_25198,N_24094,N_24770);
or U25199 (N_25199,N_24086,N_24314);
nand U25200 (N_25200,N_24814,N_24909);
and U25201 (N_25201,N_24304,N_24936);
nor U25202 (N_25202,N_24728,N_24101);
nand U25203 (N_25203,N_24344,N_24705);
xnor U25204 (N_25204,N_24367,N_24944);
or U25205 (N_25205,N_24773,N_24341);
and U25206 (N_25206,N_24642,N_24324);
and U25207 (N_25207,N_24510,N_24243);
or U25208 (N_25208,N_24200,N_24682);
or U25209 (N_25209,N_24794,N_24424);
and U25210 (N_25210,N_24262,N_24125);
nor U25211 (N_25211,N_24639,N_24720);
nor U25212 (N_25212,N_24134,N_24095);
or U25213 (N_25213,N_24984,N_24504);
nand U25214 (N_25214,N_24592,N_24275);
xor U25215 (N_25215,N_24615,N_24255);
or U25216 (N_25216,N_24945,N_24126);
or U25217 (N_25217,N_24206,N_24730);
and U25218 (N_25218,N_24890,N_24938);
xnor U25219 (N_25219,N_24046,N_24838);
xor U25220 (N_25220,N_24666,N_24800);
nor U25221 (N_25221,N_24899,N_24295);
and U25222 (N_25222,N_24121,N_24546);
and U25223 (N_25223,N_24062,N_24392);
and U25224 (N_25224,N_24604,N_24016);
nand U25225 (N_25225,N_24808,N_24952);
nor U25226 (N_25226,N_24609,N_24864);
and U25227 (N_25227,N_24879,N_24798);
or U25228 (N_25228,N_24727,N_24193);
xnor U25229 (N_25229,N_24823,N_24659);
and U25230 (N_25230,N_24306,N_24999);
nand U25231 (N_25231,N_24934,N_24204);
and U25232 (N_25232,N_24047,N_24636);
nor U25233 (N_25233,N_24566,N_24054);
xnor U25234 (N_25234,N_24147,N_24110);
nand U25235 (N_25235,N_24928,N_24067);
or U25236 (N_25236,N_24221,N_24216);
and U25237 (N_25237,N_24567,N_24282);
or U25238 (N_25238,N_24198,N_24494);
xor U25239 (N_25239,N_24307,N_24071);
and U25240 (N_25240,N_24169,N_24959);
or U25241 (N_25241,N_24393,N_24122);
or U25242 (N_25242,N_24513,N_24073);
or U25243 (N_25243,N_24750,N_24871);
and U25244 (N_25244,N_24447,N_24170);
or U25245 (N_25245,N_24428,N_24267);
and U25246 (N_25246,N_24611,N_24647);
xnor U25247 (N_25247,N_24900,N_24117);
xnor U25248 (N_25248,N_24256,N_24558);
nand U25249 (N_25249,N_24704,N_24175);
and U25250 (N_25250,N_24347,N_24155);
xnor U25251 (N_25251,N_24001,N_24248);
nand U25252 (N_25252,N_24464,N_24309);
nand U25253 (N_25253,N_24981,N_24734);
xnor U25254 (N_25254,N_24403,N_24142);
nor U25255 (N_25255,N_24410,N_24626);
or U25256 (N_25256,N_24805,N_24487);
nor U25257 (N_25257,N_24440,N_24253);
nor U25258 (N_25258,N_24378,N_24804);
or U25259 (N_25259,N_24246,N_24412);
xnor U25260 (N_25260,N_24207,N_24667);
xnor U25261 (N_25261,N_24552,N_24694);
nor U25262 (N_25262,N_24853,N_24765);
nor U25263 (N_25263,N_24030,N_24797);
nand U25264 (N_25264,N_24299,N_24070);
or U25265 (N_25265,N_24153,N_24325);
nand U25266 (N_25266,N_24632,N_24326);
and U25267 (N_25267,N_24118,N_24977);
nor U25268 (N_25268,N_24293,N_24877);
nand U25269 (N_25269,N_24132,N_24722);
xor U25270 (N_25270,N_24873,N_24937);
nand U25271 (N_25271,N_24617,N_24503);
xnor U25272 (N_25272,N_24586,N_24435);
nor U25273 (N_25273,N_24799,N_24359);
xnor U25274 (N_25274,N_24520,N_24269);
and U25275 (N_25275,N_24388,N_24565);
or U25276 (N_25276,N_24342,N_24292);
xor U25277 (N_25277,N_24629,N_24979);
or U25278 (N_25278,N_24376,N_24966);
or U25279 (N_25279,N_24511,N_24404);
or U25280 (N_25280,N_24793,N_24338);
and U25281 (N_25281,N_24534,N_24214);
nor U25282 (N_25282,N_24322,N_24651);
xor U25283 (N_25283,N_24606,N_24842);
nand U25284 (N_25284,N_24135,N_24633);
nand U25285 (N_25285,N_24851,N_24482);
or U25286 (N_25286,N_24601,N_24518);
nor U25287 (N_25287,N_24907,N_24266);
nand U25288 (N_25288,N_24733,N_24637);
xnor U25289 (N_25289,N_24492,N_24451);
xnor U25290 (N_25290,N_24622,N_24721);
nor U25291 (N_25291,N_24136,N_24151);
nor U25292 (N_25292,N_24465,N_24802);
nand U25293 (N_25293,N_24619,N_24895);
or U25294 (N_25294,N_24419,N_24272);
xnor U25295 (N_25295,N_24860,N_24752);
nand U25296 (N_25296,N_24778,N_24595);
xnor U25297 (N_25297,N_24975,N_24244);
and U25298 (N_25298,N_24531,N_24120);
nor U25299 (N_25299,N_24123,N_24641);
or U25300 (N_25300,N_24056,N_24203);
or U25301 (N_25301,N_24087,N_24029);
or U25302 (N_25302,N_24383,N_24559);
nand U25303 (N_25303,N_24349,N_24608);
and U25304 (N_25304,N_24483,N_24498);
or U25305 (N_25305,N_24076,N_24833);
nor U25306 (N_25306,N_24729,N_24241);
xor U25307 (N_25307,N_24594,N_24099);
xor U25308 (N_25308,N_24539,N_24933);
nor U25309 (N_25309,N_24957,N_24224);
nand U25310 (N_25310,N_24374,N_24152);
or U25311 (N_25311,N_24926,N_24994);
and U25312 (N_25312,N_24104,N_24665);
and U25313 (N_25313,N_24960,N_24662);
xor U25314 (N_25314,N_24782,N_24467);
xor U25315 (N_25315,N_24201,N_24919);
nand U25316 (N_25316,N_24845,N_24075);
or U25317 (N_25317,N_24710,N_24008);
nand U25318 (N_25318,N_24827,N_24514);
nand U25319 (N_25319,N_24327,N_24014);
nand U25320 (N_25320,N_24818,N_24025);
and U25321 (N_25321,N_24302,N_24497);
and U25322 (N_25322,N_24386,N_24638);
and U25323 (N_25323,N_24847,N_24478);
and U25324 (N_25324,N_24917,N_24949);
nor U25325 (N_25325,N_24407,N_24348);
and U25326 (N_25326,N_24736,N_24351);
nand U25327 (N_25327,N_24780,N_24116);
nor U25328 (N_25328,N_24105,N_24218);
or U25329 (N_25329,N_24817,N_24011);
nand U25330 (N_25330,N_24213,N_24985);
xnor U25331 (N_25331,N_24437,N_24059);
or U25332 (N_25332,N_24187,N_24974);
and U25333 (N_25333,N_24695,N_24988);
or U25334 (N_25334,N_24792,N_24409);
nor U25335 (N_25335,N_24210,N_24486);
and U25336 (N_25336,N_24616,N_24252);
and U25337 (N_25337,N_24278,N_24914);
nor U25338 (N_25338,N_24751,N_24311);
nand U25339 (N_25339,N_24040,N_24223);
nor U25340 (N_25340,N_24671,N_24784);
nor U25341 (N_25341,N_24069,N_24365);
xnor U25342 (N_25342,N_24831,N_24422);
and U25343 (N_25343,N_24399,N_24408);
and U25344 (N_25344,N_24723,N_24239);
nand U25345 (N_25345,N_24755,N_24186);
and U25346 (N_25346,N_24402,N_24107);
and U25347 (N_25347,N_24268,N_24113);
nand U25348 (N_25348,N_24902,N_24850);
nor U25349 (N_25349,N_24749,N_24114);
or U25350 (N_25350,N_24692,N_24578);
xor U25351 (N_25351,N_24891,N_24867);
xnor U25352 (N_25352,N_24082,N_24446);
and U25353 (N_25353,N_24488,N_24942);
and U25354 (N_25354,N_24737,N_24339);
nor U25355 (N_25355,N_24390,N_24019);
and U25356 (N_25356,N_24996,N_24414);
or U25357 (N_25357,N_24878,N_24209);
nand U25358 (N_25358,N_24333,N_24298);
xnor U25359 (N_25359,N_24003,N_24929);
xor U25360 (N_25360,N_24922,N_24391);
and U25361 (N_25361,N_24180,N_24048);
nor U25362 (N_25362,N_24049,N_24872);
and U25363 (N_25363,N_24603,N_24380);
xor U25364 (N_25364,N_24897,N_24772);
nor U25365 (N_25365,N_24656,N_24280);
xnor U25366 (N_25366,N_24868,N_24449);
xnor U25367 (N_25367,N_24787,N_24247);
nand U25368 (N_25368,N_24544,N_24476);
nand U25369 (N_25369,N_24777,N_24063);
xnor U25370 (N_25370,N_24884,N_24533);
or U25371 (N_25371,N_24858,N_24166);
nor U25372 (N_25372,N_24976,N_24401);
nand U25373 (N_25373,N_24812,N_24432);
and U25374 (N_25374,N_24625,N_24714);
and U25375 (N_25375,N_24904,N_24703);
or U25376 (N_25376,N_24174,N_24013);
or U25377 (N_25377,N_24000,N_24044);
nor U25378 (N_25378,N_24066,N_24719);
nand U25379 (N_25379,N_24041,N_24053);
xor U25380 (N_25380,N_24251,N_24971);
and U25381 (N_25381,N_24935,N_24108);
and U25382 (N_25382,N_24950,N_24381);
or U25383 (N_25383,N_24663,N_24161);
xor U25384 (N_25384,N_24826,N_24260);
nor U25385 (N_25385,N_24921,N_24740);
nor U25386 (N_25386,N_24058,N_24441);
and U25387 (N_25387,N_24724,N_24677);
nor U25388 (N_25388,N_24184,N_24150);
nor U25389 (N_25389,N_24589,N_24274);
or U25390 (N_25390,N_24650,N_24885);
and U25391 (N_25391,N_24664,N_24438);
or U25392 (N_25392,N_24457,N_24366);
nor U25393 (N_25393,N_24263,N_24967);
nand U25394 (N_25394,N_24162,N_24079);
nor U25395 (N_25395,N_24912,N_24869);
or U25396 (N_25396,N_24758,N_24715);
nor U25397 (N_25397,N_24993,N_24669);
and U25398 (N_25398,N_24962,N_24506);
nor U25399 (N_25399,N_24088,N_24744);
or U25400 (N_25400,N_24748,N_24179);
nand U25401 (N_25401,N_24146,N_24130);
nor U25402 (N_25402,N_24475,N_24237);
and U25403 (N_25403,N_24443,N_24157);
nand U25404 (N_25404,N_24841,N_24055);
nand U25405 (N_25405,N_24924,N_24644);
or U25406 (N_25406,N_24183,N_24708);
nor U25407 (N_25407,N_24657,N_24470);
and U25408 (N_25408,N_24254,N_24865);
or U25409 (N_25409,N_24555,N_24796);
nor U25410 (N_25410,N_24995,N_24434);
nand U25411 (N_25411,N_24236,N_24124);
xor U25412 (N_25412,N_24397,N_24163);
and U25413 (N_25413,N_24168,N_24192);
nand U25414 (N_25414,N_24536,N_24767);
xnor U25415 (N_25415,N_24832,N_24741);
nor U25416 (N_25416,N_24140,N_24990);
nor U25417 (N_25417,N_24144,N_24427);
xor U25418 (N_25418,N_24149,N_24954);
nand U25419 (N_25419,N_24474,N_24425);
or U25420 (N_25420,N_24436,N_24051);
and U25421 (N_25421,N_24083,N_24442);
and U25422 (N_25422,N_24925,N_24290);
nand U25423 (N_25423,N_24764,N_24057);
nand U25424 (N_25424,N_24389,N_24145);
nand U25425 (N_25425,N_24415,N_24951);
or U25426 (N_25426,N_24844,N_24188);
nand U25427 (N_25427,N_24830,N_24527);
nor U25428 (N_25428,N_24364,N_24713);
nor U25429 (N_25429,N_24829,N_24676);
nand U25430 (N_25430,N_24112,N_24624);
or U25431 (N_25431,N_24652,N_24965);
and U25432 (N_25432,N_24746,N_24756);
xnor U25433 (N_25433,N_24332,N_24672);
nand U25434 (N_25434,N_24548,N_24017);
or U25435 (N_25435,N_24893,N_24484);
xor U25436 (N_25436,N_24460,N_24468);
nand U25437 (N_25437,N_24461,N_24815);
nor U25438 (N_25438,N_24111,N_24481);
nand U25439 (N_25439,N_24866,N_24956);
and U25440 (N_25440,N_24289,N_24852);
or U25441 (N_25441,N_24855,N_24097);
xor U25442 (N_25442,N_24212,N_24139);
xnor U25443 (N_25443,N_24857,N_24096);
or U25444 (N_25444,N_24035,N_24060);
xnor U25445 (N_25445,N_24318,N_24883);
nand U25446 (N_25446,N_24238,N_24093);
xnor U25447 (N_25447,N_24522,N_24881);
and U25448 (N_25448,N_24023,N_24037);
and U25449 (N_25449,N_24560,N_24308);
and U25450 (N_25450,N_24668,N_24287);
nor U25451 (N_25451,N_24766,N_24450);
and U25452 (N_25452,N_24894,N_24022);
nor U25453 (N_25453,N_24452,N_24258);
nand U25454 (N_25454,N_24159,N_24479);
or U25455 (N_25455,N_24968,N_24321);
nor U25456 (N_25456,N_24165,N_24074);
or U25457 (N_25457,N_24679,N_24532);
xor U25458 (N_25458,N_24618,N_24077);
nor U25459 (N_25459,N_24271,N_24242);
nor U25460 (N_25460,N_24469,N_24329);
xnor U25461 (N_25461,N_24177,N_24007);
nand U25462 (N_25462,N_24613,N_24803);
nor U25463 (N_25463,N_24320,N_24379);
xnor U25464 (N_25464,N_24913,N_24426);
nand U25465 (N_25465,N_24065,N_24195);
xnor U25466 (N_25466,N_24834,N_24501);
and U25467 (N_25467,N_24738,N_24839);
nand U25468 (N_25468,N_24315,N_24538);
or U25469 (N_25469,N_24416,N_24776);
nor U25470 (N_25470,N_24220,N_24119);
nand U25471 (N_25471,N_24553,N_24747);
xor U25472 (N_25472,N_24806,N_24039);
nor U25473 (N_25473,N_24493,N_24779);
and U25474 (N_25474,N_24809,N_24043);
xnor U25475 (N_25475,N_24045,N_24836);
nand U25476 (N_25476,N_24420,N_24080);
nor U25477 (N_25477,N_24702,N_24471);
and U25478 (N_25478,N_24369,N_24350);
and U25479 (N_25479,N_24202,N_24572);
and U25480 (N_25480,N_24439,N_24156);
nand U25481 (N_25481,N_24918,N_24196);
nand U25482 (N_25482,N_24577,N_24849);
nand U25483 (N_25483,N_24068,N_24554);
nor U25484 (N_25484,N_24417,N_24453);
nand U25485 (N_25485,N_24882,N_24158);
nor U25486 (N_25486,N_24588,N_24178);
xor U25487 (N_25487,N_24742,N_24931);
nand U25488 (N_25488,N_24607,N_24791);
nand U25489 (N_25489,N_24129,N_24801);
nand U25490 (N_25490,N_24788,N_24257);
nor U25491 (N_25491,N_24496,N_24541);
xnor U25492 (N_25492,N_24706,N_24712);
and U25493 (N_25493,N_24371,N_24576);
or U25494 (N_25494,N_24992,N_24593);
or U25495 (N_25495,N_24106,N_24930);
nand U25496 (N_25496,N_24361,N_24328);
or U25497 (N_25497,N_24354,N_24898);
xor U25498 (N_25498,N_24563,N_24370);
nor U25499 (N_25499,N_24353,N_24288);
and U25500 (N_25500,N_24628,N_24274);
or U25501 (N_25501,N_24128,N_24618);
and U25502 (N_25502,N_24560,N_24154);
xor U25503 (N_25503,N_24916,N_24658);
xnor U25504 (N_25504,N_24674,N_24329);
and U25505 (N_25505,N_24184,N_24447);
and U25506 (N_25506,N_24935,N_24680);
nand U25507 (N_25507,N_24802,N_24766);
nor U25508 (N_25508,N_24820,N_24595);
or U25509 (N_25509,N_24738,N_24879);
and U25510 (N_25510,N_24632,N_24372);
nor U25511 (N_25511,N_24416,N_24579);
nand U25512 (N_25512,N_24001,N_24116);
or U25513 (N_25513,N_24150,N_24235);
nand U25514 (N_25514,N_24798,N_24490);
nand U25515 (N_25515,N_24434,N_24152);
nor U25516 (N_25516,N_24395,N_24610);
nand U25517 (N_25517,N_24976,N_24995);
xnor U25518 (N_25518,N_24526,N_24326);
and U25519 (N_25519,N_24442,N_24947);
nand U25520 (N_25520,N_24843,N_24983);
and U25521 (N_25521,N_24837,N_24781);
nor U25522 (N_25522,N_24553,N_24198);
xnor U25523 (N_25523,N_24774,N_24078);
and U25524 (N_25524,N_24187,N_24257);
xnor U25525 (N_25525,N_24969,N_24966);
or U25526 (N_25526,N_24857,N_24886);
and U25527 (N_25527,N_24711,N_24142);
and U25528 (N_25528,N_24757,N_24126);
and U25529 (N_25529,N_24572,N_24861);
xor U25530 (N_25530,N_24729,N_24607);
nand U25531 (N_25531,N_24686,N_24459);
or U25532 (N_25532,N_24260,N_24534);
nand U25533 (N_25533,N_24279,N_24658);
nand U25534 (N_25534,N_24149,N_24056);
nand U25535 (N_25535,N_24764,N_24337);
and U25536 (N_25536,N_24038,N_24832);
nand U25537 (N_25537,N_24909,N_24727);
nand U25538 (N_25538,N_24924,N_24780);
and U25539 (N_25539,N_24426,N_24908);
and U25540 (N_25540,N_24803,N_24776);
and U25541 (N_25541,N_24996,N_24959);
nand U25542 (N_25542,N_24316,N_24544);
nor U25543 (N_25543,N_24055,N_24089);
xnor U25544 (N_25544,N_24545,N_24561);
nor U25545 (N_25545,N_24272,N_24268);
or U25546 (N_25546,N_24289,N_24048);
xnor U25547 (N_25547,N_24746,N_24520);
nor U25548 (N_25548,N_24431,N_24077);
or U25549 (N_25549,N_24087,N_24581);
xnor U25550 (N_25550,N_24638,N_24250);
xor U25551 (N_25551,N_24284,N_24374);
nand U25552 (N_25552,N_24486,N_24967);
or U25553 (N_25553,N_24557,N_24570);
nor U25554 (N_25554,N_24421,N_24847);
and U25555 (N_25555,N_24714,N_24106);
nand U25556 (N_25556,N_24576,N_24377);
xor U25557 (N_25557,N_24052,N_24983);
xor U25558 (N_25558,N_24344,N_24738);
xnor U25559 (N_25559,N_24401,N_24684);
nand U25560 (N_25560,N_24358,N_24578);
nor U25561 (N_25561,N_24091,N_24224);
or U25562 (N_25562,N_24989,N_24787);
or U25563 (N_25563,N_24423,N_24302);
xor U25564 (N_25564,N_24637,N_24562);
nand U25565 (N_25565,N_24062,N_24439);
and U25566 (N_25566,N_24423,N_24573);
nor U25567 (N_25567,N_24909,N_24155);
xnor U25568 (N_25568,N_24242,N_24521);
xor U25569 (N_25569,N_24168,N_24600);
or U25570 (N_25570,N_24703,N_24300);
or U25571 (N_25571,N_24827,N_24451);
or U25572 (N_25572,N_24213,N_24939);
xnor U25573 (N_25573,N_24500,N_24381);
nor U25574 (N_25574,N_24223,N_24511);
nand U25575 (N_25575,N_24737,N_24841);
and U25576 (N_25576,N_24255,N_24973);
xnor U25577 (N_25577,N_24438,N_24054);
nor U25578 (N_25578,N_24734,N_24583);
xor U25579 (N_25579,N_24324,N_24380);
or U25580 (N_25580,N_24709,N_24099);
and U25581 (N_25581,N_24320,N_24100);
nand U25582 (N_25582,N_24442,N_24603);
xnor U25583 (N_25583,N_24244,N_24827);
nor U25584 (N_25584,N_24054,N_24763);
xor U25585 (N_25585,N_24124,N_24989);
xor U25586 (N_25586,N_24025,N_24530);
nand U25587 (N_25587,N_24314,N_24658);
nand U25588 (N_25588,N_24811,N_24159);
nand U25589 (N_25589,N_24982,N_24081);
xor U25590 (N_25590,N_24781,N_24510);
xor U25591 (N_25591,N_24481,N_24772);
nor U25592 (N_25592,N_24421,N_24127);
nand U25593 (N_25593,N_24714,N_24903);
xor U25594 (N_25594,N_24199,N_24160);
or U25595 (N_25595,N_24935,N_24240);
and U25596 (N_25596,N_24106,N_24302);
nand U25597 (N_25597,N_24171,N_24501);
or U25598 (N_25598,N_24811,N_24143);
or U25599 (N_25599,N_24302,N_24702);
nand U25600 (N_25600,N_24768,N_24225);
nor U25601 (N_25601,N_24801,N_24378);
and U25602 (N_25602,N_24709,N_24638);
nand U25603 (N_25603,N_24414,N_24130);
nor U25604 (N_25604,N_24913,N_24114);
nor U25605 (N_25605,N_24684,N_24261);
nand U25606 (N_25606,N_24239,N_24325);
and U25607 (N_25607,N_24098,N_24224);
xnor U25608 (N_25608,N_24038,N_24465);
or U25609 (N_25609,N_24742,N_24343);
nor U25610 (N_25610,N_24528,N_24128);
or U25611 (N_25611,N_24683,N_24640);
nand U25612 (N_25612,N_24167,N_24460);
or U25613 (N_25613,N_24237,N_24614);
nand U25614 (N_25614,N_24834,N_24446);
and U25615 (N_25615,N_24706,N_24214);
nor U25616 (N_25616,N_24957,N_24604);
nor U25617 (N_25617,N_24355,N_24848);
nand U25618 (N_25618,N_24696,N_24795);
nor U25619 (N_25619,N_24376,N_24216);
and U25620 (N_25620,N_24968,N_24524);
or U25621 (N_25621,N_24271,N_24016);
nor U25622 (N_25622,N_24560,N_24783);
and U25623 (N_25623,N_24169,N_24870);
nor U25624 (N_25624,N_24029,N_24878);
or U25625 (N_25625,N_24001,N_24162);
nor U25626 (N_25626,N_24130,N_24759);
and U25627 (N_25627,N_24071,N_24694);
xor U25628 (N_25628,N_24988,N_24517);
nand U25629 (N_25629,N_24043,N_24366);
and U25630 (N_25630,N_24761,N_24326);
xor U25631 (N_25631,N_24672,N_24797);
or U25632 (N_25632,N_24387,N_24216);
nor U25633 (N_25633,N_24208,N_24724);
and U25634 (N_25634,N_24778,N_24251);
nor U25635 (N_25635,N_24594,N_24413);
or U25636 (N_25636,N_24060,N_24745);
nand U25637 (N_25637,N_24183,N_24268);
or U25638 (N_25638,N_24105,N_24740);
or U25639 (N_25639,N_24252,N_24343);
nor U25640 (N_25640,N_24295,N_24008);
or U25641 (N_25641,N_24356,N_24251);
or U25642 (N_25642,N_24962,N_24212);
and U25643 (N_25643,N_24086,N_24005);
xor U25644 (N_25644,N_24027,N_24519);
nand U25645 (N_25645,N_24688,N_24869);
xnor U25646 (N_25646,N_24666,N_24510);
and U25647 (N_25647,N_24951,N_24763);
or U25648 (N_25648,N_24036,N_24329);
or U25649 (N_25649,N_24126,N_24484);
and U25650 (N_25650,N_24562,N_24103);
nor U25651 (N_25651,N_24737,N_24217);
nand U25652 (N_25652,N_24031,N_24488);
nor U25653 (N_25653,N_24450,N_24881);
nor U25654 (N_25654,N_24561,N_24261);
nand U25655 (N_25655,N_24974,N_24069);
or U25656 (N_25656,N_24478,N_24679);
and U25657 (N_25657,N_24592,N_24210);
or U25658 (N_25658,N_24783,N_24038);
nor U25659 (N_25659,N_24038,N_24487);
and U25660 (N_25660,N_24810,N_24808);
nand U25661 (N_25661,N_24223,N_24625);
xor U25662 (N_25662,N_24944,N_24371);
nor U25663 (N_25663,N_24939,N_24928);
nor U25664 (N_25664,N_24593,N_24605);
and U25665 (N_25665,N_24548,N_24417);
xor U25666 (N_25666,N_24845,N_24233);
nor U25667 (N_25667,N_24810,N_24616);
or U25668 (N_25668,N_24388,N_24632);
nor U25669 (N_25669,N_24820,N_24723);
xnor U25670 (N_25670,N_24729,N_24439);
or U25671 (N_25671,N_24419,N_24024);
or U25672 (N_25672,N_24650,N_24303);
xnor U25673 (N_25673,N_24622,N_24596);
xor U25674 (N_25674,N_24190,N_24973);
and U25675 (N_25675,N_24456,N_24018);
and U25676 (N_25676,N_24656,N_24580);
and U25677 (N_25677,N_24538,N_24524);
nor U25678 (N_25678,N_24985,N_24045);
nand U25679 (N_25679,N_24534,N_24615);
xor U25680 (N_25680,N_24789,N_24899);
nor U25681 (N_25681,N_24296,N_24772);
xnor U25682 (N_25682,N_24419,N_24391);
nor U25683 (N_25683,N_24186,N_24060);
nor U25684 (N_25684,N_24379,N_24196);
or U25685 (N_25685,N_24653,N_24924);
xnor U25686 (N_25686,N_24615,N_24102);
nand U25687 (N_25687,N_24161,N_24492);
nor U25688 (N_25688,N_24977,N_24748);
nor U25689 (N_25689,N_24077,N_24973);
or U25690 (N_25690,N_24661,N_24685);
nand U25691 (N_25691,N_24533,N_24457);
or U25692 (N_25692,N_24542,N_24174);
nor U25693 (N_25693,N_24131,N_24315);
xor U25694 (N_25694,N_24578,N_24118);
xnor U25695 (N_25695,N_24540,N_24513);
nor U25696 (N_25696,N_24471,N_24309);
and U25697 (N_25697,N_24972,N_24523);
or U25698 (N_25698,N_24077,N_24991);
nor U25699 (N_25699,N_24137,N_24779);
nor U25700 (N_25700,N_24674,N_24064);
xnor U25701 (N_25701,N_24825,N_24009);
xnor U25702 (N_25702,N_24693,N_24291);
nor U25703 (N_25703,N_24489,N_24025);
xor U25704 (N_25704,N_24694,N_24172);
and U25705 (N_25705,N_24765,N_24009);
nor U25706 (N_25706,N_24538,N_24408);
or U25707 (N_25707,N_24732,N_24373);
or U25708 (N_25708,N_24364,N_24250);
and U25709 (N_25709,N_24250,N_24299);
and U25710 (N_25710,N_24248,N_24907);
nor U25711 (N_25711,N_24997,N_24858);
or U25712 (N_25712,N_24958,N_24524);
or U25713 (N_25713,N_24123,N_24696);
or U25714 (N_25714,N_24600,N_24010);
and U25715 (N_25715,N_24040,N_24645);
nand U25716 (N_25716,N_24801,N_24619);
xor U25717 (N_25717,N_24309,N_24887);
or U25718 (N_25718,N_24314,N_24267);
xnor U25719 (N_25719,N_24986,N_24025);
xor U25720 (N_25720,N_24787,N_24847);
xnor U25721 (N_25721,N_24799,N_24480);
and U25722 (N_25722,N_24742,N_24440);
or U25723 (N_25723,N_24178,N_24518);
nand U25724 (N_25724,N_24102,N_24175);
nand U25725 (N_25725,N_24875,N_24892);
and U25726 (N_25726,N_24494,N_24123);
nor U25727 (N_25727,N_24103,N_24351);
xnor U25728 (N_25728,N_24517,N_24656);
nand U25729 (N_25729,N_24702,N_24160);
nor U25730 (N_25730,N_24530,N_24191);
or U25731 (N_25731,N_24136,N_24069);
xor U25732 (N_25732,N_24939,N_24474);
and U25733 (N_25733,N_24741,N_24300);
nor U25734 (N_25734,N_24685,N_24777);
xnor U25735 (N_25735,N_24167,N_24904);
xor U25736 (N_25736,N_24852,N_24314);
nor U25737 (N_25737,N_24592,N_24133);
nor U25738 (N_25738,N_24854,N_24529);
nand U25739 (N_25739,N_24396,N_24188);
nor U25740 (N_25740,N_24727,N_24410);
nor U25741 (N_25741,N_24956,N_24361);
or U25742 (N_25742,N_24785,N_24911);
xnor U25743 (N_25743,N_24949,N_24253);
or U25744 (N_25744,N_24937,N_24387);
nand U25745 (N_25745,N_24581,N_24992);
nor U25746 (N_25746,N_24937,N_24707);
nor U25747 (N_25747,N_24696,N_24632);
nor U25748 (N_25748,N_24439,N_24990);
nand U25749 (N_25749,N_24631,N_24215);
and U25750 (N_25750,N_24527,N_24794);
or U25751 (N_25751,N_24685,N_24261);
or U25752 (N_25752,N_24410,N_24619);
xor U25753 (N_25753,N_24387,N_24169);
and U25754 (N_25754,N_24863,N_24321);
or U25755 (N_25755,N_24115,N_24454);
and U25756 (N_25756,N_24949,N_24214);
xnor U25757 (N_25757,N_24111,N_24146);
and U25758 (N_25758,N_24589,N_24514);
nor U25759 (N_25759,N_24559,N_24312);
nor U25760 (N_25760,N_24128,N_24881);
and U25761 (N_25761,N_24176,N_24450);
and U25762 (N_25762,N_24331,N_24509);
nand U25763 (N_25763,N_24277,N_24799);
and U25764 (N_25764,N_24071,N_24822);
nand U25765 (N_25765,N_24437,N_24124);
xnor U25766 (N_25766,N_24978,N_24074);
nor U25767 (N_25767,N_24538,N_24949);
nor U25768 (N_25768,N_24648,N_24827);
nor U25769 (N_25769,N_24882,N_24500);
or U25770 (N_25770,N_24255,N_24757);
xnor U25771 (N_25771,N_24739,N_24930);
and U25772 (N_25772,N_24062,N_24264);
nand U25773 (N_25773,N_24181,N_24689);
and U25774 (N_25774,N_24474,N_24442);
nor U25775 (N_25775,N_24050,N_24988);
nor U25776 (N_25776,N_24495,N_24561);
nor U25777 (N_25777,N_24210,N_24570);
nor U25778 (N_25778,N_24981,N_24303);
or U25779 (N_25779,N_24455,N_24297);
nor U25780 (N_25780,N_24367,N_24608);
nor U25781 (N_25781,N_24914,N_24452);
and U25782 (N_25782,N_24903,N_24434);
nor U25783 (N_25783,N_24441,N_24384);
nor U25784 (N_25784,N_24856,N_24595);
and U25785 (N_25785,N_24206,N_24134);
and U25786 (N_25786,N_24277,N_24329);
or U25787 (N_25787,N_24383,N_24308);
nor U25788 (N_25788,N_24789,N_24302);
nand U25789 (N_25789,N_24061,N_24815);
xnor U25790 (N_25790,N_24620,N_24423);
xor U25791 (N_25791,N_24480,N_24609);
or U25792 (N_25792,N_24961,N_24971);
xnor U25793 (N_25793,N_24482,N_24558);
and U25794 (N_25794,N_24515,N_24086);
and U25795 (N_25795,N_24761,N_24638);
nor U25796 (N_25796,N_24278,N_24279);
nand U25797 (N_25797,N_24532,N_24365);
xnor U25798 (N_25798,N_24270,N_24179);
nor U25799 (N_25799,N_24119,N_24449);
nor U25800 (N_25800,N_24805,N_24510);
nand U25801 (N_25801,N_24740,N_24102);
nand U25802 (N_25802,N_24482,N_24614);
nand U25803 (N_25803,N_24865,N_24979);
and U25804 (N_25804,N_24172,N_24351);
or U25805 (N_25805,N_24722,N_24123);
and U25806 (N_25806,N_24672,N_24768);
xnor U25807 (N_25807,N_24973,N_24269);
xnor U25808 (N_25808,N_24066,N_24577);
nand U25809 (N_25809,N_24080,N_24716);
nand U25810 (N_25810,N_24188,N_24800);
or U25811 (N_25811,N_24252,N_24506);
nand U25812 (N_25812,N_24287,N_24489);
or U25813 (N_25813,N_24858,N_24104);
nor U25814 (N_25814,N_24640,N_24397);
xnor U25815 (N_25815,N_24050,N_24565);
xor U25816 (N_25816,N_24744,N_24709);
and U25817 (N_25817,N_24892,N_24077);
nor U25818 (N_25818,N_24292,N_24194);
nor U25819 (N_25819,N_24972,N_24434);
nor U25820 (N_25820,N_24728,N_24612);
xnor U25821 (N_25821,N_24255,N_24583);
and U25822 (N_25822,N_24606,N_24521);
or U25823 (N_25823,N_24613,N_24987);
or U25824 (N_25824,N_24675,N_24717);
or U25825 (N_25825,N_24012,N_24431);
nor U25826 (N_25826,N_24119,N_24775);
and U25827 (N_25827,N_24722,N_24865);
xnor U25828 (N_25828,N_24508,N_24556);
nand U25829 (N_25829,N_24933,N_24457);
and U25830 (N_25830,N_24726,N_24962);
xnor U25831 (N_25831,N_24425,N_24483);
nand U25832 (N_25832,N_24470,N_24517);
or U25833 (N_25833,N_24200,N_24687);
xnor U25834 (N_25834,N_24415,N_24361);
xor U25835 (N_25835,N_24514,N_24222);
and U25836 (N_25836,N_24977,N_24031);
nand U25837 (N_25837,N_24324,N_24927);
nor U25838 (N_25838,N_24898,N_24939);
nor U25839 (N_25839,N_24205,N_24768);
nand U25840 (N_25840,N_24110,N_24350);
nand U25841 (N_25841,N_24757,N_24264);
nor U25842 (N_25842,N_24815,N_24797);
nand U25843 (N_25843,N_24353,N_24497);
nand U25844 (N_25844,N_24849,N_24204);
nor U25845 (N_25845,N_24761,N_24774);
and U25846 (N_25846,N_24995,N_24065);
nand U25847 (N_25847,N_24717,N_24704);
or U25848 (N_25848,N_24041,N_24400);
and U25849 (N_25849,N_24358,N_24198);
or U25850 (N_25850,N_24207,N_24521);
nand U25851 (N_25851,N_24789,N_24071);
nor U25852 (N_25852,N_24775,N_24922);
nand U25853 (N_25853,N_24531,N_24201);
and U25854 (N_25854,N_24426,N_24630);
or U25855 (N_25855,N_24737,N_24232);
xor U25856 (N_25856,N_24960,N_24490);
xor U25857 (N_25857,N_24769,N_24176);
nand U25858 (N_25858,N_24430,N_24756);
and U25859 (N_25859,N_24341,N_24031);
xnor U25860 (N_25860,N_24283,N_24894);
nor U25861 (N_25861,N_24133,N_24557);
xor U25862 (N_25862,N_24040,N_24238);
nor U25863 (N_25863,N_24458,N_24904);
and U25864 (N_25864,N_24932,N_24353);
xor U25865 (N_25865,N_24951,N_24842);
nor U25866 (N_25866,N_24338,N_24767);
xor U25867 (N_25867,N_24734,N_24284);
or U25868 (N_25868,N_24941,N_24354);
xor U25869 (N_25869,N_24408,N_24960);
and U25870 (N_25870,N_24635,N_24570);
xnor U25871 (N_25871,N_24803,N_24897);
and U25872 (N_25872,N_24717,N_24911);
nand U25873 (N_25873,N_24380,N_24463);
or U25874 (N_25874,N_24661,N_24672);
xor U25875 (N_25875,N_24184,N_24880);
nor U25876 (N_25876,N_24924,N_24799);
or U25877 (N_25877,N_24388,N_24705);
xnor U25878 (N_25878,N_24614,N_24851);
nor U25879 (N_25879,N_24098,N_24921);
nor U25880 (N_25880,N_24563,N_24119);
or U25881 (N_25881,N_24554,N_24884);
nand U25882 (N_25882,N_24219,N_24937);
nor U25883 (N_25883,N_24571,N_24151);
nor U25884 (N_25884,N_24305,N_24676);
or U25885 (N_25885,N_24972,N_24023);
xnor U25886 (N_25886,N_24257,N_24577);
nand U25887 (N_25887,N_24737,N_24468);
xnor U25888 (N_25888,N_24672,N_24008);
and U25889 (N_25889,N_24695,N_24847);
xnor U25890 (N_25890,N_24794,N_24226);
nand U25891 (N_25891,N_24949,N_24071);
or U25892 (N_25892,N_24560,N_24829);
nor U25893 (N_25893,N_24661,N_24924);
nor U25894 (N_25894,N_24535,N_24607);
xnor U25895 (N_25895,N_24641,N_24578);
xor U25896 (N_25896,N_24204,N_24308);
nor U25897 (N_25897,N_24709,N_24380);
nor U25898 (N_25898,N_24327,N_24598);
nor U25899 (N_25899,N_24135,N_24996);
or U25900 (N_25900,N_24237,N_24885);
nand U25901 (N_25901,N_24845,N_24569);
xnor U25902 (N_25902,N_24502,N_24193);
xnor U25903 (N_25903,N_24549,N_24410);
and U25904 (N_25904,N_24350,N_24109);
nor U25905 (N_25905,N_24136,N_24694);
nand U25906 (N_25906,N_24961,N_24384);
xnor U25907 (N_25907,N_24826,N_24424);
nand U25908 (N_25908,N_24229,N_24534);
xor U25909 (N_25909,N_24428,N_24932);
and U25910 (N_25910,N_24837,N_24244);
nor U25911 (N_25911,N_24035,N_24311);
nand U25912 (N_25912,N_24151,N_24602);
xor U25913 (N_25913,N_24246,N_24931);
nand U25914 (N_25914,N_24486,N_24952);
xnor U25915 (N_25915,N_24606,N_24888);
nand U25916 (N_25916,N_24422,N_24270);
nor U25917 (N_25917,N_24768,N_24371);
xnor U25918 (N_25918,N_24056,N_24882);
nor U25919 (N_25919,N_24511,N_24783);
nand U25920 (N_25920,N_24831,N_24350);
nor U25921 (N_25921,N_24925,N_24443);
or U25922 (N_25922,N_24165,N_24093);
and U25923 (N_25923,N_24358,N_24001);
and U25924 (N_25924,N_24844,N_24161);
and U25925 (N_25925,N_24569,N_24614);
or U25926 (N_25926,N_24762,N_24452);
or U25927 (N_25927,N_24640,N_24743);
nor U25928 (N_25928,N_24402,N_24480);
or U25929 (N_25929,N_24364,N_24709);
nor U25930 (N_25930,N_24960,N_24838);
nand U25931 (N_25931,N_24561,N_24698);
or U25932 (N_25932,N_24261,N_24006);
or U25933 (N_25933,N_24155,N_24159);
nand U25934 (N_25934,N_24721,N_24181);
or U25935 (N_25935,N_24159,N_24567);
and U25936 (N_25936,N_24625,N_24136);
or U25937 (N_25937,N_24503,N_24547);
or U25938 (N_25938,N_24058,N_24756);
and U25939 (N_25939,N_24194,N_24053);
nor U25940 (N_25940,N_24496,N_24473);
and U25941 (N_25941,N_24168,N_24559);
nand U25942 (N_25942,N_24241,N_24035);
nor U25943 (N_25943,N_24832,N_24574);
or U25944 (N_25944,N_24218,N_24484);
nand U25945 (N_25945,N_24532,N_24445);
xor U25946 (N_25946,N_24442,N_24352);
nand U25947 (N_25947,N_24011,N_24350);
and U25948 (N_25948,N_24835,N_24779);
nand U25949 (N_25949,N_24962,N_24572);
nand U25950 (N_25950,N_24256,N_24763);
nand U25951 (N_25951,N_24118,N_24501);
xor U25952 (N_25952,N_24357,N_24048);
and U25953 (N_25953,N_24994,N_24097);
xnor U25954 (N_25954,N_24412,N_24049);
nor U25955 (N_25955,N_24577,N_24270);
nand U25956 (N_25956,N_24911,N_24799);
xor U25957 (N_25957,N_24203,N_24922);
nor U25958 (N_25958,N_24377,N_24323);
or U25959 (N_25959,N_24632,N_24955);
nor U25960 (N_25960,N_24854,N_24577);
nand U25961 (N_25961,N_24144,N_24532);
xnor U25962 (N_25962,N_24675,N_24354);
and U25963 (N_25963,N_24474,N_24062);
nand U25964 (N_25964,N_24901,N_24753);
xor U25965 (N_25965,N_24965,N_24898);
or U25966 (N_25966,N_24830,N_24170);
or U25967 (N_25967,N_24209,N_24063);
xnor U25968 (N_25968,N_24859,N_24199);
and U25969 (N_25969,N_24877,N_24552);
nand U25970 (N_25970,N_24268,N_24468);
and U25971 (N_25971,N_24661,N_24836);
xnor U25972 (N_25972,N_24768,N_24624);
and U25973 (N_25973,N_24135,N_24664);
nor U25974 (N_25974,N_24442,N_24013);
nor U25975 (N_25975,N_24499,N_24746);
xnor U25976 (N_25976,N_24109,N_24278);
xor U25977 (N_25977,N_24698,N_24016);
nor U25978 (N_25978,N_24855,N_24690);
nor U25979 (N_25979,N_24047,N_24194);
nor U25980 (N_25980,N_24808,N_24608);
and U25981 (N_25981,N_24839,N_24408);
or U25982 (N_25982,N_24177,N_24940);
and U25983 (N_25983,N_24746,N_24841);
nor U25984 (N_25984,N_24630,N_24920);
nor U25985 (N_25985,N_24152,N_24764);
nor U25986 (N_25986,N_24563,N_24598);
xor U25987 (N_25987,N_24652,N_24055);
or U25988 (N_25988,N_24049,N_24141);
nor U25989 (N_25989,N_24866,N_24951);
or U25990 (N_25990,N_24971,N_24393);
nand U25991 (N_25991,N_24655,N_24881);
nand U25992 (N_25992,N_24904,N_24570);
or U25993 (N_25993,N_24422,N_24082);
xnor U25994 (N_25994,N_24129,N_24963);
and U25995 (N_25995,N_24980,N_24969);
nand U25996 (N_25996,N_24897,N_24705);
or U25997 (N_25997,N_24277,N_24162);
nand U25998 (N_25998,N_24170,N_24182);
nor U25999 (N_25999,N_24163,N_24503);
nand U26000 (N_26000,N_25136,N_25905);
and U26001 (N_26001,N_25651,N_25412);
nand U26002 (N_26002,N_25237,N_25118);
xor U26003 (N_26003,N_25210,N_25975);
nor U26004 (N_26004,N_25413,N_25102);
and U26005 (N_26005,N_25385,N_25699);
nor U26006 (N_26006,N_25918,N_25092);
nor U26007 (N_26007,N_25979,N_25660);
or U26008 (N_26008,N_25255,N_25420);
or U26009 (N_26009,N_25222,N_25474);
or U26010 (N_26010,N_25125,N_25664);
nand U26011 (N_26011,N_25545,N_25005);
xor U26012 (N_26012,N_25151,N_25642);
xor U26013 (N_26013,N_25869,N_25688);
nor U26014 (N_26014,N_25386,N_25910);
and U26015 (N_26015,N_25819,N_25944);
or U26016 (N_26016,N_25206,N_25393);
nand U26017 (N_26017,N_25579,N_25309);
or U26018 (N_26018,N_25761,N_25695);
nor U26019 (N_26019,N_25959,N_25707);
nand U26020 (N_26020,N_25185,N_25725);
nor U26021 (N_26021,N_25552,N_25609);
nor U26022 (N_26022,N_25266,N_25229);
or U26023 (N_26023,N_25416,N_25879);
nor U26024 (N_26024,N_25328,N_25826);
nor U26025 (N_26025,N_25011,N_25339);
or U26026 (N_26026,N_25320,N_25631);
xor U26027 (N_26027,N_25949,N_25331);
nand U26028 (N_26028,N_25227,N_25506);
nor U26029 (N_26029,N_25862,N_25738);
nand U26030 (N_26030,N_25257,N_25865);
and U26031 (N_26031,N_25219,N_25265);
or U26032 (N_26032,N_25193,N_25742);
nand U26033 (N_26033,N_25499,N_25459);
nor U26034 (N_26034,N_25704,N_25403);
or U26035 (N_26035,N_25055,N_25659);
and U26036 (N_26036,N_25252,N_25716);
xor U26037 (N_26037,N_25964,N_25850);
nor U26038 (N_26038,N_25717,N_25596);
and U26039 (N_26039,N_25757,N_25358);
nand U26040 (N_26040,N_25480,N_25076);
and U26041 (N_26041,N_25890,N_25736);
xor U26042 (N_26042,N_25468,N_25566);
and U26043 (N_26043,N_25851,N_25250);
nand U26044 (N_26044,N_25685,N_25999);
or U26045 (N_26045,N_25238,N_25967);
nor U26046 (N_26046,N_25556,N_25275);
or U26047 (N_26047,N_25713,N_25251);
or U26048 (N_26048,N_25604,N_25426);
and U26049 (N_26049,N_25079,N_25876);
and U26050 (N_26050,N_25923,N_25810);
and U26051 (N_26051,N_25855,N_25772);
and U26052 (N_26052,N_25111,N_25859);
xor U26053 (N_26053,N_25505,N_25900);
and U26054 (N_26054,N_25202,N_25268);
or U26055 (N_26055,N_25560,N_25315);
nand U26056 (N_26056,N_25883,N_25470);
xnor U26057 (N_26057,N_25754,N_25313);
nor U26058 (N_26058,N_25832,N_25952);
and U26059 (N_26059,N_25798,N_25588);
nand U26060 (N_26060,N_25316,N_25849);
xor U26061 (N_26061,N_25698,N_25948);
xor U26062 (N_26062,N_25510,N_25517);
nor U26063 (N_26063,N_25198,N_25035);
and U26064 (N_26064,N_25475,N_25931);
xor U26065 (N_26065,N_25149,N_25686);
nor U26066 (N_26066,N_25308,N_25196);
and U26067 (N_26067,N_25167,N_25383);
and U26068 (N_26068,N_25260,N_25042);
or U26069 (N_26069,N_25902,N_25899);
xnor U26070 (N_26070,N_25435,N_25155);
and U26071 (N_26071,N_25954,N_25414);
xnor U26072 (N_26072,N_25981,N_25113);
nor U26073 (N_26073,N_25858,N_25710);
nor U26074 (N_26074,N_25719,N_25903);
xor U26075 (N_26075,N_25546,N_25187);
nand U26076 (N_26076,N_25683,N_25303);
xnor U26077 (N_26077,N_25771,N_25195);
or U26078 (N_26078,N_25019,N_25735);
or U26079 (N_26079,N_25289,N_25933);
xnor U26080 (N_26080,N_25008,N_25535);
and U26081 (N_26081,N_25301,N_25971);
or U26082 (N_26082,N_25992,N_25613);
nand U26083 (N_26083,N_25365,N_25796);
and U26084 (N_26084,N_25818,N_25321);
and U26085 (N_26085,N_25286,N_25569);
xnor U26086 (N_26086,N_25225,N_25681);
or U26087 (N_26087,N_25956,N_25715);
or U26088 (N_26088,N_25955,N_25188);
nand U26089 (N_26089,N_25951,N_25564);
nand U26090 (N_26090,N_25084,N_25878);
xnor U26091 (N_26091,N_25128,N_25839);
nand U26092 (N_26092,N_25075,N_25370);
nand U26093 (N_26093,N_25728,N_25082);
nand U26094 (N_26094,N_25423,N_25670);
nand U26095 (N_26095,N_25484,N_25373);
and U26096 (N_26096,N_25846,N_25354);
nand U26097 (N_26097,N_25443,N_25086);
nand U26098 (N_26098,N_25473,N_25823);
or U26099 (N_26099,N_25067,N_25993);
and U26100 (N_26100,N_25124,N_25371);
nand U26101 (N_26101,N_25091,N_25665);
nand U26102 (N_26102,N_25610,N_25132);
or U26103 (N_26103,N_25534,N_25921);
or U26104 (N_26104,N_25165,N_25802);
nand U26105 (N_26105,N_25244,N_25750);
and U26106 (N_26106,N_25840,N_25580);
nor U26107 (N_26107,N_25957,N_25848);
and U26108 (N_26108,N_25307,N_25114);
nor U26109 (N_26109,N_25319,N_25976);
nand U26110 (N_26110,N_25489,N_25197);
xnor U26111 (N_26111,N_25411,N_25372);
and U26112 (N_26112,N_25752,N_25016);
nand U26113 (N_26113,N_25392,N_25290);
or U26114 (N_26114,N_25362,N_25540);
or U26115 (N_26115,N_25432,N_25162);
and U26116 (N_26116,N_25551,N_25628);
xor U26117 (N_26117,N_25523,N_25213);
and U26118 (N_26118,N_25083,N_25504);
nor U26119 (N_26119,N_25494,N_25943);
xnor U26120 (N_26120,N_25996,N_25749);
and U26121 (N_26121,N_25936,N_25418);
xor U26122 (N_26122,N_25287,N_25778);
nand U26123 (N_26123,N_25003,N_25051);
xor U26124 (N_26124,N_25577,N_25336);
nor U26125 (N_26125,N_25602,N_25767);
or U26126 (N_26126,N_25253,N_25325);
xor U26127 (N_26127,N_25182,N_25679);
xnor U26128 (N_26128,N_25029,N_25882);
nand U26129 (N_26129,N_25820,N_25015);
nor U26130 (N_26130,N_25333,N_25929);
nand U26131 (N_26131,N_25916,N_25205);
and U26132 (N_26132,N_25740,N_25201);
nand U26133 (N_26133,N_25288,N_25199);
or U26134 (N_26134,N_25074,N_25998);
and U26135 (N_26135,N_25745,N_25984);
and U26136 (N_26136,N_25822,N_25300);
and U26137 (N_26137,N_25207,N_25421);
and U26138 (N_26138,N_25977,N_25583);
nor U26139 (N_26139,N_25396,N_25834);
and U26140 (N_26140,N_25001,N_25041);
nor U26141 (N_26141,N_25511,N_25471);
nand U26142 (N_26142,N_25060,N_25892);
or U26143 (N_26143,N_25962,N_25980);
and U26144 (N_26144,N_25166,N_25478);
nor U26145 (N_26145,N_25764,N_25747);
and U26146 (N_26146,N_25842,N_25053);
nand U26147 (N_26147,N_25490,N_25397);
nand U26148 (N_26148,N_25438,N_25753);
or U26149 (N_26149,N_25920,N_25226);
and U26150 (N_26150,N_25389,N_25142);
or U26151 (N_26151,N_25040,N_25700);
xnor U26152 (N_26152,N_25024,N_25705);
nor U26153 (N_26153,N_25284,N_25089);
nand U26154 (N_26154,N_25632,N_25110);
xnor U26155 (N_26155,N_25530,N_25326);
xnor U26156 (N_26156,N_25230,N_25827);
xor U26157 (N_26157,N_25542,N_25374);
nand U26158 (N_26158,N_25769,N_25417);
nor U26159 (N_26159,N_25756,N_25381);
nor U26160 (N_26160,N_25612,N_25746);
nand U26161 (N_26161,N_25183,N_25050);
nor U26162 (N_26162,N_25495,N_25472);
and U26163 (N_26163,N_25800,N_25486);
and U26164 (N_26164,N_25653,N_25901);
xor U26165 (N_26165,N_25158,N_25160);
nor U26166 (N_26166,N_25061,N_25805);
nand U26167 (N_26167,N_25345,N_25267);
nor U26168 (N_26168,N_25240,N_25570);
or U26169 (N_26169,N_25312,N_25018);
and U26170 (N_26170,N_25231,N_25938);
and U26171 (N_26171,N_25963,N_25871);
nor U26172 (N_26172,N_25584,N_25279);
and U26173 (N_26173,N_25550,N_25518);
nand U26174 (N_26174,N_25191,N_25232);
xnor U26175 (N_26175,N_25242,N_25821);
nor U26176 (N_26176,N_25483,N_25675);
or U26177 (N_26177,N_25965,N_25533);
nand U26178 (N_26178,N_25282,N_25452);
or U26179 (N_26179,N_25898,N_25816);
or U26180 (N_26180,N_25002,N_25112);
or U26181 (N_26181,N_25982,N_25991);
nand U26182 (N_26182,N_25406,N_25626);
nor U26183 (N_26183,N_25007,N_25776);
or U26184 (N_26184,N_25450,N_25594);
nor U26185 (N_26185,N_25678,N_25857);
xor U26186 (N_26186,N_25927,N_25448);
xor U26187 (N_26187,N_25455,N_25164);
xor U26188 (N_26188,N_25721,N_25147);
nor U26189 (N_26189,N_25513,N_25638);
and U26190 (N_26190,N_25697,N_25031);
or U26191 (N_26191,N_25507,N_25578);
xnor U26192 (N_26192,N_25152,N_25509);
or U26193 (N_26193,N_25572,N_25274);
or U26194 (N_26194,N_25378,N_25127);
and U26195 (N_26195,N_25223,N_25028);
nor U26196 (N_26196,N_25236,N_25220);
xnor U26197 (N_26197,N_25906,N_25622);
nor U26198 (N_26198,N_25937,N_25972);
and U26199 (N_26199,N_25945,N_25586);
nand U26200 (N_26200,N_25677,N_25911);
xor U26201 (N_26201,N_25794,N_25885);
and U26202 (N_26202,N_25693,N_25590);
or U26203 (N_26203,N_25669,N_25329);
and U26204 (N_26204,N_25843,N_25496);
xnor U26205 (N_26205,N_25405,N_25732);
or U26206 (N_26206,N_25817,N_25272);
nand U26207 (N_26207,N_25856,N_25743);
nor U26208 (N_26208,N_25310,N_25744);
xnor U26209 (N_26209,N_25457,N_25139);
xnor U26210 (N_26210,N_25515,N_25200);
and U26211 (N_26211,N_25658,N_25758);
xor U26212 (N_26212,N_25722,N_25741);
nor U26213 (N_26213,N_25652,N_25379);
or U26214 (N_26214,N_25481,N_25498);
xnor U26215 (N_26215,N_25332,N_25433);
and U26216 (N_26216,N_25808,N_25881);
and U26217 (N_26217,N_25718,N_25825);
or U26218 (N_26218,N_25294,N_25514);
nand U26219 (N_26219,N_25330,N_25145);
xor U26220 (N_26220,N_25595,N_25441);
nand U26221 (N_26221,N_25368,N_25787);
xnor U26222 (N_26222,N_25585,N_25607);
and U26223 (N_26223,N_25059,N_25347);
or U26224 (N_26224,N_25922,N_25000);
or U26225 (N_26225,N_25844,N_25711);
nand U26226 (N_26226,N_25046,N_25960);
and U26227 (N_26227,N_25341,N_25476);
and U26228 (N_26228,N_25235,N_25904);
or U26229 (N_26229,N_25208,N_25647);
nor U26230 (N_26230,N_25502,N_25487);
and U26231 (N_26231,N_25941,N_25360);
xor U26232 (N_26232,N_25926,N_25045);
and U26233 (N_26233,N_25968,N_25702);
and U26234 (N_26234,N_25872,N_25305);
and U26235 (N_26235,N_25215,N_25762);
or U26236 (N_26236,N_25655,N_25343);
xor U26237 (N_26237,N_25380,N_25701);
nor U26238 (N_26238,N_25121,N_25995);
or U26239 (N_26239,N_25759,N_25317);
xor U26240 (N_26240,N_25140,N_25549);
xor U26241 (N_26241,N_25465,N_25204);
and U26242 (N_26242,N_25302,N_25088);
nor U26243 (N_26243,N_25726,N_25010);
nor U26244 (N_26244,N_25430,N_25667);
and U26245 (N_26245,N_25346,N_25439);
xor U26246 (N_26246,N_25589,N_25806);
nor U26247 (N_26247,N_25344,N_25367);
and U26248 (N_26248,N_25617,N_25212);
or U26249 (N_26249,N_25841,N_25587);
nor U26250 (N_26250,N_25217,N_25168);
nand U26251 (N_26251,N_25928,N_25099);
nand U26252 (N_26252,N_25836,N_25845);
and U26253 (N_26253,N_25256,N_25179);
or U26254 (N_26254,N_25123,N_25243);
nor U26255 (N_26255,N_25668,N_25064);
xnor U26256 (N_26256,N_25134,N_25780);
or U26257 (N_26257,N_25500,N_25304);
nor U26258 (N_26258,N_25233,N_25241);
and U26259 (N_26259,N_25946,N_25097);
nand U26260 (N_26260,N_25234,N_25966);
xor U26261 (N_26261,N_25676,N_25209);
xnor U26262 (N_26262,N_25706,N_25065);
or U26263 (N_26263,N_25690,N_25571);
nor U26264 (N_26264,N_25461,N_25449);
nor U26265 (N_26265,N_25184,N_25884);
nor U26266 (N_26266,N_25627,N_25751);
nand U26267 (N_26267,N_25431,N_25391);
nor U26268 (N_26268,N_25090,N_25864);
and U26269 (N_26269,N_25625,N_25529);
nand U26270 (N_26270,N_25526,N_25190);
nand U26271 (N_26271,N_25327,N_25792);
nand U26272 (N_26272,N_25565,N_25342);
or U26273 (N_26273,N_25171,N_25763);
xnor U26274 (N_26274,N_25323,N_25833);
or U26275 (N_26275,N_25122,N_25974);
nor U26276 (N_26276,N_25352,N_25245);
nand U26277 (N_26277,N_25157,N_25755);
and U26278 (N_26278,N_25666,N_25297);
nand U26279 (N_26279,N_25643,N_25056);
and U26280 (N_26280,N_25961,N_25174);
nand U26281 (N_26281,N_25394,N_25618);
nand U26282 (N_26282,N_25043,N_25491);
nor U26283 (N_26283,N_25630,N_25852);
xnor U26284 (N_26284,N_25508,N_25004);
and U26285 (N_26285,N_25356,N_25703);
nor U26286 (N_26286,N_25692,N_25069);
nand U26287 (N_26287,N_25338,N_25285);
nor U26288 (N_26288,N_25645,N_25770);
or U26289 (N_26289,N_25674,N_25605);
xnor U26290 (N_26290,N_25034,N_25488);
xor U26291 (N_26291,N_25913,N_25314);
nand U26292 (N_26292,N_25154,N_25427);
nand U26293 (N_26293,N_25614,N_25942);
nand U26294 (N_26294,N_25646,N_25311);
nand U26295 (N_26295,N_25192,N_25657);
xnor U26296 (N_26296,N_25057,N_25072);
xnor U26297 (N_26297,N_25477,N_25654);
nand U26298 (N_26298,N_25246,N_25791);
nand U26299 (N_26299,N_25661,N_25887);
and U26300 (N_26300,N_25785,N_25860);
or U26301 (N_26301,N_25582,N_25033);
nand U26302 (N_26302,N_25137,N_25634);
and U26303 (N_26303,N_25425,N_25958);
xor U26304 (N_26304,N_25538,N_25765);
or U26305 (N_26305,N_25177,N_25989);
nor U26306 (N_26306,N_25181,N_25548);
nand U26307 (N_26307,N_25983,N_25077);
and U26308 (N_26308,N_25708,N_25847);
nor U26309 (N_26309,N_25886,N_25663);
nand U26310 (N_26310,N_25434,N_25214);
and U26311 (N_26311,N_25611,N_25880);
and U26312 (N_26312,N_25531,N_25485);
or U26313 (N_26313,N_25115,N_25335);
and U26314 (N_26314,N_25044,N_25720);
nand U26315 (N_26315,N_25429,N_25276);
nand U26316 (N_26316,N_25760,N_25953);
nor U26317 (N_26317,N_25621,N_25349);
nor U26318 (N_26318,N_25135,N_25013);
or U26319 (N_26319,N_25264,N_25422);
nand U26320 (N_26320,N_25153,N_25462);
and U26321 (N_26321,N_25078,N_25131);
xor U26322 (N_26322,N_25873,N_25175);
nand U26323 (N_26323,N_25624,N_25599);
or U26324 (N_26324,N_25896,N_25100);
and U26325 (N_26325,N_25436,N_25066);
xor U26326 (N_26326,N_25891,N_25568);
nand U26327 (N_26327,N_25442,N_25159);
or U26328 (N_26328,N_25440,N_25262);
or U26329 (N_26329,N_25247,N_25203);
and U26330 (N_26330,N_25080,N_25463);
nand U26331 (N_26331,N_25334,N_25593);
nor U26332 (N_26332,N_25133,N_25451);
nand U26333 (N_26333,N_25801,N_25789);
xor U26334 (N_26334,N_25512,N_25553);
nor U26335 (N_26335,N_25466,N_25867);
nor U26336 (N_26336,N_25039,N_25464);
xor U26337 (N_26337,N_25934,N_25493);
and U26338 (N_26338,N_25062,N_25623);
nor U26339 (N_26339,N_25444,N_25469);
nand U26340 (N_26340,N_25914,N_25375);
nand U26341 (N_26341,N_25592,N_25786);
nand U26342 (N_26342,N_25835,N_25536);
nand U26343 (N_26343,N_25635,N_25619);
or U26344 (N_26344,N_25804,N_25576);
xor U26345 (N_26345,N_25415,N_25216);
and U26346 (N_26346,N_25729,N_25454);
or U26347 (N_26347,N_25598,N_25637);
or U26348 (N_26348,N_25388,N_25293);
nor U26349 (N_26349,N_25574,N_25146);
and U26350 (N_26350,N_25012,N_25516);
nand U26351 (N_26351,N_25837,N_25603);
xor U26352 (N_26352,N_25799,N_25723);
and U26353 (N_26353,N_25988,N_25909);
nor U26354 (N_26354,N_25456,N_25492);
nand U26355 (N_26355,N_25813,N_25273);
and U26356 (N_26356,N_25528,N_25384);
or U26357 (N_26357,N_25969,N_25978);
or U26358 (N_26358,N_25912,N_25793);
or U26359 (N_26359,N_25739,N_25520);
xor U26360 (N_26360,N_25271,N_25866);
nand U26361 (N_26361,N_25254,N_25648);
nand U26362 (N_26362,N_25052,N_25877);
nand U26363 (N_26363,N_25337,N_25712);
and U26364 (N_26364,N_25156,N_25689);
nand U26365 (N_26365,N_25119,N_25795);
or U26366 (N_26366,N_25616,N_25437);
xnor U26367 (N_26367,N_25006,N_25782);
xnor U26368 (N_26368,N_25809,N_25567);
xnor U26369 (N_26369,N_25063,N_25298);
nor U26370 (N_26370,N_25357,N_25283);
nand U26371 (N_26371,N_25126,N_25355);
nor U26372 (N_26372,N_25709,N_25400);
nand U26373 (N_26373,N_25054,N_25221);
or U26374 (N_26374,N_25985,N_25460);
nand U26375 (N_26375,N_25169,N_25636);
nor U26376 (N_26376,N_25557,N_25503);
nor U26377 (N_26377,N_25875,N_25562);
and U26378 (N_26378,N_25094,N_25853);
or U26379 (N_26379,N_25037,N_25453);
xnor U26380 (N_26380,N_25522,N_25278);
nand U26381 (N_26381,N_25218,N_25779);
nand U26382 (N_26382,N_25032,N_25970);
nor U26383 (N_26383,N_25306,N_25376);
nand U26384 (N_26384,N_25684,N_25608);
or U26385 (N_26385,N_25020,N_25694);
nor U26386 (N_26386,N_25211,N_25364);
xor U26387 (N_26387,N_25138,N_25724);
or U26388 (N_26388,N_25730,N_25532);
nor U26389 (N_26389,N_25714,N_25258);
nand U26390 (N_26390,N_25893,N_25408);
and U26391 (N_26391,N_25363,N_25398);
nand U26392 (N_26392,N_25543,N_25629);
nor U26393 (N_26393,N_25009,N_25829);
nand U26394 (N_26394,N_25854,N_25095);
xor U26395 (N_26395,N_25919,N_25986);
nand U26396 (N_26396,N_25402,N_25939);
or U26397 (N_26397,N_25807,N_25924);
or U26398 (N_26398,N_25047,N_25351);
nand U26399 (N_26399,N_25527,N_25073);
and U26400 (N_26400,N_25561,N_25087);
nor U26401 (N_26401,N_25680,N_25925);
xor U26402 (N_26402,N_25682,N_25130);
nor U26403 (N_26403,N_25117,N_25537);
and U26404 (N_26404,N_25105,N_25650);
nand U26405 (N_26405,N_25525,N_25868);
nand U26406 (N_26406,N_25501,N_25048);
or U26407 (N_26407,N_25521,N_25737);
nand U26408 (N_26408,N_25777,N_25194);
and U26409 (N_26409,N_25014,N_25322);
or U26410 (N_26410,N_25458,N_25824);
xor U26411 (N_26411,N_25781,N_25103);
or U26412 (N_26412,N_25620,N_25555);
and U26413 (N_26413,N_25098,N_25591);
and U26414 (N_26414,N_25990,N_25861);
nor U26415 (N_26415,N_25120,N_25030);
xor U26416 (N_26416,N_25895,N_25559);
nor U26417 (N_26417,N_25811,N_25409);
nor U26418 (N_26418,N_25144,N_25870);
and U26419 (N_26419,N_25017,N_25539);
nand U26420 (N_26420,N_25022,N_25994);
xnor U26421 (N_26421,N_25148,N_25025);
or U26422 (N_26422,N_25143,N_25377);
nand U26423 (N_26423,N_25997,N_25382);
or U26424 (N_26424,N_25270,N_25224);
nor U26425 (N_26425,N_25831,N_25601);
xor U26426 (N_26426,N_25973,N_25324);
nor U26427 (N_26427,N_25897,N_25178);
and U26428 (N_26428,N_25812,N_25987);
nor U26429 (N_26429,N_25186,N_25068);
or U26430 (N_26430,N_25889,N_25172);
nand U26431 (N_26431,N_25830,N_25366);
and U26432 (N_26432,N_25445,N_25691);
and U26433 (N_26433,N_25269,N_25350);
xor U26434 (N_26434,N_25519,N_25150);
nand U26435 (N_26435,N_25399,N_25296);
xor U26436 (N_26436,N_25774,N_25907);
or U26437 (N_26437,N_25615,N_25874);
nand U26438 (N_26438,N_25387,N_25482);
xor U26439 (N_26439,N_25597,N_25248);
or U26440 (N_26440,N_25395,N_25673);
or U26441 (N_26441,N_25915,N_25259);
xor U26442 (N_26442,N_25239,N_25662);
xnor U26443 (N_26443,N_25106,N_25930);
nand U26444 (N_26444,N_25173,N_25544);
xor U26445 (N_26445,N_25116,N_25803);
or U26446 (N_26446,N_25581,N_25263);
nor U26447 (N_26447,N_25775,N_25606);
and U26448 (N_26448,N_25163,N_25547);
xor U26449 (N_26449,N_25467,N_25295);
and U26450 (N_26450,N_25640,N_25541);
or U26451 (N_26451,N_25348,N_25731);
xor U26452 (N_26452,N_25071,N_25291);
nor U26453 (N_26453,N_25249,N_25096);
nor U26454 (N_26454,N_25558,N_25733);
or U26455 (N_26455,N_25277,N_25081);
nor U26456 (N_26456,N_25497,N_25180);
or U26457 (N_26457,N_25639,N_25672);
xor U26458 (N_26458,N_25563,N_25108);
xor U26459 (N_26459,N_25036,N_25292);
xnor U26460 (N_26460,N_25633,N_25390);
or U26461 (N_26461,N_25940,N_25917);
xnor U26462 (N_26462,N_25107,N_25353);
xor U26463 (N_26463,N_25023,N_25404);
nand U26464 (N_26464,N_25687,N_25109);
nand U26465 (N_26465,N_25407,N_25170);
nor U26466 (N_26466,N_25734,N_25299);
xor U26467 (N_26467,N_25788,N_25021);
nand U26468 (N_26468,N_25671,N_25189);
nor U26469 (N_26469,N_25768,N_25790);
or U26470 (N_26470,N_25828,N_25554);
nor U26471 (N_26471,N_25410,N_25058);
nand U26472 (N_26472,N_25908,N_25318);
and U26473 (N_26473,N_25784,N_25093);
or U26474 (N_26474,N_25141,N_25261);
nand U26475 (N_26475,N_25026,N_25369);
xnor U26476 (N_26476,N_25524,N_25727);
or U26477 (N_26477,N_25038,N_25947);
nand U26478 (N_26478,N_25340,N_25176);
and U26479 (N_26479,N_25101,N_25656);
nand U26480 (N_26480,N_25428,N_25838);
nand U26481 (N_26481,N_25027,N_25401);
or U26482 (N_26482,N_25894,N_25575);
xor U26483 (N_26483,N_25950,N_25104);
or U26484 (N_26484,N_25696,N_25641);
or U26485 (N_26485,N_25359,N_25748);
or U26486 (N_26486,N_25773,N_25573);
nand U26487 (N_26487,N_25085,N_25649);
nand U26488 (N_26488,N_25280,N_25783);
xor U26489 (N_26489,N_25935,N_25888);
and U26490 (N_26490,N_25814,N_25932);
nand U26491 (N_26491,N_25228,N_25447);
and U26492 (N_26492,N_25129,N_25419);
xor U26493 (N_26493,N_25161,N_25766);
nor U26494 (N_26494,N_25446,N_25797);
xor U26495 (N_26495,N_25600,N_25424);
nor U26496 (N_26496,N_25644,N_25479);
nor U26497 (N_26497,N_25070,N_25049);
nor U26498 (N_26498,N_25281,N_25361);
nand U26499 (N_26499,N_25815,N_25863);
nor U26500 (N_26500,N_25540,N_25559);
and U26501 (N_26501,N_25315,N_25543);
xor U26502 (N_26502,N_25842,N_25182);
or U26503 (N_26503,N_25364,N_25295);
and U26504 (N_26504,N_25675,N_25682);
and U26505 (N_26505,N_25024,N_25561);
nand U26506 (N_26506,N_25101,N_25555);
nor U26507 (N_26507,N_25384,N_25223);
nand U26508 (N_26508,N_25720,N_25619);
nand U26509 (N_26509,N_25839,N_25833);
nand U26510 (N_26510,N_25808,N_25524);
and U26511 (N_26511,N_25361,N_25441);
nor U26512 (N_26512,N_25432,N_25525);
xnor U26513 (N_26513,N_25772,N_25258);
nand U26514 (N_26514,N_25936,N_25604);
nand U26515 (N_26515,N_25721,N_25978);
nor U26516 (N_26516,N_25109,N_25400);
nand U26517 (N_26517,N_25997,N_25935);
and U26518 (N_26518,N_25214,N_25616);
nor U26519 (N_26519,N_25674,N_25818);
nor U26520 (N_26520,N_25310,N_25994);
nand U26521 (N_26521,N_25703,N_25447);
or U26522 (N_26522,N_25125,N_25035);
nor U26523 (N_26523,N_25550,N_25880);
or U26524 (N_26524,N_25028,N_25394);
or U26525 (N_26525,N_25390,N_25384);
xnor U26526 (N_26526,N_25160,N_25622);
nand U26527 (N_26527,N_25428,N_25511);
nand U26528 (N_26528,N_25602,N_25466);
and U26529 (N_26529,N_25383,N_25605);
xor U26530 (N_26530,N_25841,N_25690);
or U26531 (N_26531,N_25491,N_25155);
nand U26532 (N_26532,N_25314,N_25797);
nor U26533 (N_26533,N_25899,N_25415);
nor U26534 (N_26534,N_25443,N_25752);
nor U26535 (N_26535,N_25699,N_25574);
xor U26536 (N_26536,N_25655,N_25003);
xnor U26537 (N_26537,N_25536,N_25094);
or U26538 (N_26538,N_25691,N_25534);
or U26539 (N_26539,N_25026,N_25455);
or U26540 (N_26540,N_25021,N_25982);
or U26541 (N_26541,N_25036,N_25172);
or U26542 (N_26542,N_25642,N_25640);
xnor U26543 (N_26543,N_25619,N_25086);
nor U26544 (N_26544,N_25646,N_25095);
or U26545 (N_26545,N_25462,N_25062);
and U26546 (N_26546,N_25262,N_25350);
or U26547 (N_26547,N_25144,N_25914);
and U26548 (N_26548,N_25634,N_25477);
and U26549 (N_26549,N_25930,N_25679);
nor U26550 (N_26550,N_25663,N_25627);
xnor U26551 (N_26551,N_25811,N_25303);
nor U26552 (N_26552,N_25493,N_25196);
and U26553 (N_26553,N_25563,N_25103);
xor U26554 (N_26554,N_25838,N_25156);
nand U26555 (N_26555,N_25394,N_25388);
or U26556 (N_26556,N_25411,N_25783);
or U26557 (N_26557,N_25355,N_25182);
and U26558 (N_26558,N_25208,N_25603);
nor U26559 (N_26559,N_25543,N_25926);
and U26560 (N_26560,N_25954,N_25857);
nand U26561 (N_26561,N_25243,N_25573);
xor U26562 (N_26562,N_25730,N_25750);
and U26563 (N_26563,N_25818,N_25573);
xor U26564 (N_26564,N_25697,N_25374);
nor U26565 (N_26565,N_25787,N_25804);
nor U26566 (N_26566,N_25407,N_25193);
or U26567 (N_26567,N_25469,N_25615);
and U26568 (N_26568,N_25349,N_25213);
nor U26569 (N_26569,N_25367,N_25947);
nor U26570 (N_26570,N_25161,N_25974);
xor U26571 (N_26571,N_25619,N_25096);
nand U26572 (N_26572,N_25886,N_25200);
nand U26573 (N_26573,N_25927,N_25053);
xor U26574 (N_26574,N_25343,N_25667);
or U26575 (N_26575,N_25857,N_25849);
nand U26576 (N_26576,N_25939,N_25071);
or U26577 (N_26577,N_25474,N_25144);
and U26578 (N_26578,N_25128,N_25753);
xnor U26579 (N_26579,N_25116,N_25945);
nand U26580 (N_26580,N_25912,N_25382);
and U26581 (N_26581,N_25934,N_25725);
xnor U26582 (N_26582,N_25133,N_25252);
or U26583 (N_26583,N_25380,N_25526);
nor U26584 (N_26584,N_25353,N_25963);
nand U26585 (N_26585,N_25314,N_25980);
nor U26586 (N_26586,N_25635,N_25186);
nand U26587 (N_26587,N_25109,N_25355);
or U26588 (N_26588,N_25032,N_25403);
nor U26589 (N_26589,N_25826,N_25465);
nand U26590 (N_26590,N_25681,N_25831);
xor U26591 (N_26591,N_25134,N_25046);
xnor U26592 (N_26592,N_25706,N_25834);
nand U26593 (N_26593,N_25571,N_25420);
nand U26594 (N_26594,N_25545,N_25133);
and U26595 (N_26595,N_25671,N_25505);
nor U26596 (N_26596,N_25966,N_25191);
nand U26597 (N_26597,N_25118,N_25861);
nor U26598 (N_26598,N_25347,N_25656);
xnor U26599 (N_26599,N_25415,N_25543);
xor U26600 (N_26600,N_25821,N_25263);
and U26601 (N_26601,N_25449,N_25282);
or U26602 (N_26602,N_25814,N_25012);
xor U26603 (N_26603,N_25699,N_25407);
and U26604 (N_26604,N_25224,N_25654);
nand U26605 (N_26605,N_25405,N_25396);
nor U26606 (N_26606,N_25989,N_25147);
and U26607 (N_26607,N_25518,N_25162);
nor U26608 (N_26608,N_25411,N_25490);
or U26609 (N_26609,N_25329,N_25211);
or U26610 (N_26610,N_25847,N_25936);
or U26611 (N_26611,N_25965,N_25125);
xnor U26612 (N_26612,N_25568,N_25128);
and U26613 (N_26613,N_25594,N_25348);
nor U26614 (N_26614,N_25004,N_25415);
nand U26615 (N_26615,N_25117,N_25251);
xnor U26616 (N_26616,N_25624,N_25333);
xnor U26617 (N_26617,N_25997,N_25741);
and U26618 (N_26618,N_25980,N_25935);
nand U26619 (N_26619,N_25438,N_25234);
and U26620 (N_26620,N_25568,N_25925);
nor U26621 (N_26621,N_25080,N_25945);
and U26622 (N_26622,N_25937,N_25741);
and U26623 (N_26623,N_25028,N_25971);
and U26624 (N_26624,N_25850,N_25555);
or U26625 (N_26625,N_25231,N_25777);
nor U26626 (N_26626,N_25964,N_25436);
and U26627 (N_26627,N_25380,N_25691);
and U26628 (N_26628,N_25937,N_25112);
nor U26629 (N_26629,N_25367,N_25676);
or U26630 (N_26630,N_25204,N_25093);
xor U26631 (N_26631,N_25497,N_25920);
nor U26632 (N_26632,N_25079,N_25341);
or U26633 (N_26633,N_25896,N_25594);
and U26634 (N_26634,N_25497,N_25696);
nor U26635 (N_26635,N_25274,N_25081);
and U26636 (N_26636,N_25484,N_25791);
and U26637 (N_26637,N_25358,N_25713);
or U26638 (N_26638,N_25985,N_25156);
and U26639 (N_26639,N_25581,N_25201);
or U26640 (N_26640,N_25822,N_25667);
xnor U26641 (N_26641,N_25194,N_25916);
nand U26642 (N_26642,N_25870,N_25861);
xor U26643 (N_26643,N_25812,N_25266);
nand U26644 (N_26644,N_25472,N_25769);
nor U26645 (N_26645,N_25383,N_25077);
nand U26646 (N_26646,N_25610,N_25301);
nand U26647 (N_26647,N_25032,N_25451);
or U26648 (N_26648,N_25151,N_25402);
nand U26649 (N_26649,N_25367,N_25511);
nor U26650 (N_26650,N_25581,N_25380);
or U26651 (N_26651,N_25403,N_25745);
and U26652 (N_26652,N_25829,N_25289);
nand U26653 (N_26653,N_25610,N_25102);
nand U26654 (N_26654,N_25744,N_25547);
and U26655 (N_26655,N_25125,N_25645);
nor U26656 (N_26656,N_25998,N_25899);
xnor U26657 (N_26657,N_25079,N_25836);
and U26658 (N_26658,N_25342,N_25987);
xnor U26659 (N_26659,N_25574,N_25881);
or U26660 (N_26660,N_25528,N_25569);
or U26661 (N_26661,N_25660,N_25363);
xor U26662 (N_26662,N_25319,N_25225);
nor U26663 (N_26663,N_25413,N_25590);
nand U26664 (N_26664,N_25360,N_25604);
nor U26665 (N_26665,N_25199,N_25365);
nand U26666 (N_26666,N_25742,N_25632);
nor U26667 (N_26667,N_25348,N_25209);
nand U26668 (N_26668,N_25752,N_25954);
nand U26669 (N_26669,N_25413,N_25380);
xor U26670 (N_26670,N_25017,N_25368);
nor U26671 (N_26671,N_25519,N_25959);
or U26672 (N_26672,N_25571,N_25611);
nor U26673 (N_26673,N_25884,N_25679);
and U26674 (N_26674,N_25303,N_25436);
or U26675 (N_26675,N_25680,N_25462);
and U26676 (N_26676,N_25767,N_25412);
and U26677 (N_26677,N_25272,N_25101);
and U26678 (N_26678,N_25445,N_25053);
nor U26679 (N_26679,N_25649,N_25202);
or U26680 (N_26680,N_25604,N_25770);
nor U26681 (N_26681,N_25103,N_25626);
and U26682 (N_26682,N_25375,N_25962);
and U26683 (N_26683,N_25248,N_25459);
nor U26684 (N_26684,N_25396,N_25119);
nor U26685 (N_26685,N_25619,N_25324);
xor U26686 (N_26686,N_25832,N_25018);
xnor U26687 (N_26687,N_25083,N_25692);
and U26688 (N_26688,N_25005,N_25144);
nand U26689 (N_26689,N_25541,N_25859);
xor U26690 (N_26690,N_25005,N_25410);
nand U26691 (N_26691,N_25838,N_25361);
or U26692 (N_26692,N_25353,N_25358);
xnor U26693 (N_26693,N_25044,N_25716);
nor U26694 (N_26694,N_25932,N_25459);
and U26695 (N_26695,N_25044,N_25881);
or U26696 (N_26696,N_25158,N_25892);
and U26697 (N_26697,N_25984,N_25214);
nor U26698 (N_26698,N_25395,N_25640);
nor U26699 (N_26699,N_25998,N_25643);
or U26700 (N_26700,N_25942,N_25633);
nand U26701 (N_26701,N_25377,N_25891);
nand U26702 (N_26702,N_25368,N_25531);
nand U26703 (N_26703,N_25916,N_25746);
and U26704 (N_26704,N_25119,N_25123);
xnor U26705 (N_26705,N_25386,N_25771);
and U26706 (N_26706,N_25598,N_25292);
and U26707 (N_26707,N_25617,N_25974);
xor U26708 (N_26708,N_25611,N_25517);
xor U26709 (N_26709,N_25125,N_25253);
and U26710 (N_26710,N_25447,N_25582);
and U26711 (N_26711,N_25553,N_25879);
or U26712 (N_26712,N_25288,N_25147);
nand U26713 (N_26713,N_25089,N_25685);
or U26714 (N_26714,N_25182,N_25350);
nand U26715 (N_26715,N_25574,N_25758);
nand U26716 (N_26716,N_25725,N_25113);
nor U26717 (N_26717,N_25922,N_25911);
nand U26718 (N_26718,N_25067,N_25464);
xnor U26719 (N_26719,N_25987,N_25513);
or U26720 (N_26720,N_25344,N_25350);
xnor U26721 (N_26721,N_25407,N_25700);
xor U26722 (N_26722,N_25476,N_25364);
nor U26723 (N_26723,N_25520,N_25578);
nand U26724 (N_26724,N_25396,N_25012);
or U26725 (N_26725,N_25917,N_25371);
nor U26726 (N_26726,N_25535,N_25032);
and U26727 (N_26727,N_25129,N_25472);
nand U26728 (N_26728,N_25221,N_25749);
xor U26729 (N_26729,N_25529,N_25709);
nor U26730 (N_26730,N_25931,N_25349);
nor U26731 (N_26731,N_25990,N_25773);
xor U26732 (N_26732,N_25498,N_25172);
nor U26733 (N_26733,N_25148,N_25142);
nand U26734 (N_26734,N_25943,N_25673);
xnor U26735 (N_26735,N_25130,N_25921);
nor U26736 (N_26736,N_25210,N_25576);
xnor U26737 (N_26737,N_25048,N_25391);
and U26738 (N_26738,N_25475,N_25585);
or U26739 (N_26739,N_25349,N_25112);
nor U26740 (N_26740,N_25127,N_25545);
nor U26741 (N_26741,N_25143,N_25911);
nor U26742 (N_26742,N_25302,N_25815);
nor U26743 (N_26743,N_25795,N_25384);
nor U26744 (N_26744,N_25395,N_25424);
and U26745 (N_26745,N_25714,N_25991);
nor U26746 (N_26746,N_25254,N_25405);
xor U26747 (N_26747,N_25175,N_25061);
nor U26748 (N_26748,N_25871,N_25304);
nor U26749 (N_26749,N_25044,N_25435);
nor U26750 (N_26750,N_25768,N_25383);
nor U26751 (N_26751,N_25930,N_25484);
xor U26752 (N_26752,N_25782,N_25348);
nor U26753 (N_26753,N_25056,N_25987);
or U26754 (N_26754,N_25636,N_25605);
and U26755 (N_26755,N_25708,N_25985);
or U26756 (N_26756,N_25877,N_25277);
and U26757 (N_26757,N_25434,N_25048);
and U26758 (N_26758,N_25880,N_25824);
xor U26759 (N_26759,N_25746,N_25658);
and U26760 (N_26760,N_25729,N_25430);
or U26761 (N_26761,N_25369,N_25783);
nor U26762 (N_26762,N_25383,N_25920);
nand U26763 (N_26763,N_25123,N_25471);
xnor U26764 (N_26764,N_25687,N_25690);
and U26765 (N_26765,N_25755,N_25986);
or U26766 (N_26766,N_25179,N_25037);
xor U26767 (N_26767,N_25638,N_25257);
xor U26768 (N_26768,N_25512,N_25067);
nor U26769 (N_26769,N_25068,N_25395);
nand U26770 (N_26770,N_25654,N_25404);
and U26771 (N_26771,N_25845,N_25347);
nand U26772 (N_26772,N_25145,N_25069);
and U26773 (N_26773,N_25659,N_25331);
or U26774 (N_26774,N_25078,N_25963);
xnor U26775 (N_26775,N_25470,N_25430);
and U26776 (N_26776,N_25802,N_25890);
nor U26777 (N_26777,N_25050,N_25835);
or U26778 (N_26778,N_25516,N_25489);
nor U26779 (N_26779,N_25088,N_25835);
nor U26780 (N_26780,N_25712,N_25174);
nor U26781 (N_26781,N_25265,N_25412);
nand U26782 (N_26782,N_25259,N_25383);
and U26783 (N_26783,N_25339,N_25916);
nand U26784 (N_26784,N_25841,N_25017);
and U26785 (N_26785,N_25893,N_25463);
nor U26786 (N_26786,N_25828,N_25879);
xor U26787 (N_26787,N_25703,N_25419);
xnor U26788 (N_26788,N_25255,N_25530);
nand U26789 (N_26789,N_25807,N_25013);
xnor U26790 (N_26790,N_25266,N_25928);
or U26791 (N_26791,N_25677,N_25745);
xor U26792 (N_26792,N_25734,N_25218);
xnor U26793 (N_26793,N_25907,N_25638);
and U26794 (N_26794,N_25363,N_25771);
nor U26795 (N_26795,N_25953,N_25406);
nor U26796 (N_26796,N_25580,N_25912);
or U26797 (N_26797,N_25870,N_25383);
xor U26798 (N_26798,N_25254,N_25510);
xor U26799 (N_26799,N_25414,N_25291);
and U26800 (N_26800,N_25726,N_25773);
xor U26801 (N_26801,N_25444,N_25274);
or U26802 (N_26802,N_25698,N_25131);
and U26803 (N_26803,N_25319,N_25482);
nor U26804 (N_26804,N_25274,N_25518);
nor U26805 (N_26805,N_25835,N_25588);
nor U26806 (N_26806,N_25800,N_25909);
and U26807 (N_26807,N_25973,N_25148);
and U26808 (N_26808,N_25019,N_25135);
nor U26809 (N_26809,N_25161,N_25529);
nor U26810 (N_26810,N_25332,N_25886);
nor U26811 (N_26811,N_25687,N_25890);
or U26812 (N_26812,N_25476,N_25721);
and U26813 (N_26813,N_25715,N_25391);
xnor U26814 (N_26814,N_25233,N_25774);
nor U26815 (N_26815,N_25002,N_25055);
nand U26816 (N_26816,N_25171,N_25388);
or U26817 (N_26817,N_25276,N_25458);
xnor U26818 (N_26818,N_25250,N_25365);
or U26819 (N_26819,N_25255,N_25315);
or U26820 (N_26820,N_25439,N_25545);
or U26821 (N_26821,N_25713,N_25065);
nand U26822 (N_26822,N_25362,N_25534);
nor U26823 (N_26823,N_25481,N_25545);
and U26824 (N_26824,N_25851,N_25185);
nor U26825 (N_26825,N_25232,N_25653);
nor U26826 (N_26826,N_25054,N_25322);
or U26827 (N_26827,N_25121,N_25162);
nor U26828 (N_26828,N_25616,N_25876);
or U26829 (N_26829,N_25579,N_25001);
or U26830 (N_26830,N_25053,N_25258);
nand U26831 (N_26831,N_25805,N_25735);
and U26832 (N_26832,N_25599,N_25489);
nor U26833 (N_26833,N_25376,N_25147);
xnor U26834 (N_26834,N_25646,N_25309);
xor U26835 (N_26835,N_25431,N_25215);
nor U26836 (N_26836,N_25200,N_25736);
and U26837 (N_26837,N_25936,N_25427);
xnor U26838 (N_26838,N_25035,N_25825);
and U26839 (N_26839,N_25446,N_25128);
or U26840 (N_26840,N_25435,N_25307);
nor U26841 (N_26841,N_25340,N_25869);
nand U26842 (N_26842,N_25219,N_25251);
and U26843 (N_26843,N_25312,N_25948);
nor U26844 (N_26844,N_25479,N_25676);
and U26845 (N_26845,N_25343,N_25950);
xnor U26846 (N_26846,N_25544,N_25049);
and U26847 (N_26847,N_25568,N_25221);
nor U26848 (N_26848,N_25815,N_25767);
and U26849 (N_26849,N_25218,N_25180);
xnor U26850 (N_26850,N_25224,N_25814);
nand U26851 (N_26851,N_25629,N_25497);
and U26852 (N_26852,N_25434,N_25741);
nor U26853 (N_26853,N_25723,N_25325);
nor U26854 (N_26854,N_25386,N_25148);
nand U26855 (N_26855,N_25241,N_25104);
or U26856 (N_26856,N_25566,N_25336);
xor U26857 (N_26857,N_25549,N_25766);
or U26858 (N_26858,N_25827,N_25342);
and U26859 (N_26859,N_25721,N_25675);
xnor U26860 (N_26860,N_25634,N_25614);
nor U26861 (N_26861,N_25439,N_25909);
or U26862 (N_26862,N_25731,N_25814);
nand U26863 (N_26863,N_25764,N_25878);
and U26864 (N_26864,N_25742,N_25207);
nand U26865 (N_26865,N_25202,N_25031);
or U26866 (N_26866,N_25185,N_25355);
nand U26867 (N_26867,N_25103,N_25165);
nand U26868 (N_26868,N_25036,N_25267);
xor U26869 (N_26869,N_25580,N_25810);
and U26870 (N_26870,N_25193,N_25478);
xnor U26871 (N_26871,N_25551,N_25959);
or U26872 (N_26872,N_25941,N_25074);
nand U26873 (N_26873,N_25574,N_25307);
or U26874 (N_26874,N_25042,N_25611);
nand U26875 (N_26875,N_25210,N_25395);
or U26876 (N_26876,N_25159,N_25955);
and U26877 (N_26877,N_25967,N_25710);
or U26878 (N_26878,N_25864,N_25299);
or U26879 (N_26879,N_25666,N_25762);
and U26880 (N_26880,N_25529,N_25659);
nor U26881 (N_26881,N_25135,N_25807);
nand U26882 (N_26882,N_25441,N_25359);
nand U26883 (N_26883,N_25426,N_25904);
xor U26884 (N_26884,N_25463,N_25692);
nand U26885 (N_26885,N_25563,N_25602);
xnor U26886 (N_26886,N_25721,N_25232);
xor U26887 (N_26887,N_25952,N_25983);
nand U26888 (N_26888,N_25541,N_25429);
or U26889 (N_26889,N_25163,N_25003);
nor U26890 (N_26890,N_25590,N_25905);
nand U26891 (N_26891,N_25041,N_25936);
nor U26892 (N_26892,N_25381,N_25800);
and U26893 (N_26893,N_25388,N_25678);
and U26894 (N_26894,N_25389,N_25469);
nor U26895 (N_26895,N_25828,N_25759);
or U26896 (N_26896,N_25413,N_25126);
xor U26897 (N_26897,N_25870,N_25883);
and U26898 (N_26898,N_25617,N_25559);
xnor U26899 (N_26899,N_25947,N_25146);
and U26900 (N_26900,N_25806,N_25267);
nor U26901 (N_26901,N_25855,N_25146);
nand U26902 (N_26902,N_25338,N_25470);
nand U26903 (N_26903,N_25469,N_25448);
nor U26904 (N_26904,N_25947,N_25290);
and U26905 (N_26905,N_25629,N_25490);
and U26906 (N_26906,N_25655,N_25656);
nand U26907 (N_26907,N_25687,N_25680);
or U26908 (N_26908,N_25217,N_25502);
xnor U26909 (N_26909,N_25180,N_25840);
xnor U26910 (N_26910,N_25253,N_25855);
nor U26911 (N_26911,N_25147,N_25075);
and U26912 (N_26912,N_25699,N_25994);
and U26913 (N_26913,N_25486,N_25845);
or U26914 (N_26914,N_25460,N_25060);
or U26915 (N_26915,N_25033,N_25505);
nor U26916 (N_26916,N_25779,N_25248);
or U26917 (N_26917,N_25803,N_25836);
nor U26918 (N_26918,N_25346,N_25975);
nor U26919 (N_26919,N_25296,N_25347);
and U26920 (N_26920,N_25239,N_25092);
and U26921 (N_26921,N_25474,N_25694);
nor U26922 (N_26922,N_25432,N_25664);
nand U26923 (N_26923,N_25867,N_25320);
or U26924 (N_26924,N_25638,N_25814);
or U26925 (N_26925,N_25634,N_25313);
or U26926 (N_26926,N_25616,N_25849);
nor U26927 (N_26927,N_25092,N_25758);
xor U26928 (N_26928,N_25035,N_25384);
and U26929 (N_26929,N_25980,N_25183);
or U26930 (N_26930,N_25922,N_25934);
nand U26931 (N_26931,N_25097,N_25167);
nor U26932 (N_26932,N_25420,N_25650);
nand U26933 (N_26933,N_25554,N_25952);
and U26934 (N_26934,N_25325,N_25426);
nor U26935 (N_26935,N_25729,N_25632);
or U26936 (N_26936,N_25114,N_25924);
xnor U26937 (N_26937,N_25392,N_25546);
nand U26938 (N_26938,N_25910,N_25032);
or U26939 (N_26939,N_25700,N_25827);
nand U26940 (N_26940,N_25987,N_25472);
nor U26941 (N_26941,N_25429,N_25267);
and U26942 (N_26942,N_25503,N_25999);
nor U26943 (N_26943,N_25337,N_25107);
xor U26944 (N_26944,N_25860,N_25815);
nand U26945 (N_26945,N_25806,N_25240);
and U26946 (N_26946,N_25183,N_25058);
nand U26947 (N_26947,N_25300,N_25380);
and U26948 (N_26948,N_25295,N_25954);
nor U26949 (N_26949,N_25918,N_25689);
or U26950 (N_26950,N_25004,N_25431);
or U26951 (N_26951,N_25358,N_25063);
nand U26952 (N_26952,N_25501,N_25659);
nor U26953 (N_26953,N_25221,N_25771);
nor U26954 (N_26954,N_25631,N_25103);
nand U26955 (N_26955,N_25483,N_25073);
or U26956 (N_26956,N_25758,N_25910);
and U26957 (N_26957,N_25998,N_25096);
xnor U26958 (N_26958,N_25755,N_25341);
or U26959 (N_26959,N_25197,N_25573);
nor U26960 (N_26960,N_25433,N_25622);
nor U26961 (N_26961,N_25668,N_25485);
and U26962 (N_26962,N_25604,N_25448);
xnor U26963 (N_26963,N_25592,N_25351);
xor U26964 (N_26964,N_25211,N_25213);
xnor U26965 (N_26965,N_25105,N_25909);
or U26966 (N_26966,N_25675,N_25729);
xor U26967 (N_26967,N_25159,N_25163);
or U26968 (N_26968,N_25851,N_25957);
xor U26969 (N_26969,N_25046,N_25292);
nor U26970 (N_26970,N_25315,N_25123);
xnor U26971 (N_26971,N_25651,N_25152);
nand U26972 (N_26972,N_25523,N_25180);
nand U26973 (N_26973,N_25450,N_25535);
nor U26974 (N_26974,N_25261,N_25139);
and U26975 (N_26975,N_25097,N_25433);
xor U26976 (N_26976,N_25529,N_25819);
nand U26977 (N_26977,N_25137,N_25623);
xnor U26978 (N_26978,N_25582,N_25347);
nand U26979 (N_26979,N_25138,N_25906);
and U26980 (N_26980,N_25998,N_25670);
xor U26981 (N_26981,N_25155,N_25686);
nor U26982 (N_26982,N_25205,N_25383);
xor U26983 (N_26983,N_25513,N_25371);
nand U26984 (N_26984,N_25733,N_25350);
xor U26985 (N_26985,N_25467,N_25601);
or U26986 (N_26986,N_25098,N_25524);
nand U26987 (N_26987,N_25485,N_25239);
and U26988 (N_26988,N_25070,N_25374);
nor U26989 (N_26989,N_25512,N_25591);
nand U26990 (N_26990,N_25574,N_25590);
or U26991 (N_26991,N_25011,N_25188);
nor U26992 (N_26992,N_25916,N_25020);
nand U26993 (N_26993,N_25241,N_25484);
xor U26994 (N_26994,N_25141,N_25657);
nor U26995 (N_26995,N_25174,N_25400);
nor U26996 (N_26996,N_25375,N_25433);
or U26997 (N_26997,N_25435,N_25514);
xnor U26998 (N_26998,N_25156,N_25165);
nand U26999 (N_26999,N_25774,N_25330);
nand U27000 (N_27000,N_26588,N_26986);
or U27001 (N_27001,N_26328,N_26060);
or U27002 (N_27002,N_26168,N_26812);
nor U27003 (N_27003,N_26739,N_26323);
xor U27004 (N_27004,N_26552,N_26380);
and U27005 (N_27005,N_26308,N_26867);
or U27006 (N_27006,N_26128,N_26260);
nand U27007 (N_27007,N_26881,N_26572);
xor U27008 (N_27008,N_26004,N_26205);
xor U27009 (N_27009,N_26997,N_26605);
nor U27010 (N_27010,N_26575,N_26777);
or U27011 (N_27011,N_26428,N_26754);
and U27012 (N_27012,N_26946,N_26611);
or U27013 (N_27013,N_26884,N_26906);
nor U27014 (N_27014,N_26318,N_26793);
nor U27015 (N_27015,N_26087,N_26163);
nand U27016 (N_27016,N_26885,N_26374);
xor U27017 (N_27017,N_26621,N_26689);
and U27018 (N_27018,N_26847,N_26320);
or U27019 (N_27019,N_26315,N_26731);
nand U27020 (N_27020,N_26039,N_26051);
and U27021 (N_27021,N_26435,N_26031);
and U27022 (N_27022,N_26147,N_26782);
nand U27023 (N_27023,N_26755,N_26512);
xor U27024 (N_27024,N_26618,N_26942);
nand U27025 (N_27025,N_26167,N_26337);
and U27026 (N_27026,N_26693,N_26698);
and U27027 (N_27027,N_26898,N_26985);
xnor U27028 (N_27028,N_26598,N_26427);
xnor U27029 (N_27029,N_26336,N_26834);
or U27030 (N_27030,N_26525,N_26854);
and U27031 (N_27031,N_26983,N_26647);
xor U27032 (N_27032,N_26543,N_26891);
nand U27033 (N_27033,N_26437,N_26599);
xor U27034 (N_27034,N_26827,N_26720);
nand U27035 (N_27035,N_26562,N_26631);
and U27036 (N_27036,N_26027,N_26638);
nand U27037 (N_27037,N_26651,N_26722);
nand U27038 (N_27038,N_26510,N_26893);
nand U27039 (N_27039,N_26800,N_26186);
nand U27040 (N_27040,N_26515,N_26653);
xor U27041 (N_27041,N_26623,N_26862);
or U27042 (N_27042,N_26565,N_26998);
and U27043 (N_27043,N_26046,N_26106);
xnor U27044 (N_27044,N_26369,N_26379);
and U27045 (N_27045,N_26724,N_26803);
nor U27046 (N_27046,N_26982,N_26035);
and U27047 (N_27047,N_26444,N_26700);
or U27048 (N_27048,N_26430,N_26467);
and U27049 (N_27049,N_26970,N_26249);
or U27050 (N_27050,N_26246,N_26578);
or U27051 (N_27051,N_26784,N_26357);
xor U27052 (N_27052,N_26963,N_26936);
nand U27053 (N_27053,N_26386,N_26872);
nor U27054 (N_27054,N_26445,N_26492);
or U27055 (N_27055,N_26240,N_26393);
nand U27056 (N_27056,N_26539,N_26686);
or U27057 (N_27057,N_26877,N_26414);
nand U27058 (N_27058,N_26814,N_26583);
or U27059 (N_27059,N_26619,N_26704);
nor U27060 (N_27060,N_26028,N_26497);
nand U27061 (N_27061,N_26150,N_26110);
or U27062 (N_27062,N_26557,N_26820);
and U27063 (N_27063,N_26289,N_26351);
nor U27064 (N_27064,N_26387,N_26682);
or U27065 (N_27065,N_26865,N_26711);
nor U27066 (N_27066,N_26158,N_26918);
and U27067 (N_27067,N_26262,N_26441);
and U27068 (N_27068,N_26825,N_26394);
nand U27069 (N_27069,N_26071,N_26391);
or U27070 (N_27070,N_26330,N_26355);
nand U27071 (N_27071,N_26836,N_26426);
nand U27072 (N_27072,N_26758,N_26398);
or U27073 (N_27073,N_26453,N_26573);
nand U27074 (N_27074,N_26074,N_26894);
or U27075 (N_27075,N_26607,N_26170);
xor U27076 (N_27076,N_26532,N_26833);
or U27077 (N_27077,N_26053,N_26574);
nor U27078 (N_27078,N_26674,N_26592);
xnor U27079 (N_27079,N_26630,N_26745);
nor U27080 (N_27080,N_26063,N_26223);
and U27081 (N_27081,N_26596,N_26818);
xor U27082 (N_27082,N_26587,N_26786);
xnor U27083 (N_27083,N_26145,N_26256);
nand U27084 (N_27084,N_26645,N_26920);
xnor U27085 (N_27085,N_26734,N_26113);
and U27086 (N_27086,N_26669,N_26171);
nor U27087 (N_27087,N_26247,N_26736);
or U27088 (N_27088,N_26601,N_26826);
xnor U27089 (N_27089,N_26368,N_26684);
and U27090 (N_27090,N_26644,N_26547);
nor U27091 (N_27091,N_26132,N_26399);
xnor U27092 (N_27092,N_26635,N_26560);
xnor U27093 (N_27093,N_26474,N_26189);
and U27094 (N_27094,N_26646,N_26903);
nand U27095 (N_27095,N_26513,N_26664);
and U27096 (N_27096,N_26855,N_26889);
nand U27097 (N_27097,N_26781,N_26420);
nand U27098 (N_27098,N_26727,N_26079);
nor U27099 (N_27099,N_26500,N_26987);
or U27100 (N_27100,N_26962,N_26549);
xor U27101 (N_27101,N_26406,N_26602);
and U27102 (N_27102,N_26233,N_26415);
xor U27103 (N_27103,N_26359,N_26966);
xor U27104 (N_27104,N_26904,N_26251);
xnor U27105 (N_27105,N_26400,N_26707);
and U27106 (N_27106,N_26665,N_26412);
or U27107 (N_27107,N_26397,N_26200);
or U27108 (N_27108,N_26291,N_26934);
nor U27109 (N_27109,N_26327,N_26579);
nand U27110 (N_27110,N_26551,N_26125);
xnor U27111 (N_27111,N_26211,N_26012);
and U27112 (N_27112,N_26114,N_26177);
or U27113 (N_27113,N_26312,N_26124);
and U27114 (N_27114,N_26527,N_26805);
xnor U27115 (N_27115,N_26851,N_26639);
or U27116 (N_27116,N_26356,N_26643);
xnor U27117 (N_27117,N_26570,N_26569);
and U27118 (N_27118,N_26038,N_26191);
xor U27119 (N_27119,N_26155,N_26442);
nor U27120 (N_27120,N_26221,N_26788);
or U27121 (N_27121,N_26058,N_26238);
and U27122 (N_27122,N_26488,N_26384);
xor U27123 (N_27123,N_26296,N_26350);
xnor U27124 (N_27124,N_26600,N_26105);
nand U27125 (N_27125,N_26571,N_26123);
nor U27126 (N_27126,N_26477,N_26436);
xnor U27127 (N_27127,N_26870,N_26556);
nand U27128 (N_27128,N_26801,N_26534);
and U27129 (N_27129,N_26287,N_26075);
or U27130 (N_27130,N_26694,N_26952);
nor U27131 (N_27131,N_26844,N_26264);
or U27132 (N_27132,N_26448,N_26773);
or U27133 (N_27133,N_26005,N_26779);
and U27134 (N_27134,N_26370,N_26797);
xor U27135 (N_27135,N_26710,N_26258);
xnor U27136 (N_27136,N_26136,N_26438);
and U27137 (N_27137,N_26452,N_26971);
or U27138 (N_27138,N_26222,N_26650);
or U27139 (N_27139,N_26135,N_26590);
nor U27140 (N_27140,N_26196,N_26770);
and U27141 (N_27141,N_26678,N_26730);
nor U27142 (N_27142,N_26142,N_26838);
or U27143 (N_27143,N_26849,N_26279);
nand U27144 (N_27144,N_26115,N_26659);
or U27145 (N_27145,N_26916,N_26187);
and U27146 (N_27146,N_26042,N_26895);
xnor U27147 (N_27147,N_26926,N_26133);
nand U27148 (N_27148,N_26540,N_26879);
nand U27149 (N_27149,N_26157,N_26082);
or U27150 (N_27150,N_26768,N_26991);
or U27151 (N_27151,N_26741,N_26511);
or U27152 (N_27152,N_26056,N_26482);
or U27153 (N_27153,N_26306,N_26810);
or U27154 (N_27154,N_26544,N_26129);
xnor U27155 (N_27155,N_26976,N_26914);
nor U27156 (N_27156,N_26748,N_26974);
xor U27157 (N_27157,N_26446,N_26790);
xnor U27158 (N_27158,N_26047,N_26696);
nand U27159 (N_27159,N_26109,N_26830);
nor U27160 (N_27160,N_26888,N_26813);
and U27161 (N_27161,N_26964,N_26747);
xor U27162 (N_27162,N_26016,N_26385);
nor U27163 (N_27163,N_26595,N_26229);
xor U27164 (N_27164,N_26626,N_26176);
xnor U27165 (N_27165,N_26604,N_26506);
nor U27166 (N_27166,N_26712,N_26507);
or U27167 (N_27167,N_26494,N_26283);
or U27168 (N_27168,N_26950,N_26390);
xor U27169 (N_27169,N_26358,N_26036);
and U27170 (N_27170,N_26897,N_26609);
nand U27171 (N_27171,N_26806,N_26403);
or U27172 (N_27172,N_26190,N_26072);
nand U27173 (N_27173,N_26978,N_26218);
or U27174 (N_27174,N_26099,N_26363);
nor U27175 (N_27175,N_26050,N_26945);
and U27176 (N_27176,N_26006,N_26947);
or U27177 (N_27177,N_26178,N_26089);
xor U27178 (N_27178,N_26495,N_26613);
nand U27179 (N_27179,N_26761,N_26941);
nor U27180 (N_27180,N_26160,N_26086);
nor U27181 (N_27181,N_26973,N_26226);
or U27182 (N_27182,N_26902,N_26044);
and U27183 (N_27183,N_26681,N_26993);
xor U27184 (N_27184,N_26301,N_26470);
xnor U27185 (N_27185,N_26269,N_26034);
xor U27186 (N_27186,N_26714,N_26709);
and U27187 (N_27187,N_26487,N_26371);
xor U27188 (N_27188,N_26628,N_26622);
nor U27189 (N_27189,N_26017,N_26325);
or U27190 (N_27190,N_26553,N_26422);
nor U27191 (N_27191,N_26673,N_26546);
and U27192 (N_27192,N_26667,N_26764);
and U27193 (N_27193,N_26091,N_26181);
nor U27194 (N_27194,N_26994,N_26413);
and U27195 (N_27195,N_26666,N_26843);
xnor U27196 (N_27196,N_26835,N_26057);
nor U27197 (N_27197,N_26410,N_26880);
and U27198 (N_27198,N_26995,N_26210);
or U27199 (N_27199,N_26848,N_26498);
and U27200 (N_27200,N_26085,N_26425);
or U27201 (N_27201,N_26496,N_26567);
xnor U27202 (N_27202,N_26118,N_26732);
and U27203 (N_27203,N_26802,N_26933);
nand U27204 (N_27204,N_26915,N_26514);
nor U27205 (N_27205,N_26185,N_26081);
or U27206 (N_27206,N_26454,N_26152);
nor U27207 (N_27207,N_26791,N_26029);
nor U27208 (N_27208,N_26783,N_26120);
and U27209 (N_27209,N_26852,N_26996);
and U27210 (N_27210,N_26938,N_26586);
and U27211 (N_27211,N_26990,N_26676);
nand U27212 (N_27212,N_26340,N_26767);
and U27213 (N_27213,N_26013,N_26148);
nor U27214 (N_27214,N_26365,N_26295);
xor U27215 (N_27215,N_26929,N_26615);
and U27216 (N_27216,N_26939,N_26416);
nor U27217 (N_27217,N_26408,N_26753);
or U27218 (N_27218,N_26321,N_26354);
or U27219 (N_27219,N_26695,N_26577);
and U27220 (N_27220,N_26434,N_26585);
and U27221 (N_27221,N_26280,N_26526);
nor U27222 (N_27222,N_26775,N_26332);
nor U27223 (N_27223,N_26112,N_26288);
or U27224 (N_27224,N_26429,N_26899);
nand U27225 (N_27225,N_26153,N_26648);
and U27226 (N_27226,N_26780,N_26396);
nor U27227 (N_27227,N_26743,N_26491);
nand U27228 (N_27228,N_26887,N_26863);
and U27229 (N_27229,N_26772,N_26204);
xor U27230 (N_27230,N_26959,N_26180);
nor U27231 (N_27231,N_26878,N_26164);
xor U27232 (N_27232,N_26433,N_26203);
or U27233 (N_27233,N_26138,N_26377);
nor U27234 (N_27234,N_26401,N_26041);
or U27235 (N_27235,N_26339,N_26000);
or U27236 (N_27236,N_26307,N_26440);
nand U27237 (N_27237,N_26236,N_26584);
or U27238 (N_27238,N_26531,N_26194);
xor U27239 (N_27239,N_26616,N_26956);
nor U27240 (N_27240,N_26746,N_26612);
nor U27241 (N_27241,N_26424,N_26271);
or U27242 (N_27242,N_26088,N_26451);
nor U27243 (N_27243,N_26930,N_26431);
nor U27244 (N_27244,N_26054,N_26411);
and U27245 (N_27245,N_26311,N_26554);
or U27246 (N_27246,N_26980,N_26119);
and U27247 (N_27247,N_26636,N_26738);
and U27248 (N_27248,N_26943,N_26458);
xor U27249 (N_27249,N_26591,N_26760);
nand U27250 (N_27250,N_26011,N_26671);
or U27251 (N_27251,N_26537,N_26824);
and U27252 (N_27252,N_26095,N_26293);
nand U27253 (N_27253,N_26972,N_26999);
xor U27254 (N_27254,N_26217,N_26703);
xor U27255 (N_27255,N_26008,N_26733);
or U27256 (N_27256,N_26582,N_26921);
and U27257 (N_27257,N_26309,N_26466);
nor U27258 (N_27258,N_26680,N_26750);
nand U27259 (N_27259,N_26846,N_26984);
or U27260 (N_27260,N_26310,N_26209);
and U27261 (N_27261,N_26093,N_26388);
nor U27262 (N_27262,N_26742,N_26502);
or U27263 (N_27263,N_26699,N_26524);
or U27264 (N_27264,N_26961,N_26407);
xor U27265 (N_27265,N_26277,N_26473);
or U27266 (N_27266,N_26227,N_26395);
nand U27267 (N_27267,N_26338,N_26449);
and U27268 (N_27268,N_26907,N_26771);
and U27269 (N_27269,N_26317,N_26183);
nor U27270 (N_27270,N_26104,N_26561);
and U27271 (N_27271,N_26326,N_26098);
nand U27272 (N_27272,N_26232,N_26642);
xnor U27273 (N_27273,N_26333,N_26030);
nand U27274 (N_27274,N_26206,N_26228);
nor U27275 (N_27275,N_26603,N_26284);
xnor U27276 (N_27276,N_26874,N_26859);
or U27277 (N_27277,N_26706,N_26062);
or U27278 (N_27278,N_26342,N_26463);
nor U27279 (N_27279,N_26542,N_26624);
nand U27280 (N_27280,N_26461,N_26392);
or U27281 (N_27281,N_26958,N_26558);
nand U27282 (N_27282,N_26559,N_26480);
and U27283 (N_27283,N_26068,N_26548);
nor U27284 (N_27284,N_26024,N_26977);
nand U27285 (N_27285,N_26179,N_26154);
nand U27286 (N_27286,N_26725,N_26715);
and U27287 (N_27287,N_26021,N_26439);
and U27288 (N_27288,N_26541,N_26485);
nand U27289 (N_27289,N_26381,N_26932);
xnor U27290 (N_27290,N_26637,N_26464);
and U27291 (N_27291,N_26829,N_26744);
nor U27292 (N_27292,N_26762,N_26166);
and U27293 (N_27293,N_26608,N_26346);
or U27294 (N_27294,N_26382,N_26324);
xnor U27295 (N_27295,N_26364,N_26319);
nand U27296 (N_27296,N_26979,N_26216);
xor U27297 (N_27297,N_26242,N_26188);
nor U27298 (N_27298,N_26286,N_26675);
and U27299 (N_27299,N_26316,N_26362);
nand U27300 (N_27300,N_26503,N_26655);
nand U27301 (N_27301,N_26208,N_26841);
nand U27302 (N_27302,N_26064,N_26641);
nand U27303 (N_27303,N_26617,N_26685);
nor U27304 (N_27304,N_26003,N_26234);
and U27305 (N_27305,N_26043,N_26343);
nand U27306 (N_27306,N_26953,N_26007);
and U27307 (N_27307,N_26490,N_26019);
nand U27308 (N_27308,N_26049,N_26352);
xor U27309 (N_27309,N_26302,N_26632);
or U27310 (N_27310,N_26923,N_26789);
nand U27311 (N_27311,N_26219,N_26065);
xnor U27312 (N_27312,N_26530,N_26581);
and U27313 (N_27313,N_26861,N_26735);
and U27314 (N_27314,N_26873,N_26871);
xnor U27315 (N_27315,N_26597,N_26245);
xnor U27316 (N_27316,N_26061,N_26729);
or U27317 (N_27317,N_26025,N_26896);
nor U27318 (N_27318,N_26248,N_26202);
nor U27319 (N_27319,N_26182,N_26130);
nor U27320 (N_27320,N_26564,N_26668);
nor U27321 (N_27321,N_26383,N_26949);
and U27322 (N_27322,N_26823,N_26432);
or U27323 (N_27323,N_26697,N_26716);
nor U27324 (N_27324,N_26169,N_26886);
nor U27325 (N_27325,N_26298,N_26968);
nand U27326 (N_27326,N_26528,N_26184);
xor U27327 (N_27327,N_26140,N_26928);
or U27328 (N_27328,N_26192,N_26869);
or U27329 (N_27329,N_26917,N_26721);
or U27330 (N_27330,N_26389,N_26523);
nand U27331 (N_27331,N_26522,N_26975);
nor U27332 (N_27332,N_26214,N_26468);
nor U27333 (N_27333,N_26931,N_26139);
nand U27334 (N_27334,N_26201,N_26672);
and U27335 (N_27335,N_26225,N_26335);
nor U27336 (N_27336,N_26014,N_26001);
or U27337 (N_27337,N_26417,N_26197);
nor U27338 (N_27338,N_26536,N_26864);
nor U27339 (N_27339,N_26508,N_26483);
or U27340 (N_27340,N_26144,N_26493);
and U27341 (N_27341,N_26077,N_26078);
xnor U27342 (N_27342,N_26811,N_26831);
nor U27343 (N_27343,N_26103,N_26032);
or U27344 (N_27344,N_26804,N_26045);
or U27345 (N_27345,N_26402,N_26465);
xor U27346 (N_27346,N_26111,N_26278);
and U27347 (N_27347,N_26349,N_26076);
or U27348 (N_27348,N_26662,N_26663);
xor U27349 (N_27349,N_26692,N_26719);
and U27350 (N_27350,N_26244,N_26372);
or U27351 (N_27351,N_26765,N_26285);
or U27352 (N_27352,N_26842,N_26272);
and U27353 (N_27353,N_26084,N_26143);
xor U27354 (N_27354,N_26022,N_26489);
xnor U27355 (N_27355,N_26740,N_26718);
xor U27356 (N_27356,N_26471,N_26231);
and U27357 (N_27357,N_26594,N_26299);
or U27358 (N_27358,N_26101,N_26273);
or U27359 (N_27359,N_26876,N_26215);
or U27360 (N_27360,N_26701,N_26083);
xnor U27361 (N_27361,N_26457,N_26499);
or U27362 (N_27362,N_26965,N_26267);
xor U27363 (N_27363,N_26281,N_26620);
xnor U27364 (N_27364,N_26199,N_26728);
xor U27365 (N_27365,N_26717,N_26660);
nand U27366 (N_27366,N_26450,N_26243);
xnor U27367 (N_27367,N_26066,N_26010);
or U27368 (N_27368,N_26988,N_26347);
xnor U27369 (N_27369,N_26459,N_26937);
or U27370 (N_27370,N_26769,N_26796);
xnor U27371 (N_27371,N_26348,N_26213);
and U27372 (N_27372,N_26935,N_26069);
xor U27373 (N_27373,N_26275,N_26992);
nor U27374 (N_27374,N_26606,N_26419);
xor U27375 (N_27375,N_26020,N_26486);
xor U27376 (N_27376,N_26052,N_26509);
nand U27377 (N_27377,N_26787,N_26625);
nand U27378 (N_27378,N_26478,N_26067);
and U27379 (N_27379,N_26883,N_26795);
xor U27380 (N_27380,N_26241,N_26331);
or U27381 (N_27381,N_26860,N_26839);
and U27382 (N_27382,N_26274,N_26856);
xor U27383 (N_27383,N_26094,N_26520);
nor U27384 (N_27384,N_26505,N_26550);
and U27385 (N_27385,N_26265,N_26948);
nor U27386 (N_27386,N_26766,N_26837);
xor U27387 (N_27387,N_26353,N_26195);
xnor U27388 (N_27388,N_26792,N_26033);
or U27389 (N_27389,N_26175,N_26096);
xor U27390 (N_27390,N_26957,N_26361);
xor U27391 (N_27391,N_26304,N_26670);
nor U27392 (N_27392,N_26303,N_26108);
or U27393 (N_27393,N_26633,N_26519);
nor U27394 (N_27394,N_26752,N_26845);
xnor U27395 (N_27395,N_26018,N_26640);
nor U27396 (N_27396,N_26162,N_26819);
xor U27397 (N_27397,N_26922,N_26951);
or U27398 (N_27398,N_26516,N_26455);
nor U27399 (N_27399,N_26266,N_26763);
and U27400 (N_27400,N_26322,N_26418);
or U27401 (N_27401,N_26460,N_26373);
nor U27402 (N_27402,N_26305,N_26905);
and U27403 (N_27403,N_26344,N_26944);
nand U27404 (N_27404,N_26759,N_26866);
xnor U27405 (N_27405,N_26652,N_26174);
xnor U27406 (N_27406,N_26568,N_26954);
or U27407 (N_27407,N_26375,N_26479);
or U27408 (N_27408,N_26149,N_26593);
nor U27409 (N_27409,N_26737,N_26127);
nor U27410 (N_27410,N_26405,N_26092);
or U27411 (N_27411,N_26073,N_26858);
xnor U27412 (N_27412,N_26252,N_26723);
or U27413 (N_27413,N_26751,N_26037);
nor U27414 (N_27414,N_26255,N_26239);
nor U27415 (N_27415,N_26367,N_26015);
xor U27416 (N_27416,N_26237,N_26421);
nand U27417 (N_27417,N_26475,N_26250);
nor U27418 (N_27418,N_26981,N_26313);
and U27419 (N_27419,N_26469,N_26580);
nor U27420 (N_27420,N_26097,N_26687);
and U27421 (N_27421,N_26259,N_26297);
nor U27422 (N_27422,N_26634,N_26100);
nor U27423 (N_27423,N_26808,N_26055);
or U27424 (N_27424,N_26472,N_26009);
or U27425 (N_27425,N_26121,N_26749);
or U27426 (N_27426,N_26913,N_26023);
or U27427 (N_27427,N_26235,N_26161);
xor U27428 (N_27428,N_26253,N_26816);
or U27429 (N_27429,N_26040,N_26576);
and U27430 (N_27430,N_26334,N_26026);
and U27431 (N_27431,N_26654,N_26757);
nor U27432 (N_27432,N_26809,N_26345);
and U27433 (N_27433,N_26156,N_26165);
or U27434 (N_27434,N_26159,N_26261);
nand U27435 (N_27435,N_26137,N_26868);
and U27436 (N_27436,N_26141,N_26927);
nand U27437 (N_27437,N_26679,N_26535);
nor U27438 (N_27438,N_26798,N_26756);
nor U27439 (N_27439,N_26967,N_26409);
nor U27440 (N_27440,N_26443,N_26126);
nand U27441 (N_27441,N_26882,N_26230);
or U27442 (N_27442,N_26048,N_26300);
xnor U27443 (N_27443,N_26924,N_26713);
nor U27444 (N_27444,N_26538,N_26456);
nor U27445 (N_27445,N_26122,N_26447);
and U27446 (N_27446,N_26910,N_26799);
nand U27447 (N_27447,N_26989,N_26940);
nor U27448 (N_27448,N_26151,N_26090);
xnor U27449 (N_27449,N_26521,N_26909);
xnor U27450 (N_27450,N_26070,N_26134);
xnor U27451 (N_27451,N_26360,N_26294);
nand U27452 (N_27452,N_26821,N_26875);
nor U27453 (N_27453,N_26059,N_26815);
nand U27454 (N_27454,N_26224,N_26908);
and U27455 (N_27455,N_26726,N_26504);
and U27456 (N_27456,N_26629,N_26683);
or U27457 (N_27457,N_26254,N_26545);
and U27458 (N_27458,N_26901,N_26193);
nor U27459 (N_27459,N_26131,N_26517);
xor U27460 (N_27460,N_26476,N_26146);
nor U27461 (N_27461,N_26778,N_26850);
nand U27462 (N_27462,N_26840,N_26627);
or U27463 (N_27463,N_26292,N_26366);
and U27464 (N_27464,N_26501,N_26658);
or U27465 (N_27465,N_26807,N_26969);
nand U27466 (N_27466,N_26708,N_26614);
and U27467 (N_27467,N_26900,N_26832);
nand U27468 (N_27468,N_26116,N_26002);
and U27469 (N_27469,N_26198,N_26649);
xor U27470 (N_27470,N_26785,N_26817);
nand U27471 (N_27471,N_26107,N_26314);
or U27472 (N_27472,N_26566,N_26563);
nand U27473 (N_27473,N_26117,N_26207);
xnor U27474 (N_27474,N_26376,N_26688);
xnor U27475 (N_27475,N_26378,N_26341);
and U27476 (N_27476,N_26657,N_26705);
xor U27477 (N_27477,N_26919,N_26890);
and U27478 (N_27478,N_26960,N_26276);
or U27479 (N_27479,N_26462,N_26656);
nor U27480 (N_27480,N_26853,N_26555);
nand U27481 (N_27481,N_26404,N_26270);
nor U27482 (N_27482,N_26911,N_26172);
or U27483 (N_27483,N_26828,N_26484);
xor U27484 (N_27484,N_26955,N_26080);
nand U27485 (N_27485,N_26690,N_26329);
and U27486 (N_27486,N_26912,N_26290);
nor U27487 (N_27487,N_26794,N_26857);
xor U27488 (N_27488,N_26925,N_26892);
nor U27489 (N_27489,N_26529,N_26774);
xor U27490 (N_27490,N_26268,N_26610);
or U27491 (N_27491,N_26220,N_26677);
nand U27492 (N_27492,N_26102,N_26518);
nor U27493 (N_27493,N_26691,N_26776);
nor U27494 (N_27494,N_26661,N_26173);
nand U27495 (N_27495,N_26257,N_26481);
xnor U27496 (N_27496,N_26282,N_26822);
xor U27497 (N_27497,N_26589,N_26212);
nor U27498 (N_27498,N_26702,N_26423);
and U27499 (N_27499,N_26533,N_26263);
and U27500 (N_27500,N_26123,N_26524);
or U27501 (N_27501,N_26785,N_26346);
or U27502 (N_27502,N_26476,N_26355);
nand U27503 (N_27503,N_26901,N_26352);
xor U27504 (N_27504,N_26888,N_26421);
xor U27505 (N_27505,N_26049,N_26090);
nand U27506 (N_27506,N_26690,N_26750);
xor U27507 (N_27507,N_26051,N_26470);
nor U27508 (N_27508,N_26089,N_26388);
or U27509 (N_27509,N_26569,N_26191);
xor U27510 (N_27510,N_26347,N_26329);
nor U27511 (N_27511,N_26470,N_26478);
nand U27512 (N_27512,N_26478,N_26409);
nor U27513 (N_27513,N_26936,N_26223);
nand U27514 (N_27514,N_26318,N_26392);
xor U27515 (N_27515,N_26649,N_26877);
nand U27516 (N_27516,N_26134,N_26616);
xnor U27517 (N_27517,N_26212,N_26499);
nand U27518 (N_27518,N_26085,N_26468);
xor U27519 (N_27519,N_26465,N_26265);
xnor U27520 (N_27520,N_26200,N_26195);
nor U27521 (N_27521,N_26003,N_26960);
xnor U27522 (N_27522,N_26198,N_26457);
nor U27523 (N_27523,N_26936,N_26087);
nor U27524 (N_27524,N_26889,N_26636);
nand U27525 (N_27525,N_26992,N_26086);
nor U27526 (N_27526,N_26543,N_26003);
nand U27527 (N_27527,N_26320,N_26865);
or U27528 (N_27528,N_26403,N_26790);
xnor U27529 (N_27529,N_26539,N_26598);
and U27530 (N_27530,N_26295,N_26873);
or U27531 (N_27531,N_26525,N_26454);
and U27532 (N_27532,N_26529,N_26207);
and U27533 (N_27533,N_26966,N_26397);
nor U27534 (N_27534,N_26211,N_26482);
and U27535 (N_27535,N_26295,N_26558);
or U27536 (N_27536,N_26371,N_26954);
or U27537 (N_27537,N_26698,N_26437);
xnor U27538 (N_27538,N_26109,N_26469);
or U27539 (N_27539,N_26877,N_26540);
nand U27540 (N_27540,N_26176,N_26260);
nand U27541 (N_27541,N_26887,N_26840);
or U27542 (N_27542,N_26615,N_26916);
and U27543 (N_27543,N_26352,N_26585);
nand U27544 (N_27544,N_26110,N_26620);
and U27545 (N_27545,N_26356,N_26621);
nor U27546 (N_27546,N_26736,N_26186);
and U27547 (N_27547,N_26187,N_26035);
or U27548 (N_27548,N_26711,N_26420);
nor U27549 (N_27549,N_26532,N_26303);
nand U27550 (N_27550,N_26916,N_26814);
nor U27551 (N_27551,N_26548,N_26135);
and U27552 (N_27552,N_26989,N_26305);
nand U27553 (N_27553,N_26027,N_26195);
or U27554 (N_27554,N_26523,N_26696);
and U27555 (N_27555,N_26796,N_26120);
or U27556 (N_27556,N_26089,N_26091);
nor U27557 (N_27557,N_26922,N_26334);
or U27558 (N_27558,N_26601,N_26046);
xor U27559 (N_27559,N_26315,N_26810);
nor U27560 (N_27560,N_26696,N_26489);
nand U27561 (N_27561,N_26661,N_26964);
and U27562 (N_27562,N_26479,N_26873);
nor U27563 (N_27563,N_26181,N_26283);
nor U27564 (N_27564,N_26124,N_26867);
and U27565 (N_27565,N_26261,N_26709);
and U27566 (N_27566,N_26337,N_26149);
nand U27567 (N_27567,N_26502,N_26286);
and U27568 (N_27568,N_26826,N_26408);
and U27569 (N_27569,N_26435,N_26583);
xor U27570 (N_27570,N_26161,N_26100);
and U27571 (N_27571,N_26167,N_26971);
or U27572 (N_27572,N_26587,N_26842);
or U27573 (N_27573,N_26426,N_26260);
nand U27574 (N_27574,N_26569,N_26472);
xnor U27575 (N_27575,N_26854,N_26159);
or U27576 (N_27576,N_26688,N_26731);
nand U27577 (N_27577,N_26406,N_26146);
nand U27578 (N_27578,N_26823,N_26211);
or U27579 (N_27579,N_26014,N_26518);
xor U27580 (N_27580,N_26593,N_26694);
nor U27581 (N_27581,N_26809,N_26466);
and U27582 (N_27582,N_26096,N_26890);
nand U27583 (N_27583,N_26885,N_26456);
xnor U27584 (N_27584,N_26390,N_26812);
xnor U27585 (N_27585,N_26605,N_26958);
or U27586 (N_27586,N_26757,N_26085);
nor U27587 (N_27587,N_26467,N_26806);
or U27588 (N_27588,N_26442,N_26686);
nor U27589 (N_27589,N_26583,N_26476);
and U27590 (N_27590,N_26095,N_26798);
nand U27591 (N_27591,N_26208,N_26330);
nand U27592 (N_27592,N_26445,N_26807);
and U27593 (N_27593,N_26561,N_26356);
or U27594 (N_27594,N_26054,N_26612);
and U27595 (N_27595,N_26480,N_26364);
nor U27596 (N_27596,N_26970,N_26303);
or U27597 (N_27597,N_26017,N_26963);
xor U27598 (N_27598,N_26897,N_26922);
nor U27599 (N_27599,N_26874,N_26361);
nor U27600 (N_27600,N_26369,N_26345);
nand U27601 (N_27601,N_26078,N_26781);
or U27602 (N_27602,N_26780,N_26436);
nand U27603 (N_27603,N_26231,N_26496);
xnor U27604 (N_27604,N_26052,N_26161);
or U27605 (N_27605,N_26320,N_26976);
or U27606 (N_27606,N_26335,N_26791);
or U27607 (N_27607,N_26476,N_26147);
xnor U27608 (N_27608,N_26981,N_26336);
xnor U27609 (N_27609,N_26002,N_26609);
nor U27610 (N_27610,N_26555,N_26667);
or U27611 (N_27611,N_26599,N_26367);
nor U27612 (N_27612,N_26713,N_26453);
and U27613 (N_27613,N_26929,N_26720);
and U27614 (N_27614,N_26697,N_26080);
nand U27615 (N_27615,N_26693,N_26960);
and U27616 (N_27616,N_26425,N_26408);
xnor U27617 (N_27617,N_26202,N_26852);
xor U27618 (N_27618,N_26358,N_26471);
or U27619 (N_27619,N_26472,N_26088);
and U27620 (N_27620,N_26018,N_26747);
nor U27621 (N_27621,N_26277,N_26225);
xnor U27622 (N_27622,N_26129,N_26204);
nand U27623 (N_27623,N_26661,N_26241);
or U27624 (N_27624,N_26673,N_26004);
nor U27625 (N_27625,N_26241,N_26364);
and U27626 (N_27626,N_26798,N_26605);
or U27627 (N_27627,N_26011,N_26523);
and U27628 (N_27628,N_26049,N_26568);
or U27629 (N_27629,N_26047,N_26466);
or U27630 (N_27630,N_26133,N_26744);
and U27631 (N_27631,N_26992,N_26388);
xnor U27632 (N_27632,N_26550,N_26733);
nor U27633 (N_27633,N_26469,N_26821);
xor U27634 (N_27634,N_26523,N_26551);
and U27635 (N_27635,N_26913,N_26645);
and U27636 (N_27636,N_26781,N_26719);
and U27637 (N_27637,N_26807,N_26667);
and U27638 (N_27638,N_26166,N_26707);
nor U27639 (N_27639,N_26457,N_26314);
xnor U27640 (N_27640,N_26019,N_26440);
xor U27641 (N_27641,N_26943,N_26211);
and U27642 (N_27642,N_26431,N_26457);
and U27643 (N_27643,N_26029,N_26211);
and U27644 (N_27644,N_26521,N_26687);
nor U27645 (N_27645,N_26294,N_26450);
nor U27646 (N_27646,N_26798,N_26217);
nor U27647 (N_27647,N_26093,N_26197);
nor U27648 (N_27648,N_26038,N_26130);
or U27649 (N_27649,N_26095,N_26397);
nand U27650 (N_27650,N_26181,N_26012);
and U27651 (N_27651,N_26240,N_26138);
xor U27652 (N_27652,N_26683,N_26388);
and U27653 (N_27653,N_26051,N_26199);
or U27654 (N_27654,N_26186,N_26129);
or U27655 (N_27655,N_26005,N_26003);
and U27656 (N_27656,N_26300,N_26841);
xor U27657 (N_27657,N_26773,N_26771);
nor U27658 (N_27658,N_26801,N_26304);
nand U27659 (N_27659,N_26296,N_26093);
or U27660 (N_27660,N_26547,N_26403);
nand U27661 (N_27661,N_26350,N_26561);
or U27662 (N_27662,N_26183,N_26711);
or U27663 (N_27663,N_26967,N_26546);
nand U27664 (N_27664,N_26160,N_26787);
and U27665 (N_27665,N_26888,N_26199);
or U27666 (N_27666,N_26564,N_26990);
nand U27667 (N_27667,N_26442,N_26126);
and U27668 (N_27668,N_26284,N_26713);
and U27669 (N_27669,N_26357,N_26629);
nor U27670 (N_27670,N_26007,N_26677);
nand U27671 (N_27671,N_26405,N_26883);
nand U27672 (N_27672,N_26389,N_26948);
nand U27673 (N_27673,N_26266,N_26163);
or U27674 (N_27674,N_26132,N_26878);
and U27675 (N_27675,N_26702,N_26676);
xnor U27676 (N_27676,N_26102,N_26115);
nand U27677 (N_27677,N_26628,N_26512);
or U27678 (N_27678,N_26993,N_26815);
and U27679 (N_27679,N_26790,N_26541);
or U27680 (N_27680,N_26213,N_26022);
nand U27681 (N_27681,N_26781,N_26121);
nand U27682 (N_27682,N_26881,N_26511);
nor U27683 (N_27683,N_26483,N_26320);
or U27684 (N_27684,N_26612,N_26401);
and U27685 (N_27685,N_26963,N_26860);
nor U27686 (N_27686,N_26348,N_26303);
xor U27687 (N_27687,N_26564,N_26357);
nand U27688 (N_27688,N_26025,N_26746);
and U27689 (N_27689,N_26980,N_26814);
xnor U27690 (N_27690,N_26485,N_26311);
and U27691 (N_27691,N_26444,N_26101);
nor U27692 (N_27692,N_26539,N_26736);
xnor U27693 (N_27693,N_26771,N_26276);
nand U27694 (N_27694,N_26067,N_26289);
and U27695 (N_27695,N_26522,N_26331);
nor U27696 (N_27696,N_26481,N_26277);
nor U27697 (N_27697,N_26470,N_26164);
and U27698 (N_27698,N_26812,N_26871);
nand U27699 (N_27699,N_26413,N_26936);
nor U27700 (N_27700,N_26537,N_26154);
or U27701 (N_27701,N_26233,N_26915);
nand U27702 (N_27702,N_26278,N_26313);
and U27703 (N_27703,N_26950,N_26488);
or U27704 (N_27704,N_26483,N_26982);
xor U27705 (N_27705,N_26368,N_26074);
or U27706 (N_27706,N_26055,N_26659);
nor U27707 (N_27707,N_26739,N_26883);
nand U27708 (N_27708,N_26569,N_26930);
nand U27709 (N_27709,N_26896,N_26354);
or U27710 (N_27710,N_26368,N_26822);
or U27711 (N_27711,N_26523,N_26530);
and U27712 (N_27712,N_26131,N_26757);
nand U27713 (N_27713,N_26623,N_26727);
nand U27714 (N_27714,N_26616,N_26426);
nor U27715 (N_27715,N_26551,N_26949);
and U27716 (N_27716,N_26361,N_26311);
nand U27717 (N_27717,N_26304,N_26696);
xnor U27718 (N_27718,N_26031,N_26356);
nor U27719 (N_27719,N_26627,N_26124);
nand U27720 (N_27720,N_26823,N_26073);
nand U27721 (N_27721,N_26097,N_26343);
nand U27722 (N_27722,N_26236,N_26467);
and U27723 (N_27723,N_26040,N_26575);
xnor U27724 (N_27724,N_26176,N_26668);
nand U27725 (N_27725,N_26432,N_26651);
and U27726 (N_27726,N_26552,N_26064);
or U27727 (N_27727,N_26989,N_26430);
and U27728 (N_27728,N_26836,N_26547);
nor U27729 (N_27729,N_26671,N_26782);
or U27730 (N_27730,N_26150,N_26884);
or U27731 (N_27731,N_26191,N_26070);
and U27732 (N_27732,N_26647,N_26020);
or U27733 (N_27733,N_26660,N_26124);
and U27734 (N_27734,N_26934,N_26447);
xor U27735 (N_27735,N_26139,N_26827);
and U27736 (N_27736,N_26143,N_26080);
or U27737 (N_27737,N_26514,N_26100);
nor U27738 (N_27738,N_26126,N_26549);
and U27739 (N_27739,N_26347,N_26251);
xor U27740 (N_27740,N_26990,N_26542);
or U27741 (N_27741,N_26744,N_26012);
and U27742 (N_27742,N_26496,N_26453);
nor U27743 (N_27743,N_26054,N_26851);
or U27744 (N_27744,N_26664,N_26620);
and U27745 (N_27745,N_26014,N_26150);
or U27746 (N_27746,N_26192,N_26370);
nand U27747 (N_27747,N_26217,N_26981);
nor U27748 (N_27748,N_26662,N_26892);
nor U27749 (N_27749,N_26000,N_26772);
nor U27750 (N_27750,N_26758,N_26448);
xnor U27751 (N_27751,N_26592,N_26506);
nand U27752 (N_27752,N_26086,N_26514);
nor U27753 (N_27753,N_26662,N_26456);
nor U27754 (N_27754,N_26533,N_26537);
xor U27755 (N_27755,N_26227,N_26063);
and U27756 (N_27756,N_26335,N_26046);
or U27757 (N_27757,N_26938,N_26485);
or U27758 (N_27758,N_26791,N_26172);
xor U27759 (N_27759,N_26644,N_26098);
or U27760 (N_27760,N_26994,N_26224);
and U27761 (N_27761,N_26985,N_26476);
or U27762 (N_27762,N_26739,N_26135);
nor U27763 (N_27763,N_26033,N_26634);
and U27764 (N_27764,N_26510,N_26251);
xor U27765 (N_27765,N_26491,N_26885);
xor U27766 (N_27766,N_26790,N_26494);
and U27767 (N_27767,N_26559,N_26267);
and U27768 (N_27768,N_26399,N_26676);
or U27769 (N_27769,N_26435,N_26106);
nand U27770 (N_27770,N_26470,N_26362);
nor U27771 (N_27771,N_26192,N_26490);
and U27772 (N_27772,N_26801,N_26077);
and U27773 (N_27773,N_26724,N_26998);
nand U27774 (N_27774,N_26137,N_26862);
xnor U27775 (N_27775,N_26753,N_26741);
or U27776 (N_27776,N_26797,N_26250);
or U27777 (N_27777,N_26400,N_26391);
and U27778 (N_27778,N_26275,N_26657);
nand U27779 (N_27779,N_26542,N_26749);
or U27780 (N_27780,N_26703,N_26445);
nand U27781 (N_27781,N_26109,N_26826);
xnor U27782 (N_27782,N_26967,N_26676);
nor U27783 (N_27783,N_26444,N_26135);
or U27784 (N_27784,N_26952,N_26386);
nand U27785 (N_27785,N_26791,N_26493);
nand U27786 (N_27786,N_26503,N_26215);
nor U27787 (N_27787,N_26386,N_26867);
xnor U27788 (N_27788,N_26589,N_26929);
nor U27789 (N_27789,N_26505,N_26850);
nand U27790 (N_27790,N_26601,N_26814);
and U27791 (N_27791,N_26750,N_26506);
nor U27792 (N_27792,N_26347,N_26192);
nor U27793 (N_27793,N_26937,N_26381);
nand U27794 (N_27794,N_26050,N_26614);
or U27795 (N_27795,N_26018,N_26398);
nand U27796 (N_27796,N_26544,N_26843);
nand U27797 (N_27797,N_26587,N_26924);
nor U27798 (N_27798,N_26520,N_26135);
xor U27799 (N_27799,N_26528,N_26713);
and U27800 (N_27800,N_26404,N_26637);
nand U27801 (N_27801,N_26321,N_26993);
xnor U27802 (N_27802,N_26805,N_26090);
and U27803 (N_27803,N_26006,N_26801);
or U27804 (N_27804,N_26818,N_26851);
or U27805 (N_27805,N_26424,N_26750);
and U27806 (N_27806,N_26858,N_26448);
nor U27807 (N_27807,N_26839,N_26599);
nor U27808 (N_27808,N_26254,N_26318);
nor U27809 (N_27809,N_26144,N_26968);
nor U27810 (N_27810,N_26077,N_26227);
and U27811 (N_27811,N_26300,N_26832);
xnor U27812 (N_27812,N_26147,N_26391);
and U27813 (N_27813,N_26554,N_26947);
nand U27814 (N_27814,N_26379,N_26423);
nand U27815 (N_27815,N_26341,N_26044);
nand U27816 (N_27816,N_26684,N_26010);
or U27817 (N_27817,N_26206,N_26770);
or U27818 (N_27818,N_26671,N_26065);
nor U27819 (N_27819,N_26748,N_26594);
xor U27820 (N_27820,N_26813,N_26412);
and U27821 (N_27821,N_26964,N_26026);
and U27822 (N_27822,N_26110,N_26422);
nor U27823 (N_27823,N_26613,N_26816);
xnor U27824 (N_27824,N_26656,N_26204);
nand U27825 (N_27825,N_26609,N_26590);
and U27826 (N_27826,N_26991,N_26788);
and U27827 (N_27827,N_26613,N_26580);
and U27828 (N_27828,N_26663,N_26001);
nand U27829 (N_27829,N_26653,N_26346);
or U27830 (N_27830,N_26166,N_26819);
or U27831 (N_27831,N_26665,N_26513);
nor U27832 (N_27832,N_26724,N_26837);
nand U27833 (N_27833,N_26454,N_26642);
xor U27834 (N_27834,N_26358,N_26636);
or U27835 (N_27835,N_26473,N_26245);
or U27836 (N_27836,N_26845,N_26924);
nand U27837 (N_27837,N_26131,N_26075);
xnor U27838 (N_27838,N_26984,N_26775);
xor U27839 (N_27839,N_26156,N_26155);
nand U27840 (N_27840,N_26915,N_26163);
xnor U27841 (N_27841,N_26603,N_26503);
and U27842 (N_27842,N_26577,N_26329);
nor U27843 (N_27843,N_26897,N_26401);
nand U27844 (N_27844,N_26502,N_26859);
xor U27845 (N_27845,N_26319,N_26141);
nor U27846 (N_27846,N_26274,N_26780);
nor U27847 (N_27847,N_26526,N_26542);
and U27848 (N_27848,N_26537,N_26648);
nor U27849 (N_27849,N_26687,N_26045);
nor U27850 (N_27850,N_26774,N_26021);
or U27851 (N_27851,N_26459,N_26651);
or U27852 (N_27852,N_26746,N_26618);
or U27853 (N_27853,N_26068,N_26103);
and U27854 (N_27854,N_26348,N_26885);
and U27855 (N_27855,N_26313,N_26785);
xnor U27856 (N_27856,N_26106,N_26946);
and U27857 (N_27857,N_26684,N_26629);
or U27858 (N_27858,N_26033,N_26650);
nand U27859 (N_27859,N_26989,N_26158);
nand U27860 (N_27860,N_26528,N_26247);
or U27861 (N_27861,N_26603,N_26677);
xor U27862 (N_27862,N_26514,N_26787);
or U27863 (N_27863,N_26508,N_26764);
or U27864 (N_27864,N_26442,N_26056);
and U27865 (N_27865,N_26530,N_26215);
or U27866 (N_27866,N_26695,N_26190);
nand U27867 (N_27867,N_26966,N_26487);
or U27868 (N_27868,N_26245,N_26776);
xnor U27869 (N_27869,N_26077,N_26170);
nor U27870 (N_27870,N_26987,N_26728);
nor U27871 (N_27871,N_26093,N_26348);
or U27872 (N_27872,N_26182,N_26058);
nor U27873 (N_27873,N_26855,N_26207);
and U27874 (N_27874,N_26647,N_26592);
xor U27875 (N_27875,N_26883,N_26401);
and U27876 (N_27876,N_26065,N_26376);
xor U27877 (N_27877,N_26341,N_26911);
nand U27878 (N_27878,N_26003,N_26352);
or U27879 (N_27879,N_26031,N_26436);
xor U27880 (N_27880,N_26473,N_26108);
nor U27881 (N_27881,N_26748,N_26655);
xnor U27882 (N_27882,N_26627,N_26228);
nand U27883 (N_27883,N_26372,N_26357);
or U27884 (N_27884,N_26748,N_26612);
nor U27885 (N_27885,N_26655,N_26431);
and U27886 (N_27886,N_26256,N_26320);
or U27887 (N_27887,N_26171,N_26116);
xor U27888 (N_27888,N_26829,N_26157);
xnor U27889 (N_27889,N_26674,N_26409);
and U27890 (N_27890,N_26745,N_26543);
nand U27891 (N_27891,N_26491,N_26393);
nand U27892 (N_27892,N_26736,N_26404);
xor U27893 (N_27893,N_26494,N_26734);
nand U27894 (N_27894,N_26958,N_26255);
xnor U27895 (N_27895,N_26290,N_26644);
or U27896 (N_27896,N_26494,N_26061);
nand U27897 (N_27897,N_26839,N_26513);
xor U27898 (N_27898,N_26140,N_26613);
nand U27899 (N_27899,N_26720,N_26495);
nand U27900 (N_27900,N_26576,N_26148);
xor U27901 (N_27901,N_26951,N_26516);
nor U27902 (N_27902,N_26310,N_26424);
or U27903 (N_27903,N_26866,N_26757);
nand U27904 (N_27904,N_26577,N_26364);
nand U27905 (N_27905,N_26074,N_26570);
xor U27906 (N_27906,N_26072,N_26519);
and U27907 (N_27907,N_26291,N_26738);
nor U27908 (N_27908,N_26895,N_26166);
nand U27909 (N_27909,N_26719,N_26537);
nand U27910 (N_27910,N_26241,N_26868);
xor U27911 (N_27911,N_26105,N_26873);
or U27912 (N_27912,N_26700,N_26281);
or U27913 (N_27913,N_26037,N_26310);
and U27914 (N_27914,N_26754,N_26852);
and U27915 (N_27915,N_26945,N_26898);
nor U27916 (N_27916,N_26971,N_26341);
nor U27917 (N_27917,N_26715,N_26928);
and U27918 (N_27918,N_26163,N_26292);
and U27919 (N_27919,N_26071,N_26532);
xor U27920 (N_27920,N_26089,N_26460);
xor U27921 (N_27921,N_26954,N_26976);
xnor U27922 (N_27922,N_26666,N_26051);
nor U27923 (N_27923,N_26619,N_26512);
nor U27924 (N_27924,N_26343,N_26631);
and U27925 (N_27925,N_26674,N_26705);
xnor U27926 (N_27926,N_26645,N_26158);
nand U27927 (N_27927,N_26727,N_26333);
and U27928 (N_27928,N_26021,N_26434);
nand U27929 (N_27929,N_26023,N_26651);
nand U27930 (N_27930,N_26556,N_26831);
or U27931 (N_27931,N_26065,N_26117);
nor U27932 (N_27932,N_26575,N_26451);
xnor U27933 (N_27933,N_26177,N_26715);
or U27934 (N_27934,N_26862,N_26262);
xor U27935 (N_27935,N_26899,N_26370);
or U27936 (N_27936,N_26497,N_26308);
or U27937 (N_27937,N_26192,N_26901);
nand U27938 (N_27938,N_26411,N_26507);
nor U27939 (N_27939,N_26806,N_26897);
xor U27940 (N_27940,N_26264,N_26188);
and U27941 (N_27941,N_26024,N_26180);
and U27942 (N_27942,N_26179,N_26577);
xor U27943 (N_27943,N_26801,N_26348);
xor U27944 (N_27944,N_26340,N_26410);
nor U27945 (N_27945,N_26731,N_26503);
or U27946 (N_27946,N_26022,N_26454);
and U27947 (N_27947,N_26648,N_26084);
and U27948 (N_27948,N_26846,N_26607);
or U27949 (N_27949,N_26907,N_26117);
xor U27950 (N_27950,N_26212,N_26469);
nor U27951 (N_27951,N_26383,N_26456);
nand U27952 (N_27952,N_26006,N_26509);
nor U27953 (N_27953,N_26281,N_26123);
and U27954 (N_27954,N_26897,N_26573);
nand U27955 (N_27955,N_26051,N_26830);
nand U27956 (N_27956,N_26450,N_26637);
xor U27957 (N_27957,N_26494,N_26053);
nand U27958 (N_27958,N_26359,N_26760);
nand U27959 (N_27959,N_26632,N_26662);
nand U27960 (N_27960,N_26826,N_26545);
nor U27961 (N_27961,N_26079,N_26928);
and U27962 (N_27962,N_26780,N_26943);
or U27963 (N_27963,N_26764,N_26918);
xor U27964 (N_27964,N_26626,N_26820);
nand U27965 (N_27965,N_26836,N_26160);
nor U27966 (N_27966,N_26186,N_26891);
and U27967 (N_27967,N_26563,N_26026);
nor U27968 (N_27968,N_26158,N_26490);
nor U27969 (N_27969,N_26988,N_26992);
and U27970 (N_27970,N_26616,N_26125);
nor U27971 (N_27971,N_26324,N_26822);
or U27972 (N_27972,N_26282,N_26825);
xnor U27973 (N_27973,N_26465,N_26366);
xnor U27974 (N_27974,N_26227,N_26580);
nand U27975 (N_27975,N_26057,N_26298);
nor U27976 (N_27976,N_26402,N_26509);
xor U27977 (N_27977,N_26554,N_26388);
or U27978 (N_27978,N_26425,N_26988);
xnor U27979 (N_27979,N_26347,N_26229);
xnor U27980 (N_27980,N_26767,N_26711);
and U27981 (N_27981,N_26061,N_26148);
or U27982 (N_27982,N_26915,N_26830);
or U27983 (N_27983,N_26072,N_26209);
or U27984 (N_27984,N_26290,N_26305);
nor U27985 (N_27985,N_26363,N_26178);
xor U27986 (N_27986,N_26931,N_26291);
xnor U27987 (N_27987,N_26716,N_26345);
or U27988 (N_27988,N_26842,N_26694);
or U27989 (N_27989,N_26843,N_26692);
or U27990 (N_27990,N_26197,N_26202);
or U27991 (N_27991,N_26667,N_26907);
nand U27992 (N_27992,N_26046,N_26964);
xor U27993 (N_27993,N_26327,N_26074);
or U27994 (N_27994,N_26204,N_26480);
nand U27995 (N_27995,N_26853,N_26790);
or U27996 (N_27996,N_26183,N_26117);
nand U27997 (N_27997,N_26216,N_26360);
xnor U27998 (N_27998,N_26993,N_26773);
xnor U27999 (N_27999,N_26775,N_26903);
and U28000 (N_28000,N_27319,N_27829);
nor U28001 (N_28001,N_27109,N_27653);
nor U28002 (N_28002,N_27224,N_27197);
nand U28003 (N_28003,N_27294,N_27359);
or U28004 (N_28004,N_27409,N_27688);
nand U28005 (N_28005,N_27933,N_27735);
or U28006 (N_28006,N_27843,N_27292);
nor U28007 (N_28007,N_27942,N_27578);
nand U28008 (N_28008,N_27181,N_27958);
and U28009 (N_28009,N_27943,N_27463);
xor U28010 (N_28010,N_27650,N_27733);
xnor U28011 (N_28011,N_27862,N_27477);
nand U28012 (N_28012,N_27821,N_27452);
nor U28013 (N_28013,N_27972,N_27362);
nor U28014 (N_28014,N_27125,N_27119);
xor U28015 (N_28015,N_27510,N_27937);
xor U28016 (N_28016,N_27651,N_27701);
nor U28017 (N_28017,N_27217,N_27657);
nor U28018 (N_28018,N_27456,N_27929);
nor U28019 (N_28019,N_27711,N_27526);
or U28020 (N_28020,N_27654,N_27345);
nand U28021 (N_28021,N_27503,N_27955);
and U28022 (N_28022,N_27455,N_27435);
and U28023 (N_28023,N_27137,N_27535);
xor U28024 (N_28024,N_27870,N_27133);
nand U28025 (N_28025,N_27306,N_27171);
xnor U28026 (N_28026,N_27176,N_27480);
or U28027 (N_28027,N_27996,N_27403);
nor U28028 (N_28028,N_27911,N_27537);
nand U28029 (N_28029,N_27961,N_27719);
nor U28030 (N_28030,N_27396,N_27582);
or U28031 (N_28031,N_27844,N_27038);
xor U28032 (N_28032,N_27631,N_27177);
nand U28033 (N_28033,N_27635,N_27431);
and U28034 (N_28034,N_27371,N_27614);
nand U28035 (N_28035,N_27694,N_27853);
nand U28036 (N_28036,N_27041,N_27900);
or U28037 (N_28037,N_27325,N_27671);
nor U28038 (N_28038,N_27336,N_27784);
nand U28039 (N_28039,N_27548,N_27953);
nand U28040 (N_28040,N_27069,N_27395);
and U28041 (N_28041,N_27246,N_27000);
and U28042 (N_28042,N_27233,N_27028);
and U28043 (N_28043,N_27804,N_27358);
xnor U28044 (N_28044,N_27831,N_27825);
or U28045 (N_28045,N_27085,N_27814);
or U28046 (N_28046,N_27930,N_27433);
or U28047 (N_28047,N_27718,N_27956);
xor U28048 (N_28048,N_27150,N_27196);
or U28049 (N_28049,N_27785,N_27502);
nand U28050 (N_28050,N_27778,N_27194);
and U28051 (N_28051,N_27732,N_27188);
nor U28052 (N_28052,N_27507,N_27430);
and U28053 (N_28053,N_27628,N_27994);
nand U28054 (N_28054,N_27418,N_27615);
nand U28055 (N_28055,N_27968,N_27494);
nand U28056 (N_28056,N_27415,N_27794);
nand U28057 (N_28057,N_27066,N_27461);
and U28058 (N_28058,N_27216,N_27474);
and U28059 (N_28059,N_27258,N_27849);
or U28060 (N_28060,N_27774,N_27343);
and U28061 (N_28061,N_27779,N_27979);
xor U28062 (N_28062,N_27159,N_27847);
or U28063 (N_28063,N_27812,N_27394);
and U28064 (N_28064,N_27334,N_27245);
and U28065 (N_28065,N_27790,N_27886);
nand U28066 (N_28066,N_27126,N_27006);
and U28067 (N_28067,N_27218,N_27272);
xnor U28068 (N_28068,N_27656,N_27724);
nor U28069 (N_28069,N_27570,N_27748);
or U28070 (N_28070,N_27554,N_27758);
nand U28071 (N_28071,N_27750,N_27161);
and U28072 (N_28072,N_27964,N_27939);
xnor U28073 (N_28073,N_27341,N_27786);
xor U28074 (N_28074,N_27305,N_27860);
or U28075 (N_28075,N_27330,N_27211);
nand U28076 (N_28076,N_27247,N_27948);
xor U28077 (N_28077,N_27068,N_27664);
nand U28078 (N_28078,N_27026,N_27117);
xor U28079 (N_28079,N_27367,N_27749);
or U28080 (N_28080,N_27293,N_27714);
nand U28081 (N_28081,N_27031,N_27589);
and U28082 (N_28082,N_27542,N_27110);
and U28083 (N_28083,N_27282,N_27202);
nand U28084 (N_28084,N_27030,N_27514);
nor U28085 (N_28085,N_27529,N_27501);
nor U28086 (N_28086,N_27241,N_27976);
or U28087 (N_28087,N_27666,N_27407);
or U28088 (N_28088,N_27989,N_27867);
xnor U28089 (N_28089,N_27723,N_27162);
nand U28090 (N_28090,N_27284,N_27412);
nand U28091 (N_28091,N_27070,N_27824);
nor U28092 (N_28092,N_27127,N_27571);
xor U28093 (N_28093,N_27564,N_27486);
or U28094 (N_28094,N_27576,N_27385);
xnor U28095 (N_28095,N_27873,N_27665);
or U28096 (N_28096,N_27339,N_27121);
nand U28097 (N_28097,N_27903,N_27620);
nor U28098 (N_28098,N_27781,N_27184);
and U28099 (N_28099,N_27250,N_27473);
nand U28100 (N_28100,N_27256,N_27260);
or U28101 (N_28101,N_27116,N_27344);
or U28102 (N_28102,N_27215,N_27295);
xnor U28103 (N_28103,N_27533,N_27267);
xnor U28104 (N_28104,N_27562,N_27601);
nor U28105 (N_28105,N_27550,N_27335);
and U28106 (N_28106,N_27500,N_27077);
or U28107 (N_28107,N_27259,N_27050);
nor U28108 (N_28108,N_27329,N_27802);
xor U28109 (N_28109,N_27003,N_27840);
and U28110 (N_28110,N_27591,N_27228);
xnor U28111 (N_28111,N_27826,N_27190);
nor U28112 (N_28112,N_27690,N_27275);
nor U28113 (N_28113,N_27982,N_27475);
xnor U28114 (N_28114,N_27199,N_27042);
or U28115 (N_28115,N_27419,N_27609);
nor U28116 (N_28116,N_27348,N_27149);
or U28117 (N_28117,N_27519,N_27096);
nor U28118 (N_28118,N_27206,N_27745);
or U28119 (N_28119,N_27365,N_27071);
nand U28120 (N_28120,N_27593,N_27299);
and U28121 (N_28121,N_27018,N_27846);
nor U28122 (N_28122,N_27285,N_27816);
xnor U28123 (N_28123,N_27044,N_27327);
nand U28124 (N_28124,N_27630,N_27516);
nand U28125 (N_28125,N_27771,N_27905);
xor U28126 (N_28126,N_27361,N_27378);
and U28127 (N_28127,N_27321,N_27819);
nand U28128 (N_28128,N_27434,N_27495);
nand U28129 (N_28129,N_27225,N_27416);
nor U28130 (N_28130,N_27020,N_27283);
and U28131 (N_28131,N_27424,N_27296);
nand U28132 (N_28132,N_27699,N_27600);
and U28133 (N_28133,N_27737,N_27698);
nor U28134 (N_28134,N_27356,N_27675);
nand U28135 (N_28135,N_27298,N_27744);
xnor U28136 (N_28136,N_27895,N_27466);
xnor U28137 (N_28137,N_27552,N_27405);
nand U28138 (N_28138,N_27059,N_27048);
nand U28139 (N_28139,N_27357,N_27122);
or U28140 (N_28140,N_27565,N_27730);
xnor U28141 (N_28141,N_27072,N_27106);
or U28142 (N_28142,N_27450,N_27114);
nor U28143 (N_28143,N_27896,N_27757);
xor U28144 (N_28144,N_27780,N_27637);
xnor U28145 (N_28145,N_27108,N_27276);
or U28146 (N_28146,N_27483,N_27426);
or U28147 (N_28147,N_27521,N_27340);
and U28148 (N_28148,N_27981,N_27083);
xnor U28149 (N_28149,N_27793,N_27097);
xor U28150 (N_28150,N_27414,N_27890);
nand U28151 (N_28151,N_27249,N_27420);
or U28152 (N_28152,N_27852,N_27488);
xor U28153 (N_28153,N_27153,N_27878);
xor U28154 (N_28154,N_27875,N_27363);
or U28155 (N_28155,N_27054,N_27012);
and U28156 (N_28156,N_27879,N_27248);
or U28157 (N_28157,N_27705,N_27709);
or U28158 (N_28158,N_27314,N_27173);
or U28159 (N_28159,N_27324,N_27621);
nand U28160 (N_28160,N_27629,N_27147);
nand U28161 (N_28161,N_27198,N_27987);
nand U28162 (N_28162,N_27627,N_27478);
nor U28163 (N_28163,N_27471,N_27373);
or U28164 (N_28164,N_27617,N_27892);
or U28165 (N_28165,N_27062,N_27392);
and U28166 (N_28166,N_27261,N_27597);
and U28167 (N_28167,N_27644,N_27207);
nand U28168 (N_28168,N_27763,N_27103);
xnor U28169 (N_28169,N_27947,N_27985);
or U28170 (N_28170,N_27855,N_27192);
xor U28171 (N_28171,N_27935,N_27884);
nor U28172 (N_28172,N_27220,N_27271);
and U28173 (N_28173,N_27320,N_27752);
xnor U28174 (N_28174,N_27406,N_27820);
nor U28175 (N_28175,N_27156,N_27914);
nor U28176 (N_28176,N_27596,N_27386);
nor U28177 (N_28177,N_27756,N_27663);
xnor U28178 (N_28178,N_27379,N_27166);
nor U28179 (N_28179,N_27287,N_27230);
or U28180 (N_28180,N_27047,N_27269);
xor U28181 (N_28181,N_27767,N_27772);
nor U28182 (N_28182,N_27610,N_27572);
nand U28183 (N_28183,N_27584,N_27801);
and U28184 (N_28184,N_27897,N_27616);
nor U28185 (N_28185,N_27755,N_27333);
and U28186 (N_28186,N_27061,N_27859);
nor U28187 (N_28187,N_27795,N_27557);
and U28188 (N_28188,N_27008,N_27787);
nand U28189 (N_28189,N_27612,N_27015);
nor U28190 (N_28190,N_27936,N_27525);
nor U28191 (N_28191,N_27925,N_27010);
nand U28192 (N_28192,N_27204,N_27799);
and U28193 (N_28193,N_27618,N_27439);
nor U28194 (N_28194,N_27446,N_27203);
and U28195 (N_28195,N_27811,N_27684);
nor U28196 (N_28196,N_27851,N_27963);
nand U28197 (N_28197,N_27476,N_27291);
nor U28198 (N_28198,N_27236,N_27809);
nor U28199 (N_28199,N_27586,N_27423);
xor U28200 (N_28200,N_27100,N_27641);
and U28201 (N_28201,N_27729,N_27286);
xor U28202 (N_28202,N_27876,N_27155);
or U28203 (N_28203,N_27965,N_27857);
and U28204 (N_28204,N_27574,N_27832);
nand U28205 (N_28205,N_27101,N_27214);
and U28206 (N_28206,N_27978,N_27798);
or U28207 (N_28207,N_27034,N_27702);
xor U28208 (N_28208,N_27946,N_27370);
nand U28209 (N_28209,N_27229,N_27354);
or U28210 (N_28210,N_27076,N_27393);
nor U28211 (N_28211,N_27513,N_27761);
and U28212 (N_28212,N_27064,N_27080);
or U28213 (N_28213,N_27093,N_27374);
or U28214 (N_28214,N_27776,N_27265);
nor U28215 (N_28215,N_27874,N_27099);
or U28216 (N_28216,N_27950,N_27567);
or U28217 (N_28217,N_27797,N_27753);
or U28218 (N_28218,N_27687,N_27511);
nor U28219 (N_28219,N_27998,N_27604);
and U28220 (N_28220,N_27997,N_27530);
and U28221 (N_28221,N_27545,N_27556);
or U28222 (N_28222,N_27493,N_27850);
nor U28223 (N_28223,N_27845,N_27029);
nand U28224 (N_28224,N_27743,N_27364);
xor U28225 (N_28225,N_27445,N_27993);
or U28226 (N_28226,N_27052,N_27634);
or U28227 (N_28227,N_27973,N_27470);
xor U28228 (N_28228,N_27063,N_27595);
and U28229 (N_28229,N_27736,N_27769);
nand U28230 (N_28230,N_27402,N_27135);
xnor U28231 (N_28231,N_27760,N_27509);
and U28232 (N_28232,N_27536,N_27580);
and U28233 (N_28233,N_27527,N_27540);
or U28234 (N_28234,N_27401,N_27682);
xnor U28235 (N_28235,N_27678,N_27278);
and U28236 (N_28236,N_27893,N_27167);
or U28237 (N_28237,N_27436,N_27971);
nand U28238 (N_28238,N_27390,N_27924);
nor U28239 (N_28239,N_27661,N_27722);
nor U28240 (N_28240,N_27254,N_27607);
and U28241 (N_28241,N_27951,N_27504);
nor U28242 (N_28242,N_27346,N_27738);
nor U28243 (N_28243,N_27623,N_27531);
xnor U28244 (N_28244,N_27277,N_27288);
nand U28245 (N_28245,N_27871,N_27399);
xnor U28246 (N_28246,N_27734,N_27468);
nand U28247 (N_28247,N_27464,N_27090);
nor U28248 (N_28248,N_27704,N_27583);
nor U28249 (N_28249,N_27636,N_27309);
xnor U28250 (N_28250,N_27219,N_27417);
nor U28251 (N_28251,N_27916,N_27124);
nand U28252 (N_28252,N_27238,N_27193);
nand U28253 (N_28253,N_27791,N_27413);
and U28254 (N_28254,N_27592,N_27005);
and U28255 (N_28255,N_27479,N_27086);
nor U28256 (N_28256,N_27342,N_27146);
xor U28257 (N_28257,N_27983,N_27581);
and U28258 (N_28258,N_27541,N_27622);
nor U28259 (N_28259,N_27569,N_27649);
nand U28260 (N_28260,N_27765,N_27624);
or U28261 (N_28261,N_27775,N_27381);
or U28262 (N_28262,N_27459,N_27759);
nand U28263 (N_28263,N_27462,N_27648);
xnor U28264 (N_28264,N_27279,N_27970);
nand U28265 (N_28265,N_27561,N_27932);
xor U28266 (N_28266,N_27172,N_27588);
xor U28267 (N_28267,N_27355,N_27088);
and U28268 (N_28268,N_27404,N_27270);
xor U28269 (N_28269,N_27175,N_27195);
or U28270 (N_28270,N_27280,N_27301);
nor U28271 (N_28271,N_27725,N_27858);
nand U28272 (N_28272,N_27662,N_27465);
and U28273 (N_28273,N_27123,N_27762);
nor U28274 (N_28274,N_27366,N_27881);
and U28275 (N_28275,N_27508,N_27001);
nor U28276 (N_28276,N_27717,N_27836);
xor U28277 (N_28277,N_27449,N_27136);
and U28278 (N_28278,N_27244,N_27553);
and U28279 (N_28279,N_27318,N_27922);
nor U28280 (N_28280,N_27024,N_27689);
xnor U28281 (N_28281,N_27655,N_27647);
or U28282 (N_28282,N_27290,N_27923);
and U28283 (N_28283,N_27907,N_27212);
and U28284 (N_28284,N_27497,N_27766);
xor U28285 (N_28285,N_27865,N_27491);
or U28286 (N_28286,N_27695,N_27023);
and U28287 (N_28287,N_27817,N_27075);
or U28288 (N_28288,N_27864,N_27611);
and U28289 (N_28289,N_27053,N_27777);
or U28290 (N_28290,N_27658,N_27512);
nand U28291 (N_28291,N_27739,N_27073);
nor U28292 (N_28292,N_27598,N_27693);
and U28293 (N_28293,N_27178,N_27489);
or U28294 (N_28294,N_27303,N_27016);
xnor U28295 (N_28295,N_27132,N_27917);
nand U28296 (N_28296,N_27457,N_27443);
or U28297 (N_28297,N_27672,N_27021);
and U28298 (N_28298,N_27255,N_27563);
nor U28299 (N_28299,N_27208,N_27913);
nor U28300 (N_28300,N_27677,N_27049);
nor U28301 (N_28301,N_27506,N_27482);
nand U28302 (N_28302,N_27326,N_27861);
or U28303 (N_28303,N_27170,N_27440);
or U28304 (N_28304,N_27349,N_27013);
or U28305 (N_28305,N_27585,N_27667);
or U28306 (N_28306,N_27713,N_27544);
nor U28307 (N_28307,N_27528,N_27460);
or U28308 (N_28308,N_27988,N_27242);
or U28309 (N_28309,N_27043,N_27888);
or U28310 (N_28310,N_27148,N_27837);
or U28311 (N_28311,N_27539,N_27742);
nor U28312 (N_28312,N_27496,N_27681);
and U28313 (N_28313,N_27154,N_27619);
nor U28314 (N_28314,N_27594,N_27789);
or U28315 (N_28315,N_27331,N_27398);
nor U28316 (N_28316,N_27113,N_27646);
nor U28317 (N_28317,N_27558,N_27613);
nor U28318 (N_28318,N_27057,N_27095);
or U28319 (N_28319,N_27764,N_27067);
nand U28320 (N_28320,N_27222,N_27268);
nand U28321 (N_28321,N_27828,N_27880);
and U28322 (N_28322,N_27518,N_27633);
or U28323 (N_28323,N_27140,N_27454);
or U28324 (N_28324,N_27037,N_27143);
xnor U28325 (N_28325,N_27263,N_27388);
and U28326 (N_28326,N_27902,N_27046);
nor U28327 (N_28327,N_27686,N_27863);
nor U28328 (N_28328,N_27543,N_27472);
and U28329 (N_28329,N_27669,N_27891);
nor U28330 (N_28330,N_27523,N_27727);
xor U28331 (N_28331,N_27920,N_27603);
or U28332 (N_28332,N_27918,N_27901);
xnor U28333 (N_28333,N_27573,N_27183);
and U28334 (N_28334,N_27009,N_27683);
or U28335 (N_28335,N_27894,N_27898);
and U28336 (N_28336,N_27338,N_27209);
or U28337 (N_28337,N_27185,N_27975);
nor U28338 (N_28338,N_27856,N_27118);
and U28339 (N_28339,N_27027,N_27115);
nand U28340 (N_28340,N_27899,N_27350);
nand U28341 (N_28341,N_27397,N_27266);
or U28342 (N_28342,N_27969,N_27237);
nand U28343 (N_28343,N_27376,N_27036);
nand U28344 (N_28344,N_27347,N_27866);
or U28345 (N_28345,N_27954,N_27952);
xnor U28346 (N_28346,N_27626,N_27643);
xor U28347 (N_28347,N_27297,N_27882);
nor U28348 (N_28348,N_27094,N_27264);
nor U28349 (N_28349,N_27164,N_27389);
or U28350 (N_28350,N_27692,N_27382);
xnor U28351 (N_28351,N_27927,N_27427);
nand U28352 (N_28352,N_27962,N_27223);
and U28353 (N_28353,N_27142,N_27231);
or U28354 (N_28354,N_27668,N_27235);
and U28355 (N_28355,N_27712,N_27011);
or U28356 (N_28356,N_27375,N_27065);
nor U28357 (N_28357,N_27377,N_27940);
xor U28358 (N_28358,N_27599,N_27670);
or U28359 (N_28359,N_27708,N_27007);
nand U28360 (N_28360,N_27239,N_27908);
nand U28361 (N_28361,N_27869,N_27251);
nand U28362 (N_28362,N_27841,N_27796);
and U28363 (N_28363,N_27602,N_27240);
or U28364 (N_28364,N_27180,N_27524);
and U28365 (N_28365,N_27673,N_27107);
and U28366 (N_28366,N_27391,N_27906);
nand U28367 (N_28367,N_27490,N_27437);
nand U28368 (N_28368,N_27685,N_27642);
nor U28369 (N_28369,N_27141,N_27575);
or U28370 (N_28370,N_27337,N_27017);
xnor U28371 (N_28371,N_27660,N_27442);
and U28372 (N_28372,N_27104,N_27977);
xor U28373 (N_28373,N_27716,N_27084);
or U28374 (N_28374,N_27138,N_27566);
and U28375 (N_28375,N_27408,N_27715);
or U28376 (N_28376,N_27014,N_27747);
nand U28377 (N_28377,N_27352,N_27441);
or U28378 (N_28378,N_27990,N_27205);
nand U28379 (N_28379,N_27606,N_27081);
xor U28380 (N_28380,N_27720,N_27966);
xnor U28381 (N_28381,N_27960,N_27411);
nor U28382 (N_28382,N_27422,N_27429);
nor U28383 (N_28383,N_27974,N_27191);
or U28384 (N_28384,N_27485,N_27274);
or U28385 (N_28385,N_27721,N_27425);
or U28386 (N_28386,N_27004,N_27885);
and U28387 (N_28387,N_27830,N_27487);
nand U28388 (N_28388,N_27889,N_27517);
nor U28389 (N_28389,N_27060,N_27999);
nand U28390 (N_28390,N_27421,N_27481);
or U28391 (N_28391,N_27316,N_27931);
xor U28392 (N_28392,N_27243,N_27726);
xnor U28393 (N_28393,N_27788,N_27332);
xor U28394 (N_28394,N_27130,N_27751);
xnor U28395 (N_28395,N_27823,N_27696);
nand U28396 (N_28396,N_27174,N_27838);
nor U28397 (N_28397,N_27547,N_27055);
nor U28398 (N_28398,N_27098,N_27967);
nor U28399 (N_28399,N_27213,N_27515);
xnor U28400 (N_28400,N_27144,N_27492);
and U28401 (N_28401,N_27555,N_27451);
or U28402 (N_28402,N_27078,N_27549);
or U28403 (N_28403,N_27674,N_27089);
xor U28404 (N_28404,N_27679,N_27639);
or U28405 (N_28405,N_27587,N_27625);
xor U28406 (N_28406,N_27520,N_27815);
or U28407 (N_28407,N_27728,N_27169);
xnor U28408 (N_28408,N_27221,N_27315);
xor U28409 (N_28409,N_27210,N_27919);
nor U28410 (N_28410,N_27498,N_27458);
nor U28411 (N_28411,N_27313,N_27105);
xor U28412 (N_28412,N_27447,N_27102);
nand U28413 (N_28413,N_27152,N_27058);
or U28414 (N_28414,N_27827,N_27438);
nor U28415 (N_28415,N_27157,N_27910);
nor U28416 (N_28416,N_27934,N_27792);
or U28417 (N_28417,N_27770,N_27035);
nor U28418 (N_28418,N_27710,N_27002);
or U28419 (N_28419,N_27145,N_27201);
xor U28420 (N_28420,N_27731,N_27469);
xnor U28421 (N_28421,N_27383,N_27868);
nand U28422 (N_28422,N_27323,N_27995);
xnor U28423 (N_28423,N_27448,N_27986);
or U28424 (N_28424,N_27833,N_27444);
xnor U28425 (N_28425,N_27308,N_27045);
nand U28426 (N_28426,N_27168,N_27281);
and U28427 (N_28427,N_27453,N_27707);
or U28428 (N_28428,N_27252,N_27112);
nor U28429 (N_28429,N_27959,N_27056);
or U28430 (N_28430,N_27074,N_27659);
or U28431 (N_28431,N_27803,N_27992);
or U28432 (N_28432,N_27703,N_27428);
nor U28433 (N_28433,N_27782,N_27310);
and U28434 (N_28434,N_27040,N_27151);
nor U28435 (N_28435,N_27312,N_27915);
nand U28436 (N_28436,N_27033,N_27351);
xnor U28437 (N_28437,N_27697,N_27091);
or U28438 (N_28438,N_27706,N_27945);
xor U28439 (N_28439,N_27944,N_27652);
xor U28440 (N_28440,N_27307,N_27467);
nor U28441 (N_28441,N_27019,N_27740);
or U28442 (N_28442,N_27590,N_27700);
or U28443 (N_28443,N_27608,N_27991);
xor U28444 (N_28444,N_27773,N_27300);
and U28445 (N_28445,N_27568,N_27111);
and U28446 (N_28446,N_27848,N_27822);
nand U28447 (N_28447,N_27921,N_27546);
or U28448 (N_28448,N_27025,N_27186);
nor U28449 (N_28449,N_27768,N_27928);
or U28450 (N_28450,N_27806,N_27505);
xor U28451 (N_28451,N_27082,N_27234);
nor U28452 (N_28452,N_27805,N_27980);
or U28453 (N_28453,N_27328,N_27092);
nor U28454 (N_28454,N_27165,N_27400);
nand U28455 (N_28455,N_27926,N_27800);
or U28456 (N_28456,N_27560,N_27410);
nor U28457 (N_28457,N_27368,N_27842);
xor U28458 (N_28458,N_27754,N_27179);
or U28459 (N_28459,N_27534,N_27807);
and U28460 (N_28460,N_27160,N_27360);
and U28461 (N_28461,N_27691,N_27387);
nor U28462 (N_28462,N_27128,N_27484);
nor U28463 (N_28463,N_27741,N_27079);
nor U28464 (N_28464,N_27051,N_27808);
and U28465 (N_28465,N_27499,N_27532);
nand U28466 (N_28466,N_27632,N_27227);
and U28467 (N_28467,N_27984,N_27158);
nor U28468 (N_28468,N_27783,N_27605);
nand U28469 (N_28469,N_27134,N_27834);
or U28470 (N_28470,N_27854,N_27189);
and U28471 (N_28471,N_27818,N_27163);
xnor U28472 (N_28472,N_27087,N_27579);
and U28473 (N_28473,N_27559,N_27273);
nand U28474 (N_28474,N_27680,N_27432);
and U28475 (N_28475,N_27129,N_27941);
xnor U28476 (N_28476,N_27289,N_27813);
nor U28477 (N_28477,N_27384,N_27302);
or U28478 (N_28478,N_27949,N_27904);
nor U28479 (N_28479,N_27304,N_27676);
xnor U28480 (N_28480,N_27369,N_27746);
xnor U28481 (N_28481,N_27883,N_27311);
or U28482 (N_28482,N_27638,N_27938);
nor U28483 (N_28483,N_27551,N_27131);
nor U28484 (N_28484,N_27577,N_27810);
nor U28485 (N_28485,N_27182,N_27022);
and U28486 (N_28486,N_27957,N_27322);
and U28487 (N_28487,N_27380,N_27232);
nor U28488 (N_28488,N_27909,N_27262);
and U28489 (N_28489,N_27839,N_27912);
or U28490 (N_28490,N_27835,N_27253);
xnor U28491 (N_28491,N_27887,N_27187);
nor U28492 (N_28492,N_27522,N_27317);
or U28493 (N_28493,N_27645,N_27032);
nand U28494 (N_28494,N_27640,N_27372);
nand U28495 (N_28495,N_27257,N_27120);
xnor U28496 (N_28496,N_27872,N_27200);
nand U28497 (N_28497,N_27877,N_27353);
xor U28498 (N_28498,N_27039,N_27139);
and U28499 (N_28499,N_27226,N_27538);
xnor U28500 (N_28500,N_27623,N_27393);
xnor U28501 (N_28501,N_27559,N_27966);
nand U28502 (N_28502,N_27793,N_27055);
xor U28503 (N_28503,N_27446,N_27589);
and U28504 (N_28504,N_27329,N_27222);
xnor U28505 (N_28505,N_27808,N_27246);
and U28506 (N_28506,N_27265,N_27275);
nand U28507 (N_28507,N_27836,N_27423);
nor U28508 (N_28508,N_27409,N_27491);
xnor U28509 (N_28509,N_27375,N_27043);
nand U28510 (N_28510,N_27972,N_27657);
and U28511 (N_28511,N_27593,N_27540);
or U28512 (N_28512,N_27173,N_27692);
or U28513 (N_28513,N_27585,N_27852);
xnor U28514 (N_28514,N_27352,N_27925);
or U28515 (N_28515,N_27159,N_27800);
or U28516 (N_28516,N_27383,N_27936);
and U28517 (N_28517,N_27861,N_27975);
nor U28518 (N_28518,N_27811,N_27626);
or U28519 (N_28519,N_27642,N_27636);
nand U28520 (N_28520,N_27569,N_27605);
nor U28521 (N_28521,N_27123,N_27989);
nor U28522 (N_28522,N_27006,N_27953);
and U28523 (N_28523,N_27141,N_27849);
and U28524 (N_28524,N_27732,N_27898);
xnor U28525 (N_28525,N_27911,N_27306);
nand U28526 (N_28526,N_27595,N_27940);
and U28527 (N_28527,N_27556,N_27436);
nand U28528 (N_28528,N_27822,N_27877);
nor U28529 (N_28529,N_27552,N_27336);
or U28530 (N_28530,N_27384,N_27139);
nand U28531 (N_28531,N_27692,N_27875);
xnor U28532 (N_28532,N_27563,N_27824);
xnor U28533 (N_28533,N_27745,N_27318);
nor U28534 (N_28534,N_27470,N_27026);
nor U28535 (N_28535,N_27105,N_27722);
nand U28536 (N_28536,N_27118,N_27969);
nand U28537 (N_28537,N_27189,N_27040);
and U28538 (N_28538,N_27478,N_27425);
xor U28539 (N_28539,N_27071,N_27555);
nand U28540 (N_28540,N_27748,N_27104);
or U28541 (N_28541,N_27084,N_27693);
nand U28542 (N_28542,N_27935,N_27699);
nand U28543 (N_28543,N_27033,N_27305);
nor U28544 (N_28544,N_27563,N_27724);
nor U28545 (N_28545,N_27017,N_27728);
nor U28546 (N_28546,N_27071,N_27007);
nor U28547 (N_28547,N_27551,N_27919);
nor U28548 (N_28548,N_27344,N_27933);
nor U28549 (N_28549,N_27452,N_27093);
or U28550 (N_28550,N_27557,N_27238);
or U28551 (N_28551,N_27020,N_27623);
xnor U28552 (N_28552,N_27418,N_27649);
nor U28553 (N_28553,N_27373,N_27806);
and U28554 (N_28554,N_27803,N_27287);
nand U28555 (N_28555,N_27104,N_27056);
xor U28556 (N_28556,N_27664,N_27930);
nor U28557 (N_28557,N_27043,N_27923);
nand U28558 (N_28558,N_27789,N_27298);
and U28559 (N_28559,N_27891,N_27081);
xnor U28560 (N_28560,N_27730,N_27646);
nand U28561 (N_28561,N_27706,N_27307);
nand U28562 (N_28562,N_27739,N_27484);
and U28563 (N_28563,N_27724,N_27296);
xnor U28564 (N_28564,N_27660,N_27835);
nand U28565 (N_28565,N_27946,N_27402);
or U28566 (N_28566,N_27478,N_27510);
and U28567 (N_28567,N_27827,N_27267);
and U28568 (N_28568,N_27778,N_27457);
nand U28569 (N_28569,N_27995,N_27640);
and U28570 (N_28570,N_27543,N_27951);
xor U28571 (N_28571,N_27090,N_27057);
xor U28572 (N_28572,N_27226,N_27448);
nand U28573 (N_28573,N_27590,N_27502);
nand U28574 (N_28574,N_27074,N_27345);
or U28575 (N_28575,N_27244,N_27899);
nand U28576 (N_28576,N_27579,N_27118);
xnor U28577 (N_28577,N_27668,N_27595);
or U28578 (N_28578,N_27752,N_27376);
xor U28579 (N_28579,N_27505,N_27544);
nand U28580 (N_28580,N_27367,N_27825);
and U28581 (N_28581,N_27640,N_27298);
xnor U28582 (N_28582,N_27794,N_27037);
nand U28583 (N_28583,N_27706,N_27762);
nor U28584 (N_28584,N_27217,N_27151);
xnor U28585 (N_28585,N_27057,N_27117);
and U28586 (N_28586,N_27174,N_27858);
or U28587 (N_28587,N_27740,N_27528);
xnor U28588 (N_28588,N_27418,N_27687);
nor U28589 (N_28589,N_27539,N_27573);
or U28590 (N_28590,N_27046,N_27115);
nand U28591 (N_28591,N_27908,N_27621);
and U28592 (N_28592,N_27904,N_27620);
nor U28593 (N_28593,N_27483,N_27410);
xor U28594 (N_28594,N_27319,N_27769);
nand U28595 (N_28595,N_27800,N_27744);
nor U28596 (N_28596,N_27481,N_27546);
and U28597 (N_28597,N_27906,N_27773);
xor U28598 (N_28598,N_27939,N_27170);
or U28599 (N_28599,N_27625,N_27881);
or U28600 (N_28600,N_27742,N_27608);
or U28601 (N_28601,N_27610,N_27344);
nand U28602 (N_28602,N_27614,N_27919);
or U28603 (N_28603,N_27572,N_27224);
and U28604 (N_28604,N_27368,N_27125);
or U28605 (N_28605,N_27876,N_27311);
nor U28606 (N_28606,N_27657,N_27990);
xnor U28607 (N_28607,N_27571,N_27573);
and U28608 (N_28608,N_27336,N_27641);
or U28609 (N_28609,N_27199,N_27235);
nor U28610 (N_28610,N_27644,N_27460);
nor U28611 (N_28611,N_27744,N_27322);
nor U28612 (N_28612,N_27885,N_27981);
or U28613 (N_28613,N_27484,N_27985);
nand U28614 (N_28614,N_27656,N_27219);
nand U28615 (N_28615,N_27863,N_27748);
and U28616 (N_28616,N_27265,N_27842);
nor U28617 (N_28617,N_27175,N_27027);
or U28618 (N_28618,N_27307,N_27989);
nor U28619 (N_28619,N_27789,N_27479);
or U28620 (N_28620,N_27031,N_27617);
nor U28621 (N_28621,N_27330,N_27566);
and U28622 (N_28622,N_27828,N_27561);
xor U28623 (N_28623,N_27010,N_27368);
nor U28624 (N_28624,N_27110,N_27817);
xor U28625 (N_28625,N_27561,N_27093);
xnor U28626 (N_28626,N_27144,N_27591);
and U28627 (N_28627,N_27683,N_27320);
nor U28628 (N_28628,N_27247,N_27827);
and U28629 (N_28629,N_27379,N_27414);
and U28630 (N_28630,N_27237,N_27372);
and U28631 (N_28631,N_27372,N_27456);
or U28632 (N_28632,N_27785,N_27390);
and U28633 (N_28633,N_27213,N_27970);
nand U28634 (N_28634,N_27807,N_27223);
nor U28635 (N_28635,N_27754,N_27103);
nand U28636 (N_28636,N_27214,N_27651);
nand U28637 (N_28637,N_27678,N_27513);
nor U28638 (N_28638,N_27865,N_27423);
nand U28639 (N_28639,N_27873,N_27861);
xor U28640 (N_28640,N_27665,N_27589);
or U28641 (N_28641,N_27989,N_27505);
or U28642 (N_28642,N_27073,N_27225);
xnor U28643 (N_28643,N_27305,N_27826);
xnor U28644 (N_28644,N_27444,N_27231);
xnor U28645 (N_28645,N_27137,N_27648);
and U28646 (N_28646,N_27042,N_27859);
or U28647 (N_28647,N_27867,N_27623);
xnor U28648 (N_28648,N_27671,N_27443);
xnor U28649 (N_28649,N_27837,N_27324);
and U28650 (N_28650,N_27594,N_27407);
nand U28651 (N_28651,N_27955,N_27105);
or U28652 (N_28652,N_27735,N_27711);
nor U28653 (N_28653,N_27216,N_27508);
nand U28654 (N_28654,N_27924,N_27563);
or U28655 (N_28655,N_27221,N_27033);
nand U28656 (N_28656,N_27577,N_27691);
nor U28657 (N_28657,N_27637,N_27227);
and U28658 (N_28658,N_27745,N_27232);
and U28659 (N_28659,N_27777,N_27484);
xnor U28660 (N_28660,N_27537,N_27965);
nor U28661 (N_28661,N_27285,N_27693);
or U28662 (N_28662,N_27973,N_27531);
nor U28663 (N_28663,N_27495,N_27921);
xor U28664 (N_28664,N_27543,N_27006);
xor U28665 (N_28665,N_27821,N_27050);
nor U28666 (N_28666,N_27766,N_27650);
nand U28667 (N_28667,N_27623,N_27563);
and U28668 (N_28668,N_27062,N_27634);
xor U28669 (N_28669,N_27785,N_27426);
or U28670 (N_28670,N_27988,N_27357);
xor U28671 (N_28671,N_27630,N_27910);
nand U28672 (N_28672,N_27741,N_27873);
xor U28673 (N_28673,N_27043,N_27705);
xor U28674 (N_28674,N_27156,N_27638);
xor U28675 (N_28675,N_27013,N_27273);
nor U28676 (N_28676,N_27326,N_27958);
or U28677 (N_28677,N_27260,N_27791);
and U28678 (N_28678,N_27115,N_27441);
xor U28679 (N_28679,N_27202,N_27872);
nand U28680 (N_28680,N_27561,N_27513);
xnor U28681 (N_28681,N_27170,N_27980);
and U28682 (N_28682,N_27883,N_27386);
xor U28683 (N_28683,N_27692,N_27311);
and U28684 (N_28684,N_27693,N_27743);
and U28685 (N_28685,N_27944,N_27167);
or U28686 (N_28686,N_27681,N_27527);
or U28687 (N_28687,N_27456,N_27145);
xor U28688 (N_28688,N_27719,N_27846);
nor U28689 (N_28689,N_27421,N_27539);
or U28690 (N_28690,N_27832,N_27423);
and U28691 (N_28691,N_27772,N_27633);
and U28692 (N_28692,N_27452,N_27949);
nand U28693 (N_28693,N_27715,N_27579);
and U28694 (N_28694,N_27233,N_27150);
and U28695 (N_28695,N_27837,N_27528);
nor U28696 (N_28696,N_27037,N_27803);
xnor U28697 (N_28697,N_27986,N_27200);
nor U28698 (N_28698,N_27534,N_27499);
xor U28699 (N_28699,N_27323,N_27337);
xnor U28700 (N_28700,N_27041,N_27158);
or U28701 (N_28701,N_27155,N_27011);
nor U28702 (N_28702,N_27938,N_27026);
or U28703 (N_28703,N_27588,N_27672);
nor U28704 (N_28704,N_27901,N_27583);
or U28705 (N_28705,N_27949,N_27741);
and U28706 (N_28706,N_27089,N_27555);
nor U28707 (N_28707,N_27176,N_27444);
and U28708 (N_28708,N_27015,N_27132);
nand U28709 (N_28709,N_27717,N_27203);
nand U28710 (N_28710,N_27657,N_27050);
xnor U28711 (N_28711,N_27260,N_27412);
nor U28712 (N_28712,N_27284,N_27989);
nor U28713 (N_28713,N_27455,N_27408);
and U28714 (N_28714,N_27528,N_27948);
nand U28715 (N_28715,N_27221,N_27095);
nor U28716 (N_28716,N_27234,N_27998);
nor U28717 (N_28717,N_27685,N_27855);
and U28718 (N_28718,N_27634,N_27018);
xnor U28719 (N_28719,N_27859,N_27849);
or U28720 (N_28720,N_27311,N_27955);
nor U28721 (N_28721,N_27485,N_27044);
xnor U28722 (N_28722,N_27760,N_27428);
xor U28723 (N_28723,N_27410,N_27629);
or U28724 (N_28724,N_27722,N_27777);
or U28725 (N_28725,N_27148,N_27801);
or U28726 (N_28726,N_27166,N_27593);
xnor U28727 (N_28727,N_27009,N_27968);
and U28728 (N_28728,N_27221,N_27552);
or U28729 (N_28729,N_27267,N_27170);
or U28730 (N_28730,N_27161,N_27539);
and U28731 (N_28731,N_27356,N_27742);
xor U28732 (N_28732,N_27689,N_27286);
and U28733 (N_28733,N_27686,N_27218);
nor U28734 (N_28734,N_27510,N_27848);
and U28735 (N_28735,N_27792,N_27823);
nand U28736 (N_28736,N_27563,N_27610);
xnor U28737 (N_28737,N_27416,N_27022);
or U28738 (N_28738,N_27911,N_27230);
or U28739 (N_28739,N_27663,N_27065);
or U28740 (N_28740,N_27569,N_27796);
nor U28741 (N_28741,N_27325,N_27027);
nor U28742 (N_28742,N_27330,N_27866);
or U28743 (N_28743,N_27656,N_27104);
or U28744 (N_28744,N_27148,N_27540);
nor U28745 (N_28745,N_27931,N_27659);
and U28746 (N_28746,N_27191,N_27639);
nand U28747 (N_28747,N_27037,N_27054);
nand U28748 (N_28748,N_27224,N_27901);
or U28749 (N_28749,N_27768,N_27332);
nand U28750 (N_28750,N_27333,N_27434);
xnor U28751 (N_28751,N_27791,N_27853);
and U28752 (N_28752,N_27679,N_27505);
and U28753 (N_28753,N_27815,N_27951);
xnor U28754 (N_28754,N_27635,N_27172);
nor U28755 (N_28755,N_27085,N_27932);
nand U28756 (N_28756,N_27453,N_27127);
and U28757 (N_28757,N_27125,N_27686);
and U28758 (N_28758,N_27176,N_27630);
and U28759 (N_28759,N_27184,N_27632);
xor U28760 (N_28760,N_27718,N_27842);
or U28761 (N_28761,N_27400,N_27019);
nand U28762 (N_28762,N_27117,N_27077);
and U28763 (N_28763,N_27449,N_27198);
and U28764 (N_28764,N_27796,N_27719);
or U28765 (N_28765,N_27259,N_27252);
xnor U28766 (N_28766,N_27851,N_27365);
xnor U28767 (N_28767,N_27823,N_27586);
or U28768 (N_28768,N_27860,N_27167);
xnor U28769 (N_28769,N_27706,N_27366);
nand U28770 (N_28770,N_27975,N_27503);
nor U28771 (N_28771,N_27154,N_27344);
nor U28772 (N_28772,N_27621,N_27234);
or U28773 (N_28773,N_27234,N_27252);
nor U28774 (N_28774,N_27809,N_27113);
or U28775 (N_28775,N_27350,N_27537);
xnor U28776 (N_28776,N_27803,N_27634);
or U28777 (N_28777,N_27122,N_27841);
or U28778 (N_28778,N_27564,N_27496);
or U28779 (N_28779,N_27220,N_27337);
xor U28780 (N_28780,N_27509,N_27476);
nand U28781 (N_28781,N_27204,N_27167);
or U28782 (N_28782,N_27923,N_27635);
nand U28783 (N_28783,N_27439,N_27589);
nor U28784 (N_28784,N_27112,N_27561);
and U28785 (N_28785,N_27742,N_27569);
and U28786 (N_28786,N_27903,N_27276);
and U28787 (N_28787,N_27013,N_27733);
or U28788 (N_28788,N_27069,N_27526);
xor U28789 (N_28789,N_27791,N_27491);
nor U28790 (N_28790,N_27825,N_27719);
nor U28791 (N_28791,N_27759,N_27726);
xnor U28792 (N_28792,N_27441,N_27801);
xnor U28793 (N_28793,N_27966,N_27702);
and U28794 (N_28794,N_27177,N_27457);
nand U28795 (N_28795,N_27370,N_27842);
xnor U28796 (N_28796,N_27332,N_27381);
xnor U28797 (N_28797,N_27721,N_27697);
nor U28798 (N_28798,N_27685,N_27946);
or U28799 (N_28799,N_27768,N_27626);
or U28800 (N_28800,N_27852,N_27185);
nand U28801 (N_28801,N_27467,N_27321);
nor U28802 (N_28802,N_27955,N_27167);
or U28803 (N_28803,N_27310,N_27150);
xor U28804 (N_28804,N_27600,N_27824);
nor U28805 (N_28805,N_27393,N_27652);
and U28806 (N_28806,N_27360,N_27487);
and U28807 (N_28807,N_27541,N_27980);
or U28808 (N_28808,N_27041,N_27740);
xnor U28809 (N_28809,N_27034,N_27686);
and U28810 (N_28810,N_27061,N_27376);
or U28811 (N_28811,N_27228,N_27674);
xnor U28812 (N_28812,N_27923,N_27554);
and U28813 (N_28813,N_27805,N_27197);
nand U28814 (N_28814,N_27570,N_27992);
nand U28815 (N_28815,N_27891,N_27271);
or U28816 (N_28816,N_27781,N_27483);
and U28817 (N_28817,N_27868,N_27494);
nand U28818 (N_28818,N_27759,N_27582);
nor U28819 (N_28819,N_27516,N_27205);
nand U28820 (N_28820,N_27773,N_27679);
and U28821 (N_28821,N_27442,N_27094);
xnor U28822 (N_28822,N_27850,N_27229);
nor U28823 (N_28823,N_27630,N_27048);
nand U28824 (N_28824,N_27024,N_27590);
or U28825 (N_28825,N_27258,N_27490);
nand U28826 (N_28826,N_27446,N_27430);
nand U28827 (N_28827,N_27788,N_27558);
and U28828 (N_28828,N_27225,N_27598);
nor U28829 (N_28829,N_27025,N_27258);
or U28830 (N_28830,N_27332,N_27695);
xnor U28831 (N_28831,N_27749,N_27259);
nand U28832 (N_28832,N_27693,N_27038);
nand U28833 (N_28833,N_27180,N_27305);
and U28834 (N_28834,N_27260,N_27881);
and U28835 (N_28835,N_27795,N_27599);
nand U28836 (N_28836,N_27788,N_27782);
and U28837 (N_28837,N_27731,N_27459);
nand U28838 (N_28838,N_27855,N_27678);
nand U28839 (N_28839,N_27580,N_27883);
nor U28840 (N_28840,N_27908,N_27965);
xnor U28841 (N_28841,N_27506,N_27996);
and U28842 (N_28842,N_27616,N_27972);
or U28843 (N_28843,N_27176,N_27575);
or U28844 (N_28844,N_27088,N_27495);
nand U28845 (N_28845,N_27532,N_27603);
and U28846 (N_28846,N_27486,N_27357);
or U28847 (N_28847,N_27273,N_27009);
nor U28848 (N_28848,N_27594,N_27309);
and U28849 (N_28849,N_27174,N_27701);
nand U28850 (N_28850,N_27427,N_27734);
or U28851 (N_28851,N_27988,N_27658);
and U28852 (N_28852,N_27644,N_27478);
nor U28853 (N_28853,N_27118,N_27788);
or U28854 (N_28854,N_27085,N_27970);
xor U28855 (N_28855,N_27456,N_27063);
nand U28856 (N_28856,N_27697,N_27273);
and U28857 (N_28857,N_27377,N_27602);
nor U28858 (N_28858,N_27135,N_27047);
or U28859 (N_28859,N_27222,N_27154);
and U28860 (N_28860,N_27116,N_27103);
nor U28861 (N_28861,N_27627,N_27320);
or U28862 (N_28862,N_27975,N_27208);
xnor U28863 (N_28863,N_27034,N_27248);
or U28864 (N_28864,N_27924,N_27062);
nand U28865 (N_28865,N_27659,N_27819);
and U28866 (N_28866,N_27491,N_27280);
nand U28867 (N_28867,N_27345,N_27050);
and U28868 (N_28868,N_27251,N_27573);
xor U28869 (N_28869,N_27965,N_27369);
xor U28870 (N_28870,N_27925,N_27203);
xor U28871 (N_28871,N_27286,N_27032);
and U28872 (N_28872,N_27247,N_27648);
and U28873 (N_28873,N_27579,N_27757);
xnor U28874 (N_28874,N_27659,N_27837);
nand U28875 (N_28875,N_27180,N_27693);
nor U28876 (N_28876,N_27314,N_27955);
or U28877 (N_28877,N_27690,N_27415);
or U28878 (N_28878,N_27624,N_27343);
and U28879 (N_28879,N_27230,N_27261);
or U28880 (N_28880,N_27160,N_27866);
nand U28881 (N_28881,N_27833,N_27554);
xor U28882 (N_28882,N_27762,N_27692);
nand U28883 (N_28883,N_27002,N_27070);
xor U28884 (N_28884,N_27494,N_27852);
or U28885 (N_28885,N_27277,N_27728);
and U28886 (N_28886,N_27858,N_27452);
and U28887 (N_28887,N_27178,N_27086);
xnor U28888 (N_28888,N_27357,N_27844);
xor U28889 (N_28889,N_27039,N_27141);
xnor U28890 (N_28890,N_27524,N_27947);
nor U28891 (N_28891,N_27470,N_27656);
or U28892 (N_28892,N_27437,N_27452);
nor U28893 (N_28893,N_27807,N_27139);
nor U28894 (N_28894,N_27751,N_27994);
or U28895 (N_28895,N_27918,N_27967);
nor U28896 (N_28896,N_27117,N_27133);
and U28897 (N_28897,N_27911,N_27873);
nor U28898 (N_28898,N_27482,N_27598);
and U28899 (N_28899,N_27050,N_27850);
and U28900 (N_28900,N_27012,N_27502);
and U28901 (N_28901,N_27968,N_27987);
nand U28902 (N_28902,N_27787,N_27076);
or U28903 (N_28903,N_27054,N_27579);
or U28904 (N_28904,N_27100,N_27087);
xor U28905 (N_28905,N_27824,N_27411);
nand U28906 (N_28906,N_27747,N_27910);
or U28907 (N_28907,N_27277,N_27434);
nand U28908 (N_28908,N_27092,N_27656);
nor U28909 (N_28909,N_27880,N_27131);
nor U28910 (N_28910,N_27959,N_27627);
nor U28911 (N_28911,N_27289,N_27181);
or U28912 (N_28912,N_27283,N_27212);
xor U28913 (N_28913,N_27245,N_27359);
nor U28914 (N_28914,N_27638,N_27845);
xor U28915 (N_28915,N_27563,N_27140);
nor U28916 (N_28916,N_27260,N_27003);
xnor U28917 (N_28917,N_27947,N_27884);
xor U28918 (N_28918,N_27546,N_27989);
or U28919 (N_28919,N_27302,N_27619);
or U28920 (N_28920,N_27229,N_27199);
and U28921 (N_28921,N_27399,N_27590);
nand U28922 (N_28922,N_27580,N_27863);
and U28923 (N_28923,N_27488,N_27802);
nor U28924 (N_28924,N_27483,N_27592);
or U28925 (N_28925,N_27755,N_27818);
nand U28926 (N_28926,N_27967,N_27104);
xnor U28927 (N_28927,N_27719,N_27357);
and U28928 (N_28928,N_27301,N_27400);
nand U28929 (N_28929,N_27029,N_27986);
and U28930 (N_28930,N_27270,N_27717);
and U28931 (N_28931,N_27577,N_27890);
xor U28932 (N_28932,N_27934,N_27287);
or U28933 (N_28933,N_27798,N_27086);
nor U28934 (N_28934,N_27357,N_27142);
and U28935 (N_28935,N_27879,N_27727);
or U28936 (N_28936,N_27959,N_27262);
xnor U28937 (N_28937,N_27534,N_27142);
and U28938 (N_28938,N_27403,N_27076);
xor U28939 (N_28939,N_27690,N_27978);
nand U28940 (N_28940,N_27629,N_27194);
xnor U28941 (N_28941,N_27818,N_27745);
nor U28942 (N_28942,N_27317,N_27874);
xor U28943 (N_28943,N_27805,N_27361);
and U28944 (N_28944,N_27613,N_27454);
or U28945 (N_28945,N_27186,N_27735);
xor U28946 (N_28946,N_27258,N_27662);
or U28947 (N_28947,N_27632,N_27775);
xnor U28948 (N_28948,N_27624,N_27352);
nand U28949 (N_28949,N_27031,N_27256);
nand U28950 (N_28950,N_27976,N_27843);
nor U28951 (N_28951,N_27395,N_27297);
nand U28952 (N_28952,N_27835,N_27513);
and U28953 (N_28953,N_27444,N_27055);
and U28954 (N_28954,N_27146,N_27587);
and U28955 (N_28955,N_27752,N_27870);
nand U28956 (N_28956,N_27954,N_27823);
nor U28957 (N_28957,N_27085,N_27538);
and U28958 (N_28958,N_27182,N_27737);
and U28959 (N_28959,N_27502,N_27401);
nand U28960 (N_28960,N_27457,N_27085);
nand U28961 (N_28961,N_27256,N_27570);
nand U28962 (N_28962,N_27362,N_27345);
and U28963 (N_28963,N_27217,N_27843);
nor U28964 (N_28964,N_27749,N_27673);
and U28965 (N_28965,N_27041,N_27386);
xnor U28966 (N_28966,N_27982,N_27176);
and U28967 (N_28967,N_27222,N_27915);
or U28968 (N_28968,N_27343,N_27869);
and U28969 (N_28969,N_27593,N_27835);
nand U28970 (N_28970,N_27162,N_27592);
nor U28971 (N_28971,N_27198,N_27187);
and U28972 (N_28972,N_27357,N_27798);
and U28973 (N_28973,N_27963,N_27447);
nand U28974 (N_28974,N_27904,N_27314);
xor U28975 (N_28975,N_27929,N_27485);
nor U28976 (N_28976,N_27611,N_27008);
xor U28977 (N_28977,N_27835,N_27109);
xnor U28978 (N_28978,N_27229,N_27767);
or U28979 (N_28979,N_27541,N_27241);
and U28980 (N_28980,N_27097,N_27906);
and U28981 (N_28981,N_27900,N_27420);
or U28982 (N_28982,N_27280,N_27162);
and U28983 (N_28983,N_27106,N_27289);
or U28984 (N_28984,N_27632,N_27281);
or U28985 (N_28985,N_27754,N_27735);
nor U28986 (N_28986,N_27098,N_27240);
nand U28987 (N_28987,N_27536,N_27370);
nand U28988 (N_28988,N_27137,N_27243);
nor U28989 (N_28989,N_27544,N_27968);
nand U28990 (N_28990,N_27241,N_27610);
xor U28991 (N_28991,N_27300,N_27297);
nor U28992 (N_28992,N_27351,N_27070);
xnor U28993 (N_28993,N_27566,N_27477);
or U28994 (N_28994,N_27387,N_27530);
nand U28995 (N_28995,N_27533,N_27099);
or U28996 (N_28996,N_27412,N_27604);
nand U28997 (N_28997,N_27551,N_27279);
nand U28998 (N_28998,N_27711,N_27878);
and U28999 (N_28999,N_27494,N_27727);
nand U29000 (N_29000,N_28787,N_28417);
and U29001 (N_29001,N_28026,N_28355);
xor U29002 (N_29002,N_28699,N_28428);
xnor U29003 (N_29003,N_28583,N_28304);
xnor U29004 (N_29004,N_28277,N_28205);
or U29005 (N_29005,N_28182,N_28259);
or U29006 (N_29006,N_28169,N_28528);
nor U29007 (N_29007,N_28204,N_28935);
or U29008 (N_29008,N_28704,N_28109);
nor U29009 (N_29009,N_28911,N_28043);
or U29010 (N_29010,N_28585,N_28751);
and U29011 (N_29011,N_28083,N_28061);
and U29012 (N_29012,N_28166,N_28076);
or U29013 (N_29013,N_28489,N_28488);
xnor U29014 (N_29014,N_28587,N_28668);
or U29015 (N_29015,N_28900,N_28721);
xnor U29016 (N_29016,N_28118,N_28392);
nor U29017 (N_29017,N_28505,N_28176);
nand U29018 (N_29018,N_28734,N_28031);
and U29019 (N_29019,N_28020,N_28716);
xnor U29020 (N_29020,N_28363,N_28336);
xnor U29021 (N_29021,N_28389,N_28689);
xnor U29022 (N_29022,N_28448,N_28881);
and U29023 (N_29023,N_28939,N_28074);
nor U29024 (N_29024,N_28374,N_28762);
or U29025 (N_29025,N_28062,N_28605);
or U29026 (N_29026,N_28930,N_28027);
xor U29027 (N_29027,N_28603,N_28616);
xor U29028 (N_29028,N_28570,N_28940);
and U29029 (N_29029,N_28179,N_28743);
and U29030 (N_29030,N_28303,N_28321);
nand U29031 (N_29031,N_28576,N_28287);
or U29032 (N_29032,N_28608,N_28101);
nor U29033 (N_29033,N_28424,N_28157);
and U29034 (N_29034,N_28974,N_28927);
nand U29035 (N_29035,N_28969,N_28993);
nor U29036 (N_29036,N_28727,N_28331);
xor U29037 (N_29037,N_28238,N_28347);
or U29038 (N_29038,N_28046,N_28218);
or U29039 (N_29039,N_28341,N_28460);
nand U29040 (N_29040,N_28311,N_28418);
nand U29041 (N_29041,N_28194,N_28151);
nor U29042 (N_29042,N_28013,N_28917);
or U29043 (N_29043,N_28507,N_28367);
or U29044 (N_29044,N_28469,N_28495);
and U29045 (N_29045,N_28518,N_28636);
xor U29046 (N_29046,N_28849,N_28910);
and U29047 (N_29047,N_28593,N_28122);
nor U29048 (N_29048,N_28954,N_28464);
xor U29049 (N_29049,N_28901,N_28768);
nor U29050 (N_29050,N_28419,N_28113);
and U29051 (N_29051,N_28802,N_28577);
nor U29052 (N_29052,N_28695,N_28415);
and U29053 (N_29053,N_28683,N_28730);
nor U29054 (N_29054,N_28024,N_28407);
or U29055 (N_29055,N_28688,N_28823);
and U29056 (N_29056,N_28792,N_28813);
xnor U29057 (N_29057,N_28081,N_28627);
xnor U29058 (N_29058,N_28245,N_28388);
nand U29059 (N_29059,N_28895,N_28788);
xor U29060 (N_29060,N_28423,N_28868);
or U29061 (N_29061,N_28160,N_28095);
or U29062 (N_29062,N_28738,N_28509);
and U29063 (N_29063,N_28353,N_28493);
nand U29064 (N_29064,N_28834,N_28998);
or U29065 (N_29065,N_28421,N_28427);
xor U29066 (N_29066,N_28105,N_28379);
xor U29067 (N_29067,N_28299,N_28758);
xor U29068 (N_29068,N_28565,N_28847);
or U29069 (N_29069,N_28200,N_28440);
nor U29070 (N_29070,N_28618,N_28432);
nand U29071 (N_29071,N_28386,N_28425);
nor U29072 (N_29072,N_28836,N_28997);
nor U29073 (N_29073,N_28922,N_28138);
or U29074 (N_29074,N_28181,N_28712);
and U29075 (N_29075,N_28978,N_28461);
nor U29076 (N_29076,N_28556,N_28199);
or U29077 (N_29077,N_28560,N_28725);
xor U29078 (N_29078,N_28862,N_28152);
nor U29079 (N_29079,N_28284,N_28017);
or U29080 (N_29080,N_28305,N_28498);
and U29081 (N_29081,N_28288,N_28529);
or U29082 (N_29082,N_28850,N_28808);
xor U29083 (N_29083,N_28091,N_28533);
or U29084 (N_29084,N_28400,N_28470);
and U29085 (N_29085,N_28637,N_28812);
nor U29086 (N_29086,N_28028,N_28579);
nor U29087 (N_29087,N_28621,N_28350);
nand U29088 (N_29088,N_28669,N_28785);
xnor U29089 (N_29089,N_28821,N_28972);
and U29090 (N_29090,N_28269,N_28744);
xor U29091 (N_29091,N_28263,N_28896);
nor U29092 (N_29092,N_28652,N_28686);
xnor U29093 (N_29093,N_28144,N_28296);
nand U29094 (N_29094,N_28855,N_28692);
and U29095 (N_29095,N_28511,N_28237);
nand U29096 (N_29096,N_28970,N_28146);
nor U29097 (N_29097,N_28883,N_28080);
nand U29098 (N_29098,N_28430,N_28597);
xnor U29099 (N_29099,N_28368,N_28713);
or U29100 (N_29100,N_28980,N_28624);
nor U29101 (N_29101,N_28575,N_28063);
nor U29102 (N_29102,N_28025,N_28767);
xnor U29103 (N_29103,N_28796,N_28480);
or U29104 (N_29104,N_28444,N_28957);
nor U29105 (N_29105,N_28958,N_28348);
or U29106 (N_29106,N_28354,N_28441);
or U29107 (N_29107,N_28410,N_28333);
nand U29108 (N_29108,N_28312,N_28822);
or U29109 (N_29109,N_28646,N_28362);
nor U29110 (N_29110,N_28403,N_28859);
nand U29111 (N_29111,N_28573,N_28451);
or U29112 (N_29112,N_28258,N_28516);
and U29113 (N_29113,N_28369,N_28359);
nor U29114 (N_29114,N_28842,N_28938);
nand U29115 (N_29115,N_28019,N_28309);
or U29116 (N_29116,N_28248,N_28745);
and U29117 (N_29117,N_28915,N_28924);
xor U29118 (N_29118,N_28236,N_28942);
and U29119 (N_29119,N_28562,N_28703);
or U29120 (N_29120,N_28462,N_28875);
nor U29121 (N_29121,N_28933,N_28890);
or U29122 (N_29122,N_28051,N_28054);
nand U29123 (N_29123,N_28398,N_28860);
or U29124 (N_29124,N_28319,N_28222);
nand U29125 (N_29125,N_28082,N_28771);
nand U29126 (N_29126,N_28065,N_28376);
or U29127 (N_29127,N_28750,N_28474);
or U29128 (N_29128,N_28271,N_28142);
nor U29129 (N_29129,N_28190,N_28588);
nor U29130 (N_29130,N_28657,N_28919);
nand U29131 (N_29131,N_28292,N_28711);
nor U29132 (N_29132,N_28861,N_28783);
xnor U29133 (N_29133,N_28521,N_28983);
xnor U29134 (N_29134,N_28756,N_28781);
nand U29135 (N_29135,N_28690,N_28965);
xor U29136 (N_29136,N_28174,N_28261);
nor U29137 (N_29137,N_28596,N_28675);
xnor U29138 (N_29138,N_28365,N_28092);
nand U29139 (N_29139,N_28945,N_28156);
or U29140 (N_29140,N_28749,N_28231);
and U29141 (N_29141,N_28210,N_28232);
and U29142 (N_29142,N_28943,N_28035);
xnor U29143 (N_29143,N_28888,N_28235);
nand U29144 (N_29144,N_28439,N_28385);
and U29145 (N_29145,N_28931,N_28530);
or U29146 (N_29146,N_28681,N_28346);
or U29147 (N_29147,N_28519,N_28634);
or U29148 (N_29148,N_28837,N_28022);
xnor U29149 (N_29149,N_28276,N_28793);
xor U29150 (N_29150,N_28542,N_28622);
or U29151 (N_29151,N_28684,N_28056);
and U29152 (N_29152,N_28584,N_28406);
and U29153 (N_29153,N_28093,N_28696);
nor U29154 (N_29154,N_28196,N_28589);
nand U29155 (N_29155,N_28777,N_28548);
xor U29156 (N_29156,N_28453,N_28662);
or U29157 (N_29157,N_28250,N_28459);
xor U29158 (N_29158,N_28798,N_28630);
nor U29159 (N_29159,N_28857,N_28650);
xor U29160 (N_29160,N_28393,N_28302);
nand U29161 (N_29161,N_28178,N_28731);
or U29162 (N_29162,N_28396,N_28714);
xnor U29163 (N_29163,N_28926,N_28908);
xor U29164 (N_29164,N_28639,N_28254);
and U29165 (N_29165,N_28670,N_28158);
nor U29166 (N_29166,N_28854,N_28666);
nor U29167 (N_29167,N_28497,N_28592);
xor U29168 (N_29168,N_28682,N_28549);
nand U29169 (N_29169,N_28955,N_28937);
nand U29170 (N_29170,N_28989,N_28000);
nor U29171 (N_29171,N_28499,N_28060);
and U29172 (N_29172,N_28437,N_28329);
and U29173 (N_29173,N_28332,N_28753);
nand U29174 (N_29174,N_28594,N_28201);
nor U29175 (N_29175,N_28840,N_28984);
nor U29176 (N_29176,N_28343,N_28960);
or U29177 (N_29177,N_28825,N_28534);
or U29178 (N_29178,N_28315,N_28918);
or U29179 (N_29179,N_28571,N_28220);
nand U29180 (N_29180,N_28923,N_28119);
or U29181 (N_29181,N_28366,N_28177);
or U29182 (N_29182,N_28411,N_28852);
or U29183 (N_29183,N_28987,N_28841);
nor U29184 (N_29184,N_28230,N_28981);
or U29185 (N_29185,N_28496,N_28795);
and U29186 (N_29186,N_28759,N_28314);
nand U29187 (N_29187,N_28635,N_28401);
xor U29188 (N_29188,N_28452,N_28904);
and U29189 (N_29189,N_28255,N_28525);
and U29190 (N_29190,N_28766,N_28252);
nor U29191 (N_29191,N_28442,N_28257);
and U29192 (N_29192,N_28877,N_28293);
xnor U29193 (N_29193,N_28936,N_28757);
nor U29194 (N_29194,N_28660,N_28267);
or U29195 (N_29195,N_28242,N_28701);
nor U29196 (N_29196,N_28322,N_28550);
and U29197 (N_29197,N_28752,N_28088);
xor U29198 (N_29198,N_28578,N_28274);
and U29199 (N_29199,N_28905,N_28044);
or U29200 (N_29200,N_28773,N_28941);
nor U29201 (N_29201,N_28186,N_28833);
and U29202 (N_29202,N_28869,N_28463);
and U29203 (N_29203,N_28581,N_28643);
or U29204 (N_29204,N_28818,N_28626);
nand U29205 (N_29205,N_28640,N_28582);
or U29206 (N_29206,N_28990,N_28104);
nand U29207 (N_29207,N_28717,N_28914);
and U29208 (N_29208,N_28420,N_28010);
or U29209 (N_29209,N_28283,N_28988);
or U29210 (N_29210,N_28098,N_28475);
and U29211 (N_29211,N_28566,N_28619);
nand U29212 (N_29212,N_28364,N_28246);
nand U29213 (N_29213,N_28677,N_28953);
nand U29214 (N_29214,N_28503,N_28121);
xnor U29215 (N_29215,N_28599,N_28223);
xor U29216 (N_29216,N_28002,N_28510);
or U29217 (N_29217,N_28794,N_28951);
or U29218 (N_29218,N_28541,N_28378);
nor U29219 (N_29219,N_28185,N_28115);
xor U29220 (N_29220,N_28819,N_28815);
nor U29221 (N_29221,N_28048,N_28478);
xnor U29222 (N_29222,N_28382,N_28371);
and U29223 (N_29223,N_28195,N_28645);
xnor U29224 (N_29224,N_28431,N_28213);
and U29225 (N_29225,N_28967,N_28372);
xnor U29226 (N_29226,N_28553,N_28995);
nor U29227 (N_29227,N_28617,N_28625);
and U29228 (N_29228,N_28710,N_28206);
or U29229 (N_29229,N_28191,N_28748);
or U29230 (N_29230,N_28467,N_28127);
nand U29231 (N_29231,N_28700,N_28663);
nor U29232 (N_29232,N_28806,N_28728);
nor U29233 (N_29233,N_28632,N_28673);
nand U29234 (N_29234,N_28897,N_28828);
nor U29235 (N_29235,N_28159,N_28527);
or U29236 (N_29236,N_28898,N_28886);
nor U29237 (N_29237,N_28800,N_28057);
nor U29238 (N_29238,N_28887,N_28239);
nor U29239 (N_29239,N_28014,N_28784);
or U29240 (N_29240,N_28391,N_28172);
nor U29241 (N_29241,N_28522,N_28128);
xor U29242 (N_29242,N_28340,N_28535);
nor U29243 (N_29243,N_28208,N_28047);
and U29244 (N_29244,N_28789,N_28233);
xor U29245 (N_29245,N_28099,N_28906);
or U29246 (N_29246,N_28135,N_28672);
nor U29247 (N_29247,N_28066,N_28724);
xor U29248 (N_29248,N_28033,N_28572);
or U29249 (N_29249,N_28243,N_28435);
nor U29250 (N_29250,N_28880,N_28568);
or U29251 (N_29251,N_28810,N_28107);
or U29252 (N_29252,N_28380,N_28387);
or U29253 (N_29253,N_28740,N_28709);
nor U29254 (N_29254,N_28183,N_28648);
and U29255 (N_29255,N_28003,N_28273);
or U29256 (N_29256,N_28811,N_28718);
or U29257 (N_29257,N_28532,N_28885);
or U29258 (N_29258,N_28702,N_28545);
nor U29259 (N_29259,N_28733,N_28449);
or U29260 (N_29260,N_28558,N_28851);
and U29261 (N_29261,N_28438,N_28665);
nor U29262 (N_29262,N_28286,N_28045);
and U29263 (N_29263,N_28275,N_28502);
or U29264 (N_29264,N_28486,N_28244);
nor U29265 (N_29265,N_28656,N_28538);
nor U29266 (N_29266,N_28306,N_28112);
or U29267 (N_29267,N_28563,N_28039);
nor U29268 (N_29268,N_28858,N_28832);
nand U29269 (N_29269,N_28465,N_28772);
nor U29270 (N_29270,N_28994,N_28075);
nand U29271 (N_29271,N_28433,N_28468);
or U29272 (N_29272,N_28591,N_28472);
or U29273 (N_29273,N_28466,N_28780);
and U29274 (N_29274,N_28059,N_28876);
xor U29275 (N_29275,N_28884,N_28557);
or U29276 (N_29276,N_28012,N_28167);
xor U29277 (N_29277,N_28586,N_28999);
and U29278 (N_29278,N_28456,N_28547);
or U29279 (N_29279,N_28069,N_28327);
nor U29280 (N_29280,N_28394,N_28755);
nor U29281 (N_29281,N_28086,N_28085);
xnor U29282 (N_29282,N_28590,N_28778);
nor U29283 (N_29283,N_28087,N_28030);
xor U29284 (N_29284,N_28878,N_28279);
xnor U29285 (N_29285,N_28604,N_28889);
nor U29286 (N_29286,N_28126,N_28925);
and U29287 (N_29287,N_28517,N_28377);
xnor U29288 (N_29288,N_28829,N_28893);
or U29289 (N_29289,N_28153,N_28328);
and U29290 (N_29290,N_28154,N_28356);
xnor U29291 (N_29291,N_28602,N_28264);
or U29292 (N_29292,N_28843,N_28073);
or U29293 (N_29293,N_28187,N_28402);
nor U29294 (N_29294,N_28982,N_28149);
xnor U29295 (N_29295,N_28803,N_28620);
nand U29296 (N_29296,N_28839,N_28612);
nand U29297 (N_29297,N_28053,N_28976);
or U29298 (N_29298,N_28217,N_28316);
and U29299 (N_29299,N_28872,N_28150);
or U29300 (N_29300,N_28455,N_28330);
nand U29301 (N_29301,N_28959,N_28077);
xor U29302 (N_29302,N_28058,N_28977);
or U29303 (N_29303,N_28021,N_28506);
or U29304 (N_29304,N_28776,N_28963);
xor U29305 (N_29305,N_28985,N_28546);
nor U29306 (N_29306,N_28551,N_28055);
xnor U29307 (N_29307,N_28644,N_28317);
nand U29308 (N_29308,N_28633,N_28947);
nand U29309 (N_29309,N_28826,N_28848);
xor U29310 (N_29310,N_28479,N_28909);
nor U29311 (N_29311,N_28193,N_28814);
nand U29312 (N_29312,N_28623,N_28552);
or U29313 (N_29313,N_28323,N_28416);
or U29314 (N_29314,N_28189,N_28342);
nor U29315 (N_29315,N_28240,N_28735);
nor U29316 (N_29316,N_28383,N_28214);
nand U29317 (N_29317,N_28746,N_28034);
nand U29318 (N_29318,N_28671,N_28471);
nor U29319 (N_29319,N_28397,N_28009);
xor U29320 (N_29320,N_28764,N_28447);
and U29321 (N_29321,N_28129,N_28674);
nor U29322 (N_29322,N_28490,N_28761);
and U29323 (N_29323,N_28268,N_28697);
or U29324 (N_29324,N_28485,N_28050);
or U29325 (N_29325,N_28865,N_28395);
nor U29326 (N_29326,N_28229,N_28638);
xor U29327 (N_29327,N_28100,N_28520);
nand U29328 (N_29328,N_28197,N_28732);
nor U29329 (N_29329,N_28477,N_28687);
and U29330 (N_29330,N_28540,N_28171);
or U29331 (N_29331,N_28907,N_28120);
nand U29332 (N_29332,N_28831,N_28147);
and U29333 (N_29333,N_28032,N_28873);
or U29334 (N_29334,N_28698,N_28291);
or U29335 (N_29335,N_28531,N_28096);
nand U29336 (N_29336,N_28537,N_28763);
and U29337 (N_29337,N_28145,N_28301);
xor U29338 (N_29338,N_28116,N_28443);
and U29339 (N_29339,N_28289,N_28155);
xor U29340 (N_29340,N_28337,N_28726);
nand U29341 (N_29341,N_28864,N_28559);
nand U29342 (N_29342,N_28790,N_28856);
or U29343 (N_29343,N_28184,N_28114);
or U29344 (N_29344,N_28102,N_28655);
nand U29345 (N_29345,N_28791,N_28760);
nand U29346 (N_29346,N_28262,N_28729);
and U29347 (N_29347,N_28979,N_28870);
and U29348 (N_29348,N_28770,N_28253);
and U29349 (N_29349,N_28132,N_28008);
xnor U29350 (N_29350,N_28631,N_28708);
nor U29351 (N_29351,N_28816,N_28804);
nor U29352 (N_29352,N_28137,N_28281);
nand U29353 (N_29353,N_28294,N_28405);
xnor U29354 (N_29354,N_28140,N_28600);
nor U29355 (N_29355,N_28966,N_28226);
and U29356 (N_29356,N_28500,N_28139);
nand U29357 (N_29357,N_28295,N_28601);
nor U29358 (N_29358,N_28015,N_28260);
nor U29359 (N_29359,N_28280,N_28741);
nand U29360 (N_29360,N_28029,N_28962);
xor U29361 (N_29361,N_28647,N_28384);
xnor U29362 (N_29362,N_28318,N_28125);
nand U29363 (N_29363,N_28426,N_28487);
nor U29364 (N_29364,N_28004,N_28799);
nand U29365 (N_29365,N_28338,N_28929);
xor U29366 (N_29366,N_28554,N_28824);
or U29367 (N_29367,N_28006,N_28765);
or U29368 (N_29368,N_28345,N_28946);
nor U29369 (N_29369,N_28412,N_28298);
nand U29370 (N_29370,N_28606,N_28266);
and U29371 (N_29371,N_28921,N_28747);
or U29372 (N_29372,N_28801,N_28409);
nand U29373 (N_29373,N_28251,N_28564);
nor U29374 (N_29374,N_28971,N_28052);
nand U29375 (N_29375,N_28361,N_28163);
or U29376 (N_29376,N_28706,N_28968);
or U29377 (N_29377,N_28515,N_28899);
nor U29378 (N_29378,N_28344,N_28580);
xor U29379 (N_29379,N_28956,N_28221);
nor U29380 (N_29380,N_28664,N_28739);
nand U29381 (N_29381,N_28106,N_28016);
and U29382 (N_29382,N_28705,N_28595);
nand U29383 (N_29383,N_28040,N_28863);
and U29384 (N_29384,N_28508,N_28133);
and U29385 (N_29385,N_28404,N_28207);
nand U29386 (N_29386,N_28598,N_28903);
nor U29387 (N_29387,N_28422,N_28042);
nor U29388 (N_29388,N_28693,N_28209);
and U29389 (N_29389,N_28513,N_28320);
and U29390 (N_29390,N_28180,N_28334);
and U29391 (N_29391,N_28991,N_28124);
and U29392 (N_29392,N_28524,N_28285);
xnor U29393 (N_29393,N_28846,N_28103);
and U29394 (N_29394,N_28641,N_28996);
nand U29395 (N_29395,N_28018,N_28555);
or U29396 (N_29396,N_28501,N_28504);
xnor U29397 (N_29397,N_28992,N_28227);
nor U29398 (N_29398,N_28916,N_28481);
or U29399 (N_29399,N_28543,N_28676);
nand U29400 (N_29400,N_28574,N_28934);
and U29401 (N_29401,N_28173,N_28871);
and U29402 (N_29402,N_28786,N_28961);
xnor U29403 (N_29403,N_28290,N_28313);
nand U29404 (N_29404,N_28131,N_28715);
xor U29405 (N_29405,N_28078,N_28613);
xnor U29406 (N_29406,N_28975,N_28413);
and U29407 (N_29407,N_28835,N_28272);
nor U29408 (N_29408,N_28457,N_28228);
and U29409 (N_29409,N_28458,N_28782);
nand U29410 (N_29410,N_28891,N_28807);
nand U29411 (N_29411,N_28064,N_28162);
nand U29412 (N_29412,N_28720,N_28454);
nor U29413 (N_29413,N_28165,N_28308);
nand U29414 (N_29414,N_28491,N_28882);
nor U29415 (N_29415,N_28234,N_28300);
nand U29416 (N_29416,N_28754,N_28079);
xnor U29417 (N_29417,N_28429,N_28526);
and U29418 (N_29418,N_28324,N_28068);
nor U29419 (N_29419,N_28198,N_28202);
xnor U29420 (N_29420,N_28492,N_28049);
nand U29421 (N_29421,N_28774,N_28007);
nand U29422 (N_29422,N_28607,N_28041);
nor U29423 (N_29423,N_28838,N_28070);
or U29424 (N_29424,N_28360,N_28651);
nand U29425 (N_29425,N_28775,N_28216);
or U29426 (N_29426,N_28071,N_28659);
and U29427 (N_29427,N_28215,N_28005);
or U29428 (N_29428,N_28110,N_28866);
xnor U29429 (N_29429,N_28928,N_28892);
nor U29430 (N_29430,N_28445,N_28111);
xnor U29431 (N_29431,N_28023,N_28001);
nand U29432 (N_29432,N_28879,N_28797);
nor U29433 (N_29433,N_28370,N_28414);
and U29434 (N_29434,N_28408,N_28143);
and U29435 (N_29435,N_28326,N_28544);
nor U29436 (N_29436,N_28736,N_28707);
or U29437 (N_29437,N_28037,N_28357);
and U29438 (N_29438,N_28844,N_28874);
xnor U29439 (N_29439,N_28256,N_28117);
and U29440 (N_29440,N_28628,N_28536);
or U29441 (N_29441,N_28307,N_28067);
xnor U29442 (N_29442,N_28270,N_28436);
nand U29443 (N_29443,N_28373,N_28450);
xnor U29444 (N_29444,N_28642,N_28225);
nor U29445 (N_29445,N_28483,N_28212);
or U29446 (N_29446,N_28952,N_28912);
or U29447 (N_29447,N_28282,N_28446);
xnor U29448 (N_29448,N_28986,N_28192);
nor U29449 (N_29449,N_28161,N_28779);
xnor U29450 (N_29450,N_28678,N_28894);
nand U29451 (N_29451,N_28950,N_28949);
and U29452 (N_29452,N_28691,N_28661);
xnor U29453 (N_29453,N_28611,N_28203);
and U29454 (N_29454,N_28352,N_28278);
xor U29455 (N_29455,N_28737,N_28809);
or U29456 (N_29456,N_28108,N_28390);
or U29457 (N_29457,N_28609,N_28523);
xor U29458 (N_29458,N_28141,N_28539);
nor U29459 (N_29459,N_28094,N_28399);
or U29460 (N_29460,N_28038,N_28948);
nand U29461 (N_29461,N_28723,N_28827);
nand U29462 (N_29462,N_28484,N_28339);
or U29463 (N_29463,N_28168,N_28920);
nor U29464 (N_29464,N_28090,N_28349);
nor U29465 (N_29465,N_28973,N_28667);
nor U29466 (N_29466,N_28820,N_28211);
xnor U29467 (N_29467,N_28561,N_28310);
nor U29468 (N_29468,N_28134,N_28694);
or U29469 (N_29469,N_28494,N_28944);
xnor U29470 (N_29470,N_28805,N_28170);
and U29471 (N_29471,N_28722,N_28653);
or U29472 (N_29472,N_28247,N_28476);
xor U29473 (N_29473,N_28381,N_28649);
or U29474 (N_29474,N_28902,N_28482);
nand U29475 (N_29475,N_28742,N_28514);
nor U29476 (N_29476,N_28325,N_28658);
or U29477 (N_29477,N_28615,N_28679);
nor U29478 (N_29478,N_28769,N_28867);
nand U29479 (N_29479,N_28297,N_28148);
nor U29480 (N_29480,N_28845,N_28249);
nor U29481 (N_29481,N_28685,N_28097);
nor U29482 (N_29482,N_28719,N_28680);
and U29483 (N_29483,N_28853,N_28175);
nor U29484 (N_29484,N_28123,N_28567);
nor U29485 (N_29485,N_28036,N_28136);
xnor U29486 (N_29486,N_28375,N_28614);
or U29487 (N_29487,N_28830,N_28932);
or U29488 (N_29488,N_28164,N_28434);
nand U29489 (N_29489,N_28817,N_28913);
or U29490 (N_29490,N_28084,N_28241);
nor U29491 (N_29491,N_28130,N_28629);
or U29492 (N_29492,N_28654,N_28473);
nor U29493 (N_29493,N_28335,N_28219);
xnor U29494 (N_29494,N_28011,N_28089);
xnor U29495 (N_29495,N_28569,N_28358);
or U29496 (N_29496,N_28512,N_28610);
nand U29497 (N_29497,N_28072,N_28188);
or U29498 (N_29498,N_28964,N_28224);
or U29499 (N_29499,N_28351,N_28265);
nand U29500 (N_29500,N_28030,N_28098);
nand U29501 (N_29501,N_28443,N_28598);
nand U29502 (N_29502,N_28884,N_28780);
or U29503 (N_29503,N_28431,N_28385);
or U29504 (N_29504,N_28507,N_28639);
or U29505 (N_29505,N_28074,N_28277);
xor U29506 (N_29506,N_28749,N_28748);
xnor U29507 (N_29507,N_28093,N_28016);
nand U29508 (N_29508,N_28983,N_28322);
nor U29509 (N_29509,N_28540,N_28426);
nand U29510 (N_29510,N_28927,N_28389);
or U29511 (N_29511,N_28934,N_28923);
xor U29512 (N_29512,N_28102,N_28884);
nand U29513 (N_29513,N_28460,N_28110);
xor U29514 (N_29514,N_28766,N_28796);
nor U29515 (N_29515,N_28014,N_28043);
nor U29516 (N_29516,N_28634,N_28107);
xor U29517 (N_29517,N_28677,N_28139);
nor U29518 (N_29518,N_28279,N_28317);
and U29519 (N_29519,N_28732,N_28204);
nor U29520 (N_29520,N_28214,N_28781);
nor U29521 (N_29521,N_28991,N_28546);
nor U29522 (N_29522,N_28952,N_28090);
nand U29523 (N_29523,N_28216,N_28300);
or U29524 (N_29524,N_28089,N_28827);
and U29525 (N_29525,N_28073,N_28979);
nor U29526 (N_29526,N_28565,N_28980);
nor U29527 (N_29527,N_28350,N_28331);
xor U29528 (N_29528,N_28203,N_28352);
xnor U29529 (N_29529,N_28554,N_28711);
and U29530 (N_29530,N_28254,N_28473);
xnor U29531 (N_29531,N_28511,N_28043);
nand U29532 (N_29532,N_28279,N_28675);
xor U29533 (N_29533,N_28808,N_28843);
nor U29534 (N_29534,N_28084,N_28956);
nand U29535 (N_29535,N_28299,N_28842);
and U29536 (N_29536,N_28583,N_28191);
and U29537 (N_29537,N_28404,N_28037);
nand U29538 (N_29538,N_28890,N_28124);
or U29539 (N_29539,N_28967,N_28854);
xnor U29540 (N_29540,N_28770,N_28178);
xor U29541 (N_29541,N_28990,N_28982);
nand U29542 (N_29542,N_28548,N_28783);
xor U29543 (N_29543,N_28291,N_28042);
nand U29544 (N_29544,N_28805,N_28302);
xnor U29545 (N_29545,N_28337,N_28977);
xor U29546 (N_29546,N_28389,N_28644);
nand U29547 (N_29547,N_28569,N_28930);
nand U29548 (N_29548,N_28471,N_28353);
nor U29549 (N_29549,N_28129,N_28255);
nand U29550 (N_29550,N_28543,N_28792);
or U29551 (N_29551,N_28911,N_28372);
and U29552 (N_29552,N_28036,N_28358);
xnor U29553 (N_29553,N_28933,N_28340);
nor U29554 (N_29554,N_28235,N_28422);
nand U29555 (N_29555,N_28077,N_28252);
and U29556 (N_29556,N_28777,N_28400);
xnor U29557 (N_29557,N_28830,N_28089);
xor U29558 (N_29558,N_28837,N_28982);
nor U29559 (N_29559,N_28330,N_28748);
nor U29560 (N_29560,N_28543,N_28958);
nand U29561 (N_29561,N_28495,N_28860);
and U29562 (N_29562,N_28056,N_28502);
or U29563 (N_29563,N_28504,N_28157);
xor U29564 (N_29564,N_28762,N_28206);
nand U29565 (N_29565,N_28991,N_28317);
or U29566 (N_29566,N_28596,N_28128);
nor U29567 (N_29567,N_28008,N_28738);
nor U29568 (N_29568,N_28823,N_28642);
xor U29569 (N_29569,N_28644,N_28697);
xnor U29570 (N_29570,N_28907,N_28861);
or U29571 (N_29571,N_28236,N_28307);
nor U29572 (N_29572,N_28386,N_28014);
xor U29573 (N_29573,N_28795,N_28606);
or U29574 (N_29574,N_28444,N_28212);
nor U29575 (N_29575,N_28954,N_28121);
and U29576 (N_29576,N_28722,N_28629);
nand U29577 (N_29577,N_28518,N_28865);
and U29578 (N_29578,N_28308,N_28013);
nand U29579 (N_29579,N_28813,N_28356);
xor U29580 (N_29580,N_28382,N_28847);
nand U29581 (N_29581,N_28316,N_28436);
nor U29582 (N_29582,N_28580,N_28495);
or U29583 (N_29583,N_28933,N_28277);
xnor U29584 (N_29584,N_28918,N_28095);
nor U29585 (N_29585,N_28165,N_28011);
nand U29586 (N_29586,N_28723,N_28189);
nor U29587 (N_29587,N_28126,N_28721);
and U29588 (N_29588,N_28644,N_28416);
or U29589 (N_29589,N_28056,N_28139);
nor U29590 (N_29590,N_28337,N_28496);
nand U29591 (N_29591,N_28861,N_28722);
nor U29592 (N_29592,N_28926,N_28328);
xnor U29593 (N_29593,N_28441,N_28940);
xnor U29594 (N_29594,N_28507,N_28663);
nor U29595 (N_29595,N_28132,N_28238);
and U29596 (N_29596,N_28881,N_28359);
nor U29597 (N_29597,N_28724,N_28786);
and U29598 (N_29598,N_28542,N_28532);
nor U29599 (N_29599,N_28946,N_28943);
nor U29600 (N_29600,N_28705,N_28822);
and U29601 (N_29601,N_28006,N_28956);
and U29602 (N_29602,N_28336,N_28046);
and U29603 (N_29603,N_28010,N_28470);
nand U29604 (N_29604,N_28204,N_28444);
and U29605 (N_29605,N_28989,N_28101);
and U29606 (N_29606,N_28630,N_28370);
xor U29607 (N_29607,N_28527,N_28303);
and U29608 (N_29608,N_28017,N_28251);
xnor U29609 (N_29609,N_28265,N_28445);
nor U29610 (N_29610,N_28526,N_28868);
xor U29611 (N_29611,N_28663,N_28115);
nand U29612 (N_29612,N_28297,N_28608);
xnor U29613 (N_29613,N_28449,N_28655);
nand U29614 (N_29614,N_28581,N_28430);
and U29615 (N_29615,N_28661,N_28548);
or U29616 (N_29616,N_28882,N_28496);
and U29617 (N_29617,N_28896,N_28771);
and U29618 (N_29618,N_28645,N_28406);
xnor U29619 (N_29619,N_28217,N_28777);
nor U29620 (N_29620,N_28249,N_28992);
nand U29621 (N_29621,N_28949,N_28155);
xnor U29622 (N_29622,N_28208,N_28926);
and U29623 (N_29623,N_28587,N_28776);
or U29624 (N_29624,N_28613,N_28734);
nor U29625 (N_29625,N_28266,N_28462);
xnor U29626 (N_29626,N_28959,N_28410);
nor U29627 (N_29627,N_28342,N_28463);
nor U29628 (N_29628,N_28230,N_28709);
nor U29629 (N_29629,N_28271,N_28432);
and U29630 (N_29630,N_28614,N_28991);
or U29631 (N_29631,N_28392,N_28943);
nand U29632 (N_29632,N_28850,N_28029);
xnor U29633 (N_29633,N_28624,N_28495);
and U29634 (N_29634,N_28682,N_28531);
and U29635 (N_29635,N_28655,N_28866);
nand U29636 (N_29636,N_28308,N_28044);
nand U29637 (N_29637,N_28688,N_28910);
xnor U29638 (N_29638,N_28475,N_28424);
and U29639 (N_29639,N_28898,N_28734);
nor U29640 (N_29640,N_28219,N_28626);
nand U29641 (N_29641,N_28077,N_28034);
nand U29642 (N_29642,N_28477,N_28761);
xor U29643 (N_29643,N_28400,N_28128);
or U29644 (N_29644,N_28343,N_28252);
and U29645 (N_29645,N_28579,N_28194);
nand U29646 (N_29646,N_28879,N_28974);
or U29647 (N_29647,N_28591,N_28428);
nor U29648 (N_29648,N_28088,N_28159);
nor U29649 (N_29649,N_28196,N_28089);
or U29650 (N_29650,N_28068,N_28070);
and U29651 (N_29651,N_28533,N_28274);
and U29652 (N_29652,N_28157,N_28675);
and U29653 (N_29653,N_28311,N_28873);
nand U29654 (N_29654,N_28111,N_28154);
or U29655 (N_29655,N_28510,N_28480);
or U29656 (N_29656,N_28180,N_28784);
or U29657 (N_29657,N_28547,N_28582);
xnor U29658 (N_29658,N_28784,N_28930);
and U29659 (N_29659,N_28051,N_28335);
xnor U29660 (N_29660,N_28575,N_28529);
nor U29661 (N_29661,N_28672,N_28374);
xor U29662 (N_29662,N_28761,N_28062);
or U29663 (N_29663,N_28354,N_28824);
xor U29664 (N_29664,N_28442,N_28395);
or U29665 (N_29665,N_28807,N_28814);
or U29666 (N_29666,N_28801,N_28005);
or U29667 (N_29667,N_28761,N_28704);
nand U29668 (N_29668,N_28506,N_28294);
nor U29669 (N_29669,N_28637,N_28571);
nand U29670 (N_29670,N_28126,N_28256);
xor U29671 (N_29671,N_28836,N_28028);
xnor U29672 (N_29672,N_28448,N_28650);
or U29673 (N_29673,N_28577,N_28534);
or U29674 (N_29674,N_28591,N_28736);
nor U29675 (N_29675,N_28637,N_28596);
nand U29676 (N_29676,N_28265,N_28200);
or U29677 (N_29677,N_28447,N_28593);
xnor U29678 (N_29678,N_28088,N_28454);
nor U29679 (N_29679,N_28087,N_28369);
nand U29680 (N_29680,N_28408,N_28367);
nand U29681 (N_29681,N_28166,N_28092);
nand U29682 (N_29682,N_28712,N_28586);
nor U29683 (N_29683,N_28081,N_28988);
and U29684 (N_29684,N_28913,N_28743);
nand U29685 (N_29685,N_28375,N_28797);
and U29686 (N_29686,N_28287,N_28842);
or U29687 (N_29687,N_28453,N_28533);
or U29688 (N_29688,N_28450,N_28928);
nor U29689 (N_29689,N_28343,N_28841);
nor U29690 (N_29690,N_28279,N_28895);
or U29691 (N_29691,N_28666,N_28724);
or U29692 (N_29692,N_28979,N_28014);
nand U29693 (N_29693,N_28057,N_28732);
and U29694 (N_29694,N_28805,N_28147);
and U29695 (N_29695,N_28296,N_28959);
and U29696 (N_29696,N_28860,N_28143);
or U29697 (N_29697,N_28124,N_28448);
and U29698 (N_29698,N_28045,N_28857);
and U29699 (N_29699,N_28554,N_28377);
nand U29700 (N_29700,N_28974,N_28514);
nor U29701 (N_29701,N_28803,N_28372);
or U29702 (N_29702,N_28052,N_28907);
nor U29703 (N_29703,N_28825,N_28340);
or U29704 (N_29704,N_28365,N_28588);
xnor U29705 (N_29705,N_28490,N_28759);
xnor U29706 (N_29706,N_28275,N_28024);
nand U29707 (N_29707,N_28525,N_28128);
and U29708 (N_29708,N_28661,N_28962);
xor U29709 (N_29709,N_28377,N_28068);
nand U29710 (N_29710,N_28953,N_28972);
xnor U29711 (N_29711,N_28480,N_28973);
nor U29712 (N_29712,N_28629,N_28340);
nor U29713 (N_29713,N_28750,N_28049);
and U29714 (N_29714,N_28474,N_28060);
nor U29715 (N_29715,N_28198,N_28932);
and U29716 (N_29716,N_28606,N_28413);
nor U29717 (N_29717,N_28306,N_28095);
or U29718 (N_29718,N_28353,N_28284);
xnor U29719 (N_29719,N_28666,N_28159);
and U29720 (N_29720,N_28708,N_28683);
or U29721 (N_29721,N_28416,N_28346);
nor U29722 (N_29722,N_28251,N_28193);
and U29723 (N_29723,N_28619,N_28268);
xnor U29724 (N_29724,N_28913,N_28919);
and U29725 (N_29725,N_28679,N_28065);
and U29726 (N_29726,N_28742,N_28718);
nor U29727 (N_29727,N_28881,N_28369);
nor U29728 (N_29728,N_28790,N_28254);
nor U29729 (N_29729,N_28708,N_28935);
or U29730 (N_29730,N_28821,N_28515);
nor U29731 (N_29731,N_28266,N_28622);
xnor U29732 (N_29732,N_28880,N_28494);
xnor U29733 (N_29733,N_28562,N_28308);
xor U29734 (N_29734,N_28165,N_28477);
nor U29735 (N_29735,N_28290,N_28223);
nor U29736 (N_29736,N_28866,N_28965);
nand U29737 (N_29737,N_28374,N_28593);
or U29738 (N_29738,N_28050,N_28490);
nor U29739 (N_29739,N_28108,N_28609);
nor U29740 (N_29740,N_28844,N_28885);
and U29741 (N_29741,N_28147,N_28883);
nor U29742 (N_29742,N_28541,N_28346);
nand U29743 (N_29743,N_28189,N_28558);
nor U29744 (N_29744,N_28215,N_28611);
nor U29745 (N_29745,N_28260,N_28834);
nand U29746 (N_29746,N_28234,N_28177);
nor U29747 (N_29747,N_28133,N_28370);
and U29748 (N_29748,N_28602,N_28020);
or U29749 (N_29749,N_28219,N_28652);
nand U29750 (N_29750,N_28312,N_28401);
nor U29751 (N_29751,N_28140,N_28467);
nor U29752 (N_29752,N_28928,N_28454);
xnor U29753 (N_29753,N_28673,N_28668);
nand U29754 (N_29754,N_28656,N_28902);
nor U29755 (N_29755,N_28446,N_28522);
xor U29756 (N_29756,N_28200,N_28960);
and U29757 (N_29757,N_28269,N_28923);
nor U29758 (N_29758,N_28427,N_28518);
xor U29759 (N_29759,N_28303,N_28143);
nand U29760 (N_29760,N_28225,N_28882);
or U29761 (N_29761,N_28316,N_28799);
xor U29762 (N_29762,N_28303,N_28880);
nand U29763 (N_29763,N_28396,N_28040);
xnor U29764 (N_29764,N_28216,N_28194);
or U29765 (N_29765,N_28069,N_28158);
nor U29766 (N_29766,N_28361,N_28430);
nor U29767 (N_29767,N_28383,N_28931);
nor U29768 (N_29768,N_28230,N_28188);
nand U29769 (N_29769,N_28615,N_28039);
nand U29770 (N_29770,N_28718,N_28600);
nand U29771 (N_29771,N_28597,N_28153);
xor U29772 (N_29772,N_28314,N_28472);
xnor U29773 (N_29773,N_28329,N_28624);
nor U29774 (N_29774,N_28452,N_28061);
xnor U29775 (N_29775,N_28704,N_28808);
nand U29776 (N_29776,N_28740,N_28880);
or U29777 (N_29777,N_28786,N_28449);
xor U29778 (N_29778,N_28687,N_28119);
or U29779 (N_29779,N_28358,N_28144);
and U29780 (N_29780,N_28842,N_28158);
nor U29781 (N_29781,N_28248,N_28570);
and U29782 (N_29782,N_28385,N_28719);
xnor U29783 (N_29783,N_28450,N_28370);
nor U29784 (N_29784,N_28601,N_28917);
nand U29785 (N_29785,N_28089,N_28239);
xor U29786 (N_29786,N_28526,N_28658);
nor U29787 (N_29787,N_28828,N_28680);
and U29788 (N_29788,N_28693,N_28792);
nand U29789 (N_29789,N_28647,N_28238);
and U29790 (N_29790,N_28181,N_28707);
or U29791 (N_29791,N_28854,N_28840);
or U29792 (N_29792,N_28656,N_28459);
nor U29793 (N_29793,N_28139,N_28897);
nand U29794 (N_29794,N_28308,N_28039);
and U29795 (N_29795,N_28506,N_28869);
and U29796 (N_29796,N_28665,N_28320);
or U29797 (N_29797,N_28745,N_28771);
or U29798 (N_29798,N_28342,N_28959);
xnor U29799 (N_29799,N_28300,N_28634);
nor U29800 (N_29800,N_28145,N_28174);
and U29801 (N_29801,N_28538,N_28027);
and U29802 (N_29802,N_28960,N_28998);
nor U29803 (N_29803,N_28794,N_28204);
nand U29804 (N_29804,N_28047,N_28908);
nor U29805 (N_29805,N_28123,N_28722);
or U29806 (N_29806,N_28107,N_28158);
or U29807 (N_29807,N_28078,N_28426);
or U29808 (N_29808,N_28521,N_28805);
nor U29809 (N_29809,N_28301,N_28827);
xor U29810 (N_29810,N_28770,N_28132);
nor U29811 (N_29811,N_28078,N_28259);
or U29812 (N_29812,N_28012,N_28892);
xor U29813 (N_29813,N_28999,N_28735);
or U29814 (N_29814,N_28726,N_28200);
and U29815 (N_29815,N_28168,N_28407);
nand U29816 (N_29816,N_28591,N_28010);
or U29817 (N_29817,N_28840,N_28311);
nand U29818 (N_29818,N_28628,N_28017);
and U29819 (N_29819,N_28409,N_28141);
nor U29820 (N_29820,N_28834,N_28627);
nor U29821 (N_29821,N_28695,N_28597);
or U29822 (N_29822,N_28597,N_28166);
nand U29823 (N_29823,N_28564,N_28417);
nor U29824 (N_29824,N_28246,N_28854);
and U29825 (N_29825,N_28320,N_28349);
nor U29826 (N_29826,N_28117,N_28325);
xor U29827 (N_29827,N_28144,N_28632);
nand U29828 (N_29828,N_28582,N_28369);
nor U29829 (N_29829,N_28646,N_28005);
xor U29830 (N_29830,N_28248,N_28782);
and U29831 (N_29831,N_28996,N_28084);
nand U29832 (N_29832,N_28102,N_28486);
and U29833 (N_29833,N_28497,N_28110);
nor U29834 (N_29834,N_28945,N_28485);
and U29835 (N_29835,N_28952,N_28588);
and U29836 (N_29836,N_28421,N_28385);
xor U29837 (N_29837,N_28812,N_28339);
or U29838 (N_29838,N_28026,N_28807);
nand U29839 (N_29839,N_28795,N_28987);
or U29840 (N_29840,N_28680,N_28117);
xnor U29841 (N_29841,N_28314,N_28221);
and U29842 (N_29842,N_28457,N_28485);
xor U29843 (N_29843,N_28701,N_28423);
or U29844 (N_29844,N_28527,N_28996);
nor U29845 (N_29845,N_28957,N_28435);
nand U29846 (N_29846,N_28478,N_28990);
or U29847 (N_29847,N_28884,N_28689);
xor U29848 (N_29848,N_28977,N_28454);
or U29849 (N_29849,N_28960,N_28465);
nor U29850 (N_29850,N_28188,N_28351);
or U29851 (N_29851,N_28285,N_28821);
and U29852 (N_29852,N_28559,N_28077);
and U29853 (N_29853,N_28759,N_28783);
xnor U29854 (N_29854,N_28342,N_28550);
or U29855 (N_29855,N_28462,N_28654);
nor U29856 (N_29856,N_28755,N_28034);
or U29857 (N_29857,N_28296,N_28350);
nor U29858 (N_29858,N_28689,N_28645);
nor U29859 (N_29859,N_28065,N_28159);
xor U29860 (N_29860,N_28856,N_28090);
nor U29861 (N_29861,N_28573,N_28636);
nand U29862 (N_29862,N_28202,N_28011);
and U29863 (N_29863,N_28338,N_28915);
nor U29864 (N_29864,N_28850,N_28974);
nor U29865 (N_29865,N_28700,N_28981);
nand U29866 (N_29866,N_28234,N_28038);
nand U29867 (N_29867,N_28269,N_28028);
or U29868 (N_29868,N_28432,N_28884);
nand U29869 (N_29869,N_28190,N_28107);
and U29870 (N_29870,N_28537,N_28826);
xor U29871 (N_29871,N_28229,N_28027);
nand U29872 (N_29872,N_28245,N_28355);
xor U29873 (N_29873,N_28674,N_28666);
nand U29874 (N_29874,N_28169,N_28634);
and U29875 (N_29875,N_28605,N_28112);
xor U29876 (N_29876,N_28175,N_28832);
xnor U29877 (N_29877,N_28541,N_28207);
nand U29878 (N_29878,N_28993,N_28780);
or U29879 (N_29879,N_28010,N_28621);
or U29880 (N_29880,N_28260,N_28211);
xnor U29881 (N_29881,N_28710,N_28640);
nor U29882 (N_29882,N_28845,N_28814);
nor U29883 (N_29883,N_28462,N_28460);
or U29884 (N_29884,N_28728,N_28316);
or U29885 (N_29885,N_28066,N_28709);
or U29886 (N_29886,N_28778,N_28245);
nand U29887 (N_29887,N_28311,N_28910);
and U29888 (N_29888,N_28509,N_28374);
xor U29889 (N_29889,N_28881,N_28338);
nor U29890 (N_29890,N_28782,N_28670);
nand U29891 (N_29891,N_28671,N_28489);
nand U29892 (N_29892,N_28581,N_28217);
nand U29893 (N_29893,N_28143,N_28331);
nor U29894 (N_29894,N_28436,N_28859);
or U29895 (N_29895,N_28333,N_28165);
xor U29896 (N_29896,N_28205,N_28256);
xor U29897 (N_29897,N_28435,N_28476);
and U29898 (N_29898,N_28266,N_28459);
or U29899 (N_29899,N_28929,N_28667);
nor U29900 (N_29900,N_28818,N_28432);
and U29901 (N_29901,N_28686,N_28178);
and U29902 (N_29902,N_28108,N_28185);
nand U29903 (N_29903,N_28100,N_28016);
or U29904 (N_29904,N_28919,N_28002);
nor U29905 (N_29905,N_28874,N_28713);
xor U29906 (N_29906,N_28457,N_28420);
nand U29907 (N_29907,N_28793,N_28911);
and U29908 (N_29908,N_28880,N_28258);
xnor U29909 (N_29909,N_28204,N_28917);
and U29910 (N_29910,N_28141,N_28035);
nor U29911 (N_29911,N_28807,N_28753);
xnor U29912 (N_29912,N_28023,N_28839);
nor U29913 (N_29913,N_28119,N_28393);
xnor U29914 (N_29914,N_28353,N_28814);
or U29915 (N_29915,N_28800,N_28764);
nor U29916 (N_29916,N_28184,N_28295);
nand U29917 (N_29917,N_28609,N_28976);
nand U29918 (N_29918,N_28705,N_28442);
and U29919 (N_29919,N_28288,N_28303);
nand U29920 (N_29920,N_28316,N_28147);
nand U29921 (N_29921,N_28004,N_28891);
or U29922 (N_29922,N_28717,N_28467);
or U29923 (N_29923,N_28058,N_28103);
nor U29924 (N_29924,N_28678,N_28083);
or U29925 (N_29925,N_28481,N_28089);
nand U29926 (N_29926,N_28098,N_28072);
nand U29927 (N_29927,N_28480,N_28683);
nor U29928 (N_29928,N_28762,N_28550);
or U29929 (N_29929,N_28610,N_28014);
and U29930 (N_29930,N_28831,N_28241);
nor U29931 (N_29931,N_28421,N_28978);
xor U29932 (N_29932,N_28955,N_28635);
nand U29933 (N_29933,N_28948,N_28908);
or U29934 (N_29934,N_28636,N_28784);
nor U29935 (N_29935,N_28386,N_28153);
xnor U29936 (N_29936,N_28869,N_28868);
or U29937 (N_29937,N_28196,N_28308);
and U29938 (N_29938,N_28189,N_28846);
nand U29939 (N_29939,N_28111,N_28633);
or U29940 (N_29940,N_28258,N_28124);
xor U29941 (N_29941,N_28287,N_28475);
xor U29942 (N_29942,N_28945,N_28565);
xnor U29943 (N_29943,N_28618,N_28599);
or U29944 (N_29944,N_28404,N_28731);
or U29945 (N_29945,N_28366,N_28826);
xor U29946 (N_29946,N_28367,N_28946);
nor U29947 (N_29947,N_28569,N_28183);
nor U29948 (N_29948,N_28042,N_28302);
nand U29949 (N_29949,N_28955,N_28028);
or U29950 (N_29950,N_28710,N_28337);
xor U29951 (N_29951,N_28028,N_28424);
xnor U29952 (N_29952,N_28457,N_28546);
and U29953 (N_29953,N_28470,N_28486);
and U29954 (N_29954,N_28276,N_28417);
nor U29955 (N_29955,N_28434,N_28107);
and U29956 (N_29956,N_28469,N_28181);
xnor U29957 (N_29957,N_28307,N_28746);
or U29958 (N_29958,N_28648,N_28342);
nand U29959 (N_29959,N_28015,N_28755);
nor U29960 (N_29960,N_28501,N_28162);
nor U29961 (N_29961,N_28725,N_28661);
nor U29962 (N_29962,N_28841,N_28753);
or U29963 (N_29963,N_28121,N_28841);
and U29964 (N_29964,N_28296,N_28577);
or U29965 (N_29965,N_28397,N_28904);
xor U29966 (N_29966,N_28549,N_28227);
or U29967 (N_29967,N_28631,N_28085);
xor U29968 (N_29968,N_28264,N_28243);
and U29969 (N_29969,N_28062,N_28944);
nand U29970 (N_29970,N_28226,N_28891);
nand U29971 (N_29971,N_28587,N_28044);
or U29972 (N_29972,N_28892,N_28624);
nor U29973 (N_29973,N_28805,N_28173);
and U29974 (N_29974,N_28695,N_28890);
nand U29975 (N_29975,N_28945,N_28599);
or U29976 (N_29976,N_28447,N_28245);
and U29977 (N_29977,N_28863,N_28293);
nor U29978 (N_29978,N_28946,N_28690);
xnor U29979 (N_29979,N_28300,N_28009);
nor U29980 (N_29980,N_28243,N_28589);
nor U29981 (N_29981,N_28199,N_28251);
nor U29982 (N_29982,N_28702,N_28108);
and U29983 (N_29983,N_28236,N_28680);
or U29984 (N_29984,N_28248,N_28866);
or U29985 (N_29985,N_28411,N_28929);
nor U29986 (N_29986,N_28678,N_28018);
or U29987 (N_29987,N_28621,N_28827);
and U29988 (N_29988,N_28907,N_28019);
and U29989 (N_29989,N_28224,N_28646);
or U29990 (N_29990,N_28653,N_28775);
nand U29991 (N_29991,N_28072,N_28531);
nand U29992 (N_29992,N_28198,N_28239);
xor U29993 (N_29993,N_28919,N_28601);
xor U29994 (N_29994,N_28822,N_28411);
nand U29995 (N_29995,N_28841,N_28213);
or U29996 (N_29996,N_28379,N_28024);
or U29997 (N_29997,N_28967,N_28579);
or U29998 (N_29998,N_28933,N_28458);
nor U29999 (N_29999,N_28917,N_28563);
nand U30000 (N_30000,N_29929,N_29633);
nand U30001 (N_30001,N_29172,N_29907);
nor U30002 (N_30002,N_29819,N_29161);
or U30003 (N_30003,N_29806,N_29669);
nor U30004 (N_30004,N_29079,N_29538);
and U30005 (N_30005,N_29371,N_29195);
nor U30006 (N_30006,N_29096,N_29511);
xnor U30007 (N_30007,N_29299,N_29621);
nor U30008 (N_30008,N_29211,N_29736);
nand U30009 (N_30009,N_29137,N_29495);
nor U30010 (N_30010,N_29175,N_29998);
nor U30011 (N_30011,N_29198,N_29729);
xnor U30012 (N_30012,N_29493,N_29710);
xnor U30013 (N_30013,N_29178,N_29758);
and U30014 (N_30014,N_29537,N_29273);
nor U30015 (N_30015,N_29242,N_29999);
xnor U30016 (N_30016,N_29612,N_29312);
or U30017 (N_30017,N_29001,N_29958);
nor U30018 (N_30018,N_29107,N_29858);
nor U30019 (N_30019,N_29184,N_29580);
or U30020 (N_30020,N_29038,N_29446);
or U30021 (N_30021,N_29237,N_29264);
and U30022 (N_30022,N_29465,N_29798);
xor U30023 (N_30023,N_29123,N_29149);
xnor U30024 (N_30024,N_29368,N_29268);
nor U30025 (N_30025,N_29704,N_29221);
nor U30026 (N_30026,N_29277,N_29201);
nor U30027 (N_30027,N_29048,N_29434);
xor U30028 (N_30028,N_29988,N_29638);
and U30029 (N_30029,N_29564,N_29678);
and U30030 (N_30030,N_29406,N_29063);
or U30031 (N_30031,N_29786,N_29481);
and U30032 (N_30032,N_29934,N_29711);
or U30033 (N_30033,N_29046,N_29941);
and U30034 (N_30034,N_29218,N_29088);
xor U30035 (N_30035,N_29724,N_29730);
or U30036 (N_30036,N_29637,N_29336);
and U30037 (N_30037,N_29008,N_29219);
or U30038 (N_30038,N_29895,N_29940);
xnor U30039 (N_30039,N_29438,N_29015);
and U30040 (N_30040,N_29106,N_29668);
nand U30041 (N_30041,N_29192,N_29332);
nor U30042 (N_30042,N_29548,N_29270);
xnor U30043 (N_30043,N_29334,N_29304);
nand U30044 (N_30044,N_29550,N_29810);
and U30045 (N_30045,N_29631,N_29333);
nor U30046 (N_30046,N_29171,N_29418);
nand U30047 (N_30047,N_29040,N_29595);
nor U30048 (N_30048,N_29148,N_29413);
xnor U30049 (N_30049,N_29759,N_29900);
nand U30050 (N_30050,N_29365,N_29712);
nor U30051 (N_30051,N_29665,N_29426);
nor U30052 (N_30052,N_29177,N_29379);
xnor U30053 (N_30053,N_29142,N_29878);
nor U30054 (N_30054,N_29214,N_29340);
or U30055 (N_30055,N_29582,N_29656);
nor U30056 (N_30056,N_29473,N_29628);
nand U30057 (N_30057,N_29479,N_29186);
nor U30058 (N_30058,N_29714,N_29540);
or U30059 (N_30059,N_29374,N_29154);
and U30060 (N_30060,N_29609,N_29357);
or U30061 (N_30061,N_29830,N_29667);
or U30062 (N_30062,N_29728,N_29429);
nand U30063 (N_30063,N_29308,N_29743);
or U30064 (N_30064,N_29098,N_29875);
nand U30065 (N_30065,N_29187,N_29838);
and U30066 (N_30066,N_29698,N_29771);
nor U30067 (N_30067,N_29833,N_29501);
nor U30068 (N_30068,N_29660,N_29859);
nand U30069 (N_30069,N_29155,N_29468);
or U30070 (N_30070,N_29984,N_29132);
or U30071 (N_30071,N_29947,N_29459);
nand U30072 (N_30072,N_29715,N_29274);
nor U30073 (N_30073,N_29347,N_29938);
or U30074 (N_30074,N_29824,N_29441);
nand U30075 (N_30075,N_29247,N_29167);
nand U30076 (N_30076,N_29065,N_29885);
nand U30077 (N_30077,N_29381,N_29975);
nor U30078 (N_30078,N_29395,N_29645);
xnor U30079 (N_30079,N_29185,N_29653);
xnor U30080 (N_30080,N_29352,N_29007);
or U30081 (N_30081,N_29593,N_29639);
nand U30082 (N_30082,N_29453,N_29574);
or U30083 (N_30083,N_29809,N_29752);
and U30084 (N_30084,N_29452,N_29377);
xor U30085 (N_30085,N_29706,N_29544);
nor U30086 (N_30086,N_29145,N_29579);
and U30087 (N_30087,N_29094,N_29541);
nand U30088 (N_30088,N_29422,N_29045);
xor U30089 (N_30089,N_29419,N_29363);
nor U30090 (N_30090,N_29217,N_29222);
and U30091 (N_30091,N_29694,N_29671);
nand U30092 (N_30092,N_29158,N_29474);
xor U30093 (N_30093,N_29234,N_29269);
or U30094 (N_30094,N_29647,N_29971);
nor U30095 (N_30095,N_29284,N_29525);
and U30096 (N_30096,N_29071,N_29014);
or U30097 (N_30097,N_29839,N_29405);
or U30098 (N_30098,N_29262,N_29613);
nand U30099 (N_30099,N_29636,N_29910);
or U30100 (N_30100,N_29753,N_29361);
xor U30101 (N_30101,N_29303,N_29616);
and U30102 (N_30102,N_29103,N_29233);
and U30103 (N_30103,N_29112,N_29762);
and U30104 (N_30104,N_29049,N_29510);
or U30105 (N_30105,N_29913,N_29569);
nand U30106 (N_30106,N_29527,N_29925);
or U30107 (N_30107,N_29995,N_29433);
nor U30108 (N_30108,N_29436,N_29399);
and U30109 (N_30109,N_29089,N_29487);
and U30110 (N_30110,N_29116,N_29006);
nand U30111 (N_30111,N_29129,N_29298);
nor U30112 (N_30112,N_29200,N_29632);
nand U30113 (N_30113,N_29985,N_29174);
nand U30114 (N_30114,N_29119,N_29834);
nor U30115 (N_30115,N_29283,N_29323);
nand U30116 (N_30116,N_29981,N_29029);
and U30117 (N_30117,N_29111,N_29570);
and U30118 (N_30118,N_29781,N_29605);
nand U30119 (N_30119,N_29393,N_29249);
nand U30120 (N_30120,N_29402,N_29165);
xnor U30121 (N_30121,N_29814,N_29004);
xor U30122 (N_30122,N_29757,N_29542);
xnor U30123 (N_30123,N_29607,N_29194);
nand U30124 (N_30124,N_29850,N_29276);
nand U30125 (N_30125,N_29944,N_29017);
or U30126 (N_30126,N_29254,N_29733);
nor U30127 (N_30127,N_29560,N_29231);
or U30128 (N_30128,N_29568,N_29414);
or U30129 (N_30129,N_29403,N_29488);
nand U30130 (N_30130,N_29326,N_29589);
nand U30131 (N_30131,N_29735,N_29412);
xnor U30132 (N_30132,N_29444,N_29756);
and U30133 (N_30133,N_29914,N_29275);
and U30134 (N_30134,N_29904,N_29416);
nor U30135 (N_30135,N_29902,N_29421);
nand U30136 (N_30136,N_29070,N_29443);
nor U30137 (N_30137,N_29372,N_29024);
and U30138 (N_30138,N_29003,N_29844);
nand U30139 (N_30139,N_29257,N_29294);
xor U30140 (N_30140,N_29673,N_29974);
xor U30141 (N_30141,N_29573,N_29448);
and U30142 (N_30142,N_29871,N_29597);
or U30143 (N_30143,N_29250,N_29193);
nor U30144 (N_30144,N_29445,N_29462);
nor U30145 (N_30145,N_29311,N_29518);
and U30146 (N_30146,N_29770,N_29396);
nor U30147 (N_30147,N_29266,N_29338);
or U30148 (N_30148,N_29253,N_29846);
and U30149 (N_30149,N_29457,N_29500);
xor U30150 (N_30150,N_29239,N_29091);
xnor U30151 (N_30151,N_29788,N_29783);
nor U30152 (N_30152,N_29815,N_29558);
or U30153 (N_30153,N_29203,N_29033);
and U30154 (N_30154,N_29061,N_29562);
nor U30155 (N_30155,N_29872,N_29932);
and U30156 (N_30156,N_29853,N_29800);
xnor U30157 (N_30157,N_29695,N_29220);
or U30158 (N_30158,N_29686,N_29880);
nor U30159 (N_30159,N_29258,N_29751);
xor U30160 (N_30160,N_29288,N_29471);
xor U30161 (N_30161,N_29847,N_29476);
or U30162 (N_30162,N_29344,N_29851);
or U30163 (N_30163,N_29674,N_29320);
xnor U30164 (N_30164,N_29764,N_29852);
nor U30165 (N_30165,N_29391,N_29987);
and U30166 (N_30166,N_29328,N_29078);
nand U30167 (N_30167,N_29967,N_29108);
or U30168 (N_30168,N_29962,N_29489);
xnor U30169 (N_30169,N_29528,N_29069);
and U30170 (N_30170,N_29627,N_29169);
and U30171 (N_30171,N_29390,N_29845);
and U30172 (N_30172,N_29105,N_29989);
and U30173 (N_30173,N_29747,N_29207);
nor U30174 (N_30174,N_29230,N_29292);
nand U30175 (N_30175,N_29848,N_29077);
and U30176 (N_30176,N_29901,N_29497);
xnor U30177 (N_30177,N_29397,N_29888);
nor U30178 (N_30178,N_29050,N_29491);
nor U30179 (N_30179,N_29725,N_29652);
or U30180 (N_30180,N_29212,N_29521);
or U30181 (N_30181,N_29869,N_29930);
nand U30182 (N_30182,N_29480,N_29252);
and U30183 (N_30183,N_29547,N_29028);
or U30184 (N_30184,N_29796,N_29963);
or U30185 (N_30185,N_29583,N_29530);
or U30186 (N_30186,N_29509,N_29191);
nand U30187 (N_30187,N_29622,N_29196);
and U30188 (N_30188,N_29842,N_29013);
xor U30189 (N_30189,N_29255,N_29654);
nand U30190 (N_30190,N_29949,N_29456);
xor U30191 (N_30191,N_29586,N_29532);
xor U30192 (N_30192,N_29310,N_29978);
nor U30193 (N_30193,N_29055,N_29097);
nand U30194 (N_30194,N_29437,N_29227);
nor U30195 (N_30195,N_29507,N_29359);
and U30196 (N_30196,N_29209,N_29829);
or U30197 (N_30197,N_29047,N_29110);
nor U30198 (N_30198,N_29716,N_29064);
or U30199 (N_30199,N_29517,N_29068);
and U30200 (N_30200,N_29820,N_29943);
or U30201 (N_30201,N_29290,N_29401);
nand U30202 (N_30202,N_29857,N_29778);
nor U30203 (N_30203,N_29058,N_29703);
xnor U30204 (N_30204,N_29140,N_29713);
and U30205 (N_30205,N_29442,N_29021);
or U30206 (N_30206,N_29279,N_29225);
nand U30207 (N_30207,N_29828,N_29862);
or U30208 (N_30208,N_29486,N_29120);
and U30209 (N_30209,N_29346,N_29982);
xor U30210 (N_30210,N_29976,N_29827);
nor U30211 (N_30211,N_29494,N_29546);
or U30212 (N_30212,N_29794,N_29331);
nand U30213 (N_30213,N_29926,N_29977);
xnor U30214 (N_30214,N_29409,N_29319);
or U30215 (N_30215,N_29650,N_29166);
and U30216 (N_30216,N_29012,N_29923);
nor U30217 (N_30217,N_29832,N_29935);
xor U30218 (N_30218,N_29018,N_29036);
xnor U30219 (N_30219,N_29953,N_29629);
nor U30220 (N_30220,N_29937,N_29555);
nand U30221 (N_30221,N_29948,N_29305);
nor U30222 (N_30222,N_29229,N_29520);
or U30223 (N_30223,N_29818,N_29883);
and U30224 (N_30224,N_29327,N_29043);
or U30225 (N_30225,N_29460,N_29378);
xnor U30226 (N_30226,N_29927,N_29911);
or U30227 (N_30227,N_29676,N_29408);
or U30228 (N_30228,N_29490,N_29080);
nor U30229 (N_30229,N_29278,N_29567);
nor U30230 (N_30230,N_29643,N_29435);
or U30231 (N_30231,N_29354,N_29738);
or U30232 (N_30232,N_29610,N_29826);
or U30233 (N_30233,N_29960,N_29246);
nor U30234 (N_30234,N_29228,N_29150);
xnor U30235 (N_30235,N_29990,N_29243);
xor U30236 (N_30236,N_29866,N_29876);
xnor U30237 (N_30237,N_29113,N_29956);
or U30238 (N_30238,N_29614,N_29640);
nor U30239 (N_30239,N_29691,N_29626);
nor U30240 (N_30240,N_29179,N_29973);
nor U30241 (N_30241,N_29646,N_29594);
nor U30242 (N_30242,N_29223,N_29325);
and U30243 (N_30243,N_29513,N_29463);
nand U30244 (N_30244,N_29649,N_29514);
nand U30245 (N_30245,N_29461,N_29536);
xor U30246 (N_30246,N_29141,N_29916);
or U30247 (N_30247,N_29519,N_29804);
nor U30248 (N_30248,N_29469,N_29625);
xnor U30249 (N_30249,N_29075,N_29543);
or U30250 (N_30250,N_29240,N_29767);
nor U30251 (N_30251,N_29915,N_29924);
nand U30252 (N_30252,N_29604,N_29019);
or U30253 (N_30253,N_29727,N_29950);
xor U30254 (N_30254,N_29590,N_29611);
nand U30255 (N_30255,N_29182,N_29251);
nand U30256 (N_30256,N_29600,N_29765);
or U30257 (N_30257,N_29076,N_29856);
xnor U30258 (N_30258,N_29657,N_29799);
or U30259 (N_30259,N_29921,N_29159);
and U30260 (N_30260,N_29143,N_29744);
nor U30261 (N_30261,N_29306,N_29084);
nor U30262 (N_30262,N_29533,N_29210);
nand U30263 (N_30263,N_29109,N_29700);
or U30264 (N_30264,N_29134,N_29267);
or U30265 (N_30265,N_29034,N_29183);
nor U30266 (N_30266,N_29282,N_29369);
or U30267 (N_30267,N_29271,N_29873);
xor U30268 (N_30268,N_29585,N_29300);
nor U30269 (N_30269,N_29572,N_29843);
nand U30270 (N_30270,N_29606,N_29085);
or U30271 (N_30271,N_29118,N_29245);
nand U30272 (N_30272,N_29531,N_29659);
or U30273 (N_30273,N_29499,N_29717);
nor U30274 (N_30274,N_29086,N_29483);
xnor U30275 (N_30275,N_29529,N_29959);
nor U30276 (N_30276,N_29877,N_29782);
and U30277 (N_30277,N_29933,N_29072);
and U30278 (N_30278,N_29411,N_29054);
nor U30279 (N_30279,N_29708,N_29400);
xnor U30280 (N_30280,N_29115,N_29905);
nand U30281 (N_30281,N_29746,N_29919);
nand U30282 (N_30282,N_29451,N_29503);
xor U30283 (N_30283,N_29389,N_29741);
and U30284 (N_30284,N_29942,N_29887);
xnor U30285 (N_30285,N_29152,N_29351);
and U30286 (N_30286,N_29057,N_29260);
nor U30287 (N_30287,N_29188,N_29502);
and U30288 (N_30288,N_29232,N_29440);
xor U30289 (N_30289,N_29394,N_29101);
nand U30290 (N_30290,N_29670,N_29144);
and U30291 (N_30291,N_29053,N_29592);
nand U30292 (N_30292,N_29742,N_29983);
nand U30293 (N_30293,N_29126,N_29130);
nor U30294 (N_30294,N_29428,N_29367);
or U30295 (N_30295,N_29335,N_29176);
xor U30296 (N_30296,N_29163,N_29749);
nor U30297 (N_30297,N_29404,N_29472);
nor U30298 (N_30298,N_29970,N_29748);
xor U30299 (N_30299,N_29138,N_29965);
nand U30300 (N_30300,N_29690,N_29601);
nor U30301 (N_30301,N_29863,N_29577);
nor U30302 (N_30302,N_29566,N_29791);
nor U30303 (N_30303,N_29993,N_29860);
nand U30304 (N_30304,N_29512,N_29787);
nand U30305 (N_30305,N_29807,N_29350);
xor U30306 (N_30306,N_29624,N_29127);
or U30307 (N_30307,N_29563,N_29726);
or U30308 (N_30308,N_29370,N_29615);
nor U30309 (N_30309,N_29994,N_29755);
nand U30310 (N_30310,N_29296,N_29321);
or U30311 (N_30311,N_29467,N_29802);
or U30312 (N_30312,N_29215,N_29897);
or U30313 (N_30313,N_29032,N_29432);
or U30314 (N_30314,N_29343,N_29881);
nor U30315 (N_30315,N_29893,N_29383);
or U30316 (N_30316,N_29651,N_29868);
nand U30317 (N_30317,N_29737,N_29630);
or U30318 (N_30318,N_29516,N_29526);
xnor U30319 (N_30319,N_29324,N_29458);
and U30320 (N_30320,N_29693,N_29552);
nand U30321 (N_30321,N_29153,N_29202);
xor U30322 (N_30322,N_29557,N_29482);
and U30323 (N_30323,N_29156,N_29505);
nor U30324 (N_30324,N_29882,N_29979);
nor U30325 (N_30325,N_29297,N_29889);
or U30326 (N_30326,N_29576,N_29855);
xnor U30327 (N_30327,N_29301,N_29385);
nor U30328 (N_30328,N_29362,N_29092);
and U30329 (N_30329,N_29235,N_29470);
or U30330 (N_30330,N_29884,N_29823);
and U30331 (N_30331,N_29801,N_29151);
and U30332 (N_30332,N_29173,N_29886);
nand U30333 (N_30333,N_29330,N_29339);
and U30334 (N_30334,N_29244,N_29025);
and U30335 (N_30335,N_29634,N_29162);
nand U30336 (N_30336,N_29685,N_29104);
or U30337 (N_30337,N_29890,N_29992);
nand U30338 (N_30338,N_29287,N_29635);
nand U30339 (N_30339,N_29062,N_29591);
and U30340 (N_30340,N_29874,N_29355);
xor U30341 (N_30341,N_29599,N_29803);
nand U30342 (N_30342,N_29122,N_29447);
xnor U30343 (N_30343,N_29504,N_29709);
xnor U30344 (N_30344,N_29011,N_29295);
xnor U30345 (N_30345,N_29754,N_29506);
and U30346 (N_30346,N_29785,N_29811);
nand U30347 (N_30347,N_29051,N_29955);
xnor U30348 (N_30348,N_29835,N_29816);
and U30349 (N_30349,N_29204,N_29131);
xnor U30350 (N_30350,N_29587,N_29358);
and U30351 (N_30351,N_29750,N_29966);
and U30352 (N_30352,N_29454,N_29341);
nor U30353 (N_30353,N_29722,N_29697);
nand U30354 (N_30354,N_29095,N_29831);
or U30355 (N_30355,N_29415,N_29052);
and U30356 (N_30356,N_29619,N_29545);
xor U30357 (N_30357,N_29475,N_29812);
or U30358 (N_30358,N_29766,N_29909);
nor U30359 (N_30359,N_29996,N_29197);
xnor U30360 (N_30360,N_29492,N_29696);
nor U30361 (N_30361,N_29661,N_29216);
and U30362 (N_30362,N_29898,N_29565);
nor U30363 (N_30363,N_29997,N_29224);
and U30364 (N_30364,N_29688,N_29917);
and U30365 (N_30365,N_29102,N_29961);
nor U30366 (N_30366,N_29684,N_29208);
nand U30367 (N_30367,N_29164,N_29681);
nand U30368 (N_30368,N_29618,N_29496);
nand U30369 (N_30369,N_29005,N_29281);
xor U30370 (N_30370,N_29980,N_29817);
nand U30371 (N_30371,N_29146,N_29663);
and U30372 (N_30372,N_29865,N_29879);
nor U30373 (N_30373,N_29559,N_29206);
xor U30374 (N_30374,N_29236,N_29009);
and U30375 (N_30375,N_29719,N_29608);
nor U30376 (N_30376,N_29042,N_29464);
xor U30377 (N_30377,N_29135,N_29318);
nor U30378 (N_30378,N_29023,N_29672);
or U30379 (N_30379,N_29792,N_29867);
nand U30380 (N_30380,N_29180,N_29439);
and U30381 (N_30381,N_29342,N_29302);
xnor U30382 (N_30382,N_29662,N_29136);
nand U30383 (N_30383,N_29648,N_29316);
nor U30384 (N_30384,N_29083,N_29664);
and U30385 (N_30385,N_29087,N_29322);
or U30386 (N_30386,N_29620,N_29314);
and U30387 (N_30387,N_29384,N_29675);
xor U30388 (N_30388,N_29170,N_29484);
xnor U30389 (N_30389,N_29366,N_29745);
and U30390 (N_30390,N_29705,N_29387);
xnor U30391 (N_30391,N_29692,N_29936);
and U30392 (N_30392,N_29360,N_29160);
nor U30393 (N_30393,N_29082,N_29680);
or U30394 (N_30394,N_29329,N_29952);
xnor U30395 (N_30395,N_29825,N_29721);
and U30396 (N_30396,N_29337,N_29066);
xnor U30397 (N_30397,N_29734,N_29683);
or U30398 (N_30398,N_29485,N_29002);
nor U30399 (N_30399,N_29272,N_29739);
or U30400 (N_30400,N_29259,N_29117);
nor U30401 (N_30401,N_29309,N_29289);
nor U30402 (N_30402,N_29761,N_29912);
and U30403 (N_30403,N_29073,N_29808);
or U30404 (N_30404,N_29317,N_29939);
nand U30405 (N_30405,N_29918,N_29522);
and U30406 (N_30406,N_29836,N_29598);
nand U30407 (N_30407,N_29382,N_29658);
and U30408 (N_30408,N_29392,N_29718);
nand U30409 (N_30409,N_29922,N_29773);
xor U30410 (N_30410,N_29906,N_29081);
xor U30411 (N_30411,N_29945,N_29037);
nand U30412 (N_30412,N_29093,N_29407);
nand U30413 (N_30413,N_29199,N_29951);
xnor U30414 (N_30414,N_29285,N_29682);
nand U30415 (N_30415,N_29265,N_29139);
nand U30416 (N_30416,N_29508,N_29280);
xnor U30417 (N_30417,N_29090,N_29478);
or U30418 (N_30418,N_29964,N_29039);
or U30419 (N_30419,N_29784,N_29455);
or U30420 (N_30420,N_29731,N_29779);
xor U30421 (N_30421,N_29022,N_29854);
nand U30422 (N_30422,N_29291,N_29790);
or U30423 (N_30423,N_29797,N_29026);
nor U30424 (N_30424,N_29687,N_29315);
nand U30425 (N_30425,N_29813,N_29553);
nor U30426 (N_30426,N_29364,N_29263);
nor U30427 (N_30427,N_29133,N_29205);
nand U30428 (N_30428,N_29427,N_29972);
or U30429 (N_30429,N_29010,N_29549);
xor U30430 (N_30430,N_29124,N_29641);
xor U30431 (N_30431,N_29899,N_29016);
and U30432 (N_30432,N_29841,N_29060);
nor U30433 (N_30433,N_29466,N_29313);
nand U30434 (N_30434,N_29450,N_29157);
xnor U30435 (N_30435,N_29891,N_29189);
nor U30436 (N_30436,N_29256,N_29892);
xor U30437 (N_30437,N_29373,N_29128);
and U30438 (N_30438,N_29410,N_29720);
or U30439 (N_30439,N_29789,N_29701);
nor U30440 (N_30440,N_29777,N_29732);
nand U30441 (N_30441,N_29449,N_29760);
nor U30442 (N_30442,N_29954,N_29398);
nand U30443 (N_30443,N_29181,N_29059);
and U30444 (N_30444,N_29534,N_29293);
xor U30445 (N_30445,N_29099,N_29423);
and U30446 (N_30446,N_29515,N_29840);
nor U30447 (N_30447,N_29793,N_29498);
or U30448 (N_30448,N_29896,N_29584);
nand U30449 (N_30449,N_29775,N_29596);
and U30450 (N_30450,N_29030,N_29417);
xor U30451 (N_30451,N_29702,N_29356);
nand U30452 (N_30452,N_29388,N_29805);
or U30453 (N_30453,N_29780,N_29535);
xnor U30454 (N_30454,N_29677,N_29986);
or U30455 (N_30455,N_29226,N_29957);
or U30456 (N_30456,N_29539,N_29772);
and U30457 (N_30457,N_29617,N_29100);
nor U30458 (N_30458,N_29523,N_29776);
nor U30459 (N_30459,N_29849,N_29286);
nand U30460 (N_30460,N_29307,N_29699);
nor U30461 (N_30461,N_29931,N_29238);
or U30462 (N_30462,N_29561,N_29578);
and U30463 (N_30463,N_29348,N_29000);
nor U30464 (N_30464,N_29261,N_29723);
xor U30465 (N_30465,N_29020,N_29035);
xnor U30466 (N_30466,N_29147,N_29424);
nand U30467 (N_30467,N_29679,N_29588);
nor U30468 (N_30468,N_29074,N_29991);
nor U30469 (N_30469,N_29689,N_29837);
nor U30470 (N_30470,N_29556,N_29375);
or U30471 (N_30471,N_29248,N_29213);
or U30472 (N_30472,N_29027,N_29795);
and U30473 (N_30473,N_29928,N_29121);
or U30474 (N_30474,N_29581,N_29864);
or U30475 (N_30475,N_29769,N_29190);
nand U30476 (N_30476,N_29386,N_29114);
nand U30477 (N_30477,N_29524,N_29551);
or U30478 (N_30478,N_29623,N_29376);
or U30479 (N_30479,N_29946,N_29740);
nand U30480 (N_30480,N_29655,N_29920);
nand U30481 (N_30481,N_29380,N_29125);
xnor U30482 (N_30482,N_29894,N_29642);
nand U30483 (N_30483,N_29969,N_29861);
nor U30484 (N_30484,N_29554,N_29420);
nor U30485 (N_30485,N_29707,N_29031);
or U30486 (N_30486,N_29602,N_29044);
or U30487 (N_30487,N_29431,N_29774);
nand U30488 (N_30488,N_29763,N_29821);
xor U30489 (N_30489,N_29644,N_29870);
nor U30490 (N_30490,N_29477,N_29908);
nand U30491 (N_30491,N_29603,N_29903);
and U30492 (N_30492,N_29353,N_29056);
nor U30493 (N_30493,N_29575,N_29067);
xnor U30494 (N_30494,N_29571,N_29168);
nor U30495 (N_30495,N_29345,N_29041);
or U30496 (N_30496,N_29822,N_29768);
and U30497 (N_30497,N_29666,N_29430);
and U30498 (N_30498,N_29349,N_29425);
nand U30499 (N_30499,N_29241,N_29968);
nor U30500 (N_30500,N_29509,N_29566);
or U30501 (N_30501,N_29082,N_29583);
xor U30502 (N_30502,N_29995,N_29965);
xor U30503 (N_30503,N_29218,N_29508);
and U30504 (N_30504,N_29036,N_29455);
or U30505 (N_30505,N_29017,N_29789);
nand U30506 (N_30506,N_29831,N_29247);
or U30507 (N_30507,N_29013,N_29141);
and U30508 (N_30508,N_29550,N_29768);
xor U30509 (N_30509,N_29497,N_29507);
and U30510 (N_30510,N_29371,N_29879);
nand U30511 (N_30511,N_29438,N_29561);
and U30512 (N_30512,N_29678,N_29442);
and U30513 (N_30513,N_29746,N_29186);
nand U30514 (N_30514,N_29174,N_29571);
or U30515 (N_30515,N_29681,N_29231);
nand U30516 (N_30516,N_29253,N_29022);
or U30517 (N_30517,N_29141,N_29658);
xnor U30518 (N_30518,N_29280,N_29905);
nand U30519 (N_30519,N_29486,N_29038);
nand U30520 (N_30520,N_29007,N_29023);
or U30521 (N_30521,N_29746,N_29146);
or U30522 (N_30522,N_29551,N_29897);
xor U30523 (N_30523,N_29841,N_29286);
or U30524 (N_30524,N_29893,N_29990);
nor U30525 (N_30525,N_29266,N_29524);
and U30526 (N_30526,N_29888,N_29362);
nor U30527 (N_30527,N_29633,N_29812);
nand U30528 (N_30528,N_29000,N_29848);
and U30529 (N_30529,N_29931,N_29462);
or U30530 (N_30530,N_29425,N_29904);
nor U30531 (N_30531,N_29262,N_29457);
xor U30532 (N_30532,N_29926,N_29146);
and U30533 (N_30533,N_29587,N_29406);
and U30534 (N_30534,N_29892,N_29043);
nand U30535 (N_30535,N_29392,N_29235);
nand U30536 (N_30536,N_29566,N_29883);
and U30537 (N_30537,N_29645,N_29107);
and U30538 (N_30538,N_29726,N_29239);
nand U30539 (N_30539,N_29348,N_29159);
or U30540 (N_30540,N_29162,N_29429);
xor U30541 (N_30541,N_29420,N_29377);
or U30542 (N_30542,N_29370,N_29081);
and U30543 (N_30543,N_29082,N_29312);
and U30544 (N_30544,N_29507,N_29380);
nor U30545 (N_30545,N_29521,N_29199);
nor U30546 (N_30546,N_29030,N_29412);
or U30547 (N_30547,N_29011,N_29230);
nor U30548 (N_30548,N_29078,N_29781);
or U30549 (N_30549,N_29520,N_29580);
nand U30550 (N_30550,N_29632,N_29109);
xnor U30551 (N_30551,N_29903,N_29745);
nor U30552 (N_30552,N_29937,N_29514);
or U30553 (N_30553,N_29188,N_29038);
xor U30554 (N_30554,N_29632,N_29352);
nor U30555 (N_30555,N_29017,N_29799);
nor U30556 (N_30556,N_29643,N_29469);
or U30557 (N_30557,N_29514,N_29638);
nand U30558 (N_30558,N_29557,N_29757);
and U30559 (N_30559,N_29831,N_29893);
nand U30560 (N_30560,N_29781,N_29324);
nor U30561 (N_30561,N_29417,N_29011);
xor U30562 (N_30562,N_29644,N_29265);
nor U30563 (N_30563,N_29585,N_29836);
nand U30564 (N_30564,N_29828,N_29960);
and U30565 (N_30565,N_29099,N_29044);
xnor U30566 (N_30566,N_29704,N_29695);
nor U30567 (N_30567,N_29610,N_29719);
nor U30568 (N_30568,N_29234,N_29922);
nand U30569 (N_30569,N_29547,N_29579);
and U30570 (N_30570,N_29449,N_29539);
xnor U30571 (N_30571,N_29213,N_29839);
and U30572 (N_30572,N_29004,N_29687);
xnor U30573 (N_30573,N_29964,N_29320);
xnor U30574 (N_30574,N_29679,N_29806);
or U30575 (N_30575,N_29526,N_29249);
and U30576 (N_30576,N_29345,N_29607);
nand U30577 (N_30577,N_29253,N_29799);
nor U30578 (N_30578,N_29704,N_29886);
nand U30579 (N_30579,N_29682,N_29134);
nand U30580 (N_30580,N_29087,N_29110);
nand U30581 (N_30581,N_29002,N_29491);
nor U30582 (N_30582,N_29871,N_29381);
and U30583 (N_30583,N_29549,N_29050);
or U30584 (N_30584,N_29850,N_29554);
nor U30585 (N_30585,N_29555,N_29999);
nor U30586 (N_30586,N_29139,N_29449);
xnor U30587 (N_30587,N_29220,N_29555);
or U30588 (N_30588,N_29583,N_29024);
nor U30589 (N_30589,N_29014,N_29779);
xnor U30590 (N_30590,N_29456,N_29151);
nor U30591 (N_30591,N_29349,N_29026);
or U30592 (N_30592,N_29100,N_29079);
nor U30593 (N_30593,N_29559,N_29133);
nor U30594 (N_30594,N_29944,N_29563);
xor U30595 (N_30595,N_29454,N_29096);
and U30596 (N_30596,N_29756,N_29237);
nand U30597 (N_30597,N_29385,N_29755);
xor U30598 (N_30598,N_29907,N_29945);
nand U30599 (N_30599,N_29374,N_29470);
nor U30600 (N_30600,N_29232,N_29437);
xnor U30601 (N_30601,N_29359,N_29041);
xnor U30602 (N_30602,N_29089,N_29430);
nand U30603 (N_30603,N_29331,N_29728);
nand U30604 (N_30604,N_29301,N_29022);
xnor U30605 (N_30605,N_29594,N_29917);
nand U30606 (N_30606,N_29974,N_29517);
and U30607 (N_30607,N_29658,N_29939);
xor U30608 (N_30608,N_29339,N_29214);
nand U30609 (N_30609,N_29187,N_29703);
and U30610 (N_30610,N_29614,N_29946);
nand U30611 (N_30611,N_29966,N_29544);
xnor U30612 (N_30612,N_29741,N_29859);
or U30613 (N_30613,N_29723,N_29373);
nand U30614 (N_30614,N_29875,N_29491);
and U30615 (N_30615,N_29379,N_29836);
nand U30616 (N_30616,N_29333,N_29585);
and U30617 (N_30617,N_29814,N_29098);
or U30618 (N_30618,N_29263,N_29874);
nor U30619 (N_30619,N_29950,N_29818);
and U30620 (N_30620,N_29188,N_29091);
nor U30621 (N_30621,N_29156,N_29908);
or U30622 (N_30622,N_29848,N_29020);
and U30623 (N_30623,N_29274,N_29785);
xnor U30624 (N_30624,N_29334,N_29550);
and U30625 (N_30625,N_29854,N_29859);
or U30626 (N_30626,N_29890,N_29510);
or U30627 (N_30627,N_29261,N_29628);
xor U30628 (N_30628,N_29872,N_29343);
xnor U30629 (N_30629,N_29215,N_29743);
nor U30630 (N_30630,N_29523,N_29188);
nand U30631 (N_30631,N_29966,N_29014);
nor U30632 (N_30632,N_29018,N_29577);
or U30633 (N_30633,N_29034,N_29418);
nor U30634 (N_30634,N_29264,N_29336);
and U30635 (N_30635,N_29570,N_29148);
or U30636 (N_30636,N_29820,N_29076);
nor U30637 (N_30637,N_29669,N_29200);
nand U30638 (N_30638,N_29356,N_29134);
xnor U30639 (N_30639,N_29493,N_29629);
xor U30640 (N_30640,N_29579,N_29174);
nor U30641 (N_30641,N_29832,N_29848);
nor U30642 (N_30642,N_29993,N_29400);
and U30643 (N_30643,N_29791,N_29960);
nor U30644 (N_30644,N_29983,N_29592);
nor U30645 (N_30645,N_29553,N_29593);
and U30646 (N_30646,N_29951,N_29870);
or U30647 (N_30647,N_29938,N_29312);
or U30648 (N_30648,N_29131,N_29401);
or U30649 (N_30649,N_29388,N_29970);
xnor U30650 (N_30650,N_29853,N_29500);
nand U30651 (N_30651,N_29430,N_29051);
xor U30652 (N_30652,N_29718,N_29457);
or U30653 (N_30653,N_29407,N_29346);
nand U30654 (N_30654,N_29277,N_29996);
or U30655 (N_30655,N_29279,N_29028);
nor U30656 (N_30656,N_29222,N_29749);
nand U30657 (N_30657,N_29191,N_29729);
xnor U30658 (N_30658,N_29785,N_29161);
and U30659 (N_30659,N_29049,N_29952);
xnor U30660 (N_30660,N_29388,N_29229);
and U30661 (N_30661,N_29422,N_29223);
nor U30662 (N_30662,N_29885,N_29307);
nand U30663 (N_30663,N_29054,N_29705);
nand U30664 (N_30664,N_29428,N_29518);
nand U30665 (N_30665,N_29409,N_29071);
nor U30666 (N_30666,N_29167,N_29408);
nor U30667 (N_30667,N_29061,N_29409);
or U30668 (N_30668,N_29363,N_29369);
xor U30669 (N_30669,N_29439,N_29323);
nor U30670 (N_30670,N_29763,N_29150);
and U30671 (N_30671,N_29384,N_29895);
or U30672 (N_30672,N_29233,N_29248);
nand U30673 (N_30673,N_29674,N_29905);
or U30674 (N_30674,N_29870,N_29040);
or U30675 (N_30675,N_29017,N_29645);
and U30676 (N_30676,N_29689,N_29082);
nor U30677 (N_30677,N_29104,N_29263);
and U30678 (N_30678,N_29737,N_29615);
nand U30679 (N_30679,N_29817,N_29186);
xor U30680 (N_30680,N_29901,N_29239);
and U30681 (N_30681,N_29253,N_29362);
nand U30682 (N_30682,N_29372,N_29685);
or U30683 (N_30683,N_29814,N_29712);
nor U30684 (N_30684,N_29165,N_29550);
xnor U30685 (N_30685,N_29147,N_29558);
nor U30686 (N_30686,N_29958,N_29148);
nand U30687 (N_30687,N_29419,N_29194);
nor U30688 (N_30688,N_29977,N_29001);
and U30689 (N_30689,N_29686,N_29462);
xnor U30690 (N_30690,N_29783,N_29638);
nand U30691 (N_30691,N_29226,N_29815);
nor U30692 (N_30692,N_29495,N_29800);
xor U30693 (N_30693,N_29261,N_29031);
nor U30694 (N_30694,N_29298,N_29829);
xor U30695 (N_30695,N_29076,N_29492);
xor U30696 (N_30696,N_29747,N_29938);
and U30697 (N_30697,N_29771,N_29246);
and U30698 (N_30698,N_29199,N_29242);
xor U30699 (N_30699,N_29614,N_29950);
or U30700 (N_30700,N_29362,N_29333);
nand U30701 (N_30701,N_29220,N_29926);
nor U30702 (N_30702,N_29822,N_29871);
nand U30703 (N_30703,N_29312,N_29687);
xor U30704 (N_30704,N_29666,N_29691);
and U30705 (N_30705,N_29674,N_29342);
and U30706 (N_30706,N_29321,N_29931);
nand U30707 (N_30707,N_29510,N_29123);
xor U30708 (N_30708,N_29885,N_29402);
xor U30709 (N_30709,N_29269,N_29228);
and U30710 (N_30710,N_29396,N_29720);
nand U30711 (N_30711,N_29562,N_29391);
xnor U30712 (N_30712,N_29278,N_29755);
and U30713 (N_30713,N_29392,N_29520);
and U30714 (N_30714,N_29027,N_29385);
xnor U30715 (N_30715,N_29894,N_29694);
xnor U30716 (N_30716,N_29666,N_29535);
nor U30717 (N_30717,N_29250,N_29217);
or U30718 (N_30718,N_29907,N_29666);
and U30719 (N_30719,N_29190,N_29588);
nor U30720 (N_30720,N_29204,N_29289);
nand U30721 (N_30721,N_29943,N_29648);
nand U30722 (N_30722,N_29181,N_29211);
nor U30723 (N_30723,N_29163,N_29461);
or U30724 (N_30724,N_29102,N_29037);
nor U30725 (N_30725,N_29295,N_29456);
or U30726 (N_30726,N_29479,N_29108);
or U30727 (N_30727,N_29694,N_29255);
and U30728 (N_30728,N_29838,N_29611);
and U30729 (N_30729,N_29105,N_29437);
and U30730 (N_30730,N_29930,N_29761);
or U30731 (N_30731,N_29475,N_29695);
or U30732 (N_30732,N_29490,N_29084);
nand U30733 (N_30733,N_29907,N_29583);
and U30734 (N_30734,N_29930,N_29350);
xor U30735 (N_30735,N_29828,N_29202);
nand U30736 (N_30736,N_29857,N_29672);
and U30737 (N_30737,N_29566,N_29167);
nor U30738 (N_30738,N_29833,N_29713);
xor U30739 (N_30739,N_29934,N_29024);
and U30740 (N_30740,N_29963,N_29175);
nand U30741 (N_30741,N_29238,N_29557);
nor U30742 (N_30742,N_29941,N_29719);
or U30743 (N_30743,N_29426,N_29575);
xnor U30744 (N_30744,N_29653,N_29791);
and U30745 (N_30745,N_29185,N_29735);
nor U30746 (N_30746,N_29904,N_29955);
nand U30747 (N_30747,N_29885,N_29445);
nand U30748 (N_30748,N_29021,N_29832);
nor U30749 (N_30749,N_29425,N_29897);
and U30750 (N_30750,N_29368,N_29777);
nor U30751 (N_30751,N_29280,N_29564);
nand U30752 (N_30752,N_29191,N_29263);
or U30753 (N_30753,N_29205,N_29157);
or U30754 (N_30754,N_29305,N_29140);
nand U30755 (N_30755,N_29575,N_29648);
nand U30756 (N_30756,N_29028,N_29340);
nand U30757 (N_30757,N_29182,N_29087);
xnor U30758 (N_30758,N_29337,N_29116);
nor U30759 (N_30759,N_29604,N_29306);
nand U30760 (N_30760,N_29447,N_29003);
nand U30761 (N_30761,N_29266,N_29010);
xnor U30762 (N_30762,N_29753,N_29784);
and U30763 (N_30763,N_29344,N_29178);
xor U30764 (N_30764,N_29416,N_29079);
or U30765 (N_30765,N_29730,N_29606);
nand U30766 (N_30766,N_29433,N_29654);
or U30767 (N_30767,N_29844,N_29675);
or U30768 (N_30768,N_29150,N_29515);
or U30769 (N_30769,N_29854,N_29379);
nand U30770 (N_30770,N_29027,N_29109);
nor U30771 (N_30771,N_29581,N_29748);
nor U30772 (N_30772,N_29429,N_29827);
nor U30773 (N_30773,N_29818,N_29033);
nor U30774 (N_30774,N_29079,N_29058);
nor U30775 (N_30775,N_29806,N_29556);
nand U30776 (N_30776,N_29694,N_29860);
and U30777 (N_30777,N_29311,N_29737);
nand U30778 (N_30778,N_29411,N_29955);
or U30779 (N_30779,N_29956,N_29848);
nor U30780 (N_30780,N_29119,N_29372);
xnor U30781 (N_30781,N_29506,N_29264);
nor U30782 (N_30782,N_29121,N_29259);
xnor U30783 (N_30783,N_29283,N_29722);
nor U30784 (N_30784,N_29901,N_29708);
xnor U30785 (N_30785,N_29978,N_29783);
and U30786 (N_30786,N_29304,N_29400);
nor U30787 (N_30787,N_29687,N_29591);
or U30788 (N_30788,N_29985,N_29561);
or U30789 (N_30789,N_29068,N_29408);
or U30790 (N_30790,N_29103,N_29424);
xnor U30791 (N_30791,N_29897,N_29133);
or U30792 (N_30792,N_29862,N_29186);
nand U30793 (N_30793,N_29892,N_29625);
nor U30794 (N_30794,N_29241,N_29001);
and U30795 (N_30795,N_29509,N_29959);
or U30796 (N_30796,N_29016,N_29371);
or U30797 (N_30797,N_29384,N_29974);
xor U30798 (N_30798,N_29826,N_29474);
nand U30799 (N_30799,N_29929,N_29308);
and U30800 (N_30800,N_29102,N_29832);
nand U30801 (N_30801,N_29592,N_29847);
nand U30802 (N_30802,N_29910,N_29558);
nand U30803 (N_30803,N_29285,N_29157);
xnor U30804 (N_30804,N_29024,N_29051);
xnor U30805 (N_30805,N_29303,N_29942);
nor U30806 (N_30806,N_29108,N_29421);
xor U30807 (N_30807,N_29733,N_29626);
xnor U30808 (N_30808,N_29686,N_29908);
and U30809 (N_30809,N_29434,N_29870);
xor U30810 (N_30810,N_29042,N_29374);
or U30811 (N_30811,N_29953,N_29288);
and U30812 (N_30812,N_29886,N_29319);
nor U30813 (N_30813,N_29650,N_29596);
or U30814 (N_30814,N_29324,N_29944);
xor U30815 (N_30815,N_29509,N_29320);
nand U30816 (N_30816,N_29776,N_29712);
or U30817 (N_30817,N_29225,N_29435);
xnor U30818 (N_30818,N_29911,N_29916);
nand U30819 (N_30819,N_29960,N_29304);
and U30820 (N_30820,N_29051,N_29976);
nor U30821 (N_30821,N_29290,N_29066);
nor U30822 (N_30822,N_29488,N_29430);
or U30823 (N_30823,N_29644,N_29628);
and U30824 (N_30824,N_29095,N_29535);
and U30825 (N_30825,N_29153,N_29077);
nand U30826 (N_30826,N_29193,N_29864);
and U30827 (N_30827,N_29374,N_29398);
or U30828 (N_30828,N_29555,N_29363);
and U30829 (N_30829,N_29181,N_29804);
or U30830 (N_30830,N_29271,N_29499);
nand U30831 (N_30831,N_29169,N_29413);
xnor U30832 (N_30832,N_29490,N_29463);
nor U30833 (N_30833,N_29435,N_29757);
xnor U30834 (N_30834,N_29933,N_29288);
and U30835 (N_30835,N_29278,N_29840);
nor U30836 (N_30836,N_29907,N_29927);
xor U30837 (N_30837,N_29735,N_29047);
and U30838 (N_30838,N_29739,N_29449);
and U30839 (N_30839,N_29781,N_29140);
nor U30840 (N_30840,N_29658,N_29380);
nand U30841 (N_30841,N_29875,N_29013);
or U30842 (N_30842,N_29174,N_29822);
nor U30843 (N_30843,N_29644,N_29684);
nand U30844 (N_30844,N_29518,N_29646);
xnor U30845 (N_30845,N_29891,N_29210);
nor U30846 (N_30846,N_29898,N_29852);
nand U30847 (N_30847,N_29798,N_29714);
nor U30848 (N_30848,N_29420,N_29668);
or U30849 (N_30849,N_29398,N_29470);
nand U30850 (N_30850,N_29283,N_29494);
nand U30851 (N_30851,N_29988,N_29062);
or U30852 (N_30852,N_29587,N_29083);
nand U30853 (N_30853,N_29983,N_29197);
nand U30854 (N_30854,N_29291,N_29523);
and U30855 (N_30855,N_29171,N_29314);
xnor U30856 (N_30856,N_29298,N_29716);
nor U30857 (N_30857,N_29448,N_29273);
and U30858 (N_30858,N_29761,N_29181);
or U30859 (N_30859,N_29976,N_29031);
or U30860 (N_30860,N_29260,N_29753);
nor U30861 (N_30861,N_29503,N_29292);
nand U30862 (N_30862,N_29352,N_29658);
or U30863 (N_30863,N_29530,N_29857);
and U30864 (N_30864,N_29477,N_29798);
nor U30865 (N_30865,N_29278,N_29216);
nand U30866 (N_30866,N_29528,N_29288);
or U30867 (N_30867,N_29587,N_29656);
nor U30868 (N_30868,N_29654,N_29171);
xor U30869 (N_30869,N_29891,N_29465);
and U30870 (N_30870,N_29276,N_29431);
xnor U30871 (N_30871,N_29139,N_29613);
xor U30872 (N_30872,N_29487,N_29898);
nor U30873 (N_30873,N_29714,N_29066);
and U30874 (N_30874,N_29264,N_29598);
and U30875 (N_30875,N_29930,N_29369);
nor U30876 (N_30876,N_29924,N_29315);
xnor U30877 (N_30877,N_29925,N_29436);
nand U30878 (N_30878,N_29495,N_29125);
or U30879 (N_30879,N_29525,N_29594);
xor U30880 (N_30880,N_29351,N_29568);
xnor U30881 (N_30881,N_29681,N_29436);
nor U30882 (N_30882,N_29828,N_29000);
xnor U30883 (N_30883,N_29274,N_29203);
xor U30884 (N_30884,N_29034,N_29892);
nand U30885 (N_30885,N_29173,N_29677);
xnor U30886 (N_30886,N_29383,N_29384);
or U30887 (N_30887,N_29867,N_29755);
xor U30888 (N_30888,N_29207,N_29517);
or U30889 (N_30889,N_29997,N_29090);
and U30890 (N_30890,N_29925,N_29359);
xnor U30891 (N_30891,N_29668,N_29649);
nand U30892 (N_30892,N_29921,N_29162);
or U30893 (N_30893,N_29120,N_29553);
xor U30894 (N_30894,N_29673,N_29229);
nor U30895 (N_30895,N_29049,N_29829);
nor U30896 (N_30896,N_29265,N_29336);
or U30897 (N_30897,N_29122,N_29090);
nand U30898 (N_30898,N_29696,N_29895);
and U30899 (N_30899,N_29139,N_29587);
xor U30900 (N_30900,N_29403,N_29649);
xor U30901 (N_30901,N_29040,N_29021);
nor U30902 (N_30902,N_29825,N_29204);
or U30903 (N_30903,N_29079,N_29856);
nor U30904 (N_30904,N_29446,N_29680);
nor U30905 (N_30905,N_29934,N_29762);
and U30906 (N_30906,N_29372,N_29055);
and U30907 (N_30907,N_29921,N_29246);
nand U30908 (N_30908,N_29374,N_29325);
nand U30909 (N_30909,N_29254,N_29258);
nand U30910 (N_30910,N_29859,N_29739);
or U30911 (N_30911,N_29331,N_29327);
and U30912 (N_30912,N_29217,N_29220);
nor U30913 (N_30913,N_29234,N_29792);
nor U30914 (N_30914,N_29366,N_29309);
nand U30915 (N_30915,N_29042,N_29393);
or U30916 (N_30916,N_29310,N_29127);
and U30917 (N_30917,N_29390,N_29272);
or U30918 (N_30918,N_29167,N_29411);
and U30919 (N_30919,N_29649,N_29719);
and U30920 (N_30920,N_29850,N_29375);
or U30921 (N_30921,N_29026,N_29703);
or U30922 (N_30922,N_29612,N_29847);
nor U30923 (N_30923,N_29209,N_29063);
nand U30924 (N_30924,N_29220,N_29290);
and U30925 (N_30925,N_29106,N_29256);
or U30926 (N_30926,N_29021,N_29253);
nor U30927 (N_30927,N_29417,N_29115);
nand U30928 (N_30928,N_29645,N_29474);
nor U30929 (N_30929,N_29233,N_29486);
nor U30930 (N_30930,N_29829,N_29343);
nand U30931 (N_30931,N_29274,N_29805);
nor U30932 (N_30932,N_29781,N_29828);
or U30933 (N_30933,N_29661,N_29619);
xor U30934 (N_30934,N_29541,N_29375);
and U30935 (N_30935,N_29074,N_29207);
nor U30936 (N_30936,N_29529,N_29836);
nor U30937 (N_30937,N_29888,N_29026);
xor U30938 (N_30938,N_29248,N_29856);
or U30939 (N_30939,N_29151,N_29049);
nand U30940 (N_30940,N_29516,N_29275);
or U30941 (N_30941,N_29967,N_29081);
nor U30942 (N_30942,N_29813,N_29855);
or U30943 (N_30943,N_29442,N_29279);
and U30944 (N_30944,N_29712,N_29479);
or U30945 (N_30945,N_29967,N_29148);
or U30946 (N_30946,N_29810,N_29185);
and U30947 (N_30947,N_29429,N_29928);
nor U30948 (N_30948,N_29812,N_29058);
nand U30949 (N_30949,N_29128,N_29481);
or U30950 (N_30950,N_29524,N_29366);
or U30951 (N_30951,N_29006,N_29806);
xnor U30952 (N_30952,N_29023,N_29674);
xnor U30953 (N_30953,N_29235,N_29122);
and U30954 (N_30954,N_29706,N_29799);
or U30955 (N_30955,N_29721,N_29085);
or U30956 (N_30956,N_29879,N_29029);
nand U30957 (N_30957,N_29922,N_29501);
nand U30958 (N_30958,N_29361,N_29492);
or U30959 (N_30959,N_29332,N_29002);
and U30960 (N_30960,N_29851,N_29540);
and U30961 (N_30961,N_29915,N_29895);
and U30962 (N_30962,N_29386,N_29420);
and U30963 (N_30963,N_29969,N_29255);
xor U30964 (N_30964,N_29669,N_29538);
nor U30965 (N_30965,N_29456,N_29730);
and U30966 (N_30966,N_29593,N_29273);
nor U30967 (N_30967,N_29471,N_29119);
and U30968 (N_30968,N_29385,N_29435);
xor U30969 (N_30969,N_29891,N_29640);
or U30970 (N_30970,N_29946,N_29848);
nand U30971 (N_30971,N_29621,N_29014);
xnor U30972 (N_30972,N_29076,N_29588);
and U30973 (N_30973,N_29644,N_29776);
xnor U30974 (N_30974,N_29371,N_29606);
nor U30975 (N_30975,N_29352,N_29202);
or U30976 (N_30976,N_29859,N_29974);
and U30977 (N_30977,N_29579,N_29066);
or U30978 (N_30978,N_29106,N_29742);
xor U30979 (N_30979,N_29437,N_29539);
or U30980 (N_30980,N_29075,N_29903);
xor U30981 (N_30981,N_29044,N_29364);
nor U30982 (N_30982,N_29233,N_29159);
and U30983 (N_30983,N_29333,N_29975);
nor U30984 (N_30984,N_29690,N_29895);
nor U30985 (N_30985,N_29831,N_29732);
xnor U30986 (N_30986,N_29269,N_29917);
and U30987 (N_30987,N_29007,N_29627);
xnor U30988 (N_30988,N_29644,N_29865);
nor U30989 (N_30989,N_29681,N_29213);
xor U30990 (N_30990,N_29850,N_29773);
xnor U30991 (N_30991,N_29850,N_29011);
xor U30992 (N_30992,N_29647,N_29979);
or U30993 (N_30993,N_29372,N_29258);
or U30994 (N_30994,N_29195,N_29443);
nor U30995 (N_30995,N_29722,N_29833);
nor U30996 (N_30996,N_29157,N_29427);
nand U30997 (N_30997,N_29594,N_29996);
nor U30998 (N_30998,N_29002,N_29401);
xnor U30999 (N_30999,N_29198,N_29661);
xor U31000 (N_31000,N_30538,N_30399);
nand U31001 (N_31001,N_30986,N_30710);
nor U31002 (N_31002,N_30900,N_30184);
nand U31003 (N_31003,N_30932,N_30702);
or U31004 (N_31004,N_30099,N_30653);
xnor U31005 (N_31005,N_30031,N_30460);
nand U31006 (N_31006,N_30470,N_30020);
nand U31007 (N_31007,N_30004,N_30782);
xor U31008 (N_31008,N_30283,N_30927);
xor U31009 (N_31009,N_30976,N_30656);
or U31010 (N_31010,N_30618,N_30621);
nor U31011 (N_31011,N_30585,N_30831);
and U31012 (N_31012,N_30473,N_30925);
nor U31013 (N_31013,N_30069,N_30661);
xnor U31014 (N_31014,N_30134,N_30689);
xnor U31015 (N_31015,N_30378,N_30504);
and U31016 (N_31016,N_30561,N_30809);
and U31017 (N_31017,N_30597,N_30302);
and U31018 (N_31018,N_30784,N_30558);
nor U31019 (N_31019,N_30033,N_30388);
nor U31020 (N_31020,N_30598,N_30658);
and U31021 (N_31021,N_30731,N_30848);
nor U31022 (N_31022,N_30748,N_30619);
or U31023 (N_31023,N_30596,N_30912);
nand U31024 (N_31024,N_30592,N_30531);
xor U31025 (N_31025,N_30352,N_30959);
nand U31026 (N_31026,N_30040,N_30508);
or U31027 (N_31027,N_30447,N_30157);
or U31028 (N_31028,N_30001,N_30591);
nor U31029 (N_31029,N_30210,N_30933);
xnor U31030 (N_31030,N_30572,N_30586);
nand U31031 (N_31031,N_30016,N_30027);
nor U31032 (N_31032,N_30814,N_30244);
nand U31033 (N_31033,N_30650,N_30622);
xor U31034 (N_31034,N_30002,N_30061);
or U31035 (N_31035,N_30593,N_30499);
nand U31036 (N_31036,N_30118,N_30454);
and U31037 (N_31037,N_30633,N_30091);
xnor U31038 (N_31038,N_30541,N_30347);
and U31039 (N_31039,N_30300,N_30173);
and U31040 (N_31040,N_30233,N_30349);
xnor U31041 (N_31041,N_30837,N_30924);
nand U31042 (N_31042,N_30567,N_30296);
or U31043 (N_31043,N_30018,N_30594);
or U31044 (N_31044,N_30902,N_30429);
nand U31045 (N_31045,N_30497,N_30998);
nand U31046 (N_31046,N_30711,N_30866);
or U31047 (N_31047,N_30863,N_30030);
nand U31048 (N_31048,N_30323,N_30212);
xnor U31049 (N_31049,N_30439,N_30330);
nand U31050 (N_31050,N_30791,N_30771);
or U31051 (N_31051,N_30444,N_30076);
or U31052 (N_31052,N_30741,N_30403);
and U31053 (N_31053,N_30105,N_30843);
nand U31054 (N_31054,N_30326,N_30487);
and U31055 (N_31055,N_30333,N_30951);
nor U31056 (N_31056,N_30495,N_30742);
xnor U31057 (N_31057,N_30207,N_30097);
xnor U31058 (N_31058,N_30509,N_30582);
nor U31059 (N_31059,N_30434,N_30915);
or U31060 (N_31060,N_30433,N_30974);
xnor U31061 (N_31061,N_30073,N_30305);
nand U31062 (N_31062,N_30777,N_30894);
or U31063 (N_31063,N_30198,N_30611);
and U31064 (N_31064,N_30634,N_30461);
or U31065 (N_31065,N_30587,N_30936);
and U31066 (N_31066,N_30723,N_30035);
xor U31067 (N_31067,N_30138,N_30211);
or U31068 (N_31068,N_30026,N_30750);
nor U31069 (N_31069,N_30287,N_30778);
nor U31070 (N_31070,N_30801,N_30730);
nand U31071 (N_31071,N_30607,N_30223);
nor U31072 (N_31072,N_30215,N_30146);
or U31073 (N_31073,N_30638,N_30871);
and U31074 (N_31074,N_30518,N_30695);
xor U31075 (N_31075,N_30590,N_30328);
or U31076 (N_31076,N_30680,N_30588);
nor U31077 (N_31077,N_30535,N_30180);
xor U31078 (N_31078,N_30379,N_30017);
nor U31079 (N_31079,N_30910,N_30918);
and U31080 (N_31080,N_30732,N_30267);
xnor U31081 (N_31081,N_30816,N_30214);
nor U31082 (N_31082,N_30103,N_30421);
nor U31083 (N_31083,N_30235,N_30325);
and U31084 (N_31084,N_30032,N_30839);
xnor U31085 (N_31085,N_30054,N_30112);
or U31086 (N_31086,N_30978,N_30553);
and U31087 (N_31087,N_30288,N_30868);
xnor U31088 (N_31088,N_30892,N_30746);
and U31089 (N_31089,N_30224,N_30997);
xnor U31090 (N_31090,N_30941,N_30011);
or U31091 (N_31091,N_30056,N_30667);
nor U31092 (N_31092,N_30606,N_30392);
and U31093 (N_31093,N_30756,N_30274);
nand U31094 (N_31094,N_30983,N_30458);
xnor U31095 (N_31095,N_30089,N_30232);
xor U31096 (N_31096,N_30623,N_30317);
and U31097 (N_31097,N_30007,N_30303);
nand U31098 (N_31098,N_30948,N_30298);
and U31099 (N_31099,N_30257,N_30337);
and U31100 (N_31100,N_30525,N_30284);
and U31101 (N_31101,N_30278,N_30540);
and U31102 (N_31102,N_30336,N_30425);
nor U31103 (N_31103,N_30218,N_30861);
and U31104 (N_31104,N_30808,N_30909);
xor U31105 (N_31105,N_30763,N_30166);
and U31106 (N_31106,N_30740,N_30921);
and U31107 (N_31107,N_30744,N_30811);
nand U31108 (N_31108,N_30208,N_30152);
and U31109 (N_31109,N_30188,N_30327);
nor U31110 (N_31110,N_30869,N_30367);
nand U31111 (N_31111,N_30281,N_30136);
or U31112 (N_31112,N_30199,N_30562);
nor U31113 (N_31113,N_30943,N_30480);
xor U31114 (N_31114,N_30329,N_30041);
and U31115 (N_31115,N_30766,N_30551);
nor U31116 (N_31116,N_30654,N_30456);
nand U31117 (N_31117,N_30788,N_30301);
or U31118 (N_31118,N_30123,N_30971);
xor U31119 (N_31119,N_30269,N_30859);
nor U31120 (N_31120,N_30187,N_30050);
or U31121 (N_31121,N_30800,N_30545);
or U31122 (N_31122,N_30673,N_30872);
or U31123 (N_31123,N_30911,N_30320);
and U31124 (N_31124,N_30128,N_30645);
and U31125 (N_31125,N_30878,N_30722);
and U31126 (N_31126,N_30580,N_30898);
nor U31127 (N_31127,N_30792,N_30940);
nand U31128 (N_31128,N_30491,N_30729);
xor U31129 (N_31129,N_30039,N_30088);
xor U31130 (N_31130,N_30981,N_30227);
xnor U31131 (N_31131,N_30524,N_30749);
nor U31132 (N_31132,N_30725,N_30954);
xor U31133 (N_31133,N_30094,N_30849);
or U31134 (N_31134,N_30687,N_30490);
and U31135 (N_31135,N_30409,N_30609);
xnor U31136 (N_31136,N_30143,N_30698);
xnor U31137 (N_31137,N_30700,N_30979);
xnor U31138 (N_31138,N_30944,N_30679);
nand U31139 (N_31139,N_30957,N_30398);
nor U31140 (N_31140,N_30534,N_30290);
nor U31141 (N_31141,N_30471,N_30884);
and U31142 (N_31142,N_30360,N_30437);
nor U31143 (N_31143,N_30841,N_30907);
xnor U31144 (N_31144,N_30405,N_30441);
and U31145 (N_31145,N_30570,N_30922);
nand U31146 (N_31146,N_30221,N_30798);
or U31147 (N_31147,N_30824,N_30108);
and U31148 (N_31148,N_30579,N_30334);
nand U31149 (N_31149,N_30034,N_30289);
nor U31150 (N_31150,N_30457,N_30404);
nor U31151 (N_31151,N_30662,N_30131);
xor U31152 (N_31152,N_30282,N_30393);
xnor U31153 (N_31153,N_30029,N_30319);
nor U31154 (N_31154,N_30547,N_30202);
xnor U31155 (N_31155,N_30905,N_30158);
or U31156 (N_31156,N_30716,N_30400);
and U31157 (N_31157,N_30096,N_30028);
nand U31158 (N_31158,N_30669,N_30697);
nand U31159 (N_31159,N_30391,N_30197);
nand U31160 (N_31160,N_30293,N_30324);
nor U31161 (N_31161,N_30494,N_30557);
or U31162 (N_31162,N_30543,N_30739);
or U31163 (N_31163,N_30726,N_30307);
and U31164 (N_31164,N_30764,N_30847);
nand U31165 (N_31165,N_30394,N_30414);
xor U31166 (N_31166,N_30502,N_30620);
xnor U31167 (N_31167,N_30164,N_30203);
nor U31168 (N_31168,N_30605,N_30046);
nand U31169 (N_31169,N_30501,N_30266);
xnor U31170 (N_31170,N_30528,N_30365);
nor U31171 (N_31171,N_30485,N_30610);
xor U31172 (N_31172,N_30830,N_30265);
or U31173 (N_31173,N_30436,N_30757);
and U31174 (N_31174,N_30649,N_30375);
or U31175 (N_31175,N_30196,N_30310);
and U31176 (N_31176,N_30745,N_30366);
and U31177 (N_31177,N_30260,N_30171);
and U31178 (N_31178,N_30464,N_30044);
xnor U31179 (N_31179,N_30381,N_30646);
and U31180 (N_31180,N_30036,N_30345);
and U31181 (N_31181,N_30362,N_30364);
nor U31182 (N_31182,N_30920,N_30038);
and U31183 (N_31183,N_30111,N_30230);
nor U31184 (N_31184,N_30413,N_30760);
nor U31185 (N_31185,N_30956,N_30820);
nand U31186 (N_31186,N_30191,N_30251);
nor U31187 (N_31187,N_30758,N_30150);
xor U31188 (N_31188,N_30879,N_30126);
nand U31189 (N_31189,N_30172,N_30708);
xnor U31190 (N_31190,N_30955,N_30459);
or U31191 (N_31191,N_30870,N_30176);
nand U31192 (N_31192,N_30886,N_30442);
xor U31193 (N_31193,N_30238,N_30013);
nand U31194 (N_31194,N_30179,N_30684);
nor U31195 (N_31195,N_30245,N_30086);
nand U31196 (N_31196,N_30867,N_30468);
nor U31197 (N_31197,N_30613,N_30821);
or U31198 (N_31198,N_30942,N_30559);
and U31199 (N_31199,N_30735,N_30904);
or U31200 (N_31200,N_30930,N_30544);
nand U31201 (N_31201,N_30410,N_30259);
or U31202 (N_31202,N_30566,N_30068);
and U31203 (N_31203,N_30642,N_30229);
nand U31204 (N_31204,N_30492,N_30774);
and U31205 (N_31205,N_30721,N_30488);
xnor U31206 (N_31206,N_30342,N_30339);
nor U31207 (N_31207,N_30626,N_30236);
xor U31208 (N_31208,N_30472,N_30926);
xor U31209 (N_31209,N_30556,N_30916);
xnor U31210 (N_31210,N_30104,N_30996);
nand U31211 (N_31211,N_30635,N_30408);
nand U31212 (N_31212,N_30864,N_30548);
nor U31213 (N_31213,N_30734,N_30019);
nor U31214 (N_31214,N_30009,N_30617);
nand U31215 (N_31215,N_30133,N_30827);
nor U31216 (N_31216,N_30092,N_30406);
nor U31217 (N_31217,N_30549,N_30162);
xnor U31218 (N_31218,N_30563,N_30200);
and U31219 (N_31219,N_30880,N_30875);
xnor U31220 (N_31220,N_30383,N_30844);
and U31221 (N_31221,N_30124,N_30081);
or U31222 (N_31222,N_30718,N_30573);
or U31223 (N_31223,N_30415,N_30629);
and U31224 (N_31224,N_30463,N_30489);
or U31225 (N_31225,N_30674,N_30308);
xnor U31226 (N_31226,N_30812,N_30947);
nand U31227 (N_31227,N_30411,N_30681);
and U31228 (N_31228,N_30690,N_30115);
nor U31229 (N_31229,N_30291,N_30507);
and U31230 (N_31230,N_30555,N_30751);
and U31231 (N_31231,N_30024,N_30512);
or U31232 (N_31232,N_30484,N_30407);
and U31233 (N_31233,N_30255,N_30966);
and U31234 (N_31234,N_30603,N_30008);
or U31235 (N_31235,N_30789,N_30438);
or U31236 (N_31236,N_30706,N_30874);
and U31237 (N_31237,N_30676,N_30520);
xor U31238 (N_31238,N_30891,N_30987);
or U31239 (N_31239,N_30466,N_30813);
and U31240 (N_31240,N_30242,N_30641);
nor U31241 (N_31241,N_30084,N_30005);
and U31242 (N_31242,N_30015,N_30513);
and U31243 (N_31243,N_30539,N_30220);
or U31244 (N_31244,N_30988,N_30059);
nor U31245 (N_31245,N_30206,N_30095);
and U31246 (N_31246,N_30935,N_30455);
nor U31247 (N_31247,N_30853,N_30523);
or U31248 (N_31248,N_30469,N_30420);
or U31249 (N_31249,N_30560,N_30982);
xnor U31250 (N_31250,N_30738,N_30350);
or U31251 (N_31251,N_30834,N_30139);
and U31252 (N_31252,N_30733,N_30479);
nand U31253 (N_31253,N_30737,N_30724);
nor U31254 (N_31254,N_30893,N_30787);
xor U31255 (N_31255,N_30209,N_30589);
xor U31256 (N_31256,N_30806,N_30648);
or U31257 (N_31257,N_30604,N_30883);
xor U31258 (N_31258,N_30072,N_30496);
nor U31259 (N_31259,N_30249,N_30006);
and U31260 (N_31260,N_30804,N_30102);
nor U31261 (N_31261,N_30928,N_30636);
xnor U31262 (N_31262,N_30493,N_30803);
and U31263 (N_31263,N_30145,N_30314);
and U31264 (N_31264,N_30219,N_30991);
and U31265 (N_31265,N_30082,N_30775);
nand U31266 (N_31266,N_30704,N_30992);
xor U31267 (N_31267,N_30614,N_30647);
and U31268 (N_31268,N_30682,N_30299);
or U31269 (N_31269,N_30968,N_30752);
nor U31270 (N_31270,N_30478,N_30885);
nand U31271 (N_31271,N_30385,N_30231);
nor U31272 (N_31272,N_30990,N_30273);
nand U31273 (N_31273,N_30678,N_30577);
and U31274 (N_31274,N_30204,N_30402);
nand U31275 (N_31275,N_30802,N_30422);
nand U31276 (N_31276,N_30130,N_30773);
and U31277 (N_31277,N_30177,N_30783);
nand U31278 (N_31278,N_30051,N_30554);
nor U31279 (N_31279,N_30141,N_30475);
or U31280 (N_31280,N_30688,N_30213);
or U31281 (N_31281,N_30829,N_30228);
or U31282 (N_31282,N_30160,N_30873);
xnor U31283 (N_31283,N_30728,N_30828);
and U31284 (N_31284,N_30003,N_30952);
and U31285 (N_31285,N_30963,N_30655);
or U31286 (N_31286,N_30795,N_30984);
xor U31287 (N_31287,N_30881,N_30243);
or U31288 (N_31288,N_30753,N_30845);
nor U31289 (N_31289,N_30192,N_30465);
or U31290 (N_31290,N_30677,N_30368);
and U31291 (N_31291,N_30755,N_30964);
xor U31292 (N_31292,N_30581,N_30306);
xor U31293 (N_31293,N_30759,N_30309);
and U31294 (N_31294,N_30840,N_30651);
xor U31295 (N_31295,N_30876,N_30346);
nand U31296 (N_31296,N_30021,N_30268);
nor U31297 (N_31297,N_30012,N_30318);
and U31298 (N_31298,N_30810,N_30078);
xor U31299 (N_31299,N_30970,N_30359);
xnor U31300 (N_31300,N_30125,N_30637);
and U31301 (N_31301,N_30226,N_30969);
xor U31302 (N_31302,N_30999,N_30819);
or U31303 (N_31303,N_30776,N_30522);
or U31304 (N_31304,N_30659,N_30793);
xor U31305 (N_31305,N_30022,N_30106);
xnor U31306 (N_31306,N_30113,N_30790);
nor U31307 (N_31307,N_30440,N_30432);
xnor U31308 (N_31308,N_30174,N_30505);
and U31309 (N_31309,N_30780,N_30154);
or U31310 (N_31310,N_30550,N_30395);
nor U31311 (N_31311,N_30363,N_30053);
or U31312 (N_31312,N_30857,N_30178);
or U31313 (N_31313,N_30510,N_30043);
nor U31314 (N_31314,N_30252,N_30836);
and U31315 (N_31315,N_30396,N_30374);
xnor U31316 (N_31316,N_30356,N_30696);
xnor U31317 (N_31317,N_30114,N_30877);
nor U31318 (N_31318,N_30060,N_30657);
and U31319 (N_31319,N_30216,N_30527);
nand U31320 (N_31320,N_30946,N_30361);
xor U31321 (N_31321,N_30170,N_30132);
nand U31322 (N_31322,N_30822,N_30616);
nand U31323 (N_31323,N_30085,N_30093);
nand U31324 (N_31324,N_30424,N_30565);
or U31325 (N_31325,N_30090,N_30511);
nor U31326 (N_31326,N_30761,N_30435);
nor U31327 (N_31327,N_30358,N_30153);
nor U31328 (N_31328,N_30474,N_30312);
and U31329 (N_31329,N_30823,N_30973);
and U31330 (N_31330,N_30825,N_30427);
xor U31331 (N_31331,N_30772,N_30014);
or U31332 (N_31332,N_30486,N_30167);
nand U31333 (N_31333,N_30913,N_30770);
xor U31334 (N_31334,N_30344,N_30338);
nand U31335 (N_31335,N_30923,N_30185);
xnor U31336 (N_31336,N_30142,N_30860);
nand U31337 (N_31337,N_30727,N_30483);
and U31338 (N_31338,N_30304,N_30934);
xor U31339 (N_31339,N_30058,N_30369);
or U31340 (N_31340,N_30109,N_30332);
xor U31341 (N_31341,N_30382,N_30272);
nor U31342 (N_31342,N_30663,N_30190);
and U31343 (N_31343,N_30075,N_30275);
and U31344 (N_31344,N_30256,N_30376);
or U31345 (N_31345,N_30234,N_30107);
and U31346 (N_31346,N_30887,N_30516);
xnor U31347 (N_31347,N_30165,N_30895);
nand U31348 (N_31348,N_30205,N_30767);
and U31349 (N_31349,N_30953,N_30343);
nor U31350 (N_31350,N_30189,N_30785);
nor U31351 (N_31351,N_30140,N_30720);
nor U31352 (N_31352,N_30071,N_30451);
nor U31353 (N_31353,N_30949,N_30818);
nand U31354 (N_31354,N_30295,N_30937);
xnor U31355 (N_31355,N_30335,N_30660);
or U31356 (N_31356,N_30416,N_30010);
nor U31357 (N_31357,N_30253,N_30799);
nor U31358 (N_31358,N_30584,N_30715);
nand U31359 (N_31359,N_30627,N_30671);
nand U31360 (N_31360,N_30506,N_30498);
or U31361 (N_31361,N_30717,N_30575);
nor U31362 (N_31362,N_30246,N_30262);
nor U31363 (N_31363,N_30062,N_30693);
nand U31364 (N_31364,N_30643,N_30297);
nor U31365 (N_31365,N_30418,N_30612);
and U31366 (N_31366,N_30431,N_30533);
xor U31367 (N_31367,N_30351,N_30101);
or U31368 (N_31368,N_30117,N_30048);
or U31369 (N_31369,N_30797,N_30552);
xor U31370 (N_31370,N_30993,N_30628);
xnor U31371 (N_31371,N_30569,N_30079);
or U31372 (N_31372,N_30201,N_30529);
and U31373 (N_31373,N_30666,N_30248);
nand U31374 (N_31374,N_30514,N_30699);
or U31375 (N_31375,N_30270,N_30754);
and U31376 (N_31376,N_30386,N_30279);
nand U31377 (N_31377,N_30159,N_30193);
nand U31378 (N_31378,N_30786,N_30736);
nand U31379 (N_31379,N_30217,N_30652);
or U31380 (N_31380,N_30779,N_30664);
nand U31381 (N_31381,N_30049,N_30063);
and U31382 (N_31382,N_30322,N_30070);
nor U31383 (N_31383,N_30945,N_30965);
nand U31384 (N_31384,N_30526,N_30430);
nor U31385 (N_31385,N_30137,N_30897);
nor U31386 (N_31386,N_30692,N_30929);
nand U31387 (N_31387,N_30975,N_30568);
nor U31388 (N_31388,N_30631,N_30453);
xor U31389 (N_31389,N_30276,N_30833);
and U31390 (N_31390,N_30443,N_30835);
and U31391 (N_31391,N_30707,N_30271);
xor U31392 (N_31392,N_30045,N_30083);
or U31393 (N_31393,N_30277,N_30481);
nand U31394 (N_31394,N_30316,N_30181);
xor U31395 (N_31395,N_30148,N_30852);
xor U31396 (N_31396,N_30862,N_30331);
nor U31397 (N_31397,N_30670,N_30914);
nand U31398 (N_31398,N_30175,N_30321);
or U31399 (N_31399,N_30147,N_30578);
or U31400 (N_31400,N_30858,N_30691);
nand U31401 (N_31401,N_30292,N_30149);
nand U31402 (N_31402,N_30675,N_30477);
nand U31403 (N_31403,N_30100,N_30452);
nand U31404 (N_31404,N_30239,N_30794);
and U31405 (N_31405,N_30254,N_30890);
nor U31406 (N_31406,N_30960,N_30889);
and U31407 (N_31407,N_30450,N_30632);
and U31408 (N_31408,N_30426,N_30462);
nand U31409 (N_31409,N_30194,N_30602);
nand U31410 (N_31410,N_30264,N_30195);
xnor U31411 (N_31411,N_30151,N_30805);
nand U31412 (N_31412,N_30931,N_30476);
and U31413 (N_31413,N_30354,N_30583);
and U31414 (N_31414,N_30313,N_30576);
xnor U31415 (N_31415,N_30135,N_30709);
xor U31416 (N_31416,N_30057,N_30564);
nor U31417 (N_31417,N_30542,N_30161);
or U31418 (N_31418,N_30448,N_30064);
nand U31419 (N_31419,N_30025,N_30169);
xnor U31420 (N_31420,N_30939,N_30000);
and U31421 (N_31421,N_30615,N_30377);
xor U31422 (N_31422,N_30419,N_30155);
or U31423 (N_31423,N_30994,N_30023);
and U31424 (N_31424,N_30537,N_30080);
or U31425 (N_31425,N_30762,N_30919);
or U31426 (N_31426,N_30258,N_30624);
and U31427 (N_31427,N_30644,N_30599);
or U31428 (N_31428,N_30672,N_30445);
or U31429 (N_31429,N_30713,N_30144);
or U31430 (N_31430,N_30851,N_30817);
or U31431 (N_31431,N_30182,N_30694);
nor U31432 (N_31432,N_30116,N_30630);
nand U31433 (N_31433,N_30888,N_30401);
and U31434 (N_31434,N_30743,N_30985);
nand U31435 (N_31435,N_30850,N_30247);
xnor U31436 (N_31436,N_30972,N_30768);
and U31437 (N_31437,N_30428,N_30705);
and U31438 (N_31438,N_30384,N_30390);
nand U31439 (N_31439,N_30348,N_30962);
or U31440 (N_31440,N_30380,N_30037);
and U31441 (N_31441,N_30519,N_30899);
or U31442 (N_31442,N_30719,N_30482);
or U31443 (N_31443,N_30357,N_30412);
nand U31444 (N_31444,N_30515,N_30842);
or U31445 (N_31445,N_30237,N_30156);
nor U31446 (N_31446,N_30608,N_30855);
xor U31447 (N_31447,N_30906,N_30241);
nand U31448 (N_31448,N_30340,N_30449);
nand U31449 (N_31449,N_30120,N_30521);
or U31450 (N_31450,N_30668,N_30882);
nand U31451 (N_31451,N_30077,N_30372);
or U31452 (N_31452,N_30536,N_30854);
nor U31453 (N_31453,N_30055,N_30856);
or U31454 (N_31454,N_30532,N_30446);
nand U31455 (N_31455,N_30765,N_30371);
and U31456 (N_31456,N_30355,N_30423);
nor U31457 (N_31457,N_30961,N_30665);
and U31458 (N_31458,N_30261,N_30896);
nor U31459 (N_31459,N_30389,N_30685);
or U31460 (N_31460,N_30168,N_30640);
and U31461 (N_31461,N_30353,N_30683);
nor U31462 (N_31462,N_30995,N_30280);
and U31463 (N_31463,N_30250,N_30121);
xnor U31464 (N_31464,N_30703,N_30285);
nor U31465 (N_31465,N_30294,N_30625);
or U31466 (N_31466,N_30315,N_30222);
nand U31467 (N_31467,N_30815,N_30917);
or U31468 (N_31468,N_30286,N_30832);
xor U31469 (N_31469,N_30574,N_30938);
xor U31470 (N_31470,N_30714,N_30047);
or U31471 (N_31471,N_30980,N_30781);
and U31472 (N_31472,N_30122,N_30119);
xnor U31473 (N_31473,N_30183,N_30546);
and U31474 (N_31474,N_30747,N_30163);
nand U31475 (N_31475,N_30067,N_30052);
xor U31476 (N_31476,N_30517,N_30311);
nand U31477 (N_31477,N_30571,N_30826);
nor U31478 (N_31478,N_30397,N_30065);
and U31479 (N_31479,N_30530,N_30639);
xnor U31480 (N_31480,N_30967,N_30807);
or U31481 (N_31481,N_30686,N_30467);
xnor U31482 (N_31482,N_30417,N_30908);
xnor U31483 (N_31483,N_30186,N_30769);
or U31484 (N_31484,N_30601,N_30865);
nand U31485 (N_31485,N_30950,N_30989);
or U31486 (N_31486,N_30503,N_30701);
nand U31487 (N_31487,N_30098,N_30373);
xnor U31488 (N_31488,N_30958,N_30903);
and U31489 (N_31489,N_30846,N_30838);
or U31490 (N_31490,N_30600,N_30387);
or U31491 (N_31491,N_30341,N_30370);
xor U31492 (N_31492,N_30977,N_30901);
nand U31493 (N_31493,N_30127,N_30595);
xnor U31494 (N_31494,N_30042,N_30263);
nand U31495 (N_31495,N_30240,N_30074);
and U31496 (N_31496,N_30129,N_30066);
nor U31497 (N_31497,N_30500,N_30796);
and U31498 (N_31498,N_30225,N_30110);
xnor U31499 (N_31499,N_30087,N_30712);
and U31500 (N_31500,N_30159,N_30859);
or U31501 (N_31501,N_30679,N_30456);
and U31502 (N_31502,N_30237,N_30311);
or U31503 (N_31503,N_30380,N_30553);
or U31504 (N_31504,N_30009,N_30969);
nor U31505 (N_31505,N_30096,N_30446);
and U31506 (N_31506,N_30505,N_30059);
nor U31507 (N_31507,N_30581,N_30370);
nand U31508 (N_31508,N_30533,N_30542);
or U31509 (N_31509,N_30680,N_30657);
and U31510 (N_31510,N_30575,N_30461);
nand U31511 (N_31511,N_30846,N_30878);
xor U31512 (N_31512,N_30634,N_30725);
nand U31513 (N_31513,N_30323,N_30707);
and U31514 (N_31514,N_30119,N_30089);
xor U31515 (N_31515,N_30045,N_30356);
nor U31516 (N_31516,N_30107,N_30469);
nand U31517 (N_31517,N_30525,N_30429);
xor U31518 (N_31518,N_30795,N_30417);
or U31519 (N_31519,N_30451,N_30329);
and U31520 (N_31520,N_30286,N_30398);
and U31521 (N_31521,N_30578,N_30825);
xnor U31522 (N_31522,N_30619,N_30689);
xor U31523 (N_31523,N_30094,N_30143);
nand U31524 (N_31524,N_30504,N_30478);
xor U31525 (N_31525,N_30535,N_30728);
nand U31526 (N_31526,N_30789,N_30064);
nor U31527 (N_31527,N_30133,N_30596);
and U31528 (N_31528,N_30560,N_30519);
and U31529 (N_31529,N_30323,N_30815);
or U31530 (N_31530,N_30440,N_30300);
nand U31531 (N_31531,N_30368,N_30238);
nor U31532 (N_31532,N_30754,N_30732);
nand U31533 (N_31533,N_30369,N_30119);
nor U31534 (N_31534,N_30125,N_30948);
or U31535 (N_31535,N_30018,N_30619);
nand U31536 (N_31536,N_30560,N_30842);
nor U31537 (N_31537,N_30297,N_30919);
or U31538 (N_31538,N_30225,N_30740);
or U31539 (N_31539,N_30036,N_30057);
or U31540 (N_31540,N_30838,N_30309);
and U31541 (N_31541,N_30251,N_30512);
nor U31542 (N_31542,N_30601,N_30069);
or U31543 (N_31543,N_30091,N_30559);
nand U31544 (N_31544,N_30407,N_30962);
or U31545 (N_31545,N_30389,N_30226);
xor U31546 (N_31546,N_30525,N_30256);
nor U31547 (N_31547,N_30788,N_30397);
or U31548 (N_31548,N_30378,N_30532);
or U31549 (N_31549,N_30037,N_30310);
nor U31550 (N_31550,N_30436,N_30655);
or U31551 (N_31551,N_30368,N_30159);
nand U31552 (N_31552,N_30524,N_30556);
nand U31553 (N_31553,N_30386,N_30511);
xnor U31554 (N_31554,N_30132,N_30326);
and U31555 (N_31555,N_30976,N_30994);
xnor U31556 (N_31556,N_30719,N_30581);
nor U31557 (N_31557,N_30449,N_30847);
nor U31558 (N_31558,N_30589,N_30814);
nand U31559 (N_31559,N_30504,N_30241);
or U31560 (N_31560,N_30743,N_30874);
and U31561 (N_31561,N_30075,N_30553);
xor U31562 (N_31562,N_30170,N_30568);
nor U31563 (N_31563,N_30480,N_30084);
nand U31564 (N_31564,N_30982,N_30039);
nor U31565 (N_31565,N_30683,N_30773);
nor U31566 (N_31566,N_30281,N_30396);
xor U31567 (N_31567,N_30709,N_30306);
or U31568 (N_31568,N_30772,N_30624);
and U31569 (N_31569,N_30678,N_30305);
nor U31570 (N_31570,N_30414,N_30542);
nand U31571 (N_31571,N_30847,N_30455);
or U31572 (N_31572,N_30511,N_30033);
xor U31573 (N_31573,N_30597,N_30578);
nand U31574 (N_31574,N_30025,N_30097);
nand U31575 (N_31575,N_30083,N_30889);
nor U31576 (N_31576,N_30029,N_30393);
xnor U31577 (N_31577,N_30924,N_30945);
nor U31578 (N_31578,N_30886,N_30657);
and U31579 (N_31579,N_30175,N_30409);
nand U31580 (N_31580,N_30820,N_30546);
or U31581 (N_31581,N_30401,N_30487);
nand U31582 (N_31582,N_30889,N_30354);
nand U31583 (N_31583,N_30147,N_30830);
xnor U31584 (N_31584,N_30526,N_30972);
xor U31585 (N_31585,N_30068,N_30814);
xor U31586 (N_31586,N_30143,N_30679);
nor U31587 (N_31587,N_30773,N_30378);
nand U31588 (N_31588,N_30541,N_30588);
or U31589 (N_31589,N_30201,N_30803);
and U31590 (N_31590,N_30943,N_30633);
xor U31591 (N_31591,N_30996,N_30287);
or U31592 (N_31592,N_30434,N_30137);
or U31593 (N_31593,N_30447,N_30118);
or U31594 (N_31594,N_30607,N_30592);
or U31595 (N_31595,N_30628,N_30491);
or U31596 (N_31596,N_30154,N_30931);
or U31597 (N_31597,N_30250,N_30499);
or U31598 (N_31598,N_30205,N_30510);
or U31599 (N_31599,N_30367,N_30576);
nand U31600 (N_31600,N_30027,N_30817);
nand U31601 (N_31601,N_30171,N_30786);
nand U31602 (N_31602,N_30866,N_30435);
nand U31603 (N_31603,N_30038,N_30171);
nand U31604 (N_31604,N_30506,N_30320);
nand U31605 (N_31605,N_30442,N_30468);
nor U31606 (N_31606,N_30840,N_30681);
xor U31607 (N_31607,N_30814,N_30532);
xor U31608 (N_31608,N_30118,N_30459);
or U31609 (N_31609,N_30804,N_30023);
nor U31610 (N_31610,N_30486,N_30056);
or U31611 (N_31611,N_30271,N_30554);
nand U31612 (N_31612,N_30897,N_30213);
xnor U31613 (N_31613,N_30845,N_30836);
xnor U31614 (N_31614,N_30700,N_30916);
xnor U31615 (N_31615,N_30428,N_30537);
or U31616 (N_31616,N_30758,N_30296);
nand U31617 (N_31617,N_30788,N_30071);
and U31618 (N_31618,N_30632,N_30242);
nor U31619 (N_31619,N_30292,N_30706);
xor U31620 (N_31620,N_30617,N_30653);
nor U31621 (N_31621,N_30174,N_30191);
nand U31622 (N_31622,N_30016,N_30807);
nand U31623 (N_31623,N_30712,N_30390);
nand U31624 (N_31624,N_30042,N_30130);
nor U31625 (N_31625,N_30543,N_30220);
nor U31626 (N_31626,N_30205,N_30684);
nand U31627 (N_31627,N_30015,N_30160);
nand U31628 (N_31628,N_30207,N_30346);
xnor U31629 (N_31629,N_30069,N_30298);
and U31630 (N_31630,N_30043,N_30316);
xor U31631 (N_31631,N_30122,N_30244);
and U31632 (N_31632,N_30184,N_30148);
or U31633 (N_31633,N_30636,N_30446);
nand U31634 (N_31634,N_30165,N_30581);
or U31635 (N_31635,N_30687,N_30377);
or U31636 (N_31636,N_30232,N_30568);
nand U31637 (N_31637,N_30599,N_30686);
xnor U31638 (N_31638,N_30363,N_30289);
nor U31639 (N_31639,N_30546,N_30427);
or U31640 (N_31640,N_30787,N_30759);
xnor U31641 (N_31641,N_30640,N_30492);
and U31642 (N_31642,N_30014,N_30659);
nand U31643 (N_31643,N_30308,N_30649);
xor U31644 (N_31644,N_30135,N_30256);
and U31645 (N_31645,N_30988,N_30707);
xnor U31646 (N_31646,N_30790,N_30400);
or U31647 (N_31647,N_30318,N_30963);
nand U31648 (N_31648,N_30384,N_30290);
nor U31649 (N_31649,N_30903,N_30852);
nor U31650 (N_31650,N_30180,N_30515);
xnor U31651 (N_31651,N_30292,N_30093);
nor U31652 (N_31652,N_30303,N_30434);
and U31653 (N_31653,N_30249,N_30938);
nor U31654 (N_31654,N_30889,N_30128);
and U31655 (N_31655,N_30124,N_30000);
or U31656 (N_31656,N_30953,N_30488);
or U31657 (N_31657,N_30135,N_30058);
nor U31658 (N_31658,N_30971,N_30177);
nand U31659 (N_31659,N_30426,N_30056);
xnor U31660 (N_31660,N_30618,N_30429);
nor U31661 (N_31661,N_30613,N_30734);
nor U31662 (N_31662,N_30729,N_30576);
and U31663 (N_31663,N_30083,N_30046);
nand U31664 (N_31664,N_30690,N_30346);
xor U31665 (N_31665,N_30187,N_30992);
or U31666 (N_31666,N_30180,N_30245);
and U31667 (N_31667,N_30236,N_30233);
xnor U31668 (N_31668,N_30660,N_30642);
nor U31669 (N_31669,N_30369,N_30008);
or U31670 (N_31670,N_30218,N_30585);
and U31671 (N_31671,N_30545,N_30785);
nor U31672 (N_31672,N_30729,N_30281);
nor U31673 (N_31673,N_30512,N_30782);
xor U31674 (N_31674,N_30620,N_30680);
xnor U31675 (N_31675,N_30458,N_30368);
or U31676 (N_31676,N_30086,N_30029);
nand U31677 (N_31677,N_30714,N_30036);
nor U31678 (N_31678,N_30811,N_30083);
nor U31679 (N_31679,N_30505,N_30176);
or U31680 (N_31680,N_30848,N_30207);
nand U31681 (N_31681,N_30638,N_30181);
and U31682 (N_31682,N_30614,N_30604);
xnor U31683 (N_31683,N_30309,N_30442);
nor U31684 (N_31684,N_30606,N_30276);
nor U31685 (N_31685,N_30428,N_30891);
xnor U31686 (N_31686,N_30875,N_30066);
and U31687 (N_31687,N_30558,N_30352);
or U31688 (N_31688,N_30286,N_30088);
xnor U31689 (N_31689,N_30626,N_30121);
xor U31690 (N_31690,N_30171,N_30643);
xor U31691 (N_31691,N_30346,N_30622);
or U31692 (N_31692,N_30242,N_30975);
or U31693 (N_31693,N_30099,N_30289);
or U31694 (N_31694,N_30697,N_30419);
xnor U31695 (N_31695,N_30207,N_30241);
nand U31696 (N_31696,N_30216,N_30620);
and U31697 (N_31697,N_30590,N_30994);
nor U31698 (N_31698,N_30889,N_30151);
or U31699 (N_31699,N_30485,N_30307);
xnor U31700 (N_31700,N_30483,N_30768);
nand U31701 (N_31701,N_30431,N_30566);
or U31702 (N_31702,N_30465,N_30696);
nor U31703 (N_31703,N_30556,N_30219);
nor U31704 (N_31704,N_30367,N_30604);
nor U31705 (N_31705,N_30324,N_30008);
and U31706 (N_31706,N_30231,N_30623);
and U31707 (N_31707,N_30096,N_30845);
or U31708 (N_31708,N_30515,N_30653);
nor U31709 (N_31709,N_30190,N_30645);
nor U31710 (N_31710,N_30553,N_30032);
and U31711 (N_31711,N_30304,N_30262);
nor U31712 (N_31712,N_30079,N_30437);
nor U31713 (N_31713,N_30506,N_30222);
or U31714 (N_31714,N_30193,N_30536);
xor U31715 (N_31715,N_30043,N_30049);
nor U31716 (N_31716,N_30375,N_30345);
nor U31717 (N_31717,N_30686,N_30117);
and U31718 (N_31718,N_30283,N_30861);
nor U31719 (N_31719,N_30414,N_30871);
nand U31720 (N_31720,N_30432,N_30964);
or U31721 (N_31721,N_30235,N_30553);
nand U31722 (N_31722,N_30981,N_30141);
nor U31723 (N_31723,N_30641,N_30903);
or U31724 (N_31724,N_30738,N_30429);
or U31725 (N_31725,N_30236,N_30926);
nand U31726 (N_31726,N_30060,N_30416);
nand U31727 (N_31727,N_30177,N_30299);
and U31728 (N_31728,N_30504,N_30985);
xor U31729 (N_31729,N_30785,N_30288);
or U31730 (N_31730,N_30251,N_30040);
nand U31731 (N_31731,N_30138,N_30253);
xor U31732 (N_31732,N_30304,N_30826);
nor U31733 (N_31733,N_30838,N_30422);
and U31734 (N_31734,N_30924,N_30022);
or U31735 (N_31735,N_30452,N_30367);
and U31736 (N_31736,N_30589,N_30925);
nor U31737 (N_31737,N_30309,N_30967);
nand U31738 (N_31738,N_30210,N_30561);
or U31739 (N_31739,N_30474,N_30528);
nand U31740 (N_31740,N_30178,N_30911);
nand U31741 (N_31741,N_30896,N_30761);
nor U31742 (N_31742,N_30359,N_30336);
nor U31743 (N_31743,N_30111,N_30330);
nand U31744 (N_31744,N_30199,N_30537);
nand U31745 (N_31745,N_30380,N_30880);
and U31746 (N_31746,N_30677,N_30439);
xor U31747 (N_31747,N_30290,N_30971);
xor U31748 (N_31748,N_30352,N_30633);
nor U31749 (N_31749,N_30221,N_30487);
nor U31750 (N_31750,N_30683,N_30380);
xor U31751 (N_31751,N_30639,N_30178);
or U31752 (N_31752,N_30274,N_30767);
nor U31753 (N_31753,N_30348,N_30014);
nand U31754 (N_31754,N_30579,N_30314);
or U31755 (N_31755,N_30204,N_30060);
xor U31756 (N_31756,N_30456,N_30172);
xor U31757 (N_31757,N_30981,N_30850);
or U31758 (N_31758,N_30552,N_30566);
nor U31759 (N_31759,N_30399,N_30189);
or U31760 (N_31760,N_30420,N_30884);
xor U31761 (N_31761,N_30294,N_30134);
nor U31762 (N_31762,N_30701,N_30554);
or U31763 (N_31763,N_30542,N_30976);
nand U31764 (N_31764,N_30459,N_30467);
or U31765 (N_31765,N_30906,N_30496);
or U31766 (N_31766,N_30146,N_30930);
or U31767 (N_31767,N_30591,N_30056);
or U31768 (N_31768,N_30811,N_30631);
and U31769 (N_31769,N_30968,N_30271);
and U31770 (N_31770,N_30916,N_30344);
xor U31771 (N_31771,N_30543,N_30748);
nand U31772 (N_31772,N_30785,N_30536);
xor U31773 (N_31773,N_30538,N_30436);
xnor U31774 (N_31774,N_30709,N_30891);
and U31775 (N_31775,N_30972,N_30290);
or U31776 (N_31776,N_30953,N_30228);
nor U31777 (N_31777,N_30453,N_30701);
and U31778 (N_31778,N_30660,N_30400);
nor U31779 (N_31779,N_30278,N_30455);
nor U31780 (N_31780,N_30198,N_30478);
xnor U31781 (N_31781,N_30192,N_30461);
and U31782 (N_31782,N_30219,N_30597);
or U31783 (N_31783,N_30233,N_30729);
nor U31784 (N_31784,N_30197,N_30260);
nor U31785 (N_31785,N_30514,N_30336);
nor U31786 (N_31786,N_30740,N_30308);
nor U31787 (N_31787,N_30220,N_30258);
nand U31788 (N_31788,N_30222,N_30773);
nor U31789 (N_31789,N_30642,N_30581);
or U31790 (N_31790,N_30763,N_30206);
xnor U31791 (N_31791,N_30405,N_30840);
nand U31792 (N_31792,N_30140,N_30248);
nor U31793 (N_31793,N_30563,N_30633);
nor U31794 (N_31794,N_30946,N_30435);
or U31795 (N_31795,N_30007,N_30618);
nand U31796 (N_31796,N_30680,N_30036);
nor U31797 (N_31797,N_30094,N_30741);
nor U31798 (N_31798,N_30760,N_30526);
and U31799 (N_31799,N_30296,N_30516);
xor U31800 (N_31800,N_30238,N_30859);
nand U31801 (N_31801,N_30134,N_30438);
and U31802 (N_31802,N_30346,N_30531);
and U31803 (N_31803,N_30617,N_30949);
or U31804 (N_31804,N_30877,N_30408);
or U31805 (N_31805,N_30294,N_30732);
nor U31806 (N_31806,N_30889,N_30844);
and U31807 (N_31807,N_30976,N_30597);
xnor U31808 (N_31808,N_30046,N_30713);
or U31809 (N_31809,N_30894,N_30221);
and U31810 (N_31810,N_30535,N_30662);
and U31811 (N_31811,N_30617,N_30715);
nand U31812 (N_31812,N_30987,N_30882);
nor U31813 (N_31813,N_30206,N_30969);
or U31814 (N_31814,N_30290,N_30724);
xor U31815 (N_31815,N_30325,N_30291);
or U31816 (N_31816,N_30851,N_30215);
xor U31817 (N_31817,N_30424,N_30473);
and U31818 (N_31818,N_30551,N_30104);
nor U31819 (N_31819,N_30256,N_30035);
or U31820 (N_31820,N_30595,N_30596);
and U31821 (N_31821,N_30218,N_30373);
xnor U31822 (N_31822,N_30659,N_30789);
nor U31823 (N_31823,N_30164,N_30882);
nor U31824 (N_31824,N_30587,N_30682);
or U31825 (N_31825,N_30488,N_30179);
nor U31826 (N_31826,N_30455,N_30529);
nand U31827 (N_31827,N_30706,N_30328);
nor U31828 (N_31828,N_30571,N_30574);
nand U31829 (N_31829,N_30754,N_30509);
nor U31830 (N_31830,N_30063,N_30802);
xnor U31831 (N_31831,N_30592,N_30890);
or U31832 (N_31832,N_30423,N_30346);
xor U31833 (N_31833,N_30543,N_30913);
xnor U31834 (N_31834,N_30276,N_30632);
or U31835 (N_31835,N_30165,N_30833);
nand U31836 (N_31836,N_30238,N_30213);
nand U31837 (N_31837,N_30873,N_30987);
and U31838 (N_31838,N_30189,N_30670);
or U31839 (N_31839,N_30121,N_30562);
and U31840 (N_31840,N_30184,N_30373);
xnor U31841 (N_31841,N_30186,N_30488);
or U31842 (N_31842,N_30400,N_30582);
nand U31843 (N_31843,N_30639,N_30004);
and U31844 (N_31844,N_30678,N_30399);
nor U31845 (N_31845,N_30859,N_30436);
nor U31846 (N_31846,N_30916,N_30236);
and U31847 (N_31847,N_30928,N_30402);
nand U31848 (N_31848,N_30524,N_30940);
and U31849 (N_31849,N_30078,N_30881);
or U31850 (N_31850,N_30876,N_30238);
and U31851 (N_31851,N_30389,N_30918);
xor U31852 (N_31852,N_30613,N_30760);
and U31853 (N_31853,N_30441,N_30679);
nand U31854 (N_31854,N_30315,N_30152);
and U31855 (N_31855,N_30140,N_30607);
nand U31856 (N_31856,N_30626,N_30954);
nor U31857 (N_31857,N_30774,N_30151);
or U31858 (N_31858,N_30996,N_30538);
and U31859 (N_31859,N_30233,N_30026);
and U31860 (N_31860,N_30788,N_30128);
and U31861 (N_31861,N_30613,N_30773);
or U31862 (N_31862,N_30833,N_30517);
or U31863 (N_31863,N_30667,N_30422);
or U31864 (N_31864,N_30855,N_30406);
xnor U31865 (N_31865,N_30264,N_30818);
nor U31866 (N_31866,N_30592,N_30394);
nor U31867 (N_31867,N_30122,N_30469);
nand U31868 (N_31868,N_30102,N_30709);
nand U31869 (N_31869,N_30638,N_30458);
nor U31870 (N_31870,N_30278,N_30100);
nand U31871 (N_31871,N_30033,N_30687);
nor U31872 (N_31872,N_30455,N_30686);
nor U31873 (N_31873,N_30298,N_30354);
or U31874 (N_31874,N_30819,N_30097);
xnor U31875 (N_31875,N_30957,N_30141);
xor U31876 (N_31876,N_30752,N_30523);
xnor U31877 (N_31877,N_30606,N_30585);
nand U31878 (N_31878,N_30451,N_30923);
xor U31879 (N_31879,N_30216,N_30256);
or U31880 (N_31880,N_30454,N_30642);
nand U31881 (N_31881,N_30619,N_30702);
or U31882 (N_31882,N_30087,N_30093);
or U31883 (N_31883,N_30755,N_30398);
or U31884 (N_31884,N_30157,N_30487);
nor U31885 (N_31885,N_30651,N_30978);
and U31886 (N_31886,N_30957,N_30230);
nand U31887 (N_31887,N_30826,N_30590);
nor U31888 (N_31888,N_30496,N_30330);
and U31889 (N_31889,N_30499,N_30350);
or U31890 (N_31890,N_30484,N_30292);
nor U31891 (N_31891,N_30243,N_30392);
nor U31892 (N_31892,N_30493,N_30796);
nand U31893 (N_31893,N_30441,N_30049);
xor U31894 (N_31894,N_30211,N_30481);
nand U31895 (N_31895,N_30827,N_30975);
nand U31896 (N_31896,N_30709,N_30571);
or U31897 (N_31897,N_30333,N_30644);
nor U31898 (N_31898,N_30347,N_30929);
xor U31899 (N_31899,N_30261,N_30426);
nor U31900 (N_31900,N_30659,N_30352);
nor U31901 (N_31901,N_30977,N_30083);
nand U31902 (N_31902,N_30547,N_30926);
xor U31903 (N_31903,N_30404,N_30281);
nand U31904 (N_31904,N_30650,N_30739);
nand U31905 (N_31905,N_30458,N_30830);
and U31906 (N_31906,N_30773,N_30131);
and U31907 (N_31907,N_30113,N_30364);
or U31908 (N_31908,N_30805,N_30251);
and U31909 (N_31909,N_30048,N_30776);
and U31910 (N_31910,N_30667,N_30624);
xnor U31911 (N_31911,N_30121,N_30248);
xor U31912 (N_31912,N_30386,N_30878);
nor U31913 (N_31913,N_30823,N_30571);
xnor U31914 (N_31914,N_30883,N_30236);
and U31915 (N_31915,N_30314,N_30757);
and U31916 (N_31916,N_30125,N_30055);
xor U31917 (N_31917,N_30446,N_30589);
xor U31918 (N_31918,N_30927,N_30478);
nor U31919 (N_31919,N_30135,N_30339);
xnor U31920 (N_31920,N_30277,N_30540);
nor U31921 (N_31921,N_30397,N_30103);
or U31922 (N_31922,N_30884,N_30497);
xor U31923 (N_31923,N_30319,N_30097);
and U31924 (N_31924,N_30957,N_30675);
xor U31925 (N_31925,N_30925,N_30997);
nand U31926 (N_31926,N_30159,N_30944);
nand U31927 (N_31927,N_30767,N_30018);
or U31928 (N_31928,N_30939,N_30351);
or U31929 (N_31929,N_30864,N_30968);
nand U31930 (N_31930,N_30450,N_30781);
and U31931 (N_31931,N_30006,N_30625);
xor U31932 (N_31932,N_30239,N_30883);
xnor U31933 (N_31933,N_30681,N_30234);
or U31934 (N_31934,N_30511,N_30370);
nor U31935 (N_31935,N_30652,N_30242);
and U31936 (N_31936,N_30347,N_30049);
nand U31937 (N_31937,N_30302,N_30389);
or U31938 (N_31938,N_30317,N_30435);
xor U31939 (N_31939,N_30531,N_30132);
xnor U31940 (N_31940,N_30649,N_30884);
and U31941 (N_31941,N_30425,N_30490);
nor U31942 (N_31942,N_30964,N_30307);
nor U31943 (N_31943,N_30816,N_30991);
nand U31944 (N_31944,N_30973,N_30769);
nand U31945 (N_31945,N_30105,N_30848);
nand U31946 (N_31946,N_30271,N_30895);
xor U31947 (N_31947,N_30796,N_30250);
nand U31948 (N_31948,N_30172,N_30451);
and U31949 (N_31949,N_30510,N_30347);
and U31950 (N_31950,N_30948,N_30615);
nand U31951 (N_31951,N_30386,N_30532);
xnor U31952 (N_31952,N_30374,N_30169);
xnor U31953 (N_31953,N_30007,N_30995);
xnor U31954 (N_31954,N_30855,N_30078);
nor U31955 (N_31955,N_30446,N_30693);
or U31956 (N_31956,N_30308,N_30499);
xor U31957 (N_31957,N_30282,N_30033);
nand U31958 (N_31958,N_30324,N_30311);
and U31959 (N_31959,N_30138,N_30292);
xnor U31960 (N_31960,N_30897,N_30402);
nor U31961 (N_31961,N_30602,N_30538);
and U31962 (N_31962,N_30803,N_30714);
or U31963 (N_31963,N_30545,N_30480);
nand U31964 (N_31964,N_30208,N_30872);
and U31965 (N_31965,N_30710,N_30829);
nor U31966 (N_31966,N_30518,N_30847);
nand U31967 (N_31967,N_30327,N_30001);
or U31968 (N_31968,N_30744,N_30326);
nor U31969 (N_31969,N_30640,N_30515);
or U31970 (N_31970,N_30582,N_30497);
or U31971 (N_31971,N_30451,N_30111);
or U31972 (N_31972,N_30303,N_30394);
or U31973 (N_31973,N_30879,N_30950);
nor U31974 (N_31974,N_30252,N_30273);
nand U31975 (N_31975,N_30139,N_30163);
nand U31976 (N_31976,N_30487,N_30223);
or U31977 (N_31977,N_30741,N_30735);
nand U31978 (N_31978,N_30444,N_30704);
xor U31979 (N_31979,N_30526,N_30677);
nand U31980 (N_31980,N_30187,N_30359);
and U31981 (N_31981,N_30523,N_30742);
and U31982 (N_31982,N_30608,N_30314);
and U31983 (N_31983,N_30594,N_30702);
xnor U31984 (N_31984,N_30974,N_30120);
nor U31985 (N_31985,N_30956,N_30972);
nor U31986 (N_31986,N_30104,N_30665);
nor U31987 (N_31987,N_30620,N_30262);
nor U31988 (N_31988,N_30841,N_30402);
xnor U31989 (N_31989,N_30818,N_30406);
nand U31990 (N_31990,N_30058,N_30242);
xor U31991 (N_31991,N_30138,N_30818);
or U31992 (N_31992,N_30875,N_30300);
xnor U31993 (N_31993,N_30676,N_30370);
and U31994 (N_31994,N_30420,N_30688);
nand U31995 (N_31995,N_30729,N_30763);
and U31996 (N_31996,N_30910,N_30588);
and U31997 (N_31997,N_30601,N_30267);
nand U31998 (N_31998,N_30725,N_30005);
xnor U31999 (N_31999,N_30262,N_30250);
and U32000 (N_32000,N_31070,N_31489);
nor U32001 (N_32001,N_31916,N_31439);
or U32002 (N_32002,N_31761,N_31780);
xnor U32003 (N_32003,N_31305,N_31948);
or U32004 (N_32004,N_31859,N_31038);
nor U32005 (N_32005,N_31694,N_31179);
xnor U32006 (N_32006,N_31455,N_31901);
and U32007 (N_32007,N_31639,N_31704);
nand U32008 (N_32008,N_31309,N_31363);
nor U32009 (N_32009,N_31827,N_31477);
and U32010 (N_32010,N_31880,N_31036);
nor U32011 (N_32011,N_31722,N_31004);
and U32012 (N_32012,N_31401,N_31096);
and U32013 (N_32013,N_31529,N_31003);
xnor U32014 (N_32014,N_31440,N_31119);
nand U32015 (N_32015,N_31760,N_31559);
nor U32016 (N_32016,N_31166,N_31613);
nand U32017 (N_32017,N_31875,N_31226);
or U32018 (N_32018,N_31131,N_31876);
or U32019 (N_32019,N_31350,N_31207);
nand U32020 (N_32020,N_31777,N_31246);
nand U32021 (N_32021,N_31746,N_31375);
nand U32022 (N_32022,N_31597,N_31755);
xor U32023 (N_32023,N_31532,N_31826);
and U32024 (N_32024,N_31302,N_31648);
xor U32025 (N_32025,N_31514,N_31173);
nand U32026 (N_32026,N_31900,N_31194);
nand U32027 (N_32027,N_31998,N_31579);
xnor U32028 (N_32028,N_31595,N_31729);
nand U32029 (N_32029,N_31797,N_31787);
nor U32030 (N_32030,N_31599,N_31376);
nand U32031 (N_32031,N_31971,N_31655);
nand U32032 (N_32032,N_31300,N_31565);
nand U32033 (N_32033,N_31237,N_31621);
and U32034 (N_32034,N_31978,N_31877);
xor U32035 (N_32035,N_31538,N_31594);
and U32036 (N_32036,N_31351,N_31750);
or U32037 (N_32037,N_31804,N_31645);
and U32038 (N_32038,N_31820,N_31806);
nand U32039 (N_32039,N_31123,N_31284);
or U32040 (N_32040,N_31537,N_31148);
nor U32041 (N_32041,N_31331,N_31835);
nand U32042 (N_32042,N_31719,N_31083);
xnor U32043 (N_32043,N_31470,N_31261);
nor U32044 (N_32044,N_31685,N_31551);
nor U32045 (N_32045,N_31362,N_31915);
and U32046 (N_32046,N_31651,N_31442);
nand U32047 (N_32047,N_31019,N_31423);
or U32048 (N_32048,N_31609,N_31979);
or U32049 (N_32049,N_31385,N_31243);
nor U32050 (N_32050,N_31073,N_31566);
nand U32051 (N_32051,N_31554,N_31333);
nand U32052 (N_32052,N_31451,N_31002);
nand U32053 (N_32053,N_31549,N_31850);
and U32054 (N_32054,N_31980,N_31910);
nand U32055 (N_32055,N_31136,N_31710);
nand U32056 (N_32056,N_31545,N_31782);
and U32057 (N_32057,N_31281,N_31151);
nand U32058 (N_32058,N_31367,N_31593);
or U32059 (N_32059,N_31318,N_31052);
or U32060 (N_32060,N_31010,N_31196);
and U32061 (N_32061,N_31964,N_31487);
nand U32062 (N_32062,N_31042,N_31301);
or U32063 (N_32063,N_31713,N_31637);
or U32064 (N_32064,N_31057,N_31034);
nor U32065 (N_32065,N_31898,N_31178);
nor U32066 (N_32066,N_31149,N_31156);
nor U32067 (N_32067,N_31033,N_31563);
xor U32068 (N_32068,N_31252,N_31622);
or U32069 (N_32069,N_31348,N_31795);
or U32070 (N_32070,N_31502,N_31773);
xor U32071 (N_32071,N_31814,N_31957);
or U32072 (N_32072,N_31186,N_31408);
and U32073 (N_32073,N_31051,N_31976);
nor U32074 (N_32074,N_31672,N_31221);
nand U32075 (N_32075,N_31698,N_31330);
nand U32076 (N_32076,N_31654,N_31749);
or U32077 (N_32077,N_31743,N_31521);
nor U32078 (N_32078,N_31108,N_31269);
and U32079 (N_32079,N_31839,N_31786);
and U32080 (N_32080,N_31724,N_31426);
nor U32081 (N_32081,N_31356,N_31906);
nand U32082 (N_32082,N_31265,N_31630);
xor U32083 (N_32083,N_31693,N_31050);
xnor U32084 (N_32084,N_31282,N_31918);
xor U32085 (N_32085,N_31843,N_31093);
xnor U32086 (N_32086,N_31696,N_31168);
xnor U32087 (N_32087,N_31295,N_31646);
or U32088 (N_32088,N_31319,N_31954);
and U32089 (N_32089,N_31378,N_31241);
or U32090 (N_32090,N_31857,N_31412);
or U32091 (N_32091,N_31361,N_31965);
or U32092 (N_32092,N_31347,N_31960);
nor U32093 (N_32093,N_31867,N_31837);
xor U32094 (N_32094,N_31799,N_31636);
or U32095 (N_32095,N_31175,N_31270);
or U32096 (N_32096,N_31303,N_31862);
nand U32097 (N_32097,N_31009,N_31882);
nand U32098 (N_32098,N_31045,N_31308);
nand U32099 (N_32099,N_31046,N_31417);
and U32100 (N_32100,N_31572,N_31774);
nor U32101 (N_32101,N_31267,N_31222);
or U32102 (N_32102,N_31851,N_31526);
nand U32103 (N_32103,N_31977,N_31808);
xor U32104 (N_32104,N_31399,N_31500);
nor U32105 (N_32105,N_31776,N_31001);
nand U32106 (N_32106,N_31642,N_31829);
xnor U32107 (N_32107,N_31856,N_31955);
nor U32108 (N_32108,N_31200,N_31381);
or U32109 (N_32109,N_31137,N_31264);
xnor U32110 (N_32110,N_31533,N_31111);
xor U32111 (N_32111,N_31199,N_31943);
or U32112 (N_32112,N_31371,N_31732);
xor U32113 (N_32113,N_31225,N_31629);
nor U32114 (N_32114,N_31031,N_31480);
or U32115 (N_32115,N_31436,N_31778);
or U32116 (N_32116,N_31763,N_31388);
nand U32117 (N_32117,N_31012,N_31546);
or U32118 (N_32118,N_31063,N_31678);
nand U32119 (N_32119,N_31280,N_31247);
nand U32120 (N_32120,N_31803,N_31848);
nand U32121 (N_32121,N_31996,N_31967);
nand U32122 (N_32122,N_31790,N_31326);
nand U32123 (N_32123,N_31372,N_31525);
nor U32124 (N_32124,N_31413,N_31499);
or U32125 (N_32125,N_31968,N_31468);
xnor U32126 (N_32126,N_31716,N_31970);
nand U32127 (N_32127,N_31531,N_31974);
and U32128 (N_32128,N_31368,N_31158);
xor U32129 (N_32129,N_31712,N_31890);
and U32130 (N_32130,N_31479,N_31140);
or U32131 (N_32131,N_31788,N_31422);
or U32132 (N_32132,N_31509,N_31129);
and U32133 (N_32133,N_31485,N_31634);
xor U32134 (N_32134,N_31335,N_31193);
nor U32135 (N_32135,N_31759,N_31201);
xor U32136 (N_32136,N_31204,N_31972);
and U32137 (N_32137,N_31752,N_31234);
nor U32138 (N_32138,N_31107,N_31170);
and U32139 (N_32139,N_31153,N_31407);
and U32140 (N_32140,N_31411,N_31410);
and U32141 (N_32141,N_31091,N_31292);
nor U32142 (N_32142,N_31902,N_31147);
and U32143 (N_32143,N_31400,N_31576);
nor U32144 (N_32144,N_31506,N_31056);
and U32145 (N_32145,N_31962,N_31619);
xor U32146 (N_32146,N_31067,N_31816);
xor U32147 (N_32147,N_31585,N_31662);
nand U32148 (N_32148,N_31739,N_31557);
or U32149 (N_32149,N_31114,N_31517);
nor U32150 (N_32150,N_31233,N_31064);
xor U32151 (N_32151,N_31891,N_31329);
xor U32152 (N_32152,N_31103,N_31727);
or U32153 (N_32153,N_31668,N_31404);
xnor U32154 (N_32154,N_31471,N_31665);
nor U32155 (N_32155,N_31128,N_31578);
nor U32156 (N_32156,N_31605,N_31275);
nand U32157 (N_32157,N_31323,N_31087);
and U32158 (N_32158,N_31187,N_31475);
and U32159 (N_32159,N_31438,N_31311);
or U32160 (N_32160,N_31986,N_31680);
and U32161 (N_32161,N_31659,N_31952);
nor U32162 (N_32162,N_31124,N_31035);
and U32163 (N_32163,N_31562,N_31903);
nand U32164 (N_32164,N_31062,N_31737);
xnor U32165 (N_32165,N_31789,N_31205);
nand U32166 (N_32166,N_31165,N_31592);
nor U32167 (N_32167,N_31598,N_31098);
or U32168 (N_32168,N_31109,N_31897);
xor U32169 (N_32169,N_31567,N_31105);
and U32170 (N_32170,N_31516,N_31540);
nand U32171 (N_32171,N_31337,N_31374);
nand U32172 (N_32172,N_31238,N_31547);
nor U32173 (N_32173,N_31853,N_31306);
nor U32174 (N_32174,N_31380,N_31709);
nor U32175 (N_32175,N_31415,N_31245);
nor U32176 (N_32176,N_31458,N_31092);
nor U32177 (N_32177,N_31060,N_31766);
and U32178 (N_32178,N_31771,N_31044);
nor U32179 (N_32179,N_31811,N_31365);
nand U32180 (N_32180,N_31478,N_31581);
or U32181 (N_32181,N_31821,N_31048);
or U32182 (N_32182,N_31498,N_31825);
nor U32183 (N_32183,N_31818,N_31617);
xnor U32184 (N_32184,N_31913,N_31633);
nand U32185 (N_32185,N_31728,N_31176);
and U32186 (N_32186,N_31679,N_31503);
nor U32187 (N_32187,N_31707,N_31346);
xnor U32188 (N_32188,N_31874,N_31892);
or U32189 (N_32189,N_31390,N_31208);
xnor U32190 (N_32190,N_31961,N_31030);
and U32191 (N_32191,N_31435,N_31932);
nand U32192 (N_32192,N_31753,N_31177);
nand U32193 (N_32193,N_31911,N_31941);
or U32194 (N_32194,N_31250,N_31150);
xnor U32195 (N_32195,N_31386,N_31936);
xnor U32196 (N_32196,N_31467,N_31523);
or U32197 (N_32197,N_31686,N_31614);
nor U32198 (N_32198,N_31834,N_31039);
nor U32199 (N_32199,N_31740,N_31772);
nor U32200 (N_32200,N_31784,N_31588);
xnor U32201 (N_32201,N_31658,N_31992);
nor U32202 (N_32202,N_31403,N_31026);
and U32203 (N_32203,N_31344,N_31883);
or U32204 (N_32204,N_31249,N_31449);
nor U32205 (N_32205,N_31975,N_31623);
and U32206 (N_32206,N_31494,N_31914);
nor U32207 (N_32207,N_31930,N_31603);
xor U32208 (N_32208,N_31457,N_31764);
or U32209 (N_32209,N_31765,N_31625);
nor U32210 (N_32210,N_31230,N_31555);
and U32211 (N_32211,N_31813,N_31474);
nand U32212 (N_32212,N_31299,N_31022);
xnor U32213 (N_32213,N_31610,N_31711);
or U32214 (N_32214,N_31626,N_31076);
and U32215 (N_32215,N_31917,N_31574);
xor U32216 (N_32216,N_31453,N_31184);
or U32217 (N_32217,N_31181,N_31987);
nand U32218 (N_32218,N_31058,N_31973);
nand U32219 (N_32219,N_31700,N_31121);
nand U32220 (N_32220,N_31798,N_31419);
or U32221 (N_32221,N_31154,N_31486);
nor U32222 (N_32222,N_31869,N_31312);
and U32223 (N_32223,N_31416,N_31427);
xnor U32224 (N_32224,N_31615,N_31815);
or U32225 (N_32225,N_31653,N_31879);
nand U32226 (N_32226,N_31216,N_31699);
or U32227 (N_32227,N_31783,N_31522);
or U32228 (N_32228,N_31520,N_31735);
nor U32229 (N_32229,N_31504,N_31756);
nor U32230 (N_32230,N_31604,N_31667);
or U32231 (N_32231,N_31242,N_31608);
xor U32232 (N_32232,N_31054,N_31473);
nor U32233 (N_32233,N_31370,N_31643);
nand U32234 (N_32234,N_31469,N_31259);
nand U32235 (N_32235,N_31355,N_31963);
and U32236 (N_32236,N_31923,N_31999);
xnor U32237 (N_32237,N_31369,N_31988);
or U32238 (N_32238,N_31432,N_31223);
xor U32239 (N_32239,N_31144,N_31511);
xor U32240 (N_32240,N_31908,N_31845);
or U32241 (N_32241,N_31985,N_31842);
nor U32242 (N_32242,N_31501,N_31738);
nand U32243 (N_32243,N_31320,N_31840);
nand U32244 (N_32244,N_31767,N_31327);
and U32245 (N_32245,N_31692,N_31113);
or U32246 (N_32246,N_31213,N_31674);
nor U32247 (N_32247,N_31733,N_31420);
nand U32248 (N_32248,N_31425,N_31159);
xor U32249 (N_32249,N_31138,N_31907);
or U32250 (N_32250,N_31656,N_31552);
or U32251 (N_32251,N_31582,N_31112);
nor U32252 (N_32252,N_31933,N_31244);
and U32253 (N_32253,N_31239,N_31338);
xnor U32254 (N_32254,N_31530,N_31807);
nor U32255 (N_32255,N_31887,N_31452);
or U32256 (N_32256,N_31990,N_31488);
or U32257 (N_32257,N_31518,N_31627);
nand U32258 (N_32258,N_31612,N_31997);
nand U32259 (N_32259,N_31336,N_31444);
xnor U32260 (N_32260,N_31705,N_31454);
nand U32261 (N_32261,N_31189,N_31548);
and U32262 (N_32262,N_31027,N_31995);
or U32263 (N_32263,N_31029,N_31324);
or U32264 (N_32264,N_31736,N_31926);
xnor U32265 (N_32265,N_31198,N_31663);
xnor U32266 (N_32266,N_31586,N_31854);
and U32267 (N_32267,N_31947,N_31424);
or U32268 (N_32268,N_31535,N_31919);
or U32269 (N_32269,N_31993,N_31228);
nand U32270 (N_32270,N_31888,N_31358);
and U32271 (N_32271,N_31490,N_31456);
nor U32272 (N_32272,N_31157,N_31934);
xor U32273 (N_32273,N_31695,N_31065);
and U32274 (N_32274,N_31041,N_31102);
or U32275 (N_32275,N_31345,N_31717);
nor U32276 (N_32276,N_31448,N_31215);
or U32277 (N_32277,N_31644,N_31602);
nand U32278 (N_32278,N_31421,N_31145);
nor U32279 (N_32279,N_31071,N_31895);
nor U32280 (N_32280,N_31254,N_31379);
nor U32281 (N_32281,N_31018,N_31081);
and U32282 (N_32282,N_31013,N_31794);
or U32283 (N_32283,N_31163,N_31687);
and U32284 (N_32284,N_31288,N_31681);
or U32285 (N_32285,N_31409,N_31550);
nor U32286 (N_32286,N_31074,N_31394);
nand U32287 (N_32287,N_31864,N_31796);
or U32288 (N_32288,N_31231,N_31573);
and U32289 (N_32289,N_31191,N_31089);
or U32290 (N_32290,N_31758,N_31638);
or U32291 (N_32291,N_31949,N_31274);
nor U32292 (N_32292,N_31095,N_31289);
nor U32293 (N_32293,N_31536,N_31053);
and U32294 (N_32294,N_31757,N_31446);
or U32295 (N_32295,N_31349,N_31684);
xnor U32296 (N_32296,N_31310,N_31236);
nor U32297 (N_32297,N_31190,N_31754);
and U32298 (N_32298,N_31387,N_31428);
and U32299 (N_32299,N_31868,N_31258);
or U32300 (N_32300,N_31953,N_31037);
or U32301 (N_32301,N_31162,N_31366);
nand U32302 (N_32302,N_31675,N_31904);
nand U32303 (N_32303,N_31217,N_31496);
or U32304 (N_32304,N_31211,N_31575);
xor U32305 (N_32305,N_31384,N_31110);
nand U32306 (N_32306,N_31748,N_31775);
or U32307 (N_32307,N_31855,N_31544);
nand U32308 (N_32308,N_31618,N_31115);
or U32309 (N_32309,N_31650,N_31541);
and U32310 (N_32310,N_31912,N_31689);
nand U32311 (N_32311,N_31133,N_31169);
nand U32312 (N_32312,N_31209,N_31688);
and U32313 (N_32313,N_31515,N_31606);
nor U32314 (N_32314,N_31182,N_31460);
xnor U32315 (N_32315,N_31800,N_31463);
nor U32316 (N_32316,N_31072,N_31430);
and U32317 (N_32317,N_31373,N_31769);
xor U32318 (N_32318,N_31106,N_31703);
nand U32319 (N_32319,N_31382,N_31647);
xor U32320 (N_32320,N_31059,N_31127);
nor U32321 (N_32321,N_31313,N_31929);
nor U32322 (N_32322,N_31669,N_31793);
and U32323 (N_32323,N_31398,N_31383);
xor U32324 (N_32324,N_31744,N_31583);
nand U32325 (N_32325,N_31043,N_31801);
xnor U32326 (N_32326,N_31878,N_31564);
and U32327 (N_32327,N_31212,N_31090);
or U32328 (N_32328,N_31008,N_31871);
and U32329 (N_32329,N_31286,N_31360);
xnor U32330 (N_32330,N_31982,N_31852);
nand U32331 (N_32331,N_31276,N_31377);
and U32332 (N_32332,N_31075,N_31886);
or U32333 (N_32333,N_31884,N_31393);
nor U32334 (N_32334,N_31991,N_31364);
nand U32335 (N_32335,N_31924,N_31958);
nor U32336 (N_32336,N_31339,N_31134);
nor U32337 (N_32337,N_31005,N_31616);
nand U32338 (N_32338,N_31745,N_31484);
or U32339 (N_32339,N_31392,N_31872);
or U32340 (N_32340,N_31863,N_31465);
or U32341 (N_32341,N_31495,N_31751);
nand U32342 (N_32342,N_31402,N_31905);
xor U32343 (N_32343,N_31120,N_31160);
and U32344 (N_32344,N_31922,N_31691);
and U32345 (N_32345,N_31192,N_31861);
or U32346 (N_32346,N_31251,N_31741);
nor U32347 (N_32347,N_31047,N_31406);
nor U32348 (N_32348,N_31589,N_31321);
nor U32349 (N_32349,N_31255,N_31040);
nand U32350 (N_32350,N_31011,N_31632);
and U32351 (N_32351,N_31701,N_31202);
and U32352 (N_32352,N_31220,N_31352);
or U32353 (N_32353,N_31690,N_31984);
nor U32354 (N_32354,N_31085,N_31620);
and U32355 (N_32355,N_31257,N_31726);
and U32356 (N_32356,N_31519,N_31718);
and U32357 (N_32357,N_31611,N_31141);
xor U32358 (N_32358,N_31206,N_31260);
nand U32359 (N_32359,N_31328,N_31395);
nand U32360 (N_32360,N_31024,N_31556);
xnor U32361 (N_32361,N_31505,N_31000);
or U32362 (N_32362,N_31833,N_31527);
xnor U32363 (N_32363,N_31940,N_31088);
nand U32364 (N_32364,N_31015,N_31715);
nand U32365 (N_32365,N_31277,N_31860);
xnor U32366 (N_32366,N_31673,N_31077);
or U32367 (N_32367,N_31812,N_31683);
nand U32368 (N_32368,N_31253,N_31791);
xnor U32369 (N_32369,N_31293,N_31441);
nor U32370 (N_32370,N_31285,N_31635);
or U32371 (N_32371,N_31294,N_31023);
nand U32372 (N_32372,N_31482,N_31894);
nor U32373 (N_32373,N_31342,N_31291);
xnor U32374 (N_32374,N_31100,N_31459);
xor U32375 (N_32375,N_31779,N_31104);
and U32376 (N_32376,N_31762,N_31101);
nor U32377 (N_32377,N_31725,N_31132);
nor U32378 (N_32378,N_31849,N_31570);
nand U32379 (N_32379,N_31126,N_31055);
nor U32380 (N_32380,N_31560,N_31601);
nor U32381 (N_32381,N_31889,N_31049);
and U32382 (N_32382,N_31823,N_31476);
nand U32383 (N_32383,N_31297,N_31677);
nor U32384 (N_32384,N_31510,N_31927);
or U32385 (N_32385,N_31817,N_31097);
nand U32386 (N_32386,N_31099,N_31893);
nor U32387 (N_32387,N_31227,N_31641);
xnor U32388 (N_32388,N_31028,N_31171);
or U32389 (N_32389,N_31079,N_31624);
or U32390 (N_32390,N_31706,N_31657);
nand U32391 (N_32391,N_31844,N_31481);
nand U32392 (N_32392,N_31587,N_31483);
or U32393 (N_32393,N_31032,N_31188);
nand U32394 (N_32394,N_31433,N_31956);
nand U32395 (N_32395,N_31836,N_31969);
xor U32396 (N_32396,N_31240,N_31865);
xor U32397 (N_32397,N_31304,N_31183);
or U32398 (N_32398,N_31224,N_31290);
nand U32399 (N_32399,N_31061,N_31938);
nand U32400 (N_32400,N_31273,N_31946);
or U32401 (N_32401,N_31661,N_31822);
nor U32402 (N_32402,N_31828,N_31322);
xnor U32403 (N_32403,N_31069,N_31571);
or U32404 (N_32404,N_31135,N_31450);
and U32405 (N_32405,N_31298,N_31405);
or U32406 (N_32406,N_31287,N_31870);
xor U32407 (N_32407,N_31508,N_31832);
nor U32408 (N_32408,N_31078,N_31130);
and U32409 (N_32409,N_31434,N_31939);
nand U32410 (N_32410,N_31266,N_31966);
xnor U32411 (N_32411,N_31640,N_31590);
nand U32412 (N_32412,N_31841,N_31279);
nand U32413 (N_32413,N_31283,N_31730);
and U32414 (N_32414,N_31944,N_31017);
nand U32415 (N_32415,N_31125,N_31343);
and U32416 (N_32416,N_31180,N_31676);
nand U32417 (N_32417,N_31447,N_31080);
nor U32418 (N_32418,N_31117,N_31950);
nand U32419 (N_32419,N_31553,N_31942);
nor U32420 (N_32420,N_31466,N_31307);
or U32421 (N_32421,N_31146,N_31768);
nand U32422 (N_32422,N_31278,N_31866);
xnor U32423 (N_32423,N_31805,N_31397);
and U32424 (N_32424,N_31445,N_31210);
and U32425 (N_32425,N_31528,N_31920);
or U32426 (N_32426,N_31219,N_31139);
nand U32427 (N_32427,N_31316,N_31981);
nand U32428 (N_32428,N_31086,N_31167);
xor U32429 (N_32429,N_31607,N_31195);
or U32430 (N_32430,N_31831,N_31025);
and U32431 (N_32431,N_31389,N_31649);
and U32432 (N_32432,N_31568,N_31007);
or U32433 (N_32433,N_31983,N_31155);
and U32434 (N_32434,N_31512,N_31315);
nor U32435 (N_32435,N_31340,N_31164);
nor U32436 (N_32436,N_31357,N_31858);
and U32437 (N_32437,N_31491,N_31172);
xor U32438 (N_32438,N_31271,N_31909);
nand U32439 (N_32439,N_31142,N_31185);
or U32440 (N_32440,N_31885,N_31359);
nor U32441 (N_32441,N_31232,N_31561);
and U32442 (N_32442,N_31558,N_31174);
nand U32443 (N_32443,N_31731,N_31945);
xnor U32444 (N_32444,N_31770,N_31596);
nand U32445 (N_32445,N_31994,N_31122);
nand U32446 (N_32446,N_31666,N_31896);
or U32447 (N_32447,N_31116,N_31016);
xor U32448 (N_32448,N_31391,N_31396);
or U32449 (N_32449,N_31702,N_31660);
and U32450 (N_32450,N_31810,N_31152);
xnor U32451 (N_32451,N_31235,N_31325);
or U32452 (N_32452,N_31317,N_31203);
xnor U32453 (N_32453,N_31682,N_31792);
xor U32454 (N_32454,N_31584,N_31937);
nor U32455 (N_32455,N_31118,N_31899);
or U32456 (N_32456,N_31925,N_31747);
and U32457 (N_32457,N_31989,N_31781);
or U32458 (N_32458,N_31951,N_31577);
xnor U32459 (N_32459,N_31268,N_31472);
nor U32460 (N_32460,N_31020,N_31262);
or U32461 (N_32461,N_31492,N_31734);
nand U32462 (N_32462,N_31631,N_31873);
nor U32463 (N_32463,N_31539,N_31341);
nand U32464 (N_32464,N_31809,N_31229);
xor U32465 (N_32465,N_31524,N_31824);
nor U32466 (N_32466,N_31464,N_31670);
xnor U32467 (N_32467,N_31014,N_31600);
and U32468 (N_32468,N_31664,N_31143);
nor U32469 (N_32469,N_31819,N_31720);
and U32470 (N_32470,N_31543,N_31256);
xor U32471 (N_32471,N_31332,N_31742);
nor U32472 (N_32472,N_31006,N_31785);
nor U32473 (N_32473,N_31353,N_31921);
xnor U32474 (N_32474,N_31714,N_31721);
and U32475 (N_32475,N_31697,N_31263);
and U32476 (N_32476,N_31272,N_31429);
nand U32477 (N_32477,N_31161,N_31354);
and U32478 (N_32478,N_31959,N_31628);
nand U32479 (N_32479,N_31542,N_31847);
nor U32480 (N_32480,N_31493,N_31437);
or U32481 (N_32481,N_31443,N_31094);
nand U32482 (N_32482,N_31068,N_31431);
xnor U32483 (N_32483,N_31334,N_31928);
or U32484 (N_32484,N_31084,N_31802);
nor U32485 (N_32485,N_31534,N_31708);
or U32486 (N_32486,N_31569,N_31507);
xor U32487 (N_32487,N_31462,N_31418);
nand U32488 (N_32488,N_31935,N_31838);
xor U32489 (N_32489,N_31671,N_31214);
and U32490 (N_32490,N_31218,N_31197);
and U32491 (N_32491,N_31846,N_31497);
xor U32492 (N_32492,N_31248,N_31931);
or U32493 (N_32493,N_31513,N_31881);
or U32494 (N_32494,N_31066,N_31414);
nand U32495 (N_32495,N_31314,N_31296);
and U32496 (N_32496,N_31652,N_31580);
nand U32497 (N_32497,N_31723,N_31830);
and U32498 (N_32498,N_31082,N_31021);
xnor U32499 (N_32499,N_31461,N_31591);
and U32500 (N_32500,N_31432,N_31031);
nand U32501 (N_32501,N_31748,N_31489);
nand U32502 (N_32502,N_31794,N_31545);
and U32503 (N_32503,N_31414,N_31231);
and U32504 (N_32504,N_31058,N_31149);
and U32505 (N_32505,N_31520,N_31287);
xor U32506 (N_32506,N_31060,N_31351);
xor U32507 (N_32507,N_31014,N_31394);
and U32508 (N_32508,N_31884,N_31550);
nand U32509 (N_32509,N_31185,N_31886);
nand U32510 (N_32510,N_31913,N_31415);
xor U32511 (N_32511,N_31268,N_31193);
xnor U32512 (N_32512,N_31268,N_31187);
or U32513 (N_32513,N_31055,N_31940);
xnor U32514 (N_32514,N_31159,N_31527);
or U32515 (N_32515,N_31262,N_31353);
nand U32516 (N_32516,N_31363,N_31531);
nand U32517 (N_32517,N_31918,N_31448);
xor U32518 (N_32518,N_31493,N_31389);
xor U32519 (N_32519,N_31627,N_31084);
or U32520 (N_32520,N_31159,N_31174);
nand U32521 (N_32521,N_31935,N_31395);
and U32522 (N_32522,N_31717,N_31865);
nor U32523 (N_32523,N_31538,N_31123);
and U32524 (N_32524,N_31588,N_31187);
xnor U32525 (N_32525,N_31100,N_31058);
and U32526 (N_32526,N_31550,N_31596);
nand U32527 (N_32527,N_31406,N_31416);
and U32528 (N_32528,N_31704,N_31750);
or U32529 (N_32529,N_31512,N_31283);
nand U32530 (N_32530,N_31120,N_31951);
xor U32531 (N_32531,N_31382,N_31202);
or U32532 (N_32532,N_31967,N_31021);
or U32533 (N_32533,N_31556,N_31686);
or U32534 (N_32534,N_31724,N_31551);
or U32535 (N_32535,N_31673,N_31274);
or U32536 (N_32536,N_31722,N_31892);
nand U32537 (N_32537,N_31288,N_31103);
xor U32538 (N_32538,N_31363,N_31889);
xor U32539 (N_32539,N_31146,N_31569);
nand U32540 (N_32540,N_31825,N_31455);
nand U32541 (N_32541,N_31754,N_31210);
nor U32542 (N_32542,N_31246,N_31966);
xor U32543 (N_32543,N_31361,N_31288);
xor U32544 (N_32544,N_31096,N_31730);
nor U32545 (N_32545,N_31644,N_31893);
nand U32546 (N_32546,N_31482,N_31717);
xnor U32547 (N_32547,N_31798,N_31420);
and U32548 (N_32548,N_31341,N_31177);
xnor U32549 (N_32549,N_31445,N_31076);
nand U32550 (N_32550,N_31127,N_31472);
and U32551 (N_32551,N_31084,N_31651);
nor U32552 (N_32552,N_31774,N_31126);
and U32553 (N_32553,N_31714,N_31356);
nand U32554 (N_32554,N_31339,N_31018);
xnor U32555 (N_32555,N_31542,N_31830);
nand U32556 (N_32556,N_31299,N_31556);
and U32557 (N_32557,N_31366,N_31406);
or U32558 (N_32558,N_31403,N_31381);
nor U32559 (N_32559,N_31445,N_31270);
and U32560 (N_32560,N_31414,N_31757);
nor U32561 (N_32561,N_31069,N_31227);
nor U32562 (N_32562,N_31051,N_31364);
and U32563 (N_32563,N_31508,N_31352);
or U32564 (N_32564,N_31658,N_31274);
or U32565 (N_32565,N_31329,N_31508);
xor U32566 (N_32566,N_31096,N_31382);
or U32567 (N_32567,N_31469,N_31992);
nand U32568 (N_32568,N_31556,N_31984);
or U32569 (N_32569,N_31690,N_31049);
nor U32570 (N_32570,N_31947,N_31989);
nand U32571 (N_32571,N_31481,N_31257);
xnor U32572 (N_32572,N_31650,N_31774);
and U32573 (N_32573,N_31275,N_31122);
xnor U32574 (N_32574,N_31021,N_31232);
nand U32575 (N_32575,N_31880,N_31446);
and U32576 (N_32576,N_31447,N_31992);
or U32577 (N_32577,N_31745,N_31464);
and U32578 (N_32578,N_31232,N_31894);
xnor U32579 (N_32579,N_31593,N_31414);
nand U32580 (N_32580,N_31159,N_31553);
or U32581 (N_32581,N_31131,N_31656);
or U32582 (N_32582,N_31382,N_31170);
and U32583 (N_32583,N_31526,N_31240);
nand U32584 (N_32584,N_31504,N_31921);
nand U32585 (N_32585,N_31228,N_31234);
nand U32586 (N_32586,N_31369,N_31696);
nand U32587 (N_32587,N_31123,N_31586);
and U32588 (N_32588,N_31457,N_31164);
xor U32589 (N_32589,N_31402,N_31339);
xnor U32590 (N_32590,N_31192,N_31450);
nor U32591 (N_32591,N_31817,N_31393);
xor U32592 (N_32592,N_31725,N_31070);
xnor U32593 (N_32593,N_31346,N_31833);
nor U32594 (N_32594,N_31640,N_31756);
or U32595 (N_32595,N_31684,N_31366);
nor U32596 (N_32596,N_31819,N_31420);
or U32597 (N_32597,N_31413,N_31246);
nor U32598 (N_32598,N_31768,N_31502);
nor U32599 (N_32599,N_31614,N_31239);
xnor U32600 (N_32600,N_31489,N_31207);
nor U32601 (N_32601,N_31836,N_31917);
nor U32602 (N_32602,N_31204,N_31739);
xnor U32603 (N_32603,N_31882,N_31703);
or U32604 (N_32604,N_31586,N_31110);
nand U32605 (N_32605,N_31779,N_31797);
nand U32606 (N_32606,N_31626,N_31928);
or U32607 (N_32607,N_31302,N_31945);
xor U32608 (N_32608,N_31648,N_31558);
or U32609 (N_32609,N_31967,N_31434);
and U32610 (N_32610,N_31800,N_31022);
xnor U32611 (N_32611,N_31443,N_31021);
nand U32612 (N_32612,N_31289,N_31337);
and U32613 (N_32613,N_31267,N_31522);
and U32614 (N_32614,N_31616,N_31741);
xor U32615 (N_32615,N_31940,N_31605);
xor U32616 (N_32616,N_31775,N_31005);
or U32617 (N_32617,N_31979,N_31675);
nor U32618 (N_32618,N_31123,N_31987);
xnor U32619 (N_32619,N_31449,N_31807);
or U32620 (N_32620,N_31094,N_31038);
and U32621 (N_32621,N_31728,N_31952);
nor U32622 (N_32622,N_31745,N_31856);
or U32623 (N_32623,N_31089,N_31483);
and U32624 (N_32624,N_31301,N_31919);
and U32625 (N_32625,N_31491,N_31690);
xor U32626 (N_32626,N_31996,N_31870);
nor U32627 (N_32627,N_31044,N_31993);
nor U32628 (N_32628,N_31795,N_31960);
or U32629 (N_32629,N_31889,N_31457);
nor U32630 (N_32630,N_31364,N_31816);
nor U32631 (N_32631,N_31549,N_31951);
and U32632 (N_32632,N_31492,N_31697);
xnor U32633 (N_32633,N_31657,N_31917);
or U32634 (N_32634,N_31109,N_31689);
nand U32635 (N_32635,N_31164,N_31362);
xnor U32636 (N_32636,N_31656,N_31417);
nor U32637 (N_32637,N_31312,N_31007);
or U32638 (N_32638,N_31511,N_31160);
xnor U32639 (N_32639,N_31947,N_31868);
and U32640 (N_32640,N_31326,N_31299);
nor U32641 (N_32641,N_31039,N_31217);
nand U32642 (N_32642,N_31565,N_31333);
xor U32643 (N_32643,N_31193,N_31123);
or U32644 (N_32644,N_31594,N_31688);
nor U32645 (N_32645,N_31549,N_31464);
xor U32646 (N_32646,N_31836,N_31495);
xor U32647 (N_32647,N_31708,N_31981);
xor U32648 (N_32648,N_31656,N_31880);
xnor U32649 (N_32649,N_31262,N_31735);
or U32650 (N_32650,N_31704,N_31139);
and U32651 (N_32651,N_31849,N_31763);
or U32652 (N_32652,N_31680,N_31883);
and U32653 (N_32653,N_31614,N_31472);
and U32654 (N_32654,N_31463,N_31326);
or U32655 (N_32655,N_31562,N_31482);
or U32656 (N_32656,N_31470,N_31680);
nor U32657 (N_32657,N_31257,N_31819);
nor U32658 (N_32658,N_31120,N_31079);
and U32659 (N_32659,N_31949,N_31745);
or U32660 (N_32660,N_31562,N_31797);
or U32661 (N_32661,N_31044,N_31576);
and U32662 (N_32662,N_31771,N_31710);
nand U32663 (N_32663,N_31502,N_31229);
nand U32664 (N_32664,N_31919,N_31085);
xor U32665 (N_32665,N_31126,N_31977);
and U32666 (N_32666,N_31557,N_31524);
or U32667 (N_32667,N_31588,N_31284);
nor U32668 (N_32668,N_31500,N_31876);
nand U32669 (N_32669,N_31090,N_31169);
and U32670 (N_32670,N_31789,N_31044);
xor U32671 (N_32671,N_31509,N_31277);
and U32672 (N_32672,N_31854,N_31237);
nor U32673 (N_32673,N_31084,N_31111);
xor U32674 (N_32674,N_31905,N_31595);
xnor U32675 (N_32675,N_31002,N_31878);
and U32676 (N_32676,N_31605,N_31838);
and U32677 (N_32677,N_31068,N_31623);
nor U32678 (N_32678,N_31547,N_31876);
or U32679 (N_32679,N_31091,N_31514);
xnor U32680 (N_32680,N_31182,N_31759);
nand U32681 (N_32681,N_31709,N_31255);
nor U32682 (N_32682,N_31936,N_31024);
nand U32683 (N_32683,N_31605,N_31127);
xor U32684 (N_32684,N_31598,N_31023);
or U32685 (N_32685,N_31646,N_31064);
nor U32686 (N_32686,N_31492,N_31020);
xor U32687 (N_32687,N_31409,N_31194);
nand U32688 (N_32688,N_31410,N_31902);
or U32689 (N_32689,N_31597,N_31420);
nand U32690 (N_32690,N_31370,N_31586);
xor U32691 (N_32691,N_31199,N_31081);
xnor U32692 (N_32692,N_31772,N_31831);
nor U32693 (N_32693,N_31420,N_31415);
or U32694 (N_32694,N_31841,N_31982);
and U32695 (N_32695,N_31049,N_31094);
nand U32696 (N_32696,N_31859,N_31146);
nand U32697 (N_32697,N_31422,N_31583);
nor U32698 (N_32698,N_31550,N_31454);
or U32699 (N_32699,N_31163,N_31323);
and U32700 (N_32700,N_31380,N_31856);
nor U32701 (N_32701,N_31407,N_31541);
or U32702 (N_32702,N_31991,N_31726);
nor U32703 (N_32703,N_31510,N_31421);
or U32704 (N_32704,N_31721,N_31645);
or U32705 (N_32705,N_31025,N_31948);
xor U32706 (N_32706,N_31474,N_31705);
and U32707 (N_32707,N_31300,N_31089);
nor U32708 (N_32708,N_31395,N_31027);
or U32709 (N_32709,N_31790,N_31592);
nand U32710 (N_32710,N_31031,N_31557);
or U32711 (N_32711,N_31763,N_31112);
or U32712 (N_32712,N_31235,N_31135);
and U32713 (N_32713,N_31494,N_31230);
or U32714 (N_32714,N_31190,N_31691);
or U32715 (N_32715,N_31968,N_31999);
and U32716 (N_32716,N_31458,N_31997);
xnor U32717 (N_32717,N_31838,N_31109);
and U32718 (N_32718,N_31407,N_31943);
nor U32719 (N_32719,N_31162,N_31074);
or U32720 (N_32720,N_31906,N_31897);
nand U32721 (N_32721,N_31900,N_31599);
nor U32722 (N_32722,N_31518,N_31204);
nor U32723 (N_32723,N_31488,N_31703);
and U32724 (N_32724,N_31800,N_31728);
or U32725 (N_32725,N_31210,N_31244);
and U32726 (N_32726,N_31426,N_31867);
nand U32727 (N_32727,N_31471,N_31724);
xor U32728 (N_32728,N_31104,N_31684);
and U32729 (N_32729,N_31118,N_31145);
and U32730 (N_32730,N_31171,N_31553);
or U32731 (N_32731,N_31523,N_31485);
and U32732 (N_32732,N_31449,N_31234);
nor U32733 (N_32733,N_31257,N_31203);
xor U32734 (N_32734,N_31435,N_31956);
or U32735 (N_32735,N_31004,N_31902);
and U32736 (N_32736,N_31977,N_31204);
nand U32737 (N_32737,N_31378,N_31184);
nor U32738 (N_32738,N_31236,N_31755);
xnor U32739 (N_32739,N_31849,N_31654);
nand U32740 (N_32740,N_31438,N_31026);
and U32741 (N_32741,N_31004,N_31112);
and U32742 (N_32742,N_31846,N_31897);
nor U32743 (N_32743,N_31885,N_31871);
and U32744 (N_32744,N_31698,N_31800);
or U32745 (N_32745,N_31944,N_31611);
xnor U32746 (N_32746,N_31252,N_31986);
nand U32747 (N_32747,N_31788,N_31727);
and U32748 (N_32748,N_31310,N_31231);
xor U32749 (N_32749,N_31315,N_31526);
or U32750 (N_32750,N_31127,N_31071);
nand U32751 (N_32751,N_31098,N_31127);
or U32752 (N_32752,N_31539,N_31639);
xor U32753 (N_32753,N_31433,N_31414);
or U32754 (N_32754,N_31226,N_31073);
nor U32755 (N_32755,N_31777,N_31345);
nor U32756 (N_32756,N_31525,N_31477);
xnor U32757 (N_32757,N_31016,N_31656);
or U32758 (N_32758,N_31526,N_31117);
and U32759 (N_32759,N_31966,N_31309);
and U32760 (N_32760,N_31445,N_31305);
and U32761 (N_32761,N_31071,N_31489);
and U32762 (N_32762,N_31489,N_31284);
nor U32763 (N_32763,N_31146,N_31753);
nand U32764 (N_32764,N_31709,N_31303);
xor U32765 (N_32765,N_31532,N_31120);
or U32766 (N_32766,N_31198,N_31820);
nand U32767 (N_32767,N_31714,N_31057);
nor U32768 (N_32768,N_31273,N_31448);
and U32769 (N_32769,N_31356,N_31625);
nand U32770 (N_32770,N_31061,N_31328);
nand U32771 (N_32771,N_31487,N_31221);
nor U32772 (N_32772,N_31202,N_31169);
nor U32773 (N_32773,N_31025,N_31000);
xnor U32774 (N_32774,N_31774,N_31590);
and U32775 (N_32775,N_31510,N_31365);
nor U32776 (N_32776,N_31910,N_31432);
or U32777 (N_32777,N_31037,N_31547);
or U32778 (N_32778,N_31839,N_31926);
nor U32779 (N_32779,N_31733,N_31700);
and U32780 (N_32780,N_31688,N_31722);
or U32781 (N_32781,N_31325,N_31051);
nand U32782 (N_32782,N_31197,N_31600);
xnor U32783 (N_32783,N_31925,N_31456);
or U32784 (N_32784,N_31257,N_31235);
and U32785 (N_32785,N_31781,N_31467);
nor U32786 (N_32786,N_31893,N_31883);
and U32787 (N_32787,N_31185,N_31607);
xor U32788 (N_32788,N_31255,N_31135);
nor U32789 (N_32789,N_31859,N_31351);
xnor U32790 (N_32790,N_31130,N_31037);
and U32791 (N_32791,N_31958,N_31752);
xnor U32792 (N_32792,N_31725,N_31013);
xor U32793 (N_32793,N_31843,N_31076);
xor U32794 (N_32794,N_31225,N_31380);
nand U32795 (N_32795,N_31395,N_31029);
xor U32796 (N_32796,N_31200,N_31574);
and U32797 (N_32797,N_31627,N_31193);
and U32798 (N_32798,N_31394,N_31787);
nand U32799 (N_32799,N_31662,N_31301);
and U32800 (N_32800,N_31577,N_31903);
nand U32801 (N_32801,N_31184,N_31958);
xor U32802 (N_32802,N_31509,N_31037);
nor U32803 (N_32803,N_31150,N_31349);
nor U32804 (N_32804,N_31264,N_31804);
nand U32805 (N_32805,N_31954,N_31894);
nor U32806 (N_32806,N_31080,N_31004);
nand U32807 (N_32807,N_31148,N_31634);
xor U32808 (N_32808,N_31774,N_31429);
nor U32809 (N_32809,N_31477,N_31309);
or U32810 (N_32810,N_31393,N_31455);
nand U32811 (N_32811,N_31913,N_31733);
nor U32812 (N_32812,N_31571,N_31303);
nand U32813 (N_32813,N_31226,N_31897);
nand U32814 (N_32814,N_31495,N_31372);
nand U32815 (N_32815,N_31932,N_31569);
or U32816 (N_32816,N_31547,N_31829);
and U32817 (N_32817,N_31248,N_31542);
nand U32818 (N_32818,N_31858,N_31090);
nand U32819 (N_32819,N_31715,N_31801);
or U32820 (N_32820,N_31973,N_31662);
or U32821 (N_32821,N_31060,N_31999);
or U32822 (N_32822,N_31500,N_31823);
and U32823 (N_32823,N_31943,N_31803);
nand U32824 (N_32824,N_31766,N_31760);
and U32825 (N_32825,N_31527,N_31930);
nor U32826 (N_32826,N_31759,N_31082);
xnor U32827 (N_32827,N_31527,N_31719);
xor U32828 (N_32828,N_31397,N_31734);
or U32829 (N_32829,N_31337,N_31977);
xor U32830 (N_32830,N_31722,N_31107);
nor U32831 (N_32831,N_31798,N_31973);
nor U32832 (N_32832,N_31155,N_31391);
or U32833 (N_32833,N_31307,N_31892);
or U32834 (N_32834,N_31087,N_31859);
or U32835 (N_32835,N_31613,N_31029);
nand U32836 (N_32836,N_31072,N_31994);
nor U32837 (N_32837,N_31629,N_31535);
or U32838 (N_32838,N_31384,N_31584);
nand U32839 (N_32839,N_31465,N_31187);
xnor U32840 (N_32840,N_31079,N_31099);
xor U32841 (N_32841,N_31607,N_31653);
nor U32842 (N_32842,N_31558,N_31217);
nor U32843 (N_32843,N_31770,N_31446);
xnor U32844 (N_32844,N_31201,N_31251);
or U32845 (N_32845,N_31782,N_31818);
nand U32846 (N_32846,N_31160,N_31249);
nor U32847 (N_32847,N_31063,N_31257);
xor U32848 (N_32848,N_31501,N_31657);
or U32849 (N_32849,N_31109,N_31183);
nor U32850 (N_32850,N_31891,N_31503);
xor U32851 (N_32851,N_31343,N_31111);
xor U32852 (N_32852,N_31058,N_31863);
nand U32853 (N_32853,N_31358,N_31174);
xor U32854 (N_32854,N_31127,N_31724);
and U32855 (N_32855,N_31253,N_31709);
nor U32856 (N_32856,N_31281,N_31584);
or U32857 (N_32857,N_31477,N_31251);
nor U32858 (N_32858,N_31795,N_31141);
and U32859 (N_32859,N_31953,N_31859);
xnor U32860 (N_32860,N_31418,N_31292);
nor U32861 (N_32861,N_31169,N_31432);
nor U32862 (N_32862,N_31880,N_31196);
and U32863 (N_32863,N_31690,N_31788);
or U32864 (N_32864,N_31686,N_31867);
and U32865 (N_32865,N_31455,N_31122);
xnor U32866 (N_32866,N_31902,N_31736);
and U32867 (N_32867,N_31237,N_31123);
or U32868 (N_32868,N_31735,N_31959);
or U32869 (N_32869,N_31634,N_31102);
xnor U32870 (N_32870,N_31494,N_31125);
xor U32871 (N_32871,N_31310,N_31719);
nand U32872 (N_32872,N_31323,N_31826);
nand U32873 (N_32873,N_31177,N_31010);
and U32874 (N_32874,N_31890,N_31733);
nor U32875 (N_32875,N_31732,N_31286);
and U32876 (N_32876,N_31883,N_31828);
nor U32877 (N_32877,N_31214,N_31821);
nand U32878 (N_32878,N_31257,N_31760);
and U32879 (N_32879,N_31968,N_31092);
or U32880 (N_32880,N_31209,N_31095);
nand U32881 (N_32881,N_31571,N_31186);
nand U32882 (N_32882,N_31977,N_31023);
nand U32883 (N_32883,N_31078,N_31591);
xnor U32884 (N_32884,N_31060,N_31143);
nand U32885 (N_32885,N_31239,N_31826);
nor U32886 (N_32886,N_31185,N_31709);
nor U32887 (N_32887,N_31669,N_31176);
xnor U32888 (N_32888,N_31091,N_31114);
nor U32889 (N_32889,N_31583,N_31705);
or U32890 (N_32890,N_31332,N_31734);
or U32891 (N_32891,N_31812,N_31769);
or U32892 (N_32892,N_31263,N_31162);
and U32893 (N_32893,N_31009,N_31845);
or U32894 (N_32894,N_31076,N_31487);
nor U32895 (N_32895,N_31075,N_31235);
or U32896 (N_32896,N_31110,N_31447);
xnor U32897 (N_32897,N_31199,N_31569);
xnor U32898 (N_32898,N_31903,N_31718);
or U32899 (N_32899,N_31452,N_31830);
xnor U32900 (N_32900,N_31565,N_31068);
and U32901 (N_32901,N_31843,N_31892);
or U32902 (N_32902,N_31303,N_31581);
xor U32903 (N_32903,N_31494,N_31074);
xor U32904 (N_32904,N_31916,N_31600);
xor U32905 (N_32905,N_31199,N_31007);
nand U32906 (N_32906,N_31178,N_31020);
xor U32907 (N_32907,N_31206,N_31907);
xnor U32908 (N_32908,N_31543,N_31559);
nand U32909 (N_32909,N_31951,N_31474);
xnor U32910 (N_32910,N_31537,N_31523);
xor U32911 (N_32911,N_31313,N_31268);
or U32912 (N_32912,N_31391,N_31591);
xor U32913 (N_32913,N_31210,N_31340);
and U32914 (N_32914,N_31238,N_31887);
xnor U32915 (N_32915,N_31447,N_31902);
and U32916 (N_32916,N_31462,N_31271);
and U32917 (N_32917,N_31549,N_31887);
xnor U32918 (N_32918,N_31301,N_31181);
nor U32919 (N_32919,N_31651,N_31403);
xnor U32920 (N_32920,N_31120,N_31395);
or U32921 (N_32921,N_31654,N_31267);
or U32922 (N_32922,N_31423,N_31036);
nor U32923 (N_32923,N_31328,N_31048);
xnor U32924 (N_32924,N_31130,N_31956);
xor U32925 (N_32925,N_31788,N_31702);
nor U32926 (N_32926,N_31480,N_31015);
or U32927 (N_32927,N_31029,N_31211);
and U32928 (N_32928,N_31806,N_31935);
and U32929 (N_32929,N_31590,N_31661);
nor U32930 (N_32930,N_31547,N_31683);
nor U32931 (N_32931,N_31289,N_31805);
and U32932 (N_32932,N_31435,N_31136);
nand U32933 (N_32933,N_31159,N_31572);
and U32934 (N_32934,N_31434,N_31372);
or U32935 (N_32935,N_31840,N_31953);
nor U32936 (N_32936,N_31947,N_31906);
or U32937 (N_32937,N_31533,N_31197);
or U32938 (N_32938,N_31351,N_31617);
and U32939 (N_32939,N_31171,N_31627);
xor U32940 (N_32940,N_31794,N_31972);
and U32941 (N_32941,N_31392,N_31341);
or U32942 (N_32942,N_31573,N_31211);
or U32943 (N_32943,N_31020,N_31742);
nand U32944 (N_32944,N_31016,N_31401);
or U32945 (N_32945,N_31676,N_31825);
nand U32946 (N_32946,N_31082,N_31083);
and U32947 (N_32947,N_31505,N_31437);
or U32948 (N_32948,N_31984,N_31417);
and U32949 (N_32949,N_31731,N_31110);
xnor U32950 (N_32950,N_31530,N_31457);
xor U32951 (N_32951,N_31840,N_31820);
xnor U32952 (N_32952,N_31152,N_31071);
or U32953 (N_32953,N_31265,N_31145);
xor U32954 (N_32954,N_31241,N_31799);
nor U32955 (N_32955,N_31014,N_31341);
nand U32956 (N_32956,N_31772,N_31273);
xnor U32957 (N_32957,N_31028,N_31834);
nand U32958 (N_32958,N_31784,N_31193);
or U32959 (N_32959,N_31250,N_31950);
and U32960 (N_32960,N_31714,N_31879);
and U32961 (N_32961,N_31655,N_31576);
and U32962 (N_32962,N_31912,N_31114);
nand U32963 (N_32963,N_31705,N_31844);
nor U32964 (N_32964,N_31434,N_31842);
and U32965 (N_32965,N_31840,N_31738);
nand U32966 (N_32966,N_31409,N_31591);
nor U32967 (N_32967,N_31302,N_31528);
nor U32968 (N_32968,N_31259,N_31991);
nor U32969 (N_32969,N_31792,N_31509);
xnor U32970 (N_32970,N_31095,N_31940);
or U32971 (N_32971,N_31320,N_31816);
nor U32972 (N_32972,N_31871,N_31971);
xor U32973 (N_32973,N_31797,N_31234);
or U32974 (N_32974,N_31143,N_31848);
and U32975 (N_32975,N_31541,N_31115);
and U32976 (N_32976,N_31368,N_31195);
nor U32977 (N_32977,N_31902,N_31435);
nand U32978 (N_32978,N_31178,N_31685);
or U32979 (N_32979,N_31874,N_31057);
and U32980 (N_32980,N_31670,N_31359);
or U32981 (N_32981,N_31416,N_31645);
xor U32982 (N_32982,N_31521,N_31215);
nand U32983 (N_32983,N_31976,N_31714);
xor U32984 (N_32984,N_31558,N_31184);
and U32985 (N_32985,N_31634,N_31145);
or U32986 (N_32986,N_31342,N_31221);
or U32987 (N_32987,N_31517,N_31030);
nand U32988 (N_32988,N_31219,N_31035);
and U32989 (N_32989,N_31161,N_31626);
nand U32990 (N_32990,N_31168,N_31470);
and U32991 (N_32991,N_31481,N_31639);
nor U32992 (N_32992,N_31681,N_31616);
and U32993 (N_32993,N_31263,N_31105);
or U32994 (N_32994,N_31351,N_31336);
nand U32995 (N_32995,N_31860,N_31572);
nand U32996 (N_32996,N_31380,N_31193);
nand U32997 (N_32997,N_31525,N_31943);
and U32998 (N_32998,N_31748,N_31524);
nand U32999 (N_32999,N_31879,N_31500);
nand U33000 (N_33000,N_32765,N_32991);
nor U33001 (N_33001,N_32619,N_32156);
xor U33002 (N_33002,N_32287,N_32898);
and U33003 (N_33003,N_32075,N_32425);
nand U33004 (N_33004,N_32072,N_32048);
or U33005 (N_33005,N_32598,N_32269);
xnor U33006 (N_33006,N_32512,N_32874);
nor U33007 (N_33007,N_32664,N_32102);
or U33008 (N_33008,N_32870,N_32310);
and U33009 (N_33009,N_32777,N_32291);
and U33010 (N_33010,N_32375,N_32641);
or U33011 (N_33011,N_32669,N_32470);
xor U33012 (N_33012,N_32240,N_32423);
xnor U33013 (N_33013,N_32361,N_32886);
nand U33014 (N_33014,N_32280,N_32185);
nor U33015 (N_33015,N_32562,N_32579);
xor U33016 (N_33016,N_32553,N_32924);
xnor U33017 (N_33017,N_32289,N_32057);
or U33018 (N_33018,N_32172,N_32390);
nor U33019 (N_33019,N_32037,N_32929);
or U33020 (N_33020,N_32138,N_32322);
nand U33021 (N_33021,N_32903,N_32087);
xor U33022 (N_33022,N_32735,N_32392);
nand U33023 (N_33023,N_32752,N_32412);
xnor U33024 (N_33024,N_32521,N_32586);
nor U33025 (N_33025,N_32159,N_32200);
xor U33026 (N_33026,N_32980,N_32839);
nor U33027 (N_33027,N_32356,N_32011);
xor U33028 (N_33028,N_32443,N_32733);
nor U33029 (N_33029,N_32565,N_32342);
and U33030 (N_33030,N_32576,N_32943);
or U33031 (N_33031,N_32042,N_32056);
or U33032 (N_33032,N_32052,N_32177);
and U33033 (N_33033,N_32370,N_32064);
or U33034 (N_33034,N_32357,N_32348);
xnor U33035 (N_33035,N_32007,N_32848);
or U33036 (N_33036,N_32725,N_32999);
nor U33037 (N_33037,N_32808,N_32580);
nor U33038 (N_33038,N_32825,N_32374);
and U33039 (N_33039,N_32006,N_32000);
xor U33040 (N_33040,N_32083,N_32678);
xor U33041 (N_33041,N_32648,N_32601);
and U33042 (N_33042,N_32104,N_32414);
nor U33043 (N_33043,N_32230,N_32837);
or U33044 (N_33044,N_32549,N_32933);
xnor U33045 (N_33045,N_32749,N_32594);
nand U33046 (N_33046,N_32398,N_32629);
and U33047 (N_33047,N_32140,N_32389);
or U33048 (N_33048,N_32846,N_32306);
and U33049 (N_33049,N_32282,N_32341);
nand U33050 (N_33050,N_32950,N_32518);
and U33051 (N_33051,N_32090,N_32986);
nand U33052 (N_33052,N_32192,N_32936);
nand U33053 (N_33053,N_32712,N_32859);
nand U33054 (N_33054,N_32040,N_32570);
xnor U33055 (N_33055,N_32184,N_32440);
or U33056 (N_33056,N_32054,N_32876);
or U33057 (N_33057,N_32401,N_32106);
and U33058 (N_33058,N_32729,N_32433);
and U33059 (N_33059,N_32131,N_32290);
or U33060 (N_33060,N_32609,N_32147);
or U33061 (N_33061,N_32274,N_32315);
and U33062 (N_33062,N_32649,N_32481);
xor U33063 (N_33063,N_32365,N_32456);
xnor U33064 (N_33064,N_32119,N_32126);
nand U33065 (N_33065,N_32016,N_32703);
xnor U33066 (N_33066,N_32647,N_32221);
or U33067 (N_33067,N_32850,N_32904);
nand U33068 (N_33068,N_32421,N_32039);
and U33069 (N_33069,N_32428,N_32128);
nand U33070 (N_33070,N_32841,N_32308);
xnor U33071 (N_33071,N_32536,N_32533);
or U33072 (N_33072,N_32668,N_32127);
nor U33073 (N_33073,N_32393,N_32731);
or U33074 (N_33074,N_32275,N_32782);
nand U33075 (N_33075,N_32797,N_32860);
and U33076 (N_33076,N_32084,N_32381);
or U33077 (N_33077,N_32989,N_32100);
nand U33078 (N_33078,N_32014,N_32441);
nor U33079 (N_33079,N_32867,N_32092);
nand U33080 (N_33080,N_32820,N_32962);
nand U33081 (N_33081,N_32191,N_32169);
and U33082 (N_33082,N_32754,N_32646);
nor U33083 (N_33083,N_32852,N_32742);
nor U33084 (N_33084,N_32815,N_32208);
xnor U33085 (N_33085,N_32271,N_32511);
or U33086 (N_33086,N_32931,N_32260);
or U33087 (N_33087,N_32427,N_32717);
nand U33088 (N_33088,N_32432,N_32460);
nor U33089 (N_33089,N_32636,N_32951);
xnor U33090 (N_33090,N_32843,N_32885);
nand U33091 (N_33091,N_32327,N_32288);
or U33092 (N_33092,N_32158,N_32034);
and U33093 (N_33093,N_32363,N_32968);
nor U33094 (N_33094,N_32803,N_32910);
and U33095 (N_33095,N_32150,N_32170);
xor U33096 (N_33096,N_32482,N_32205);
xor U33097 (N_33097,N_32845,N_32495);
nand U33098 (N_33098,N_32545,N_32935);
xor U33099 (N_33099,N_32018,N_32779);
nor U33100 (N_33100,N_32701,N_32137);
nand U33101 (N_33101,N_32789,N_32771);
and U33102 (N_33102,N_32466,N_32343);
or U33103 (N_33103,N_32748,N_32584);
or U33104 (N_33104,N_32151,N_32108);
and U33105 (N_33105,N_32661,N_32746);
xor U33106 (N_33106,N_32118,N_32738);
and U33107 (N_33107,N_32004,N_32613);
nand U33108 (N_33108,N_32251,N_32892);
nand U33109 (N_33109,N_32996,N_32812);
and U33110 (N_33110,N_32409,N_32146);
and U33111 (N_33111,N_32921,N_32141);
nor U33112 (N_33112,N_32875,N_32798);
nor U33113 (N_33113,N_32133,N_32539);
or U33114 (N_33114,N_32399,N_32901);
or U33115 (N_33115,N_32659,N_32228);
or U33116 (N_33116,N_32872,N_32165);
xor U33117 (N_33117,N_32662,N_32162);
and U33118 (N_33118,N_32074,N_32956);
or U33119 (N_33119,N_32091,N_32047);
and U33120 (N_33120,N_32199,N_32344);
xor U33121 (N_33121,N_32416,N_32321);
nor U33122 (N_33122,N_32853,N_32272);
and U33123 (N_33123,N_32655,N_32088);
and U33124 (N_33124,N_32589,N_32225);
nand U33125 (N_33125,N_32086,N_32181);
xor U33126 (N_33126,N_32005,N_32773);
nand U33127 (N_33127,N_32372,N_32948);
and U33128 (N_33128,N_32216,N_32802);
xor U33129 (N_33129,N_32266,N_32385);
xnor U33130 (N_33130,N_32713,N_32605);
or U33131 (N_33131,N_32834,N_32303);
nand U33132 (N_33132,N_32050,N_32890);
nor U33133 (N_33133,N_32476,N_32621);
xnor U33134 (N_33134,N_32667,N_32194);
and U33135 (N_33135,N_32596,N_32542);
and U33136 (N_33136,N_32193,N_32821);
nor U33137 (N_33137,N_32679,N_32743);
xor U33138 (N_33138,N_32695,N_32707);
xor U33139 (N_33139,N_32334,N_32059);
or U33140 (N_33140,N_32069,N_32665);
and U33141 (N_33141,N_32350,N_32093);
or U33142 (N_33142,N_32213,N_32568);
nand U33143 (N_33143,N_32774,N_32043);
and U33144 (N_33144,N_32550,N_32012);
or U33145 (N_33145,N_32581,N_32198);
nand U33146 (N_33146,N_32279,N_32541);
nor U33147 (N_33147,N_32379,N_32492);
nor U33148 (N_33148,N_32299,N_32544);
nor U33149 (N_33149,N_32071,N_32168);
and U33150 (N_33150,N_32967,N_32257);
and U33151 (N_33151,N_32805,N_32630);
xnor U33152 (N_33152,N_32760,N_32359);
or U33153 (N_33153,N_32215,N_32858);
and U33154 (N_33154,N_32455,N_32167);
nor U33155 (N_33155,N_32281,N_32292);
and U33156 (N_33156,N_32709,N_32095);
and U33157 (N_33157,N_32196,N_32548);
and U33158 (N_33158,N_32757,N_32947);
nand U33159 (N_33159,N_32801,N_32672);
and U33160 (N_33160,N_32654,N_32937);
nand U33161 (N_33161,N_32889,N_32340);
nand U33162 (N_33162,N_32716,N_32631);
nor U33163 (N_33163,N_32608,N_32582);
or U33164 (N_33164,N_32547,N_32293);
xor U33165 (N_33165,N_32998,N_32786);
nor U33166 (N_33166,N_32276,N_32404);
nor U33167 (N_33167,N_32992,N_32391);
nor U33168 (N_33168,N_32132,N_32461);
and U33169 (N_33169,N_32189,N_32987);
xnor U33170 (N_33170,N_32690,N_32830);
and U33171 (N_33171,N_32247,N_32273);
nand U33172 (N_33172,N_32572,N_32335);
nand U33173 (N_33173,N_32974,N_32496);
nand U33174 (N_33174,N_32239,N_32448);
and U33175 (N_33175,N_32526,N_32491);
and U33176 (N_33176,N_32096,N_32683);
or U33177 (N_33177,N_32978,N_32229);
or U33178 (N_33178,N_32109,N_32810);
or U33179 (N_33179,N_32587,N_32866);
and U33180 (N_33180,N_32174,N_32122);
nand U33181 (N_33181,N_32231,N_32278);
xor U33182 (N_33182,N_32979,N_32559);
nor U33183 (N_33183,N_32130,N_32957);
nand U33184 (N_33184,N_32032,N_32333);
and U33185 (N_33185,N_32178,N_32499);
xnor U33186 (N_33186,N_32224,N_32796);
and U33187 (N_33187,N_32915,N_32573);
and U33188 (N_33188,N_32793,N_32599);
and U33189 (N_33189,N_32975,N_32489);
and U33190 (N_33190,N_32684,N_32855);
or U33191 (N_33191,N_32563,N_32912);
or U33192 (N_33192,N_32245,N_32360);
nand U33193 (N_33193,N_32882,N_32479);
nand U33194 (N_33194,N_32136,N_32248);
nand U33195 (N_33195,N_32403,N_32653);
nor U33196 (N_33196,N_32101,N_32525);
nor U33197 (N_33197,N_32745,N_32263);
and U33198 (N_33198,N_32420,N_32597);
nand U33199 (N_33199,N_32602,N_32909);
xor U33200 (N_33200,N_32769,N_32807);
and U33201 (N_33201,N_32395,N_32612);
and U33202 (N_33202,N_32065,N_32804);
nor U33203 (N_33203,N_32993,N_32741);
nor U33204 (N_33204,N_32614,N_32277);
xor U33205 (N_33205,N_32405,N_32791);
nor U33206 (N_33206,N_32710,N_32604);
xnor U33207 (N_33207,N_32444,N_32723);
nand U33208 (N_33208,N_32676,N_32354);
and U33209 (N_33209,N_32784,N_32187);
or U33210 (N_33210,N_32061,N_32705);
and U33211 (N_33211,N_32182,N_32829);
nand U33212 (N_33212,N_32049,N_32055);
and U33213 (N_33213,N_32487,N_32700);
nand U33214 (N_33214,N_32766,N_32861);
nor U33215 (N_33215,N_32941,N_32258);
and U33216 (N_33216,N_32211,N_32418);
and U33217 (N_33217,N_32387,N_32736);
and U33218 (N_33218,N_32887,N_32561);
xor U33219 (N_33219,N_32917,N_32494);
and U33220 (N_33220,N_32790,N_32347);
or U33221 (N_33221,N_32483,N_32063);
nand U33222 (N_33222,N_32380,N_32256);
nor U33223 (N_33223,N_32658,N_32082);
nor U33224 (N_33224,N_32367,N_32485);
and U33225 (N_33225,N_32787,N_32894);
xnor U33226 (N_33226,N_32566,N_32893);
xnor U33227 (N_33227,N_32402,N_32554);
nand U33228 (N_33228,N_32650,N_32595);
or U33229 (N_33229,N_32515,N_32001);
xor U33230 (N_33230,N_32973,N_32827);
nor U33231 (N_33231,N_32788,N_32711);
nand U33232 (N_33232,N_32166,N_32017);
and U33233 (N_33233,N_32611,N_32066);
xor U33234 (N_33234,N_32715,N_32783);
or U33235 (N_33235,N_32437,N_32657);
nand U33236 (N_33236,N_32204,N_32776);
and U33237 (N_33237,N_32366,N_32750);
xnor U33238 (N_33238,N_32180,N_32878);
or U33239 (N_33239,N_32134,N_32397);
and U33240 (N_33240,N_32013,N_32552);
and U33241 (N_33241,N_32352,N_32593);
and U33242 (N_33242,N_32164,N_32210);
and U33243 (N_33243,N_32522,N_32111);
or U33244 (N_33244,N_32129,N_32505);
xnor U33245 (N_33245,N_32994,N_32966);
and U33246 (N_33246,N_32249,N_32519);
nand U33247 (N_33247,N_32934,N_32517);
and U33248 (N_33248,N_32945,N_32895);
or U33249 (N_33249,N_32625,N_32537);
or U33250 (N_33250,N_32763,N_32530);
xnor U33251 (N_33251,N_32107,N_32478);
or U33252 (N_33252,N_32632,N_32120);
and U33253 (N_33253,N_32863,N_32417);
or U33254 (N_33254,N_32145,N_32949);
and U33255 (N_33255,N_32458,N_32472);
or U33256 (N_33256,N_32410,N_32152);
nand U33257 (N_33257,N_32908,N_32227);
nand U33258 (N_33258,N_32471,N_32447);
nand U33259 (N_33259,N_32044,N_32985);
and U33260 (N_33260,N_32035,N_32692);
or U33261 (N_33261,N_32755,N_32828);
or U33262 (N_33262,N_32675,N_32197);
xor U33263 (N_33263,N_32179,N_32311);
nor U33264 (N_33264,N_32693,N_32488);
or U33265 (N_33265,N_32474,N_32265);
or U33266 (N_33266,N_32098,N_32330);
nor U33267 (N_33267,N_32038,N_32160);
or U33268 (N_33268,N_32510,N_32454);
nor U33269 (N_33269,N_32284,N_32241);
and U33270 (N_33270,N_32450,N_32349);
or U33271 (N_33271,N_32833,N_32585);
and U33272 (N_33272,N_32826,N_32965);
or U33273 (N_33273,N_32928,N_32514);
nand U33274 (N_33274,N_32564,N_32911);
xor U33275 (N_33275,N_32794,N_32500);
and U33276 (N_33276,N_32824,N_32883);
xor U33277 (N_33277,N_32524,N_32857);
nor U33278 (N_33278,N_32747,N_32816);
nor U33279 (N_33279,N_32645,N_32639);
or U33280 (N_33280,N_32332,N_32702);
xor U33281 (N_33281,N_32637,N_32123);
and U33282 (N_33282,N_32324,N_32105);
or U33283 (N_33283,N_32400,N_32135);
xnor U33284 (N_33284,N_32546,N_32983);
or U33285 (N_33285,N_32767,N_32527);
nand U33286 (N_33286,N_32730,N_32296);
nand U33287 (N_33287,N_32963,N_32237);
or U33288 (N_33288,N_32900,N_32681);
nor U33289 (N_33289,N_32480,N_32226);
or U33290 (N_33290,N_32305,N_32881);
or U33291 (N_33291,N_32558,N_32078);
or U33292 (N_33292,N_32484,N_32531);
nor U33293 (N_33293,N_32529,N_32436);
xnor U33294 (N_33294,N_32355,N_32382);
or U33295 (N_33295,N_32714,N_32319);
or U33296 (N_33296,N_32666,N_32242);
nor U33297 (N_33297,N_32551,N_32261);
or U33298 (N_33298,N_32486,N_32663);
nand U33299 (N_33299,N_32214,N_32502);
and U33300 (N_33300,N_32737,N_32523);
xor U33301 (N_33301,N_32756,N_32503);
nor U33302 (N_33302,N_32888,N_32698);
nand U33303 (N_33303,N_32694,N_32590);
and U33304 (N_33304,N_32058,N_32339);
and U33305 (N_33305,N_32640,N_32961);
or U33306 (N_33306,N_32781,N_32429);
nand U33307 (N_33307,N_32024,N_32799);
or U33308 (N_33308,N_32677,N_32383);
nor U33309 (N_33309,N_32338,N_32353);
nand U33310 (N_33310,N_32699,N_32865);
nor U33311 (N_33311,N_32188,N_32997);
nor U33312 (N_33312,N_32445,N_32682);
and U33313 (N_33313,N_32691,N_32408);
xnor U33314 (N_33314,N_32610,N_32015);
xor U33315 (N_33315,N_32836,N_32688);
xor U33316 (N_33316,N_32097,N_32651);
or U33317 (N_33317,N_32616,N_32028);
nor U33318 (N_33318,N_32577,N_32940);
and U33319 (N_33319,N_32173,N_32642);
xnor U33320 (N_33320,N_32153,N_32206);
nand U33321 (N_33321,N_32452,N_32617);
nand U33322 (N_33322,N_32062,N_32516);
nand U33323 (N_33323,N_32685,N_32744);
nor U33324 (N_33324,N_32233,N_32376);
or U33325 (N_33325,N_32218,N_32114);
and U33326 (N_33326,N_32932,N_32507);
nand U33327 (N_33327,N_32222,N_32680);
and U33328 (N_33328,N_32369,N_32195);
and U33329 (N_33329,N_32202,N_32923);
or U33330 (N_33330,N_32673,N_32721);
xor U33331 (N_33331,N_32068,N_32465);
nor U33332 (N_33332,N_32972,N_32080);
xnor U33333 (N_33333,N_32907,N_32364);
or U33334 (N_33334,N_32085,N_32656);
or U33335 (N_33335,N_32926,N_32922);
nor U33336 (N_33336,N_32081,N_32426);
nand U33337 (N_33337,N_32154,N_32023);
and U33338 (N_33338,N_32176,N_32021);
nand U33339 (N_33339,N_32920,N_32124);
or U33340 (N_33340,N_32217,N_32325);
nand U33341 (N_33341,N_32161,N_32792);
nand U33342 (N_33342,N_32751,N_32368);
and U33343 (N_33343,N_32430,N_32406);
and U33344 (N_33344,N_32847,N_32424);
or U33345 (N_33345,N_32183,N_32722);
or U33346 (N_33346,N_32283,N_32142);
or U33347 (N_33347,N_32764,N_32990);
nor U33348 (N_33348,N_32493,N_32734);
or U33349 (N_33349,N_32868,N_32844);
or U33350 (N_33350,N_32396,N_32556);
nor U33351 (N_33351,N_32033,N_32328);
and U33352 (N_33352,N_32704,N_32906);
xor U33353 (N_33353,N_32253,N_32030);
nor U33354 (N_33354,N_32144,N_32520);
xor U33355 (N_33355,N_32877,N_32995);
or U33356 (N_33356,N_32411,N_32557);
or U33357 (N_33357,N_32022,N_32795);
xnor U33358 (N_33358,N_32508,N_32067);
nor U33359 (N_33359,N_32025,N_32378);
xor U33360 (N_33360,N_32575,N_32660);
or U33361 (N_33361,N_32267,N_32317);
xor U33362 (N_33362,N_32019,N_32316);
and U33363 (N_33363,N_32234,N_32125);
and U33364 (N_33364,N_32175,N_32652);
and U33365 (N_33365,N_32954,N_32800);
nor U33366 (N_33366,N_32304,N_32008);
nor U33367 (N_33367,N_32121,N_32607);
or U33368 (N_33368,N_32823,N_32313);
nand U33369 (N_33369,N_32026,N_32294);
nor U33370 (N_33370,N_32449,N_32252);
xor U33371 (N_33371,N_32362,N_32009);
or U33372 (N_33372,N_32560,N_32930);
nand U33373 (N_33373,N_32501,N_32384);
and U33374 (N_33374,N_32849,N_32209);
or U33375 (N_33375,N_32838,N_32988);
nand U33376 (N_33376,N_32431,N_32295);
nand U33377 (N_33377,N_32076,N_32905);
xor U33378 (N_33378,N_32373,N_32806);
nand U33379 (N_33379,N_32891,N_32538);
xor U33380 (N_33380,N_32944,N_32902);
nor U33381 (N_33381,N_32627,N_32785);
nor U33382 (N_33382,N_32583,N_32854);
and U33383 (N_33383,N_32761,N_32475);
xor U33384 (N_33384,N_32116,N_32186);
xor U33385 (N_33385,N_32259,N_32244);
xor U33386 (N_33386,N_32451,N_32077);
xor U33387 (N_33387,N_32053,N_32255);
nand U33388 (N_33388,N_32413,N_32236);
or U33389 (N_33389,N_32262,N_32535);
nor U33390 (N_33390,N_32171,N_32318);
and U33391 (N_33391,N_32143,N_32506);
nor U33392 (N_33392,N_32051,N_32036);
nor U33393 (N_33393,N_32407,N_32264);
and U33394 (N_33394,N_32643,N_32623);
and U33395 (N_33395,N_32155,N_32633);
xnor U33396 (N_33396,N_32323,N_32331);
nand U33397 (N_33397,N_32298,N_32442);
nand U33398 (N_33398,N_32626,N_32916);
xor U33399 (N_33399,N_32758,N_32588);
or U33400 (N_33400,N_32578,N_32286);
or U33401 (N_33401,N_32969,N_32148);
xnor U33402 (N_33402,N_32981,N_32113);
and U33403 (N_33403,N_32163,N_32439);
nand U33404 (N_33404,N_32919,N_32842);
nand U33405 (N_33405,N_32003,N_32073);
nand U33406 (N_33406,N_32768,N_32726);
xnor U33407 (N_33407,N_32314,N_32320);
xnor U33408 (N_33408,N_32345,N_32635);
nor U33409 (N_33409,N_32953,N_32309);
nor U33410 (N_33410,N_32670,N_32099);
xor U33411 (N_33411,N_32307,N_32959);
nor U33412 (N_33412,N_32775,N_32045);
and U33413 (N_33413,N_32232,N_32982);
nand U33414 (N_33414,N_32094,N_32567);
xnor U33415 (N_33415,N_32438,N_32899);
nor U33416 (N_33416,N_32706,N_32238);
nand U33417 (N_33417,N_32115,N_32002);
nand U33418 (N_33418,N_32201,N_32939);
or U33419 (N_33419,N_32540,N_32624);
and U33420 (N_33420,N_32831,N_32918);
xnor U33421 (N_33421,N_32459,N_32346);
xnor U33422 (N_33422,N_32606,N_32634);
or U33423 (N_33423,N_32856,N_32984);
xnor U33424 (N_33424,N_32873,N_32600);
or U33425 (N_33425,N_32089,N_32778);
nor U33426 (N_33426,N_32027,N_32117);
and U33427 (N_33427,N_32814,N_32351);
and U33428 (N_33428,N_32913,N_32780);
xnor U33429 (N_33429,N_32386,N_32638);
and U33430 (N_33430,N_32498,N_32762);
nor U33431 (N_33431,N_32528,N_32103);
or U33432 (N_33432,N_32468,N_32070);
xor U33433 (N_33433,N_32840,N_32671);
or U33434 (N_33434,N_32336,N_32832);
xor U33435 (N_33435,N_32727,N_32811);
nor U33436 (N_33436,N_32463,N_32270);
and U33437 (N_33437,N_32689,N_32880);
or U33438 (N_33438,N_32628,N_32235);
xor U33439 (N_33439,N_32010,N_32708);
and U33440 (N_33440,N_32509,N_32534);
and U33441 (N_33441,N_32246,N_32358);
and U33442 (N_33442,N_32543,N_32592);
or U33443 (N_33443,N_32835,N_32976);
nand U33444 (N_33444,N_32818,N_32457);
or U33445 (N_33445,N_32819,N_32955);
or U33446 (N_33446,N_32817,N_32477);
xor U33447 (N_33447,N_32719,N_32207);
nand U33448 (N_33448,N_32809,N_32371);
nand U33449 (N_33449,N_32925,N_32869);
nand U33450 (N_33450,N_32337,N_32490);
nor U33451 (N_33451,N_32434,N_32469);
xnor U33452 (N_33452,N_32914,N_32896);
nand U33453 (N_33453,N_32739,N_32724);
and U33454 (N_33454,N_32112,N_32759);
nor U33455 (N_33455,N_32219,N_32312);
nand U33456 (N_33456,N_32753,N_32977);
xnor U33457 (N_33457,N_32946,N_32952);
xnor U33458 (N_33458,N_32927,N_32453);
and U33459 (N_33459,N_32718,N_32326);
and U33460 (N_33460,N_32574,N_32697);
and U33461 (N_33461,N_32190,N_32394);
xor U33462 (N_33462,N_32467,N_32728);
or U33463 (N_33463,N_32110,N_32302);
or U33464 (N_33464,N_32970,N_32422);
nor U33465 (N_33465,N_32020,N_32591);
nor U33466 (N_33466,N_32212,N_32419);
nand U33467 (N_33467,N_32740,N_32250);
xnor U33468 (N_33468,N_32686,N_32571);
nand U33469 (N_33469,N_32938,N_32615);
and U33470 (N_33470,N_32732,N_32862);
nand U33471 (N_33471,N_32060,N_32220);
nand U33472 (N_33472,N_32964,N_32464);
and U33473 (N_33473,N_32243,N_32268);
nand U33474 (N_33474,N_32446,N_32388);
and U33475 (N_33475,N_32555,N_32473);
xor U33476 (N_33476,N_32772,N_32674);
xor U33477 (N_33477,N_32687,N_32958);
xor U33478 (N_33478,N_32139,N_32435);
or U33479 (N_33479,N_32377,N_32620);
or U33480 (N_33480,N_32254,N_32031);
or U33481 (N_33481,N_32462,N_32644);
nand U33482 (N_33482,N_32871,N_32879);
or U33483 (N_33483,N_32622,N_32149);
nand U33484 (N_33484,N_32960,N_32569);
nand U33485 (N_33485,N_32300,N_32864);
xor U33486 (N_33486,N_32203,N_32297);
xor U33487 (N_33487,N_32029,N_32513);
xor U33488 (N_33488,N_32415,N_32770);
or U33489 (N_33489,N_32504,N_32720);
and U33490 (N_33490,N_32696,N_32942);
xor U33491 (N_33491,N_32603,N_32884);
and U33492 (N_33492,N_32822,N_32851);
or U33493 (N_33493,N_32532,N_32157);
or U33494 (N_33494,N_32079,N_32897);
xnor U33495 (N_33495,N_32301,N_32618);
or U33496 (N_33496,N_32046,N_32813);
or U33497 (N_33497,N_32223,N_32497);
nor U33498 (N_33498,N_32285,N_32971);
or U33499 (N_33499,N_32329,N_32041);
nor U33500 (N_33500,N_32607,N_32340);
xnor U33501 (N_33501,N_32845,N_32521);
nand U33502 (N_33502,N_32144,N_32838);
and U33503 (N_33503,N_32235,N_32878);
xor U33504 (N_33504,N_32849,N_32419);
or U33505 (N_33505,N_32261,N_32705);
and U33506 (N_33506,N_32466,N_32536);
nor U33507 (N_33507,N_32959,N_32522);
xnor U33508 (N_33508,N_32133,N_32276);
nand U33509 (N_33509,N_32822,N_32279);
and U33510 (N_33510,N_32507,N_32824);
nor U33511 (N_33511,N_32916,N_32533);
nor U33512 (N_33512,N_32372,N_32735);
and U33513 (N_33513,N_32708,N_32322);
xor U33514 (N_33514,N_32345,N_32775);
or U33515 (N_33515,N_32514,N_32891);
or U33516 (N_33516,N_32076,N_32069);
or U33517 (N_33517,N_32009,N_32426);
and U33518 (N_33518,N_32449,N_32042);
nand U33519 (N_33519,N_32282,N_32305);
or U33520 (N_33520,N_32506,N_32946);
nor U33521 (N_33521,N_32870,N_32209);
and U33522 (N_33522,N_32703,N_32061);
or U33523 (N_33523,N_32162,N_32661);
nor U33524 (N_33524,N_32774,N_32528);
or U33525 (N_33525,N_32580,N_32983);
and U33526 (N_33526,N_32077,N_32445);
and U33527 (N_33527,N_32838,N_32458);
nand U33528 (N_33528,N_32161,N_32976);
and U33529 (N_33529,N_32223,N_32999);
nor U33530 (N_33530,N_32164,N_32872);
nand U33531 (N_33531,N_32538,N_32093);
and U33532 (N_33532,N_32820,N_32679);
and U33533 (N_33533,N_32243,N_32361);
nand U33534 (N_33534,N_32362,N_32022);
xnor U33535 (N_33535,N_32159,N_32117);
nor U33536 (N_33536,N_32771,N_32119);
or U33537 (N_33537,N_32991,N_32706);
nor U33538 (N_33538,N_32586,N_32556);
nor U33539 (N_33539,N_32491,N_32474);
nor U33540 (N_33540,N_32086,N_32974);
and U33541 (N_33541,N_32534,N_32797);
nand U33542 (N_33542,N_32058,N_32884);
and U33543 (N_33543,N_32514,N_32475);
and U33544 (N_33544,N_32078,N_32995);
and U33545 (N_33545,N_32635,N_32629);
nor U33546 (N_33546,N_32701,N_32062);
nor U33547 (N_33547,N_32340,N_32422);
nor U33548 (N_33548,N_32540,N_32461);
or U33549 (N_33549,N_32948,N_32436);
and U33550 (N_33550,N_32343,N_32173);
xnor U33551 (N_33551,N_32981,N_32183);
nand U33552 (N_33552,N_32830,N_32182);
or U33553 (N_33553,N_32623,N_32654);
nand U33554 (N_33554,N_32649,N_32619);
or U33555 (N_33555,N_32035,N_32647);
or U33556 (N_33556,N_32288,N_32727);
nand U33557 (N_33557,N_32989,N_32475);
nor U33558 (N_33558,N_32448,N_32334);
nor U33559 (N_33559,N_32042,N_32873);
nor U33560 (N_33560,N_32699,N_32020);
and U33561 (N_33561,N_32987,N_32749);
or U33562 (N_33562,N_32283,N_32485);
and U33563 (N_33563,N_32611,N_32162);
nand U33564 (N_33564,N_32669,N_32416);
nor U33565 (N_33565,N_32993,N_32472);
nand U33566 (N_33566,N_32776,N_32299);
nor U33567 (N_33567,N_32648,N_32768);
nor U33568 (N_33568,N_32727,N_32621);
or U33569 (N_33569,N_32608,N_32871);
nor U33570 (N_33570,N_32492,N_32613);
nand U33571 (N_33571,N_32649,N_32477);
xor U33572 (N_33572,N_32130,N_32147);
or U33573 (N_33573,N_32161,N_32002);
or U33574 (N_33574,N_32438,N_32686);
nand U33575 (N_33575,N_32744,N_32085);
nor U33576 (N_33576,N_32880,N_32497);
and U33577 (N_33577,N_32277,N_32509);
nor U33578 (N_33578,N_32230,N_32333);
and U33579 (N_33579,N_32530,N_32205);
xor U33580 (N_33580,N_32377,N_32118);
nor U33581 (N_33581,N_32126,N_32477);
and U33582 (N_33582,N_32330,N_32915);
nor U33583 (N_33583,N_32292,N_32867);
and U33584 (N_33584,N_32225,N_32289);
and U33585 (N_33585,N_32086,N_32970);
nand U33586 (N_33586,N_32080,N_32575);
nor U33587 (N_33587,N_32037,N_32889);
or U33588 (N_33588,N_32880,N_32151);
and U33589 (N_33589,N_32082,N_32524);
or U33590 (N_33590,N_32226,N_32458);
and U33591 (N_33591,N_32777,N_32902);
and U33592 (N_33592,N_32793,N_32753);
or U33593 (N_33593,N_32025,N_32070);
nand U33594 (N_33594,N_32413,N_32642);
nand U33595 (N_33595,N_32168,N_32506);
nand U33596 (N_33596,N_32424,N_32846);
nand U33597 (N_33597,N_32697,N_32817);
and U33598 (N_33598,N_32999,N_32595);
and U33599 (N_33599,N_32372,N_32421);
and U33600 (N_33600,N_32619,N_32199);
xor U33601 (N_33601,N_32571,N_32440);
xor U33602 (N_33602,N_32541,N_32745);
nor U33603 (N_33603,N_32690,N_32116);
nor U33604 (N_33604,N_32366,N_32393);
or U33605 (N_33605,N_32773,N_32958);
xnor U33606 (N_33606,N_32778,N_32158);
nand U33607 (N_33607,N_32917,N_32837);
and U33608 (N_33608,N_32719,N_32807);
nor U33609 (N_33609,N_32219,N_32429);
xor U33610 (N_33610,N_32681,N_32534);
nor U33611 (N_33611,N_32493,N_32158);
nand U33612 (N_33612,N_32013,N_32695);
or U33613 (N_33613,N_32476,N_32978);
or U33614 (N_33614,N_32456,N_32604);
and U33615 (N_33615,N_32450,N_32688);
nand U33616 (N_33616,N_32971,N_32458);
and U33617 (N_33617,N_32437,N_32129);
xnor U33618 (N_33618,N_32002,N_32227);
nor U33619 (N_33619,N_32279,N_32936);
nor U33620 (N_33620,N_32986,N_32824);
nand U33621 (N_33621,N_32378,N_32885);
nand U33622 (N_33622,N_32049,N_32300);
and U33623 (N_33623,N_32922,N_32910);
nor U33624 (N_33624,N_32157,N_32387);
nand U33625 (N_33625,N_32401,N_32866);
or U33626 (N_33626,N_32817,N_32776);
and U33627 (N_33627,N_32468,N_32238);
and U33628 (N_33628,N_32132,N_32928);
and U33629 (N_33629,N_32381,N_32008);
nand U33630 (N_33630,N_32821,N_32474);
nand U33631 (N_33631,N_32191,N_32248);
nor U33632 (N_33632,N_32008,N_32553);
nand U33633 (N_33633,N_32437,N_32276);
or U33634 (N_33634,N_32886,N_32851);
nor U33635 (N_33635,N_32632,N_32210);
or U33636 (N_33636,N_32162,N_32372);
nor U33637 (N_33637,N_32894,N_32828);
nor U33638 (N_33638,N_32281,N_32836);
xor U33639 (N_33639,N_32369,N_32999);
nand U33640 (N_33640,N_32523,N_32853);
xnor U33641 (N_33641,N_32436,N_32070);
and U33642 (N_33642,N_32883,N_32960);
or U33643 (N_33643,N_32028,N_32768);
and U33644 (N_33644,N_32107,N_32163);
nor U33645 (N_33645,N_32597,N_32559);
nand U33646 (N_33646,N_32610,N_32214);
nand U33647 (N_33647,N_32244,N_32300);
nor U33648 (N_33648,N_32706,N_32584);
nor U33649 (N_33649,N_32327,N_32542);
and U33650 (N_33650,N_32266,N_32828);
xor U33651 (N_33651,N_32829,N_32208);
nand U33652 (N_33652,N_32495,N_32537);
nor U33653 (N_33653,N_32493,N_32690);
xnor U33654 (N_33654,N_32216,N_32460);
and U33655 (N_33655,N_32087,N_32394);
and U33656 (N_33656,N_32449,N_32578);
xor U33657 (N_33657,N_32318,N_32890);
or U33658 (N_33658,N_32281,N_32405);
xnor U33659 (N_33659,N_32122,N_32095);
nand U33660 (N_33660,N_32268,N_32991);
xor U33661 (N_33661,N_32117,N_32195);
and U33662 (N_33662,N_32174,N_32085);
or U33663 (N_33663,N_32877,N_32937);
or U33664 (N_33664,N_32188,N_32688);
nor U33665 (N_33665,N_32681,N_32549);
xnor U33666 (N_33666,N_32461,N_32071);
or U33667 (N_33667,N_32761,N_32605);
nand U33668 (N_33668,N_32380,N_32884);
xor U33669 (N_33669,N_32498,N_32377);
and U33670 (N_33670,N_32671,N_32360);
nand U33671 (N_33671,N_32834,N_32045);
xor U33672 (N_33672,N_32299,N_32723);
nand U33673 (N_33673,N_32538,N_32002);
or U33674 (N_33674,N_32169,N_32773);
nor U33675 (N_33675,N_32886,N_32029);
xor U33676 (N_33676,N_32473,N_32718);
nor U33677 (N_33677,N_32002,N_32399);
or U33678 (N_33678,N_32363,N_32422);
or U33679 (N_33679,N_32482,N_32226);
and U33680 (N_33680,N_32910,N_32509);
xnor U33681 (N_33681,N_32270,N_32613);
and U33682 (N_33682,N_32296,N_32044);
nand U33683 (N_33683,N_32184,N_32382);
nor U33684 (N_33684,N_32042,N_32040);
nand U33685 (N_33685,N_32689,N_32123);
nor U33686 (N_33686,N_32377,N_32300);
or U33687 (N_33687,N_32790,N_32108);
xor U33688 (N_33688,N_32138,N_32868);
or U33689 (N_33689,N_32189,N_32420);
xnor U33690 (N_33690,N_32518,N_32194);
xnor U33691 (N_33691,N_32320,N_32123);
and U33692 (N_33692,N_32218,N_32502);
nand U33693 (N_33693,N_32349,N_32818);
xnor U33694 (N_33694,N_32499,N_32333);
or U33695 (N_33695,N_32407,N_32244);
xor U33696 (N_33696,N_32585,N_32834);
xor U33697 (N_33697,N_32160,N_32753);
nor U33698 (N_33698,N_32366,N_32638);
or U33699 (N_33699,N_32516,N_32544);
nand U33700 (N_33700,N_32819,N_32202);
and U33701 (N_33701,N_32185,N_32385);
xor U33702 (N_33702,N_32215,N_32243);
and U33703 (N_33703,N_32635,N_32529);
nor U33704 (N_33704,N_32044,N_32851);
and U33705 (N_33705,N_32668,N_32598);
xor U33706 (N_33706,N_32416,N_32853);
nand U33707 (N_33707,N_32500,N_32467);
xor U33708 (N_33708,N_32193,N_32485);
and U33709 (N_33709,N_32452,N_32875);
nand U33710 (N_33710,N_32356,N_32670);
nor U33711 (N_33711,N_32081,N_32921);
or U33712 (N_33712,N_32397,N_32352);
and U33713 (N_33713,N_32114,N_32539);
and U33714 (N_33714,N_32799,N_32852);
nor U33715 (N_33715,N_32358,N_32146);
and U33716 (N_33716,N_32454,N_32701);
and U33717 (N_33717,N_32746,N_32017);
xor U33718 (N_33718,N_32045,N_32255);
or U33719 (N_33719,N_32625,N_32304);
xor U33720 (N_33720,N_32848,N_32990);
or U33721 (N_33721,N_32699,N_32134);
nand U33722 (N_33722,N_32175,N_32830);
nor U33723 (N_33723,N_32367,N_32351);
xor U33724 (N_33724,N_32271,N_32164);
nand U33725 (N_33725,N_32143,N_32773);
or U33726 (N_33726,N_32110,N_32486);
xor U33727 (N_33727,N_32787,N_32182);
nand U33728 (N_33728,N_32460,N_32888);
or U33729 (N_33729,N_32166,N_32467);
xor U33730 (N_33730,N_32304,N_32083);
and U33731 (N_33731,N_32605,N_32942);
nor U33732 (N_33732,N_32796,N_32117);
and U33733 (N_33733,N_32003,N_32789);
nand U33734 (N_33734,N_32558,N_32307);
xnor U33735 (N_33735,N_32877,N_32228);
nand U33736 (N_33736,N_32247,N_32412);
nor U33737 (N_33737,N_32860,N_32372);
nand U33738 (N_33738,N_32565,N_32260);
nand U33739 (N_33739,N_32505,N_32650);
xor U33740 (N_33740,N_32246,N_32457);
xor U33741 (N_33741,N_32019,N_32038);
nor U33742 (N_33742,N_32081,N_32861);
nor U33743 (N_33743,N_32926,N_32095);
xnor U33744 (N_33744,N_32844,N_32446);
xor U33745 (N_33745,N_32727,N_32992);
and U33746 (N_33746,N_32314,N_32860);
or U33747 (N_33747,N_32188,N_32176);
and U33748 (N_33748,N_32014,N_32651);
nor U33749 (N_33749,N_32688,N_32509);
nor U33750 (N_33750,N_32562,N_32274);
nand U33751 (N_33751,N_32004,N_32012);
xor U33752 (N_33752,N_32685,N_32112);
nor U33753 (N_33753,N_32131,N_32209);
xnor U33754 (N_33754,N_32658,N_32706);
or U33755 (N_33755,N_32561,N_32261);
or U33756 (N_33756,N_32010,N_32993);
or U33757 (N_33757,N_32202,N_32891);
xor U33758 (N_33758,N_32946,N_32273);
nand U33759 (N_33759,N_32270,N_32049);
and U33760 (N_33760,N_32521,N_32170);
or U33761 (N_33761,N_32911,N_32816);
xor U33762 (N_33762,N_32406,N_32312);
and U33763 (N_33763,N_32442,N_32384);
and U33764 (N_33764,N_32114,N_32670);
xor U33765 (N_33765,N_32062,N_32850);
xnor U33766 (N_33766,N_32897,N_32557);
and U33767 (N_33767,N_32531,N_32631);
xnor U33768 (N_33768,N_32264,N_32126);
nand U33769 (N_33769,N_32504,N_32703);
or U33770 (N_33770,N_32037,N_32132);
or U33771 (N_33771,N_32062,N_32694);
nor U33772 (N_33772,N_32991,N_32774);
nand U33773 (N_33773,N_32370,N_32938);
nor U33774 (N_33774,N_32548,N_32785);
nor U33775 (N_33775,N_32826,N_32933);
nor U33776 (N_33776,N_32105,N_32834);
nor U33777 (N_33777,N_32506,N_32136);
and U33778 (N_33778,N_32085,N_32925);
and U33779 (N_33779,N_32658,N_32093);
nor U33780 (N_33780,N_32315,N_32906);
and U33781 (N_33781,N_32925,N_32199);
xor U33782 (N_33782,N_32487,N_32959);
and U33783 (N_33783,N_32478,N_32233);
xnor U33784 (N_33784,N_32970,N_32446);
or U33785 (N_33785,N_32108,N_32581);
xnor U33786 (N_33786,N_32092,N_32963);
and U33787 (N_33787,N_32867,N_32938);
nand U33788 (N_33788,N_32871,N_32373);
or U33789 (N_33789,N_32943,N_32767);
nand U33790 (N_33790,N_32125,N_32381);
xnor U33791 (N_33791,N_32311,N_32713);
nand U33792 (N_33792,N_32052,N_32692);
nor U33793 (N_33793,N_32933,N_32010);
or U33794 (N_33794,N_32566,N_32005);
or U33795 (N_33795,N_32779,N_32237);
or U33796 (N_33796,N_32335,N_32170);
or U33797 (N_33797,N_32916,N_32364);
nand U33798 (N_33798,N_32543,N_32453);
nand U33799 (N_33799,N_32342,N_32830);
nand U33800 (N_33800,N_32721,N_32277);
or U33801 (N_33801,N_32678,N_32861);
or U33802 (N_33802,N_32371,N_32353);
nand U33803 (N_33803,N_32059,N_32187);
nand U33804 (N_33804,N_32872,N_32925);
xor U33805 (N_33805,N_32155,N_32172);
nor U33806 (N_33806,N_32287,N_32017);
nor U33807 (N_33807,N_32178,N_32919);
and U33808 (N_33808,N_32088,N_32125);
and U33809 (N_33809,N_32792,N_32965);
and U33810 (N_33810,N_32179,N_32301);
or U33811 (N_33811,N_32809,N_32793);
or U33812 (N_33812,N_32555,N_32934);
xnor U33813 (N_33813,N_32990,N_32708);
xnor U33814 (N_33814,N_32307,N_32062);
and U33815 (N_33815,N_32769,N_32185);
nand U33816 (N_33816,N_32684,N_32112);
xnor U33817 (N_33817,N_32081,N_32159);
xor U33818 (N_33818,N_32831,N_32378);
or U33819 (N_33819,N_32805,N_32243);
nor U33820 (N_33820,N_32715,N_32296);
nand U33821 (N_33821,N_32569,N_32140);
nand U33822 (N_33822,N_32474,N_32355);
or U33823 (N_33823,N_32444,N_32819);
nor U33824 (N_33824,N_32026,N_32273);
nor U33825 (N_33825,N_32991,N_32462);
xnor U33826 (N_33826,N_32162,N_32628);
and U33827 (N_33827,N_32345,N_32268);
nand U33828 (N_33828,N_32315,N_32207);
nor U33829 (N_33829,N_32368,N_32048);
nor U33830 (N_33830,N_32656,N_32740);
xnor U33831 (N_33831,N_32320,N_32436);
or U33832 (N_33832,N_32535,N_32849);
or U33833 (N_33833,N_32748,N_32535);
xor U33834 (N_33834,N_32880,N_32412);
nand U33835 (N_33835,N_32378,N_32211);
xnor U33836 (N_33836,N_32451,N_32402);
nand U33837 (N_33837,N_32347,N_32806);
nor U33838 (N_33838,N_32766,N_32688);
xnor U33839 (N_33839,N_32608,N_32522);
or U33840 (N_33840,N_32170,N_32300);
nor U33841 (N_33841,N_32215,N_32492);
nand U33842 (N_33842,N_32847,N_32205);
xnor U33843 (N_33843,N_32186,N_32223);
nand U33844 (N_33844,N_32273,N_32049);
nor U33845 (N_33845,N_32300,N_32390);
or U33846 (N_33846,N_32453,N_32547);
and U33847 (N_33847,N_32499,N_32411);
xnor U33848 (N_33848,N_32974,N_32319);
and U33849 (N_33849,N_32036,N_32366);
or U33850 (N_33850,N_32254,N_32927);
and U33851 (N_33851,N_32977,N_32166);
nor U33852 (N_33852,N_32961,N_32656);
nand U33853 (N_33853,N_32728,N_32245);
nor U33854 (N_33854,N_32316,N_32775);
nand U33855 (N_33855,N_32294,N_32634);
xnor U33856 (N_33856,N_32988,N_32284);
nand U33857 (N_33857,N_32187,N_32818);
nand U33858 (N_33858,N_32206,N_32664);
or U33859 (N_33859,N_32684,N_32822);
nor U33860 (N_33860,N_32600,N_32571);
nor U33861 (N_33861,N_32891,N_32567);
or U33862 (N_33862,N_32631,N_32237);
xnor U33863 (N_33863,N_32852,N_32869);
or U33864 (N_33864,N_32991,N_32274);
and U33865 (N_33865,N_32559,N_32339);
or U33866 (N_33866,N_32733,N_32269);
and U33867 (N_33867,N_32851,N_32507);
and U33868 (N_33868,N_32911,N_32806);
nor U33869 (N_33869,N_32705,N_32519);
and U33870 (N_33870,N_32962,N_32357);
nor U33871 (N_33871,N_32352,N_32223);
nand U33872 (N_33872,N_32975,N_32384);
and U33873 (N_33873,N_32509,N_32118);
and U33874 (N_33874,N_32453,N_32714);
nor U33875 (N_33875,N_32318,N_32250);
nor U33876 (N_33876,N_32908,N_32350);
and U33877 (N_33877,N_32297,N_32199);
nor U33878 (N_33878,N_32581,N_32453);
and U33879 (N_33879,N_32722,N_32276);
nor U33880 (N_33880,N_32855,N_32742);
or U33881 (N_33881,N_32702,N_32414);
xor U33882 (N_33882,N_32985,N_32040);
or U33883 (N_33883,N_32032,N_32472);
or U33884 (N_33884,N_32494,N_32448);
nand U33885 (N_33885,N_32283,N_32640);
nor U33886 (N_33886,N_32436,N_32229);
and U33887 (N_33887,N_32551,N_32733);
nor U33888 (N_33888,N_32256,N_32257);
nand U33889 (N_33889,N_32835,N_32941);
nand U33890 (N_33890,N_32495,N_32572);
or U33891 (N_33891,N_32637,N_32313);
xor U33892 (N_33892,N_32594,N_32085);
and U33893 (N_33893,N_32101,N_32040);
xnor U33894 (N_33894,N_32039,N_32126);
or U33895 (N_33895,N_32375,N_32764);
xor U33896 (N_33896,N_32253,N_32770);
nand U33897 (N_33897,N_32944,N_32899);
xor U33898 (N_33898,N_32112,N_32870);
or U33899 (N_33899,N_32839,N_32081);
nand U33900 (N_33900,N_32766,N_32877);
or U33901 (N_33901,N_32197,N_32356);
nor U33902 (N_33902,N_32872,N_32712);
and U33903 (N_33903,N_32711,N_32659);
nor U33904 (N_33904,N_32899,N_32073);
nor U33905 (N_33905,N_32999,N_32334);
nor U33906 (N_33906,N_32199,N_32623);
and U33907 (N_33907,N_32294,N_32337);
or U33908 (N_33908,N_32529,N_32110);
xnor U33909 (N_33909,N_32238,N_32831);
nor U33910 (N_33910,N_32254,N_32387);
nor U33911 (N_33911,N_32782,N_32333);
and U33912 (N_33912,N_32399,N_32422);
nor U33913 (N_33913,N_32241,N_32649);
nor U33914 (N_33914,N_32798,N_32665);
or U33915 (N_33915,N_32286,N_32335);
or U33916 (N_33916,N_32371,N_32126);
xor U33917 (N_33917,N_32928,N_32632);
and U33918 (N_33918,N_32645,N_32765);
or U33919 (N_33919,N_32182,N_32177);
xnor U33920 (N_33920,N_32485,N_32476);
nand U33921 (N_33921,N_32415,N_32954);
or U33922 (N_33922,N_32840,N_32409);
xnor U33923 (N_33923,N_32641,N_32152);
nor U33924 (N_33924,N_32050,N_32948);
xor U33925 (N_33925,N_32232,N_32094);
nor U33926 (N_33926,N_32177,N_32233);
xor U33927 (N_33927,N_32003,N_32919);
and U33928 (N_33928,N_32366,N_32713);
and U33929 (N_33929,N_32746,N_32950);
and U33930 (N_33930,N_32940,N_32614);
or U33931 (N_33931,N_32527,N_32557);
nor U33932 (N_33932,N_32820,N_32516);
and U33933 (N_33933,N_32265,N_32691);
xnor U33934 (N_33934,N_32453,N_32708);
and U33935 (N_33935,N_32952,N_32686);
xnor U33936 (N_33936,N_32926,N_32302);
or U33937 (N_33937,N_32687,N_32834);
nor U33938 (N_33938,N_32837,N_32102);
and U33939 (N_33939,N_32173,N_32921);
nand U33940 (N_33940,N_32171,N_32748);
and U33941 (N_33941,N_32690,N_32193);
nor U33942 (N_33942,N_32680,N_32082);
nor U33943 (N_33943,N_32841,N_32201);
or U33944 (N_33944,N_32873,N_32753);
or U33945 (N_33945,N_32005,N_32801);
xnor U33946 (N_33946,N_32176,N_32401);
xor U33947 (N_33947,N_32782,N_32242);
nand U33948 (N_33948,N_32870,N_32219);
and U33949 (N_33949,N_32376,N_32312);
nand U33950 (N_33950,N_32056,N_32165);
nor U33951 (N_33951,N_32159,N_32398);
and U33952 (N_33952,N_32444,N_32607);
and U33953 (N_33953,N_32352,N_32418);
xor U33954 (N_33954,N_32212,N_32822);
nand U33955 (N_33955,N_32781,N_32316);
nor U33956 (N_33956,N_32308,N_32046);
or U33957 (N_33957,N_32041,N_32961);
xor U33958 (N_33958,N_32424,N_32861);
or U33959 (N_33959,N_32591,N_32723);
nand U33960 (N_33960,N_32037,N_32116);
xnor U33961 (N_33961,N_32534,N_32538);
and U33962 (N_33962,N_32274,N_32674);
and U33963 (N_33963,N_32134,N_32273);
nand U33964 (N_33964,N_32599,N_32847);
and U33965 (N_33965,N_32424,N_32552);
nor U33966 (N_33966,N_32426,N_32667);
and U33967 (N_33967,N_32802,N_32505);
xnor U33968 (N_33968,N_32111,N_32957);
or U33969 (N_33969,N_32037,N_32978);
nor U33970 (N_33970,N_32433,N_32248);
nor U33971 (N_33971,N_32222,N_32215);
xnor U33972 (N_33972,N_32546,N_32818);
or U33973 (N_33973,N_32651,N_32976);
xnor U33974 (N_33974,N_32029,N_32509);
nand U33975 (N_33975,N_32279,N_32803);
and U33976 (N_33976,N_32990,N_32340);
nor U33977 (N_33977,N_32103,N_32701);
nor U33978 (N_33978,N_32601,N_32752);
nand U33979 (N_33979,N_32196,N_32308);
nand U33980 (N_33980,N_32891,N_32157);
nor U33981 (N_33981,N_32827,N_32129);
or U33982 (N_33982,N_32665,N_32189);
nand U33983 (N_33983,N_32691,N_32925);
or U33984 (N_33984,N_32942,N_32882);
and U33985 (N_33985,N_32453,N_32622);
or U33986 (N_33986,N_32489,N_32573);
xor U33987 (N_33987,N_32177,N_32735);
and U33988 (N_33988,N_32467,N_32126);
nor U33989 (N_33989,N_32876,N_32810);
nand U33990 (N_33990,N_32330,N_32026);
nand U33991 (N_33991,N_32457,N_32108);
nand U33992 (N_33992,N_32472,N_32573);
and U33993 (N_33993,N_32864,N_32140);
xor U33994 (N_33994,N_32888,N_32174);
and U33995 (N_33995,N_32775,N_32485);
nand U33996 (N_33996,N_32652,N_32633);
nor U33997 (N_33997,N_32334,N_32525);
nor U33998 (N_33998,N_32716,N_32721);
or U33999 (N_33999,N_32957,N_32109);
and U34000 (N_34000,N_33458,N_33525);
or U34001 (N_34001,N_33705,N_33621);
nand U34002 (N_34002,N_33051,N_33637);
nand U34003 (N_34003,N_33822,N_33745);
or U34004 (N_34004,N_33395,N_33563);
nand U34005 (N_34005,N_33918,N_33583);
nor U34006 (N_34006,N_33842,N_33562);
nor U34007 (N_34007,N_33509,N_33193);
nand U34008 (N_34008,N_33283,N_33472);
and U34009 (N_34009,N_33712,N_33826);
nor U34010 (N_34010,N_33612,N_33076);
nand U34011 (N_34011,N_33270,N_33451);
or U34012 (N_34012,N_33470,N_33956);
or U34013 (N_34013,N_33486,N_33915);
xor U34014 (N_34014,N_33813,N_33540);
nand U34015 (N_34015,N_33875,N_33805);
and U34016 (N_34016,N_33972,N_33827);
xor U34017 (N_34017,N_33992,N_33169);
nand U34018 (N_34018,N_33232,N_33476);
xor U34019 (N_34019,N_33917,N_33181);
and U34020 (N_34020,N_33921,N_33494);
nor U34021 (N_34021,N_33715,N_33057);
or U34022 (N_34022,N_33359,N_33198);
nand U34023 (N_34023,N_33686,N_33244);
or U34024 (N_34024,N_33610,N_33774);
nand U34025 (N_34025,N_33250,N_33024);
or U34026 (N_34026,N_33424,N_33041);
nor U34027 (N_34027,N_33381,N_33350);
nor U34028 (N_34028,N_33134,N_33707);
nand U34029 (N_34029,N_33659,N_33197);
nand U34030 (N_34030,N_33256,N_33086);
nor U34031 (N_34031,N_33434,N_33599);
nand U34032 (N_34032,N_33518,N_33721);
and U34033 (N_34033,N_33653,N_33087);
or U34034 (N_34034,N_33243,N_33904);
xor U34035 (N_34035,N_33015,N_33454);
xor U34036 (N_34036,N_33406,N_33431);
nor U34037 (N_34037,N_33655,N_33186);
nand U34038 (N_34038,N_33772,N_33098);
nor U34039 (N_34039,N_33988,N_33668);
nor U34040 (N_34040,N_33611,N_33142);
or U34041 (N_34041,N_33515,N_33366);
or U34042 (N_34042,N_33965,N_33009);
xnor U34043 (N_34043,N_33025,N_33122);
and U34044 (N_34044,N_33558,N_33464);
xor U34045 (N_34045,N_33478,N_33561);
and U34046 (N_34046,N_33764,N_33274);
and U34047 (N_34047,N_33370,N_33364);
nor U34048 (N_34048,N_33940,N_33786);
xor U34049 (N_34049,N_33297,N_33045);
xor U34050 (N_34050,N_33631,N_33264);
nand U34051 (N_34051,N_33908,N_33436);
and U34052 (N_34052,N_33731,N_33097);
nor U34053 (N_34053,N_33639,N_33996);
or U34054 (N_34054,N_33156,N_33688);
xnor U34055 (N_34055,N_33132,N_33717);
and U34056 (N_34056,N_33167,N_33199);
nand U34057 (N_34057,N_33962,N_33835);
nor U34058 (N_34058,N_33204,N_33006);
nand U34059 (N_34059,N_33517,N_33588);
nand U34060 (N_34060,N_33897,N_33994);
xnor U34061 (N_34061,N_33691,N_33229);
xor U34062 (N_34062,N_33175,N_33855);
xor U34063 (N_34063,N_33834,N_33031);
and U34064 (N_34064,N_33234,N_33579);
nor U34065 (N_34065,N_33184,N_33516);
nor U34066 (N_34066,N_33023,N_33866);
xor U34067 (N_34067,N_33874,N_33766);
and U34068 (N_34068,N_33352,N_33439);
xor U34069 (N_34069,N_33849,N_33000);
nand U34070 (N_34070,N_33791,N_33168);
or U34071 (N_34071,N_33943,N_33238);
xor U34072 (N_34072,N_33730,N_33047);
nand U34073 (N_34073,N_33339,N_33795);
nor U34074 (N_34074,N_33262,N_33550);
or U34075 (N_34075,N_33582,N_33081);
xor U34076 (N_34076,N_33094,N_33755);
or U34077 (N_34077,N_33614,N_33480);
nand U34078 (N_34078,N_33475,N_33662);
xnor U34079 (N_34079,N_33393,N_33372);
nand U34080 (N_34080,N_33684,N_33012);
xnor U34081 (N_34081,N_33208,N_33895);
nand U34082 (N_34082,N_33548,N_33288);
and U34083 (N_34083,N_33195,N_33459);
and U34084 (N_34084,N_33894,N_33964);
nand U34085 (N_34085,N_33983,N_33280);
nand U34086 (N_34086,N_33898,N_33819);
xor U34087 (N_34087,N_33419,N_33117);
nand U34088 (N_34088,N_33798,N_33541);
and U34089 (N_34089,N_33481,N_33971);
or U34090 (N_34090,N_33001,N_33130);
nand U34091 (N_34091,N_33353,N_33360);
nand U34092 (N_34092,N_33846,N_33151);
nor U34093 (N_34093,N_33733,N_33106);
nand U34094 (N_34094,N_33467,N_33398);
and U34095 (N_34095,N_33066,N_33387);
xor U34096 (N_34096,N_33881,N_33260);
and U34097 (N_34097,N_33604,N_33585);
nand U34098 (N_34098,N_33811,N_33946);
or U34099 (N_34099,N_33149,N_33258);
xor U34100 (N_34100,N_33865,N_33375);
nand U34101 (N_34101,N_33211,N_33746);
or U34102 (N_34102,N_33643,N_33060);
and U34103 (N_34103,N_33871,N_33756);
nand U34104 (N_34104,N_33088,N_33416);
and U34105 (N_34105,N_33951,N_33650);
and U34106 (N_34106,N_33050,N_33037);
or U34107 (N_34107,N_33796,N_33008);
and U34108 (N_34108,N_33010,N_33404);
and U34109 (N_34109,N_33083,N_33433);
or U34110 (N_34110,N_33413,N_33137);
and U34111 (N_34111,N_33335,N_33602);
nor U34112 (N_34112,N_33292,N_33929);
nand U34113 (N_34113,N_33285,N_33299);
nand U34114 (N_34114,N_33327,N_33544);
or U34115 (N_34115,N_33128,N_33435);
or U34116 (N_34116,N_33392,N_33160);
nand U34117 (N_34117,N_33155,N_33036);
or U34118 (N_34118,N_33374,N_33950);
nor U34119 (N_34119,N_33944,N_33751);
nand U34120 (N_34120,N_33841,N_33832);
or U34121 (N_34121,N_33030,N_33565);
xnor U34122 (N_34122,N_33221,N_33447);
nand U34123 (N_34123,N_33963,N_33159);
or U34124 (N_34124,N_33456,N_33560);
or U34125 (N_34125,N_33601,N_33933);
nor U34126 (N_34126,N_33263,N_33147);
or U34127 (N_34127,N_33093,N_33089);
and U34128 (N_34128,N_33213,N_33308);
xor U34129 (N_34129,N_33889,N_33830);
and U34130 (N_34130,N_33616,N_33411);
nand U34131 (N_34131,N_33183,N_33491);
or U34132 (N_34132,N_33729,N_33354);
and U34133 (N_34133,N_33864,N_33109);
nor U34134 (N_34134,N_33329,N_33559);
or U34135 (N_34135,N_33649,N_33719);
nand U34136 (N_34136,N_33514,N_33222);
and U34137 (N_34137,N_33104,N_33629);
nor U34138 (N_34138,N_33551,N_33131);
nand U34139 (N_34139,N_33018,N_33936);
and U34140 (N_34140,N_33291,N_33461);
and U34141 (N_34141,N_33276,N_33091);
nor U34142 (N_34142,N_33824,N_33342);
and U34143 (N_34143,N_33882,N_33888);
xor U34144 (N_34144,N_33513,N_33337);
and U34145 (N_34145,N_33430,N_33926);
xor U34146 (N_34146,N_33646,N_33334);
nor U34147 (N_34147,N_33574,N_33293);
nor U34148 (N_34148,N_33836,N_33343);
xor U34149 (N_34149,N_33537,N_33654);
and U34150 (N_34150,N_33900,N_33325);
or U34151 (N_34151,N_33931,N_33444);
nand U34152 (N_34152,N_33749,N_33272);
xnor U34153 (N_34153,N_33483,N_33991);
nor U34154 (N_34154,N_33641,N_33538);
and U34155 (N_34155,N_33512,N_33355);
and U34156 (N_34156,N_33448,N_33273);
and U34157 (N_34157,N_33687,N_33150);
and U34158 (N_34158,N_33027,N_33403);
xor U34159 (N_34159,N_33368,N_33862);
or U34160 (N_34160,N_33787,N_33676);
xor U34161 (N_34161,N_33196,N_33125);
xnor U34162 (N_34162,N_33744,N_33205);
nand U34163 (N_34163,N_33529,N_33628);
xnor U34164 (N_34164,N_33870,N_33178);
and U34165 (N_34165,N_33911,N_33271);
xor U34166 (N_34166,N_33408,N_33941);
xnor U34167 (N_34167,N_33703,N_33177);
and U34168 (N_34168,N_33879,N_33054);
or U34169 (N_34169,N_33575,N_33215);
xnor U34170 (N_34170,N_33652,N_33477);
and U34171 (N_34171,N_33697,N_33982);
and U34172 (N_34172,N_33453,N_33939);
or U34173 (N_34173,N_33927,N_33121);
xor U34174 (N_34174,N_33407,N_33938);
or U34175 (N_34175,N_33975,N_33973);
and U34176 (N_34176,N_33068,N_33752);
xnor U34177 (N_34177,N_33500,N_33999);
nor U34178 (N_34178,N_33591,N_33598);
xor U34179 (N_34179,N_33564,N_33157);
nand U34180 (N_34180,N_33397,N_33666);
or U34181 (N_34181,N_33976,N_33425);
or U34182 (N_34182,N_33217,N_33555);
xor U34183 (N_34183,N_33499,N_33362);
nand U34184 (N_34184,N_33739,N_33671);
xnor U34185 (N_34185,N_33985,N_33576);
and U34186 (N_34186,N_33804,N_33203);
nor U34187 (N_34187,N_33053,N_33124);
nand U34188 (N_34188,N_33742,N_33401);
nor U34189 (N_34189,N_33332,N_33942);
and U34190 (N_34190,N_33016,N_33810);
or U34191 (N_34191,N_33896,N_33105);
nor U34192 (N_34192,N_33584,N_33771);
nand U34193 (N_34193,N_33573,N_33148);
nor U34194 (N_34194,N_33361,N_33954);
nand U34195 (N_34195,N_33903,N_33455);
xor U34196 (N_34196,N_33872,N_33071);
nor U34197 (N_34197,N_33781,N_33702);
xnor U34198 (N_34198,N_33007,N_33063);
and U34199 (N_34199,N_33290,N_33901);
xnor U34200 (N_34200,N_33239,N_33286);
or U34201 (N_34201,N_33535,N_33748);
nor U34202 (N_34202,N_33298,N_33984);
nor U34203 (N_34203,N_33663,N_33161);
xor U34204 (N_34204,N_33549,N_33185);
nor U34205 (N_34205,N_33626,N_33017);
nand U34206 (N_34206,N_33907,N_33331);
and U34207 (N_34207,N_33158,N_33837);
nor U34208 (N_34208,N_33289,N_33038);
nand U34209 (N_34209,N_33987,N_33556);
xor U34210 (N_34210,N_33369,N_33613);
nand U34211 (N_34211,N_33333,N_33466);
nor U34212 (N_34212,N_33252,N_33957);
or U34213 (N_34213,N_33219,N_33661);
xnor U34214 (N_34214,N_33279,N_33807);
and U34215 (N_34215,N_33390,N_33210);
nor U34216 (N_34216,N_33145,N_33140);
xnor U34217 (N_34217,N_33426,N_33974);
or U34218 (N_34218,N_33765,N_33539);
and U34219 (N_34219,N_33979,N_33523);
and U34220 (N_34220,N_33101,N_33821);
or U34221 (N_34221,N_33487,N_33039);
and U34222 (N_34222,N_33667,N_33776);
xnor U34223 (N_34223,N_33496,N_33617);
xnor U34224 (N_34224,N_33528,N_33577);
or U34225 (N_34225,N_33783,N_33020);
or U34226 (N_34226,N_33571,N_33747);
nand U34227 (N_34227,N_33314,N_33287);
nand U34228 (N_34228,N_33315,N_33880);
xor U34229 (N_34229,N_33580,N_33869);
xnor U34230 (N_34230,N_33868,N_33200);
nand U34231 (N_34231,N_33304,N_33019);
nand U34232 (N_34232,N_33302,N_33254);
and U34233 (N_34233,N_33495,N_33055);
and U34234 (N_34234,N_33511,N_33249);
xor U34235 (N_34235,N_33968,N_33534);
xor U34236 (N_34236,N_33592,N_33768);
nand U34237 (N_34237,N_33711,N_33754);
nand U34238 (N_34238,N_33346,N_33013);
nand U34239 (N_34239,N_33422,N_33554);
xnor U34240 (N_34240,N_33990,N_33127);
xnor U34241 (N_34241,N_33236,N_33852);
nor U34242 (N_34242,N_33376,N_33520);
xnor U34243 (N_34243,N_33048,N_33072);
nand U34244 (N_34244,N_33845,N_33625);
xnor U34245 (N_34245,N_33531,N_33165);
nor U34246 (N_34246,N_33493,N_33947);
or U34247 (N_34247,N_33202,N_33075);
xor U34248 (N_34248,N_33113,N_33788);
nand U34249 (N_34249,N_33174,N_33624);
nor U34250 (N_34250,N_33913,N_33553);
nand U34251 (N_34251,N_33138,N_33797);
and U34252 (N_34252,N_33473,N_33860);
or U34253 (N_34253,N_33838,N_33700);
xnor U34254 (N_34254,N_33522,N_33328);
or U34255 (N_34255,N_33032,N_33677);
or U34256 (N_34256,N_33420,N_33449);
nor U34257 (N_34257,N_33318,N_33620);
nand U34258 (N_34258,N_33833,N_33126);
or U34259 (N_34259,N_33418,N_33469);
xnor U34260 (N_34260,N_33463,N_33718);
nor U34261 (N_34261,N_33465,N_33034);
xor U34262 (N_34262,N_33778,N_33022);
and U34263 (N_34263,N_33503,N_33490);
xnor U34264 (N_34264,N_33103,N_33692);
nand U34265 (N_34265,N_33693,N_33672);
and U34266 (N_34266,N_33853,N_33741);
nand U34267 (N_34267,N_33740,N_33658);
and U34268 (N_34268,N_33266,N_33726);
nand U34269 (N_34269,N_33521,N_33118);
xor U34270 (N_34270,N_33884,N_33502);
xor U34271 (N_34271,N_33042,N_33295);
nand U34272 (N_34272,N_33173,N_33510);
and U34273 (N_34273,N_33306,N_33878);
xor U34274 (N_34274,N_33877,N_33237);
and U34275 (N_34275,N_33135,N_33762);
nand U34276 (N_34276,N_33568,N_33934);
xnor U34277 (N_34277,N_33587,N_33187);
nand U34278 (N_34278,N_33303,N_33710);
nand U34279 (N_34279,N_33077,N_33674);
or U34280 (N_34280,N_33259,N_33044);
nand U34281 (N_34281,N_33636,N_33770);
nor U34282 (N_34282,N_33861,N_33527);
nand U34283 (N_34283,N_33714,N_33801);
xor U34284 (N_34284,N_33052,N_33114);
or U34285 (N_34285,N_33247,N_33600);
nor U34286 (N_34286,N_33231,N_33367);
or U34287 (N_34287,N_33644,N_33107);
xor U34288 (N_34288,N_33952,N_33396);
and U34289 (N_34289,N_33316,N_33507);
and U34290 (N_34290,N_33257,N_33474);
xor U34291 (N_34291,N_33763,N_33312);
xnor U34292 (N_34292,N_33920,N_33794);
and U34293 (N_34293,N_33640,N_33526);
and U34294 (N_34294,N_33338,N_33737);
and U34295 (N_34295,N_33136,N_33958);
nor U34296 (N_34296,N_33542,N_33123);
and U34297 (N_34297,N_33698,N_33980);
nand U34298 (N_34298,N_33630,N_33981);
and U34299 (N_34299,N_33504,N_33102);
nand U34300 (N_34300,N_33978,N_33948);
xor U34301 (N_34301,N_33163,N_33246);
nor U34302 (N_34302,N_33995,N_33026);
or U34303 (N_34303,N_33240,N_33402);
or U34304 (N_34304,N_33767,N_33384);
and U34305 (N_34305,N_33326,N_33716);
xnor U34306 (N_34306,N_33371,N_33074);
nor U34307 (N_34307,N_33817,N_33594);
nor U34308 (N_34308,N_33021,N_33660);
nor U34309 (N_34309,N_33388,N_33603);
nand U34310 (N_34310,N_33307,N_33910);
nor U34311 (N_34311,N_33758,N_33632);
xor U34312 (N_34312,N_33269,N_33753);
nor U34313 (N_34313,N_33058,N_33450);
nor U34314 (N_34314,N_33645,N_33428);
and U34315 (N_34315,N_33615,N_33146);
xnor U34316 (N_34316,N_33356,N_33176);
and U34317 (N_34317,N_33363,N_33680);
nor U34318 (N_34318,N_33092,N_33380);
nand U34319 (N_34319,N_33207,N_33998);
and U34320 (N_34320,N_33873,N_33152);
or U34321 (N_34321,N_33530,N_33241);
xnor U34322 (N_34322,N_33191,N_33648);
xnor U34323 (N_34323,N_33412,N_33497);
nand U34324 (N_34324,N_33133,N_33228);
nor U34325 (N_34325,N_33593,N_33341);
nand U34326 (N_34326,N_33235,N_33789);
nor U34327 (N_34327,N_33357,N_33932);
nand U34328 (N_34328,N_33002,N_33410);
nor U34329 (N_34329,N_33966,N_33062);
or U34330 (N_34330,N_33844,N_33890);
nor U34331 (N_34331,N_33669,N_33803);
or U34332 (N_34332,N_33281,N_33399);
nor U34333 (N_34333,N_33162,N_33386);
nand U34334 (N_34334,N_33622,N_33154);
nor U34335 (N_34335,N_33040,N_33035);
or U34336 (N_34336,N_33993,N_33850);
nand U34337 (N_34337,N_33095,N_33863);
xnor U34338 (N_34338,N_33482,N_33432);
nand U34339 (N_34339,N_33442,N_33441);
nor U34340 (N_34340,N_33647,N_33633);
nor U34341 (N_34341,N_33119,N_33893);
or U34342 (N_34342,N_33634,N_33679);
xnor U34343 (N_34343,N_33701,N_33638);
nor U34344 (N_34344,N_33347,N_33699);
xor U34345 (N_34345,N_33642,N_33440);
and U34346 (N_34346,N_33265,N_33665);
nand U34347 (N_34347,N_33414,N_33245);
nor U34348 (N_34348,N_33166,N_33856);
and U34349 (N_34349,N_33732,N_33618);
nand U34350 (N_34350,N_33906,N_33519);
or U34351 (N_34351,N_33489,N_33282);
and U34352 (N_34352,N_33959,N_33311);
and U34353 (N_34353,N_33912,N_33351);
nand U34354 (N_34354,N_33570,N_33823);
and U34355 (N_34355,N_33536,N_33348);
nor U34356 (N_34356,N_33268,N_33253);
nand U34357 (N_34357,N_33713,N_33049);
nand U34358 (N_34358,N_33777,N_33816);
or U34359 (N_34359,N_33004,N_33623);
xnor U34360 (N_34360,N_33589,N_33858);
nand U34361 (N_34361,N_33736,N_33949);
or U34362 (N_34362,N_33319,N_33111);
or U34363 (N_34363,N_33383,N_33251);
xor U34364 (N_34364,N_33082,N_33782);
and U34365 (N_34365,N_33100,N_33902);
nand U34366 (N_34366,N_33139,N_33809);
or U34367 (N_34367,N_33596,N_33854);
and U34368 (N_34368,N_33033,N_33761);
nand U34369 (N_34369,N_33545,N_33505);
nand U34370 (N_34370,N_33792,N_33278);
nor U34371 (N_34371,N_33843,N_33067);
nand U34372 (N_34372,N_33829,N_33064);
or U34373 (N_34373,N_33859,N_33552);
nand U34374 (N_34374,N_33743,N_33061);
xor U34375 (N_34375,N_33799,N_33738);
or U34376 (N_34376,N_33673,N_33883);
nor U34377 (N_34377,N_33313,N_33802);
nand U34378 (N_34378,N_33080,N_33887);
nand U34379 (N_34379,N_33378,N_33675);
nor U34380 (N_34380,N_33656,N_33317);
nand U34381 (N_34381,N_33720,N_33694);
nand U34382 (N_34382,N_33590,N_33619);
xor U34383 (N_34383,N_33899,N_33501);
xnor U34384 (N_34384,N_33696,N_33218);
nor U34385 (N_34385,N_33336,N_33182);
xor U34386 (N_34386,N_33471,N_33201);
nor U34387 (N_34387,N_33848,N_33479);
nand U34388 (N_34388,N_33345,N_33977);
nand U34389 (N_34389,N_33206,N_33567);
nor U34390 (N_34390,N_33970,N_33417);
xnor U34391 (N_34391,N_33759,N_33989);
and U34392 (N_34392,N_33115,N_33808);
nor U34393 (N_34393,N_33891,N_33581);
nand U34394 (N_34394,N_33379,N_33391);
or U34395 (N_34395,N_33230,N_33373);
and U34396 (N_34396,N_33242,N_33757);
or U34397 (N_34397,N_33233,N_33457);
nor U34398 (N_34398,N_33043,N_33427);
xnor U34399 (N_34399,N_33172,N_33828);
nor U34400 (N_34400,N_33179,N_33725);
xor U34401 (N_34401,N_33144,N_33320);
nand U34402 (N_34402,N_33011,N_33586);
nand U34403 (N_34403,N_33790,N_33831);
nand U34404 (N_34404,N_33909,N_33309);
nor U34405 (N_34405,N_33324,N_33508);
and U34406 (N_34406,N_33769,N_33704);
and U34407 (N_34407,N_33484,N_33377);
and U34408 (N_34408,N_33867,N_33227);
xnor U34409 (N_34409,N_33815,N_33664);
and U34410 (N_34410,N_33557,N_33141);
or U34411 (N_34411,N_33394,N_33546);
or U34412 (N_34412,N_33305,N_33967);
or U34413 (N_34413,N_33682,N_33248);
xnor U34414 (N_34414,N_33690,N_33005);
xnor U34415 (N_34415,N_33170,N_33986);
and U34416 (N_34416,N_33171,N_33775);
nand U34417 (N_34417,N_33209,N_33079);
and U34418 (N_34418,N_33090,N_33651);
and U34419 (N_34419,N_33812,N_33547);
xnor U34420 (N_34420,N_33190,N_33773);
xor U34421 (N_34421,N_33785,N_33825);
nand U34422 (N_34422,N_33468,N_33597);
nand U34423 (N_34423,N_33533,N_33935);
and U34424 (N_34424,N_33116,N_33277);
nand U34425 (N_34425,N_33275,N_33216);
nand U34426 (N_34426,N_33188,N_33930);
or U34427 (N_34427,N_33685,N_33344);
nand U34428 (N_34428,N_33498,N_33084);
and U34429 (N_34429,N_33727,N_33806);
nand U34430 (N_34430,N_33919,N_33485);
nand U34431 (N_34431,N_33953,N_33296);
or U34432 (N_34432,N_33607,N_33922);
nor U34433 (N_34433,N_33153,N_33445);
or U34434 (N_34434,N_33840,N_33572);
xnor U34435 (N_34435,N_33543,N_33595);
or U34436 (N_34436,N_33180,N_33892);
xnor U34437 (N_34437,N_33925,N_33857);
nand U34438 (N_34438,N_33678,N_33321);
nor U34439 (N_34439,N_33421,N_33189);
xnor U34440 (N_34440,N_33506,N_33784);
or U34441 (N_34441,N_33609,N_33820);
xor U34442 (N_34442,N_33800,N_33488);
nand U34443 (N_34443,N_33524,N_33708);
or U34444 (N_34444,N_33429,N_33143);
xor U34445 (N_34445,N_33750,N_33294);
and U34446 (N_34446,N_33847,N_33460);
and U34447 (N_34447,N_33945,N_33657);
nand U34448 (N_34448,N_33267,N_33069);
nand U34449 (N_34449,N_33192,N_33452);
nand U34450 (N_34450,N_33608,N_33885);
and U34451 (N_34451,N_33937,N_33300);
nand U34452 (N_34452,N_33194,N_33224);
or U34453 (N_34453,N_33358,N_33214);
nor U34454 (N_34454,N_33112,N_33108);
xnor U34455 (N_34455,N_33365,N_33323);
nor U34456 (N_34456,N_33310,N_33627);
xor U34457 (N_34457,N_33014,N_33029);
xnor U34458 (N_34458,N_33492,N_33997);
xor U34459 (N_34459,N_33851,N_33322);
nor U34460 (N_34460,N_33923,N_33400);
nor U34461 (N_34461,N_33261,N_33056);
nor U34462 (N_34462,N_33096,N_33120);
or U34463 (N_34463,N_33226,N_33389);
and U34464 (N_34464,N_33003,N_33164);
nand U34465 (N_34465,N_33735,N_33955);
nand U34466 (N_34466,N_33670,N_33681);
nand U34467 (N_34467,N_33078,N_33073);
xor U34468 (N_34468,N_33220,N_33129);
nor U34469 (N_34469,N_33578,N_33340);
or U34470 (N_34470,N_33689,N_33779);
and U34471 (N_34471,N_33914,N_33695);
nor U34472 (N_34472,N_33409,N_33349);
or U34473 (N_34473,N_33070,N_33110);
or U34474 (N_34474,N_33709,N_33446);
nand U34475 (N_34475,N_33099,N_33059);
nand U34476 (N_34476,N_33065,N_33223);
nor U34477 (N_34477,N_33928,N_33437);
nand U34478 (N_34478,N_33722,N_33960);
or U34479 (N_34479,N_33606,N_33635);
or U34480 (N_34480,N_33330,N_33569);
nand U34481 (N_34481,N_33405,N_33438);
nor U34482 (N_34482,N_33212,N_33462);
xor U34483 (N_34483,N_33706,N_33839);
and U34484 (N_34484,N_33255,N_33724);
and U34485 (N_34485,N_33969,N_33046);
xor U34486 (N_34486,N_33605,N_33723);
and U34487 (N_34487,N_33566,N_33382);
nand U34488 (N_34488,N_33683,N_33905);
and U34489 (N_34489,N_33532,N_33728);
and U34490 (N_34490,N_33085,N_33760);
xnor U34491 (N_34491,N_33876,N_33818);
or U34492 (N_34492,N_33443,N_33284);
xor U34493 (N_34493,N_33814,N_33415);
or U34494 (N_34494,N_33886,N_33225);
nor U34495 (N_34495,N_33793,N_33385);
or U34496 (N_34496,N_33916,N_33961);
or U34497 (N_34497,N_33780,N_33734);
or U34498 (N_34498,N_33423,N_33301);
and U34499 (N_34499,N_33028,N_33924);
xor U34500 (N_34500,N_33078,N_33859);
nor U34501 (N_34501,N_33009,N_33539);
xor U34502 (N_34502,N_33316,N_33180);
nor U34503 (N_34503,N_33158,N_33940);
nand U34504 (N_34504,N_33908,N_33313);
and U34505 (N_34505,N_33530,N_33657);
or U34506 (N_34506,N_33095,N_33671);
or U34507 (N_34507,N_33822,N_33087);
nand U34508 (N_34508,N_33845,N_33564);
xnor U34509 (N_34509,N_33785,N_33675);
nand U34510 (N_34510,N_33356,N_33753);
or U34511 (N_34511,N_33102,N_33157);
nor U34512 (N_34512,N_33771,N_33053);
xor U34513 (N_34513,N_33309,N_33665);
or U34514 (N_34514,N_33368,N_33828);
or U34515 (N_34515,N_33283,N_33418);
nor U34516 (N_34516,N_33190,N_33845);
or U34517 (N_34517,N_33261,N_33778);
nor U34518 (N_34518,N_33112,N_33582);
nand U34519 (N_34519,N_33358,N_33368);
or U34520 (N_34520,N_33102,N_33154);
nand U34521 (N_34521,N_33942,N_33124);
xor U34522 (N_34522,N_33195,N_33991);
nand U34523 (N_34523,N_33060,N_33597);
nor U34524 (N_34524,N_33289,N_33890);
nand U34525 (N_34525,N_33849,N_33269);
nand U34526 (N_34526,N_33393,N_33777);
nand U34527 (N_34527,N_33596,N_33673);
nor U34528 (N_34528,N_33736,N_33143);
xor U34529 (N_34529,N_33496,N_33823);
and U34530 (N_34530,N_33521,N_33190);
nor U34531 (N_34531,N_33187,N_33361);
or U34532 (N_34532,N_33992,N_33429);
xor U34533 (N_34533,N_33210,N_33140);
and U34534 (N_34534,N_33246,N_33289);
nor U34535 (N_34535,N_33033,N_33383);
and U34536 (N_34536,N_33108,N_33974);
xnor U34537 (N_34537,N_33607,N_33725);
nand U34538 (N_34538,N_33633,N_33352);
xor U34539 (N_34539,N_33437,N_33628);
nand U34540 (N_34540,N_33281,N_33961);
or U34541 (N_34541,N_33788,N_33696);
and U34542 (N_34542,N_33004,N_33213);
xnor U34543 (N_34543,N_33667,N_33443);
or U34544 (N_34544,N_33390,N_33774);
xnor U34545 (N_34545,N_33725,N_33321);
or U34546 (N_34546,N_33359,N_33154);
xor U34547 (N_34547,N_33240,N_33431);
nor U34548 (N_34548,N_33088,N_33887);
and U34549 (N_34549,N_33068,N_33547);
xnor U34550 (N_34550,N_33922,N_33985);
nand U34551 (N_34551,N_33216,N_33806);
nor U34552 (N_34552,N_33500,N_33558);
and U34553 (N_34553,N_33098,N_33646);
and U34554 (N_34554,N_33975,N_33086);
nand U34555 (N_34555,N_33790,N_33819);
xor U34556 (N_34556,N_33565,N_33307);
and U34557 (N_34557,N_33110,N_33297);
xnor U34558 (N_34558,N_33520,N_33176);
nand U34559 (N_34559,N_33532,N_33398);
xor U34560 (N_34560,N_33022,N_33298);
nand U34561 (N_34561,N_33017,N_33185);
nand U34562 (N_34562,N_33617,N_33346);
nand U34563 (N_34563,N_33617,N_33671);
or U34564 (N_34564,N_33813,N_33680);
xor U34565 (N_34565,N_33261,N_33465);
xnor U34566 (N_34566,N_33833,N_33685);
nand U34567 (N_34567,N_33253,N_33215);
nor U34568 (N_34568,N_33508,N_33372);
nand U34569 (N_34569,N_33184,N_33955);
xnor U34570 (N_34570,N_33904,N_33962);
xor U34571 (N_34571,N_33646,N_33975);
xnor U34572 (N_34572,N_33181,N_33643);
nand U34573 (N_34573,N_33933,N_33831);
nor U34574 (N_34574,N_33994,N_33421);
nand U34575 (N_34575,N_33698,N_33926);
and U34576 (N_34576,N_33396,N_33311);
or U34577 (N_34577,N_33064,N_33408);
xnor U34578 (N_34578,N_33414,N_33843);
and U34579 (N_34579,N_33087,N_33652);
xor U34580 (N_34580,N_33125,N_33363);
or U34581 (N_34581,N_33100,N_33805);
nand U34582 (N_34582,N_33934,N_33750);
nor U34583 (N_34583,N_33247,N_33432);
nand U34584 (N_34584,N_33360,N_33086);
and U34585 (N_34585,N_33009,N_33112);
or U34586 (N_34586,N_33091,N_33999);
or U34587 (N_34587,N_33180,N_33612);
nor U34588 (N_34588,N_33060,N_33502);
and U34589 (N_34589,N_33776,N_33918);
xor U34590 (N_34590,N_33128,N_33591);
nor U34591 (N_34591,N_33415,N_33578);
nand U34592 (N_34592,N_33082,N_33187);
or U34593 (N_34593,N_33683,N_33812);
nand U34594 (N_34594,N_33911,N_33357);
nor U34595 (N_34595,N_33163,N_33073);
and U34596 (N_34596,N_33524,N_33926);
nand U34597 (N_34597,N_33282,N_33958);
or U34598 (N_34598,N_33432,N_33525);
nor U34599 (N_34599,N_33374,N_33848);
and U34600 (N_34600,N_33997,N_33125);
nand U34601 (N_34601,N_33494,N_33142);
nor U34602 (N_34602,N_33414,N_33573);
nor U34603 (N_34603,N_33041,N_33417);
nor U34604 (N_34604,N_33152,N_33429);
nor U34605 (N_34605,N_33158,N_33981);
nor U34606 (N_34606,N_33868,N_33603);
nor U34607 (N_34607,N_33119,N_33676);
or U34608 (N_34608,N_33918,N_33915);
xnor U34609 (N_34609,N_33917,N_33721);
or U34610 (N_34610,N_33009,N_33399);
nor U34611 (N_34611,N_33146,N_33080);
or U34612 (N_34612,N_33863,N_33402);
nand U34613 (N_34613,N_33746,N_33730);
and U34614 (N_34614,N_33471,N_33525);
nor U34615 (N_34615,N_33366,N_33827);
or U34616 (N_34616,N_33452,N_33754);
nor U34617 (N_34617,N_33563,N_33562);
nand U34618 (N_34618,N_33032,N_33911);
xor U34619 (N_34619,N_33669,N_33724);
or U34620 (N_34620,N_33919,N_33042);
nand U34621 (N_34621,N_33727,N_33367);
xnor U34622 (N_34622,N_33674,N_33113);
or U34623 (N_34623,N_33642,N_33861);
or U34624 (N_34624,N_33991,N_33521);
nand U34625 (N_34625,N_33370,N_33201);
or U34626 (N_34626,N_33461,N_33389);
xor U34627 (N_34627,N_33752,N_33403);
nor U34628 (N_34628,N_33818,N_33450);
nand U34629 (N_34629,N_33706,N_33229);
xnor U34630 (N_34630,N_33707,N_33556);
or U34631 (N_34631,N_33058,N_33164);
nor U34632 (N_34632,N_33118,N_33409);
xnor U34633 (N_34633,N_33831,N_33532);
nand U34634 (N_34634,N_33349,N_33597);
and U34635 (N_34635,N_33368,N_33497);
xor U34636 (N_34636,N_33787,N_33034);
or U34637 (N_34637,N_33387,N_33573);
xnor U34638 (N_34638,N_33153,N_33904);
nor U34639 (N_34639,N_33623,N_33497);
nand U34640 (N_34640,N_33228,N_33045);
xnor U34641 (N_34641,N_33224,N_33003);
nand U34642 (N_34642,N_33987,N_33711);
nand U34643 (N_34643,N_33593,N_33229);
or U34644 (N_34644,N_33913,N_33759);
nand U34645 (N_34645,N_33594,N_33960);
xor U34646 (N_34646,N_33964,N_33304);
nand U34647 (N_34647,N_33635,N_33057);
xnor U34648 (N_34648,N_33247,N_33672);
xnor U34649 (N_34649,N_33279,N_33981);
or U34650 (N_34650,N_33491,N_33911);
xor U34651 (N_34651,N_33249,N_33018);
and U34652 (N_34652,N_33649,N_33776);
or U34653 (N_34653,N_33622,N_33760);
xnor U34654 (N_34654,N_33555,N_33742);
nor U34655 (N_34655,N_33902,N_33275);
xor U34656 (N_34656,N_33069,N_33940);
or U34657 (N_34657,N_33737,N_33211);
xnor U34658 (N_34658,N_33501,N_33965);
xnor U34659 (N_34659,N_33538,N_33478);
nor U34660 (N_34660,N_33351,N_33475);
nor U34661 (N_34661,N_33760,N_33063);
or U34662 (N_34662,N_33543,N_33431);
nand U34663 (N_34663,N_33167,N_33070);
nand U34664 (N_34664,N_33527,N_33187);
or U34665 (N_34665,N_33698,N_33934);
nor U34666 (N_34666,N_33490,N_33279);
or U34667 (N_34667,N_33537,N_33366);
or U34668 (N_34668,N_33864,N_33222);
nor U34669 (N_34669,N_33764,N_33530);
nand U34670 (N_34670,N_33074,N_33544);
or U34671 (N_34671,N_33447,N_33573);
nor U34672 (N_34672,N_33070,N_33844);
and U34673 (N_34673,N_33577,N_33248);
or U34674 (N_34674,N_33412,N_33301);
nor U34675 (N_34675,N_33447,N_33916);
and U34676 (N_34676,N_33700,N_33944);
nor U34677 (N_34677,N_33625,N_33926);
nor U34678 (N_34678,N_33809,N_33864);
xnor U34679 (N_34679,N_33581,N_33726);
or U34680 (N_34680,N_33131,N_33453);
and U34681 (N_34681,N_33285,N_33372);
and U34682 (N_34682,N_33645,N_33687);
xor U34683 (N_34683,N_33454,N_33353);
and U34684 (N_34684,N_33140,N_33035);
nand U34685 (N_34685,N_33834,N_33822);
nand U34686 (N_34686,N_33177,N_33639);
nand U34687 (N_34687,N_33323,N_33576);
nand U34688 (N_34688,N_33413,N_33712);
and U34689 (N_34689,N_33472,N_33619);
and U34690 (N_34690,N_33165,N_33124);
nand U34691 (N_34691,N_33628,N_33644);
xnor U34692 (N_34692,N_33015,N_33811);
or U34693 (N_34693,N_33149,N_33301);
nor U34694 (N_34694,N_33332,N_33718);
xor U34695 (N_34695,N_33079,N_33163);
and U34696 (N_34696,N_33148,N_33850);
nand U34697 (N_34697,N_33864,N_33909);
xnor U34698 (N_34698,N_33784,N_33314);
or U34699 (N_34699,N_33409,N_33079);
xnor U34700 (N_34700,N_33163,N_33997);
nor U34701 (N_34701,N_33260,N_33253);
and U34702 (N_34702,N_33060,N_33133);
nor U34703 (N_34703,N_33578,N_33700);
nand U34704 (N_34704,N_33256,N_33228);
nor U34705 (N_34705,N_33681,N_33062);
xor U34706 (N_34706,N_33867,N_33150);
nand U34707 (N_34707,N_33023,N_33320);
or U34708 (N_34708,N_33765,N_33713);
nor U34709 (N_34709,N_33650,N_33382);
or U34710 (N_34710,N_33776,N_33088);
nand U34711 (N_34711,N_33574,N_33097);
and U34712 (N_34712,N_33630,N_33934);
or U34713 (N_34713,N_33572,N_33730);
nand U34714 (N_34714,N_33419,N_33678);
nand U34715 (N_34715,N_33522,N_33947);
nor U34716 (N_34716,N_33393,N_33970);
or U34717 (N_34717,N_33178,N_33846);
or U34718 (N_34718,N_33788,N_33496);
nand U34719 (N_34719,N_33707,N_33143);
or U34720 (N_34720,N_33391,N_33764);
and U34721 (N_34721,N_33988,N_33821);
xnor U34722 (N_34722,N_33723,N_33209);
or U34723 (N_34723,N_33497,N_33688);
or U34724 (N_34724,N_33712,N_33119);
nand U34725 (N_34725,N_33638,N_33750);
nor U34726 (N_34726,N_33575,N_33627);
nor U34727 (N_34727,N_33848,N_33866);
or U34728 (N_34728,N_33611,N_33665);
or U34729 (N_34729,N_33166,N_33958);
or U34730 (N_34730,N_33106,N_33201);
xnor U34731 (N_34731,N_33586,N_33064);
nand U34732 (N_34732,N_33612,N_33831);
or U34733 (N_34733,N_33716,N_33704);
nor U34734 (N_34734,N_33306,N_33164);
xnor U34735 (N_34735,N_33416,N_33379);
and U34736 (N_34736,N_33543,N_33063);
or U34737 (N_34737,N_33191,N_33529);
nand U34738 (N_34738,N_33520,N_33239);
xor U34739 (N_34739,N_33938,N_33102);
nor U34740 (N_34740,N_33742,N_33606);
nand U34741 (N_34741,N_33455,N_33171);
and U34742 (N_34742,N_33578,N_33576);
nand U34743 (N_34743,N_33094,N_33305);
nor U34744 (N_34744,N_33396,N_33684);
xor U34745 (N_34745,N_33790,N_33766);
and U34746 (N_34746,N_33552,N_33064);
and U34747 (N_34747,N_33811,N_33751);
or U34748 (N_34748,N_33704,N_33901);
xnor U34749 (N_34749,N_33635,N_33540);
nand U34750 (N_34750,N_33166,N_33211);
nor U34751 (N_34751,N_33950,N_33960);
or U34752 (N_34752,N_33959,N_33168);
or U34753 (N_34753,N_33236,N_33004);
nand U34754 (N_34754,N_33909,N_33291);
xor U34755 (N_34755,N_33229,N_33267);
and U34756 (N_34756,N_33545,N_33821);
and U34757 (N_34757,N_33517,N_33537);
xor U34758 (N_34758,N_33483,N_33106);
nor U34759 (N_34759,N_33263,N_33957);
xor U34760 (N_34760,N_33084,N_33671);
xor U34761 (N_34761,N_33335,N_33331);
nand U34762 (N_34762,N_33844,N_33271);
nand U34763 (N_34763,N_33299,N_33926);
or U34764 (N_34764,N_33649,N_33204);
xor U34765 (N_34765,N_33153,N_33494);
and U34766 (N_34766,N_33031,N_33097);
nor U34767 (N_34767,N_33859,N_33886);
nand U34768 (N_34768,N_33054,N_33081);
nand U34769 (N_34769,N_33308,N_33795);
nor U34770 (N_34770,N_33013,N_33218);
or U34771 (N_34771,N_33767,N_33010);
xor U34772 (N_34772,N_33602,N_33089);
xor U34773 (N_34773,N_33737,N_33018);
or U34774 (N_34774,N_33539,N_33114);
xnor U34775 (N_34775,N_33201,N_33553);
nand U34776 (N_34776,N_33854,N_33821);
or U34777 (N_34777,N_33803,N_33326);
and U34778 (N_34778,N_33723,N_33642);
nand U34779 (N_34779,N_33183,N_33874);
and U34780 (N_34780,N_33896,N_33223);
nor U34781 (N_34781,N_33379,N_33323);
and U34782 (N_34782,N_33009,N_33232);
nand U34783 (N_34783,N_33033,N_33742);
nand U34784 (N_34784,N_33949,N_33087);
and U34785 (N_34785,N_33858,N_33021);
and U34786 (N_34786,N_33188,N_33652);
or U34787 (N_34787,N_33789,N_33362);
xor U34788 (N_34788,N_33521,N_33172);
or U34789 (N_34789,N_33429,N_33972);
and U34790 (N_34790,N_33138,N_33173);
or U34791 (N_34791,N_33346,N_33685);
nand U34792 (N_34792,N_33222,N_33003);
and U34793 (N_34793,N_33632,N_33249);
and U34794 (N_34794,N_33622,N_33143);
nor U34795 (N_34795,N_33212,N_33011);
nand U34796 (N_34796,N_33864,N_33517);
or U34797 (N_34797,N_33877,N_33324);
or U34798 (N_34798,N_33797,N_33323);
and U34799 (N_34799,N_33789,N_33493);
xor U34800 (N_34800,N_33223,N_33441);
nor U34801 (N_34801,N_33605,N_33128);
nor U34802 (N_34802,N_33719,N_33658);
nor U34803 (N_34803,N_33334,N_33645);
xor U34804 (N_34804,N_33292,N_33306);
and U34805 (N_34805,N_33617,N_33521);
and U34806 (N_34806,N_33416,N_33493);
and U34807 (N_34807,N_33864,N_33407);
and U34808 (N_34808,N_33444,N_33008);
or U34809 (N_34809,N_33021,N_33801);
nand U34810 (N_34810,N_33001,N_33713);
or U34811 (N_34811,N_33724,N_33541);
and U34812 (N_34812,N_33441,N_33262);
xor U34813 (N_34813,N_33172,N_33474);
nor U34814 (N_34814,N_33063,N_33811);
or U34815 (N_34815,N_33207,N_33906);
nand U34816 (N_34816,N_33728,N_33430);
and U34817 (N_34817,N_33285,N_33716);
nor U34818 (N_34818,N_33346,N_33365);
or U34819 (N_34819,N_33908,N_33911);
or U34820 (N_34820,N_33847,N_33346);
xnor U34821 (N_34821,N_33910,N_33082);
or U34822 (N_34822,N_33896,N_33064);
nand U34823 (N_34823,N_33316,N_33089);
xnor U34824 (N_34824,N_33810,N_33614);
xor U34825 (N_34825,N_33353,N_33905);
nand U34826 (N_34826,N_33494,N_33787);
and U34827 (N_34827,N_33917,N_33664);
nand U34828 (N_34828,N_33776,N_33350);
nand U34829 (N_34829,N_33028,N_33180);
xnor U34830 (N_34830,N_33354,N_33826);
xnor U34831 (N_34831,N_33518,N_33376);
xnor U34832 (N_34832,N_33619,N_33764);
nor U34833 (N_34833,N_33125,N_33418);
or U34834 (N_34834,N_33554,N_33398);
nand U34835 (N_34835,N_33605,N_33047);
nand U34836 (N_34836,N_33740,N_33898);
or U34837 (N_34837,N_33752,N_33746);
nand U34838 (N_34838,N_33317,N_33602);
and U34839 (N_34839,N_33013,N_33947);
nor U34840 (N_34840,N_33208,N_33003);
or U34841 (N_34841,N_33931,N_33423);
xor U34842 (N_34842,N_33615,N_33570);
and U34843 (N_34843,N_33831,N_33311);
or U34844 (N_34844,N_33912,N_33706);
nor U34845 (N_34845,N_33440,N_33496);
xnor U34846 (N_34846,N_33362,N_33033);
nor U34847 (N_34847,N_33014,N_33593);
or U34848 (N_34848,N_33735,N_33450);
xnor U34849 (N_34849,N_33961,N_33789);
nor U34850 (N_34850,N_33667,N_33213);
nor U34851 (N_34851,N_33578,N_33617);
nand U34852 (N_34852,N_33068,N_33869);
nand U34853 (N_34853,N_33477,N_33038);
or U34854 (N_34854,N_33000,N_33983);
and U34855 (N_34855,N_33492,N_33014);
and U34856 (N_34856,N_33560,N_33010);
nor U34857 (N_34857,N_33240,N_33610);
and U34858 (N_34858,N_33713,N_33743);
xnor U34859 (N_34859,N_33399,N_33177);
and U34860 (N_34860,N_33797,N_33960);
xor U34861 (N_34861,N_33653,N_33765);
nor U34862 (N_34862,N_33067,N_33871);
nand U34863 (N_34863,N_33191,N_33201);
xnor U34864 (N_34864,N_33375,N_33861);
nor U34865 (N_34865,N_33589,N_33779);
and U34866 (N_34866,N_33652,N_33531);
nand U34867 (N_34867,N_33744,N_33317);
xnor U34868 (N_34868,N_33253,N_33094);
nor U34869 (N_34869,N_33881,N_33058);
nor U34870 (N_34870,N_33590,N_33832);
nor U34871 (N_34871,N_33236,N_33279);
xor U34872 (N_34872,N_33078,N_33962);
and U34873 (N_34873,N_33494,N_33468);
and U34874 (N_34874,N_33896,N_33360);
nand U34875 (N_34875,N_33833,N_33626);
nand U34876 (N_34876,N_33348,N_33137);
nor U34877 (N_34877,N_33162,N_33280);
or U34878 (N_34878,N_33109,N_33499);
nand U34879 (N_34879,N_33103,N_33541);
or U34880 (N_34880,N_33216,N_33622);
nand U34881 (N_34881,N_33403,N_33311);
and U34882 (N_34882,N_33398,N_33004);
nand U34883 (N_34883,N_33312,N_33243);
nand U34884 (N_34884,N_33418,N_33849);
nand U34885 (N_34885,N_33597,N_33592);
xor U34886 (N_34886,N_33302,N_33115);
and U34887 (N_34887,N_33903,N_33229);
nand U34888 (N_34888,N_33403,N_33654);
nor U34889 (N_34889,N_33668,N_33317);
or U34890 (N_34890,N_33934,N_33457);
nor U34891 (N_34891,N_33714,N_33750);
nor U34892 (N_34892,N_33560,N_33123);
nand U34893 (N_34893,N_33954,N_33739);
nand U34894 (N_34894,N_33740,N_33453);
and U34895 (N_34895,N_33495,N_33284);
xnor U34896 (N_34896,N_33557,N_33435);
nor U34897 (N_34897,N_33212,N_33102);
nor U34898 (N_34898,N_33263,N_33358);
and U34899 (N_34899,N_33450,N_33831);
or U34900 (N_34900,N_33322,N_33604);
nand U34901 (N_34901,N_33959,N_33717);
nand U34902 (N_34902,N_33918,N_33316);
nand U34903 (N_34903,N_33940,N_33064);
nor U34904 (N_34904,N_33005,N_33984);
and U34905 (N_34905,N_33071,N_33310);
nor U34906 (N_34906,N_33113,N_33810);
or U34907 (N_34907,N_33913,N_33459);
or U34908 (N_34908,N_33190,N_33125);
and U34909 (N_34909,N_33670,N_33748);
and U34910 (N_34910,N_33946,N_33491);
xnor U34911 (N_34911,N_33190,N_33013);
or U34912 (N_34912,N_33824,N_33198);
nor U34913 (N_34913,N_33456,N_33546);
xor U34914 (N_34914,N_33038,N_33048);
and U34915 (N_34915,N_33920,N_33091);
nand U34916 (N_34916,N_33890,N_33676);
and U34917 (N_34917,N_33492,N_33857);
or U34918 (N_34918,N_33148,N_33989);
nor U34919 (N_34919,N_33361,N_33038);
nand U34920 (N_34920,N_33631,N_33358);
xor U34921 (N_34921,N_33860,N_33650);
or U34922 (N_34922,N_33198,N_33622);
or U34923 (N_34923,N_33957,N_33258);
nor U34924 (N_34924,N_33362,N_33133);
xnor U34925 (N_34925,N_33459,N_33033);
nor U34926 (N_34926,N_33100,N_33634);
nand U34927 (N_34927,N_33402,N_33426);
and U34928 (N_34928,N_33182,N_33298);
xnor U34929 (N_34929,N_33777,N_33454);
nor U34930 (N_34930,N_33348,N_33341);
and U34931 (N_34931,N_33298,N_33734);
nand U34932 (N_34932,N_33356,N_33190);
and U34933 (N_34933,N_33948,N_33579);
nor U34934 (N_34934,N_33970,N_33165);
nor U34935 (N_34935,N_33984,N_33106);
and U34936 (N_34936,N_33482,N_33757);
nand U34937 (N_34937,N_33090,N_33991);
and U34938 (N_34938,N_33842,N_33411);
or U34939 (N_34939,N_33684,N_33632);
xor U34940 (N_34940,N_33929,N_33827);
xnor U34941 (N_34941,N_33070,N_33352);
nand U34942 (N_34942,N_33375,N_33410);
or U34943 (N_34943,N_33041,N_33665);
nor U34944 (N_34944,N_33469,N_33146);
nor U34945 (N_34945,N_33864,N_33503);
and U34946 (N_34946,N_33285,N_33605);
nor U34947 (N_34947,N_33557,N_33768);
or U34948 (N_34948,N_33190,N_33249);
nor U34949 (N_34949,N_33021,N_33865);
nor U34950 (N_34950,N_33048,N_33372);
and U34951 (N_34951,N_33014,N_33704);
nor U34952 (N_34952,N_33386,N_33079);
nand U34953 (N_34953,N_33510,N_33111);
nand U34954 (N_34954,N_33430,N_33673);
nor U34955 (N_34955,N_33401,N_33906);
nand U34956 (N_34956,N_33550,N_33899);
xnor U34957 (N_34957,N_33241,N_33136);
nand U34958 (N_34958,N_33487,N_33444);
or U34959 (N_34959,N_33931,N_33364);
nand U34960 (N_34960,N_33694,N_33821);
nand U34961 (N_34961,N_33933,N_33940);
and U34962 (N_34962,N_33963,N_33720);
or U34963 (N_34963,N_33237,N_33341);
and U34964 (N_34964,N_33376,N_33077);
nand U34965 (N_34965,N_33299,N_33001);
xor U34966 (N_34966,N_33844,N_33878);
xnor U34967 (N_34967,N_33553,N_33569);
or U34968 (N_34968,N_33261,N_33121);
xor U34969 (N_34969,N_33321,N_33016);
nor U34970 (N_34970,N_33399,N_33481);
nand U34971 (N_34971,N_33044,N_33616);
nor U34972 (N_34972,N_33340,N_33954);
nor U34973 (N_34973,N_33625,N_33492);
nand U34974 (N_34974,N_33792,N_33402);
nor U34975 (N_34975,N_33053,N_33166);
xnor U34976 (N_34976,N_33470,N_33409);
xor U34977 (N_34977,N_33276,N_33089);
nor U34978 (N_34978,N_33755,N_33407);
and U34979 (N_34979,N_33224,N_33736);
nand U34980 (N_34980,N_33607,N_33927);
nor U34981 (N_34981,N_33437,N_33527);
xnor U34982 (N_34982,N_33694,N_33483);
and U34983 (N_34983,N_33040,N_33395);
nand U34984 (N_34984,N_33316,N_33242);
nor U34985 (N_34985,N_33570,N_33125);
xor U34986 (N_34986,N_33043,N_33104);
or U34987 (N_34987,N_33101,N_33474);
xor U34988 (N_34988,N_33544,N_33902);
or U34989 (N_34989,N_33353,N_33703);
nor U34990 (N_34990,N_33654,N_33297);
xor U34991 (N_34991,N_33468,N_33230);
nand U34992 (N_34992,N_33449,N_33026);
nor U34993 (N_34993,N_33365,N_33012);
or U34994 (N_34994,N_33336,N_33594);
xnor U34995 (N_34995,N_33714,N_33560);
xnor U34996 (N_34996,N_33148,N_33426);
nor U34997 (N_34997,N_33311,N_33284);
nand U34998 (N_34998,N_33667,N_33391);
and U34999 (N_34999,N_33841,N_33354);
nand U35000 (N_35000,N_34156,N_34553);
xor U35001 (N_35001,N_34678,N_34082);
nor U35002 (N_35002,N_34196,N_34513);
or U35003 (N_35003,N_34387,N_34781);
or U35004 (N_35004,N_34654,N_34242);
or U35005 (N_35005,N_34042,N_34707);
xnor U35006 (N_35006,N_34577,N_34225);
or U35007 (N_35007,N_34580,N_34686);
xor U35008 (N_35008,N_34552,N_34471);
xor U35009 (N_35009,N_34323,N_34711);
and U35010 (N_35010,N_34232,N_34938);
nor U35011 (N_35011,N_34639,N_34438);
nand U35012 (N_35012,N_34987,N_34761);
and U35013 (N_35013,N_34192,N_34485);
or U35014 (N_35014,N_34853,N_34182);
nor U35015 (N_35015,N_34036,N_34754);
or U35016 (N_35016,N_34628,N_34330);
nor U35017 (N_35017,N_34619,N_34429);
and U35018 (N_35018,N_34501,N_34664);
nand U35019 (N_35019,N_34331,N_34335);
nand U35020 (N_35020,N_34772,N_34475);
xnor U35021 (N_35021,N_34727,N_34187);
and U35022 (N_35022,N_34883,N_34773);
nor U35023 (N_35023,N_34821,N_34329);
nor U35024 (N_35024,N_34464,N_34339);
nand U35025 (N_35025,N_34027,N_34663);
xor U35026 (N_35026,N_34923,N_34684);
nor U35027 (N_35027,N_34842,N_34794);
or U35028 (N_35028,N_34249,N_34836);
or U35029 (N_35029,N_34364,N_34197);
xor U35030 (N_35030,N_34290,N_34723);
nand U35031 (N_35031,N_34532,N_34109);
and U35032 (N_35032,N_34140,N_34291);
and U35033 (N_35033,N_34277,N_34827);
xnor U35034 (N_35034,N_34798,N_34385);
or U35035 (N_35035,N_34789,N_34714);
or U35036 (N_35036,N_34436,N_34159);
nand U35037 (N_35037,N_34598,N_34815);
nand U35038 (N_35038,N_34698,N_34076);
nand U35039 (N_35039,N_34776,N_34336);
and U35040 (N_35040,N_34944,N_34765);
and U35041 (N_35041,N_34165,N_34747);
nand U35042 (N_35042,N_34056,N_34763);
nor U35043 (N_35043,N_34072,N_34790);
and U35044 (N_35044,N_34869,N_34729);
xnor U35045 (N_35045,N_34832,N_34312);
nand U35046 (N_35046,N_34411,N_34541);
nand U35047 (N_35047,N_34749,N_34007);
and U35048 (N_35048,N_34468,N_34648);
xnor U35049 (N_35049,N_34680,N_34492);
or U35050 (N_35050,N_34049,N_34732);
xor U35051 (N_35051,N_34777,N_34131);
xnor U35052 (N_35052,N_34300,N_34612);
nand U35053 (N_35053,N_34644,N_34251);
or U35054 (N_35054,N_34181,N_34606);
nand U35055 (N_35055,N_34117,N_34637);
or U35056 (N_35056,N_34880,N_34284);
and U35057 (N_35057,N_34378,N_34063);
xor U35058 (N_35058,N_34615,N_34672);
nand U35059 (N_35059,N_34093,N_34751);
nor U35060 (N_35060,N_34488,N_34636);
nor U35061 (N_35061,N_34050,N_34122);
or U35062 (N_35062,N_34922,N_34124);
nor U35063 (N_35063,N_34793,N_34588);
nor U35064 (N_35064,N_34755,N_34914);
and U35065 (N_35065,N_34688,N_34893);
or U35066 (N_35066,N_34660,N_34014);
nor U35067 (N_35067,N_34595,N_34162);
or U35068 (N_35068,N_34040,N_34432);
nor U35069 (N_35069,N_34110,N_34956);
nor U35070 (N_35070,N_34209,N_34293);
and U35071 (N_35071,N_34877,N_34490);
xnor U35072 (N_35072,N_34795,N_34143);
nor U35073 (N_35073,N_34825,N_34902);
and U35074 (N_35074,N_34415,N_34961);
xor U35075 (N_35075,N_34292,N_34951);
or U35076 (N_35076,N_34417,N_34434);
or U35077 (N_35077,N_34622,N_34910);
xor U35078 (N_35078,N_34274,N_34788);
nand U35079 (N_35079,N_34246,N_34837);
and U35080 (N_35080,N_34942,N_34442);
or U35081 (N_35081,N_34955,N_34279);
nor U35082 (N_35082,N_34097,N_34351);
xnor U35083 (N_35083,N_34271,N_34889);
or U35084 (N_35084,N_34618,N_34972);
nand U35085 (N_35085,N_34431,N_34028);
nor U35086 (N_35086,N_34430,N_34587);
and U35087 (N_35087,N_34086,N_34753);
or U35088 (N_35088,N_34807,N_34183);
and U35089 (N_35089,N_34633,N_34486);
nor U35090 (N_35090,N_34210,N_34758);
nor U35091 (N_35091,N_34802,N_34400);
nand U35092 (N_35092,N_34689,N_34964);
and U35093 (N_35093,N_34326,N_34605);
xor U35094 (N_35094,N_34797,N_34787);
xnor U35095 (N_35095,N_34613,N_34157);
and U35096 (N_35096,N_34597,N_34084);
xnor U35097 (N_35097,N_34349,N_34937);
nand U35098 (N_35098,N_34523,N_34665);
or U35099 (N_35099,N_34362,N_34778);
or U35100 (N_35100,N_34898,N_34656);
or U35101 (N_35101,N_34693,N_34016);
nand U35102 (N_35102,N_34200,N_34748);
xor U35103 (N_35103,N_34382,N_34238);
or U35104 (N_35104,N_34670,N_34509);
and U35105 (N_35105,N_34325,N_34064);
or U35106 (N_35106,N_34283,N_34444);
and U35107 (N_35107,N_34575,N_34959);
nand U35108 (N_35108,N_34950,N_34104);
nor U35109 (N_35109,N_34224,N_34834);
xor U35110 (N_35110,N_34518,N_34854);
nor U35111 (N_35111,N_34258,N_34307);
xor U35112 (N_35112,N_34390,N_34929);
nor U35113 (N_35113,N_34551,N_34774);
and U35114 (N_35114,N_34590,N_34900);
nor U35115 (N_35115,N_34847,N_34879);
and U35116 (N_35116,N_34531,N_34055);
and U35117 (N_35117,N_34616,N_34180);
xor U35118 (N_35118,N_34596,N_34971);
nand U35119 (N_35119,N_34516,N_34739);
nand U35120 (N_35120,N_34736,N_34039);
xnor U35121 (N_35121,N_34495,N_34667);
nand U35122 (N_35122,N_34319,N_34303);
and U35123 (N_35123,N_34174,N_34918);
nor U35124 (N_35124,N_34463,N_34690);
xor U35125 (N_35125,N_34999,N_34533);
xnor U35126 (N_35126,N_34735,N_34134);
nand U35127 (N_35127,N_34559,N_34626);
and U35128 (N_35128,N_34476,N_34422);
or U35129 (N_35129,N_34398,N_34306);
xor U35130 (N_35130,N_34374,N_34170);
or U35131 (N_35131,N_34101,N_34768);
or U35132 (N_35132,N_34738,N_34890);
nor U35133 (N_35133,N_34592,N_34960);
or U35134 (N_35134,N_34546,N_34296);
nor U35135 (N_35135,N_34130,N_34453);
nor U35136 (N_35136,N_34421,N_34333);
xor U35137 (N_35137,N_34158,N_34188);
and U35138 (N_35138,N_34945,N_34231);
nand U35139 (N_35139,N_34993,N_34321);
and U35140 (N_35140,N_34557,N_34322);
nand U35141 (N_35141,N_34457,N_34583);
nand U35142 (N_35142,N_34874,N_34947);
nor U35143 (N_35143,N_34791,N_34909);
or U35144 (N_35144,N_34066,N_34345);
or U35145 (N_35145,N_34658,N_34169);
or U35146 (N_35146,N_34282,N_34975);
nand U35147 (N_35147,N_34870,N_34178);
nor U35148 (N_35148,N_34816,N_34675);
xnor U35149 (N_35149,N_34047,N_34695);
nor U35150 (N_35150,N_34425,N_34010);
or U35151 (N_35151,N_34734,N_34383);
nor U35152 (N_35152,N_34548,N_34722);
or U35153 (N_35153,N_34653,N_34479);
or U35154 (N_35154,N_34058,N_34657);
nand U35155 (N_35155,N_34315,N_34885);
xor U35156 (N_35156,N_34671,N_34343);
xor U35157 (N_35157,N_34480,N_34921);
nand U35158 (N_35158,N_34439,N_34091);
nand U35159 (N_35159,N_34594,N_34891);
xnor U35160 (N_35160,N_34135,N_34585);
and U35161 (N_35161,N_34514,N_34524);
nor U35162 (N_35162,N_34403,N_34054);
xor U35163 (N_35163,N_34340,N_34865);
nor U35164 (N_35164,N_34230,N_34511);
or U35165 (N_35165,N_34369,N_34413);
xor U35166 (N_35166,N_34830,N_34604);
or U35167 (N_35167,N_34525,N_34447);
xnor U35168 (N_35168,N_34085,N_34234);
nor U35169 (N_35169,N_34493,N_34172);
xnor U35170 (N_35170,N_34388,N_34717);
nand U35171 (N_35171,N_34308,N_34166);
nor U35172 (N_35172,N_34543,N_34652);
nand U35173 (N_35173,N_34219,N_34146);
and U35174 (N_35174,N_34077,N_34168);
nor U35175 (N_35175,N_34244,N_34127);
nor U35176 (N_35176,N_34268,N_34997);
xor U35177 (N_35177,N_34337,N_34263);
and U35178 (N_35178,N_34932,N_34133);
nand U35179 (N_35179,N_34507,N_34191);
xnor U35180 (N_35180,N_34705,N_34676);
and U35181 (N_35181,N_34487,N_34840);
nand U35182 (N_35182,N_34931,N_34875);
and U35183 (N_35183,N_34068,N_34470);
nor U35184 (N_35184,N_34469,N_34083);
and U35185 (N_35185,N_34038,N_34372);
or U35186 (N_35186,N_34863,N_34184);
or U35187 (N_35187,N_34683,N_34119);
nand U35188 (N_35188,N_34905,N_34835);
nand U35189 (N_35189,N_34145,N_34685);
or U35190 (N_35190,N_34659,N_34895);
nor U35191 (N_35191,N_34572,N_34574);
or U35192 (N_35192,N_34356,N_34701);
nor U35193 (N_35193,N_34269,N_34692);
and U35194 (N_35194,N_34102,N_34245);
nor U35195 (N_35195,N_34173,N_34227);
nand U35196 (N_35196,N_34946,N_34582);
and U35197 (N_35197,N_34212,N_34304);
or U35198 (N_35198,N_34995,N_34309);
nand U35199 (N_35199,N_34149,N_34046);
nor U35200 (N_35200,N_34297,N_34650);
xnor U35201 (N_35201,N_34281,N_34370);
and U35202 (N_35202,N_34478,N_34189);
xnor U35203 (N_35203,N_34745,N_34011);
and U35204 (N_35204,N_34108,N_34779);
nand U35205 (N_35205,N_34060,N_34631);
and U35206 (N_35206,N_34395,N_34092);
or U35207 (N_35207,N_34820,N_34477);
xnor U35208 (N_35208,N_34073,N_34861);
or U35209 (N_35209,N_34289,N_34573);
and U35210 (N_35210,N_34229,N_34979);
xnor U35211 (N_35211,N_34142,N_34967);
xor U35212 (N_35212,N_34549,N_34030);
nand U35213 (N_35213,N_34610,N_34884);
nor U35214 (N_35214,N_34617,N_34517);
xor U35215 (N_35215,N_34756,N_34868);
or U35216 (N_35216,N_34892,N_34872);
nor U35217 (N_35217,N_34752,N_34241);
and U35218 (N_35218,N_34409,N_34535);
nand U35219 (N_35219,N_34796,N_34265);
nand U35220 (N_35220,N_34826,N_34858);
nand U35221 (N_35221,N_34601,N_34784);
and U35222 (N_35222,N_34114,N_34744);
xor U35223 (N_35223,N_34953,N_34498);
xor U35224 (N_35224,N_34965,N_34473);
and U35225 (N_35225,N_34090,N_34031);
nand U35226 (N_35226,N_34609,N_34371);
or U35227 (N_35227,N_34213,N_34405);
nand U35228 (N_35228,N_34482,N_34264);
nor U35229 (N_35229,N_34916,N_34095);
and U35230 (N_35230,N_34221,N_34402);
nand U35231 (N_35231,N_34125,N_34275);
or U35232 (N_35232,N_34406,N_34298);
and U35233 (N_35233,N_34079,N_34974);
xor U35234 (N_35234,N_34222,N_34668);
nand U35235 (N_35235,N_34044,N_34233);
nand U35236 (N_35236,N_34504,N_34638);
and U35237 (N_35237,N_34545,N_34278);
nand U35238 (N_35238,N_34299,N_34699);
or U35239 (N_35239,N_34332,N_34903);
nor U35240 (N_35240,N_34542,N_34150);
xor U35241 (N_35241,N_34919,N_34726);
or U35242 (N_35242,N_34771,N_34742);
nand U35243 (N_35243,N_34259,N_34088);
nand U35244 (N_35244,N_34560,N_34757);
nand U35245 (N_35245,N_34065,N_34908);
or U35246 (N_35246,N_34005,N_34075);
xor U35247 (N_35247,N_34750,N_34970);
nand U35248 (N_35248,N_34941,N_34556);
and U35249 (N_35249,N_34725,N_34448);
or U35250 (N_35250,N_34240,N_34966);
nor U35251 (N_35251,N_34009,N_34508);
or U35252 (N_35252,N_34139,N_34161);
and U35253 (N_35253,N_34202,N_34899);
and U35254 (N_35254,N_34160,N_34579);
and U35255 (N_35255,N_34106,N_34074);
nor U35256 (N_35256,N_34871,N_34045);
or U35257 (N_35257,N_34380,N_34379);
and U35258 (N_35258,N_34334,N_34026);
or U35259 (N_35259,N_34355,N_34148);
xor U35260 (N_35260,N_34239,N_34254);
and U35261 (N_35261,N_34452,N_34977);
nor U35262 (N_35262,N_34414,N_34408);
and U35263 (N_35263,N_34973,N_34099);
nand U35264 (N_35264,N_34926,N_34539);
nand U35265 (N_35265,N_34123,N_34800);
nand U35266 (N_35266,N_34113,N_34569);
nand U35267 (N_35267,N_34152,N_34410);
or U35268 (N_35268,N_34841,N_34731);
nand U35269 (N_35269,N_34554,N_34994);
xnor U35270 (N_35270,N_34581,N_34248);
nor U35271 (N_35271,N_34691,N_34949);
nand U35272 (N_35272,N_34043,N_34939);
nand U35273 (N_35273,N_34352,N_34250);
or U35274 (N_35274,N_34002,N_34235);
nand U35275 (N_35275,N_34866,N_34911);
and U35276 (N_35276,N_34568,N_34623);
and U35277 (N_35277,N_34702,N_34985);
nor U35278 (N_35278,N_34620,N_34270);
and U35279 (N_35279,N_34584,N_34012);
xnor U35280 (N_35280,N_34906,N_34828);
and U35281 (N_35281,N_34983,N_34635);
nand U35282 (N_35282,N_34103,N_34489);
xor U35283 (N_35283,N_34608,N_34855);
nor U35284 (N_35284,N_34454,N_34600);
or U35285 (N_35285,N_34019,N_34645);
or U35286 (N_35286,N_34285,N_34673);
nand U35287 (N_35287,N_34314,N_34358);
or U35288 (N_35288,N_34037,N_34603);
nor U35289 (N_35289,N_34424,N_34474);
nand U35290 (N_35290,N_34770,N_34353);
xor U35291 (N_35291,N_34220,N_34697);
nor U35292 (N_35292,N_34137,N_34562);
nor U35293 (N_35293,N_34833,N_34775);
nor U35294 (N_35294,N_34208,N_34144);
nor U35295 (N_35295,N_34810,N_34522);
nor U35296 (N_35296,N_34443,N_34976);
nor U35297 (N_35297,N_34132,N_34185);
xor U35298 (N_35298,N_34217,N_34435);
or U35299 (N_35299,N_34565,N_34367);
nand U35300 (N_35300,N_34324,N_34365);
xnor U35301 (N_35301,N_34341,N_34786);
or U35302 (N_35302,N_34710,N_34769);
nor U35303 (N_35303,N_34704,N_34497);
and U35304 (N_35304,N_34401,N_34021);
nor U35305 (N_35305,N_34121,N_34035);
nor U35306 (N_35306,N_34743,N_34625);
and U35307 (N_35307,N_34393,N_34116);
xnor U35308 (N_35308,N_34151,N_34118);
nor U35309 (N_35309,N_34766,N_34175);
or U35310 (N_35310,N_34968,N_34243);
nand U35311 (N_35311,N_34377,N_34437);
or U35312 (N_35312,N_34375,N_34376);
xor U35313 (N_35313,N_34544,N_34211);
or U35314 (N_35314,N_34759,N_34915);
xnor U35315 (N_35315,N_34978,N_34481);
and U35316 (N_35316,N_34857,N_34018);
and U35317 (N_35317,N_34733,N_34805);
nand U35318 (N_35318,N_34996,N_34015);
nand U35319 (N_35319,N_34201,N_34839);
xor U35320 (N_35320,N_34611,N_34740);
nand U35321 (N_35321,N_34661,N_34466);
xnor U35322 (N_35322,N_34897,N_34706);
nor U35323 (N_35323,N_34989,N_34589);
nor U35324 (N_35324,N_34404,N_34730);
and U35325 (N_35325,N_34936,N_34984);
nor U35326 (N_35326,N_34228,N_34320);
nor U35327 (N_35327,N_34780,N_34257);
xnor U35328 (N_35328,N_34179,N_34029);
or U35329 (N_35329,N_34520,N_34593);
nand U35330 (N_35330,N_34943,N_34363);
xnor U35331 (N_35331,N_34540,N_34602);
or U35332 (N_35332,N_34359,N_34503);
nand U35333 (N_35333,N_34318,N_34008);
and U35334 (N_35334,N_34261,N_34718);
and U35335 (N_35335,N_34845,N_34500);
nor U35336 (N_35336,N_34896,N_34838);
xnor U35337 (N_35337,N_34071,N_34061);
and U35338 (N_35338,N_34920,N_34822);
xnor U35339 (N_35339,N_34694,N_34154);
nand U35340 (N_35340,N_34316,N_34817);
nor U35341 (N_35341,N_34782,N_34621);
or U35342 (N_35342,N_34630,N_34098);
nor U35343 (N_35343,N_34647,N_34527);
xor U35344 (N_35344,N_34427,N_34538);
or U35345 (N_35345,N_34327,N_34505);
nor U35346 (N_35346,N_34467,N_34338);
or U35347 (N_35347,N_34934,N_34247);
nand U35348 (N_35348,N_34223,N_34566);
nand U35349 (N_35349,N_34128,N_34806);
and U35350 (N_35350,N_34824,N_34886);
nor U35351 (N_35351,N_34164,N_34397);
or U35352 (N_35352,N_34426,N_34465);
and U35353 (N_35353,N_34273,N_34925);
and U35354 (N_35354,N_34801,N_34843);
nand U35355 (N_35355,N_34360,N_34381);
or U35356 (N_35356,N_34253,N_34591);
nand U35357 (N_35357,N_34041,N_34111);
xnor U35358 (N_35358,N_34862,N_34214);
nand U35359 (N_35359,N_34537,N_34687);
and U35360 (N_35360,N_34440,N_34399);
nand U35361 (N_35361,N_34059,N_34823);
xnor U35362 (N_35362,N_34347,N_34785);
nand U35363 (N_35363,N_34199,N_34696);
nand U35364 (N_35364,N_34962,N_34311);
and U35365 (N_35365,N_34831,N_34762);
xor U35366 (N_35366,N_34190,N_34679);
or U35367 (N_35367,N_34887,N_34003);
nand U35368 (N_35368,N_34901,N_34814);
nor U35369 (N_35369,N_34033,N_34709);
or U35370 (N_35370,N_34286,N_34389);
nor U35371 (N_35371,N_34195,N_34963);
nand U35372 (N_35372,N_34491,N_34651);
nand U35373 (N_35373,N_34515,N_34856);
or U35374 (N_35374,N_34930,N_34528);
and U35375 (N_35375,N_34153,N_34700);
nand U35376 (N_35376,N_34981,N_34081);
nand U35377 (N_35377,N_34563,N_34100);
and U35378 (N_35378,N_34419,N_34808);
or U35379 (N_35379,N_34681,N_34715);
nand U35380 (N_35380,N_34519,N_34373);
and U35381 (N_35381,N_34724,N_34713);
nor U35382 (N_35382,N_34020,N_34423);
nand U35383 (N_35383,N_34034,N_34506);
nand U35384 (N_35384,N_34940,N_34407);
and U35385 (N_35385,N_34811,N_34643);
or U35386 (N_35386,N_34952,N_34057);
nand U35387 (N_35387,N_34428,N_34147);
and U35388 (N_35388,N_34207,N_34913);
xnor U35389 (N_35389,N_34708,N_34361);
nor U35390 (N_35390,N_34716,N_34529);
nor U35391 (N_35391,N_34459,N_34864);
nand U35392 (N_35392,N_34412,N_34813);
nor U35393 (N_35393,N_34462,N_34669);
or U35394 (N_35394,N_34888,N_34555);
nand U35395 (N_35395,N_34394,N_34305);
nor U35396 (N_35396,N_34080,N_34112);
or U35397 (N_35397,N_34416,N_34067);
xor U35398 (N_35398,N_34069,N_34236);
and U35399 (N_35399,N_34001,N_34460);
or U35400 (N_35400,N_34138,N_34053);
nand U35401 (N_35401,N_34004,N_34662);
and U35402 (N_35402,N_34873,N_34215);
nor U35403 (N_35403,N_34627,N_34969);
and U35404 (N_35404,N_34819,N_34570);
nor U35405 (N_35405,N_34120,N_34070);
nand U35406 (N_35406,N_34812,N_34578);
nor U35407 (N_35407,N_34629,N_34876);
and U35408 (N_35408,N_34666,N_34483);
nor U35409 (N_35409,N_34927,N_34530);
xnor U35410 (N_35410,N_34859,N_34255);
xor U35411 (N_35411,N_34115,N_34860);
or U35412 (N_35412,N_34494,N_34721);
and U35413 (N_35413,N_34107,N_34256);
nor U35414 (N_35414,N_34576,N_34799);
or U35415 (N_35415,N_34640,N_34302);
nor U35416 (N_35416,N_34342,N_34655);
and U35417 (N_35417,N_34194,N_34547);
nand U35418 (N_35418,N_34882,N_34386);
nor U35419 (N_35419,N_34176,N_34392);
nand U35420 (N_35420,N_34129,N_34163);
or U35421 (N_35421,N_34632,N_34052);
or U35422 (N_35422,N_34992,N_34287);
or U35423 (N_35423,N_34461,N_34456);
nand U35424 (N_35424,N_34867,N_34472);
and U35425 (N_35425,N_34746,N_34048);
or U35426 (N_35426,N_34288,N_34198);
or U35427 (N_35427,N_34998,N_34193);
or U35428 (N_35428,N_34928,N_34032);
xor U35429 (N_35429,N_34105,N_34023);
nor U35430 (N_35430,N_34451,N_34348);
xor U35431 (N_35431,N_34350,N_34136);
and U35432 (N_35432,N_34512,N_34022);
or U35433 (N_35433,N_34096,N_34171);
and U35434 (N_35434,N_34804,N_34792);
nor U35435 (N_35435,N_34366,N_34006);
and U35436 (N_35436,N_34499,N_34450);
xnor U35437 (N_35437,N_34155,N_34561);
and U35438 (N_35438,N_34988,N_34586);
and U35439 (N_35439,N_34958,N_34301);
nand U35440 (N_35440,N_34186,N_34599);
nand U35441 (N_35441,N_34441,N_34013);
nor U35442 (N_35442,N_34935,N_34809);
and U35443 (N_35443,N_34317,N_34986);
nand U35444 (N_35444,N_34368,N_34310);
nand U35445 (N_35445,N_34094,N_34571);
and U35446 (N_35446,N_34737,N_34267);
or U35447 (N_35447,N_34141,N_34829);
and U35448 (N_35448,N_34078,N_34924);
xnor U35449 (N_35449,N_34907,N_34328);
and U35450 (N_35450,N_34990,N_34204);
or U35451 (N_35451,N_34849,N_34852);
and U35452 (N_35452,N_34677,N_34550);
or U35453 (N_35453,N_34917,N_34357);
and U35454 (N_35454,N_34760,N_34354);
and U35455 (N_35455,N_34894,N_34484);
xor U35456 (N_35456,N_34624,N_34719);
xor U35457 (N_35457,N_34954,N_34433);
or U35458 (N_35458,N_34272,N_34458);
nor U35459 (N_35459,N_34912,N_34294);
nor U35460 (N_35460,N_34496,N_34205);
nor U35461 (N_35461,N_34521,N_34646);
nand U35462 (N_35462,N_34017,N_34089);
or U35463 (N_35463,N_34051,N_34266);
and U35464 (N_35464,N_34764,N_34649);
nor U35465 (N_35465,N_34844,N_34177);
or U35466 (N_35466,N_34510,N_34502);
and U35467 (N_35467,N_34260,N_34087);
nand U35468 (N_35468,N_34262,N_34980);
nand U35469 (N_35469,N_34558,N_34904);
or U35470 (N_35470,N_34526,N_34682);
nor U35471 (N_35471,N_34881,N_34720);
nand U35472 (N_35472,N_34534,N_34280);
xnor U35473 (N_35473,N_34384,N_34741);
or U35474 (N_35474,N_34252,N_34216);
nor U35475 (N_35475,N_34536,N_34313);
or U35476 (N_35476,N_34767,N_34455);
and U35477 (N_35477,N_34848,N_34295);
xor U35478 (N_35478,N_34126,N_34062);
or U35479 (N_35479,N_34564,N_34206);
nand U35480 (N_35480,N_34991,N_34218);
nand U35481 (N_35481,N_34641,N_34025);
nand U35482 (N_35482,N_34674,N_34420);
nand U35483 (N_35483,N_34851,N_34982);
xnor U35484 (N_35484,N_34446,N_34818);
or U35485 (N_35485,N_34567,N_34344);
xnor U35486 (N_35486,N_34203,N_34418);
or U35487 (N_35487,N_34396,N_34728);
nor U35488 (N_35488,N_34634,N_34642);
or U35489 (N_35489,N_34237,N_34449);
and U35490 (N_35490,N_34850,N_34024);
nand U35491 (N_35491,N_34614,N_34000);
nor U35492 (N_35492,N_34703,N_34226);
nor U35493 (N_35493,N_34783,N_34391);
nor U35494 (N_35494,N_34878,N_34346);
nor U35495 (N_35495,N_34803,N_34948);
nor U35496 (N_35496,N_34607,N_34957);
and U35497 (N_35497,N_34846,N_34933);
xnor U35498 (N_35498,N_34167,N_34276);
nand U35499 (N_35499,N_34712,N_34445);
nor U35500 (N_35500,N_34053,N_34740);
nor U35501 (N_35501,N_34680,N_34946);
nand U35502 (N_35502,N_34753,N_34816);
or U35503 (N_35503,N_34710,N_34536);
or U35504 (N_35504,N_34148,N_34287);
xor U35505 (N_35505,N_34564,N_34187);
nand U35506 (N_35506,N_34274,N_34201);
and U35507 (N_35507,N_34106,N_34213);
xor U35508 (N_35508,N_34368,N_34051);
nand U35509 (N_35509,N_34341,N_34342);
nor U35510 (N_35510,N_34409,N_34589);
nor U35511 (N_35511,N_34325,N_34450);
and U35512 (N_35512,N_34212,N_34677);
and U35513 (N_35513,N_34300,N_34454);
and U35514 (N_35514,N_34502,N_34647);
nand U35515 (N_35515,N_34348,N_34006);
nand U35516 (N_35516,N_34155,N_34929);
nand U35517 (N_35517,N_34271,N_34269);
and U35518 (N_35518,N_34559,N_34793);
nor U35519 (N_35519,N_34009,N_34457);
or U35520 (N_35520,N_34179,N_34219);
xor U35521 (N_35521,N_34364,N_34077);
xor U35522 (N_35522,N_34430,N_34545);
xor U35523 (N_35523,N_34054,N_34526);
xnor U35524 (N_35524,N_34914,N_34640);
and U35525 (N_35525,N_34421,N_34949);
nand U35526 (N_35526,N_34059,N_34545);
or U35527 (N_35527,N_34553,N_34235);
or U35528 (N_35528,N_34061,N_34977);
and U35529 (N_35529,N_34772,N_34146);
and U35530 (N_35530,N_34664,N_34818);
and U35531 (N_35531,N_34903,N_34910);
and U35532 (N_35532,N_34752,N_34175);
nor U35533 (N_35533,N_34491,N_34576);
xor U35534 (N_35534,N_34736,N_34394);
nor U35535 (N_35535,N_34045,N_34275);
nand U35536 (N_35536,N_34733,N_34601);
or U35537 (N_35537,N_34579,N_34027);
nand U35538 (N_35538,N_34965,N_34282);
xnor U35539 (N_35539,N_34257,N_34974);
and U35540 (N_35540,N_34131,N_34077);
or U35541 (N_35541,N_34123,N_34214);
nor U35542 (N_35542,N_34456,N_34966);
xor U35543 (N_35543,N_34078,N_34997);
xor U35544 (N_35544,N_34062,N_34812);
and U35545 (N_35545,N_34848,N_34125);
or U35546 (N_35546,N_34398,N_34562);
xnor U35547 (N_35547,N_34071,N_34973);
or U35548 (N_35548,N_34263,N_34231);
and U35549 (N_35549,N_34749,N_34791);
nand U35550 (N_35550,N_34616,N_34032);
nand U35551 (N_35551,N_34304,N_34687);
xor U35552 (N_35552,N_34101,N_34811);
nand U35553 (N_35553,N_34460,N_34018);
and U35554 (N_35554,N_34868,N_34426);
or U35555 (N_35555,N_34168,N_34276);
nor U35556 (N_35556,N_34168,N_34791);
or U35557 (N_35557,N_34105,N_34421);
nor U35558 (N_35558,N_34318,N_34247);
nand U35559 (N_35559,N_34034,N_34889);
and U35560 (N_35560,N_34215,N_34876);
nand U35561 (N_35561,N_34654,N_34492);
nor U35562 (N_35562,N_34979,N_34606);
nand U35563 (N_35563,N_34994,N_34049);
nand U35564 (N_35564,N_34455,N_34929);
and U35565 (N_35565,N_34751,N_34215);
nor U35566 (N_35566,N_34767,N_34688);
and U35567 (N_35567,N_34292,N_34345);
or U35568 (N_35568,N_34402,N_34883);
nor U35569 (N_35569,N_34485,N_34557);
and U35570 (N_35570,N_34818,N_34673);
xnor U35571 (N_35571,N_34218,N_34984);
or U35572 (N_35572,N_34295,N_34332);
xnor U35573 (N_35573,N_34625,N_34067);
nor U35574 (N_35574,N_34137,N_34102);
nor U35575 (N_35575,N_34535,N_34691);
nand U35576 (N_35576,N_34483,N_34213);
or U35577 (N_35577,N_34716,N_34581);
or U35578 (N_35578,N_34950,N_34051);
and U35579 (N_35579,N_34607,N_34160);
xor U35580 (N_35580,N_34330,N_34601);
nor U35581 (N_35581,N_34284,N_34848);
or U35582 (N_35582,N_34706,N_34506);
and U35583 (N_35583,N_34725,N_34918);
and U35584 (N_35584,N_34086,N_34383);
nor U35585 (N_35585,N_34812,N_34828);
and U35586 (N_35586,N_34620,N_34266);
or U35587 (N_35587,N_34370,N_34662);
nor U35588 (N_35588,N_34193,N_34111);
or U35589 (N_35589,N_34946,N_34612);
xor U35590 (N_35590,N_34243,N_34639);
nand U35591 (N_35591,N_34050,N_34071);
xnor U35592 (N_35592,N_34745,N_34004);
xor U35593 (N_35593,N_34656,N_34650);
or U35594 (N_35594,N_34724,N_34118);
or U35595 (N_35595,N_34818,N_34240);
nand U35596 (N_35596,N_34370,N_34259);
nand U35597 (N_35597,N_34421,N_34028);
or U35598 (N_35598,N_34640,N_34219);
xor U35599 (N_35599,N_34565,N_34493);
nor U35600 (N_35600,N_34177,N_34464);
or U35601 (N_35601,N_34417,N_34265);
or U35602 (N_35602,N_34878,N_34661);
and U35603 (N_35603,N_34577,N_34267);
nor U35604 (N_35604,N_34240,N_34065);
and U35605 (N_35605,N_34502,N_34779);
and U35606 (N_35606,N_34276,N_34093);
or U35607 (N_35607,N_34286,N_34479);
nor U35608 (N_35608,N_34668,N_34211);
xor U35609 (N_35609,N_34130,N_34278);
and U35610 (N_35610,N_34808,N_34907);
xnor U35611 (N_35611,N_34065,N_34789);
xnor U35612 (N_35612,N_34089,N_34366);
nor U35613 (N_35613,N_34236,N_34243);
or U35614 (N_35614,N_34478,N_34654);
xor U35615 (N_35615,N_34186,N_34645);
xor U35616 (N_35616,N_34755,N_34857);
xnor U35617 (N_35617,N_34835,N_34414);
or U35618 (N_35618,N_34295,N_34585);
xnor U35619 (N_35619,N_34442,N_34070);
nand U35620 (N_35620,N_34212,N_34216);
and U35621 (N_35621,N_34991,N_34940);
nor U35622 (N_35622,N_34685,N_34548);
nand U35623 (N_35623,N_34493,N_34532);
and U35624 (N_35624,N_34528,N_34345);
xnor U35625 (N_35625,N_34892,N_34906);
and U35626 (N_35626,N_34948,N_34228);
xnor U35627 (N_35627,N_34432,N_34881);
nand U35628 (N_35628,N_34496,N_34407);
or U35629 (N_35629,N_34013,N_34776);
or U35630 (N_35630,N_34005,N_34163);
or U35631 (N_35631,N_34236,N_34404);
or U35632 (N_35632,N_34030,N_34843);
nor U35633 (N_35633,N_34764,N_34775);
nor U35634 (N_35634,N_34804,N_34989);
nand U35635 (N_35635,N_34284,N_34016);
nand U35636 (N_35636,N_34847,N_34528);
nor U35637 (N_35637,N_34842,N_34071);
and U35638 (N_35638,N_34205,N_34945);
or U35639 (N_35639,N_34296,N_34708);
nand U35640 (N_35640,N_34084,N_34920);
xor U35641 (N_35641,N_34211,N_34343);
and U35642 (N_35642,N_34634,N_34614);
or U35643 (N_35643,N_34958,N_34744);
nor U35644 (N_35644,N_34188,N_34413);
and U35645 (N_35645,N_34179,N_34708);
nor U35646 (N_35646,N_34694,N_34027);
or U35647 (N_35647,N_34127,N_34084);
xnor U35648 (N_35648,N_34922,N_34489);
or U35649 (N_35649,N_34421,N_34256);
nand U35650 (N_35650,N_34062,N_34875);
xnor U35651 (N_35651,N_34948,N_34860);
xnor U35652 (N_35652,N_34502,N_34914);
and U35653 (N_35653,N_34133,N_34870);
or U35654 (N_35654,N_34109,N_34350);
nand U35655 (N_35655,N_34417,N_34235);
and U35656 (N_35656,N_34761,N_34608);
or U35657 (N_35657,N_34462,N_34597);
nor U35658 (N_35658,N_34293,N_34257);
nor U35659 (N_35659,N_34275,N_34026);
xnor U35660 (N_35660,N_34930,N_34995);
nand U35661 (N_35661,N_34374,N_34284);
or U35662 (N_35662,N_34176,N_34437);
nor U35663 (N_35663,N_34660,N_34212);
nor U35664 (N_35664,N_34544,N_34479);
and U35665 (N_35665,N_34671,N_34401);
and U35666 (N_35666,N_34625,N_34379);
xor U35667 (N_35667,N_34689,N_34274);
or U35668 (N_35668,N_34650,N_34040);
nand U35669 (N_35669,N_34528,N_34364);
xnor U35670 (N_35670,N_34783,N_34489);
and U35671 (N_35671,N_34088,N_34890);
nand U35672 (N_35672,N_34008,N_34158);
or U35673 (N_35673,N_34869,N_34412);
xor U35674 (N_35674,N_34554,N_34929);
xor U35675 (N_35675,N_34611,N_34664);
nor U35676 (N_35676,N_34102,N_34684);
or U35677 (N_35677,N_34958,N_34258);
xnor U35678 (N_35678,N_34100,N_34250);
xnor U35679 (N_35679,N_34587,N_34544);
nand U35680 (N_35680,N_34920,N_34950);
and U35681 (N_35681,N_34850,N_34588);
nor U35682 (N_35682,N_34742,N_34504);
or U35683 (N_35683,N_34355,N_34904);
nand U35684 (N_35684,N_34117,N_34200);
and U35685 (N_35685,N_34938,N_34313);
xnor U35686 (N_35686,N_34024,N_34493);
xnor U35687 (N_35687,N_34310,N_34132);
or U35688 (N_35688,N_34853,N_34501);
xor U35689 (N_35689,N_34492,N_34044);
and U35690 (N_35690,N_34129,N_34890);
xor U35691 (N_35691,N_34359,N_34160);
and U35692 (N_35692,N_34027,N_34056);
and U35693 (N_35693,N_34308,N_34385);
and U35694 (N_35694,N_34454,N_34414);
nand U35695 (N_35695,N_34485,N_34872);
nand U35696 (N_35696,N_34491,N_34867);
xnor U35697 (N_35697,N_34063,N_34960);
nor U35698 (N_35698,N_34905,N_34770);
nor U35699 (N_35699,N_34236,N_34870);
or U35700 (N_35700,N_34872,N_34338);
nand U35701 (N_35701,N_34201,N_34882);
nand U35702 (N_35702,N_34812,N_34140);
nand U35703 (N_35703,N_34499,N_34524);
nand U35704 (N_35704,N_34341,N_34228);
xor U35705 (N_35705,N_34682,N_34949);
xnor U35706 (N_35706,N_34791,N_34614);
nand U35707 (N_35707,N_34508,N_34162);
and U35708 (N_35708,N_34367,N_34478);
nor U35709 (N_35709,N_34674,N_34917);
or U35710 (N_35710,N_34654,N_34502);
and U35711 (N_35711,N_34730,N_34793);
xnor U35712 (N_35712,N_34375,N_34636);
nand U35713 (N_35713,N_34298,N_34138);
and U35714 (N_35714,N_34912,N_34755);
nor U35715 (N_35715,N_34790,N_34111);
or U35716 (N_35716,N_34522,N_34641);
and U35717 (N_35717,N_34699,N_34763);
or U35718 (N_35718,N_34916,N_34251);
nand U35719 (N_35719,N_34390,N_34956);
xnor U35720 (N_35720,N_34837,N_34699);
nand U35721 (N_35721,N_34822,N_34465);
xnor U35722 (N_35722,N_34752,N_34231);
xnor U35723 (N_35723,N_34509,N_34149);
and U35724 (N_35724,N_34733,N_34498);
and U35725 (N_35725,N_34541,N_34323);
nor U35726 (N_35726,N_34502,N_34361);
and U35727 (N_35727,N_34426,N_34271);
and U35728 (N_35728,N_34227,N_34074);
nor U35729 (N_35729,N_34124,N_34783);
or U35730 (N_35730,N_34849,N_34442);
xnor U35731 (N_35731,N_34857,N_34142);
xor U35732 (N_35732,N_34720,N_34595);
and U35733 (N_35733,N_34291,N_34221);
xor U35734 (N_35734,N_34439,N_34879);
nor U35735 (N_35735,N_34544,N_34866);
nand U35736 (N_35736,N_34489,N_34011);
nor U35737 (N_35737,N_34067,N_34905);
xnor U35738 (N_35738,N_34749,N_34866);
nor U35739 (N_35739,N_34333,N_34638);
nand U35740 (N_35740,N_34963,N_34590);
xnor U35741 (N_35741,N_34739,N_34875);
and U35742 (N_35742,N_34783,N_34097);
xnor U35743 (N_35743,N_34111,N_34448);
nand U35744 (N_35744,N_34312,N_34457);
nor U35745 (N_35745,N_34608,N_34639);
nand U35746 (N_35746,N_34510,N_34046);
and U35747 (N_35747,N_34925,N_34185);
nor U35748 (N_35748,N_34187,N_34595);
or U35749 (N_35749,N_34744,N_34464);
nand U35750 (N_35750,N_34568,N_34413);
xnor U35751 (N_35751,N_34026,N_34349);
or U35752 (N_35752,N_34709,N_34167);
xnor U35753 (N_35753,N_34488,N_34522);
or U35754 (N_35754,N_34176,N_34017);
xor U35755 (N_35755,N_34996,N_34966);
and U35756 (N_35756,N_34206,N_34175);
xor U35757 (N_35757,N_34848,N_34310);
nor U35758 (N_35758,N_34307,N_34750);
nor U35759 (N_35759,N_34809,N_34430);
nor U35760 (N_35760,N_34086,N_34376);
nor U35761 (N_35761,N_34343,N_34687);
nor U35762 (N_35762,N_34693,N_34813);
xor U35763 (N_35763,N_34218,N_34655);
nand U35764 (N_35764,N_34258,N_34689);
xor U35765 (N_35765,N_34409,N_34027);
xnor U35766 (N_35766,N_34462,N_34479);
or U35767 (N_35767,N_34768,N_34032);
nor U35768 (N_35768,N_34092,N_34554);
nand U35769 (N_35769,N_34567,N_34410);
and U35770 (N_35770,N_34662,N_34993);
nand U35771 (N_35771,N_34681,N_34677);
xnor U35772 (N_35772,N_34746,N_34141);
nor U35773 (N_35773,N_34866,N_34795);
or U35774 (N_35774,N_34659,N_34480);
or U35775 (N_35775,N_34843,N_34537);
xor U35776 (N_35776,N_34783,N_34537);
nor U35777 (N_35777,N_34985,N_34830);
nand U35778 (N_35778,N_34597,N_34268);
nand U35779 (N_35779,N_34594,N_34222);
or U35780 (N_35780,N_34948,N_34452);
and U35781 (N_35781,N_34161,N_34457);
nand U35782 (N_35782,N_34499,N_34463);
xnor U35783 (N_35783,N_34671,N_34054);
or U35784 (N_35784,N_34682,N_34535);
nor U35785 (N_35785,N_34450,N_34455);
or U35786 (N_35786,N_34932,N_34240);
nor U35787 (N_35787,N_34681,N_34895);
xnor U35788 (N_35788,N_34287,N_34178);
nand U35789 (N_35789,N_34150,N_34915);
nor U35790 (N_35790,N_34237,N_34217);
nand U35791 (N_35791,N_34581,N_34353);
nand U35792 (N_35792,N_34866,N_34593);
and U35793 (N_35793,N_34718,N_34369);
xnor U35794 (N_35794,N_34326,N_34359);
or U35795 (N_35795,N_34669,N_34239);
nand U35796 (N_35796,N_34606,N_34423);
nor U35797 (N_35797,N_34524,N_34799);
or U35798 (N_35798,N_34537,N_34463);
or U35799 (N_35799,N_34073,N_34552);
xor U35800 (N_35800,N_34072,N_34738);
or U35801 (N_35801,N_34302,N_34312);
and U35802 (N_35802,N_34505,N_34043);
nand U35803 (N_35803,N_34297,N_34867);
nand U35804 (N_35804,N_34476,N_34119);
or U35805 (N_35805,N_34653,N_34733);
and U35806 (N_35806,N_34560,N_34086);
nor U35807 (N_35807,N_34438,N_34013);
and U35808 (N_35808,N_34045,N_34610);
and U35809 (N_35809,N_34321,N_34529);
nor U35810 (N_35810,N_34283,N_34113);
nand U35811 (N_35811,N_34894,N_34744);
nand U35812 (N_35812,N_34725,N_34473);
nor U35813 (N_35813,N_34639,N_34754);
xor U35814 (N_35814,N_34268,N_34595);
and U35815 (N_35815,N_34706,N_34989);
nand U35816 (N_35816,N_34580,N_34633);
or U35817 (N_35817,N_34720,N_34631);
or U35818 (N_35818,N_34197,N_34762);
or U35819 (N_35819,N_34878,N_34145);
or U35820 (N_35820,N_34125,N_34091);
nand U35821 (N_35821,N_34902,N_34422);
nor U35822 (N_35822,N_34421,N_34950);
or U35823 (N_35823,N_34160,N_34393);
and U35824 (N_35824,N_34584,N_34159);
or U35825 (N_35825,N_34987,N_34537);
nor U35826 (N_35826,N_34045,N_34824);
nor U35827 (N_35827,N_34223,N_34392);
nor U35828 (N_35828,N_34979,N_34360);
or U35829 (N_35829,N_34670,N_34167);
xnor U35830 (N_35830,N_34594,N_34073);
and U35831 (N_35831,N_34409,N_34691);
nor U35832 (N_35832,N_34082,N_34989);
nor U35833 (N_35833,N_34326,N_34133);
nand U35834 (N_35834,N_34619,N_34301);
and U35835 (N_35835,N_34342,N_34258);
nor U35836 (N_35836,N_34386,N_34743);
nor U35837 (N_35837,N_34455,N_34504);
nand U35838 (N_35838,N_34163,N_34167);
and U35839 (N_35839,N_34083,N_34421);
or U35840 (N_35840,N_34103,N_34345);
xor U35841 (N_35841,N_34911,N_34817);
and U35842 (N_35842,N_34644,N_34960);
nand U35843 (N_35843,N_34596,N_34654);
and U35844 (N_35844,N_34540,N_34046);
or U35845 (N_35845,N_34461,N_34996);
nor U35846 (N_35846,N_34734,N_34225);
nand U35847 (N_35847,N_34121,N_34917);
nand U35848 (N_35848,N_34636,N_34338);
xor U35849 (N_35849,N_34221,N_34985);
xor U35850 (N_35850,N_34166,N_34668);
nand U35851 (N_35851,N_34168,N_34553);
or U35852 (N_35852,N_34942,N_34630);
nand U35853 (N_35853,N_34919,N_34909);
nor U35854 (N_35854,N_34234,N_34004);
and U35855 (N_35855,N_34167,N_34527);
nor U35856 (N_35856,N_34573,N_34304);
or U35857 (N_35857,N_34355,N_34172);
and U35858 (N_35858,N_34310,N_34298);
nor U35859 (N_35859,N_34799,N_34866);
xnor U35860 (N_35860,N_34610,N_34348);
xor U35861 (N_35861,N_34639,N_34808);
nand U35862 (N_35862,N_34710,N_34718);
nand U35863 (N_35863,N_34729,N_34602);
or U35864 (N_35864,N_34180,N_34774);
nand U35865 (N_35865,N_34055,N_34556);
and U35866 (N_35866,N_34793,N_34862);
nor U35867 (N_35867,N_34557,N_34148);
nor U35868 (N_35868,N_34290,N_34075);
nor U35869 (N_35869,N_34724,N_34458);
or U35870 (N_35870,N_34279,N_34926);
xor U35871 (N_35871,N_34976,N_34438);
or U35872 (N_35872,N_34815,N_34386);
and U35873 (N_35873,N_34917,N_34096);
xnor U35874 (N_35874,N_34336,N_34008);
xor U35875 (N_35875,N_34845,N_34131);
nand U35876 (N_35876,N_34841,N_34026);
nor U35877 (N_35877,N_34710,N_34041);
nor U35878 (N_35878,N_34584,N_34085);
and U35879 (N_35879,N_34864,N_34691);
nand U35880 (N_35880,N_34943,N_34556);
and U35881 (N_35881,N_34439,N_34415);
nand U35882 (N_35882,N_34722,N_34242);
nor U35883 (N_35883,N_34579,N_34134);
and U35884 (N_35884,N_34489,N_34829);
nand U35885 (N_35885,N_34296,N_34721);
xnor U35886 (N_35886,N_34614,N_34152);
or U35887 (N_35887,N_34779,N_34261);
and U35888 (N_35888,N_34036,N_34466);
xnor U35889 (N_35889,N_34312,N_34888);
xor U35890 (N_35890,N_34058,N_34950);
and U35891 (N_35891,N_34390,N_34573);
nand U35892 (N_35892,N_34579,N_34795);
nor U35893 (N_35893,N_34763,N_34046);
and U35894 (N_35894,N_34113,N_34971);
nor U35895 (N_35895,N_34767,N_34552);
or U35896 (N_35896,N_34390,N_34397);
xor U35897 (N_35897,N_34436,N_34467);
xor U35898 (N_35898,N_34344,N_34455);
or U35899 (N_35899,N_34556,N_34073);
and U35900 (N_35900,N_34783,N_34329);
and U35901 (N_35901,N_34921,N_34596);
xnor U35902 (N_35902,N_34681,N_34741);
xor U35903 (N_35903,N_34492,N_34168);
and U35904 (N_35904,N_34314,N_34914);
or U35905 (N_35905,N_34444,N_34988);
xnor U35906 (N_35906,N_34974,N_34990);
nor U35907 (N_35907,N_34620,N_34600);
xor U35908 (N_35908,N_34186,N_34880);
xnor U35909 (N_35909,N_34172,N_34241);
nand U35910 (N_35910,N_34259,N_34408);
xor U35911 (N_35911,N_34936,N_34159);
nor U35912 (N_35912,N_34107,N_34517);
and U35913 (N_35913,N_34809,N_34528);
nor U35914 (N_35914,N_34308,N_34853);
nor U35915 (N_35915,N_34903,N_34069);
or U35916 (N_35916,N_34734,N_34415);
xnor U35917 (N_35917,N_34420,N_34245);
or U35918 (N_35918,N_34185,N_34959);
and U35919 (N_35919,N_34480,N_34375);
nand U35920 (N_35920,N_34478,N_34703);
nand U35921 (N_35921,N_34457,N_34754);
or U35922 (N_35922,N_34545,N_34596);
nor U35923 (N_35923,N_34584,N_34265);
nand U35924 (N_35924,N_34383,N_34958);
or U35925 (N_35925,N_34444,N_34945);
nand U35926 (N_35926,N_34088,N_34584);
or U35927 (N_35927,N_34307,N_34264);
xnor U35928 (N_35928,N_34425,N_34660);
nor U35929 (N_35929,N_34322,N_34718);
nor U35930 (N_35930,N_34951,N_34707);
or U35931 (N_35931,N_34708,N_34141);
nor U35932 (N_35932,N_34448,N_34692);
xnor U35933 (N_35933,N_34582,N_34157);
and U35934 (N_35934,N_34273,N_34858);
and U35935 (N_35935,N_34777,N_34957);
nor U35936 (N_35936,N_34862,N_34305);
and U35937 (N_35937,N_34626,N_34024);
nand U35938 (N_35938,N_34206,N_34151);
nand U35939 (N_35939,N_34507,N_34619);
xor U35940 (N_35940,N_34522,N_34588);
and U35941 (N_35941,N_34466,N_34568);
or U35942 (N_35942,N_34778,N_34811);
xor U35943 (N_35943,N_34483,N_34627);
or U35944 (N_35944,N_34215,N_34450);
or U35945 (N_35945,N_34494,N_34326);
nand U35946 (N_35946,N_34626,N_34720);
nor U35947 (N_35947,N_34576,N_34144);
nor U35948 (N_35948,N_34795,N_34042);
nor U35949 (N_35949,N_34393,N_34093);
and U35950 (N_35950,N_34999,N_34360);
xnor U35951 (N_35951,N_34961,N_34847);
and U35952 (N_35952,N_34911,N_34469);
xnor U35953 (N_35953,N_34659,N_34992);
or U35954 (N_35954,N_34182,N_34156);
xnor U35955 (N_35955,N_34560,N_34865);
nand U35956 (N_35956,N_34812,N_34248);
nand U35957 (N_35957,N_34746,N_34008);
and U35958 (N_35958,N_34762,N_34244);
nand U35959 (N_35959,N_34766,N_34055);
nor U35960 (N_35960,N_34101,N_34702);
nand U35961 (N_35961,N_34030,N_34588);
nand U35962 (N_35962,N_34284,N_34380);
xnor U35963 (N_35963,N_34713,N_34885);
or U35964 (N_35964,N_34491,N_34280);
nand U35965 (N_35965,N_34391,N_34936);
nand U35966 (N_35966,N_34772,N_34855);
xnor U35967 (N_35967,N_34724,N_34013);
nor U35968 (N_35968,N_34826,N_34145);
nor U35969 (N_35969,N_34739,N_34302);
and U35970 (N_35970,N_34674,N_34327);
xnor U35971 (N_35971,N_34114,N_34047);
and U35972 (N_35972,N_34165,N_34133);
or U35973 (N_35973,N_34719,N_34229);
xor U35974 (N_35974,N_34332,N_34086);
nor U35975 (N_35975,N_34667,N_34502);
nand U35976 (N_35976,N_34061,N_34201);
and U35977 (N_35977,N_34783,N_34399);
nand U35978 (N_35978,N_34087,N_34494);
and U35979 (N_35979,N_34505,N_34873);
nand U35980 (N_35980,N_34344,N_34151);
nand U35981 (N_35981,N_34033,N_34458);
and U35982 (N_35982,N_34560,N_34280);
nor U35983 (N_35983,N_34100,N_34748);
or U35984 (N_35984,N_34701,N_34789);
and U35985 (N_35985,N_34460,N_34668);
xor U35986 (N_35986,N_34905,N_34886);
or U35987 (N_35987,N_34093,N_34324);
or U35988 (N_35988,N_34366,N_34413);
or U35989 (N_35989,N_34776,N_34334);
or U35990 (N_35990,N_34987,N_34146);
xnor U35991 (N_35991,N_34343,N_34069);
nor U35992 (N_35992,N_34023,N_34463);
nor U35993 (N_35993,N_34162,N_34762);
or U35994 (N_35994,N_34447,N_34901);
nand U35995 (N_35995,N_34861,N_34789);
nand U35996 (N_35996,N_34801,N_34295);
nand U35997 (N_35997,N_34556,N_34258);
nor U35998 (N_35998,N_34437,N_34458);
or U35999 (N_35999,N_34345,N_34948);
and U36000 (N_36000,N_35674,N_35978);
nor U36001 (N_36001,N_35092,N_35561);
or U36002 (N_36002,N_35793,N_35559);
nand U36003 (N_36003,N_35741,N_35280);
nor U36004 (N_36004,N_35831,N_35524);
xor U36005 (N_36005,N_35214,N_35351);
xnor U36006 (N_36006,N_35700,N_35985);
nand U36007 (N_36007,N_35344,N_35303);
and U36008 (N_36008,N_35274,N_35260);
nor U36009 (N_36009,N_35382,N_35939);
xor U36010 (N_36010,N_35299,N_35654);
xnor U36011 (N_36011,N_35589,N_35965);
or U36012 (N_36012,N_35149,N_35249);
nand U36013 (N_36013,N_35539,N_35708);
or U36014 (N_36014,N_35431,N_35864);
nand U36015 (N_36015,N_35750,N_35563);
nor U36016 (N_36016,N_35161,N_35399);
and U36017 (N_36017,N_35309,N_35088);
nand U36018 (N_36018,N_35284,N_35197);
nor U36019 (N_36019,N_35325,N_35501);
or U36020 (N_36020,N_35361,N_35115);
nor U36021 (N_36021,N_35835,N_35843);
and U36022 (N_36022,N_35160,N_35279);
or U36023 (N_36023,N_35701,N_35335);
and U36024 (N_36024,N_35729,N_35637);
nand U36025 (N_36025,N_35518,N_35560);
or U36026 (N_36026,N_35986,N_35075);
xnor U36027 (N_36027,N_35136,N_35592);
or U36028 (N_36028,N_35267,N_35053);
or U36029 (N_36029,N_35934,N_35362);
and U36030 (N_36030,N_35709,N_35899);
xnor U36031 (N_36031,N_35508,N_35929);
or U36032 (N_36032,N_35544,N_35801);
or U36033 (N_36033,N_35275,N_35246);
xnor U36034 (N_36034,N_35871,N_35973);
and U36035 (N_36035,N_35412,N_35721);
xnor U36036 (N_36036,N_35911,N_35270);
and U36037 (N_36037,N_35591,N_35924);
and U36038 (N_36038,N_35919,N_35133);
nand U36039 (N_36039,N_35210,N_35635);
xnor U36040 (N_36040,N_35828,N_35014);
and U36041 (N_36041,N_35522,N_35660);
and U36042 (N_36042,N_35254,N_35857);
nor U36043 (N_36043,N_35407,N_35672);
or U36044 (N_36044,N_35538,N_35966);
nor U36045 (N_36045,N_35314,N_35029);
nor U36046 (N_36046,N_35536,N_35153);
or U36047 (N_36047,N_35620,N_35177);
xor U36048 (N_36048,N_35002,N_35706);
and U36049 (N_36049,N_35077,N_35818);
or U36050 (N_36050,N_35349,N_35675);
nor U36051 (N_36051,N_35669,N_35456);
nor U36052 (N_36052,N_35446,N_35403);
or U36053 (N_36053,N_35528,N_35912);
xnor U36054 (N_36054,N_35594,N_35521);
nand U36055 (N_36055,N_35994,N_35435);
nor U36056 (N_36056,N_35356,N_35063);
nor U36057 (N_36057,N_35469,N_35111);
or U36058 (N_36058,N_35240,N_35781);
nor U36059 (N_36059,N_35744,N_35507);
xnor U36060 (N_36060,N_35121,N_35439);
nor U36061 (N_36061,N_35350,N_35113);
and U36062 (N_36062,N_35287,N_35099);
xor U36063 (N_36063,N_35814,N_35168);
nand U36064 (N_36064,N_35505,N_35941);
and U36065 (N_36065,N_35148,N_35320);
or U36066 (N_36066,N_35200,N_35804);
nand U36067 (N_36067,N_35948,N_35735);
or U36068 (N_36068,N_35970,N_35787);
nor U36069 (N_36069,N_35156,N_35618);
and U36070 (N_36070,N_35346,N_35603);
and U36071 (N_36071,N_35112,N_35100);
nor U36072 (N_36072,N_35341,N_35656);
or U36073 (N_36073,N_35328,N_35250);
xor U36074 (N_36074,N_35738,N_35042);
nand U36075 (N_36075,N_35208,N_35850);
xnor U36076 (N_36076,N_35535,N_35488);
nand U36077 (N_36077,N_35760,N_35598);
or U36078 (N_36078,N_35622,N_35379);
xor U36079 (N_36079,N_35454,N_35822);
and U36080 (N_36080,N_35480,N_35895);
xor U36081 (N_36081,N_35523,N_35339);
nand U36082 (N_36082,N_35228,N_35234);
xnor U36083 (N_36083,N_35266,N_35043);
xnor U36084 (N_36084,N_35155,N_35131);
nor U36085 (N_36085,N_35259,N_35185);
or U36086 (N_36086,N_35789,N_35906);
nor U36087 (N_36087,N_35323,N_35613);
xnor U36088 (N_36088,N_35510,N_35791);
or U36089 (N_36089,N_35282,N_35186);
nand U36090 (N_36090,N_35837,N_35064);
nand U36091 (N_36091,N_35332,N_35542);
nor U36092 (N_36092,N_35394,N_35663);
nor U36093 (N_36093,N_35355,N_35227);
xnor U36094 (N_36094,N_35225,N_35632);
and U36095 (N_36095,N_35852,N_35474);
nor U36096 (N_36096,N_35462,N_35874);
and U36097 (N_36097,N_35684,N_35055);
nor U36098 (N_36098,N_35441,N_35008);
nor U36099 (N_36099,N_35506,N_35812);
nand U36100 (N_36100,N_35103,N_35450);
xnor U36101 (N_36101,N_35152,N_35704);
and U36102 (N_36102,N_35979,N_35913);
nand U36103 (N_36103,N_35364,N_35726);
xor U36104 (N_36104,N_35774,N_35809);
and U36105 (N_36105,N_35612,N_35993);
nor U36106 (N_36106,N_35342,N_35269);
nor U36107 (N_36107,N_35337,N_35223);
nor U36108 (N_36108,N_35253,N_35447);
nand U36109 (N_36109,N_35090,N_35476);
nor U36110 (N_36110,N_35557,N_35652);
or U36111 (N_36111,N_35116,N_35036);
or U36112 (N_36112,N_35537,N_35723);
and U36113 (N_36113,N_35098,N_35517);
nor U36114 (N_36114,N_35384,N_35806);
xor U36115 (N_36115,N_35238,N_35262);
and U36116 (N_36116,N_35666,N_35854);
or U36117 (N_36117,N_35917,N_35128);
and U36118 (N_36118,N_35138,N_35766);
or U36119 (N_36119,N_35207,N_35398);
xnor U36120 (N_36120,N_35532,N_35513);
nand U36121 (N_36121,N_35509,N_35132);
nand U36122 (N_36122,N_35243,N_35264);
or U36123 (N_36123,N_35213,N_35671);
nor U36124 (N_36124,N_35910,N_35759);
xor U36125 (N_36125,N_35037,N_35556);
xor U36126 (N_36126,N_35658,N_35989);
nor U36127 (N_36127,N_35107,N_35526);
and U36128 (N_36128,N_35377,N_35338);
nor U36129 (N_36129,N_35391,N_35554);
nor U36130 (N_36130,N_35720,N_35171);
xnor U36131 (N_36131,N_35129,N_35315);
nor U36132 (N_36132,N_35836,N_35527);
and U36133 (N_36133,N_35548,N_35963);
or U36134 (N_36134,N_35834,N_35703);
nor U36135 (N_36135,N_35661,N_35493);
nor U36136 (N_36136,N_35956,N_35184);
nand U36137 (N_36137,N_35739,N_35761);
and U36138 (N_36138,N_35491,N_35048);
nand U36139 (N_36139,N_35035,N_35124);
or U36140 (N_36140,N_35397,N_35794);
nand U36141 (N_36141,N_35023,N_35367);
nor U36142 (N_36142,N_35875,N_35888);
nor U36143 (N_36143,N_35558,N_35841);
nor U36144 (N_36144,N_35304,N_35743);
nand U36145 (N_36145,N_35330,N_35736);
nand U36146 (N_36146,N_35707,N_35363);
nand U36147 (N_36147,N_35714,N_35856);
nor U36148 (N_36148,N_35236,N_35926);
nand U36149 (N_36149,N_35215,N_35577);
and U36150 (N_36150,N_35365,N_35353);
nand U36151 (N_36151,N_35749,N_35768);
nand U36152 (N_36152,N_35907,N_35872);
nand U36153 (N_36153,N_35685,N_35500);
nor U36154 (N_36154,N_35277,N_35316);
nand U36155 (N_36155,N_35764,N_35553);
or U36156 (N_36156,N_35595,N_35347);
nand U36157 (N_36157,N_35529,N_35614);
xnor U36158 (N_36158,N_35392,N_35845);
or U36159 (N_36159,N_35555,N_35619);
xor U36160 (N_36160,N_35593,N_35503);
xnor U36161 (N_36161,N_35626,N_35960);
or U36162 (N_36162,N_35470,N_35376);
nand U36163 (N_36163,N_35085,N_35943);
xor U36164 (N_36164,N_35826,N_35004);
and U36165 (N_36165,N_35808,N_35418);
and U36166 (N_36166,N_35786,N_35640);
nand U36167 (N_36167,N_35081,N_35853);
nand U36168 (N_36168,N_35725,N_35942);
nand U36169 (N_36169,N_35256,N_35796);
and U36170 (N_36170,N_35080,N_35642);
nor U36171 (N_36171,N_35031,N_35032);
nor U36172 (N_36172,N_35784,N_35172);
nand U36173 (N_36173,N_35052,N_35731);
and U36174 (N_36174,N_35740,N_35457);
and U36175 (N_36175,N_35992,N_35013);
nor U36176 (N_36176,N_35352,N_35058);
or U36177 (N_36177,N_35778,N_35649);
xor U36178 (N_36178,N_35991,N_35512);
and U36179 (N_36179,N_35423,N_35000);
and U36180 (N_36180,N_35990,N_35083);
and U36181 (N_36181,N_35844,N_35463);
nand U36182 (N_36182,N_35079,N_35516);
nor U36183 (N_36183,N_35466,N_35478);
or U36184 (N_36184,N_35533,N_35590);
nand U36185 (N_36185,N_35584,N_35623);
and U36186 (N_36186,N_35908,N_35422);
nor U36187 (N_36187,N_35045,N_35027);
xnor U36188 (N_36188,N_35378,N_35777);
nor U36189 (N_36189,N_35746,N_35434);
xnor U36190 (N_36190,N_35567,N_35763);
nand U36191 (N_36191,N_35101,N_35310);
and U36192 (N_36192,N_35157,N_35540);
nor U36193 (N_36193,N_35798,N_35292);
and U36194 (N_36194,N_35278,N_35813);
nand U36195 (N_36195,N_35041,N_35572);
nor U36196 (N_36196,N_35628,N_35940);
xnor U36197 (N_36197,N_35388,N_35962);
xor U36198 (N_36198,N_35018,N_35847);
and U36199 (N_36199,N_35455,N_35110);
xnor U36200 (N_36200,N_35530,N_35242);
xor U36201 (N_36201,N_35792,N_35492);
xor U36202 (N_36202,N_35247,N_35040);
and U36203 (N_36203,N_35829,N_35717);
nor U36204 (N_36204,N_35015,N_35147);
and U36205 (N_36205,N_35587,N_35406);
xnor U36206 (N_36206,N_35733,N_35302);
nand U36207 (N_36207,N_35961,N_35034);
and U36208 (N_36208,N_35862,N_35430);
or U36209 (N_36209,N_35050,N_35024);
nand U36210 (N_36210,N_35150,N_35449);
nand U36211 (N_36211,N_35046,N_35641);
nor U36212 (N_36212,N_35458,N_35281);
or U36213 (N_36213,N_35017,N_35481);
nor U36214 (N_36214,N_35196,N_35424);
nor U36215 (N_36215,N_35217,N_35866);
xnor U36216 (N_36216,N_35596,N_35779);
nand U36217 (N_36217,N_35071,N_35633);
and U36218 (N_36218,N_35915,N_35769);
nand U36219 (N_36219,N_35239,N_35459);
nand U36220 (N_36220,N_35636,N_35404);
nor U36221 (N_36221,N_35819,N_35415);
xor U36222 (N_36222,N_35576,N_35627);
xnor U36223 (N_36223,N_35105,N_35194);
nand U36224 (N_36224,N_35882,N_35117);
nand U36225 (N_36225,N_35473,N_35125);
and U36226 (N_36226,N_35935,N_35802);
nand U36227 (N_36227,N_35127,N_35520);
nand U36228 (N_36228,N_35231,N_35625);
and U36229 (N_36229,N_35451,N_35889);
nor U36230 (N_36230,N_35693,N_35319);
xnor U36231 (N_36231,N_35711,N_35732);
nor U36232 (N_36232,N_35839,N_35562);
or U36233 (N_36233,N_35673,N_35601);
nor U36234 (N_36234,N_35198,N_35780);
nand U36235 (N_36235,N_35123,N_35629);
or U36236 (N_36236,N_35305,N_35583);
xor U36237 (N_36237,N_35057,N_35930);
nand U36238 (N_36238,N_35475,N_35334);
nor U36239 (N_36239,N_35848,N_35464);
xnor U36240 (N_36240,N_35348,N_35914);
nor U36241 (N_36241,N_35519,N_35324);
nor U36242 (N_36242,N_35321,N_35062);
nor U36243 (N_36243,N_35887,N_35409);
nor U36244 (N_36244,N_35797,N_35585);
nand U36245 (N_36245,N_35599,N_35010);
or U36246 (N_36246,N_35897,N_35235);
or U36247 (N_36247,N_35145,N_35465);
nor U36248 (N_36248,N_35263,N_35662);
xor U36249 (N_36249,N_35868,N_35216);
or U36250 (N_36250,N_35187,N_35343);
xor U36251 (N_36251,N_35011,N_35790);
xnor U36252 (N_36252,N_35631,N_35087);
nand U36253 (N_36253,N_35479,N_35682);
nand U36254 (N_36254,N_35968,N_35477);
nor U36255 (N_36255,N_35710,N_35573);
nand U36256 (N_36256,N_35322,N_35816);
or U36257 (N_36257,N_35932,N_35949);
and U36258 (N_36258,N_35047,N_35855);
or U36259 (N_36259,N_35676,N_35163);
and U36260 (N_36260,N_35821,N_35368);
nor U36261 (N_36261,N_35974,N_35006);
xor U36262 (N_36262,N_35443,N_35691);
nand U36263 (N_36263,N_35289,N_35565);
or U36264 (N_36264,N_35490,N_35118);
xnor U36265 (N_36265,N_35432,N_35953);
or U36266 (N_36266,N_35211,N_35879);
or U36267 (N_36267,N_35624,N_35074);
nand U36268 (N_36268,N_35830,N_35531);
nor U36269 (N_36269,N_35089,N_35617);
or U36270 (N_36270,N_35715,N_35905);
nor U36271 (N_36271,N_35609,N_35433);
or U36272 (N_36272,N_35402,N_35904);
or U36273 (N_36273,N_35301,N_35987);
or U36274 (N_36274,N_35201,N_35358);
nor U36275 (N_36275,N_35241,N_35020);
or U36276 (N_36276,N_35698,N_35615);
nor U36277 (N_36277,N_35389,N_35810);
xnor U36278 (N_36278,N_35748,N_35271);
xnor U36279 (N_36279,N_35069,N_35630);
nor U36280 (N_36280,N_35140,N_35142);
xor U36281 (N_36281,N_35051,N_35976);
and U36282 (N_36282,N_35762,N_35203);
nand U36283 (N_36283,N_35393,N_35078);
nand U36284 (N_36284,N_35182,N_35775);
and U36285 (N_36285,N_35702,N_35485);
xnor U36286 (N_36286,N_35245,N_35019);
or U36287 (N_36287,N_35219,N_35419);
nor U36288 (N_36288,N_35056,N_35568);
nor U36289 (N_36289,N_35084,N_35771);
or U36290 (N_36290,N_35952,N_35833);
nor U36291 (N_36291,N_35580,N_35805);
and U36292 (N_36292,N_35916,N_35114);
nand U36293 (N_36293,N_35144,N_35073);
nor U36294 (N_36294,N_35413,N_35898);
or U36295 (N_36295,N_35104,N_35547);
xor U36296 (N_36296,N_35995,N_35224);
and U36297 (N_36297,N_35712,N_35578);
xor U36298 (N_36298,N_35442,N_35697);
or U36299 (N_36299,N_35143,N_35947);
or U36300 (N_36300,N_35497,N_35727);
nor U36301 (N_36301,N_35918,N_35471);
nor U36302 (N_36302,N_35166,N_35678);
and U36303 (N_36303,N_35385,N_35865);
nand U36304 (N_36304,N_35803,N_35881);
nand U36305 (N_36305,N_35755,N_35967);
or U36306 (N_36306,N_35807,N_35651);
and U36307 (N_36307,N_35815,N_35340);
or U36308 (N_36308,N_35255,N_35767);
nor U36309 (N_36309,N_35983,N_35677);
and U36310 (N_36310,N_35181,N_35718);
xor U36311 (N_36311,N_35753,N_35102);
nor U36312 (N_36312,N_35938,N_35639);
or U36313 (N_36313,N_35646,N_35689);
nor U36314 (N_36314,N_35896,N_35728);
xor U36315 (N_36315,N_35005,N_35094);
nor U36316 (N_36316,N_35846,N_35648);
xor U36317 (N_36317,N_35373,N_35489);
nor U36318 (N_36318,N_35411,N_35416);
or U36319 (N_36319,N_35795,N_35179);
nand U36320 (N_36320,N_35261,N_35173);
xor U36321 (N_36321,N_35838,N_35167);
nand U36322 (N_36322,N_35944,N_35007);
xnor U36323 (N_36323,N_35716,N_35878);
nand U36324 (N_36324,N_35931,N_35997);
and U36325 (N_36325,N_35824,N_35296);
nor U36326 (N_36326,N_35574,N_35730);
xnor U36327 (N_36327,N_35467,N_35039);
nand U36328 (N_36328,N_35082,N_35445);
and U36329 (N_36329,N_35683,N_35437);
and U36330 (N_36330,N_35668,N_35146);
and U36331 (N_36331,N_35022,N_35400);
nor U36332 (N_36332,N_35487,N_35582);
and U36333 (N_36333,N_35988,N_35072);
nor U36334 (N_36334,N_35842,N_35164);
nand U36335 (N_36335,N_35958,N_35108);
nand U36336 (N_36336,N_35311,N_35823);
xnor U36337 (N_36337,N_35647,N_35306);
nor U36338 (N_36338,N_35566,N_35884);
and U36339 (N_36339,N_35095,N_35499);
xor U36340 (N_36340,N_35681,N_35811);
and U36341 (N_36341,N_35066,N_35345);
nor U36342 (N_36342,N_35390,N_35425);
nand U36343 (N_36343,N_35130,N_35616);
nand U36344 (N_36344,N_35751,N_35386);
nand U36345 (N_36345,N_35543,N_35901);
nor U36346 (N_36346,N_35183,N_35109);
or U36347 (N_36347,N_35162,N_35610);
nand U36348 (N_36348,N_35065,N_35248);
nor U36349 (N_36349,N_35307,N_35581);
nand U36350 (N_36350,N_35608,N_35230);
nor U36351 (N_36351,N_35644,N_35067);
and U36352 (N_36352,N_35141,N_35199);
and U36353 (N_36353,N_35954,N_35998);
xnor U36354 (N_36354,N_35251,N_35189);
or U36355 (N_36355,N_35936,N_35885);
and U36356 (N_36356,N_35495,N_35093);
nor U36357 (N_36357,N_35859,N_35575);
and U36358 (N_36358,N_35607,N_35354);
nand U36359 (N_36359,N_35486,N_35695);
nor U36360 (N_36360,N_35232,N_35694);
nand U36361 (N_36361,N_35193,N_35176);
nand U36362 (N_36362,N_35139,N_35785);
nor U36363 (N_36363,N_35427,N_35832);
nand U36364 (N_36364,N_35496,N_35667);
nor U36365 (N_36365,N_35817,N_35545);
and U36366 (N_36366,N_35461,N_35175);
nor U36367 (N_36367,N_35927,N_35745);
or U36368 (N_36368,N_35283,N_35514);
xnor U36369 (N_36369,N_35605,N_35326);
and U36370 (N_36370,N_35588,N_35511);
xor U36371 (N_36371,N_35525,N_35754);
nor U36372 (N_36372,N_35068,N_35169);
xor U36373 (N_36373,N_35426,N_35849);
nor U36374 (N_36374,N_35028,N_35969);
nand U36375 (N_36375,N_35611,N_35650);
or U36376 (N_36376,N_35097,N_35191);
nor U36377 (N_36377,N_35120,N_35170);
and U36378 (N_36378,N_35880,N_35417);
xnor U36379 (N_36379,N_35776,N_35922);
xnor U36380 (N_36380,N_35655,N_35229);
nor U36381 (N_36381,N_35374,N_35291);
nor U36382 (N_36382,N_35381,N_35851);
nand U36383 (N_36383,N_35964,N_35030);
and U36384 (N_36384,N_35016,N_35498);
nand U36385 (N_36385,N_35329,N_35747);
xnor U36386 (N_36386,N_35076,N_35453);
nor U36387 (N_36387,N_35165,N_35135);
or U36388 (N_36388,N_35980,N_35244);
or U36389 (N_36389,N_35258,N_35686);
nor U36390 (N_36390,N_35012,N_35396);
and U36391 (N_36391,N_35634,N_35549);
or U36392 (N_36392,N_35122,N_35886);
or U36393 (N_36393,N_35395,N_35327);
and U36394 (N_36394,N_35059,N_35765);
and U36395 (N_36395,N_35272,N_35758);
xnor U36396 (N_36396,N_35188,N_35318);
nand U36397 (N_36397,N_35946,N_35428);
and U36398 (N_36398,N_35602,N_35312);
xor U36399 (N_36399,N_35692,N_35220);
or U36400 (N_36400,N_35273,N_35552);
nor U36401 (N_36401,N_35502,N_35863);
and U36402 (N_36402,N_35752,N_35981);
xnor U36403 (N_36403,N_35414,N_35840);
and U36404 (N_36404,N_35909,N_35600);
nor U36405 (N_36405,N_35288,N_35570);
or U36406 (N_36406,N_35719,N_35799);
and U36407 (N_36407,N_35444,N_35222);
or U36408 (N_36408,N_35772,N_35333);
nor U36409 (N_36409,N_35383,N_35001);
nand U36410 (N_36410,N_35928,N_35026);
nand U36411 (N_36411,N_35257,N_35670);
nor U36412 (N_36412,N_35180,N_35061);
nor U36413 (N_36413,N_35541,N_35482);
nand U36414 (N_36414,N_35827,N_35579);
or U36415 (N_36415,N_35756,N_35298);
nand U36416 (N_36416,N_35192,N_35820);
xor U36417 (N_36417,N_35504,N_35060);
nor U36418 (N_36418,N_35860,N_35713);
nand U36419 (N_36419,N_35757,N_35371);
or U36420 (N_36420,N_35945,N_35921);
nand U36421 (N_36421,N_35452,N_35205);
nor U36422 (N_36422,N_35891,N_35773);
xor U36423 (N_36423,N_35360,N_35687);
and U36424 (N_36424,N_35550,N_35472);
nand U36425 (N_36425,N_35086,N_35657);
nor U36426 (N_36426,N_35265,N_35468);
or U36427 (N_36427,N_35999,N_35900);
or U36428 (N_36428,N_35366,N_35460);
or U36429 (N_36429,N_35070,N_35902);
nor U36430 (N_36430,N_35483,N_35044);
nand U36431 (N_36431,N_35923,N_35038);
nand U36432 (N_36432,N_35604,N_35951);
nor U36433 (N_36433,N_35159,N_35586);
and U36434 (N_36434,N_35876,N_35408);
nor U36435 (N_36435,N_35903,N_35151);
nand U36436 (N_36436,N_35955,N_35861);
xnor U36437 (N_36437,N_35950,N_35195);
nand U36438 (N_36438,N_35405,N_35770);
or U36439 (N_36439,N_35870,N_35858);
and U36440 (N_36440,N_35734,N_35096);
nor U36441 (N_36441,N_35448,N_35883);
or U36442 (N_36442,N_35285,N_35137);
or U36443 (N_36443,N_35372,N_35977);
nor U36444 (N_36444,N_35664,N_35959);
nand U36445 (N_36445,N_35920,N_35894);
nor U36446 (N_36446,N_35420,N_35276);
or U36447 (N_36447,N_35982,N_35003);
or U36448 (N_36448,N_35290,N_35551);
or U36449 (N_36449,N_35233,N_35933);
or U36450 (N_36450,N_35515,N_35690);
nand U36451 (N_36451,N_35534,N_35438);
nor U36452 (N_36452,N_35021,N_35054);
or U36453 (N_36453,N_35890,N_35401);
and U36454 (N_36454,N_35696,N_35724);
nor U36455 (N_36455,N_35436,N_35025);
xnor U36456 (N_36456,N_35606,N_35209);
and U36457 (N_36457,N_35571,N_35877);
nor U36458 (N_36458,N_35869,N_35178);
or U36459 (N_36459,N_35380,N_35218);
nand U36460 (N_36460,N_35722,N_35484);
nand U36461 (N_36461,N_35126,N_35440);
nor U36462 (N_36462,N_35782,N_35317);
xnor U36463 (N_36463,N_35638,N_35737);
nand U36464 (N_36464,N_35679,N_35984);
nand U36465 (N_36465,N_35331,N_35410);
nor U36466 (N_36466,N_35294,N_35336);
nand U36467 (N_36467,N_35300,N_35680);
or U36468 (N_36468,N_35705,N_35653);
nor U36469 (N_36469,N_35174,N_35825);
nor U36470 (N_36470,N_35212,N_35357);
xor U36471 (N_36471,N_35546,N_35190);
xor U36472 (N_36472,N_35788,N_35049);
or U36473 (N_36473,N_35033,N_35621);
nand U36474 (N_36474,N_35645,N_35699);
nor U36475 (N_36475,N_35375,N_35783);
nand U36476 (N_36476,N_35421,N_35206);
or U36477 (N_36477,N_35268,N_35800);
nand U36478 (N_36478,N_35204,N_35867);
xnor U36479 (N_36479,N_35742,N_35971);
nor U36480 (N_36480,N_35569,N_35369);
nand U36481 (N_36481,N_35221,N_35370);
nor U36482 (N_36482,N_35106,N_35134);
nand U36483 (N_36483,N_35494,N_35158);
nor U36484 (N_36484,N_35892,N_35996);
nor U36485 (N_36485,N_35564,N_35154);
nor U36486 (N_36486,N_35688,N_35009);
xor U36487 (N_36487,N_35643,N_35308);
xnor U36488 (N_36488,N_35873,N_35286);
xnor U36489 (N_36489,N_35359,N_35202);
xnor U36490 (N_36490,N_35429,N_35119);
nand U36491 (N_36491,N_35295,N_35226);
xnor U36492 (N_36492,N_35597,N_35659);
or U36493 (N_36493,N_35091,N_35293);
nand U36494 (N_36494,N_35237,N_35665);
or U36495 (N_36495,N_35957,N_35975);
and U36496 (N_36496,N_35387,N_35937);
and U36497 (N_36497,N_35313,N_35252);
or U36498 (N_36498,N_35972,N_35893);
or U36499 (N_36499,N_35925,N_35297);
and U36500 (N_36500,N_35529,N_35057);
or U36501 (N_36501,N_35477,N_35344);
and U36502 (N_36502,N_35521,N_35148);
nand U36503 (N_36503,N_35797,N_35266);
nor U36504 (N_36504,N_35490,N_35471);
nor U36505 (N_36505,N_35979,N_35217);
nand U36506 (N_36506,N_35337,N_35934);
xor U36507 (N_36507,N_35269,N_35488);
or U36508 (N_36508,N_35858,N_35456);
nor U36509 (N_36509,N_35718,N_35149);
xor U36510 (N_36510,N_35226,N_35718);
and U36511 (N_36511,N_35208,N_35377);
and U36512 (N_36512,N_35098,N_35683);
nand U36513 (N_36513,N_35088,N_35625);
and U36514 (N_36514,N_35651,N_35624);
nor U36515 (N_36515,N_35273,N_35969);
and U36516 (N_36516,N_35410,N_35612);
xnor U36517 (N_36517,N_35653,N_35467);
nand U36518 (N_36518,N_35607,N_35946);
or U36519 (N_36519,N_35926,N_35555);
xor U36520 (N_36520,N_35935,N_35222);
xor U36521 (N_36521,N_35707,N_35459);
and U36522 (N_36522,N_35236,N_35580);
and U36523 (N_36523,N_35823,N_35080);
nor U36524 (N_36524,N_35373,N_35125);
or U36525 (N_36525,N_35066,N_35159);
nor U36526 (N_36526,N_35714,N_35146);
nand U36527 (N_36527,N_35813,N_35474);
or U36528 (N_36528,N_35383,N_35480);
nor U36529 (N_36529,N_35551,N_35145);
or U36530 (N_36530,N_35326,N_35169);
nand U36531 (N_36531,N_35546,N_35239);
nor U36532 (N_36532,N_35376,N_35039);
nand U36533 (N_36533,N_35288,N_35304);
and U36534 (N_36534,N_35961,N_35896);
xnor U36535 (N_36535,N_35929,N_35452);
or U36536 (N_36536,N_35393,N_35796);
or U36537 (N_36537,N_35003,N_35019);
and U36538 (N_36538,N_35879,N_35107);
nor U36539 (N_36539,N_35251,N_35403);
nand U36540 (N_36540,N_35473,N_35986);
nand U36541 (N_36541,N_35675,N_35665);
nand U36542 (N_36542,N_35861,N_35590);
or U36543 (N_36543,N_35694,N_35261);
nand U36544 (N_36544,N_35877,N_35911);
and U36545 (N_36545,N_35683,N_35939);
nand U36546 (N_36546,N_35203,N_35244);
and U36547 (N_36547,N_35620,N_35602);
nand U36548 (N_36548,N_35749,N_35714);
or U36549 (N_36549,N_35583,N_35753);
nor U36550 (N_36550,N_35331,N_35193);
nand U36551 (N_36551,N_35516,N_35265);
nor U36552 (N_36552,N_35305,N_35121);
and U36553 (N_36553,N_35251,N_35538);
nand U36554 (N_36554,N_35910,N_35154);
nand U36555 (N_36555,N_35453,N_35373);
xor U36556 (N_36556,N_35933,N_35602);
xnor U36557 (N_36557,N_35484,N_35864);
xor U36558 (N_36558,N_35661,N_35275);
and U36559 (N_36559,N_35291,N_35818);
nor U36560 (N_36560,N_35908,N_35520);
and U36561 (N_36561,N_35655,N_35318);
and U36562 (N_36562,N_35037,N_35924);
xor U36563 (N_36563,N_35079,N_35034);
nand U36564 (N_36564,N_35881,N_35387);
and U36565 (N_36565,N_35614,N_35318);
and U36566 (N_36566,N_35317,N_35385);
and U36567 (N_36567,N_35314,N_35906);
or U36568 (N_36568,N_35161,N_35112);
and U36569 (N_36569,N_35941,N_35196);
nor U36570 (N_36570,N_35514,N_35542);
nor U36571 (N_36571,N_35383,N_35070);
and U36572 (N_36572,N_35143,N_35434);
nand U36573 (N_36573,N_35886,N_35363);
nor U36574 (N_36574,N_35072,N_35034);
xnor U36575 (N_36575,N_35691,N_35351);
or U36576 (N_36576,N_35428,N_35242);
or U36577 (N_36577,N_35881,N_35668);
nand U36578 (N_36578,N_35582,N_35726);
nor U36579 (N_36579,N_35265,N_35534);
xnor U36580 (N_36580,N_35934,N_35701);
nor U36581 (N_36581,N_35046,N_35237);
nand U36582 (N_36582,N_35277,N_35639);
xnor U36583 (N_36583,N_35195,N_35305);
and U36584 (N_36584,N_35034,N_35778);
nor U36585 (N_36585,N_35208,N_35808);
and U36586 (N_36586,N_35406,N_35598);
or U36587 (N_36587,N_35103,N_35720);
nand U36588 (N_36588,N_35918,N_35695);
xor U36589 (N_36589,N_35539,N_35536);
xnor U36590 (N_36590,N_35992,N_35946);
xor U36591 (N_36591,N_35516,N_35317);
and U36592 (N_36592,N_35979,N_35658);
and U36593 (N_36593,N_35512,N_35026);
nor U36594 (N_36594,N_35125,N_35930);
nor U36595 (N_36595,N_35823,N_35899);
nand U36596 (N_36596,N_35179,N_35516);
or U36597 (N_36597,N_35818,N_35781);
and U36598 (N_36598,N_35572,N_35468);
xnor U36599 (N_36599,N_35042,N_35242);
nor U36600 (N_36600,N_35040,N_35027);
or U36601 (N_36601,N_35133,N_35930);
or U36602 (N_36602,N_35719,N_35396);
xor U36603 (N_36603,N_35190,N_35115);
nor U36604 (N_36604,N_35127,N_35380);
nor U36605 (N_36605,N_35205,N_35225);
xor U36606 (N_36606,N_35365,N_35619);
or U36607 (N_36607,N_35452,N_35976);
xor U36608 (N_36608,N_35393,N_35813);
or U36609 (N_36609,N_35632,N_35066);
nor U36610 (N_36610,N_35182,N_35524);
or U36611 (N_36611,N_35739,N_35447);
and U36612 (N_36612,N_35313,N_35162);
xnor U36613 (N_36613,N_35656,N_35845);
and U36614 (N_36614,N_35738,N_35156);
or U36615 (N_36615,N_35669,N_35589);
xnor U36616 (N_36616,N_35638,N_35867);
nor U36617 (N_36617,N_35956,N_35069);
or U36618 (N_36618,N_35106,N_35798);
and U36619 (N_36619,N_35066,N_35790);
nor U36620 (N_36620,N_35825,N_35553);
and U36621 (N_36621,N_35458,N_35303);
nor U36622 (N_36622,N_35316,N_35164);
nand U36623 (N_36623,N_35307,N_35735);
xor U36624 (N_36624,N_35214,N_35350);
xnor U36625 (N_36625,N_35697,N_35924);
nand U36626 (N_36626,N_35309,N_35846);
or U36627 (N_36627,N_35161,N_35766);
xor U36628 (N_36628,N_35568,N_35589);
xor U36629 (N_36629,N_35015,N_35884);
nand U36630 (N_36630,N_35705,N_35602);
nor U36631 (N_36631,N_35571,N_35372);
or U36632 (N_36632,N_35757,N_35579);
xnor U36633 (N_36633,N_35725,N_35052);
xnor U36634 (N_36634,N_35364,N_35377);
nor U36635 (N_36635,N_35619,N_35963);
or U36636 (N_36636,N_35463,N_35967);
xor U36637 (N_36637,N_35537,N_35747);
and U36638 (N_36638,N_35401,N_35601);
nand U36639 (N_36639,N_35079,N_35071);
nand U36640 (N_36640,N_35414,N_35631);
xor U36641 (N_36641,N_35729,N_35673);
nand U36642 (N_36642,N_35345,N_35908);
nand U36643 (N_36643,N_35954,N_35104);
and U36644 (N_36644,N_35485,N_35512);
and U36645 (N_36645,N_35066,N_35627);
nand U36646 (N_36646,N_35287,N_35055);
nand U36647 (N_36647,N_35040,N_35301);
nand U36648 (N_36648,N_35470,N_35773);
nand U36649 (N_36649,N_35685,N_35342);
xor U36650 (N_36650,N_35959,N_35600);
nor U36651 (N_36651,N_35777,N_35979);
nand U36652 (N_36652,N_35493,N_35430);
nor U36653 (N_36653,N_35676,N_35540);
nor U36654 (N_36654,N_35761,N_35109);
xor U36655 (N_36655,N_35346,N_35960);
nor U36656 (N_36656,N_35927,N_35800);
nand U36657 (N_36657,N_35906,N_35839);
and U36658 (N_36658,N_35354,N_35396);
nor U36659 (N_36659,N_35219,N_35854);
nor U36660 (N_36660,N_35856,N_35611);
nor U36661 (N_36661,N_35214,N_35225);
and U36662 (N_36662,N_35342,N_35925);
and U36663 (N_36663,N_35001,N_35905);
xor U36664 (N_36664,N_35135,N_35908);
or U36665 (N_36665,N_35211,N_35187);
and U36666 (N_36666,N_35524,N_35216);
xnor U36667 (N_36667,N_35682,N_35144);
xnor U36668 (N_36668,N_35721,N_35658);
xnor U36669 (N_36669,N_35723,N_35333);
nand U36670 (N_36670,N_35218,N_35551);
nand U36671 (N_36671,N_35441,N_35114);
nor U36672 (N_36672,N_35598,N_35931);
nor U36673 (N_36673,N_35184,N_35882);
nor U36674 (N_36674,N_35898,N_35000);
and U36675 (N_36675,N_35169,N_35206);
nand U36676 (N_36676,N_35144,N_35103);
nor U36677 (N_36677,N_35523,N_35228);
nand U36678 (N_36678,N_35298,N_35934);
and U36679 (N_36679,N_35374,N_35979);
nand U36680 (N_36680,N_35038,N_35873);
or U36681 (N_36681,N_35588,N_35394);
or U36682 (N_36682,N_35539,N_35385);
and U36683 (N_36683,N_35331,N_35115);
nand U36684 (N_36684,N_35696,N_35495);
and U36685 (N_36685,N_35775,N_35470);
nand U36686 (N_36686,N_35893,N_35582);
and U36687 (N_36687,N_35170,N_35260);
nor U36688 (N_36688,N_35417,N_35864);
or U36689 (N_36689,N_35155,N_35604);
nand U36690 (N_36690,N_35416,N_35781);
nor U36691 (N_36691,N_35661,N_35900);
nand U36692 (N_36692,N_35288,N_35434);
nor U36693 (N_36693,N_35565,N_35416);
nor U36694 (N_36694,N_35287,N_35205);
and U36695 (N_36695,N_35562,N_35125);
and U36696 (N_36696,N_35824,N_35580);
xnor U36697 (N_36697,N_35504,N_35360);
and U36698 (N_36698,N_35723,N_35276);
nand U36699 (N_36699,N_35054,N_35688);
xnor U36700 (N_36700,N_35915,N_35200);
xnor U36701 (N_36701,N_35872,N_35603);
or U36702 (N_36702,N_35619,N_35821);
nor U36703 (N_36703,N_35704,N_35336);
nand U36704 (N_36704,N_35406,N_35678);
xnor U36705 (N_36705,N_35443,N_35239);
xor U36706 (N_36706,N_35677,N_35665);
nand U36707 (N_36707,N_35917,N_35367);
and U36708 (N_36708,N_35465,N_35329);
or U36709 (N_36709,N_35249,N_35068);
nor U36710 (N_36710,N_35913,N_35404);
nor U36711 (N_36711,N_35884,N_35725);
xor U36712 (N_36712,N_35127,N_35244);
nor U36713 (N_36713,N_35073,N_35014);
xnor U36714 (N_36714,N_35899,N_35446);
nor U36715 (N_36715,N_35112,N_35545);
nor U36716 (N_36716,N_35960,N_35425);
xor U36717 (N_36717,N_35500,N_35677);
or U36718 (N_36718,N_35597,N_35494);
and U36719 (N_36719,N_35411,N_35429);
or U36720 (N_36720,N_35490,N_35281);
nand U36721 (N_36721,N_35607,N_35635);
xnor U36722 (N_36722,N_35610,N_35894);
nor U36723 (N_36723,N_35173,N_35696);
or U36724 (N_36724,N_35758,N_35737);
nand U36725 (N_36725,N_35117,N_35438);
and U36726 (N_36726,N_35604,N_35067);
nand U36727 (N_36727,N_35024,N_35952);
nor U36728 (N_36728,N_35983,N_35354);
nor U36729 (N_36729,N_35332,N_35020);
xor U36730 (N_36730,N_35611,N_35194);
nor U36731 (N_36731,N_35843,N_35723);
nor U36732 (N_36732,N_35602,N_35031);
xnor U36733 (N_36733,N_35417,N_35646);
nand U36734 (N_36734,N_35354,N_35379);
nor U36735 (N_36735,N_35556,N_35728);
or U36736 (N_36736,N_35794,N_35776);
xor U36737 (N_36737,N_35900,N_35787);
xor U36738 (N_36738,N_35525,N_35212);
xor U36739 (N_36739,N_35906,N_35069);
and U36740 (N_36740,N_35069,N_35300);
nand U36741 (N_36741,N_35025,N_35330);
nand U36742 (N_36742,N_35316,N_35768);
nor U36743 (N_36743,N_35813,N_35080);
nand U36744 (N_36744,N_35999,N_35859);
or U36745 (N_36745,N_35328,N_35074);
or U36746 (N_36746,N_35554,N_35939);
and U36747 (N_36747,N_35237,N_35304);
nand U36748 (N_36748,N_35858,N_35751);
and U36749 (N_36749,N_35437,N_35570);
or U36750 (N_36750,N_35674,N_35161);
xnor U36751 (N_36751,N_35717,N_35459);
xnor U36752 (N_36752,N_35375,N_35087);
nand U36753 (N_36753,N_35879,N_35272);
or U36754 (N_36754,N_35921,N_35213);
xor U36755 (N_36755,N_35063,N_35587);
nor U36756 (N_36756,N_35683,N_35514);
nand U36757 (N_36757,N_35291,N_35937);
and U36758 (N_36758,N_35713,N_35104);
and U36759 (N_36759,N_35944,N_35053);
nor U36760 (N_36760,N_35371,N_35270);
or U36761 (N_36761,N_35870,N_35826);
and U36762 (N_36762,N_35560,N_35281);
nor U36763 (N_36763,N_35948,N_35677);
and U36764 (N_36764,N_35106,N_35456);
xor U36765 (N_36765,N_35444,N_35096);
nor U36766 (N_36766,N_35156,N_35779);
xnor U36767 (N_36767,N_35729,N_35896);
nand U36768 (N_36768,N_35121,N_35482);
nand U36769 (N_36769,N_35248,N_35672);
nand U36770 (N_36770,N_35821,N_35706);
and U36771 (N_36771,N_35803,N_35897);
nand U36772 (N_36772,N_35835,N_35623);
and U36773 (N_36773,N_35086,N_35773);
or U36774 (N_36774,N_35833,N_35236);
or U36775 (N_36775,N_35154,N_35321);
and U36776 (N_36776,N_35004,N_35849);
xor U36777 (N_36777,N_35800,N_35505);
nand U36778 (N_36778,N_35997,N_35364);
nand U36779 (N_36779,N_35745,N_35363);
xor U36780 (N_36780,N_35270,N_35655);
and U36781 (N_36781,N_35292,N_35819);
and U36782 (N_36782,N_35245,N_35790);
or U36783 (N_36783,N_35127,N_35008);
and U36784 (N_36784,N_35314,N_35549);
nand U36785 (N_36785,N_35926,N_35899);
nand U36786 (N_36786,N_35685,N_35834);
and U36787 (N_36787,N_35302,N_35692);
nor U36788 (N_36788,N_35944,N_35028);
xnor U36789 (N_36789,N_35892,N_35440);
nor U36790 (N_36790,N_35396,N_35956);
or U36791 (N_36791,N_35751,N_35609);
nand U36792 (N_36792,N_35652,N_35399);
xnor U36793 (N_36793,N_35042,N_35946);
xnor U36794 (N_36794,N_35553,N_35375);
or U36795 (N_36795,N_35796,N_35123);
or U36796 (N_36796,N_35953,N_35706);
nand U36797 (N_36797,N_35824,N_35919);
or U36798 (N_36798,N_35928,N_35456);
or U36799 (N_36799,N_35956,N_35067);
xnor U36800 (N_36800,N_35547,N_35406);
nand U36801 (N_36801,N_35248,N_35192);
or U36802 (N_36802,N_35237,N_35329);
nor U36803 (N_36803,N_35112,N_35500);
or U36804 (N_36804,N_35258,N_35209);
xnor U36805 (N_36805,N_35636,N_35604);
xor U36806 (N_36806,N_35834,N_35609);
or U36807 (N_36807,N_35449,N_35377);
nor U36808 (N_36808,N_35097,N_35872);
nor U36809 (N_36809,N_35237,N_35400);
or U36810 (N_36810,N_35026,N_35733);
nand U36811 (N_36811,N_35647,N_35011);
and U36812 (N_36812,N_35094,N_35242);
or U36813 (N_36813,N_35516,N_35205);
and U36814 (N_36814,N_35844,N_35468);
or U36815 (N_36815,N_35754,N_35846);
or U36816 (N_36816,N_35794,N_35581);
nor U36817 (N_36817,N_35693,N_35223);
or U36818 (N_36818,N_35965,N_35422);
nand U36819 (N_36819,N_35252,N_35368);
or U36820 (N_36820,N_35397,N_35462);
or U36821 (N_36821,N_35163,N_35638);
or U36822 (N_36822,N_35381,N_35667);
nand U36823 (N_36823,N_35484,N_35861);
xor U36824 (N_36824,N_35898,N_35657);
nand U36825 (N_36825,N_35428,N_35290);
xor U36826 (N_36826,N_35629,N_35945);
nand U36827 (N_36827,N_35586,N_35851);
nor U36828 (N_36828,N_35610,N_35643);
nor U36829 (N_36829,N_35673,N_35525);
or U36830 (N_36830,N_35546,N_35247);
xnor U36831 (N_36831,N_35261,N_35493);
nand U36832 (N_36832,N_35508,N_35037);
xnor U36833 (N_36833,N_35463,N_35827);
nor U36834 (N_36834,N_35124,N_35693);
xnor U36835 (N_36835,N_35809,N_35471);
nand U36836 (N_36836,N_35152,N_35916);
or U36837 (N_36837,N_35440,N_35648);
nor U36838 (N_36838,N_35662,N_35689);
xor U36839 (N_36839,N_35944,N_35739);
or U36840 (N_36840,N_35613,N_35333);
nor U36841 (N_36841,N_35046,N_35388);
and U36842 (N_36842,N_35802,N_35792);
nor U36843 (N_36843,N_35926,N_35257);
nor U36844 (N_36844,N_35918,N_35624);
nor U36845 (N_36845,N_35813,N_35800);
and U36846 (N_36846,N_35113,N_35145);
xor U36847 (N_36847,N_35663,N_35139);
or U36848 (N_36848,N_35610,N_35762);
and U36849 (N_36849,N_35478,N_35374);
and U36850 (N_36850,N_35760,N_35312);
and U36851 (N_36851,N_35051,N_35573);
and U36852 (N_36852,N_35521,N_35669);
or U36853 (N_36853,N_35688,N_35782);
and U36854 (N_36854,N_35416,N_35229);
or U36855 (N_36855,N_35752,N_35412);
xnor U36856 (N_36856,N_35556,N_35877);
nand U36857 (N_36857,N_35442,N_35187);
and U36858 (N_36858,N_35454,N_35915);
nand U36859 (N_36859,N_35686,N_35801);
or U36860 (N_36860,N_35350,N_35042);
or U36861 (N_36861,N_35666,N_35299);
xnor U36862 (N_36862,N_35664,N_35068);
xnor U36863 (N_36863,N_35465,N_35025);
nor U36864 (N_36864,N_35789,N_35150);
nand U36865 (N_36865,N_35357,N_35780);
nand U36866 (N_36866,N_35444,N_35691);
xor U36867 (N_36867,N_35758,N_35851);
or U36868 (N_36868,N_35141,N_35786);
nor U36869 (N_36869,N_35001,N_35759);
nand U36870 (N_36870,N_35028,N_35494);
xnor U36871 (N_36871,N_35813,N_35422);
nor U36872 (N_36872,N_35845,N_35619);
or U36873 (N_36873,N_35041,N_35410);
or U36874 (N_36874,N_35108,N_35327);
or U36875 (N_36875,N_35707,N_35265);
or U36876 (N_36876,N_35745,N_35015);
or U36877 (N_36877,N_35164,N_35240);
nor U36878 (N_36878,N_35272,N_35812);
and U36879 (N_36879,N_35502,N_35517);
nor U36880 (N_36880,N_35277,N_35650);
nor U36881 (N_36881,N_35809,N_35411);
and U36882 (N_36882,N_35911,N_35081);
and U36883 (N_36883,N_35495,N_35786);
xor U36884 (N_36884,N_35565,N_35807);
and U36885 (N_36885,N_35371,N_35597);
nand U36886 (N_36886,N_35184,N_35303);
and U36887 (N_36887,N_35698,N_35256);
nor U36888 (N_36888,N_35214,N_35709);
and U36889 (N_36889,N_35825,N_35658);
nand U36890 (N_36890,N_35779,N_35354);
xor U36891 (N_36891,N_35773,N_35099);
and U36892 (N_36892,N_35743,N_35074);
or U36893 (N_36893,N_35478,N_35151);
nand U36894 (N_36894,N_35256,N_35476);
and U36895 (N_36895,N_35112,N_35829);
and U36896 (N_36896,N_35203,N_35563);
nor U36897 (N_36897,N_35607,N_35792);
and U36898 (N_36898,N_35969,N_35497);
nand U36899 (N_36899,N_35932,N_35522);
nand U36900 (N_36900,N_35097,N_35946);
nand U36901 (N_36901,N_35833,N_35536);
or U36902 (N_36902,N_35470,N_35851);
nand U36903 (N_36903,N_35592,N_35865);
and U36904 (N_36904,N_35430,N_35279);
nor U36905 (N_36905,N_35136,N_35991);
xnor U36906 (N_36906,N_35506,N_35396);
and U36907 (N_36907,N_35124,N_35220);
or U36908 (N_36908,N_35715,N_35348);
and U36909 (N_36909,N_35986,N_35195);
and U36910 (N_36910,N_35954,N_35097);
and U36911 (N_36911,N_35223,N_35686);
xor U36912 (N_36912,N_35482,N_35863);
nor U36913 (N_36913,N_35951,N_35296);
or U36914 (N_36914,N_35267,N_35183);
nor U36915 (N_36915,N_35731,N_35548);
and U36916 (N_36916,N_35478,N_35501);
and U36917 (N_36917,N_35493,N_35654);
nand U36918 (N_36918,N_35449,N_35980);
nor U36919 (N_36919,N_35299,N_35203);
or U36920 (N_36920,N_35247,N_35946);
nor U36921 (N_36921,N_35244,N_35553);
nor U36922 (N_36922,N_35037,N_35122);
or U36923 (N_36923,N_35413,N_35903);
or U36924 (N_36924,N_35231,N_35923);
nand U36925 (N_36925,N_35287,N_35251);
or U36926 (N_36926,N_35079,N_35133);
nand U36927 (N_36927,N_35553,N_35550);
nor U36928 (N_36928,N_35309,N_35150);
nand U36929 (N_36929,N_35794,N_35994);
and U36930 (N_36930,N_35680,N_35858);
nor U36931 (N_36931,N_35680,N_35981);
nand U36932 (N_36932,N_35908,N_35587);
nand U36933 (N_36933,N_35029,N_35577);
nor U36934 (N_36934,N_35366,N_35386);
and U36935 (N_36935,N_35159,N_35578);
and U36936 (N_36936,N_35080,N_35231);
nor U36937 (N_36937,N_35026,N_35560);
and U36938 (N_36938,N_35829,N_35979);
nand U36939 (N_36939,N_35709,N_35269);
xor U36940 (N_36940,N_35008,N_35011);
nor U36941 (N_36941,N_35485,N_35744);
nor U36942 (N_36942,N_35529,N_35336);
xnor U36943 (N_36943,N_35586,N_35377);
xnor U36944 (N_36944,N_35736,N_35309);
or U36945 (N_36945,N_35632,N_35922);
or U36946 (N_36946,N_35613,N_35524);
or U36947 (N_36947,N_35186,N_35524);
and U36948 (N_36948,N_35220,N_35391);
or U36949 (N_36949,N_35057,N_35339);
nand U36950 (N_36950,N_35919,N_35618);
nand U36951 (N_36951,N_35117,N_35874);
and U36952 (N_36952,N_35780,N_35566);
nand U36953 (N_36953,N_35846,N_35349);
and U36954 (N_36954,N_35249,N_35288);
and U36955 (N_36955,N_35829,N_35872);
and U36956 (N_36956,N_35596,N_35242);
or U36957 (N_36957,N_35908,N_35496);
nand U36958 (N_36958,N_35077,N_35729);
xnor U36959 (N_36959,N_35176,N_35337);
and U36960 (N_36960,N_35042,N_35873);
and U36961 (N_36961,N_35124,N_35769);
xnor U36962 (N_36962,N_35725,N_35044);
nand U36963 (N_36963,N_35877,N_35025);
and U36964 (N_36964,N_35564,N_35787);
or U36965 (N_36965,N_35146,N_35789);
or U36966 (N_36966,N_35882,N_35234);
nor U36967 (N_36967,N_35743,N_35350);
nand U36968 (N_36968,N_35159,N_35074);
or U36969 (N_36969,N_35911,N_35084);
and U36970 (N_36970,N_35804,N_35749);
nand U36971 (N_36971,N_35396,N_35442);
and U36972 (N_36972,N_35793,N_35674);
xnor U36973 (N_36973,N_35584,N_35478);
xor U36974 (N_36974,N_35032,N_35965);
xnor U36975 (N_36975,N_35858,N_35953);
xor U36976 (N_36976,N_35702,N_35806);
nor U36977 (N_36977,N_35038,N_35461);
nor U36978 (N_36978,N_35028,N_35948);
nand U36979 (N_36979,N_35343,N_35394);
nand U36980 (N_36980,N_35372,N_35711);
nor U36981 (N_36981,N_35055,N_35156);
and U36982 (N_36982,N_35814,N_35215);
nor U36983 (N_36983,N_35395,N_35717);
and U36984 (N_36984,N_35942,N_35023);
or U36985 (N_36985,N_35477,N_35976);
and U36986 (N_36986,N_35626,N_35940);
nand U36987 (N_36987,N_35458,N_35497);
or U36988 (N_36988,N_35887,N_35828);
nor U36989 (N_36989,N_35021,N_35636);
xor U36990 (N_36990,N_35695,N_35546);
nand U36991 (N_36991,N_35371,N_35219);
or U36992 (N_36992,N_35759,N_35517);
nor U36993 (N_36993,N_35977,N_35148);
xnor U36994 (N_36994,N_35672,N_35859);
and U36995 (N_36995,N_35055,N_35602);
and U36996 (N_36996,N_35673,N_35568);
xor U36997 (N_36997,N_35110,N_35750);
xnor U36998 (N_36998,N_35687,N_35923);
and U36999 (N_36999,N_35995,N_35762);
nor U37000 (N_37000,N_36986,N_36039);
or U37001 (N_37001,N_36655,N_36709);
nor U37002 (N_37002,N_36406,N_36001);
or U37003 (N_37003,N_36616,N_36314);
xor U37004 (N_37004,N_36121,N_36016);
nor U37005 (N_37005,N_36831,N_36288);
and U37006 (N_37006,N_36832,N_36952);
nor U37007 (N_37007,N_36034,N_36434);
nor U37008 (N_37008,N_36094,N_36522);
or U37009 (N_37009,N_36764,N_36767);
xor U37010 (N_37010,N_36186,N_36460);
and U37011 (N_37011,N_36851,N_36752);
nor U37012 (N_37012,N_36865,N_36221);
nor U37013 (N_37013,N_36961,N_36141);
xnor U37014 (N_37014,N_36231,N_36134);
nor U37015 (N_37015,N_36159,N_36942);
and U37016 (N_37016,N_36305,N_36618);
nand U37017 (N_37017,N_36349,N_36586);
nand U37018 (N_37018,N_36276,N_36868);
xor U37019 (N_37019,N_36523,N_36418);
and U37020 (N_37020,N_36935,N_36053);
xor U37021 (N_37021,N_36949,N_36481);
and U37022 (N_37022,N_36504,N_36313);
and U37023 (N_37023,N_36341,N_36172);
xnor U37024 (N_37024,N_36720,N_36739);
nor U37025 (N_37025,N_36240,N_36369);
xnor U37026 (N_37026,N_36258,N_36363);
nor U37027 (N_37027,N_36223,N_36754);
or U37028 (N_37028,N_36042,N_36749);
or U37029 (N_37029,N_36465,N_36253);
xnor U37030 (N_37030,N_36782,N_36913);
nand U37031 (N_37031,N_36660,N_36945);
nor U37032 (N_37032,N_36807,N_36642);
or U37033 (N_37033,N_36352,N_36312);
xor U37034 (N_37034,N_36297,N_36975);
or U37035 (N_37035,N_36774,N_36862);
xor U37036 (N_37036,N_36430,N_36537);
and U37037 (N_37037,N_36023,N_36694);
nand U37038 (N_37038,N_36155,N_36948);
and U37039 (N_37039,N_36462,N_36909);
nand U37040 (N_37040,N_36714,N_36315);
nand U37041 (N_37041,N_36981,N_36735);
nor U37042 (N_37042,N_36367,N_36557);
xor U37043 (N_37043,N_36347,N_36741);
and U37044 (N_37044,N_36579,N_36968);
or U37045 (N_37045,N_36004,N_36974);
or U37046 (N_37046,N_36792,N_36959);
or U37047 (N_37047,N_36317,N_36476);
nand U37048 (N_37048,N_36753,N_36407);
nor U37049 (N_37049,N_36609,N_36489);
nor U37050 (N_37050,N_36459,N_36610);
nor U37051 (N_37051,N_36002,N_36771);
and U37052 (N_37052,N_36812,N_36860);
or U37053 (N_37053,N_36473,N_36021);
nor U37054 (N_37054,N_36561,N_36037);
nand U37055 (N_37055,N_36874,N_36378);
and U37056 (N_37056,N_36237,N_36491);
and U37057 (N_37057,N_36403,N_36553);
and U37058 (N_37058,N_36301,N_36057);
nor U37059 (N_37059,N_36259,N_36078);
xor U37060 (N_37060,N_36951,N_36166);
xnor U37061 (N_37061,N_36687,N_36116);
nor U37062 (N_37062,N_36101,N_36711);
and U37063 (N_37063,N_36992,N_36869);
or U37064 (N_37064,N_36925,N_36666);
and U37065 (N_37065,N_36806,N_36766);
and U37066 (N_37066,N_36988,N_36697);
or U37067 (N_37067,N_36559,N_36306);
or U37068 (N_37068,N_36146,N_36632);
nor U37069 (N_37069,N_36484,N_36630);
nor U37070 (N_37070,N_36379,N_36814);
nand U37071 (N_37071,N_36939,N_36052);
nand U37072 (N_37072,N_36744,N_36878);
or U37073 (N_37073,N_36490,N_36229);
and U37074 (N_37074,N_36442,N_36128);
and U37075 (N_37075,N_36117,N_36415);
and U37076 (N_37076,N_36745,N_36839);
xor U37077 (N_37077,N_36419,N_36947);
or U37078 (N_37078,N_36220,N_36692);
xor U37079 (N_37079,N_36040,N_36244);
and U37080 (N_37080,N_36092,N_36905);
or U37081 (N_37081,N_36800,N_36990);
nor U37082 (N_37082,N_36982,N_36686);
or U37083 (N_37083,N_36848,N_36989);
nor U37084 (N_37084,N_36519,N_36804);
xnor U37085 (N_37085,N_36803,N_36700);
xnor U37086 (N_37086,N_36087,N_36281);
or U37087 (N_37087,N_36396,N_36651);
nor U37088 (N_37088,N_36701,N_36929);
nor U37089 (N_37089,N_36653,N_36421);
and U37090 (N_37090,N_36728,N_36198);
nor U37091 (N_37091,N_36681,N_36693);
or U37092 (N_37092,N_36780,N_36424);
and U37093 (N_37093,N_36382,N_36012);
nor U37094 (N_37094,N_36090,N_36556);
nand U37095 (N_37095,N_36026,N_36723);
nand U37096 (N_37096,N_36420,N_36359);
xor U37097 (N_37097,N_36480,N_36167);
and U37098 (N_37098,N_36102,N_36156);
or U37099 (N_37099,N_36993,N_36309);
xor U37100 (N_37100,N_36280,N_36602);
or U37101 (N_37101,N_36902,N_36824);
xnor U37102 (N_37102,N_36818,N_36987);
and U37103 (N_37103,N_36985,N_36232);
nor U37104 (N_37104,N_36033,N_36149);
nor U37105 (N_37105,N_36154,N_36132);
and U37106 (N_37106,N_36544,N_36597);
or U37107 (N_37107,N_36938,N_36944);
or U37108 (N_37108,N_36724,N_36842);
and U37109 (N_37109,N_36150,N_36151);
and U37110 (N_37110,N_36567,N_36410);
or U37111 (N_37111,N_36010,N_36113);
nand U37112 (N_37112,N_36670,N_36950);
nand U37113 (N_37113,N_36289,N_36955);
xor U37114 (N_37114,N_36699,N_36748);
nand U37115 (N_37115,N_36546,N_36737);
nor U37116 (N_37116,N_36734,N_36717);
nor U37117 (N_37117,N_36494,N_36196);
or U37118 (N_37118,N_36177,N_36405);
xor U37119 (N_37119,N_36066,N_36520);
xnor U37120 (N_37120,N_36067,N_36552);
nor U37121 (N_37121,N_36661,N_36168);
nor U37122 (N_37122,N_36847,N_36511);
nand U37123 (N_37123,N_36174,N_36471);
nand U37124 (N_37124,N_36917,N_36370);
xor U37125 (N_37125,N_36592,N_36999);
or U37126 (N_37126,N_36696,N_36008);
or U37127 (N_37127,N_36380,N_36477);
nand U37128 (N_37128,N_36345,N_36801);
nor U37129 (N_37129,N_36227,N_36844);
or U37130 (N_37130,N_36742,N_36215);
and U37131 (N_37131,N_36608,N_36773);
or U37132 (N_37132,N_36098,N_36384);
nand U37133 (N_37133,N_36498,N_36269);
nand U37134 (N_37134,N_36123,N_36996);
or U37135 (N_37135,N_36152,N_36550);
nand U37136 (N_37136,N_36809,N_36295);
or U37137 (N_37137,N_36184,N_36136);
or U37138 (N_37138,N_36126,N_36303);
or U37139 (N_37139,N_36487,N_36643);
and U37140 (N_37140,N_36075,N_36147);
nor U37141 (N_37141,N_36542,N_36482);
or U37142 (N_37142,N_36387,N_36903);
xnor U37143 (N_37143,N_36401,N_36855);
or U37144 (N_37144,N_36083,N_36346);
and U37145 (N_37145,N_36810,N_36298);
and U37146 (N_37146,N_36680,N_36648);
nor U37147 (N_37147,N_36843,N_36617);
and U37148 (N_37148,N_36390,N_36912);
nor U37149 (N_37149,N_36320,N_36883);
nor U37150 (N_37150,N_36516,N_36589);
and U37151 (N_37151,N_36970,N_36445);
and U37152 (N_37152,N_36762,N_36572);
or U37153 (N_37153,N_36342,N_36448);
or U37154 (N_37154,N_36331,N_36943);
xnor U37155 (N_37155,N_36203,N_36130);
or U37156 (N_37156,N_36721,N_36133);
or U37157 (N_37157,N_36059,N_36351);
nor U37158 (N_37158,N_36093,N_36554);
xor U37159 (N_37159,N_36358,N_36013);
nand U37160 (N_37160,N_36428,N_36106);
and U37161 (N_37161,N_36614,N_36551);
xor U37162 (N_37162,N_36190,N_36569);
xor U37163 (N_37163,N_36983,N_36153);
nand U37164 (N_37164,N_36475,N_36907);
or U37165 (N_37165,N_36577,N_36474);
nor U37166 (N_37166,N_36636,N_36706);
nor U37167 (N_37167,N_36901,N_36765);
or U37168 (N_37168,N_36956,N_36978);
or U37169 (N_37169,N_36266,N_36251);
or U37170 (N_37170,N_36411,N_36239);
nand U37171 (N_37171,N_36045,N_36030);
and U37172 (N_37172,N_36478,N_36645);
nor U37173 (N_37173,N_36889,N_36285);
and U37174 (N_37174,N_36658,N_36796);
and U37175 (N_37175,N_36182,N_36371);
nor U37176 (N_37176,N_36563,N_36326);
nand U37177 (N_37177,N_36056,N_36743);
or U37178 (N_37178,N_36210,N_36125);
xor U37179 (N_37179,N_36712,N_36400);
or U37180 (N_37180,N_36148,N_36169);
xor U37181 (N_37181,N_36526,N_36392);
nor U37182 (N_37182,N_36388,N_36496);
xnor U37183 (N_37183,N_36751,N_36469);
nor U37184 (N_37184,N_36657,N_36256);
xnor U37185 (N_37185,N_36896,N_36025);
nor U37186 (N_37186,N_36509,N_36207);
xor U37187 (N_37187,N_36719,N_36348);
or U37188 (N_37188,N_36871,N_36437);
nor U37189 (N_37189,N_36191,N_36815);
nor U37190 (N_37190,N_36267,N_36880);
nor U37191 (N_37191,N_36833,N_36230);
xor U37192 (N_37192,N_36882,N_36973);
and U37193 (N_37193,N_36521,N_36641);
nand U37194 (N_37194,N_36789,N_36954);
xnor U37195 (N_37195,N_36081,N_36531);
xor U37196 (N_37196,N_36911,N_36838);
or U37197 (N_37197,N_36423,N_36802);
xnor U37198 (N_37198,N_36826,N_36808);
or U37199 (N_37199,N_36571,N_36338);
or U37200 (N_37200,N_36451,N_36091);
nor U37201 (N_37201,N_36273,N_36322);
nand U37202 (N_37202,N_36513,N_36786);
and U37203 (N_37203,N_36112,N_36041);
nor U37204 (N_37204,N_36394,N_36183);
xnor U37205 (N_37205,N_36138,N_36963);
nand U37206 (N_37206,N_36931,N_36208);
or U37207 (N_37207,N_36366,N_36079);
xor U37208 (N_37208,N_36248,N_36319);
nand U37209 (N_37209,N_36715,N_36866);
or U37210 (N_37210,N_36760,N_36143);
or U37211 (N_37211,N_36547,N_36967);
nand U37212 (N_37212,N_36456,N_36199);
and U37213 (N_37213,N_36540,N_36535);
nor U37214 (N_37214,N_36890,N_36536);
xnor U37215 (N_37215,N_36611,N_36690);
or U37216 (N_37216,N_36139,N_36118);
nand U37217 (N_37217,N_36647,N_36576);
or U37218 (N_37218,N_36329,N_36127);
nand U37219 (N_37219,N_36450,N_36441);
nor U37220 (N_37220,N_36213,N_36086);
or U37221 (N_37221,N_36849,N_36212);
nor U37222 (N_37222,N_36000,N_36870);
xnor U37223 (N_37223,N_36398,N_36649);
nor U37224 (N_37224,N_36055,N_36811);
nor U37225 (N_37225,N_36747,N_36738);
or U37226 (N_37226,N_36343,N_36111);
xor U37227 (N_37227,N_36044,N_36500);
or U37228 (N_37228,N_36466,N_36404);
nor U37229 (N_37229,N_36518,N_36376);
or U37230 (N_37230,N_36575,N_36971);
nor U37231 (N_37231,N_36583,N_36875);
and U37232 (N_37232,N_36667,N_36007);
nand U37233 (N_37233,N_36375,N_36180);
or U37234 (N_37234,N_36238,N_36937);
nor U37235 (N_37235,N_36588,N_36758);
or U37236 (N_37236,N_36162,N_36485);
or U37237 (N_37237,N_36129,N_36672);
nand U37238 (N_37238,N_36827,N_36181);
or U37239 (N_37239,N_36175,N_36776);
xnor U37240 (N_37240,N_36897,N_36918);
xnor U37241 (N_37241,N_36316,N_36727);
nand U37242 (N_37242,N_36791,N_36598);
nor U37243 (N_37243,N_36570,N_36444);
or U37244 (N_37244,N_36070,N_36596);
xor U37245 (N_37245,N_36708,N_36302);
nand U37246 (N_37246,N_36282,N_36612);
nand U37247 (N_37247,N_36255,N_36080);
nand U37248 (N_37248,N_36605,N_36479);
nand U37249 (N_37249,N_36095,N_36279);
xor U37250 (N_37250,N_36054,N_36492);
and U37251 (N_37251,N_36246,N_36321);
or U37252 (N_37252,N_36644,N_36005);
nand U37253 (N_37253,N_36110,N_36355);
nor U37254 (N_37254,N_36683,N_36381);
nand U37255 (N_37255,N_36027,N_36436);
or U37256 (N_37256,N_36356,N_36409);
xor U37257 (N_37257,N_36781,N_36894);
nor U37258 (N_37258,N_36032,N_36050);
or U37259 (N_37259,N_36365,N_36145);
xor U37260 (N_37260,N_36619,N_36638);
and U37261 (N_37261,N_36922,N_36599);
nand U37262 (N_37262,N_36962,N_36881);
and U37263 (N_37263,N_36071,N_36578);
or U37264 (N_37264,N_36438,N_36665);
nand U37265 (N_37265,N_36877,N_36634);
or U37266 (N_37266,N_36958,N_36488);
or U37267 (N_37267,N_36283,N_36124);
nor U37268 (N_37268,N_36733,N_36543);
xnor U37269 (N_37269,N_36646,N_36854);
or U37270 (N_37270,N_36755,N_36333);
and U37271 (N_37271,N_36443,N_36587);
and U37272 (N_37272,N_36895,N_36820);
xor U37273 (N_37273,N_36529,N_36510);
nor U37274 (N_37274,N_36417,N_36979);
or U37275 (N_37275,N_36076,N_36506);
or U37276 (N_37276,N_36472,N_36228);
nor U37277 (N_37277,N_36447,N_36233);
xnor U37278 (N_37278,N_36627,N_36822);
and U37279 (N_37279,N_36201,N_36729);
xnor U37280 (N_37280,N_36335,N_36876);
or U37281 (N_37281,N_36217,N_36620);
nand U37282 (N_37282,N_36562,N_36656);
or U37283 (N_37283,N_36703,N_36268);
nor U37284 (N_37284,N_36364,N_36674);
nand U37285 (N_37285,N_36063,N_36157);
and U37286 (N_37286,N_36750,N_36122);
xor U37287 (N_37287,N_36062,N_36691);
nand U37288 (N_37288,N_36819,N_36386);
and U37289 (N_37289,N_36402,N_36038);
and U37290 (N_37290,N_36783,N_36399);
and U37291 (N_37291,N_36304,N_36202);
or U37292 (N_37292,N_36389,N_36416);
nor U37293 (N_37293,N_36085,N_36272);
and U37294 (N_37294,N_36624,N_36639);
nand U37295 (N_37295,N_36675,N_36082);
nand U37296 (N_37296,N_36503,N_36224);
xnor U37297 (N_37297,N_36171,N_36817);
or U37298 (N_37298,N_36964,N_36486);
xnor U37299 (N_37299,N_36137,N_36470);
xor U37300 (N_37300,N_36245,N_36015);
nor U37301 (N_37301,N_36119,N_36373);
nand U37302 (N_37302,N_36391,N_36629);
nand U37303 (N_37303,N_36927,N_36236);
and U37304 (N_37304,N_36659,N_36501);
nand U37305 (N_37305,N_36216,N_36427);
or U37306 (N_37306,N_36160,N_36933);
or U37307 (N_37307,N_36024,N_36291);
nor U37308 (N_37308,N_36891,N_36798);
nand U37309 (N_37309,N_36914,N_36176);
and U37310 (N_37310,N_36710,N_36222);
or U37311 (N_37311,N_36073,N_36821);
and U37312 (N_37312,N_36863,N_36354);
and U37313 (N_37313,N_36413,N_36545);
and U37314 (N_37314,N_36775,N_36235);
or U37315 (N_37315,N_36058,N_36495);
or U37316 (N_37316,N_36794,N_36695);
nor U37317 (N_37317,N_36652,N_36274);
and U37318 (N_37318,N_36924,N_36788);
or U37319 (N_37319,N_36603,N_36287);
and U37320 (N_37320,N_36458,N_36628);
or U37321 (N_37321,N_36084,N_36932);
and U37322 (N_37322,N_36920,N_36785);
nor U37323 (N_37323,N_36270,N_36790);
or U37324 (N_37324,N_36089,N_36580);
nand U37325 (N_37325,N_36797,N_36574);
xnor U37326 (N_37326,N_36828,N_36845);
xor U37327 (N_37327,N_36185,N_36825);
and U37328 (N_37328,N_36823,N_36591);
or U37329 (N_37329,N_36682,N_36170);
xor U37330 (N_37330,N_36452,N_36707);
or U37331 (N_37331,N_36332,N_36103);
nand U37332 (N_37332,N_36408,N_36852);
nand U37333 (N_37333,N_36673,N_36558);
or U37334 (N_37334,N_36397,N_36006);
nand U37335 (N_37335,N_36197,N_36731);
xor U37336 (N_37336,N_36900,N_36412);
and U37337 (N_37337,N_36065,N_36976);
xnor U37338 (N_37338,N_36892,N_36689);
xnor U37339 (N_37339,N_36761,N_36226);
nand U37340 (N_37340,N_36068,N_36946);
xor U37341 (N_37341,N_36277,N_36858);
nor U37342 (N_37342,N_36662,N_36525);
or U37343 (N_37343,N_36449,N_36768);
or U37344 (N_37344,N_36621,N_36271);
or U37345 (N_37345,N_36568,N_36953);
nor U37346 (N_37346,N_36200,N_36679);
and U37347 (N_37347,N_36688,N_36921);
nor U37348 (N_37348,N_36361,N_36998);
nand U37349 (N_37349,N_36395,N_36770);
and U37350 (N_37350,N_36779,N_36676);
nand U37351 (N_37351,N_36584,N_36241);
xor U37352 (N_37352,N_36299,N_36581);
nor U37353 (N_37353,N_36104,N_36763);
nor U37354 (N_37354,N_36524,N_36533);
xor U37355 (N_37355,N_36009,N_36318);
or U37356 (N_37356,N_36211,N_36899);
xnor U37357 (N_37357,N_36746,N_36835);
nor U37358 (N_37358,N_36795,N_36565);
nand U37359 (N_37359,N_36637,N_36756);
and U37360 (N_37360,N_36671,N_36173);
and U37361 (N_37361,N_36515,N_36105);
xor U37362 (N_37362,N_36464,N_36541);
nor U37363 (N_37363,N_36372,N_36650);
nor U37364 (N_37364,N_36035,N_36722);
and U37365 (N_37365,N_36206,N_36736);
or U37366 (N_37366,N_36910,N_36414);
or U37367 (N_37367,N_36193,N_36249);
nor U37368 (N_37368,N_36906,N_36432);
nand U37369 (N_37369,N_36307,N_36593);
nor U37370 (N_37370,N_36772,N_36726);
nand U37371 (N_37371,N_36439,N_36218);
nand U37372 (N_37372,N_36850,N_36555);
nand U37373 (N_37373,N_36294,N_36934);
nor U37374 (N_37374,N_36926,N_36508);
nand U37375 (N_37375,N_36209,N_36904);
nor U37376 (N_37376,N_36161,N_36725);
or U37377 (N_37377,N_36108,N_36864);
and U37378 (N_37378,N_36353,N_36368);
and U37379 (N_37379,N_36426,N_36422);
or U37380 (N_37380,N_36158,N_36887);
nor U37381 (N_37381,N_36879,N_36435);
nand U37382 (N_37382,N_36457,N_36538);
nand U37383 (N_37383,N_36716,N_36626);
nor U37384 (N_37384,N_36813,N_36991);
nand U37385 (N_37385,N_36980,N_36678);
and U37386 (N_37386,N_36965,N_36995);
xnor U37387 (N_37387,N_36867,N_36327);
nand U37388 (N_37388,N_36049,N_36393);
and U37389 (N_37389,N_36142,N_36140);
nor U37390 (N_37390,N_36254,N_36204);
xnor U37391 (N_37391,N_36461,N_36195);
xor U37392 (N_37392,N_36446,N_36784);
or U37393 (N_37393,N_36777,N_36846);
or U37394 (N_37394,N_36061,N_36594);
and U37395 (N_37395,N_36296,N_36702);
and U37396 (N_37396,N_36069,N_36669);
and U37397 (N_37397,N_36960,N_36192);
nor U37398 (N_37398,N_36915,N_36957);
and U37399 (N_37399,N_36613,N_36340);
nand U37400 (N_37400,N_36357,N_36635);
nor U37401 (N_37401,N_36109,N_36250);
and U37402 (N_37402,N_36830,N_36502);
nor U37403 (N_37403,N_36360,N_36028);
and U37404 (N_37404,N_36337,N_36261);
nor U37405 (N_37405,N_36834,N_36325);
nor U37406 (N_37406,N_36977,N_36631);
nor U37407 (N_37407,N_36885,N_36595);
xnor U37408 (N_37408,N_36029,N_36969);
xnor U37409 (N_37409,N_36362,N_36793);
nor U37410 (N_37410,N_36528,N_36114);
xnor U37411 (N_37411,N_36144,N_36339);
nor U37412 (N_37412,N_36607,N_36011);
or U37413 (N_37413,N_36377,N_36205);
or U37414 (N_37414,N_36654,N_36300);
nand U37415 (N_37415,N_36097,N_36433);
or U37416 (N_37416,N_36046,N_36096);
nor U37417 (N_37417,N_36856,N_36165);
xnor U37418 (N_37418,N_36916,N_36017);
nor U37419 (N_37419,N_36385,N_36560);
nand U37420 (N_37420,N_36908,N_36625);
nor U37421 (N_37421,N_36455,N_36664);
and U37422 (N_37422,N_36077,N_36336);
nand U37423 (N_37423,N_36898,N_36532);
nand U37424 (N_37424,N_36585,N_36324);
nand U37425 (N_37425,N_36043,N_36787);
and U37426 (N_37426,N_36100,N_36454);
and U37427 (N_37427,N_36582,N_36857);
nor U37428 (N_37428,N_36997,N_36497);
nor U37429 (N_37429,N_36194,N_36265);
xnor U37430 (N_37430,N_36549,N_36219);
nor U37431 (N_37431,N_36573,N_36022);
or U37432 (N_37432,N_36468,N_36527);
or U37433 (N_37433,N_36188,N_36769);
and U37434 (N_37434,N_36684,N_36431);
nor U37435 (N_37435,N_36622,N_36292);
xnor U37436 (N_37436,N_36247,N_36264);
nand U37437 (N_37437,N_36940,N_36252);
and U37438 (N_37438,N_36120,N_36663);
xor U37439 (N_37439,N_36278,N_36047);
nand U37440 (N_37440,N_36178,N_36888);
nor U37441 (N_37441,N_36601,N_36923);
nand U37442 (N_37442,N_36051,N_36308);
xor U37443 (N_37443,N_36014,N_36512);
nor U37444 (N_37444,N_36323,N_36179);
nor U37445 (N_37445,N_36872,N_36548);
or U37446 (N_37446,N_36214,N_36837);
or U37447 (N_37447,N_36189,N_36064);
nand U37448 (N_37448,N_36383,N_36704);
xnor U37449 (N_37449,N_36293,N_36705);
nand U37450 (N_37450,N_36886,N_36099);
nand U37451 (N_37451,N_36187,N_36429);
xnor U37452 (N_37452,N_36841,N_36453);
and U37453 (N_37453,N_36685,N_36718);
or U37454 (N_37454,N_36310,N_36928);
nor U37455 (N_37455,N_36730,N_36440);
nand U37456 (N_37456,N_36615,N_36984);
nor U37457 (N_37457,N_36799,N_36163);
nor U37458 (N_37458,N_36740,N_36493);
or U37459 (N_37459,N_36290,N_36311);
or U37460 (N_37460,N_36873,N_36131);
or U37461 (N_37461,N_36816,N_36919);
nand U37462 (N_37462,N_36564,N_36107);
nor U37463 (N_37463,N_36677,N_36135);
or U37464 (N_37464,N_36941,N_36284);
or U37465 (N_37465,N_36514,N_36374);
or U37466 (N_37466,N_36590,N_36539);
xnor U37467 (N_37467,N_36805,N_36633);
nor U37468 (N_37468,N_36286,N_36225);
nor U37469 (N_37469,N_36074,N_36262);
or U37470 (N_37470,N_36328,N_36566);
nor U37471 (N_37471,N_36732,N_36275);
nor U37472 (N_37472,N_36018,N_36778);
or U37473 (N_37473,N_36713,N_36344);
xor U37474 (N_37474,N_36350,N_36164);
and U37475 (N_37475,N_36972,N_36606);
or U37476 (N_37476,N_36840,N_36019);
xor U37477 (N_37477,N_36330,N_36048);
nor U37478 (N_37478,N_36242,N_36257);
or U37479 (N_37479,N_36467,N_36668);
xor U37480 (N_37480,N_36483,N_36829);
xor U37481 (N_37481,N_36260,N_36031);
nor U37482 (N_37482,N_36930,N_36243);
nand U37483 (N_37483,N_36263,N_36499);
xor U37484 (N_37484,N_36234,N_36623);
nand U37485 (N_37485,N_36640,N_36893);
or U37486 (N_37486,N_36507,N_36425);
nor U37487 (N_37487,N_36861,N_36884);
nand U37488 (N_37488,N_36505,N_36115);
xor U37489 (N_37489,N_36600,N_36994);
nand U37490 (N_37490,N_36604,N_36334);
xnor U37491 (N_37491,N_36936,N_36020);
xnor U37492 (N_37492,N_36530,N_36534);
and U37493 (N_37493,N_36698,N_36463);
nand U37494 (N_37494,N_36853,N_36003);
or U37495 (N_37495,N_36757,N_36966);
nand U37496 (N_37496,N_36859,N_36060);
nand U37497 (N_37497,N_36088,N_36036);
xnor U37498 (N_37498,N_36836,N_36517);
nand U37499 (N_37499,N_36759,N_36072);
nor U37500 (N_37500,N_36068,N_36941);
nor U37501 (N_37501,N_36852,N_36424);
and U37502 (N_37502,N_36598,N_36810);
and U37503 (N_37503,N_36816,N_36238);
nand U37504 (N_37504,N_36340,N_36364);
nor U37505 (N_37505,N_36364,N_36412);
nand U37506 (N_37506,N_36173,N_36794);
nor U37507 (N_37507,N_36769,N_36237);
xor U37508 (N_37508,N_36864,N_36622);
nand U37509 (N_37509,N_36502,N_36733);
nor U37510 (N_37510,N_36135,N_36836);
xor U37511 (N_37511,N_36555,N_36713);
nor U37512 (N_37512,N_36856,N_36757);
nand U37513 (N_37513,N_36714,N_36397);
and U37514 (N_37514,N_36213,N_36640);
nor U37515 (N_37515,N_36315,N_36373);
and U37516 (N_37516,N_36739,N_36819);
nor U37517 (N_37517,N_36767,N_36092);
nor U37518 (N_37518,N_36481,N_36997);
nand U37519 (N_37519,N_36578,N_36612);
nor U37520 (N_37520,N_36054,N_36471);
nand U37521 (N_37521,N_36485,N_36376);
and U37522 (N_37522,N_36966,N_36140);
xor U37523 (N_37523,N_36204,N_36008);
nand U37524 (N_37524,N_36855,N_36575);
xnor U37525 (N_37525,N_36742,N_36159);
xnor U37526 (N_37526,N_36639,N_36065);
nand U37527 (N_37527,N_36471,N_36900);
nor U37528 (N_37528,N_36748,N_36732);
nor U37529 (N_37529,N_36468,N_36530);
xor U37530 (N_37530,N_36988,N_36036);
and U37531 (N_37531,N_36859,N_36340);
nor U37532 (N_37532,N_36186,N_36842);
xnor U37533 (N_37533,N_36220,N_36648);
xor U37534 (N_37534,N_36714,N_36049);
and U37535 (N_37535,N_36910,N_36804);
nand U37536 (N_37536,N_36238,N_36354);
or U37537 (N_37537,N_36618,N_36503);
nor U37538 (N_37538,N_36391,N_36890);
nand U37539 (N_37539,N_36027,N_36794);
nand U37540 (N_37540,N_36569,N_36928);
or U37541 (N_37541,N_36541,N_36485);
nand U37542 (N_37542,N_36154,N_36940);
nand U37543 (N_37543,N_36715,N_36392);
and U37544 (N_37544,N_36519,N_36407);
nand U37545 (N_37545,N_36780,N_36601);
or U37546 (N_37546,N_36041,N_36653);
and U37547 (N_37547,N_36635,N_36903);
nand U37548 (N_37548,N_36916,N_36048);
and U37549 (N_37549,N_36864,N_36012);
and U37550 (N_37550,N_36435,N_36282);
nor U37551 (N_37551,N_36591,N_36190);
xnor U37552 (N_37552,N_36867,N_36054);
or U37553 (N_37553,N_36579,N_36398);
nand U37554 (N_37554,N_36822,N_36572);
or U37555 (N_37555,N_36656,N_36394);
or U37556 (N_37556,N_36657,N_36585);
nor U37557 (N_37557,N_36458,N_36390);
nor U37558 (N_37558,N_36262,N_36461);
or U37559 (N_37559,N_36218,N_36235);
nand U37560 (N_37560,N_36810,N_36756);
and U37561 (N_37561,N_36321,N_36788);
and U37562 (N_37562,N_36523,N_36736);
nor U37563 (N_37563,N_36983,N_36832);
xnor U37564 (N_37564,N_36221,N_36467);
or U37565 (N_37565,N_36393,N_36208);
nor U37566 (N_37566,N_36218,N_36340);
or U37567 (N_37567,N_36435,N_36456);
nor U37568 (N_37568,N_36326,N_36067);
nand U37569 (N_37569,N_36144,N_36079);
or U37570 (N_37570,N_36752,N_36759);
nor U37571 (N_37571,N_36323,N_36407);
or U37572 (N_37572,N_36529,N_36159);
xnor U37573 (N_37573,N_36430,N_36290);
and U37574 (N_37574,N_36431,N_36499);
xnor U37575 (N_37575,N_36445,N_36307);
nor U37576 (N_37576,N_36988,N_36072);
or U37577 (N_37577,N_36415,N_36351);
or U37578 (N_37578,N_36045,N_36843);
nor U37579 (N_37579,N_36542,N_36760);
or U37580 (N_37580,N_36220,N_36076);
nor U37581 (N_37581,N_36752,N_36665);
and U37582 (N_37582,N_36906,N_36216);
xor U37583 (N_37583,N_36457,N_36603);
or U37584 (N_37584,N_36854,N_36824);
nand U37585 (N_37585,N_36143,N_36491);
and U37586 (N_37586,N_36207,N_36615);
and U37587 (N_37587,N_36789,N_36368);
or U37588 (N_37588,N_36934,N_36333);
nand U37589 (N_37589,N_36088,N_36602);
nor U37590 (N_37590,N_36958,N_36193);
xor U37591 (N_37591,N_36375,N_36415);
nand U37592 (N_37592,N_36888,N_36779);
nor U37593 (N_37593,N_36130,N_36915);
nand U37594 (N_37594,N_36382,N_36616);
xnor U37595 (N_37595,N_36513,N_36294);
nor U37596 (N_37596,N_36969,N_36882);
nor U37597 (N_37597,N_36204,N_36538);
nor U37598 (N_37598,N_36949,N_36242);
nor U37599 (N_37599,N_36556,N_36322);
nor U37600 (N_37600,N_36357,N_36551);
nor U37601 (N_37601,N_36781,N_36572);
xor U37602 (N_37602,N_36096,N_36603);
nor U37603 (N_37603,N_36135,N_36570);
nor U37604 (N_37604,N_36347,N_36576);
or U37605 (N_37605,N_36424,N_36001);
nor U37606 (N_37606,N_36073,N_36852);
xor U37607 (N_37607,N_36534,N_36452);
xnor U37608 (N_37608,N_36114,N_36134);
xor U37609 (N_37609,N_36821,N_36575);
xnor U37610 (N_37610,N_36069,N_36241);
and U37611 (N_37611,N_36746,N_36072);
nand U37612 (N_37612,N_36916,N_36176);
nor U37613 (N_37613,N_36545,N_36305);
nand U37614 (N_37614,N_36007,N_36880);
xnor U37615 (N_37615,N_36690,N_36046);
xnor U37616 (N_37616,N_36980,N_36116);
xor U37617 (N_37617,N_36594,N_36899);
nor U37618 (N_37618,N_36236,N_36380);
or U37619 (N_37619,N_36809,N_36241);
nor U37620 (N_37620,N_36018,N_36911);
nand U37621 (N_37621,N_36856,N_36397);
xnor U37622 (N_37622,N_36385,N_36725);
and U37623 (N_37623,N_36735,N_36953);
or U37624 (N_37624,N_36578,N_36559);
and U37625 (N_37625,N_36809,N_36567);
xor U37626 (N_37626,N_36117,N_36434);
nand U37627 (N_37627,N_36258,N_36897);
nand U37628 (N_37628,N_36552,N_36032);
nand U37629 (N_37629,N_36987,N_36028);
nor U37630 (N_37630,N_36118,N_36965);
nand U37631 (N_37631,N_36371,N_36572);
xnor U37632 (N_37632,N_36179,N_36926);
nor U37633 (N_37633,N_36427,N_36797);
and U37634 (N_37634,N_36477,N_36362);
and U37635 (N_37635,N_36904,N_36522);
nor U37636 (N_37636,N_36790,N_36201);
or U37637 (N_37637,N_36746,N_36811);
and U37638 (N_37638,N_36844,N_36944);
and U37639 (N_37639,N_36853,N_36259);
nand U37640 (N_37640,N_36828,N_36452);
or U37641 (N_37641,N_36813,N_36073);
xnor U37642 (N_37642,N_36840,N_36437);
or U37643 (N_37643,N_36052,N_36677);
or U37644 (N_37644,N_36869,N_36874);
or U37645 (N_37645,N_36154,N_36294);
xnor U37646 (N_37646,N_36514,N_36301);
nor U37647 (N_37647,N_36532,N_36383);
nor U37648 (N_37648,N_36811,N_36599);
nand U37649 (N_37649,N_36835,N_36392);
nor U37650 (N_37650,N_36294,N_36592);
nand U37651 (N_37651,N_36751,N_36264);
xnor U37652 (N_37652,N_36260,N_36524);
xnor U37653 (N_37653,N_36300,N_36026);
xnor U37654 (N_37654,N_36609,N_36404);
and U37655 (N_37655,N_36548,N_36992);
and U37656 (N_37656,N_36361,N_36183);
nand U37657 (N_37657,N_36158,N_36803);
nand U37658 (N_37658,N_36314,N_36131);
and U37659 (N_37659,N_36382,N_36669);
nor U37660 (N_37660,N_36130,N_36034);
nand U37661 (N_37661,N_36115,N_36401);
nor U37662 (N_37662,N_36294,N_36200);
nand U37663 (N_37663,N_36793,N_36337);
xor U37664 (N_37664,N_36594,N_36093);
xnor U37665 (N_37665,N_36935,N_36523);
nor U37666 (N_37666,N_36471,N_36159);
nor U37667 (N_37667,N_36495,N_36350);
nor U37668 (N_37668,N_36656,N_36269);
nand U37669 (N_37669,N_36387,N_36401);
xnor U37670 (N_37670,N_36387,N_36462);
xnor U37671 (N_37671,N_36430,N_36409);
nand U37672 (N_37672,N_36803,N_36889);
or U37673 (N_37673,N_36534,N_36627);
nand U37674 (N_37674,N_36569,N_36855);
and U37675 (N_37675,N_36472,N_36576);
or U37676 (N_37676,N_36621,N_36046);
or U37677 (N_37677,N_36142,N_36765);
xor U37678 (N_37678,N_36576,N_36492);
xor U37679 (N_37679,N_36216,N_36440);
nand U37680 (N_37680,N_36742,N_36244);
and U37681 (N_37681,N_36915,N_36657);
nor U37682 (N_37682,N_36196,N_36455);
nand U37683 (N_37683,N_36315,N_36876);
nand U37684 (N_37684,N_36870,N_36581);
or U37685 (N_37685,N_36471,N_36025);
nand U37686 (N_37686,N_36112,N_36846);
nor U37687 (N_37687,N_36209,N_36625);
xnor U37688 (N_37688,N_36323,N_36979);
or U37689 (N_37689,N_36641,N_36019);
xnor U37690 (N_37690,N_36514,N_36683);
or U37691 (N_37691,N_36185,N_36570);
xnor U37692 (N_37692,N_36986,N_36525);
nand U37693 (N_37693,N_36375,N_36003);
or U37694 (N_37694,N_36272,N_36770);
and U37695 (N_37695,N_36685,N_36049);
nor U37696 (N_37696,N_36817,N_36602);
and U37697 (N_37697,N_36601,N_36641);
nor U37698 (N_37698,N_36516,N_36254);
nand U37699 (N_37699,N_36120,N_36928);
nor U37700 (N_37700,N_36610,N_36290);
nor U37701 (N_37701,N_36873,N_36942);
and U37702 (N_37702,N_36115,N_36097);
xor U37703 (N_37703,N_36182,N_36689);
or U37704 (N_37704,N_36456,N_36116);
and U37705 (N_37705,N_36323,N_36401);
or U37706 (N_37706,N_36495,N_36132);
nor U37707 (N_37707,N_36187,N_36459);
and U37708 (N_37708,N_36780,N_36053);
xnor U37709 (N_37709,N_36959,N_36794);
or U37710 (N_37710,N_36514,N_36858);
or U37711 (N_37711,N_36737,N_36407);
xnor U37712 (N_37712,N_36312,N_36182);
or U37713 (N_37713,N_36905,N_36527);
xnor U37714 (N_37714,N_36581,N_36015);
nor U37715 (N_37715,N_36248,N_36497);
nand U37716 (N_37716,N_36963,N_36991);
or U37717 (N_37717,N_36566,N_36699);
xor U37718 (N_37718,N_36564,N_36416);
and U37719 (N_37719,N_36067,N_36261);
nand U37720 (N_37720,N_36568,N_36143);
or U37721 (N_37721,N_36048,N_36310);
nand U37722 (N_37722,N_36443,N_36719);
nor U37723 (N_37723,N_36008,N_36910);
nand U37724 (N_37724,N_36589,N_36632);
or U37725 (N_37725,N_36467,N_36264);
nor U37726 (N_37726,N_36164,N_36877);
xnor U37727 (N_37727,N_36111,N_36141);
nand U37728 (N_37728,N_36303,N_36292);
and U37729 (N_37729,N_36050,N_36725);
and U37730 (N_37730,N_36561,N_36538);
xnor U37731 (N_37731,N_36911,N_36145);
or U37732 (N_37732,N_36078,N_36613);
nand U37733 (N_37733,N_36293,N_36887);
xnor U37734 (N_37734,N_36599,N_36740);
or U37735 (N_37735,N_36212,N_36185);
or U37736 (N_37736,N_36713,N_36151);
and U37737 (N_37737,N_36168,N_36775);
nand U37738 (N_37738,N_36575,N_36425);
nand U37739 (N_37739,N_36777,N_36231);
nor U37740 (N_37740,N_36760,N_36991);
nor U37741 (N_37741,N_36672,N_36087);
nor U37742 (N_37742,N_36260,N_36634);
or U37743 (N_37743,N_36183,N_36415);
or U37744 (N_37744,N_36219,N_36597);
or U37745 (N_37745,N_36342,N_36883);
and U37746 (N_37746,N_36452,N_36039);
xor U37747 (N_37747,N_36102,N_36305);
nand U37748 (N_37748,N_36835,N_36085);
or U37749 (N_37749,N_36880,N_36712);
and U37750 (N_37750,N_36779,N_36964);
xnor U37751 (N_37751,N_36133,N_36958);
or U37752 (N_37752,N_36188,N_36197);
nor U37753 (N_37753,N_36938,N_36426);
and U37754 (N_37754,N_36680,N_36249);
and U37755 (N_37755,N_36886,N_36572);
xnor U37756 (N_37756,N_36857,N_36611);
nand U37757 (N_37757,N_36140,N_36439);
or U37758 (N_37758,N_36299,N_36432);
nor U37759 (N_37759,N_36998,N_36752);
and U37760 (N_37760,N_36001,N_36560);
nand U37761 (N_37761,N_36794,N_36396);
nand U37762 (N_37762,N_36372,N_36237);
xor U37763 (N_37763,N_36055,N_36973);
xnor U37764 (N_37764,N_36669,N_36426);
nand U37765 (N_37765,N_36699,N_36257);
xor U37766 (N_37766,N_36136,N_36935);
nand U37767 (N_37767,N_36145,N_36084);
xor U37768 (N_37768,N_36512,N_36265);
or U37769 (N_37769,N_36331,N_36343);
xor U37770 (N_37770,N_36370,N_36760);
and U37771 (N_37771,N_36066,N_36650);
xnor U37772 (N_37772,N_36587,N_36529);
xnor U37773 (N_37773,N_36430,N_36505);
nor U37774 (N_37774,N_36746,N_36297);
and U37775 (N_37775,N_36717,N_36172);
or U37776 (N_37776,N_36814,N_36401);
nor U37777 (N_37777,N_36165,N_36792);
nand U37778 (N_37778,N_36239,N_36654);
xor U37779 (N_37779,N_36723,N_36143);
or U37780 (N_37780,N_36964,N_36380);
nand U37781 (N_37781,N_36571,N_36850);
nor U37782 (N_37782,N_36482,N_36354);
or U37783 (N_37783,N_36189,N_36497);
nor U37784 (N_37784,N_36000,N_36816);
or U37785 (N_37785,N_36365,N_36056);
nand U37786 (N_37786,N_36533,N_36655);
nor U37787 (N_37787,N_36486,N_36509);
or U37788 (N_37788,N_36300,N_36952);
xor U37789 (N_37789,N_36815,N_36064);
nor U37790 (N_37790,N_36478,N_36563);
nor U37791 (N_37791,N_36812,N_36769);
xor U37792 (N_37792,N_36778,N_36455);
nand U37793 (N_37793,N_36042,N_36124);
and U37794 (N_37794,N_36514,N_36966);
or U37795 (N_37795,N_36819,N_36850);
nor U37796 (N_37796,N_36892,N_36273);
or U37797 (N_37797,N_36419,N_36902);
and U37798 (N_37798,N_36153,N_36449);
nand U37799 (N_37799,N_36042,N_36311);
or U37800 (N_37800,N_36863,N_36573);
or U37801 (N_37801,N_36429,N_36062);
and U37802 (N_37802,N_36171,N_36920);
or U37803 (N_37803,N_36692,N_36301);
nor U37804 (N_37804,N_36515,N_36115);
or U37805 (N_37805,N_36798,N_36412);
or U37806 (N_37806,N_36032,N_36419);
or U37807 (N_37807,N_36769,N_36155);
nor U37808 (N_37808,N_36888,N_36875);
xnor U37809 (N_37809,N_36951,N_36645);
or U37810 (N_37810,N_36616,N_36098);
or U37811 (N_37811,N_36155,N_36101);
or U37812 (N_37812,N_36650,N_36866);
xor U37813 (N_37813,N_36374,N_36079);
nor U37814 (N_37814,N_36617,N_36891);
or U37815 (N_37815,N_36546,N_36698);
nand U37816 (N_37816,N_36579,N_36234);
nor U37817 (N_37817,N_36907,N_36052);
nor U37818 (N_37818,N_36847,N_36092);
nand U37819 (N_37819,N_36505,N_36617);
nand U37820 (N_37820,N_36105,N_36564);
nand U37821 (N_37821,N_36684,N_36083);
nor U37822 (N_37822,N_36183,N_36138);
nor U37823 (N_37823,N_36749,N_36420);
nand U37824 (N_37824,N_36910,N_36871);
xnor U37825 (N_37825,N_36868,N_36986);
nor U37826 (N_37826,N_36647,N_36110);
or U37827 (N_37827,N_36343,N_36210);
nor U37828 (N_37828,N_36765,N_36835);
and U37829 (N_37829,N_36044,N_36085);
or U37830 (N_37830,N_36632,N_36693);
nand U37831 (N_37831,N_36172,N_36789);
xor U37832 (N_37832,N_36347,N_36352);
or U37833 (N_37833,N_36827,N_36571);
nand U37834 (N_37834,N_36462,N_36003);
or U37835 (N_37835,N_36273,N_36427);
or U37836 (N_37836,N_36619,N_36931);
and U37837 (N_37837,N_36998,N_36180);
or U37838 (N_37838,N_36352,N_36175);
nor U37839 (N_37839,N_36367,N_36536);
or U37840 (N_37840,N_36806,N_36102);
or U37841 (N_37841,N_36955,N_36373);
xor U37842 (N_37842,N_36228,N_36117);
xnor U37843 (N_37843,N_36432,N_36249);
or U37844 (N_37844,N_36598,N_36981);
nand U37845 (N_37845,N_36482,N_36700);
xor U37846 (N_37846,N_36131,N_36176);
nor U37847 (N_37847,N_36798,N_36091);
xnor U37848 (N_37848,N_36020,N_36485);
nand U37849 (N_37849,N_36775,N_36270);
or U37850 (N_37850,N_36041,N_36680);
xor U37851 (N_37851,N_36020,N_36851);
nand U37852 (N_37852,N_36794,N_36296);
nor U37853 (N_37853,N_36682,N_36109);
nor U37854 (N_37854,N_36748,N_36400);
and U37855 (N_37855,N_36601,N_36314);
xor U37856 (N_37856,N_36892,N_36087);
or U37857 (N_37857,N_36817,N_36970);
and U37858 (N_37858,N_36599,N_36490);
xor U37859 (N_37859,N_36881,N_36375);
and U37860 (N_37860,N_36209,N_36384);
nand U37861 (N_37861,N_36929,N_36435);
nor U37862 (N_37862,N_36319,N_36404);
nand U37863 (N_37863,N_36562,N_36475);
or U37864 (N_37864,N_36151,N_36317);
xor U37865 (N_37865,N_36518,N_36199);
or U37866 (N_37866,N_36903,N_36571);
nor U37867 (N_37867,N_36363,N_36954);
nor U37868 (N_37868,N_36175,N_36747);
and U37869 (N_37869,N_36001,N_36243);
xor U37870 (N_37870,N_36827,N_36165);
nand U37871 (N_37871,N_36881,N_36517);
nor U37872 (N_37872,N_36858,N_36325);
nand U37873 (N_37873,N_36006,N_36289);
nor U37874 (N_37874,N_36937,N_36790);
nand U37875 (N_37875,N_36168,N_36947);
or U37876 (N_37876,N_36270,N_36155);
nand U37877 (N_37877,N_36377,N_36416);
or U37878 (N_37878,N_36032,N_36526);
nor U37879 (N_37879,N_36784,N_36902);
nor U37880 (N_37880,N_36852,N_36151);
nand U37881 (N_37881,N_36075,N_36098);
xnor U37882 (N_37882,N_36119,N_36568);
and U37883 (N_37883,N_36844,N_36549);
nor U37884 (N_37884,N_36033,N_36754);
nor U37885 (N_37885,N_36629,N_36056);
nand U37886 (N_37886,N_36277,N_36881);
or U37887 (N_37887,N_36960,N_36141);
and U37888 (N_37888,N_36115,N_36299);
nor U37889 (N_37889,N_36776,N_36293);
and U37890 (N_37890,N_36047,N_36982);
and U37891 (N_37891,N_36703,N_36949);
and U37892 (N_37892,N_36592,N_36109);
nand U37893 (N_37893,N_36295,N_36976);
nor U37894 (N_37894,N_36511,N_36440);
and U37895 (N_37895,N_36783,N_36812);
and U37896 (N_37896,N_36629,N_36161);
xor U37897 (N_37897,N_36359,N_36234);
nand U37898 (N_37898,N_36670,N_36608);
nand U37899 (N_37899,N_36951,N_36477);
nand U37900 (N_37900,N_36741,N_36393);
nor U37901 (N_37901,N_36502,N_36625);
or U37902 (N_37902,N_36367,N_36472);
nand U37903 (N_37903,N_36577,N_36100);
xor U37904 (N_37904,N_36828,N_36860);
nand U37905 (N_37905,N_36134,N_36267);
nor U37906 (N_37906,N_36560,N_36016);
xor U37907 (N_37907,N_36143,N_36273);
and U37908 (N_37908,N_36389,N_36818);
or U37909 (N_37909,N_36007,N_36474);
xnor U37910 (N_37910,N_36389,N_36476);
and U37911 (N_37911,N_36209,N_36404);
and U37912 (N_37912,N_36614,N_36865);
nand U37913 (N_37913,N_36536,N_36760);
and U37914 (N_37914,N_36085,N_36588);
or U37915 (N_37915,N_36978,N_36921);
or U37916 (N_37916,N_36249,N_36384);
nand U37917 (N_37917,N_36580,N_36425);
or U37918 (N_37918,N_36482,N_36005);
and U37919 (N_37919,N_36878,N_36326);
or U37920 (N_37920,N_36276,N_36034);
and U37921 (N_37921,N_36482,N_36312);
and U37922 (N_37922,N_36492,N_36390);
nand U37923 (N_37923,N_36661,N_36028);
xor U37924 (N_37924,N_36786,N_36981);
and U37925 (N_37925,N_36421,N_36107);
nor U37926 (N_37926,N_36703,N_36144);
xnor U37927 (N_37927,N_36358,N_36349);
and U37928 (N_37928,N_36150,N_36381);
nor U37929 (N_37929,N_36221,N_36198);
nor U37930 (N_37930,N_36795,N_36599);
and U37931 (N_37931,N_36373,N_36060);
nand U37932 (N_37932,N_36504,N_36656);
xnor U37933 (N_37933,N_36824,N_36879);
nand U37934 (N_37934,N_36380,N_36918);
or U37935 (N_37935,N_36075,N_36535);
nand U37936 (N_37936,N_36331,N_36780);
or U37937 (N_37937,N_36146,N_36642);
nor U37938 (N_37938,N_36932,N_36839);
xor U37939 (N_37939,N_36336,N_36004);
nor U37940 (N_37940,N_36961,N_36421);
nor U37941 (N_37941,N_36029,N_36104);
xor U37942 (N_37942,N_36241,N_36526);
nor U37943 (N_37943,N_36251,N_36684);
nand U37944 (N_37944,N_36807,N_36067);
xor U37945 (N_37945,N_36712,N_36094);
or U37946 (N_37946,N_36283,N_36255);
nand U37947 (N_37947,N_36189,N_36668);
and U37948 (N_37948,N_36620,N_36975);
and U37949 (N_37949,N_36604,N_36537);
nand U37950 (N_37950,N_36950,N_36153);
nor U37951 (N_37951,N_36458,N_36574);
nand U37952 (N_37952,N_36218,N_36433);
or U37953 (N_37953,N_36993,N_36260);
nor U37954 (N_37954,N_36955,N_36816);
nor U37955 (N_37955,N_36105,N_36079);
nor U37956 (N_37956,N_36215,N_36674);
xor U37957 (N_37957,N_36315,N_36641);
xnor U37958 (N_37958,N_36235,N_36952);
nor U37959 (N_37959,N_36503,N_36039);
nor U37960 (N_37960,N_36289,N_36755);
and U37961 (N_37961,N_36334,N_36955);
nand U37962 (N_37962,N_36241,N_36144);
nand U37963 (N_37963,N_36310,N_36100);
and U37964 (N_37964,N_36269,N_36550);
xor U37965 (N_37965,N_36489,N_36937);
xor U37966 (N_37966,N_36282,N_36503);
xor U37967 (N_37967,N_36487,N_36452);
or U37968 (N_37968,N_36634,N_36052);
and U37969 (N_37969,N_36141,N_36893);
or U37970 (N_37970,N_36044,N_36061);
and U37971 (N_37971,N_36478,N_36322);
nor U37972 (N_37972,N_36760,N_36327);
nand U37973 (N_37973,N_36870,N_36140);
nor U37974 (N_37974,N_36066,N_36070);
nand U37975 (N_37975,N_36155,N_36627);
xor U37976 (N_37976,N_36875,N_36200);
nor U37977 (N_37977,N_36856,N_36530);
and U37978 (N_37978,N_36258,N_36331);
xor U37979 (N_37979,N_36269,N_36571);
and U37980 (N_37980,N_36851,N_36922);
nand U37981 (N_37981,N_36668,N_36108);
xnor U37982 (N_37982,N_36820,N_36777);
and U37983 (N_37983,N_36413,N_36353);
or U37984 (N_37984,N_36764,N_36196);
nand U37985 (N_37985,N_36931,N_36432);
xor U37986 (N_37986,N_36460,N_36345);
and U37987 (N_37987,N_36536,N_36928);
nor U37988 (N_37988,N_36882,N_36096);
xor U37989 (N_37989,N_36960,N_36522);
nor U37990 (N_37990,N_36795,N_36900);
and U37991 (N_37991,N_36043,N_36206);
nor U37992 (N_37992,N_36347,N_36593);
or U37993 (N_37993,N_36380,N_36571);
and U37994 (N_37994,N_36647,N_36877);
nand U37995 (N_37995,N_36295,N_36743);
nand U37996 (N_37996,N_36946,N_36839);
nand U37997 (N_37997,N_36540,N_36530);
or U37998 (N_37998,N_36377,N_36087);
nand U37999 (N_37999,N_36264,N_36276);
and U38000 (N_38000,N_37175,N_37934);
nor U38001 (N_38001,N_37673,N_37830);
nor U38002 (N_38002,N_37416,N_37567);
nand U38003 (N_38003,N_37014,N_37810);
and U38004 (N_38004,N_37256,N_37690);
or U38005 (N_38005,N_37277,N_37237);
xnor U38006 (N_38006,N_37676,N_37140);
xor U38007 (N_38007,N_37342,N_37825);
xnor U38008 (N_38008,N_37261,N_37247);
and U38009 (N_38009,N_37951,N_37086);
xor U38010 (N_38010,N_37976,N_37746);
nand U38011 (N_38011,N_37560,N_37414);
and U38012 (N_38012,N_37218,N_37472);
and U38013 (N_38013,N_37743,N_37204);
or U38014 (N_38014,N_37313,N_37084);
xor U38015 (N_38015,N_37519,N_37310);
nand U38016 (N_38016,N_37610,N_37868);
or U38017 (N_38017,N_37590,N_37853);
nor U38018 (N_38018,N_37052,N_37229);
nor U38019 (N_38019,N_37141,N_37019);
nor U38020 (N_38020,N_37377,N_37424);
nor U38021 (N_38021,N_37048,N_37007);
nor U38022 (N_38022,N_37902,N_37107);
nand U38023 (N_38023,N_37792,N_37079);
or U38024 (N_38024,N_37704,N_37628);
nor U38025 (N_38025,N_37153,N_37716);
nor U38026 (N_38026,N_37920,N_37136);
or U38027 (N_38027,N_37038,N_37465);
xor U38028 (N_38028,N_37003,N_37517);
and U38029 (N_38029,N_37219,N_37917);
nor U38030 (N_38030,N_37235,N_37845);
xor U38031 (N_38031,N_37466,N_37407);
nand U38032 (N_38032,N_37812,N_37334);
and U38033 (N_38033,N_37467,N_37447);
or U38034 (N_38034,N_37524,N_37448);
nand U38035 (N_38035,N_37764,N_37104);
and U38036 (N_38036,N_37809,N_37895);
nand U38037 (N_38037,N_37823,N_37374);
or U38038 (N_38038,N_37271,N_37436);
or U38039 (N_38039,N_37726,N_37609);
or U38040 (N_38040,N_37440,N_37657);
or U38041 (N_38041,N_37276,N_37139);
and U38042 (N_38042,N_37419,N_37514);
xor U38043 (N_38043,N_37523,N_37708);
and U38044 (N_38044,N_37512,N_37901);
and U38045 (N_38045,N_37026,N_37150);
xor U38046 (N_38046,N_37208,N_37011);
xor U38047 (N_38047,N_37930,N_37835);
nand U38048 (N_38048,N_37702,N_37837);
or U38049 (N_38049,N_37325,N_37827);
nand U38050 (N_38050,N_37185,N_37388);
or U38051 (N_38051,N_37586,N_37879);
xnor U38052 (N_38052,N_37263,N_37406);
or U38053 (N_38053,N_37127,N_37700);
and U38054 (N_38054,N_37497,N_37265);
nor U38055 (N_38055,N_37762,N_37987);
nor U38056 (N_38056,N_37995,N_37516);
or U38057 (N_38057,N_37329,N_37568);
nor U38058 (N_38058,N_37615,N_37710);
xnor U38059 (N_38059,N_37278,N_37577);
nand U38060 (N_38060,N_37439,N_37842);
or U38061 (N_38061,N_37890,N_37621);
nand U38062 (N_38062,N_37645,N_37705);
xnor U38063 (N_38063,N_37321,N_37148);
and U38064 (N_38064,N_37757,N_37077);
nor U38065 (N_38065,N_37967,N_37748);
or U38066 (N_38066,N_37573,N_37583);
xnor U38067 (N_38067,N_37551,N_37692);
nor U38068 (N_38068,N_37862,N_37683);
and U38069 (N_38069,N_37638,N_37396);
or U38070 (N_38070,N_37910,N_37399);
and U38071 (N_38071,N_37492,N_37822);
nor U38072 (N_38072,N_37380,N_37339);
or U38073 (N_38073,N_37163,N_37832);
and U38074 (N_38074,N_37703,N_37887);
nor U38075 (N_38075,N_37113,N_37786);
nor U38076 (N_38076,N_37979,N_37138);
nand U38077 (N_38077,N_37224,N_37859);
and U38078 (N_38078,N_37285,N_37670);
xnor U38079 (N_38079,N_37230,N_37949);
or U38080 (N_38080,N_37298,N_37427);
and U38081 (N_38081,N_37652,N_37595);
and U38082 (N_38082,N_37417,N_37999);
nor U38083 (N_38083,N_37206,N_37896);
nor U38084 (N_38084,N_37304,N_37533);
or U38085 (N_38085,N_37324,N_37565);
nor U38086 (N_38086,N_37120,N_37126);
xnor U38087 (N_38087,N_37563,N_37088);
or U38088 (N_38088,N_37787,N_37100);
or U38089 (N_38089,N_37337,N_37561);
xor U38090 (N_38090,N_37642,N_37661);
nor U38091 (N_38091,N_37927,N_37681);
or U38092 (N_38092,N_37182,N_37212);
nor U38093 (N_38093,N_37458,N_37689);
and U38094 (N_38094,N_37360,N_37446);
and U38095 (N_38095,N_37530,N_37991);
and U38096 (N_38096,N_37935,N_37784);
xnor U38097 (N_38097,N_37085,N_37198);
nand U38098 (N_38098,N_37782,N_37640);
and U38099 (N_38099,N_37831,N_37028);
and U38100 (N_38100,N_37114,N_37611);
xor U38101 (N_38101,N_37509,N_37596);
nor U38102 (N_38102,N_37623,N_37720);
xnor U38103 (N_38103,N_37555,N_37747);
and U38104 (N_38104,N_37082,N_37351);
or U38105 (N_38105,N_37286,N_37373);
nor U38106 (N_38106,N_37569,N_37103);
xor U38107 (N_38107,N_37147,N_37418);
and U38108 (N_38108,N_37860,N_37311);
or U38109 (N_38109,N_37744,N_37507);
and U38110 (N_38110,N_37105,N_37066);
nand U38111 (N_38111,N_37566,N_37149);
or U38112 (N_38112,N_37117,N_37618);
nand U38113 (N_38113,N_37391,N_37225);
nor U38114 (N_38114,N_37434,N_37207);
xor U38115 (N_38115,N_37384,N_37790);
nand U38116 (N_38116,N_37170,N_37005);
xor U38117 (N_38117,N_37733,N_37301);
nand U38118 (N_38118,N_37778,N_37932);
or U38119 (N_38119,N_37952,N_37101);
and U38120 (N_38120,N_37036,N_37588);
xor U38121 (N_38121,N_37711,N_37065);
xor U38122 (N_38122,N_37522,N_37080);
xnor U38123 (N_38123,N_37875,N_37682);
nor U38124 (N_38124,N_37480,N_37355);
or U38125 (N_38125,N_37428,N_37348);
or U38126 (N_38126,N_37366,N_37909);
or U38127 (N_38127,N_37030,N_37675);
or U38128 (N_38128,N_37582,N_37495);
xnor U38129 (N_38129,N_37940,N_37713);
nand U38130 (N_38130,N_37591,N_37023);
xnor U38131 (N_38131,N_37718,N_37272);
and U38132 (N_38132,N_37178,N_37798);
nor U38133 (N_38133,N_37693,N_37612);
xor U38134 (N_38134,N_37662,N_37193);
or U38135 (N_38135,N_37966,N_37258);
or U38136 (N_38136,N_37993,N_37972);
nand U38137 (N_38137,N_37487,N_37070);
and U38138 (N_38138,N_37404,N_37145);
xor U38139 (N_38139,N_37597,N_37505);
xor U38140 (N_38140,N_37449,N_37624);
nand U38141 (N_38141,N_37773,N_37367);
xor U38142 (N_38142,N_37903,N_37322);
xor U38143 (N_38143,N_37456,N_37699);
or U38144 (N_38144,N_37707,N_37259);
nand U38145 (N_38145,N_37075,N_37408);
xor U38146 (N_38146,N_37722,N_37071);
or U38147 (N_38147,N_37217,N_37287);
or U38148 (N_38148,N_37944,N_37946);
and U38149 (N_38149,N_37425,N_37041);
xnor U38150 (N_38150,N_37037,N_37254);
or U38151 (N_38151,N_37463,N_37980);
xnor U38152 (N_38152,N_37970,N_37984);
or U38153 (N_38153,N_37099,N_37280);
or U38154 (N_38154,N_37819,N_37841);
nand U38155 (N_38155,N_37081,N_37742);
or U38156 (N_38156,N_37755,N_37884);
nor U38157 (N_38157,N_37010,N_37251);
nand U38158 (N_38158,N_37055,N_37195);
xnor U38159 (N_38159,N_37098,N_37210);
nand U38160 (N_38160,N_37231,N_37326);
nand U38161 (N_38161,N_37132,N_37904);
or U38162 (N_38162,N_37167,N_37811);
nor U38163 (N_38163,N_37632,N_37988);
nand U38164 (N_38164,N_37110,N_37248);
or U38165 (N_38165,N_37594,N_37740);
and U38166 (N_38166,N_37386,N_37807);
or U38167 (N_38167,N_37460,N_37818);
and U38168 (N_38168,N_37154,N_37022);
and U38169 (N_38169,N_37122,N_37796);
nor U38170 (N_38170,N_37783,N_37959);
nor U38171 (N_38171,N_37851,N_37034);
or U38172 (N_38172,N_37655,N_37600);
xnor U38173 (N_38173,N_37571,N_37550);
xnor U38174 (N_38174,N_37196,N_37969);
and U38175 (N_38175,N_37027,N_37714);
or U38176 (N_38176,N_37482,N_37620);
nand U38177 (N_38177,N_37146,N_37330);
nor U38178 (N_38178,N_37474,N_37238);
and U38179 (N_38179,N_37634,N_37262);
nor U38180 (N_38180,N_37438,N_37341);
or U38181 (N_38181,N_37688,N_37605);
nor U38182 (N_38182,N_37989,N_37246);
nor U38183 (N_38183,N_37135,N_37494);
and U38184 (N_38184,N_37915,N_37299);
or U38185 (N_38185,N_37763,N_37158);
nor U38186 (N_38186,N_37776,N_37622);
nand U38187 (N_38187,N_37925,N_37157);
xnor U38188 (N_38188,N_37834,N_37270);
nand U38189 (N_38189,N_37788,N_37971);
nand U38190 (N_38190,N_37601,N_37012);
xnor U38191 (N_38191,N_37861,N_37385);
or U38192 (N_38192,N_37186,N_37671);
nor U38193 (N_38193,N_37958,N_37305);
or U38194 (N_38194,N_37712,N_37050);
xor U38195 (N_38195,N_37518,N_37177);
and U38196 (N_38196,N_37264,N_37358);
and U38197 (N_38197,N_37319,N_37227);
nand U38198 (N_38198,N_37585,N_37400);
or U38199 (N_38199,N_37803,N_37866);
xnor U38200 (N_38200,N_37111,N_37266);
and U38201 (N_38201,N_37442,N_37478);
nand U38202 (N_38202,N_37468,N_37602);
xnor U38203 (N_38203,N_37719,N_37527);
nor U38204 (N_38204,N_37043,N_37074);
nand U38205 (N_38205,N_37556,N_37473);
xnor U38206 (N_38206,N_37090,N_37947);
xnor U38207 (N_38207,N_37152,N_37357);
and U38208 (N_38208,N_37821,N_37284);
xnor U38209 (N_38209,N_37775,N_37869);
nand U38210 (N_38210,N_37816,N_37756);
nand U38211 (N_38211,N_37489,N_37189);
nand U38212 (N_38212,N_37665,N_37964);
and U38213 (N_38213,N_37617,N_37891);
or U38214 (N_38214,N_37996,N_37797);
nand U38215 (N_38215,N_37997,N_37540);
xnor U38216 (N_38216,N_37333,N_37736);
nand U38217 (N_38217,N_37922,N_37794);
nor U38218 (N_38218,N_37354,N_37921);
and U38219 (N_38219,N_37916,N_37059);
xor U38220 (N_38220,N_37883,N_37525);
and U38221 (N_38221,N_37572,N_37490);
nor U38222 (N_38222,N_37799,N_37124);
or U38223 (N_38223,N_37768,N_37128);
and U38224 (N_38224,N_37031,N_37244);
and U38225 (N_38225,N_37877,N_37240);
nor U38226 (N_38226,N_37429,N_37986);
nor U38227 (N_38227,N_37724,N_37476);
and U38228 (N_38228,N_37926,N_37411);
and U38229 (N_38229,N_37129,N_37183);
nand U38230 (N_38230,N_37598,N_37936);
nand U38231 (N_38231,N_37592,N_37331);
nand U38232 (N_38232,N_37637,N_37394);
xor U38233 (N_38233,N_37619,N_37302);
and U38234 (N_38234,N_37562,N_37542);
xor U38235 (N_38235,N_37123,N_37089);
nand U38236 (N_38236,N_37653,N_37888);
or U38237 (N_38237,N_37644,N_37593);
nor U38238 (N_38238,N_37546,N_37452);
nor U38239 (N_38239,N_37194,N_37253);
nor U38240 (N_38240,N_37353,N_37804);
or U38241 (N_38241,N_37759,N_37445);
or U38242 (N_38242,N_37214,N_37937);
or U38243 (N_38243,N_37426,N_37006);
or U38244 (N_38244,N_37383,N_37882);
nor U38245 (N_38245,N_37905,N_37291);
nor U38246 (N_38246,N_37197,N_37772);
xor U38247 (N_38247,N_37667,N_37076);
and U38248 (N_38248,N_37729,N_37543);
nand U38249 (N_38249,N_37273,N_37053);
nor U38250 (N_38250,N_37228,N_37062);
or U38251 (N_38251,N_37444,N_37063);
nor U38252 (N_38252,N_37282,N_37633);
or U38253 (N_38253,N_37395,N_37625);
or U38254 (N_38254,N_37886,N_37754);
and U38255 (N_38255,N_37791,N_37042);
xor U38256 (N_38256,N_37933,N_37045);
nor U38257 (N_38257,N_37636,N_37504);
nor U38258 (N_38258,N_37728,N_37420);
or U38259 (N_38259,N_37359,N_37626);
nand U38260 (N_38260,N_37865,N_37697);
nand U38261 (N_38261,N_37013,N_37630);
nand U38262 (N_38262,N_37343,N_37470);
xnor U38263 (N_38263,N_37381,N_37368);
nand U38264 (N_38264,N_37498,N_37469);
and U38265 (N_38265,N_37893,N_37180);
nand U38266 (N_38266,N_37092,N_37908);
and U38267 (N_38267,N_37002,N_37269);
or U38268 (N_38268,N_37375,N_37168);
and U38269 (N_38269,N_37846,N_37701);
nor U38270 (N_38270,N_37222,N_37867);
nand U38271 (N_38271,N_37898,N_37421);
nor U38272 (N_38272,N_37441,N_37142);
nor U38273 (N_38273,N_37205,N_37938);
nand U38274 (N_38274,N_37379,N_37535);
or U38275 (N_38275,N_37695,N_37292);
nor U38276 (N_38276,N_37233,N_37457);
or U38277 (N_38277,N_37900,N_37164);
or U38278 (N_38278,N_37973,N_37674);
nor U38279 (N_38279,N_37760,N_37627);
xor U38280 (N_38280,N_37844,N_37249);
or U38281 (N_38281,N_37017,N_37962);
xor U38282 (N_38282,N_37328,N_37169);
and U38283 (N_38283,N_37496,N_37539);
nor U38284 (N_38284,N_37309,N_37532);
nand U38285 (N_38285,N_37361,N_37923);
and U38286 (N_38286,N_37639,N_37047);
nor U38287 (N_38287,N_37200,N_37994);
and U38288 (N_38288,N_37554,N_37491);
nor U38289 (N_38289,N_37802,N_37793);
xnor U38290 (N_38290,N_37020,N_37838);
xnor U38291 (N_38291,N_37172,N_37409);
nor U38292 (N_38292,N_37215,N_37046);
nor U38293 (N_38293,N_37643,N_37192);
nand U38294 (N_38294,N_37413,N_37369);
or U38295 (N_38295,N_37850,N_37159);
nand U38296 (N_38296,N_37173,N_37477);
nand U38297 (N_38297,N_37236,N_37267);
nor U38298 (N_38298,N_37390,N_37151);
and U38299 (N_38299,N_37314,N_37412);
or U38300 (N_38300,N_37464,N_37067);
nand U38301 (N_38301,N_37134,N_37558);
nand U38302 (N_38302,N_37912,N_37795);
and U38303 (N_38303,N_37599,N_37587);
or U38304 (N_38304,N_37387,N_37503);
or U38305 (N_38305,N_37430,N_37422);
xnor U38306 (N_38306,N_37025,N_37370);
or U38307 (N_38307,N_37108,N_37488);
nor U38308 (N_38308,N_37907,N_37534);
nor U38309 (N_38309,N_37771,N_37574);
xor U38310 (N_38310,N_37453,N_37181);
and U38311 (N_38311,N_37484,N_37928);
or U38312 (N_38312,N_37161,N_37654);
or U38313 (N_38313,N_37435,N_37696);
xnor U38314 (N_38314,N_37650,N_37858);
xor U38315 (N_38315,N_37064,N_37345);
and U38316 (N_38316,N_37808,N_37401);
nor U38317 (N_38317,N_37631,N_37761);
nand U38318 (N_38318,N_37320,N_37854);
or U38319 (N_38319,N_37843,N_37433);
or U38320 (N_38320,N_37415,N_37255);
nor U38321 (N_38321,N_37190,N_37855);
or U38322 (N_38322,N_37275,N_37589);
and U38323 (N_38323,N_37929,N_37758);
nor U38324 (N_38324,N_37506,N_37260);
and U38325 (N_38325,N_37723,N_37243);
nor U38326 (N_38326,N_37226,N_37752);
or U38327 (N_38327,N_37829,N_37068);
xor U38328 (N_38328,N_37656,N_37093);
and U38329 (N_38329,N_37981,N_37953);
nor U38330 (N_38330,N_37564,N_37647);
or U38331 (N_38331,N_37083,N_37091);
nor U38332 (N_38332,N_37578,N_37857);
nand U38333 (N_38333,N_37500,N_37770);
xor U38334 (N_38334,N_37116,N_37061);
and U38335 (N_38335,N_37750,N_37162);
xnor U38336 (N_38336,N_37242,N_37058);
xnor U38337 (N_38337,N_37317,N_37559);
xnor U38338 (N_38338,N_37166,N_37057);
and U38339 (N_38339,N_37398,N_37121);
or U38340 (N_38340,N_37983,N_37443);
and U38341 (N_38341,N_37666,N_37717);
nand U38342 (N_38342,N_37044,N_37919);
and U38343 (N_38343,N_37118,N_37283);
or U38344 (N_38344,N_37942,N_37307);
nor U38345 (N_38345,N_37137,N_37731);
nor U38346 (N_38346,N_37423,N_37350);
xnor U38347 (N_38347,N_37687,N_37774);
xnor U38348 (N_38348,N_37364,N_37245);
or U38349 (N_38349,N_37096,N_37016);
nand U38350 (N_38350,N_37727,N_37336);
nor U38351 (N_38351,N_37913,N_37018);
or U38352 (N_38352,N_37863,N_37035);
xor U38353 (N_38353,N_37015,N_37450);
xnor U38354 (N_38354,N_37475,N_37279);
or U38355 (N_38355,N_37847,N_37538);
and U38356 (N_38356,N_37709,N_37806);
nor U38357 (N_38357,N_37779,N_37741);
nor U38358 (N_38358,N_37725,N_37739);
nor U38359 (N_38359,N_37363,N_37347);
nor U38360 (N_38360,N_37635,N_37471);
nand U38361 (N_38361,N_37213,N_37570);
nand U38362 (N_38362,N_37651,N_37906);
nand U38363 (N_38363,N_37000,N_37069);
nand U38364 (N_38364,N_37848,N_37106);
or U38365 (N_38365,N_37780,N_37397);
and U38366 (N_38366,N_37029,N_37056);
xor U38367 (N_38367,N_37785,N_37294);
nor U38368 (N_38368,N_37978,N_37297);
xnor U38369 (N_38369,N_37977,N_37998);
nand U38370 (N_38370,N_37557,N_37968);
xor U38371 (N_38371,N_37584,N_37871);
xnor U38372 (N_38372,N_37992,N_37371);
or U38373 (N_38373,N_37548,N_37293);
nand U38374 (N_38374,N_37160,N_37165);
nor U38375 (N_38375,N_37828,N_37965);
and U38376 (N_38376,N_37221,N_37686);
and U38377 (N_38377,N_37914,N_37608);
and U38378 (N_38378,N_37125,N_37308);
and U38379 (N_38379,N_37939,N_37544);
nor U38380 (N_38380,N_37840,N_37982);
or U38381 (N_38381,N_37143,N_37179);
and U38382 (N_38382,N_37049,N_37604);
and U38383 (N_38383,N_37281,N_37894);
and U38384 (N_38384,N_37493,N_37257);
nand U38385 (N_38385,N_37545,N_37032);
and U38386 (N_38386,N_37873,N_37340);
nand U38387 (N_38387,N_37431,N_37672);
nand U38388 (N_38388,N_37072,N_37510);
and U38389 (N_38389,N_37541,N_37737);
and U38390 (N_38390,N_37112,N_37303);
and U38391 (N_38391,N_37751,N_37392);
and U38392 (N_38392,N_37814,N_37677);
or U38393 (N_38393,N_37833,N_37800);
nand U38394 (N_38394,N_37389,N_37187);
xor U38395 (N_38395,N_37664,N_37201);
nand U38396 (N_38396,N_37511,N_37203);
or U38397 (N_38397,N_37911,N_37691);
or U38398 (N_38398,N_37306,N_37008);
nand U38399 (N_38399,N_37580,N_37462);
xnor U38400 (N_38400,N_37629,N_37529);
xor U38401 (N_38401,N_37892,N_37033);
nor U38402 (N_38402,N_37176,N_37119);
xor U38403 (N_38403,N_37356,N_37730);
xor U38404 (N_38404,N_37735,N_37191);
nand U38405 (N_38405,N_37547,N_37437);
or U38406 (N_38406,N_37216,N_37531);
nand U38407 (N_38407,N_37852,N_37753);
xor U38408 (N_38408,N_37715,N_37985);
and U38409 (N_38409,N_37549,N_37094);
xnor U38410 (N_38410,N_37223,N_37232);
nand U38411 (N_38411,N_37576,N_37499);
and U38412 (N_38412,N_37826,N_37220);
and U38413 (N_38413,N_37312,N_37553);
nand U38414 (N_38414,N_37694,N_37024);
or U38415 (N_38415,N_37955,N_37721);
nand U38416 (N_38416,N_37880,N_37402);
nor U38417 (N_38417,N_37945,N_37526);
nand U38418 (N_38418,N_37870,N_37485);
nand U38419 (N_38419,N_37289,N_37963);
nand U38420 (N_38420,N_37209,N_37581);
nor U38421 (N_38421,N_37184,N_37943);
nor U38422 (N_38422,N_37732,N_37767);
or U38423 (N_38423,N_37250,N_37552);
nand U38424 (N_38424,N_37097,N_37338);
and U38425 (N_38425,N_37648,N_37606);
or U38426 (N_38426,N_37521,N_37766);
nor U38427 (N_38427,N_37410,N_37528);
nor U38428 (N_38428,N_37820,N_37603);
nor U38429 (N_38429,N_37815,N_37155);
xor U38430 (N_38430,N_37508,N_37614);
xnor U38431 (N_38431,N_37513,N_37789);
nand U38432 (N_38432,N_37961,N_37613);
and U38433 (N_38433,N_37975,N_37885);
or U38434 (N_38434,N_37813,N_37461);
and U38435 (N_38435,N_37171,N_37899);
nor U38436 (N_38436,N_37706,N_37749);
nand U38437 (N_38437,N_37459,N_37202);
nor U38438 (N_38438,N_37144,N_37483);
nor U38439 (N_38439,N_37575,N_37376);
and U38440 (N_38440,N_37781,N_37054);
and U38441 (N_38441,N_37365,N_37102);
nor U38442 (N_38442,N_37188,N_37346);
or U38443 (N_38443,N_37801,N_37393);
and U38444 (N_38444,N_37156,N_37537);
and U38445 (N_38445,N_37405,N_37646);
nor U38446 (N_38446,N_37641,N_37290);
xor U38447 (N_38447,N_37680,N_37878);
nor U38448 (N_38448,N_37199,N_37864);
and U38449 (N_38449,N_37021,N_37769);
xnor U38450 (N_38450,N_37805,N_37889);
and U38451 (N_38451,N_37960,N_37954);
xor U38452 (N_38452,N_37268,N_37332);
and U38453 (N_38453,N_37536,N_37607);
nand U38454 (N_38454,N_37004,N_37300);
xnor U38455 (N_38455,N_37481,N_37378);
xnor U38456 (N_38456,N_37502,N_37455);
and U38457 (N_38457,N_37130,N_37349);
nor U38458 (N_38458,N_37881,N_37001);
nand U38459 (N_38459,N_37679,N_37352);
or U38460 (N_38460,N_37990,N_37372);
nor U38461 (N_38461,N_37234,N_37872);
nor U38462 (N_38462,N_37659,N_37288);
and U38463 (N_38463,N_37344,N_37515);
xor U38464 (N_38464,N_37941,N_37362);
xnor U38465 (N_38465,N_37403,N_37318);
nand U38466 (N_38466,N_37974,N_37296);
nor U38467 (N_38467,N_37078,N_37658);
and U38468 (N_38468,N_37432,N_37874);
xnor U38469 (N_38469,N_37738,N_37087);
xor U38470 (N_38470,N_37073,N_37252);
or U38471 (N_38471,N_37131,N_37824);
or U38472 (N_38472,N_37734,N_37060);
or U38473 (N_38473,N_37836,N_37817);
or U38474 (N_38474,N_37924,N_37323);
xor U38475 (N_38475,N_37663,N_37479);
and U38476 (N_38476,N_37876,N_37950);
or U38477 (N_38477,N_37316,N_37486);
and U38478 (N_38478,N_37918,N_37382);
and U38479 (N_38479,N_37295,N_37095);
xor U38480 (N_38480,N_37451,N_37241);
or U38481 (N_38481,N_37931,N_37698);
xor U38482 (N_38482,N_37133,N_37649);
nand U38483 (N_38483,N_37327,N_37579);
nand U38484 (N_38484,N_37040,N_37174);
and U38485 (N_38485,N_37109,N_37115);
nor U38486 (N_38486,N_37660,N_37051);
or U38487 (N_38487,N_37520,N_37777);
nand U38488 (N_38488,N_37956,N_37501);
nand U38489 (N_38489,N_37315,N_37849);
nor U38490 (N_38490,N_37669,N_37856);
nor U38491 (N_38491,N_37335,N_37684);
and U38492 (N_38492,N_37009,N_37274);
or U38493 (N_38493,N_37239,N_37765);
nor U38494 (N_38494,N_37211,N_37616);
nor U38495 (N_38495,N_37668,N_37678);
and U38496 (N_38496,N_37039,N_37957);
nand U38497 (N_38497,N_37685,N_37839);
and U38498 (N_38498,N_37948,N_37897);
nor U38499 (N_38499,N_37745,N_37454);
or U38500 (N_38500,N_37700,N_37155);
nand U38501 (N_38501,N_37830,N_37739);
xnor U38502 (N_38502,N_37123,N_37040);
nor U38503 (N_38503,N_37828,N_37387);
nand U38504 (N_38504,N_37811,N_37841);
or U38505 (N_38505,N_37115,N_37452);
nand U38506 (N_38506,N_37003,N_37375);
or U38507 (N_38507,N_37175,N_37229);
xor U38508 (N_38508,N_37264,N_37519);
and U38509 (N_38509,N_37196,N_37813);
or U38510 (N_38510,N_37968,N_37625);
xnor U38511 (N_38511,N_37042,N_37790);
or U38512 (N_38512,N_37613,N_37967);
xor U38513 (N_38513,N_37167,N_37383);
nand U38514 (N_38514,N_37422,N_37989);
or U38515 (N_38515,N_37408,N_37238);
nand U38516 (N_38516,N_37085,N_37925);
or U38517 (N_38517,N_37766,N_37504);
and U38518 (N_38518,N_37715,N_37898);
xnor U38519 (N_38519,N_37175,N_37482);
or U38520 (N_38520,N_37083,N_37611);
or U38521 (N_38521,N_37948,N_37394);
or U38522 (N_38522,N_37118,N_37889);
nor U38523 (N_38523,N_37404,N_37325);
nor U38524 (N_38524,N_37436,N_37506);
nand U38525 (N_38525,N_37535,N_37273);
or U38526 (N_38526,N_37673,N_37861);
nand U38527 (N_38527,N_37334,N_37919);
nand U38528 (N_38528,N_37101,N_37586);
nor U38529 (N_38529,N_37396,N_37157);
nor U38530 (N_38530,N_37282,N_37623);
nand U38531 (N_38531,N_37561,N_37550);
and U38532 (N_38532,N_37297,N_37739);
and U38533 (N_38533,N_37517,N_37388);
or U38534 (N_38534,N_37378,N_37707);
and U38535 (N_38535,N_37816,N_37376);
xor U38536 (N_38536,N_37148,N_37437);
nor U38537 (N_38537,N_37349,N_37937);
or U38538 (N_38538,N_37033,N_37324);
nor U38539 (N_38539,N_37836,N_37970);
xnor U38540 (N_38540,N_37007,N_37498);
and U38541 (N_38541,N_37538,N_37975);
or U38542 (N_38542,N_37332,N_37009);
or U38543 (N_38543,N_37180,N_37087);
xor U38544 (N_38544,N_37548,N_37902);
xor U38545 (N_38545,N_37357,N_37996);
nor U38546 (N_38546,N_37394,N_37275);
nor U38547 (N_38547,N_37783,N_37671);
or U38548 (N_38548,N_37071,N_37767);
xnor U38549 (N_38549,N_37671,N_37855);
and U38550 (N_38550,N_37032,N_37930);
and U38551 (N_38551,N_37373,N_37497);
nor U38552 (N_38552,N_37632,N_37668);
nand U38553 (N_38553,N_37011,N_37862);
xnor U38554 (N_38554,N_37714,N_37127);
nand U38555 (N_38555,N_37347,N_37737);
xor U38556 (N_38556,N_37811,N_37882);
or U38557 (N_38557,N_37495,N_37931);
and U38558 (N_38558,N_37759,N_37288);
or U38559 (N_38559,N_37865,N_37220);
xnor U38560 (N_38560,N_37527,N_37011);
nand U38561 (N_38561,N_37536,N_37798);
or U38562 (N_38562,N_37445,N_37226);
nand U38563 (N_38563,N_37307,N_37455);
nor U38564 (N_38564,N_37492,N_37554);
nand U38565 (N_38565,N_37247,N_37357);
nor U38566 (N_38566,N_37404,N_37410);
nor U38567 (N_38567,N_37298,N_37980);
nand U38568 (N_38568,N_37796,N_37143);
xor U38569 (N_38569,N_37238,N_37696);
xor U38570 (N_38570,N_37295,N_37980);
or U38571 (N_38571,N_37274,N_37074);
xnor U38572 (N_38572,N_37561,N_37125);
nand U38573 (N_38573,N_37215,N_37781);
nor U38574 (N_38574,N_37866,N_37359);
nor U38575 (N_38575,N_37577,N_37023);
xnor U38576 (N_38576,N_37042,N_37131);
xnor U38577 (N_38577,N_37347,N_37742);
xor U38578 (N_38578,N_37435,N_37667);
or U38579 (N_38579,N_37159,N_37967);
nand U38580 (N_38580,N_37130,N_37565);
nor U38581 (N_38581,N_37823,N_37810);
xnor U38582 (N_38582,N_37931,N_37130);
or U38583 (N_38583,N_37339,N_37746);
or U38584 (N_38584,N_37407,N_37000);
xor U38585 (N_38585,N_37015,N_37742);
and U38586 (N_38586,N_37241,N_37143);
nand U38587 (N_38587,N_37357,N_37264);
nor U38588 (N_38588,N_37301,N_37408);
nor U38589 (N_38589,N_37313,N_37570);
and U38590 (N_38590,N_37175,N_37542);
xnor U38591 (N_38591,N_37923,N_37271);
xor U38592 (N_38592,N_37980,N_37852);
and U38593 (N_38593,N_37710,N_37382);
or U38594 (N_38594,N_37755,N_37810);
nand U38595 (N_38595,N_37263,N_37139);
and U38596 (N_38596,N_37666,N_37245);
or U38597 (N_38597,N_37552,N_37026);
or U38598 (N_38598,N_37420,N_37114);
nand U38599 (N_38599,N_37768,N_37466);
xnor U38600 (N_38600,N_37896,N_37014);
nand U38601 (N_38601,N_37078,N_37720);
xnor U38602 (N_38602,N_37129,N_37416);
and U38603 (N_38603,N_37300,N_37297);
nand U38604 (N_38604,N_37193,N_37828);
nor U38605 (N_38605,N_37537,N_37311);
nand U38606 (N_38606,N_37572,N_37964);
nor U38607 (N_38607,N_37479,N_37350);
or U38608 (N_38608,N_37207,N_37843);
and U38609 (N_38609,N_37585,N_37988);
and U38610 (N_38610,N_37455,N_37733);
or U38611 (N_38611,N_37225,N_37883);
xor U38612 (N_38612,N_37857,N_37411);
and U38613 (N_38613,N_37102,N_37142);
xor U38614 (N_38614,N_37098,N_37875);
and U38615 (N_38615,N_37345,N_37808);
xor U38616 (N_38616,N_37528,N_37919);
nand U38617 (N_38617,N_37950,N_37525);
or U38618 (N_38618,N_37016,N_37729);
nand U38619 (N_38619,N_37750,N_37586);
xor U38620 (N_38620,N_37858,N_37694);
nor U38621 (N_38621,N_37572,N_37760);
nor U38622 (N_38622,N_37279,N_37673);
and U38623 (N_38623,N_37285,N_37483);
or U38624 (N_38624,N_37033,N_37874);
and U38625 (N_38625,N_37162,N_37920);
nand U38626 (N_38626,N_37855,N_37375);
nor U38627 (N_38627,N_37436,N_37418);
and U38628 (N_38628,N_37871,N_37615);
nor U38629 (N_38629,N_37362,N_37810);
nand U38630 (N_38630,N_37100,N_37419);
xnor U38631 (N_38631,N_37598,N_37640);
nand U38632 (N_38632,N_37390,N_37101);
or U38633 (N_38633,N_37369,N_37078);
xor U38634 (N_38634,N_37948,N_37719);
or U38635 (N_38635,N_37125,N_37437);
and U38636 (N_38636,N_37329,N_37192);
and U38637 (N_38637,N_37366,N_37332);
or U38638 (N_38638,N_37270,N_37390);
and U38639 (N_38639,N_37102,N_37407);
xor U38640 (N_38640,N_37423,N_37094);
and U38641 (N_38641,N_37350,N_37965);
nand U38642 (N_38642,N_37662,N_37849);
xnor U38643 (N_38643,N_37334,N_37885);
xor U38644 (N_38644,N_37645,N_37943);
or U38645 (N_38645,N_37469,N_37791);
nand U38646 (N_38646,N_37123,N_37884);
nor U38647 (N_38647,N_37003,N_37042);
xor U38648 (N_38648,N_37395,N_37382);
nand U38649 (N_38649,N_37799,N_37985);
nor U38650 (N_38650,N_37294,N_37417);
xnor U38651 (N_38651,N_37362,N_37586);
nor U38652 (N_38652,N_37428,N_37018);
nand U38653 (N_38653,N_37677,N_37093);
xor U38654 (N_38654,N_37496,N_37108);
and U38655 (N_38655,N_37280,N_37002);
and U38656 (N_38656,N_37605,N_37091);
or U38657 (N_38657,N_37273,N_37635);
nor U38658 (N_38658,N_37653,N_37974);
xnor U38659 (N_38659,N_37300,N_37191);
nand U38660 (N_38660,N_37936,N_37295);
xnor U38661 (N_38661,N_37614,N_37721);
and U38662 (N_38662,N_37117,N_37622);
and U38663 (N_38663,N_37549,N_37502);
nand U38664 (N_38664,N_37584,N_37223);
and U38665 (N_38665,N_37944,N_37467);
and U38666 (N_38666,N_37064,N_37231);
nand U38667 (N_38667,N_37629,N_37170);
xnor U38668 (N_38668,N_37138,N_37693);
nor U38669 (N_38669,N_37808,N_37557);
or U38670 (N_38670,N_37337,N_37242);
or U38671 (N_38671,N_37033,N_37273);
and U38672 (N_38672,N_37934,N_37675);
xnor U38673 (N_38673,N_37838,N_37990);
nor U38674 (N_38674,N_37159,N_37306);
or U38675 (N_38675,N_37758,N_37761);
or U38676 (N_38676,N_37017,N_37216);
or U38677 (N_38677,N_37174,N_37151);
and U38678 (N_38678,N_37626,N_37408);
nor U38679 (N_38679,N_37597,N_37660);
xor U38680 (N_38680,N_37105,N_37503);
nor U38681 (N_38681,N_37162,N_37009);
nor U38682 (N_38682,N_37998,N_37820);
or U38683 (N_38683,N_37993,N_37151);
nand U38684 (N_38684,N_37480,N_37541);
nor U38685 (N_38685,N_37795,N_37398);
or U38686 (N_38686,N_37616,N_37519);
and U38687 (N_38687,N_37858,N_37752);
nor U38688 (N_38688,N_37892,N_37019);
xnor U38689 (N_38689,N_37393,N_37882);
nand U38690 (N_38690,N_37411,N_37045);
and U38691 (N_38691,N_37912,N_37955);
xnor U38692 (N_38692,N_37221,N_37243);
nand U38693 (N_38693,N_37321,N_37227);
xnor U38694 (N_38694,N_37920,N_37352);
or U38695 (N_38695,N_37836,N_37042);
nand U38696 (N_38696,N_37265,N_37404);
xnor U38697 (N_38697,N_37508,N_37171);
and U38698 (N_38698,N_37861,N_37988);
or U38699 (N_38699,N_37730,N_37547);
xor U38700 (N_38700,N_37068,N_37041);
nand U38701 (N_38701,N_37988,N_37959);
xnor U38702 (N_38702,N_37109,N_37531);
nor U38703 (N_38703,N_37351,N_37597);
nand U38704 (N_38704,N_37974,N_37324);
or U38705 (N_38705,N_37272,N_37411);
or U38706 (N_38706,N_37352,N_37831);
nand U38707 (N_38707,N_37933,N_37635);
xor U38708 (N_38708,N_37298,N_37086);
xnor U38709 (N_38709,N_37965,N_37161);
or U38710 (N_38710,N_37474,N_37473);
or U38711 (N_38711,N_37044,N_37991);
nor U38712 (N_38712,N_37350,N_37477);
xor U38713 (N_38713,N_37108,N_37072);
nor U38714 (N_38714,N_37625,N_37386);
and U38715 (N_38715,N_37574,N_37176);
and U38716 (N_38716,N_37156,N_37803);
or U38717 (N_38717,N_37552,N_37960);
nor U38718 (N_38718,N_37028,N_37891);
nor U38719 (N_38719,N_37549,N_37067);
xor U38720 (N_38720,N_37283,N_37566);
nor U38721 (N_38721,N_37775,N_37705);
and U38722 (N_38722,N_37342,N_37783);
and U38723 (N_38723,N_37914,N_37068);
or U38724 (N_38724,N_37712,N_37440);
or U38725 (N_38725,N_37174,N_37141);
or U38726 (N_38726,N_37212,N_37113);
or U38727 (N_38727,N_37643,N_37843);
nor U38728 (N_38728,N_37543,N_37485);
or U38729 (N_38729,N_37298,N_37275);
nand U38730 (N_38730,N_37947,N_37887);
nand U38731 (N_38731,N_37556,N_37431);
or U38732 (N_38732,N_37770,N_37478);
xnor U38733 (N_38733,N_37420,N_37121);
xnor U38734 (N_38734,N_37822,N_37595);
and U38735 (N_38735,N_37830,N_37334);
xnor U38736 (N_38736,N_37381,N_37994);
or U38737 (N_38737,N_37667,N_37161);
xnor U38738 (N_38738,N_37363,N_37532);
and U38739 (N_38739,N_37162,N_37769);
and U38740 (N_38740,N_37829,N_37378);
nor U38741 (N_38741,N_37518,N_37883);
nand U38742 (N_38742,N_37361,N_37186);
nor U38743 (N_38743,N_37486,N_37958);
nand U38744 (N_38744,N_37765,N_37084);
or U38745 (N_38745,N_37377,N_37509);
xor U38746 (N_38746,N_37844,N_37927);
nand U38747 (N_38747,N_37992,N_37251);
nand U38748 (N_38748,N_37544,N_37057);
nand U38749 (N_38749,N_37375,N_37761);
or U38750 (N_38750,N_37423,N_37084);
nand U38751 (N_38751,N_37048,N_37329);
or U38752 (N_38752,N_37175,N_37426);
xnor U38753 (N_38753,N_37049,N_37726);
xor U38754 (N_38754,N_37566,N_37804);
or U38755 (N_38755,N_37343,N_37854);
or U38756 (N_38756,N_37175,N_37686);
nor U38757 (N_38757,N_37851,N_37919);
xnor U38758 (N_38758,N_37556,N_37194);
nand U38759 (N_38759,N_37231,N_37137);
and U38760 (N_38760,N_37945,N_37861);
nand U38761 (N_38761,N_37295,N_37131);
nand U38762 (N_38762,N_37002,N_37409);
nor U38763 (N_38763,N_37986,N_37864);
xor U38764 (N_38764,N_37154,N_37798);
nand U38765 (N_38765,N_37814,N_37149);
xor U38766 (N_38766,N_37236,N_37081);
nand U38767 (N_38767,N_37255,N_37925);
or U38768 (N_38768,N_37256,N_37627);
and U38769 (N_38769,N_37451,N_37108);
and U38770 (N_38770,N_37366,N_37259);
nand U38771 (N_38771,N_37353,N_37764);
nand U38772 (N_38772,N_37023,N_37598);
or U38773 (N_38773,N_37580,N_37093);
or U38774 (N_38774,N_37738,N_37246);
xnor U38775 (N_38775,N_37544,N_37255);
or U38776 (N_38776,N_37853,N_37896);
xor U38777 (N_38777,N_37047,N_37104);
xnor U38778 (N_38778,N_37435,N_37544);
nand U38779 (N_38779,N_37496,N_37162);
and U38780 (N_38780,N_37728,N_37354);
nor U38781 (N_38781,N_37563,N_37790);
nand U38782 (N_38782,N_37436,N_37447);
and U38783 (N_38783,N_37032,N_37007);
nand U38784 (N_38784,N_37256,N_37839);
nand U38785 (N_38785,N_37784,N_37662);
xor U38786 (N_38786,N_37359,N_37192);
nand U38787 (N_38787,N_37551,N_37250);
nand U38788 (N_38788,N_37769,N_37920);
nor U38789 (N_38789,N_37112,N_37658);
nor U38790 (N_38790,N_37709,N_37657);
nand U38791 (N_38791,N_37427,N_37043);
and U38792 (N_38792,N_37473,N_37993);
and U38793 (N_38793,N_37954,N_37393);
xnor U38794 (N_38794,N_37933,N_37451);
nor U38795 (N_38795,N_37033,N_37565);
or U38796 (N_38796,N_37793,N_37978);
nor U38797 (N_38797,N_37873,N_37016);
nor U38798 (N_38798,N_37750,N_37492);
or U38799 (N_38799,N_37049,N_37641);
xor U38800 (N_38800,N_37844,N_37846);
nor U38801 (N_38801,N_37398,N_37122);
or U38802 (N_38802,N_37822,N_37040);
nand U38803 (N_38803,N_37831,N_37662);
nand U38804 (N_38804,N_37910,N_37161);
or U38805 (N_38805,N_37649,N_37926);
nor U38806 (N_38806,N_37194,N_37520);
and U38807 (N_38807,N_37903,N_37026);
nor U38808 (N_38808,N_37750,N_37817);
xor U38809 (N_38809,N_37529,N_37076);
and U38810 (N_38810,N_37608,N_37463);
or U38811 (N_38811,N_37854,N_37229);
nor U38812 (N_38812,N_37964,N_37766);
or U38813 (N_38813,N_37447,N_37784);
nand U38814 (N_38814,N_37104,N_37448);
or U38815 (N_38815,N_37313,N_37669);
and U38816 (N_38816,N_37157,N_37223);
and U38817 (N_38817,N_37284,N_37314);
or U38818 (N_38818,N_37309,N_37695);
xor U38819 (N_38819,N_37636,N_37888);
or U38820 (N_38820,N_37574,N_37184);
or U38821 (N_38821,N_37201,N_37304);
and U38822 (N_38822,N_37069,N_37622);
nand U38823 (N_38823,N_37469,N_37553);
or U38824 (N_38824,N_37769,N_37899);
xnor U38825 (N_38825,N_37212,N_37917);
or U38826 (N_38826,N_37142,N_37003);
nand U38827 (N_38827,N_37646,N_37075);
xor U38828 (N_38828,N_37128,N_37637);
nor U38829 (N_38829,N_37506,N_37881);
xor U38830 (N_38830,N_37856,N_37602);
nand U38831 (N_38831,N_37063,N_37719);
and U38832 (N_38832,N_37818,N_37313);
or U38833 (N_38833,N_37654,N_37646);
or U38834 (N_38834,N_37591,N_37957);
nand U38835 (N_38835,N_37315,N_37995);
nand U38836 (N_38836,N_37613,N_37421);
nor U38837 (N_38837,N_37122,N_37446);
or U38838 (N_38838,N_37861,N_37526);
or U38839 (N_38839,N_37621,N_37880);
and U38840 (N_38840,N_37348,N_37863);
or U38841 (N_38841,N_37137,N_37196);
or U38842 (N_38842,N_37651,N_37745);
or U38843 (N_38843,N_37186,N_37289);
or U38844 (N_38844,N_37661,N_37496);
nand U38845 (N_38845,N_37979,N_37788);
xnor U38846 (N_38846,N_37475,N_37282);
nor U38847 (N_38847,N_37166,N_37566);
and U38848 (N_38848,N_37488,N_37507);
xnor U38849 (N_38849,N_37142,N_37996);
nand U38850 (N_38850,N_37514,N_37660);
nand U38851 (N_38851,N_37315,N_37109);
nand U38852 (N_38852,N_37643,N_37402);
or U38853 (N_38853,N_37238,N_37992);
nor U38854 (N_38854,N_37899,N_37392);
or U38855 (N_38855,N_37843,N_37758);
nor U38856 (N_38856,N_37529,N_37591);
or U38857 (N_38857,N_37231,N_37579);
or U38858 (N_38858,N_37024,N_37122);
xnor U38859 (N_38859,N_37939,N_37563);
or U38860 (N_38860,N_37165,N_37410);
or U38861 (N_38861,N_37826,N_37412);
and U38862 (N_38862,N_37071,N_37299);
nor U38863 (N_38863,N_37765,N_37412);
nor U38864 (N_38864,N_37038,N_37694);
nor U38865 (N_38865,N_37490,N_37602);
or U38866 (N_38866,N_37885,N_37301);
and U38867 (N_38867,N_37428,N_37655);
nand U38868 (N_38868,N_37114,N_37056);
and U38869 (N_38869,N_37007,N_37294);
and U38870 (N_38870,N_37489,N_37949);
nand U38871 (N_38871,N_37781,N_37013);
or U38872 (N_38872,N_37247,N_37974);
and U38873 (N_38873,N_37151,N_37695);
and U38874 (N_38874,N_37420,N_37597);
or U38875 (N_38875,N_37620,N_37778);
xor U38876 (N_38876,N_37583,N_37932);
xnor U38877 (N_38877,N_37991,N_37671);
and U38878 (N_38878,N_37489,N_37999);
xor U38879 (N_38879,N_37421,N_37251);
nand U38880 (N_38880,N_37560,N_37520);
xnor U38881 (N_38881,N_37440,N_37678);
or U38882 (N_38882,N_37896,N_37587);
nor U38883 (N_38883,N_37956,N_37147);
nand U38884 (N_38884,N_37929,N_37500);
nand U38885 (N_38885,N_37932,N_37371);
xnor U38886 (N_38886,N_37781,N_37391);
or U38887 (N_38887,N_37611,N_37038);
nand U38888 (N_38888,N_37017,N_37746);
or U38889 (N_38889,N_37069,N_37230);
nor U38890 (N_38890,N_37701,N_37507);
xor U38891 (N_38891,N_37205,N_37269);
nand U38892 (N_38892,N_37649,N_37827);
nor U38893 (N_38893,N_37410,N_37809);
and U38894 (N_38894,N_37823,N_37041);
nand U38895 (N_38895,N_37531,N_37999);
nor U38896 (N_38896,N_37454,N_37116);
and U38897 (N_38897,N_37332,N_37990);
xnor U38898 (N_38898,N_37953,N_37819);
nand U38899 (N_38899,N_37349,N_37528);
nand U38900 (N_38900,N_37159,N_37920);
and U38901 (N_38901,N_37020,N_37116);
or U38902 (N_38902,N_37602,N_37615);
and U38903 (N_38903,N_37116,N_37815);
or U38904 (N_38904,N_37975,N_37442);
and U38905 (N_38905,N_37850,N_37191);
nand U38906 (N_38906,N_37165,N_37710);
or U38907 (N_38907,N_37801,N_37432);
and U38908 (N_38908,N_37517,N_37847);
or U38909 (N_38909,N_37794,N_37210);
and U38910 (N_38910,N_37995,N_37501);
nor U38911 (N_38911,N_37721,N_37963);
nor U38912 (N_38912,N_37266,N_37374);
and U38913 (N_38913,N_37655,N_37773);
and U38914 (N_38914,N_37388,N_37821);
nor U38915 (N_38915,N_37377,N_37555);
or U38916 (N_38916,N_37284,N_37665);
xor U38917 (N_38917,N_37883,N_37164);
and U38918 (N_38918,N_37083,N_37277);
nand U38919 (N_38919,N_37190,N_37873);
nor U38920 (N_38920,N_37320,N_37024);
or U38921 (N_38921,N_37483,N_37695);
nor U38922 (N_38922,N_37771,N_37913);
xor U38923 (N_38923,N_37356,N_37195);
and U38924 (N_38924,N_37518,N_37224);
xor U38925 (N_38925,N_37374,N_37241);
nor U38926 (N_38926,N_37191,N_37760);
or U38927 (N_38927,N_37554,N_37906);
or U38928 (N_38928,N_37050,N_37791);
nor U38929 (N_38929,N_37929,N_37689);
nor U38930 (N_38930,N_37833,N_37477);
nor U38931 (N_38931,N_37815,N_37919);
and U38932 (N_38932,N_37428,N_37633);
or U38933 (N_38933,N_37485,N_37448);
nand U38934 (N_38934,N_37856,N_37378);
nand U38935 (N_38935,N_37123,N_37896);
and U38936 (N_38936,N_37792,N_37885);
and U38937 (N_38937,N_37867,N_37020);
xnor U38938 (N_38938,N_37198,N_37204);
and U38939 (N_38939,N_37893,N_37389);
xor U38940 (N_38940,N_37041,N_37858);
nor U38941 (N_38941,N_37025,N_37179);
and U38942 (N_38942,N_37649,N_37444);
or U38943 (N_38943,N_37587,N_37559);
nor U38944 (N_38944,N_37407,N_37606);
nor U38945 (N_38945,N_37212,N_37816);
nor U38946 (N_38946,N_37177,N_37818);
xnor U38947 (N_38947,N_37107,N_37699);
nand U38948 (N_38948,N_37453,N_37002);
xnor U38949 (N_38949,N_37742,N_37194);
nor U38950 (N_38950,N_37189,N_37944);
and U38951 (N_38951,N_37158,N_37271);
nand U38952 (N_38952,N_37504,N_37391);
nand U38953 (N_38953,N_37148,N_37133);
or U38954 (N_38954,N_37478,N_37203);
and U38955 (N_38955,N_37816,N_37179);
xnor U38956 (N_38956,N_37659,N_37863);
xnor U38957 (N_38957,N_37517,N_37443);
nand U38958 (N_38958,N_37693,N_37066);
nand U38959 (N_38959,N_37106,N_37215);
nand U38960 (N_38960,N_37530,N_37345);
xor U38961 (N_38961,N_37243,N_37701);
and U38962 (N_38962,N_37875,N_37483);
nor U38963 (N_38963,N_37879,N_37600);
nor U38964 (N_38964,N_37543,N_37892);
or U38965 (N_38965,N_37078,N_37745);
nand U38966 (N_38966,N_37855,N_37902);
and U38967 (N_38967,N_37428,N_37317);
nor U38968 (N_38968,N_37905,N_37606);
or U38969 (N_38969,N_37538,N_37174);
or U38970 (N_38970,N_37606,N_37496);
nand U38971 (N_38971,N_37081,N_37701);
nor U38972 (N_38972,N_37339,N_37349);
nand U38973 (N_38973,N_37098,N_37943);
and U38974 (N_38974,N_37480,N_37110);
and U38975 (N_38975,N_37831,N_37664);
xor U38976 (N_38976,N_37275,N_37541);
nand U38977 (N_38977,N_37442,N_37272);
nand U38978 (N_38978,N_37994,N_37886);
nand U38979 (N_38979,N_37085,N_37535);
and U38980 (N_38980,N_37502,N_37377);
xor U38981 (N_38981,N_37891,N_37670);
nor U38982 (N_38982,N_37117,N_37508);
or U38983 (N_38983,N_37869,N_37759);
nor U38984 (N_38984,N_37325,N_37677);
nor U38985 (N_38985,N_37883,N_37952);
and U38986 (N_38986,N_37693,N_37624);
nor U38987 (N_38987,N_37420,N_37991);
or U38988 (N_38988,N_37238,N_37865);
xnor U38989 (N_38989,N_37069,N_37180);
nor U38990 (N_38990,N_37612,N_37492);
nor U38991 (N_38991,N_37371,N_37043);
or U38992 (N_38992,N_37597,N_37703);
nand U38993 (N_38993,N_37419,N_37812);
and U38994 (N_38994,N_37765,N_37839);
nor U38995 (N_38995,N_37274,N_37712);
and U38996 (N_38996,N_37607,N_37994);
nor U38997 (N_38997,N_37948,N_37347);
and U38998 (N_38998,N_37221,N_37753);
nand U38999 (N_38999,N_37693,N_37982);
and U39000 (N_39000,N_38446,N_38881);
or U39001 (N_39001,N_38338,N_38123);
or U39002 (N_39002,N_38328,N_38288);
xor U39003 (N_39003,N_38139,N_38188);
and U39004 (N_39004,N_38841,N_38267);
and U39005 (N_39005,N_38804,N_38047);
and U39006 (N_39006,N_38237,N_38284);
xnor U39007 (N_39007,N_38579,N_38443);
xnor U39008 (N_39008,N_38825,N_38894);
nor U39009 (N_39009,N_38052,N_38718);
or U39010 (N_39010,N_38072,N_38993);
and U39011 (N_39011,N_38913,N_38137);
xnor U39012 (N_39012,N_38790,N_38964);
or U39013 (N_39013,N_38191,N_38310);
xnor U39014 (N_39014,N_38619,N_38426);
nor U39015 (N_39015,N_38061,N_38669);
or U39016 (N_39016,N_38253,N_38104);
or U39017 (N_39017,N_38933,N_38610);
or U39018 (N_39018,N_38517,N_38982);
and U39019 (N_39019,N_38956,N_38975);
and U39020 (N_39020,N_38043,N_38932);
xor U39021 (N_39021,N_38403,N_38616);
nor U39022 (N_39022,N_38304,N_38623);
nand U39023 (N_39023,N_38361,N_38357);
xor U39024 (N_39024,N_38375,N_38388);
nor U39025 (N_39025,N_38127,N_38971);
or U39026 (N_39026,N_38301,N_38534);
xnor U39027 (N_39027,N_38822,N_38834);
nor U39028 (N_39028,N_38800,N_38942);
or U39029 (N_39029,N_38447,N_38053);
and U39030 (N_39030,N_38210,N_38686);
nand U39031 (N_39031,N_38467,N_38239);
nand U39032 (N_39032,N_38489,N_38738);
xor U39033 (N_39033,N_38185,N_38297);
nor U39034 (N_39034,N_38787,N_38866);
nand U39035 (N_39035,N_38694,N_38549);
nor U39036 (N_39036,N_38335,N_38133);
nor U39037 (N_39037,N_38990,N_38638);
or U39038 (N_39038,N_38348,N_38459);
and U39039 (N_39039,N_38656,N_38373);
and U39040 (N_39040,N_38140,N_38155);
or U39041 (N_39041,N_38519,N_38176);
nand U39042 (N_39042,N_38878,N_38224);
nand U39043 (N_39043,N_38949,N_38608);
nand U39044 (N_39044,N_38076,N_38154);
or U39045 (N_39045,N_38423,N_38776);
or U39046 (N_39046,N_38536,N_38037);
nor U39047 (N_39047,N_38462,N_38548);
nand U39048 (N_39048,N_38230,N_38797);
and U39049 (N_39049,N_38920,N_38455);
or U39050 (N_39050,N_38680,N_38495);
xor U39051 (N_39051,N_38416,N_38067);
nand U39052 (N_39052,N_38028,N_38818);
and U39053 (N_39053,N_38095,N_38892);
and U39054 (N_39054,N_38336,N_38522);
xnor U39055 (N_39055,N_38978,N_38504);
and U39056 (N_39056,N_38621,N_38066);
xnor U39057 (N_39057,N_38168,N_38796);
nor U39058 (N_39058,N_38477,N_38624);
xor U39059 (N_39059,N_38196,N_38440);
nor U39060 (N_39060,N_38511,N_38194);
nand U39061 (N_39061,N_38986,N_38592);
nand U39062 (N_39062,N_38677,N_38442);
xnor U39063 (N_39063,N_38547,N_38100);
nor U39064 (N_39064,N_38500,N_38236);
nand U39065 (N_39065,N_38001,N_38174);
xor U39066 (N_39066,N_38998,N_38885);
and U39067 (N_39067,N_38668,N_38480);
or U39068 (N_39068,N_38979,N_38458);
or U39069 (N_39069,N_38420,N_38409);
nor U39070 (N_39070,N_38889,N_38231);
and U39071 (N_39071,N_38510,N_38456);
nand U39072 (N_39072,N_38503,N_38018);
nor U39073 (N_39073,N_38858,N_38255);
xor U39074 (N_39074,N_38419,N_38676);
nor U39075 (N_39075,N_38745,N_38784);
nand U39076 (N_39076,N_38523,N_38882);
or U39077 (N_39077,N_38763,N_38890);
xor U39078 (N_39078,N_38131,N_38098);
nor U39079 (N_39079,N_38537,N_38678);
nor U39080 (N_39080,N_38159,N_38068);
and U39081 (N_39081,N_38853,N_38380);
nand U39082 (N_39082,N_38259,N_38460);
nor U39083 (N_39083,N_38204,N_38090);
xor U39084 (N_39084,N_38976,N_38472);
nor U39085 (N_39085,N_38699,N_38124);
nor U39086 (N_39086,N_38454,N_38600);
nor U39087 (N_39087,N_38767,N_38539);
nor U39088 (N_39088,N_38257,N_38554);
nand U39089 (N_39089,N_38362,N_38349);
nand U39090 (N_39090,N_38739,N_38967);
or U39091 (N_39091,N_38648,N_38735);
or U39092 (N_39092,N_38609,N_38201);
xnor U39093 (N_39093,N_38852,N_38049);
and U39094 (N_39094,N_38453,N_38112);
nor U39095 (N_39095,N_38856,N_38938);
and U39096 (N_39096,N_38206,N_38937);
nand U39097 (N_39097,N_38376,N_38078);
xnor U39098 (N_39098,N_38602,N_38966);
xnor U39099 (N_39099,N_38642,N_38958);
and U39100 (N_39100,N_38783,N_38629);
nand U39101 (N_39101,N_38202,N_38050);
nor U39102 (N_39102,N_38550,N_38146);
nand U39103 (N_39103,N_38567,N_38228);
nor U39104 (N_39104,N_38870,N_38292);
nand U39105 (N_39105,N_38606,N_38717);
or U39106 (N_39106,N_38598,N_38492);
xor U39107 (N_39107,N_38665,N_38116);
nor U39108 (N_39108,N_38120,N_38184);
or U39109 (N_39109,N_38593,N_38973);
nor U39110 (N_39110,N_38021,N_38528);
xnor U39111 (N_39111,N_38189,N_38631);
nand U39112 (N_39112,N_38992,N_38172);
and U39113 (N_39113,N_38351,N_38160);
nor U39114 (N_39114,N_38479,N_38344);
and U39115 (N_39115,N_38429,N_38746);
and U39116 (N_39116,N_38162,N_38461);
and U39117 (N_39117,N_38003,N_38529);
nand U39118 (N_39118,N_38101,N_38035);
nand U39119 (N_39119,N_38064,N_38716);
and U39120 (N_39120,N_38538,N_38166);
and U39121 (N_39121,N_38723,N_38122);
or U39122 (N_39122,N_38947,N_38983);
xor U39123 (N_39123,N_38241,N_38082);
xnor U39124 (N_39124,N_38173,N_38293);
and U39125 (N_39125,N_38180,N_38708);
nand U39126 (N_39126,N_38125,N_38675);
nor U39127 (N_39127,N_38182,N_38613);
nor U39128 (N_39128,N_38353,N_38381);
nor U39129 (N_39129,N_38531,N_38828);
nand U39130 (N_39130,N_38209,N_38859);
nor U39131 (N_39131,N_38910,N_38187);
or U39132 (N_39132,N_38806,N_38483);
xor U39133 (N_39133,N_38099,N_38208);
nor U39134 (N_39134,N_38412,N_38743);
or U39135 (N_39135,N_38315,N_38662);
xor U39136 (N_39136,N_38004,N_38908);
and U39137 (N_39137,N_38792,N_38791);
or U39138 (N_39138,N_38476,N_38584);
and U39139 (N_39139,N_38896,N_38056);
nand U39140 (N_39140,N_38482,N_38406);
xor U39141 (N_39141,N_38617,N_38603);
and U39142 (N_39142,N_38860,N_38425);
nor U39143 (N_39143,N_38802,N_38060);
and U39144 (N_39144,N_38200,N_38820);
nor U39145 (N_39145,N_38436,N_38089);
nand U39146 (N_39146,N_38091,N_38058);
xor U39147 (N_39147,N_38046,N_38749);
or U39148 (N_39148,N_38935,N_38965);
nand U39149 (N_39149,N_38901,N_38904);
xor U39150 (N_39150,N_38819,N_38632);
and U39151 (N_39151,N_38689,N_38566);
nand U39152 (N_39152,N_38306,N_38331);
and U39153 (N_39153,N_38260,N_38151);
nor U39154 (N_39154,N_38726,N_38955);
or U39155 (N_39155,N_38719,N_38438);
xor U39156 (N_39156,N_38198,N_38785);
and U39157 (N_39157,N_38474,N_38364);
nor U39158 (N_39158,N_38478,N_38303);
nand U39159 (N_39159,N_38830,N_38002);
nand U39160 (N_39160,N_38010,N_38452);
nand U39161 (N_39161,N_38917,N_38542);
nand U39162 (N_39162,N_38660,N_38217);
xnor U39163 (N_39163,N_38826,N_38300);
nor U39164 (N_39164,N_38240,N_38827);
xor U39165 (N_39165,N_38421,N_38494);
and U39166 (N_39166,N_38696,N_38595);
nand U39167 (N_39167,N_38999,N_38755);
or U39168 (N_39168,N_38295,N_38342);
nor U39169 (N_39169,N_38872,N_38134);
and U39170 (N_39170,N_38270,N_38063);
nand U39171 (N_39171,N_38291,N_38559);
nor U39172 (N_39172,N_38324,N_38836);
and U39173 (N_39173,N_38756,N_38765);
nand U39174 (N_39174,N_38874,N_38736);
nor U39175 (N_39175,N_38574,N_38778);
nor U39176 (N_39176,N_38527,N_38450);
nand U39177 (N_39177,N_38895,N_38957);
or U39178 (N_39178,N_38972,N_38524);
nand U39179 (N_39179,N_38130,N_38410);
xnor U39180 (N_39180,N_38661,N_38244);
xnor U39181 (N_39181,N_38813,N_38158);
nand U39182 (N_39182,N_38569,N_38245);
xnor U39183 (N_39183,N_38313,N_38088);
or U39184 (N_39184,N_38604,N_38664);
and U39185 (N_39185,N_38924,N_38633);
nand U39186 (N_39186,N_38948,N_38867);
nand U39187 (N_39187,N_38383,N_38902);
nor U39188 (N_39188,N_38857,N_38590);
nand U39189 (N_39189,N_38759,N_38488);
nor U39190 (N_39190,N_38484,N_38628);
nor U39191 (N_39191,N_38521,N_38687);
nor U39192 (N_39192,N_38691,N_38252);
nor U39193 (N_39193,N_38281,N_38946);
xnor U39194 (N_39194,N_38518,N_38312);
xnor U39195 (N_39195,N_38931,N_38411);
and U39196 (N_39196,N_38286,N_38698);
nor U39197 (N_39197,N_38954,N_38216);
and U39198 (N_39198,N_38557,N_38022);
nor U39199 (N_39199,N_38263,N_38582);
xnor U39200 (N_39200,N_38246,N_38941);
nor U39201 (N_39201,N_38396,N_38287);
xnor U39202 (N_39202,N_38750,N_38769);
nand U39203 (N_39203,N_38980,N_38322);
nand U39204 (N_39204,N_38533,N_38110);
nor U39205 (N_39205,N_38085,N_38345);
and U39206 (N_39206,N_38135,N_38195);
or U39207 (N_39207,N_38535,N_38985);
nand U39208 (N_39208,N_38835,N_38865);
nor U39209 (N_39209,N_38798,N_38326);
nor U39210 (N_39210,N_38207,N_38309);
xnor U39211 (N_39211,N_38190,N_38888);
nand U39212 (N_39212,N_38473,N_38754);
nor U39213 (N_39213,N_38150,N_38741);
xnor U39214 (N_39214,N_38445,N_38171);
nand U39215 (N_39215,N_38780,N_38849);
nand U39216 (N_39216,N_38016,N_38880);
nor U39217 (N_39217,N_38212,N_38296);
xnor U39218 (N_39218,N_38760,N_38862);
or U39219 (N_39219,N_38075,N_38781);
and U39220 (N_39220,N_38684,N_38530);
nor U39221 (N_39221,N_38424,N_38658);
nor U39222 (N_39222,N_38855,N_38555);
xnor U39223 (N_39223,N_38605,N_38911);
or U39224 (N_39224,N_38485,N_38097);
nor U39225 (N_39225,N_38903,N_38563);
nor U39226 (N_39226,N_38929,N_38556);
xor U39227 (N_39227,N_38919,N_38871);
or U39228 (N_39228,N_38817,N_38928);
xor U39229 (N_39229,N_38352,N_38325);
nor U39230 (N_39230,N_38571,N_38565);
nor U39231 (N_39231,N_38747,N_38918);
or U39232 (N_39232,N_38846,N_38279);
nand U39233 (N_39233,N_38220,N_38170);
or U39234 (N_39234,N_38026,N_38508);
nand U39235 (N_39235,N_38040,N_38578);
nor U39236 (N_39236,N_38054,N_38038);
nand U39237 (N_39237,N_38392,N_38073);
and U39238 (N_39238,N_38157,N_38414);
xor U39239 (N_39239,N_38181,N_38671);
nand U39240 (N_39240,N_38464,N_38249);
and U39241 (N_39241,N_38925,N_38441);
or U39242 (N_39242,N_38627,N_38323);
or U39243 (N_39243,N_38183,N_38087);
or U39244 (N_39244,N_38430,N_38544);
or U39245 (N_39245,N_38017,N_38081);
nand U39246 (N_39246,N_38205,N_38906);
nor U39247 (N_39247,N_38121,N_38625);
nor U39248 (N_39248,N_38148,N_38553);
nor U39249 (N_39249,N_38583,N_38493);
nand U39250 (N_39250,N_38008,N_38163);
nand U39251 (N_39251,N_38332,N_38704);
xor U39252 (N_39252,N_38005,N_38359);
xnor U39253 (N_39253,N_38808,N_38027);
nand U39254 (N_39254,N_38102,N_38731);
or U39255 (N_39255,N_38444,N_38709);
nor U39256 (N_39256,N_38247,N_38681);
xnor U39257 (N_39257,N_38541,N_38900);
or U39258 (N_39258,N_38071,N_38305);
or U39259 (N_39259,N_38111,N_38115);
or U39260 (N_39260,N_38319,N_38744);
xor U39261 (N_39261,N_38014,N_38433);
nor U39262 (N_39262,N_38634,N_38831);
and U39263 (N_39263,N_38289,N_38809);
and U39264 (N_39264,N_38879,N_38690);
and U39265 (N_39265,N_38630,N_38341);
or U39266 (N_39266,N_38876,N_38587);
nand U39267 (N_39267,N_38712,N_38118);
and U39268 (N_39268,N_38875,N_38963);
nand U39269 (N_39269,N_38952,N_38823);
and U39270 (N_39270,N_38891,N_38794);
or U39271 (N_39271,N_38320,N_38706);
nor U39272 (N_39272,N_38697,N_38644);
and U39273 (N_39273,N_38996,N_38222);
xnor U39274 (N_39274,N_38657,N_38812);
nor U39275 (N_39275,N_38113,N_38211);
nor U39276 (N_39276,N_38415,N_38546);
nand U39277 (N_39277,N_38299,N_38128);
and U39278 (N_39278,N_38640,N_38055);
or U39279 (N_39279,N_38368,N_38019);
and U39280 (N_39280,N_38394,N_38393);
nor U39281 (N_39281,N_38591,N_38994);
xnor U39282 (N_39282,N_38520,N_38265);
or U39283 (N_39283,N_38023,N_38079);
nor U39284 (N_39284,N_38969,N_38144);
or U39285 (N_39285,N_38943,N_38679);
nor U39286 (N_39286,N_38084,N_38512);
nand U39287 (N_39287,N_38645,N_38693);
xor U39288 (N_39288,N_38036,N_38974);
or U39289 (N_39289,N_38734,N_38883);
nand U39290 (N_39290,N_38161,N_38275);
xor U39291 (N_39291,N_38490,N_38268);
nand U39292 (N_39292,N_38491,N_38468);
nor U39293 (N_39293,N_38803,N_38337);
or U39294 (N_39294,N_38561,N_38355);
xor U39295 (N_39295,N_38847,N_38358);
or U39296 (N_39296,N_38710,N_38080);
or U39297 (N_39297,N_38635,N_38984);
nor U39298 (N_39298,N_38514,N_38449);
or U39299 (N_39299,N_38307,N_38045);
and U39300 (N_39300,N_38317,N_38000);
nor U39301 (N_39301,N_38398,N_38096);
xnor U39302 (N_39302,N_38142,N_38432);
xnor U39303 (N_39303,N_38748,N_38033);
or U39304 (N_39304,N_38434,N_38673);
and U39305 (N_39305,N_38899,N_38810);
and U39306 (N_39306,N_38302,N_38077);
and U39307 (N_39307,N_38824,N_38861);
xnor U39308 (N_39308,N_38532,N_38149);
and U39309 (N_39309,N_38294,N_38250);
and U39310 (N_39310,N_38437,N_38721);
nand U39311 (N_39311,N_38262,N_38347);
or U39312 (N_39312,N_38959,N_38417);
or U39313 (N_39313,N_38580,N_38219);
and U39314 (N_39314,N_38877,N_38418);
nor U39315 (N_39315,N_38397,N_38400);
nor U39316 (N_39316,N_38427,N_38451);
or U39317 (N_39317,N_38218,N_38059);
and U39318 (N_39318,N_38272,N_38225);
nand U39319 (N_39319,N_38025,N_38197);
nand U39320 (N_39320,N_38030,N_38868);
xnor U39321 (N_39321,N_38379,N_38821);
or U39322 (N_39322,N_38647,N_38652);
nand U39323 (N_39323,N_38811,N_38807);
nand U39324 (N_39324,N_38020,N_38926);
nor U39325 (N_39325,N_38227,N_38363);
or U39326 (N_39326,N_38801,N_38465);
or U39327 (N_39327,N_38156,N_38042);
and U39328 (N_39328,N_38991,N_38177);
xor U39329 (N_39329,N_38667,N_38562);
nand U39330 (N_39330,N_38614,N_38581);
nand U39331 (N_39331,N_38715,N_38147);
xor U39332 (N_39332,N_38264,N_38513);
nand U39333 (N_39333,N_38006,N_38457);
xnor U39334 (N_39334,N_38525,N_38463);
or U39335 (N_39335,N_38873,N_38106);
xnor U39336 (N_39336,N_38844,N_38977);
or U39337 (N_39337,N_38031,N_38762);
xor U39338 (N_39338,N_38505,N_38793);
nor U39339 (N_39339,N_38243,N_38350);
and U39340 (N_39340,N_38597,N_38682);
or U39341 (N_39341,N_38714,N_38843);
xor U39342 (N_39342,N_38585,N_38032);
and U39343 (N_39343,N_38366,N_38271);
and U39344 (N_39344,N_38431,N_38939);
xnor U39345 (N_39345,N_38007,N_38768);
or U39346 (N_39346,N_38766,N_38655);
xor U39347 (N_39347,N_38499,N_38428);
nor U39348 (N_39348,N_38921,N_38387);
or U39349 (N_39349,N_38013,N_38953);
nand U39350 (N_39350,N_38832,N_38015);
or U39351 (N_39351,N_38316,N_38815);
and U39352 (N_39352,N_38601,N_38740);
nand U39353 (N_39353,N_38814,N_38650);
nand U39354 (N_39354,N_38024,N_38048);
and U39355 (N_39355,N_38290,N_38568);
and U39356 (N_39356,N_38466,N_38934);
nand U39357 (N_39357,N_38435,N_38695);
xnor U39358 (N_39358,N_38771,N_38269);
nand U39359 (N_39359,N_38215,N_38622);
nor U39360 (N_39360,N_38129,N_38051);
or U39361 (N_39361,N_38044,N_38961);
nor U39362 (N_39362,N_38751,N_38141);
nor U39363 (N_39363,N_38238,N_38779);
xor U39364 (N_39364,N_38654,N_38333);
xnor U39365 (N_39365,N_38107,N_38399);
xor U39366 (N_39366,N_38596,N_38649);
or U39367 (N_39367,N_38251,N_38070);
and U39368 (N_39368,N_38588,N_38258);
xnor U39369 (N_39369,N_38413,N_38936);
or U39370 (N_39370,N_38502,N_38805);
nor U39371 (N_39371,N_38775,N_38898);
nand U39372 (N_39372,N_38386,N_38930);
nand U39373 (N_39373,N_38065,N_38987);
or U39374 (N_39374,N_38753,N_38285);
nand U39375 (N_39375,N_38728,N_38688);
nand U39376 (N_39376,N_38905,N_38981);
nand U39377 (N_39377,N_38737,N_38848);
and U39378 (N_39378,N_38909,N_38448);
nand U39379 (N_39379,N_38764,N_38501);
nand U39380 (N_39380,N_38702,N_38092);
and U39381 (N_39381,N_38178,N_38496);
or U39382 (N_39382,N_38659,N_38382);
nand U39383 (N_39383,N_38321,N_38011);
or U39384 (N_39384,N_38009,N_38273);
nand U39385 (N_39385,N_38611,N_38594);
nand U39386 (N_39386,N_38666,N_38390);
xor U39387 (N_39387,N_38365,N_38839);
and U39388 (N_39388,N_38117,N_38940);
or U39389 (N_39389,N_38927,N_38221);
nor U39390 (N_39390,N_38799,N_38242);
or U39391 (N_39391,N_38229,N_38371);
xnor U39392 (N_39392,N_38816,N_38572);
xnor U39393 (N_39393,N_38497,N_38730);
xnor U39394 (N_39394,N_38761,N_38757);
nand U39395 (N_39395,N_38356,N_38469);
or U39396 (N_39396,N_38786,N_38886);
or U39397 (N_39397,N_38274,N_38915);
or U39398 (N_39398,N_38703,N_38618);
xnor U39399 (N_39399,N_38989,N_38685);
xnor U39400 (N_39400,N_38509,N_38837);
nand U39401 (N_39401,N_38850,N_38370);
xor U39402 (N_39402,N_38471,N_38651);
nand U39403 (N_39403,N_38540,N_38789);
and U39404 (N_39404,N_38108,N_38599);
nor U39405 (N_39405,N_38833,N_38869);
nor U39406 (N_39406,N_38863,N_38840);
and U39407 (N_39407,N_38670,N_38283);
xor U39408 (N_39408,N_38864,N_38152);
nand U39409 (N_39409,N_38261,N_38962);
nor U39410 (N_39410,N_38199,N_38845);
or U39411 (N_39411,N_38770,N_38041);
xor U39412 (N_39412,N_38498,N_38346);
and U39413 (N_39413,N_38829,N_38752);
or U39414 (N_39414,N_38167,N_38516);
nor U39415 (N_39415,N_38641,N_38653);
xnor U39416 (N_39416,N_38029,N_38354);
nand U39417 (N_39417,N_38378,N_38057);
nand U39418 (N_39418,N_38573,N_38277);
and U39419 (N_39419,N_38169,N_38636);
or U39420 (N_39420,N_38543,N_38062);
xnor U39421 (N_39421,N_38705,N_38589);
xor U39422 (N_39422,N_38884,N_38487);
nor U39423 (N_39423,N_38923,N_38266);
or U39424 (N_39424,N_38951,N_38012);
nor U39425 (N_39425,N_38701,N_38402);
nand U39426 (N_39426,N_38838,N_38374);
nand U39427 (N_39427,N_38069,N_38988);
or U39428 (N_39428,N_38729,N_38384);
xor U39429 (N_39429,N_38724,N_38475);
xnor U39430 (N_39430,N_38646,N_38620);
xnor U39431 (N_39431,N_38389,N_38119);
nor U39432 (N_39432,N_38742,N_38401);
and U39433 (N_39433,N_38551,N_38893);
or U39434 (N_39434,N_38254,N_38995);
xnor U39435 (N_39435,N_38782,N_38339);
or U39436 (N_39436,N_38439,N_38907);
xor U39437 (N_39437,N_38192,N_38179);
or U39438 (N_39438,N_38997,N_38772);
and U39439 (N_39439,N_38968,N_38663);
xnor U39440 (N_39440,N_38722,N_38727);
nor U39441 (N_39441,N_38109,N_38570);
and U39442 (N_39442,N_38186,N_38203);
or U39443 (N_39443,N_38575,N_38615);
and U39444 (N_39444,N_38732,N_38175);
xor U39445 (N_39445,N_38637,N_38407);
and U39446 (N_39446,N_38074,N_38234);
xor U39447 (N_39447,N_38360,N_38672);
or U39448 (N_39448,N_38506,N_38343);
nor U39449 (N_39449,N_38639,N_38643);
xor U39450 (N_39450,N_38405,N_38329);
nand U39451 (N_39451,N_38922,N_38887);
and U39452 (N_39452,N_38248,N_38233);
nor U39453 (N_39453,N_38945,N_38914);
or U39454 (N_39454,N_38114,N_38626);
or U39455 (N_39455,N_38854,N_38308);
or U39456 (N_39456,N_38132,N_38039);
xnor U39457 (N_39457,N_38960,N_38607);
and U39458 (N_39458,N_38367,N_38700);
nand U39459 (N_39459,N_38720,N_38683);
nand U39460 (N_39460,N_38372,N_38711);
xnor U39461 (N_39461,N_38481,N_38713);
nor U39462 (N_39462,N_38795,N_38034);
nand U39463 (N_39463,N_38912,N_38256);
or U39464 (N_39464,N_38094,N_38164);
nor U39465 (N_39465,N_38103,N_38897);
or U39466 (N_39466,N_38486,N_38560);
nor U39467 (N_39467,N_38944,N_38788);
nand U39468 (N_39468,N_38298,N_38733);
and U39469 (N_39469,N_38213,N_38280);
nand U39470 (N_39470,N_38404,N_38334);
nand U39471 (N_39471,N_38327,N_38318);
nand U39472 (N_39472,N_38105,N_38395);
and U39473 (N_39473,N_38558,N_38214);
nor U39474 (N_39474,N_38507,N_38577);
and U39475 (N_39475,N_38408,N_38916);
nand U39476 (N_39476,N_38232,N_38758);
and U39477 (N_39477,N_38586,N_38340);
nand U39478 (N_39478,N_38692,N_38235);
nor U39479 (N_39479,N_38377,N_38143);
xnor U39480 (N_39480,N_38422,N_38545);
nor U39481 (N_39481,N_38612,N_38950);
xor U39482 (N_39482,N_38330,N_38136);
nor U39483 (N_39483,N_38842,N_38725);
xnor U39484 (N_39484,N_38851,N_38773);
and U39485 (N_39485,N_38311,N_38126);
xor U39486 (N_39486,N_38153,N_38526);
and U39487 (N_39487,N_38707,N_38086);
and U39488 (N_39488,N_38369,N_38391);
and U39489 (N_39489,N_38226,N_38970);
or U39490 (N_39490,N_38138,N_38674);
xor U39491 (N_39491,N_38083,N_38470);
or U39492 (N_39492,N_38223,N_38093);
and U39493 (N_39493,N_38282,N_38193);
xnor U39494 (N_39494,N_38278,N_38165);
nand U39495 (N_39495,N_38552,N_38777);
and U39496 (N_39496,N_38564,N_38385);
nand U39497 (N_39497,N_38276,N_38145);
xor U39498 (N_39498,N_38314,N_38576);
or U39499 (N_39499,N_38515,N_38774);
nand U39500 (N_39500,N_38019,N_38178);
or U39501 (N_39501,N_38614,N_38312);
and U39502 (N_39502,N_38767,N_38621);
nor U39503 (N_39503,N_38799,N_38761);
and U39504 (N_39504,N_38512,N_38102);
and U39505 (N_39505,N_38339,N_38265);
xor U39506 (N_39506,N_38082,N_38222);
and U39507 (N_39507,N_38387,N_38723);
and U39508 (N_39508,N_38790,N_38725);
or U39509 (N_39509,N_38744,N_38015);
xor U39510 (N_39510,N_38422,N_38125);
nand U39511 (N_39511,N_38266,N_38633);
xor U39512 (N_39512,N_38782,N_38403);
and U39513 (N_39513,N_38199,N_38594);
nor U39514 (N_39514,N_38313,N_38910);
nand U39515 (N_39515,N_38059,N_38585);
nand U39516 (N_39516,N_38906,N_38183);
and U39517 (N_39517,N_38842,N_38437);
nor U39518 (N_39518,N_38764,N_38894);
nor U39519 (N_39519,N_38312,N_38095);
nand U39520 (N_39520,N_38675,N_38651);
xnor U39521 (N_39521,N_38451,N_38061);
and U39522 (N_39522,N_38960,N_38883);
and U39523 (N_39523,N_38043,N_38814);
nand U39524 (N_39524,N_38672,N_38860);
or U39525 (N_39525,N_38476,N_38043);
or U39526 (N_39526,N_38690,N_38212);
nand U39527 (N_39527,N_38765,N_38862);
and U39528 (N_39528,N_38338,N_38634);
nand U39529 (N_39529,N_38910,N_38048);
nand U39530 (N_39530,N_38819,N_38883);
nor U39531 (N_39531,N_38079,N_38993);
nor U39532 (N_39532,N_38713,N_38444);
xor U39533 (N_39533,N_38466,N_38864);
nor U39534 (N_39534,N_38738,N_38613);
and U39535 (N_39535,N_38519,N_38636);
or U39536 (N_39536,N_38574,N_38204);
xnor U39537 (N_39537,N_38079,N_38392);
nand U39538 (N_39538,N_38580,N_38393);
nand U39539 (N_39539,N_38024,N_38012);
nor U39540 (N_39540,N_38185,N_38638);
and U39541 (N_39541,N_38635,N_38841);
nor U39542 (N_39542,N_38643,N_38556);
xnor U39543 (N_39543,N_38603,N_38193);
or U39544 (N_39544,N_38032,N_38508);
xnor U39545 (N_39545,N_38743,N_38665);
or U39546 (N_39546,N_38052,N_38416);
and U39547 (N_39547,N_38612,N_38947);
or U39548 (N_39548,N_38745,N_38789);
or U39549 (N_39549,N_38057,N_38424);
xnor U39550 (N_39550,N_38574,N_38286);
and U39551 (N_39551,N_38043,N_38186);
and U39552 (N_39552,N_38451,N_38501);
or U39553 (N_39553,N_38815,N_38250);
nor U39554 (N_39554,N_38460,N_38372);
or U39555 (N_39555,N_38846,N_38723);
xor U39556 (N_39556,N_38116,N_38436);
nor U39557 (N_39557,N_38657,N_38176);
xnor U39558 (N_39558,N_38250,N_38133);
nor U39559 (N_39559,N_38793,N_38444);
nor U39560 (N_39560,N_38581,N_38710);
xnor U39561 (N_39561,N_38693,N_38136);
nand U39562 (N_39562,N_38015,N_38778);
nor U39563 (N_39563,N_38458,N_38709);
and U39564 (N_39564,N_38214,N_38878);
xor U39565 (N_39565,N_38810,N_38438);
nand U39566 (N_39566,N_38651,N_38760);
nand U39567 (N_39567,N_38403,N_38603);
and U39568 (N_39568,N_38249,N_38330);
or U39569 (N_39569,N_38808,N_38555);
xor U39570 (N_39570,N_38970,N_38810);
and U39571 (N_39571,N_38652,N_38036);
xor U39572 (N_39572,N_38986,N_38448);
xor U39573 (N_39573,N_38004,N_38285);
nand U39574 (N_39574,N_38408,N_38849);
and U39575 (N_39575,N_38253,N_38178);
or U39576 (N_39576,N_38740,N_38818);
nand U39577 (N_39577,N_38290,N_38141);
xor U39578 (N_39578,N_38493,N_38546);
nand U39579 (N_39579,N_38610,N_38360);
and U39580 (N_39580,N_38104,N_38928);
or U39581 (N_39581,N_38553,N_38055);
xnor U39582 (N_39582,N_38395,N_38200);
nand U39583 (N_39583,N_38614,N_38513);
nor U39584 (N_39584,N_38922,N_38135);
or U39585 (N_39585,N_38049,N_38383);
nand U39586 (N_39586,N_38566,N_38024);
or U39587 (N_39587,N_38224,N_38075);
or U39588 (N_39588,N_38636,N_38902);
and U39589 (N_39589,N_38087,N_38525);
and U39590 (N_39590,N_38841,N_38863);
nand U39591 (N_39591,N_38015,N_38564);
or U39592 (N_39592,N_38175,N_38281);
nand U39593 (N_39593,N_38903,N_38430);
xnor U39594 (N_39594,N_38150,N_38514);
xor U39595 (N_39595,N_38481,N_38585);
nor U39596 (N_39596,N_38635,N_38346);
xnor U39597 (N_39597,N_38611,N_38322);
nor U39598 (N_39598,N_38591,N_38947);
nand U39599 (N_39599,N_38366,N_38615);
xnor U39600 (N_39600,N_38064,N_38935);
nor U39601 (N_39601,N_38491,N_38074);
and U39602 (N_39602,N_38035,N_38349);
nand U39603 (N_39603,N_38110,N_38315);
or U39604 (N_39604,N_38855,N_38888);
and U39605 (N_39605,N_38262,N_38697);
and U39606 (N_39606,N_38455,N_38012);
nor U39607 (N_39607,N_38914,N_38738);
nor U39608 (N_39608,N_38261,N_38262);
xnor U39609 (N_39609,N_38755,N_38470);
xnor U39610 (N_39610,N_38511,N_38338);
and U39611 (N_39611,N_38768,N_38664);
or U39612 (N_39612,N_38961,N_38023);
or U39613 (N_39613,N_38500,N_38466);
xnor U39614 (N_39614,N_38329,N_38419);
or U39615 (N_39615,N_38497,N_38306);
and U39616 (N_39616,N_38402,N_38143);
nand U39617 (N_39617,N_38004,N_38413);
xnor U39618 (N_39618,N_38866,N_38411);
and U39619 (N_39619,N_38850,N_38160);
and U39620 (N_39620,N_38031,N_38798);
xor U39621 (N_39621,N_38846,N_38765);
or U39622 (N_39622,N_38455,N_38512);
or U39623 (N_39623,N_38641,N_38903);
and U39624 (N_39624,N_38205,N_38974);
nand U39625 (N_39625,N_38258,N_38949);
nand U39626 (N_39626,N_38681,N_38742);
xnor U39627 (N_39627,N_38741,N_38481);
nor U39628 (N_39628,N_38733,N_38746);
nand U39629 (N_39629,N_38355,N_38728);
xor U39630 (N_39630,N_38108,N_38922);
nor U39631 (N_39631,N_38735,N_38757);
and U39632 (N_39632,N_38322,N_38096);
nand U39633 (N_39633,N_38286,N_38453);
or U39634 (N_39634,N_38085,N_38534);
nand U39635 (N_39635,N_38160,N_38989);
xnor U39636 (N_39636,N_38322,N_38948);
nand U39637 (N_39637,N_38454,N_38597);
and U39638 (N_39638,N_38598,N_38426);
and U39639 (N_39639,N_38526,N_38856);
nand U39640 (N_39640,N_38592,N_38835);
xor U39641 (N_39641,N_38172,N_38689);
and U39642 (N_39642,N_38548,N_38535);
xnor U39643 (N_39643,N_38532,N_38850);
nor U39644 (N_39644,N_38207,N_38698);
xor U39645 (N_39645,N_38692,N_38519);
and U39646 (N_39646,N_38012,N_38063);
xor U39647 (N_39647,N_38217,N_38218);
or U39648 (N_39648,N_38629,N_38651);
and U39649 (N_39649,N_38996,N_38231);
nand U39650 (N_39650,N_38111,N_38227);
or U39651 (N_39651,N_38783,N_38905);
xor U39652 (N_39652,N_38539,N_38175);
nor U39653 (N_39653,N_38209,N_38763);
or U39654 (N_39654,N_38126,N_38919);
or U39655 (N_39655,N_38593,N_38262);
xnor U39656 (N_39656,N_38276,N_38493);
xnor U39657 (N_39657,N_38652,N_38157);
and U39658 (N_39658,N_38644,N_38391);
nand U39659 (N_39659,N_38826,N_38394);
or U39660 (N_39660,N_38088,N_38774);
nand U39661 (N_39661,N_38846,N_38064);
or U39662 (N_39662,N_38019,N_38125);
xnor U39663 (N_39663,N_38379,N_38043);
nand U39664 (N_39664,N_38781,N_38517);
nand U39665 (N_39665,N_38248,N_38491);
or U39666 (N_39666,N_38105,N_38416);
nand U39667 (N_39667,N_38146,N_38460);
nand U39668 (N_39668,N_38295,N_38742);
or U39669 (N_39669,N_38334,N_38198);
nand U39670 (N_39670,N_38975,N_38661);
or U39671 (N_39671,N_38304,N_38695);
or U39672 (N_39672,N_38581,N_38923);
or U39673 (N_39673,N_38072,N_38241);
or U39674 (N_39674,N_38573,N_38586);
nor U39675 (N_39675,N_38383,N_38566);
xnor U39676 (N_39676,N_38655,N_38511);
nand U39677 (N_39677,N_38101,N_38857);
or U39678 (N_39678,N_38738,N_38546);
or U39679 (N_39679,N_38176,N_38873);
xnor U39680 (N_39680,N_38441,N_38361);
nor U39681 (N_39681,N_38357,N_38504);
xor U39682 (N_39682,N_38022,N_38398);
and U39683 (N_39683,N_38467,N_38930);
and U39684 (N_39684,N_38426,N_38655);
xnor U39685 (N_39685,N_38964,N_38148);
nand U39686 (N_39686,N_38823,N_38156);
or U39687 (N_39687,N_38275,N_38764);
nand U39688 (N_39688,N_38837,N_38404);
or U39689 (N_39689,N_38694,N_38221);
nor U39690 (N_39690,N_38619,N_38097);
and U39691 (N_39691,N_38571,N_38316);
nand U39692 (N_39692,N_38673,N_38889);
nor U39693 (N_39693,N_38518,N_38128);
nand U39694 (N_39694,N_38376,N_38676);
or U39695 (N_39695,N_38755,N_38371);
xnor U39696 (N_39696,N_38880,N_38424);
nor U39697 (N_39697,N_38673,N_38283);
nand U39698 (N_39698,N_38243,N_38731);
nand U39699 (N_39699,N_38951,N_38023);
or U39700 (N_39700,N_38280,N_38620);
and U39701 (N_39701,N_38460,N_38276);
or U39702 (N_39702,N_38216,N_38362);
and U39703 (N_39703,N_38498,N_38634);
nor U39704 (N_39704,N_38011,N_38079);
or U39705 (N_39705,N_38141,N_38068);
nor U39706 (N_39706,N_38378,N_38417);
or U39707 (N_39707,N_38696,N_38473);
nand U39708 (N_39708,N_38628,N_38724);
xnor U39709 (N_39709,N_38499,N_38925);
xnor U39710 (N_39710,N_38946,N_38702);
nand U39711 (N_39711,N_38270,N_38291);
or U39712 (N_39712,N_38495,N_38413);
xor U39713 (N_39713,N_38662,N_38646);
xor U39714 (N_39714,N_38767,N_38870);
xor U39715 (N_39715,N_38148,N_38007);
nor U39716 (N_39716,N_38294,N_38340);
xor U39717 (N_39717,N_38231,N_38314);
or U39718 (N_39718,N_38731,N_38131);
and U39719 (N_39719,N_38366,N_38990);
or U39720 (N_39720,N_38770,N_38502);
or U39721 (N_39721,N_38828,N_38402);
nand U39722 (N_39722,N_38224,N_38642);
xnor U39723 (N_39723,N_38395,N_38883);
or U39724 (N_39724,N_38897,N_38702);
or U39725 (N_39725,N_38941,N_38092);
nand U39726 (N_39726,N_38128,N_38712);
xnor U39727 (N_39727,N_38702,N_38760);
and U39728 (N_39728,N_38153,N_38815);
xnor U39729 (N_39729,N_38408,N_38256);
and U39730 (N_39730,N_38925,N_38056);
nor U39731 (N_39731,N_38206,N_38606);
and U39732 (N_39732,N_38848,N_38146);
and U39733 (N_39733,N_38305,N_38628);
nand U39734 (N_39734,N_38554,N_38895);
nor U39735 (N_39735,N_38190,N_38703);
nand U39736 (N_39736,N_38645,N_38887);
xnor U39737 (N_39737,N_38711,N_38979);
nor U39738 (N_39738,N_38805,N_38236);
and U39739 (N_39739,N_38690,N_38187);
xor U39740 (N_39740,N_38393,N_38544);
xnor U39741 (N_39741,N_38715,N_38927);
or U39742 (N_39742,N_38645,N_38782);
xor U39743 (N_39743,N_38380,N_38455);
and U39744 (N_39744,N_38489,N_38172);
nor U39745 (N_39745,N_38196,N_38952);
nand U39746 (N_39746,N_38265,N_38000);
nor U39747 (N_39747,N_38960,N_38846);
xnor U39748 (N_39748,N_38561,N_38489);
nand U39749 (N_39749,N_38256,N_38290);
or U39750 (N_39750,N_38334,N_38174);
or U39751 (N_39751,N_38278,N_38633);
or U39752 (N_39752,N_38769,N_38522);
and U39753 (N_39753,N_38329,N_38220);
nor U39754 (N_39754,N_38562,N_38237);
or U39755 (N_39755,N_38239,N_38588);
and U39756 (N_39756,N_38383,N_38576);
and U39757 (N_39757,N_38057,N_38027);
xnor U39758 (N_39758,N_38259,N_38079);
xor U39759 (N_39759,N_38630,N_38690);
nand U39760 (N_39760,N_38975,N_38915);
nand U39761 (N_39761,N_38983,N_38449);
nor U39762 (N_39762,N_38815,N_38864);
xnor U39763 (N_39763,N_38516,N_38037);
nand U39764 (N_39764,N_38321,N_38360);
or U39765 (N_39765,N_38788,N_38352);
xnor U39766 (N_39766,N_38018,N_38260);
xor U39767 (N_39767,N_38599,N_38625);
nor U39768 (N_39768,N_38030,N_38205);
nor U39769 (N_39769,N_38403,N_38507);
xnor U39770 (N_39770,N_38122,N_38619);
or U39771 (N_39771,N_38513,N_38801);
xnor U39772 (N_39772,N_38347,N_38088);
nand U39773 (N_39773,N_38813,N_38862);
xor U39774 (N_39774,N_38745,N_38299);
or U39775 (N_39775,N_38592,N_38417);
or U39776 (N_39776,N_38748,N_38723);
nand U39777 (N_39777,N_38206,N_38402);
or U39778 (N_39778,N_38802,N_38050);
and U39779 (N_39779,N_38619,N_38270);
nor U39780 (N_39780,N_38670,N_38171);
nand U39781 (N_39781,N_38518,N_38631);
nor U39782 (N_39782,N_38827,N_38852);
xor U39783 (N_39783,N_38994,N_38010);
nor U39784 (N_39784,N_38056,N_38730);
xnor U39785 (N_39785,N_38645,N_38753);
nor U39786 (N_39786,N_38937,N_38892);
and U39787 (N_39787,N_38972,N_38901);
nor U39788 (N_39788,N_38079,N_38344);
xnor U39789 (N_39789,N_38053,N_38788);
nand U39790 (N_39790,N_38757,N_38452);
or U39791 (N_39791,N_38678,N_38652);
nand U39792 (N_39792,N_38216,N_38309);
or U39793 (N_39793,N_38321,N_38380);
nand U39794 (N_39794,N_38843,N_38386);
or U39795 (N_39795,N_38159,N_38316);
nand U39796 (N_39796,N_38054,N_38467);
or U39797 (N_39797,N_38118,N_38066);
or U39798 (N_39798,N_38323,N_38776);
xnor U39799 (N_39799,N_38483,N_38047);
nor U39800 (N_39800,N_38517,N_38746);
nor U39801 (N_39801,N_38751,N_38690);
or U39802 (N_39802,N_38917,N_38706);
nor U39803 (N_39803,N_38082,N_38881);
nand U39804 (N_39804,N_38824,N_38910);
nand U39805 (N_39805,N_38690,N_38843);
nand U39806 (N_39806,N_38486,N_38119);
nor U39807 (N_39807,N_38811,N_38809);
and U39808 (N_39808,N_38405,N_38225);
or U39809 (N_39809,N_38704,N_38685);
xor U39810 (N_39810,N_38385,N_38692);
nand U39811 (N_39811,N_38107,N_38029);
or U39812 (N_39812,N_38799,N_38555);
and U39813 (N_39813,N_38748,N_38689);
xor U39814 (N_39814,N_38454,N_38287);
nor U39815 (N_39815,N_38377,N_38493);
or U39816 (N_39816,N_38761,N_38925);
and U39817 (N_39817,N_38101,N_38161);
or U39818 (N_39818,N_38953,N_38788);
nand U39819 (N_39819,N_38735,N_38496);
and U39820 (N_39820,N_38803,N_38327);
nor U39821 (N_39821,N_38983,N_38939);
and U39822 (N_39822,N_38518,N_38486);
or U39823 (N_39823,N_38432,N_38204);
xnor U39824 (N_39824,N_38154,N_38371);
xor U39825 (N_39825,N_38460,N_38896);
nand U39826 (N_39826,N_38985,N_38994);
and U39827 (N_39827,N_38038,N_38549);
and U39828 (N_39828,N_38595,N_38630);
or U39829 (N_39829,N_38153,N_38965);
nand U39830 (N_39830,N_38801,N_38902);
xnor U39831 (N_39831,N_38425,N_38573);
or U39832 (N_39832,N_38806,N_38100);
or U39833 (N_39833,N_38699,N_38857);
and U39834 (N_39834,N_38999,N_38788);
nand U39835 (N_39835,N_38907,N_38298);
xor U39836 (N_39836,N_38135,N_38494);
nor U39837 (N_39837,N_38646,N_38479);
nand U39838 (N_39838,N_38042,N_38768);
xor U39839 (N_39839,N_38652,N_38965);
or U39840 (N_39840,N_38705,N_38298);
nand U39841 (N_39841,N_38802,N_38571);
or U39842 (N_39842,N_38115,N_38320);
nand U39843 (N_39843,N_38304,N_38026);
nand U39844 (N_39844,N_38671,N_38996);
xor U39845 (N_39845,N_38831,N_38648);
nor U39846 (N_39846,N_38901,N_38231);
nor U39847 (N_39847,N_38100,N_38684);
nor U39848 (N_39848,N_38937,N_38748);
nand U39849 (N_39849,N_38825,N_38054);
nor U39850 (N_39850,N_38160,N_38206);
or U39851 (N_39851,N_38440,N_38591);
and U39852 (N_39852,N_38774,N_38314);
xor U39853 (N_39853,N_38160,N_38413);
and U39854 (N_39854,N_38758,N_38083);
nor U39855 (N_39855,N_38512,N_38301);
or U39856 (N_39856,N_38083,N_38929);
nor U39857 (N_39857,N_38997,N_38364);
nand U39858 (N_39858,N_38878,N_38329);
or U39859 (N_39859,N_38247,N_38310);
and U39860 (N_39860,N_38850,N_38840);
and U39861 (N_39861,N_38496,N_38352);
or U39862 (N_39862,N_38175,N_38380);
nand U39863 (N_39863,N_38097,N_38353);
nand U39864 (N_39864,N_38079,N_38304);
or U39865 (N_39865,N_38031,N_38189);
xor U39866 (N_39866,N_38966,N_38574);
or U39867 (N_39867,N_38356,N_38005);
or U39868 (N_39868,N_38935,N_38750);
nand U39869 (N_39869,N_38849,N_38778);
and U39870 (N_39870,N_38590,N_38539);
and U39871 (N_39871,N_38822,N_38123);
xor U39872 (N_39872,N_38186,N_38996);
nand U39873 (N_39873,N_38780,N_38145);
nand U39874 (N_39874,N_38189,N_38550);
nand U39875 (N_39875,N_38272,N_38614);
nor U39876 (N_39876,N_38518,N_38967);
nand U39877 (N_39877,N_38554,N_38945);
or U39878 (N_39878,N_38683,N_38442);
nand U39879 (N_39879,N_38905,N_38067);
and U39880 (N_39880,N_38113,N_38240);
nand U39881 (N_39881,N_38943,N_38441);
xnor U39882 (N_39882,N_38799,N_38070);
nand U39883 (N_39883,N_38024,N_38522);
xnor U39884 (N_39884,N_38252,N_38147);
xor U39885 (N_39885,N_38727,N_38007);
nand U39886 (N_39886,N_38804,N_38475);
or U39887 (N_39887,N_38166,N_38919);
or U39888 (N_39888,N_38962,N_38157);
nor U39889 (N_39889,N_38398,N_38944);
xor U39890 (N_39890,N_38929,N_38223);
nor U39891 (N_39891,N_38670,N_38894);
xor U39892 (N_39892,N_38810,N_38400);
and U39893 (N_39893,N_38665,N_38192);
xor U39894 (N_39894,N_38903,N_38273);
nand U39895 (N_39895,N_38528,N_38438);
xor U39896 (N_39896,N_38918,N_38634);
nor U39897 (N_39897,N_38116,N_38024);
or U39898 (N_39898,N_38383,N_38430);
and U39899 (N_39899,N_38968,N_38741);
or U39900 (N_39900,N_38538,N_38341);
or U39901 (N_39901,N_38398,N_38629);
or U39902 (N_39902,N_38317,N_38522);
nor U39903 (N_39903,N_38424,N_38084);
nor U39904 (N_39904,N_38633,N_38447);
or U39905 (N_39905,N_38337,N_38326);
xnor U39906 (N_39906,N_38340,N_38605);
nor U39907 (N_39907,N_38787,N_38472);
and U39908 (N_39908,N_38283,N_38248);
nor U39909 (N_39909,N_38363,N_38453);
and U39910 (N_39910,N_38543,N_38493);
xnor U39911 (N_39911,N_38689,N_38952);
and U39912 (N_39912,N_38674,N_38287);
nand U39913 (N_39913,N_38964,N_38749);
xor U39914 (N_39914,N_38325,N_38011);
nand U39915 (N_39915,N_38937,N_38828);
or U39916 (N_39916,N_38126,N_38184);
nor U39917 (N_39917,N_38297,N_38243);
nor U39918 (N_39918,N_38799,N_38109);
and U39919 (N_39919,N_38755,N_38383);
or U39920 (N_39920,N_38659,N_38645);
nor U39921 (N_39921,N_38795,N_38014);
and U39922 (N_39922,N_38321,N_38437);
or U39923 (N_39923,N_38972,N_38149);
nand U39924 (N_39924,N_38212,N_38461);
and U39925 (N_39925,N_38585,N_38749);
nand U39926 (N_39926,N_38637,N_38573);
and U39927 (N_39927,N_38720,N_38297);
xnor U39928 (N_39928,N_38937,N_38182);
and U39929 (N_39929,N_38429,N_38747);
and U39930 (N_39930,N_38072,N_38929);
and U39931 (N_39931,N_38946,N_38036);
xnor U39932 (N_39932,N_38210,N_38136);
nor U39933 (N_39933,N_38137,N_38076);
xor U39934 (N_39934,N_38654,N_38343);
nand U39935 (N_39935,N_38216,N_38298);
nor U39936 (N_39936,N_38715,N_38635);
and U39937 (N_39937,N_38132,N_38420);
nor U39938 (N_39938,N_38956,N_38279);
nor U39939 (N_39939,N_38818,N_38542);
xor U39940 (N_39940,N_38156,N_38876);
or U39941 (N_39941,N_38178,N_38309);
and U39942 (N_39942,N_38266,N_38521);
or U39943 (N_39943,N_38807,N_38666);
nor U39944 (N_39944,N_38942,N_38710);
and U39945 (N_39945,N_38589,N_38668);
and U39946 (N_39946,N_38220,N_38796);
nand U39947 (N_39947,N_38840,N_38892);
and U39948 (N_39948,N_38990,N_38751);
and U39949 (N_39949,N_38358,N_38617);
and U39950 (N_39950,N_38631,N_38206);
nand U39951 (N_39951,N_38359,N_38868);
xnor U39952 (N_39952,N_38671,N_38946);
or U39953 (N_39953,N_38777,N_38241);
nor U39954 (N_39954,N_38263,N_38596);
nand U39955 (N_39955,N_38011,N_38529);
xnor U39956 (N_39956,N_38466,N_38964);
and U39957 (N_39957,N_38154,N_38541);
xnor U39958 (N_39958,N_38455,N_38604);
nand U39959 (N_39959,N_38819,N_38631);
or U39960 (N_39960,N_38720,N_38001);
nand U39961 (N_39961,N_38067,N_38052);
nor U39962 (N_39962,N_38669,N_38270);
and U39963 (N_39963,N_38118,N_38336);
or U39964 (N_39964,N_38388,N_38407);
nor U39965 (N_39965,N_38656,N_38845);
and U39966 (N_39966,N_38204,N_38203);
and U39967 (N_39967,N_38759,N_38391);
nor U39968 (N_39968,N_38735,N_38452);
nand U39969 (N_39969,N_38689,N_38447);
nor U39970 (N_39970,N_38809,N_38516);
and U39971 (N_39971,N_38217,N_38188);
xor U39972 (N_39972,N_38088,N_38696);
or U39973 (N_39973,N_38068,N_38158);
xnor U39974 (N_39974,N_38452,N_38191);
or U39975 (N_39975,N_38093,N_38438);
or U39976 (N_39976,N_38036,N_38017);
nand U39977 (N_39977,N_38026,N_38678);
or U39978 (N_39978,N_38609,N_38768);
xor U39979 (N_39979,N_38924,N_38017);
and U39980 (N_39980,N_38515,N_38789);
nor U39981 (N_39981,N_38987,N_38965);
and U39982 (N_39982,N_38057,N_38743);
and U39983 (N_39983,N_38266,N_38401);
nand U39984 (N_39984,N_38874,N_38099);
nor U39985 (N_39985,N_38286,N_38857);
xor U39986 (N_39986,N_38694,N_38919);
nor U39987 (N_39987,N_38078,N_38866);
nor U39988 (N_39988,N_38647,N_38121);
and U39989 (N_39989,N_38556,N_38261);
xor U39990 (N_39990,N_38377,N_38261);
and U39991 (N_39991,N_38800,N_38817);
nor U39992 (N_39992,N_38132,N_38005);
nor U39993 (N_39993,N_38475,N_38599);
nand U39994 (N_39994,N_38841,N_38516);
or U39995 (N_39995,N_38462,N_38020);
or U39996 (N_39996,N_38507,N_38254);
and U39997 (N_39997,N_38421,N_38955);
nand U39998 (N_39998,N_38247,N_38423);
xor U39999 (N_39999,N_38931,N_38905);
or U40000 (N_40000,N_39691,N_39489);
xnor U40001 (N_40001,N_39420,N_39758);
nor U40002 (N_40002,N_39210,N_39279);
and U40003 (N_40003,N_39817,N_39077);
or U40004 (N_40004,N_39819,N_39061);
nor U40005 (N_40005,N_39715,N_39519);
or U40006 (N_40006,N_39222,N_39269);
or U40007 (N_40007,N_39886,N_39369);
and U40008 (N_40008,N_39080,N_39426);
nor U40009 (N_40009,N_39336,N_39518);
nand U40010 (N_40010,N_39789,N_39716);
and U40011 (N_40011,N_39864,N_39233);
or U40012 (N_40012,N_39836,N_39616);
nand U40013 (N_40013,N_39938,N_39728);
or U40014 (N_40014,N_39692,N_39153);
xor U40015 (N_40015,N_39445,N_39044);
and U40016 (N_40016,N_39840,N_39257);
nor U40017 (N_40017,N_39074,N_39262);
nor U40018 (N_40018,N_39601,N_39820);
or U40019 (N_40019,N_39260,N_39376);
or U40020 (N_40020,N_39804,N_39893);
nor U40021 (N_40021,N_39413,N_39200);
or U40022 (N_40022,N_39071,N_39337);
and U40023 (N_40023,N_39742,N_39603);
nor U40024 (N_40024,N_39748,N_39435);
and U40025 (N_40025,N_39190,N_39466);
and U40026 (N_40026,N_39665,N_39122);
and U40027 (N_40027,N_39462,N_39319);
nor U40028 (N_40028,N_39261,N_39460);
xnor U40029 (N_40029,N_39575,N_39471);
nor U40030 (N_40030,N_39680,N_39750);
xor U40031 (N_40031,N_39853,N_39476);
and U40032 (N_40032,N_39069,N_39300);
or U40033 (N_40033,N_39835,N_39670);
xnor U40034 (N_40034,N_39457,N_39405);
or U40035 (N_40035,N_39366,N_39999);
nor U40036 (N_40036,N_39914,N_39009);
nor U40037 (N_40037,N_39671,N_39125);
and U40038 (N_40038,N_39059,N_39736);
or U40039 (N_40039,N_39150,N_39983);
xnor U40040 (N_40040,N_39038,N_39106);
nand U40041 (N_40041,N_39378,N_39577);
nor U40042 (N_40042,N_39424,N_39929);
xnor U40043 (N_40043,N_39121,N_39622);
xor U40044 (N_40044,N_39774,N_39375);
nand U40045 (N_40045,N_39990,N_39340);
and U40046 (N_40046,N_39267,N_39851);
and U40047 (N_40047,N_39975,N_39907);
nand U40048 (N_40048,N_39047,N_39952);
and U40049 (N_40049,N_39868,N_39097);
nor U40050 (N_40050,N_39474,N_39613);
xor U40051 (N_40051,N_39278,N_39033);
nand U40052 (N_40052,N_39625,N_39875);
or U40053 (N_40053,N_39783,N_39865);
nor U40054 (N_40054,N_39795,N_39672);
nor U40055 (N_40055,N_39530,N_39018);
and U40056 (N_40056,N_39107,N_39318);
nor U40057 (N_40057,N_39228,N_39548);
or U40058 (N_40058,N_39358,N_39640);
nand U40059 (N_40059,N_39843,N_39807);
nand U40060 (N_40060,N_39932,N_39484);
or U40061 (N_40061,N_39064,N_39141);
nand U40062 (N_40062,N_39173,N_39049);
and U40063 (N_40063,N_39645,N_39759);
nor U40064 (N_40064,N_39100,N_39646);
and U40065 (N_40065,N_39747,N_39446);
or U40066 (N_40066,N_39879,N_39172);
nand U40067 (N_40067,N_39123,N_39986);
nand U40068 (N_40068,N_39880,N_39571);
nor U40069 (N_40069,N_39197,N_39524);
nand U40070 (N_40070,N_39487,N_39315);
nor U40071 (N_40071,N_39828,N_39937);
nand U40072 (N_40072,N_39862,N_39175);
xor U40073 (N_40073,N_39612,N_39838);
and U40074 (N_40074,N_39654,N_39627);
nor U40075 (N_40075,N_39958,N_39338);
or U40076 (N_40076,N_39877,N_39598);
nand U40077 (N_40077,N_39913,N_39730);
and U40078 (N_40078,N_39634,N_39272);
xor U40079 (N_40079,N_39493,N_39270);
xor U40080 (N_40080,N_39285,N_39895);
nand U40081 (N_40081,N_39738,N_39459);
nand U40082 (N_40082,N_39762,N_39784);
nor U40083 (N_40083,N_39468,N_39442);
nor U40084 (N_40084,N_39023,N_39511);
xnor U40085 (N_40085,N_39361,N_39666);
nand U40086 (N_40086,N_39198,N_39689);
or U40087 (N_40087,N_39731,N_39970);
nor U40088 (N_40088,N_39642,N_39024);
or U40089 (N_40089,N_39096,N_39604);
nand U40090 (N_40090,N_39507,N_39635);
nand U40091 (N_40091,N_39700,N_39355);
or U40092 (N_40092,N_39771,N_39697);
xor U40093 (N_40093,N_39332,N_39707);
or U40094 (N_40094,N_39385,N_39391);
nand U40095 (N_40095,N_39720,N_39191);
xor U40096 (N_40096,N_39335,N_39246);
or U40097 (N_40097,N_39407,N_39330);
xor U40098 (N_40098,N_39718,N_39239);
or U40099 (N_40099,N_39087,N_39933);
nor U40100 (N_40100,N_39559,N_39713);
xnor U40101 (N_40101,N_39354,N_39576);
nand U40102 (N_40102,N_39786,N_39223);
or U40103 (N_40103,N_39109,N_39339);
nor U40104 (N_40104,N_39266,N_39372);
and U40105 (N_40105,N_39959,N_39972);
and U40106 (N_40106,N_39137,N_39167);
xor U40107 (N_40107,N_39360,N_39207);
xnor U40108 (N_40108,N_39485,N_39590);
nand U40109 (N_40109,N_39194,N_39565);
or U40110 (N_40110,N_39942,N_39154);
nand U40111 (N_40111,N_39093,N_39650);
nor U40112 (N_40112,N_39146,N_39637);
and U40113 (N_40113,N_39920,N_39963);
nand U40114 (N_40114,N_39142,N_39925);
nor U40115 (N_40115,N_39039,N_39132);
or U40116 (N_40116,N_39823,N_39651);
or U40117 (N_40117,N_39788,N_39714);
or U40118 (N_40118,N_39904,N_39652);
xnor U40119 (N_40119,N_39281,N_39701);
nor U40120 (N_40120,N_39866,N_39981);
or U40121 (N_40121,N_39912,N_39967);
nor U40122 (N_40122,N_39947,N_39702);
nor U40123 (N_40123,N_39854,N_39240);
and U40124 (N_40124,N_39472,N_39884);
nor U40125 (N_40125,N_39486,N_39745);
xnor U40126 (N_40126,N_39439,N_39301);
or U40127 (N_40127,N_39863,N_39169);
and U40128 (N_40128,N_39244,N_39016);
nand U40129 (N_40129,N_39082,N_39367);
or U40130 (N_40130,N_39067,N_39192);
or U40131 (N_40131,N_39328,N_39594);
or U40132 (N_40132,N_39220,N_39481);
or U40133 (N_40133,N_39325,N_39722);
or U40134 (N_40134,N_39253,N_39555);
xor U40135 (N_40135,N_39534,N_39756);
xor U40136 (N_40136,N_39248,N_39583);
nand U40137 (N_40137,N_39140,N_39615);
or U40138 (N_40138,N_39841,N_39757);
and U40139 (N_40139,N_39213,N_39461);
and U40140 (N_40140,N_39664,N_39229);
or U40141 (N_40141,N_39112,N_39569);
or U40142 (N_40142,N_39578,N_39909);
nor U40143 (N_40143,N_39363,N_39293);
or U40144 (N_40144,N_39790,N_39091);
nand U40145 (N_40145,N_39996,N_39221);
nor U40146 (N_40146,N_39948,N_39013);
xor U40147 (N_40147,N_39867,N_39626);
xnor U40148 (N_40148,N_39412,N_39582);
nor U40149 (N_40149,N_39303,N_39292);
nand U40150 (N_40150,N_39709,N_39552);
and U40151 (N_40151,N_39079,N_39860);
xor U40152 (N_40152,N_39208,N_39526);
or U40153 (N_40153,N_39900,N_39621);
nor U40154 (N_40154,N_39316,N_39195);
nand U40155 (N_40155,N_39124,N_39885);
or U40156 (N_40156,N_39170,N_39663);
nand U40157 (N_40157,N_39035,N_39247);
nor U40158 (N_40158,N_39066,N_39464);
or U40159 (N_40159,N_39547,N_39283);
or U40160 (N_40160,N_39176,N_39830);
nor U40161 (N_40161,N_39133,N_39095);
nand U40162 (N_40162,N_39139,N_39452);
nor U40163 (N_40163,N_39776,N_39961);
and U40164 (N_40164,N_39818,N_39591);
nor U40165 (N_40165,N_39500,N_39015);
nor U40166 (N_40166,N_39892,N_39595);
and U40167 (N_40167,N_39055,N_39393);
nor U40168 (N_40168,N_39902,N_39644);
nand U40169 (N_40169,N_39764,N_39373);
nor U40170 (N_40170,N_39772,N_39307);
nand U40171 (N_40171,N_39159,N_39546);
or U40172 (N_40172,N_39881,N_39168);
and U40173 (N_40173,N_39145,N_39342);
nand U40174 (N_40174,N_39374,N_39188);
and U40175 (N_40175,N_39638,N_39432);
and U40176 (N_40176,N_39014,N_39943);
nand U40177 (N_40177,N_39110,N_39988);
or U40178 (N_40178,N_39628,N_39636);
nor U40179 (N_40179,N_39660,N_39787);
xnor U40180 (N_40180,N_39703,N_39353);
nand U40181 (N_40181,N_39906,N_39538);
and U40182 (N_40182,N_39602,N_39331);
or U40183 (N_40183,N_39026,N_39888);
nand U40184 (N_40184,N_39219,N_39450);
nor U40185 (N_40185,N_39889,N_39147);
or U40186 (N_40186,N_39419,N_39314);
and U40187 (N_40187,N_39418,N_39515);
nand U40188 (N_40188,N_39781,N_39028);
or U40189 (N_40189,N_39825,N_39951);
nor U40190 (N_40190,N_39490,N_39686);
and U40191 (N_40191,N_39973,N_39550);
nand U40192 (N_40192,N_39311,N_39725);
nand U40193 (N_40193,N_39076,N_39404);
or U40194 (N_40194,N_39989,N_39099);
xor U40195 (N_40195,N_39451,N_39586);
and U40196 (N_40196,N_39971,N_39227);
xor U40197 (N_40197,N_39429,N_39679);
nand U40198 (N_40198,N_39231,N_39827);
or U40199 (N_40199,N_39966,N_39276);
and U40200 (N_40200,N_39763,N_39201);
or U40201 (N_40201,N_39072,N_39847);
or U40202 (N_40202,N_39286,N_39144);
xnor U40203 (N_40203,N_39876,N_39873);
xor U40204 (N_40204,N_39580,N_39540);
nand U40205 (N_40205,N_39858,N_39428);
and U40206 (N_40206,N_39822,N_39704);
and U40207 (N_40207,N_39667,N_39805);
and U40208 (N_40208,N_39799,N_39092);
xor U40209 (N_40209,N_39245,N_39088);
nand U40210 (N_40210,N_39225,N_39506);
or U40211 (N_40211,N_39002,N_39510);
or U40212 (N_40212,N_39127,N_39859);
xor U40213 (N_40213,N_39152,N_39415);
xnor U40214 (N_40214,N_39918,N_39006);
nand U40215 (N_40215,N_39890,N_39782);
and U40216 (N_40216,N_39870,N_39681);
and U40217 (N_40217,N_39921,N_39105);
nand U40218 (N_40218,N_39766,N_39574);
and U40219 (N_40219,N_39903,N_39045);
or U40220 (N_40220,N_39078,N_39754);
nand U40221 (N_40221,N_39299,N_39400);
nor U40222 (N_40222,N_39242,N_39196);
nand U40223 (N_40223,N_39987,N_39648);
and U40224 (N_40224,N_39941,N_39536);
nor U40225 (N_40225,N_39905,N_39206);
nand U40226 (N_40226,N_39848,N_39955);
nand U40227 (N_40227,N_39688,N_39950);
nand U40228 (N_40228,N_39304,N_39297);
nor U40229 (N_40229,N_39345,N_39183);
or U40230 (N_40230,N_39042,N_39492);
xor U40231 (N_40231,N_39641,N_39998);
nor U40232 (N_40232,N_39923,N_39148);
nand U40233 (N_40233,N_39114,N_39050);
and U40234 (N_40234,N_39698,N_39544);
or U40235 (N_40235,N_39031,N_39934);
or U40236 (N_40236,N_39824,N_39003);
nand U40237 (N_40237,N_39505,N_39268);
and U40238 (N_40238,N_39814,N_39346);
nor U40239 (N_40239,N_39632,N_39562);
or U40240 (N_40240,N_39513,N_39592);
nor U40241 (N_40241,N_39327,N_39694);
nor U40242 (N_40242,N_39726,N_39560);
and U40243 (N_40243,N_39241,N_39509);
nand U40244 (N_40244,N_39855,N_39732);
nor U40245 (N_40245,N_39273,N_39364);
and U40246 (N_40246,N_39563,N_39108);
and U40247 (N_40247,N_39037,N_39699);
xor U40248 (N_40248,N_39089,N_39517);
or U40249 (N_40249,N_39395,N_39532);
or U40250 (N_40250,N_39178,N_39527);
and U40251 (N_40251,N_39915,N_39803);
xnor U40252 (N_40252,N_39287,N_39712);
xnor U40253 (N_40253,N_39102,N_39901);
nor U40254 (N_40254,N_39496,N_39073);
nand U40255 (N_40255,N_39090,N_39554);
nand U40256 (N_40256,N_39005,N_39832);
and U40257 (N_40257,N_39690,N_39994);
or U40258 (N_40258,N_39796,N_39744);
xor U40259 (N_40259,N_39065,N_39727);
nor U40260 (N_40260,N_39589,N_39677);
xor U40261 (N_40261,N_39643,N_39440);
nor U40262 (N_40262,N_39522,N_39392);
xor U40263 (N_40263,N_39135,N_39968);
or U40264 (N_40264,N_39081,N_39349);
and U40265 (N_40265,N_39441,N_39623);
or U40266 (N_40266,N_39498,N_39166);
or U40267 (N_40267,N_39463,N_39323);
or U40268 (N_40268,N_39977,N_39070);
or U40269 (N_40269,N_39120,N_39414);
xnor U40270 (N_40270,N_39041,N_39422);
or U40271 (N_40271,N_39542,N_39992);
and U40272 (N_40272,N_39203,N_39760);
and U40273 (N_40273,N_39683,N_39734);
nand U40274 (N_40274,N_39953,N_39852);
xnor U40275 (N_40275,N_39662,N_39402);
nor U40276 (N_40276,N_39477,N_39842);
and U40277 (N_40277,N_39911,N_39309);
xor U40278 (N_40278,N_39751,N_39810);
and U40279 (N_40279,N_39030,N_39205);
and U40280 (N_40280,N_39383,N_39386);
nand U40281 (N_40281,N_39020,N_39394);
nor U40282 (N_40282,N_39593,N_39543);
nor U40283 (N_40283,N_39557,N_39249);
or U40284 (N_40284,N_39291,N_39104);
and U40285 (N_40285,N_39313,N_39011);
xor U40286 (N_40286,N_39343,N_39837);
nand U40287 (N_40287,N_39797,N_39356);
nor U40288 (N_40288,N_39379,N_39111);
or U40289 (N_40289,N_39288,N_39611);
and U40290 (N_40290,N_39978,N_39658);
or U40291 (N_40291,N_39344,N_39381);
nand U40292 (N_40292,N_39199,N_39237);
xor U40293 (N_40293,N_39465,N_39357);
and U40294 (N_40294,N_39034,N_39816);
xor U40295 (N_40295,N_39721,N_39310);
xnor U40296 (N_40296,N_39480,N_39926);
or U40297 (N_40297,N_39370,N_39036);
xor U40298 (N_40298,N_39695,N_39899);
xor U40299 (N_40299,N_39606,N_39600);
nor U40300 (N_40300,N_39408,N_39607);
and U40301 (N_40301,N_39608,N_39794);
or U40302 (N_40302,N_39957,N_39919);
xnor U40303 (N_40303,N_39693,N_39164);
or U40304 (N_40304,N_39813,N_39597);
nand U40305 (N_40305,N_39897,N_39417);
nand U40306 (N_40306,N_39617,N_39570);
xor U40307 (N_40307,N_39305,N_39553);
nor U40308 (N_40308,N_39226,N_39755);
nor U40309 (N_40309,N_39215,N_39204);
nor U40310 (N_40310,N_39054,N_39705);
nand U40311 (N_40311,N_39962,N_39639);
and U40312 (N_40312,N_39320,N_39083);
and U40313 (N_40313,N_39630,N_39334);
xnor U40314 (N_40314,N_39211,N_39746);
or U40315 (N_40315,N_39230,N_39098);
and U40316 (N_40316,N_39431,N_39785);
nor U40317 (N_40317,N_39541,N_39985);
nor U40318 (N_40318,N_39296,N_39812);
xnor U40319 (N_40319,N_39051,N_39454);
and U40320 (N_40320,N_39295,N_39368);
or U40321 (N_40321,N_39584,N_39214);
xor U40322 (N_40322,N_39321,N_39238);
xor U40323 (N_40323,N_39350,N_39528);
xnor U40324 (N_40324,N_39117,N_39741);
nand U40325 (N_40325,N_39512,N_39891);
nand U40326 (N_40326,N_39251,N_39302);
nor U40327 (N_40327,N_39850,N_39609);
or U40328 (N_40328,N_39647,N_39488);
nand U40329 (N_40329,N_39908,N_39060);
and U40330 (N_40330,N_39032,N_39619);
and U40331 (N_40331,N_39022,N_39898);
and U40332 (N_40332,N_39134,N_39217);
and U40333 (N_40333,N_39456,N_39399);
or U40334 (N_40334,N_39516,N_39052);
xnor U40335 (N_40335,N_39928,N_39421);
nor U40336 (N_40336,N_39556,N_39012);
and U40337 (N_40337,N_39004,N_39737);
nand U40338 (N_40338,N_39403,N_39371);
and U40339 (N_40339,N_39174,N_39284);
xor U40340 (N_40340,N_39735,N_39155);
nand U40341 (N_40341,N_39263,N_39927);
nand U40342 (N_40342,N_39682,N_39740);
xnor U40343 (N_40343,N_39380,N_39482);
nor U40344 (N_40344,N_39749,N_39685);
and U40345 (N_40345,N_39160,N_39444);
or U40346 (N_40346,N_39479,N_39684);
and U40347 (N_40347,N_39653,N_39218);
xnor U40348 (N_40348,N_39136,N_39483);
nor U40349 (N_40349,N_39765,N_39043);
and U40350 (N_40350,N_39533,N_39649);
or U40351 (N_40351,N_39365,N_39521);
and U40352 (N_40352,N_39294,N_39655);
or U40353 (N_40353,N_39171,N_39956);
and U40354 (N_40354,N_39277,N_39433);
or U40355 (N_40355,N_39599,N_39475);
or U40356 (N_40356,N_39008,N_39235);
nor U40357 (N_40357,N_39839,N_39068);
nand U40358 (N_40358,N_39455,N_39558);
nor U40359 (N_40359,N_39029,N_39793);
xnor U40360 (N_40360,N_39572,N_39529);
nand U40361 (N_40361,N_39306,N_39128);
nor U40362 (N_40362,N_39775,N_39409);
xnor U40363 (N_40363,N_39362,N_39676);
or U40364 (N_40364,N_39605,N_39057);
nand U40365 (N_40365,N_39499,N_39800);
nand U40366 (N_40366,N_39675,N_39878);
nor U40367 (N_40367,N_39872,N_39752);
nand U40368 (N_40368,N_39719,N_39945);
xnor U40369 (N_40369,N_39232,N_39425);
and U40370 (N_40370,N_39503,N_39007);
nor U40371 (N_40371,N_39769,N_39258);
xnor U40372 (N_40372,N_39778,N_39177);
nor U40373 (N_40373,N_39856,N_39341);
xor U40374 (N_40374,N_39857,N_39438);
nand U40375 (N_40375,N_39165,N_39523);
nor U40376 (N_40376,N_39129,N_39290);
or U40377 (N_40377,N_39779,N_39791);
and U40378 (N_40378,N_39976,N_39661);
nand U40379 (N_40379,N_39163,N_39917);
xor U40380 (N_40380,N_39668,N_39115);
or U40381 (N_40381,N_39255,N_39935);
and U40382 (N_40382,N_39243,N_39469);
nor U40383 (N_40383,N_39806,N_39656);
xnor U40384 (N_40384,N_39678,N_39001);
and U40385 (N_40385,N_39831,N_39874);
and U40386 (N_40386,N_39631,N_39845);
nor U40387 (N_40387,N_39495,N_39733);
nor U40388 (N_40388,N_39411,N_39436);
nor U40389 (N_40389,N_39922,N_39494);
xnor U40390 (N_40390,N_39473,N_39186);
nand U40391 (N_40391,N_39931,N_39618);
and U40392 (N_40392,N_39182,N_39629);
and U40393 (N_40393,N_39025,N_39596);
nand U40394 (N_40394,N_39317,N_39882);
and U40395 (N_40395,N_39549,N_39833);
nor U40396 (N_40396,N_39869,N_39377);
nor U40397 (N_40397,N_39162,N_39130);
or U40398 (N_40398,N_39777,N_39298);
and U40399 (N_40399,N_39535,N_39021);
nor U40400 (N_40400,N_39551,N_39984);
nand U40401 (N_40401,N_39780,N_39390);
xnor U40402 (N_40402,N_39430,N_39062);
and U40403 (N_40403,N_39657,N_39053);
and U40404 (N_40404,N_39940,N_39470);
nand U40405 (N_40405,N_39193,N_39252);
nor U40406 (N_40406,N_39161,N_39180);
nor U40407 (N_40407,N_39965,N_39158);
nand U40408 (N_40408,N_39113,N_39561);
and U40409 (N_40409,N_39579,N_39520);
xor U40410 (N_40410,N_39567,N_39706);
nor U40411 (N_40411,N_39761,N_39265);
or U40412 (N_40412,N_39960,N_39324);
nand U40413 (N_40413,N_39729,N_39815);
nand U40414 (N_40414,N_39116,N_39861);
xnor U40415 (N_40415,N_39808,N_39185);
nand U40416 (N_40416,N_39410,N_39620);
nand U40417 (N_40417,N_39674,N_39236);
nand U40418 (N_40418,N_39388,N_39406);
nor U40419 (N_40419,N_39119,N_39449);
xnor U40420 (N_40420,N_39181,N_39149);
xnor U40421 (N_40421,N_39504,N_39212);
or U40422 (N_40422,N_39724,N_39216);
nor U40423 (N_40423,N_39447,N_39352);
and U40424 (N_40424,N_39143,N_39673);
and U40425 (N_40425,N_39669,N_39993);
xor U40426 (N_40426,N_39058,N_39086);
and U40427 (N_40427,N_39946,N_39896);
xor U40428 (N_40428,N_39017,N_39275);
nor U40429 (N_40429,N_39514,N_39768);
or U40430 (N_40430,N_39739,N_39282);
or U40431 (N_40431,N_39202,N_39659);
or U40432 (N_40432,N_39351,N_39710);
nand U40433 (N_40433,N_39184,N_39974);
and U40434 (N_40434,N_39924,N_39254);
nand U40435 (N_40435,N_39846,N_39312);
xnor U40436 (N_40436,N_39792,N_39995);
nor U40437 (N_40437,N_39497,N_39834);
and U40438 (N_40438,N_39046,N_39401);
and U40439 (N_40439,N_39930,N_39347);
nand U40440 (N_40440,N_39770,N_39333);
nor U40441 (N_40441,N_39274,N_39743);
xor U40442 (N_40442,N_39910,N_39849);
nand U40443 (N_40443,N_39991,N_39964);
nand U40444 (N_40444,N_39936,N_39767);
or U40445 (N_40445,N_39398,N_39453);
nand U40446 (N_40446,N_39384,N_39508);
or U40447 (N_40447,N_39537,N_39587);
nand U40448 (N_40448,N_39101,N_39610);
or U40449 (N_40449,N_39063,N_39573);
or U40450 (N_40450,N_39085,N_39802);
nand U40451 (N_40451,N_39434,N_39773);
nand U40452 (N_40452,N_39491,N_39151);
or U40453 (N_40453,N_39944,N_39939);
and U40454 (N_40454,N_39883,N_39348);
nor U40455 (N_40455,N_39382,N_39437);
and U40456 (N_40456,N_39189,N_39711);
nand U40457 (N_40457,N_39040,N_39187);
nor U40458 (N_40458,N_39322,N_39256);
and U40459 (N_40459,N_39916,N_39126);
or U40460 (N_40460,N_39844,N_39250);
xnor U40461 (N_40461,N_39633,N_39209);
and U40462 (N_40462,N_39156,N_39717);
and U40463 (N_40463,N_39568,N_39954);
nor U40464 (N_40464,N_39056,N_39359);
nand U40465 (N_40465,N_39949,N_39826);
nor U40466 (N_40466,N_39753,N_39118);
nand U40467 (N_40467,N_39588,N_39396);
xor U40468 (N_40468,N_39614,N_39798);
nor U40469 (N_40469,N_39131,N_39427);
nor U40470 (N_40470,N_39969,N_39525);
or U40471 (N_40471,N_39821,N_39871);
or U40472 (N_40472,N_39389,N_39894);
nor U40473 (N_40473,N_39458,N_39010);
nor U40474 (N_40474,N_39478,N_39416);
or U40475 (N_40475,N_39075,N_39019);
nand U40476 (N_40476,N_39264,N_39501);
nor U40477 (N_40477,N_39423,N_39084);
nand U40478 (N_40478,N_39289,N_39027);
or U40479 (N_40479,N_39696,N_39138);
or U40480 (N_40480,N_39708,N_39809);
or U40481 (N_40481,N_39448,N_39980);
nor U40482 (N_40482,N_39531,N_39624);
or U40483 (N_40483,N_39581,N_39224);
and U40484 (N_40484,N_39000,N_39179);
nand U40485 (N_40485,N_39326,N_39397);
or U40486 (N_40486,N_39157,N_39271);
and U40487 (N_40487,N_39564,N_39094);
xnor U40488 (N_40488,N_39801,N_39887);
xor U40489 (N_40489,N_39997,N_39259);
nand U40490 (N_40490,N_39585,N_39539);
xnor U40491 (N_40491,N_39723,N_39234);
or U40492 (N_40492,N_39048,N_39329);
nor U40493 (N_40493,N_39502,N_39443);
and U40494 (N_40494,N_39467,N_39387);
xor U40495 (N_40495,N_39308,N_39979);
nor U40496 (N_40496,N_39545,N_39566);
xor U40497 (N_40497,N_39982,N_39687);
xnor U40498 (N_40498,N_39280,N_39829);
xor U40499 (N_40499,N_39103,N_39811);
nor U40500 (N_40500,N_39962,N_39260);
and U40501 (N_40501,N_39988,N_39912);
nor U40502 (N_40502,N_39221,N_39677);
xnor U40503 (N_40503,N_39031,N_39550);
nor U40504 (N_40504,N_39369,N_39800);
or U40505 (N_40505,N_39260,N_39255);
and U40506 (N_40506,N_39620,N_39033);
nor U40507 (N_40507,N_39475,N_39276);
nand U40508 (N_40508,N_39517,N_39009);
nand U40509 (N_40509,N_39101,N_39148);
nand U40510 (N_40510,N_39495,N_39870);
nand U40511 (N_40511,N_39302,N_39362);
and U40512 (N_40512,N_39576,N_39864);
and U40513 (N_40513,N_39116,N_39899);
xnor U40514 (N_40514,N_39093,N_39417);
nand U40515 (N_40515,N_39533,N_39237);
xnor U40516 (N_40516,N_39376,N_39547);
nor U40517 (N_40517,N_39162,N_39171);
nor U40518 (N_40518,N_39479,N_39919);
and U40519 (N_40519,N_39857,N_39384);
nand U40520 (N_40520,N_39560,N_39142);
xnor U40521 (N_40521,N_39364,N_39094);
nand U40522 (N_40522,N_39472,N_39025);
and U40523 (N_40523,N_39950,N_39480);
nor U40524 (N_40524,N_39528,N_39338);
and U40525 (N_40525,N_39177,N_39640);
nor U40526 (N_40526,N_39992,N_39690);
nor U40527 (N_40527,N_39945,N_39648);
or U40528 (N_40528,N_39504,N_39774);
and U40529 (N_40529,N_39930,N_39722);
nor U40530 (N_40530,N_39952,N_39294);
or U40531 (N_40531,N_39422,N_39732);
or U40532 (N_40532,N_39185,N_39035);
xnor U40533 (N_40533,N_39196,N_39746);
and U40534 (N_40534,N_39812,N_39972);
xnor U40535 (N_40535,N_39341,N_39013);
or U40536 (N_40536,N_39194,N_39296);
or U40537 (N_40537,N_39791,N_39489);
nand U40538 (N_40538,N_39300,N_39480);
nand U40539 (N_40539,N_39136,N_39444);
xor U40540 (N_40540,N_39756,N_39977);
xnor U40541 (N_40541,N_39645,N_39739);
xnor U40542 (N_40542,N_39844,N_39943);
nand U40543 (N_40543,N_39725,N_39603);
or U40544 (N_40544,N_39861,N_39390);
nand U40545 (N_40545,N_39119,N_39966);
xor U40546 (N_40546,N_39309,N_39652);
nand U40547 (N_40547,N_39552,N_39385);
or U40548 (N_40548,N_39236,N_39404);
and U40549 (N_40549,N_39044,N_39796);
or U40550 (N_40550,N_39300,N_39802);
xnor U40551 (N_40551,N_39992,N_39397);
xnor U40552 (N_40552,N_39576,N_39261);
nand U40553 (N_40553,N_39474,N_39750);
and U40554 (N_40554,N_39429,N_39887);
xor U40555 (N_40555,N_39422,N_39248);
xnor U40556 (N_40556,N_39206,N_39862);
nand U40557 (N_40557,N_39983,N_39615);
nand U40558 (N_40558,N_39556,N_39526);
and U40559 (N_40559,N_39302,N_39461);
xor U40560 (N_40560,N_39168,N_39272);
or U40561 (N_40561,N_39802,N_39327);
nand U40562 (N_40562,N_39819,N_39812);
nand U40563 (N_40563,N_39018,N_39398);
nand U40564 (N_40564,N_39124,N_39479);
nor U40565 (N_40565,N_39069,N_39198);
nand U40566 (N_40566,N_39743,N_39440);
nor U40567 (N_40567,N_39177,N_39153);
xor U40568 (N_40568,N_39285,N_39241);
or U40569 (N_40569,N_39003,N_39523);
nor U40570 (N_40570,N_39392,N_39294);
or U40571 (N_40571,N_39460,N_39792);
and U40572 (N_40572,N_39165,N_39362);
or U40573 (N_40573,N_39523,N_39290);
nand U40574 (N_40574,N_39167,N_39843);
nand U40575 (N_40575,N_39949,N_39985);
and U40576 (N_40576,N_39357,N_39715);
nor U40577 (N_40577,N_39058,N_39986);
and U40578 (N_40578,N_39065,N_39980);
nand U40579 (N_40579,N_39915,N_39407);
xor U40580 (N_40580,N_39584,N_39726);
xor U40581 (N_40581,N_39925,N_39837);
and U40582 (N_40582,N_39078,N_39806);
and U40583 (N_40583,N_39278,N_39685);
nor U40584 (N_40584,N_39898,N_39877);
nor U40585 (N_40585,N_39296,N_39488);
xor U40586 (N_40586,N_39681,N_39086);
or U40587 (N_40587,N_39076,N_39791);
nor U40588 (N_40588,N_39256,N_39686);
and U40589 (N_40589,N_39388,N_39803);
xnor U40590 (N_40590,N_39243,N_39042);
or U40591 (N_40591,N_39087,N_39908);
or U40592 (N_40592,N_39699,N_39190);
or U40593 (N_40593,N_39632,N_39831);
nor U40594 (N_40594,N_39778,N_39058);
nand U40595 (N_40595,N_39722,N_39062);
nand U40596 (N_40596,N_39032,N_39693);
nand U40597 (N_40597,N_39283,N_39970);
or U40598 (N_40598,N_39360,N_39530);
xnor U40599 (N_40599,N_39459,N_39315);
and U40600 (N_40600,N_39067,N_39969);
nor U40601 (N_40601,N_39295,N_39963);
or U40602 (N_40602,N_39866,N_39543);
nor U40603 (N_40603,N_39969,N_39358);
nand U40604 (N_40604,N_39416,N_39907);
nand U40605 (N_40605,N_39952,N_39151);
or U40606 (N_40606,N_39549,N_39828);
xor U40607 (N_40607,N_39152,N_39765);
nand U40608 (N_40608,N_39369,N_39544);
and U40609 (N_40609,N_39578,N_39092);
nor U40610 (N_40610,N_39439,N_39808);
or U40611 (N_40611,N_39018,N_39089);
or U40612 (N_40612,N_39400,N_39477);
or U40613 (N_40613,N_39189,N_39326);
and U40614 (N_40614,N_39719,N_39523);
xor U40615 (N_40615,N_39991,N_39844);
or U40616 (N_40616,N_39172,N_39482);
nor U40617 (N_40617,N_39961,N_39439);
xor U40618 (N_40618,N_39641,N_39762);
or U40619 (N_40619,N_39130,N_39286);
or U40620 (N_40620,N_39218,N_39529);
nand U40621 (N_40621,N_39072,N_39990);
nand U40622 (N_40622,N_39155,N_39995);
nand U40623 (N_40623,N_39281,N_39451);
or U40624 (N_40624,N_39668,N_39655);
nand U40625 (N_40625,N_39944,N_39773);
nand U40626 (N_40626,N_39640,N_39415);
nand U40627 (N_40627,N_39678,N_39393);
nand U40628 (N_40628,N_39047,N_39594);
and U40629 (N_40629,N_39198,N_39872);
or U40630 (N_40630,N_39192,N_39691);
or U40631 (N_40631,N_39239,N_39779);
nor U40632 (N_40632,N_39323,N_39903);
xor U40633 (N_40633,N_39351,N_39486);
xor U40634 (N_40634,N_39749,N_39001);
or U40635 (N_40635,N_39947,N_39133);
nand U40636 (N_40636,N_39221,N_39657);
xnor U40637 (N_40637,N_39223,N_39167);
nor U40638 (N_40638,N_39212,N_39165);
or U40639 (N_40639,N_39795,N_39817);
nand U40640 (N_40640,N_39153,N_39976);
nand U40641 (N_40641,N_39833,N_39736);
xnor U40642 (N_40642,N_39579,N_39864);
nand U40643 (N_40643,N_39997,N_39383);
and U40644 (N_40644,N_39856,N_39787);
or U40645 (N_40645,N_39534,N_39293);
nor U40646 (N_40646,N_39211,N_39915);
nor U40647 (N_40647,N_39758,N_39274);
nor U40648 (N_40648,N_39120,N_39692);
or U40649 (N_40649,N_39856,N_39022);
xnor U40650 (N_40650,N_39223,N_39946);
or U40651 (N_40651,N_39928,N_39572);
nand U40652 (N_40652,N_39816,N_39264);
xnor U40653 (N_40653,N_39742,N_39648);
nand U40654 (N_40654,N_39855,N_39619);
nand U40655 (N_40655,N_39783,N_39543);
xor U40656 (N_40656,N_39558,N_39565);
and U40657 (N_40657,N_39877,N_39349);
nand U40658 (N_40658,N_39274,N_39680);
or U40659 (N_40659,N_39986,N_39150);
nor U40660 (N_40660,N_39002,N_39412);
and U40661 (N_40661,N_39915,N_39806);
and U40662 (N_40662,N_39818,N_39530);
xnor U40663 (N_40663,N_39395,N_39936);
nor U40664 (N_40664,N_39038,N_39911);
nand U40665 (N_40665,N_39214,N_39435);
xor U40666 (N_40666,N_39931,N_39109);
xnor U40667 (N_40667,N_39592,N_39385);
nand U40668 (N_40668,N_39042,N_39444);
nor U40669 (N_40669,N_39195,N_39660);
nor U40670 (N_40670,N_39402,N_39169);
nand U40671 (N_40671,N_39634,N_39909);
or U40672 (N_40672,N_39411,N_39202);
nand U40673 (N_40673,N_39966,N_39283);
or U40674 (N_40674,N_39017,N_39485);
nor U40675 (N_40675,N_39505,N_39823);
nand U40676 (N_40676,N_39106,N_39801);
xnor U40677 (N_40677,N_39795,N_39935);
xor U40678 (N_40678,N_39930,N_39135);
nand U40679 (N_40679,N_39263,N_39308);
nor U40680 (N_40680,N_39814,N_39996);
xor U40681 (N_40681,N_39781,N_39306);
nor U40682 (N_40682,N_39978,N_39902);
xnor U40683 (N_40683,N_39462,N_39795);
xor U40684 (N_40684,N_39872,N_39028);
xnor U40685 (N_40685,N_39435,N_39502);
and U40686 (N_40686,N_39388,N_39859);
xnor U40687 (N_40687,N_39877,N_39091);
nand U40688 (N_40688,N_39951,N_39098);
xor U40689 (N_40689,N_39772,N_39154);
nand U40690 (N_40690,N_39680,N_39021);
or U40691 (N_40691,N_39631,N_39131);
nor U40692 (N_40692,N_39285,N_39730);
or U40693 (N_40693,N_39745,N_39336);
and U40694 (N_40694,N_39133,N_39252);
nand U40695 (N_40695,N_39602,N_39059);
nor U40696 (N_40696,N_39471,N_39389);
or U40697 (N_40697,N_39011,N_39574);
and U40698 (N_40698,N_39847,N_39930);
nand U40699 (N_40699,N_39143,N_39992);
nor U40700 (N_40700,N_39050,N_39566);
xnor U40701 (N_40701,N_39731,N_39026);
nand U40702 (N_40702,N_39019,N_39316);
or U40703 (N_40703,N_39125,N_39225);
or U40704 (N_40704,N_39873,N_39952);
nor U40705 (N_40705,N_39455,N_39667);
xor U40706 (N_40706,N_39122,N_39604);
and U40707 (N_40707,N_39583,N_39836);
nor U40708 (N_40708,N_39872,N_39860);
or U40709 (N_40709,N_39522,N_39225);
nor U40710 (N_40710,N_39430,N_39146);
nor U40711 (N_40711,N_39590,N_39093);
or U40712 (N_40712,N_39799,N_39360);
or U40713 (N_40713,N_39473,N_39610);
nand U40714 (N_40714,N_39385,N_39520);
nor U40715 (N_40715,N_39430,N_39057);
or U40716 (N_40716,N_39512,N_39619);
xor U40717 (N_40717,N_39579,N_39090);
and U40718 (N_40718,N_39863,N_39868);
xnor U40719 (N_40719,N_39547,N_39913);
and U40720 (N_40720,N_39384,N_39668);
or U40721 (N_40721,N_39034,N_39812);
xor U40722 (N_40722,N_39554,N_39384);
nand U40723 (N_40723,N_39264,N_39083);
nand U40724 (N_40724,N_39685,N_39946);
or U40725 (N_40725,N_39246,N_39840);
nand U40726 (N_40726,N_39454,N_39971);
xnor U40727 (N_40727,N_39961,N_39883);
or U40728 (N_40728,N_39892,N_39647);
nand U40729 (N_40729,N_39336,N_39718);
or U40730 (N_40730,N_39204,N_39930);
and U40731 (N_40731,N_39150,N_39603);
nor U40732 (N_40732,N_39167,N_39601);
xor U40733 (N_40733,N_39838,N_39680);
xor U40734 (N_40734,N_39732,N_39583);
and U40735 (N_40735,N_39524,N_39976);
nor U40736 (N_40736,N_39679,N_39508);
nand U40737 (N_40737,N_39030,N_39874);
nand U40738 (N_40738,N_39482,N_39717);
or U40739 (N_40739,N_39615,N_39517);
and U40740 (N_40740,N_39112,N_39998);
or U40741 (N_40741,N_39805,N_39711);
or U40742 (N_40742,N_39689,N_39909);
xor U40743 (N_40743,N_39399,N_39687);
and U40744 (N_40744,N_39507,N_39071);
xnor U40745 (N_40745,N_39753,N_39437);
and U40746 (N_40746,N_39741,N_39102);
or U40747 (N_40747,N_39982,N_39682);
nand U40748 (N_40748,N_39132,N_39435);
and U40749 (N_40749,N_39476,N_39756);
nand U40750 (N_40750,N_39730,N_39682);
xnor U40751 (N_40751,N_39947,N_39523);
nand U40752 (N_40752,N_39544,N_39349);
xor U40753 (N_40753,N_39774,N_39246);
nand U40754 (N_40754,N_39987,N_39657);
nand U40755 (N_40755,N_39178,N_39339);
nand U40756 (N_40756,N_39014,N_39119);
nor U40757 (N_40757,N_39288,N_39232);
xor U40758 (N_40758,N_39681,N_39784);
and U40759 (N_40759,N_39225,N_39683);
xor U40760 (N_40760,N_39009,N_39680);
or U40761 (N_40761,N_39249,N_39804);
nand U40762 (N_40762,N_39039,N_39293);
and U40763 (N_40763,N_39568,N_39363);
and U40764 (N_40764,N_39874,N_39961);
nor U40765 (N_40765,N_39956,N_39701);
or U40766 (N_40766,N_39853,N_39193);
nor U40767 (N_40767,N_39123,N_39768);
nand U40768 (N_40768,N_39242,N_39360);
or U40769 (N_40769,N_39084,N_39113);
nand U40770 (N_40770,N_39733,N_39870);
nand U40771 (N_40771,N_39283,N_39826);
nor U40772 (N_40772,N_39194,N_39516);
xor U40773 (N_40773,N_39006,N_39355);
nand U40774 (N_40774,N_39924,N_39178);
xor U40775 (N_40775,N_39591,N_39868);
nand U40776 (N_40776,N_39517,N_39909);
xor U40777 (N_40777,N_39939,N_39339);
and U40778 (N_40778,N_39895,N_39415);
nor U40779 (N_40779,N_39794,N_39790);
and U40780 (N_40780,N_39220,N_39335);
xor U40781 (N_40781,N_39690,N_39137);
xor U40782 (N_40782,N_39902,N_39012);
nor U40783 (N_40783,N_39280,N_39094);
and U40784 (N_40784,N_39401,N_39304);
and U40785 (N_40785,N_39938,N_39698);
or U40786 (N_40786,N_39236,N_39739);
xnor U40787 (N_40787,N_39138,N_39942);
nand U40788 (N_40788,N_39831,N_39533);
and U40789 (N_40789,N_39507,N_39805);
nor U40790 (N_40790,N_39805,N_39088);
and U40791 (N_40791,N_39026,N_39366);
or U40792 (N_40792,N_39231,N_39442);
xor U40793 (N_40793,N_39582,N_39474);
and U40794 (N_40794,N_39121,N_39348);
nand U40795 (N_40795,N_39281,N_39562);
or U40796 (N_40796,N_39066,N_39324);
nor U40797 (N_40797,N_39604,N_39322);
or U40798 (N_40798,N_39714,N_39458);
and U40799 (N_40799,N_39935,N_39425);
nor U40800 (N_40800,N_39924,N_39430);
and U40801 (N_40801,N_39653,N_39969);
nand U40802 (N_40802,N_39337,N_39657);
and U40803 (N_40803,N_39246,N_39401);
xor U40804 (N_40804,N_39897,N_39658);
and U40805 (N_40805,N_39144,N_39632);
nand U40806 (N_40806,N_39954,N_39247);
and U40807 (N_40807,N_39197,N_39757);
xnor U40808 (N_40808,N_39628,N_39040);
and U40809 (N_40809,N_39491,N_39790);
or U40810 (N_40810,N_39620,N_39784);
and U40811 (N_40811,N_39883,N_39268);
nand U40812 (N_40812,N_39696,N_39615);
or U40813 (N_40813,N_39782,N_39102);
nand U40814 (N_40814,N_39267,N_39766);
or U40815 (N_40815,N_39154,N_39973);
nor U40816 (N_40816,N_39182,N_39569);
nand U40817 (N_40817,N_39289,N_39167);
xor U40818 (N_40818,N_39076,N_39460);
nor U40819 (N_40819,N_39409,N_39247);
nand U40820 (N_40820,N_39381,N_39382);
or U40821 (N_40821,N_39974,N_39375);
and U40822 (N_40822,N_39961,N_39012);
and U40823 (N_40823,N_39791,N_39807);
and U40824 (N_40824,N_39597,N_39634);
xnor U40825 (N_40825,N_39183,N_39907);
nand U40826 (N_40826,N_39384,N_39129);
or U40827 (N_40827,N_39043,N_39448);
nand U40828 (N_40828,N_39897,N_39470);
and U40829 (N_40829,N_39720,N_39021);
nor U40830 (N_40830,N_39299,N_39585);
nor U40831 (N_40831,N_39466,N_39607);
nand U40832 (N_40832,N_39355,N_39994);
nand U40833 (N_40833,N_39881,N_39629);
and U40834 (N_40834,N_39737,N_39936);
nor U40835 (N_40835,N_39668,N_39564);
or U40836 (N_40836,N_39302,N_39938);
and U40837 (N_40837,N_39916,N_39381);
nand U40838 (N_40838,N_39733,N_39298);
or U40839 (N_40839,N_39151,N_39962);
nor U40840 (N_40840,N_39644,N_39452);
and U40841 (N_40841,N_39084,N_39231);
nor U40842 (N_40842,N_39321,N_39589);
xor U40843 (N_40843,N_39076,N_39308);
nand U40844 (N_40844,N_39408,N_39275);
nor U40845 (N_40845,N_39941,N_39775);
or U40846 (N_40846,N_39214,N_39447);
nand U40847 (N_40847,N_39322,N_39509);
nand U40848 (N_40848,N_39545,N_39048);
nor U40849 (N_40849,N_39349,N_39913);
nand U40850 (N_40850,N_39529,N_39034);
xor U40851 (N_40851,N_39420,N_39844);
nand U40852 (N_40852,N_39433,N_39045);
and U40853 (N_40853,N_39417,N_39968);
and U40854 (N_40854,N_39959,N_39161);
nor U40855 (N_40855,N_39928,N_39181);
nor U40856 (N_40856,N_39599,N_39550);
or U40857 (N_40857,N_39381,N_39271);
xor U40858 (N_40858,N_39760,N_39241);
nand U40859 (N_40859,N_39623,N_39221);
xor U40860 (N_40860,N_39620,N_39036);
nor U40861 (N_40861,N_39888,N_39100);
xnor U40862 (N_40862,N_39768,N_39156);
xor U40863 (N_40863,N_39310,N_39909);
nor U40864 (N_40864,N_39771,N_39104);
and U40865 (N_40865,N_39762,N_39850);
or U40866 (N_40866,N_39217,N_39011);
and U40867 (N_40867,N_39615,N_39948);
nor U40868 (N_40868,N_39468,N_39291);
xor U40869 (N_40869,N_39499,N_39452);
xor U40870 (N_40870,N_39281,N_39868);
and U40871 (N_40871,N_39664,N_39106);
nand U40872 (N_40872,N_39011,N_39635);
nor U40873 (N_40873,N_39903,N_39510);
nor U40874 (N_40874,N_39076,N_39085);
xor U40875 (N_40875,N_39788,N_39658);
nand U40876 (N_40876,N_39289,N_39094);
nor U40877 (N_40877,N_39042,N_39978);
xor U40878 (N_40878,N_39188,N_39746);
nor U40879 (N_40879,N_39228,N_39373);
nor U40880 (N_40880,N_39443,N_39405);
and U40881 (N_40881,N_39507,N_39157);
nor U40882 (N_40882,N_39729,N_39202);
or U40883 (N_40883,N_39837,N_39458);
xnor U40884 (N_40884,N_39504,N_39370);
or U40885 (N_40885,N_39566,N_39005);
xor U40886 (N_40886,N_39954,N_39597);
nor U40887 (N_40887,N_39705,N_39882);
nor U40888 (N_40888,N_39887,N_39098);
nor U40889 (N_40889,N_39988,N_39672);
or U40890 (N_40890,N_39391,N_39745);
xnor U40891 (N_40891,N_39866,N_39953);
and U40892 (N_40892,N_39654,N_39425);
or U40893 (N_40893,N_39614,N_39791);
or U40894 (N_40894,N_39873,N_39160);
nor U40895 (N_40895,N_39887,N_39351);
or U40896 (N_40896,N_39697,N_39650);
nand U40897 (N_40897,N_39702,N_39635);
nor U40898 (N_40898,N_39156,N_39638);
nor U40899 (N_40899,N_39152,N_39914);
and U40900 (N_40900,N_39422,N_39193);
nand U40901 (N_40901,N_39976,N_39961);
and U40902 (N_40902,N_39956,N_39025);
or U40903 (N_40903,N_39099,N_39283);
xnor U40904 (N_40904,N_39577,N_39675);
nor U40905 (N_40905,N_39135,N_39654);
and U40906 (N_40906,N_39469,N_39407);
and U40907 (N_40907,N_39743,N_39304);
nor U40908 (N_40908,N_39356,N_39288);
xor U40909 (N_40909,N_39139,N_39767);
xor U40910 (N_40910,N_39483,N_39152);
nor U40911 (N_40911,N_39724,N_39359);
and U40912 (N_40912,N_39587,N_39901);
nor U40913 (N_40913,N_39553,N_39878);
nor U40914 (N_40914,N_39007,N_39279);
nand U40915 (N_40915,N_39041,N_39763);
xnor U40916 (N_40916,N_39218,N_39524);
and U40917 (N_40917,N_39878,N_39143);
xnor U40918 (N_40918,N_39405,N_39191);
and U40919 (N_40919,N_39357,N_39147);
and U40920 (N_40920,N_39185,N_39037);
xor U40921 (N_40921,N_39343,N_39790);
and U40922 (N_40922,N_39823,N_39220);
or U40923 (N_40923,N_39323,N_39670);
xor U40924 (N_40924,N_39547,N_39410);
and U40925 (N_40925,N_39827,N_39133);
nand U40926 (N_40926,N_39752,N_39812);
or U40927 (N_40927,N_39449,N_39832);
nor U40928 (N_40928,N_39348,N_39784);
nor U40929 (N_40929,N_39162,N_39868);
and U40930 (N_40930,N_39602,N_39476);
nor U40931 (N_40931,N_39996,N_39588);
nand U40932 (N_40932,N_39066,N_39535);
or U40933 (N_40933,N_39080,N_39160);
nand U40934 (N_40934,N_39202,N_39707);
xor U40935 (N_40935,N_39751,N_39670);
nand U40936 (N_40936,N_39286,N_39613);
or U40937 (N_40937,N_39827,N_39173);
or U40938 (N_40938,N_39294,N_39829);
nand U40939 (N_40939,N_39689,N_39753);
and U40940 (N_40940,N_39347,N_39887);
xnor U40941 (N_40941,N_39014,N_39874);
nand U40942 (N_40942,N_39279,N_39581);
and U40943 (N_40943,N_39071,N_39766);
nor U40944 (N_40944,N_39322,N_39309);
xnor U40945 (N_40945,N_39501,N_39397);
nor U40946 (N_40946,N_39442,N_39167);
nor U40947 (N_40947,N_39368,N_39403);
nand U40948 (N_40948,N_39829,N_39675);
nor U40949 (N_40949,N_39609,N_39556);
or U40950 (N_40950,N_39169,N_39599);
or U40951 (N_40951,N_39654,N_39963);
or U40952 (N_40952,N_39175,N_39255);
nor U40953 (N_40953,N_39928,N_39660);
xnor U40954 (N_40954,N_39351,N_39321);
and U40955 (N_40955,N_39664,N_39048);
nor U40956 (N_40956,N_39133,N_39941);
and U40957 (N_40957,N_39626,N_39756);
nor U40958 (N_40958,N_39654,N_39036);
or U40959 (N_40959,N_39743,N_39012);
xor U40960 (N_40960,N_39167,N_39059);
nor U40961 (N_40961,N_39783,N_39664);
xor U40962 (N_40962,N_39175,N_39497);
xor U40963 (N_40963,N_39054,N_39326);
nand U40964 (N_40964,N_39604,N_39697);
and U40965 (N_40965,N_39262,N_39228);
and U40966 (N_40966,N_39300,N_39537);
nand U40967 (N_40967,N_39725,N_39568);
nor U40968 (N_40968,N_39005,N_39478);
or U40969 (N_40969,N_39346,N_39802);
and U40970 (N_40970,N_39578,N_39689);
nand U40971 (N_40971,N_39436,N_39327);
nor U40972 (N_40972,N_39216,N_39015);
and U40973 (N_40973,N_39516,N_39396);
nor U40974 (N_40974,N_39697,N_39370);
or U40975 (N_40975,N_39786,N_39381);
or U40976 (N_40976,N_39936,N_39961);
and U40977 (N_40977,N_39486,N_39439);
xor U40978 (N_40978,N_39463,N_39694);
xnor U40979 (N_40979,N_39606,N_39644);
or U40980 (N_40980,N_39935,N_39021);
nor U40981 (N_40981,N_39268,N_39371);
xor U40982 (N_40982,N_39368,N_39508);
nand U40983 (N_40983,N_39129,N_39161);
and U40984 (N_40984,N_39914,N_39349);
xnor U40985 (N_40985,N_39121,N_39806);
nor U40986 (N_40986,N_39205,N_39864);
or U40987 (N_40987,N_39287,N_39275);
xnor U40988 (N_40988,N_39628,N_39980);
nand U40989 (N_40989,N_39553,N_39699);
nand U40990 (N_40990,N_39218,N_39829);
nor U40991 (N_40991,N_39427,N_39920);
nand U40992 (N_40992,N_39456,N_39336);
or U40993 (N_40993,N_39063,N_39879);
nand U40994 (N_40994,N_39493,N_39791);
nand U40995 (N_40995,N_39424,N_39841);
and U40996 (N_40996,N_39604,N_39577);
nor U40997 (N_40997,N_39116,N_39787);
nor U40998 (N_40998,N_39762,N_39634);
xnor U40999 (N_40999,N_39454,N_39910);
or U41000 (N_41000,N_40697,N_40983);
or U41001 (N_41001,N_40446,N_40521);
and U41002 (N_41002,N_40613,N_40066);
xnor U41003 (N_41003,N_40702,N_40950);
and U41004 (N_41004,N_40688,N_40128);
xnor U41005 (N_41005,N_40631,N_40709);
nand U41006 (N_41006,N_40456,N_40215);
xor U41007 (N_41007,N_40899,N_40912);
nor U41008 (N_41008,N_40682,N_40550);
nand U41009 (N_41009,N_40995,N_40017);
nand U41010 (N_41010,N_40442,N_40825);
nand U41011 (N_41011,N_40587,N_40646);
or U41012 (N_41012,N_40663,N_40167);
and U41013 (N_41013,N_40810,N_40637);
or U41014 (N_41014,N_40137,N_40264);
xor U41015 (N_41015,N_40628,N_40733);
and U41016 (N_41016,N_40778,N_40857);
xor U41017 (N_41017,N_40144,N_40558);
xor U41018 (N_41018,N_40142,N_40900);
or U41019 (N_41019,N_40856,N_40422);
and U41020 (N_41020,N_40951,N_40477);
or U41021 (N_41021,N_40651,N_40716);
and U41022 (N_41022,N_40962,N_40745);
and U41023 (N_41023,N_40584,N_40107);
nand U41024 (N_41024,N_40679,N_40738);
or U41025 (N_41025,N_40618,N_40411);
xnor U41026 (N_41026,N_40540,N_40691);
nand U41027 (N_41027,N_40734,N_40546);
xnor U41028 (N_41028,N_40473,N_40140);
xor U41029 (N_41029,N_40491,N_40576);
and U41030 (N_41030,N_40133,N_40271);
and U41031 (N_41031,N_40827,N_40080);
or U41032 (N_41032,N_40764,N_40112);
nand U41033 (N_41033,N_40092,N_40580);
or U41034 (N_41034,N_40279,N_40018);
nor U41035 (N_41035,N_40314,N_40927);
or U41036 (N_41036,N_40500,N_40627);
nand U41037 (N_41037,N_40875,N_40413);
nand U41038 (N_41038,N_40042,N_40831);
nand U41039 (N_41039,N_40844,N_40743);
and U41040 (N_41040,N_40154,N_40355);
xor U41041 (N_41041,N_40737,N_40447);
or U41042 (N_41042,N_40385,N_40503);
nand U41043 (N_41043,N_40909,N_40259);
or U41044 (N_41044,N_40076,N_40883);
nor U41045 (N_41045,N_40276,N_40242);
and U41046 (N_41046,N_40805,N_40015);
xor U41047 (N_41047,N_40425,N_40678);
nor U41048 (N_41048,N_40484,N_40811);
nor U41049 (N_41049,N_40013,N_40780);
xnor U41050 (N_41050,N_40717,N_40203);
nor U41051 (N_41051,N_40729,N_40589);
nor U41052 (N_41052,N_40056,N_40954);
xnor U41053 (N_41053,N_40171,N_40762);
or U41054 (N_41054,N_40274,N_40190);
nand U41055 (N_41055,N_40519,N_40338);
xor U41056 (N_41056,N_40634,N_40380);
and U41057 (N_41057,N_40339,N_40728);
or U41058 (N_41058,N_40184,N_40861);
or U41059 (N_41059,N_40725,N_40999);
or U41060 (N_41060,N_40181,N_40358);
nor U41061 (N_41061,N_40067,N_40221);
xnor U41062 (N_41062,N_40660,N_40506);
xor U41063 (N_41063,N_40704,N_40784);
xor U41064 (N_41064,N_40465,N_40026);
nor U41065 (N_41065,N_40479,N_40330);
nor U41066 (N_41066,N_40481,N_40043);
or U41067 (N_41067,N_40516,N_40980);
or U41068 (N_41068,N_40489,N_40568);
nor U41069 (N_41069,N_40201,N_40812);
nor U41070 (N_41070,N_40654,N_40785);
and U41071 (N_41071,N_40115,N_40134);
nor U41072 (N_41072,N_40783,N_40829);
or U41073 (N_41073,N_40072,N_40369);
nand U41074 (N_41074,N_40907,N_40886);
or U41075 (N_41075,N_40905,N_40287);
xnor U41076 (N_41076,N_40126,N_40050);
xnor U41077 (N_41077,N_40932,N_40948);
nand U41078 (N_41078,N_40214,N_40735);
nand U41079 (N_41079,N_40700,N_40417);
or U41080 (N_41080,N_40485,N_40236);
nor U41081 (N_41081,N_40731,N_40541);
or U41082 (N_41082,N_40430,N_40750);
and U41083 (N_41083,N_40269,N_40437);
xnor U41084 (N_41084,N_40490,N_40097);
or U41085 (N_41085,N_40022,N_40206);
xnor U41086 (N_41086,N_40979,N_40629);
and U41087 (N_41087,N_40044,N_40977);
xor U41088 (N_41088,N_40048,N_40147);
or U41089 (N_41089,N_40244,N_40781);
nor U41090 (N_41090,N_40333,N_40551);
nor U41091 (N_41091,N_40658,N_40262);
or U41092 (N_41092,N_40397,N_40476);
and U41093 (N_41093,N_40329,N_40098);
or U41094 (N_41094,N_40925,N_40868);
and U41095 (N_41095,N_40429,N_40318);
nor U41096 (N_41096,N_40052,N_40918);
or U41097 (N_41097,N_40528,N_40258);
nand U41098 (N_41098,N_40852,N_40426);
nor U41099 (N_41099,N_40246,N_40790);
xor U41100 (N_41100,N_40690,N_40427);
or U41101 (N_41101,N_40419,N_40913);
and U41102 (N_41102,N_40607,N_40683);
xor U41103 (N_41103,N_40988,N_40420);
nand U41104 (N_41104,N_40590,N_40668);
or U41105 (N_41105,N_40170,N_40599);
or U41106 (N_41106,N_40091,N_40585);
xor U41107 (N_41107,N_40436,N_40758);
or U41108 (N_41108,N_40100,N_40266);
nand U41109 (N_41109,N_40273,N_40055);
nor U41110 (N_41110,N_40798,N_40159);
nand U41111 (N_41111,N_40227,N_40316);
xnor U41112 (N_41112,N_40030,N_40952);
nor U41113 (N_41113,N_40435,N_40803);
xor U41114 (N_41114,N_40994,N_40068);
nor U41115 (N_41115,N_40818,N_40257);
or U41116 (N_41116,N_40806,N_40480);
or U41117 (N_41117,N_40450,N_40351);
or U41118 (N_41118,N_40433,N_40808);
or U41119 (N_41119,N_40632,N_40841);
or U41120 (N_41120,N_40874,N_40768);
and U41121 (N_41121,N_40114,N_40471);
or U41122 (N_41122,N_40928,N_40822);
xor U41123 (N_41123,N_40364,N_40686);
or U41124 (N_41124,N_40915,N_40515);
xnor U41125 (N_41125,N_40574,N_40549);
xor U41126 (N_41126,N_40726,N_40843);
xor U41127 (N_41127,N_40566,N_40647);
nor U41128 (N_41128,N_40514,N_40036);
or U41129 (N_41129,N_40021,N_40347);
and U41130 (N_41130,N_40779,N_40956);
or U41131 (N_41131,N_40586,N_40310);
xnor U41132 (N_41132,N_40081,N_40908);
and U41133 (N_41133,N_40455,N_40940);
and U41134 (N_41134,N_40408,N_40636);
and U41135 (N_41135,N_40964,N_40796);
and U41136 (N_41136,N_40300,N_40366);
and U41137 (N_41137,N_40410,N_40431);
xor U41138 (N_41138,N_40807,N_40641);
nand U41139 (N_41139,N_40315,N_40493);
nor U41140 (N_41140,N_40070,N_40047);
and U41141 (N_41141,N_40020,N_40993);
nand U41142 (N_41142,N_40389,N_40039);
nor U41143 (N_41143,N_40248,N_40148);
nor U41144 (N_41144,N_40760,N_40243);
or U41145 (N_41145,N_40185,N_40602);
xor U41146 (N_41146,N_40205,N_40523);
nand U41147 (N_41147,N_40593,N_40759);
and U41148 (N_41148,N_40207,N_40530);
or U41149 (N_41149,N_40394,N_40062);
or U41150 (N_41150,N_40218,N_40307);
or U41151 (N_41151,N_40898,N_40556);
nand U41152 (N_41152,N_40910,N_40786);
nand U41153 (N_41153,N_40946,N_40612);
nand U41154 (N_41154,N_40958,N_40322);
or U41155 (N_41155,N_40714,N_40040);
or U41156 (N_41156,N_40853,N_40139);
nor U41157 (N_41157,N_40216,N_40579);
nor U41158 (N_41158,N_40101,N_40573);
nand U41159 (N_41159,N_40692,N_40858);
nand U41160 (N_41160,N_40849,N_40687);
nand U41161 (N_41161,N_40792,N_40129);
nor U41162 (N_41162,N_40019,N_40539);
and U41163 (N_41163,N_40024,N_40138);
xnor U41164 (N_41164,N_40461,N_40674);
xor U41165 (N_41165,N_40532,N_40225);
xnor U41166 (N_41166,N_40802,N_40096);
xor U41167 (N_41167,N_40014,N_40336);
or U41168 (N_41168,N_40027,N_40640);
nand U41169 (N_41169,N_40531,N_40563);
or U41170 (N_41170,N_40249,N_40031);
and U41171 (N_41171,N_40238,N_40766);
xnor U41172 (N_41172,N_40010,N_40968);
nand U41173 (N_41173,N_40596,N_40230);
or U41174 (N_41174,N_40226,N_40327);
and U41175 (N_41175,N_40053,N_40362);
xnor U41176 (N_41176,N_40575,N_40495);
nor U41177 (N_41177,N_40606,N_40404);
and U41178 (N_41178,N_40961,N_40669);
nor U41179 (N_41179,N_40189,N_40828);
or U41180 (N_41180,N_40740,N_40942);
nand U41181 (N_41181,N_40769,N_40388);
xnor U41182 (N_41182,N_40502,N_40029);
xor U41183 (N_41183,N_40793,N_40732);
nand U41184 (N_41184,N_40720,N_40835);
xor U41185 (N_41185,N_40833,N_40109);
or U41186 (N_41186,N_40296,N_40901);
nand U41187 (N_41187,N_40071,N_40008);
xor U41188 (N_41188,N_40294,N_40280);
and U41189 (N_41189,N_40125,N_40075);
xnor U41190 (N_41190,N_40188,N_40045);
and U41191 (N_41191,N_40777,N_40971);
nand U41192 (N_41192,N_40673,N_40665);
and U41193 (N_41193,N_40522,N_40923);
and U41194 (N_41194,N_40755,N_40839);
nor U41195 (N_41195,N_40416,N_40392);
or U41196 (N_41196,N_40756,N_40299);
nor U41197 (N_41197,N_40305,N_40545);
or U41198 (N_41198,N_40881,N_40840);
and U41199 (N_41199,N_40387,N_40542);
nor U41200 (N_41200,N_40200,N_40059);
nor U41201 (N_41201,N_40127,N_40559);
nor U41202 (N_41202,N_40082,N_40467);
xor U41203 (N_41203,N_40268,N_40194);
and U41204 (N_41204,N_40464,N_40869);
or U41205 (N_41205,N_40060,N_40867);
nor U41206 (N_41206,N_40535,N_40209);
xor U41207 (N_41207,N_40873,N_40644);
or U41208 (N_41208,N_40567,N_40403);
or U41209 (N_41209,N_40765,N_40588);
and U41210 (N_41210,N_40834,N_40123);
nand U41211 (N_41211,N_40512,N_40161);
xor U41212 (N_41212,N_40944,N_40855);
and U41213 (N_41213,N_40449,N_40459);
nor U41214 (N_41214,N_40228,N_40382);
or U41215 (N_41215,N_40526,N_40415);
nand U41216 (N_41216,N_40984,N_40600);
nor U41217 (N_41217,N_40789,N_40232);
and U41218 (N_41218,N_40313,N_40582);
nand U41219 (N_41219,N_40860,N_40309);
nor U41220 (N_41220,N_40730,N_40821);
nand U41221 (N_41221,N_40155,N_40157);
nand U41222 (N_41222,N_40211,N_40985);
xnor U41223 (N_41223,N_40240,N_40003);
or U41224 (N_41224,N_40847,N_40800);
and U41225 (N_41225,N_40289,N_40360);
xor U41226 (N_41226,N_40564,N_40153);
nand U41227 (N_41227,N_40872,N_40007);
and U41228 (N_41228,N_40707,N_40638);
xnor U41229 (N_41229,N_40694,N_40824);
and U41230 (N_41230,N_40866,N_40974);
nand U41231 (N_41231,N_40850,N_40444);
xnor U41232 (N_41232,N_40405,N_40335);
and U41233 (N_41233,N_40902,N_40213);
and U41234 (N_41234,N_40131,N_40443);
or U41235 (N_41235,N_40746,N_40265);
or U41236 (N_41236,N_40935,N_40933);
xnor U41237 (N_41237,N_40581,N_40604);
or U41238 (N_41238,N_40929,N_40368);
nor U41239 (N_41239,N_40592,N_40605);
xnor U41240 (N_41240,N_40428,N_40619);
or U41241 (N_41241,N_40423,N_40505);
and U41242 (N_41242,N_40281,N_40635);
nand U41243 (N_41243,N_40616,N_40418);
nand U41244 (N_41244,N_40340,N_40311);
xnor U41245 (N_41245,N_40337,N_40513);
xnor U41246 (N_41246,N_40367,N_40421);
and U41247 (N_41247,N_40891,N_40992);
nor U41248 (N_41248,N_40562,N_40290);
and U41249 (N_41249,N_40162,N_40676);
xnor U41250 (N_41250,N_40497,N_40611);
and U41251 (N_41251,N_40180,N_40931);
nor U41252 (N_41252,N_40306,N_40057);
xnor U41253 (N_41253,N_40145,N_40344);
and U41254 (N_41254,N_40684,N_40285);
or U41255 (N_41255,N_40578,N_40813);
and U41256 (N_41256,N_40174,N_40685);
nor U41257 (N_41257,N_40577,N_40488);
or U41258 (N_41258,N_40555,N_40196);
nand U41259 (N_41259,N_40445,N_40179);
and U41260 (N_41260,N_40924,N_40937);
or U41261 (N_41261,N_40199,N_40233);
nand U41262 (N_41262,N_40529,N_40492);
nand U41263 (N_41263,N_40352,N_40851);
or U41264 (N_41264,N_40698,N_40090);
and U41265 (N_41265,N_40987,N_40494);
xor U41266 (N_41266,N_40609,N_40049);
xnor U41267 (N_41267,N_40510,N_40791);
and U41268 (N_41268,N_40565,N_40699);
nor U41269 (N_41269,N_40656,N_40705);
and U41270 (N_41270,N_40160,N_40033);
and U41271 (N_41271,N_40941,N_40859);
xnor U41272 (N_41272,N_40560,N_40630);
or U41273 (N_41273,N_40263,N_40887);
nand U41274 (N_41274,N_40890,N_40106);
xor U41275 (N_41275,N_40152,N_40353);
or U41276 (N_41276,N_40086,N_40038);
and U41277 (N_41277,N_40458,N_40695);
and U41278 (N_41278,N_40595,N_40620);
or U41279 (N_41279,N_40776,N_40538);
xnor U41280 (N_41280,N_40889,N_40292);
nor U41281 (N_41281,N_40012,N_40610);
nor U41282 (N_41282,N_40922,N_40557);
nand U41283 (N_41283,N_40099,N_40965);
xnor U41284 (N_41284,N_40103,N_40659);
nor U41285 (N_41285,N_40703,N_40820);
nor U41286 (N_41286,N_40989,N_40301);
and U41287 (N_41287,N_40986,N_40543);
xnor U41288 (N_41288,N_40649,N_40753);
and U41289 (N_41289,N_40671,N_40251);
xor U41290 (N_41290,N_40711,N_40572);
or U41291 (N_41291,N_40548,N_40888);
and U41292 (N_41292,N_40440,N_40186);
xnor U41293 (N_41293,N_40727,N_40438);
nor U41294 (N_41294,N_40893,N_40848);
or U41295 (N_41295,N_40936,N_40229);
xor U41296 (N_41296,N_40016,N_40009);
nand U41297 (N_41297,N_40087,N_40452);
or U41298 (N_41298,N_40885,N_40371);
nor U41299 (N_41299,N_40970,N_40648);
and U41300 (N_41300,N_40884,N_40302);
nand U41301 (N_41301,N_40058,N_40439);
xor U41302 (N_41302,N_40463,N_40006);
nor U41303 (N_41303,N_40749,N_40104);
nor U41304 (N_41304,N_40414,N_40955);
xor U41305 (N_41305,N_40906,N_40832);
xnor U41306 (N_41306,N_40594,N_40121);
nor U41307 (N_41307,N_40914,N_40220);
and U41308 (N_41308,N_40374,N_40390);
and U41309 (N_41309,N_40094,N_40723);
and U41310 (N_41310,N_40591,N_40838);
and U41311 (N_41311,N_40454,N_40254);
and U41312 (N_41312,N_40373,N_40032);
or U41313 (N_41313,N_40136,N_40025);
nor U41314 (N_41314,N_40880,N_40303);
nand U41315 (N_41315,N_40079,N_40763);
nand U41316 (N_41316,N_40998,N_40041);
or U41317 (N_41317,N_40713,N_40633);
or U41318 (N_41318,N_40391,N_40219);
xnor U41319 (N_41319,N_40846,N_40722);
and U41320 (N_41320,N_40706,N_40298);
xnor U41321 (N_41321,N_40799,N_40308);
and U41322 (N_41322,N_40751,N_40583);
xnor U41323 (N_41323,N_40282,N_40973);
or U41324 (N_41324,N_40639,N_40653);
nor U41325 (N_41325,N_40401,N_40972);
or U41326 (N_41326,N_40356,N_40754);
xor U41327 (N_41327,N_40854,N_40934);
nand U41328 (N_41328,N_40239,N_40865);
and U41329 (N_41329,N_40177,N_40409);
nand U41330 (N_41330,N_40689,N_40113);
nand U41331 (N_41331,N_40377,N_40158);
xor U41332 (N_41332,N_40534,N_40460);
nand U41333 (N_41333,N_40911,N_40224);
xnor U41334 (N_41334,N_40132,N_40680);
xor U41335 (N_41335,N_40393,N_40278);
nor U41336 (N_41336,N_40349,N_40664);
nor U41337 (N_41337,N_40370,N_40192);
nand U41338 (N_41338,N_40553,N_40774);
nor U41339 (N_41339,N_40005,N_40354);
xor U41340 (N_41340,N_40645,N_40151);
xor U41341 (N_41341,N_40508,N_40615);
nand U41342 (N_41342,N_40172,N_40943);
nor U41343 (N_41343,N_40361,N_40363);
nor U41344 (N_41344,N_40741,N_40085);
and U41345 (N_41345,N_40498,N_40163);
nand U41346 (N_41346,N_40527,N_40434);
nor U41347 (N_41347,N_40939,N_40073);
and U41348 (N_41348,N_40814,N_40320);
nand U41349 (N_41349,N_40149,N_40701);
xnor U41350 (N_41350,N_40001,N_40501);
or U41351 (N_41351,N_40621,N_40675);
and U41352 (N_41352,N_40197,N_40662);
nand U41353 (N_41353,N_40323,N_40626);
or U41354 (N_41354,N_40569,N_40982);
nor U41355 (N_41355,N_40375,N_40864);
nor U41356 (N_41356,N_40571,N_40381);
or U41357 (N_41357,N_40625,N_40871);
nor U41358 (N_41358,N_40178,N_40379);
nor U41359 (N_41359,N_40350,N_40108);
or U41360 (N_41360,N_40334,N_40063);
xnor U41361 (N_41361,N_40836,N_40552);
and U41362 (N_41362,N_40202,N_40817);
nand U41363 (N_41363,N_40074,N_40078);
nand U41364 (N_41364,N_40195,N_40255);
and U41365 (N_41365,N_40483,N_40386);
and U41366 (N_41366,N_40823,N_40191);
and U41367 (N_41367,N_40617,N_40870);
or U41368 (N_41368,N_40231,N_40696);
and U41369 (N_41369,N_40953,N_40742);
nand U41370 (N_41370,N_40837,N_40261);
nand U41371 (N_41371,N_40949,N_40116);
and U41372 (N_41372,N_40400,N_40348);
xnor U41373 (N_41373,N_40325,N_40173);
and U41374 (N_41374,N_40921,N_40457);
and U41375 (N_41375,N_40920,N_40093);
or U41376 (N_41376,N_40710,N_40903);
nor U41377 (N_41377,N_40882,N_40667);
or U41378 (N_41378,N_40034,N_40118);
nand U41379 (N_41379,N_40441,N_40084);
or U41380 (N_41380,N_40117,N_40156);
nor U41381 (N_41381,N_40372,N_40520);
xor U41382 (N_41382,N_40150,N_40395);
and U41383 (N_41383,N_40959,N_40424);
xor U41384 (N_41384,N_40623,N_40288);
nor U41385 (N_41385,N_40250,N_40365);
nand U41386 (N_41386,N_40065,N_40878);
xnor U41387 (N_41387,N_40297,N_40319);
nor U41388 (N_41388,N_40996,N_40130);
and U41389 (N_41389,N_40462,N_40960);
nor U41390 (N_41390,N_40917,N_40896);
nand U41391 (N_41391,N_40895,N_40088);
nand U41392 (N_41392,N_40782,N_40002);
and U41393 (N_41393,N_40622,N_40198);
and U41394 (N_41394,N_40331,N_40210);
or U41395 (N_41395,N_40991,N_40715);
xnor U41396 (N_41396,N_40642,N_40432);
nand U41397 (N_41397,N_40102,N_40744);
or U41398 (N_41398,N_40222,N_40978);
nor U41399 (N_41399,N_40343,N_40772);
nor U41400 (N_41400,N_40023,N_40357);
and U41401 (N_41401,N_40143,N_40892);
xor U41402 (N_41402,N_40451,N_40724);
or U41403 (N_41403,N_40518,N_40721);
or U41404 (N_41404,N_40345,N_40894);
nor U41405 (N_41405,N_40816,N_40603);
or U41406 (N_41406,N_40862,N_40469);
xor U41407 (N_41407,N_40967,N_40509);
nor U41408 (N_41408,N_40051,N_40164);
or U41409 (N_41409,N_40655,N_40842);
nand U41410 (N_41410,N_40474,N_40146);
or U41411 (N_41411,N_40904,N_40283);
nand U41412 (N_41412,N_40597,N_40234);
or U41413 (N_41413,N_40326,N_40801);
xnor U41414 (N_41414,N_40761,N_40412);
and U41415 (N_41415,N_40035,N_40277);
or U41416 (N_41416,N_40719,N_40247);
and U41417 (N_41417,N_40757,N_40879);
and U41418 (N_41418,N_40511,N_40826);
nor U41419 (N_41419,N_40000,N_40332);
xnor U41420 (N_41420,N_40346,N_40845);
or U41421 (N_41421,N_40083,N_40773);
nor U41422 (N_41422,N_40876,N_40975);
nor U41423 (N_41423,N_40997,N_40863);
or U41424 (N_41424,N_40235,N_40804);
xor U41425 (N_41425,N_40770,N_40122);
nand U41426 (N_41426,N_40321,N_40245);
or U41427 (N_41427,N_40448,N_40598);
nor U41428 (N_41428,N_40524,N_40187);
or U41429 (N_41429,N_40681,N_40624);
nor U41430 (N_41430,N_40947,N_40237);
and U41431 (N_41431,N_40341,N_40795);
and U41432 (N_41432,N_40324,N_40208);
nor U41433 (N_41433,N_40957,N_40295);
nand U41434 (N_41434,N_40175,N_40570);
or U41435 (N_41435,N_40286,N_40767);
or U41436 (N_41436,N_40135,N_40794);
nand U41437 (N_41437,N_40089,N_40141);
xor U41438 (N_41438,N_40252,N_40124);
nor U41439 (N_41439,N_40614,N_40544);
and U41440 (N_41440,N_40652,N_40809);
xor U41441 (N_41441,N_40919,N_40657);
and U41442 (N_41442,N_40342,N_40926);
nor U41443 (N_41443,N_40110,N_40253);
nor U41444 (N_41444,N_40736,N_40396);
or U41445 (N_41445,N_40478,N_40468);
xnor U41446 (N_41446,N_40650,N_40775);
xnor U41447 (N_41447,N_40788,N_40317);
nand U41448 (N_41448,N_40990,N_40399);
xor U41449 (N_41449,N_40470,N_40739);
or U41450 (N_41450,N_40976,N_40475);
xnor U41451 (N_41451,N_40095,N_40963);
nand U41452 (N_41452,N_40407,N_40815);
xor U41453 (N_41453,N_40359,N_40028);
and U41454 (N_41454,N_40554,N_40169);
xnor U41455 (N_41455,N_40672,N_40666);
and U41456 (N_41456,N_40517,N_40830);
xnor U41457 (N_41457,N_40069,N_40312);
xnor U41458 (N_41458,N_40119,N_40561);
or U41459 (N_41459,N_40077,N_40176);
xnor U41460 (N_41460,N_40270,N_40547);
nand U41461 (N_41461,N_40111,N_40378);
xor U41462 (N_41462,N_40966,N_40748);
nor U41463 (N_41463,N_40752,N_40384);
nor U41464 (N_41464,N_40453,N_40166);
nor U41465 (N_41465,N_40677,N_40267);
and U41466 (N_41466,N_40661,N_40165);
and U41467 (N_41467,N_40718,N_40376);
or U41468 (N_41468,N_40275,N_40693);
nand U41469 (N_41469,N_40402,N_40291);
nor U41470 (N_41470,N_40537,N_40284);
nor U41471 (N_41471,N_40241,N_40223);
nand U41472 (N_41472,N_40193,N_40797);
and U41473 (N_41473,N_40643,N_40487);
nor U41474 (N_41474,N_40486,N_40819);
nor U41475 (N_41475,N_40217,N_40256);
or U41476 (N_41476,N_40533,N_40383);
xnor U41477 (N_41477,N_40601,N_40504);
nand U41478 (N_41478,N_40046,N_40272);
and U41479 (N_41479,N_40981,N_40938);
nor U41480 (N_41480,N_40182,N_40398);
nor U41481 (N_41481,N_40499,N_40293);
nor U41482 (N_41482,N_40712,N_40771);
and U41483 (N_41483,N_40120,N_40536);
nor U41484 (N_41484,N_40969,N_40168);
nand U41485 (N_41485,N_40496,N_40930);
or U41486 (N_41486,N_40260,N_40945);
nand U41487 (N_41487,N_40304,N_40916);
xor U41488 (N_41488,N_40037,N_40406);
or U41489 (N_41489,N_40507,N_40064);
xnor U41490 (N_41490,N_40670,N_40204);
nand U41491 (N_41491,N_40105,N_40054);
xor U41492 (N_41492,N_40608,N_40328);
xnor U41493 (N_41493,N_40472,N_40525);
or U41494 (N_41494,N_40897,N_40212);
xor U41495 (N_41495,N_40708,N_40466);
nor U41496 (N_41496,N_40061,N_40011);
and U41497 (N_41497,N_40482,N_40183);
and U41498 (N_41498,N_40004,N_40877);
nand U41499 (N_41499,N_40787,N_40747);
xor U41500 (N_41500,N_40047,N_40019);
or U41501 (N_41501,N_40165,N_40925);
nor U41502 (N_41502,N_40643,N_40960);
nand U41503 (N_41503,N_40269,N_40349);
nand U41504 (N_41504,N_40589,N_40531);
nand U41505 (N_41505,N_40814,N_40976);
and U41506 (N_41506,N_40300,N_40176);
and U41507 (N_41507,N_40836,N_40986);
nand U41508 (N_41508,N_40372,N_40363);
and U41509 (N_41509,N_40941,N_40803);
or U41510 (N_41510,N_40957,N_40218);
and U41511 (N_41511,N_40841,N_40169);
and U41512 (N_41512,N_40460,N_40767);
xor U41513 (N_41513,N_40067,N_40468);
nor U41514 (N_41514,N_40095,N_40115);
nor U41515 (N_41515,N_40785,N_40917);
xnor U41516 (N_41516,N_40638,N_40343);
and U41517 (N_41517,N_40863,N_40816);
nand U41518 (N_41518,N_40482,N_40702);
or U41519 (N_41519,N_40753,N_40775);
or U41520 (N_41520,N_40959,N_40065);
or U41521 (N_41521,N_40875,N_40521);
nand U41522 (N_41522,N_40573,N_40931);
nand U41523 (N_41523,N_40259,N_40903);
xnor U41524 (N_41524,N_40618,N_40661);
and U41525 (N_41525,N_40178,N_40846);
or U41526 (N_41526,N_40482,N_40923);
xnor U41527 (N_41527,N_40817,N_40874);
nand U41528 (N_41528,N_40283,N_40296);
or U41529 (N_41529,N_40578,N_40043);
nand U41530 (N_41530,N_40326,N_40901);
or U41531 (N_41531,N_40879,N_40261);
and U41532 (N_41532,N_40274,N_40428);
xnor U41533 (N_41533,N_40987,N_40382);
and U41534 (N_41534,N_40574,N_40324);
nand U41535 (N_41535,N_40075,N_40354);
and U41536 (N_41536,N_40589,N_40137);
or U41537 (N_41537,N_40505,N_40128);
nand U41538 (N_41538,N_40580,N_40188);
and U41539 (N_41539,N_40969,N_40028);
or U41540 (N_41540,N_40634,N_40413);
nand U41541 (N_41541,N_40044,N_40981);
nor U41542 (N_41542,N_40373,N_40243);
nor U41543 (N_41543,N_40617,N_40817);
or U41544 (N_41544,N_40312,N_40019);
xnor U41545 (N_41545,N_40028,N_40705);
xnor U41546 (N_41546,N_40842,N_40460);
nor U41547 (N_41547,N_40828,N_40982);
nand U41548 (N_41548,N_40964,N_40974);
nand U41549 (N_41549,N_40741,N_40998);
xnor U41550 (N_41550,N_40295,N_40176);
or U41551 (N_41551,N_40467,N_40803);
xor U41552 (N_41552,N_40696,N_40397);
xor U41553 (N_41553,N_40697,N_40286);
or U41554 (N_41554,N_40928,N_40610);
xor U41555 (N_41555,N_40516,N_40275);
and U41556 (N_41556,N_40677,N_40681);
and U41557 (N_41557,N_40026,N_40496);
and U41558 (N_41558,N_40874,N_40452);
and U41559 (N_41559,N_40391,N_40275);
nor U41560 (N_41560,N_40345,N_40348);
nor U41561 (N_41561,N_40404,N_40971);
nand U41562 (N_41562,N_40917,N_40004);
or U41563 (N_41563,N_40635,N_40518);
xnor U41564 (N_41564,N_40182,N_40121);
nand U41565 (N_41565,N_40594,N_40803);
xnor U41566 (N_41566,N_40359,N_40801);
nand U41567 (N_41567,N_40936,N_40118);
and U41568 (N_41568,N_40616,N_40765);
xnor U41569 (N_41569,N_40781,N_40932);
nand U41570 (N_41570,N_40772,N_40280);
nor U41571 (N_41571,N_40326,N_40401);
nor U41572 (N_41572,N_40816,N_40736);
xnor U41573 (N_41573,N_40213,N_40868);
xor U41574 (N_41574,N_40649,N_40916);
and U41575 (N_41575,N_40541,N_40084);
and U41576 (N_41576,N_40804,N_40785);
nor U41577 (N_41577,N_40825,N_40910);
and U41578 (N_41578,N_40657,N_40348);
and U41579 (N_41579,N_40156,N_40679);
xnor U41580 (N_41580,N_40866,N_40788);
and U41581 (N_41581,N_40643,N_40099);
xor U41582 (N_41582,N_40077,N_40902);
or U41583 (N_41583,N_40349,N_40711);
nand U41584 (N_41584,N_40605,N_40677);
xnor U41585 (N_41585,N_40243,N_40941);
nand U41586 (N_41586,N_40018,N_40334);
nor U41587 (N_41587,N_40632,N_40736);
xor U41588 (N_41588,N_40627,N_40463);
nand U41589 (N_41589,N_40731,N_40490);
xnor U41590 (N_41590,N_40787,N_40185);
or U41591 (N_41591,N_40219,N_40309);
xnor U41592 (N_41592,N_40850,N_40989);
or U41593 (N_41593,N_40719,N_40793);
nor U41594 (N_41594,N_40529,N_40272);
nand U41595 (N_41595,N_40716,N_40842);
nand U41596 (N_41596,N_40936,N_40356);
and U41597 (N_41597,N_40079,N_40378);
nand U41598 (N_41598,N_40238,N_40704);
and U41599 (N_41599,N_40076,N_40080);
xnor U41600 (N_41600,N_40066,N_40591);
nand U41601 (N_41601,N_40708,N_40225);
and U41602 (N_41602,N_40278,N_40014);
nor U41603 (N_41603,N_40742,N_40432);
nor U41604 (N_41604,N_40203,N_40109);
xnor U41605 (N_41605,N_40823,N_40737);
xor U41606 (N_41606,N_40683,N_40061);
nand U41607 (N_41607,N_40365,N_40916);
and U41608 (N_41608,N_40244,N_40895);
and U41609 (N_41609,N_40966,N_40167);
or U41610 (N_41610,N_40293,N_40165);
and U41611 (N_41611,N_40985,N_40990);
or U41612 (N_41612,N_40160,N_40657);
and U41613 (N_41613,N_40118,N_40532);
nand U41614 (N_41614,N_40771,N_40181);
nor U41615 (N_41615,N_40255,N_40845);
nor U41616 (N_41616,N_40489,N_40642);
nand U41617 (N_41617,N_40702,N_40657);
xnor U41618 (N_41618,N_40738,N_40412);
nand U41619 (N_41619,N_40179,N_40430);
xnor U41620 (N_41620,N_40887,N_40072);
and U41621 (N_41621,N_40527,N_40862);
nor U41622 (N_41622,N_40863,N_40973);
or U41623 (N_41623,N_40933,N_40938);
nor U41624 (N_41624,N_40233,N_40290);
xnor U41625 (N_41625,N_40604,N_40511);
or U41626 (N_41626,N_40465,N_40908);
and U41627 (N_41627,N_40890,N_40657);
nor U41628 (N_41628,N_40115,N_40255);
nor U41629 (N_41629,N_40645,N_40177);
nor U41630 (N_41630,N_40635,N_40222);
nand U41631 (N_41631,N_40791,N_40292);
and U41632 (N_41632,N_40568,N_40773);
nand U41633 (N_41633,N_40357,N_40430);
nor U41634 (N_41634,N_40980,N_40104);
xor U41635 (N_41635,N_40919,N_40644);
or U41636 (N_41636,N_40229,N_40233);
nor U41637 (N_41637,N_40779,N_40896);
nand U41638 (N_41638,N_40235,N_40770);
xor U41639 (N_41639,N_40171,N_40519);
xor U41640 (N_41640,N_40359,N_40138);
xnor U41641 (N_41641,N_40127,N_40721);
nor U41642 (N_41642,N_40166,N_40097);
xor U41643 (N_41643,N_40236,N_40262);
nand U41644 (N_41644,N_40473,N_40728);
nand U41645 (N_41645,N_40969,N_40414);
nor U41646 (N_41646,N_40635,N_40474);
and U41647 (N_41647,N_40053,N_40852);
nand U41648 (N_41648,N_40418,N_40854);
xor U41649 (N_41649,N_40332,N_40817);
nor U41650 (N_41650,N_40003,N_40314);
xnor U41651 (N_41651,N_40894,N_40984);
xnor U41652 (N_41652,N_40829,N_40533);
nor U41653 (N_41653,N_40333,N_40720);
xnor U41654 (N_41654,N_40060,N_40795);
nor U41655 (N_41655,N_40613,N_40050);
and U41656 (N_41656,N_40871,N_40132);
xnor U41657 (N_41657,N_40035,N_40310);
and U41658 (N_41658,N_40107,N_40185);
and U41659 (N_41659,N_40687,N_40147);
xor U41660 (N_41660,N_40362,N_40347);
and U41661 (N_41661,N_40410,N_40813);
xnor U41662 (N_41662,N_40482,N_40839);
and U41663 (N_41663,N_40797,N_40590);
xnor U41664 (N_41664,N_40014,N_40121);
nor U41665 (N_41665,N_40978,N_40498);
nor U41666 (N_41666,N_40862,N_40765);
or U41667 (N_41667,N_40786,N_40224);
and U41668 (N_41668,N_40998,N_40521);
and U41669 (N_41669,N_40877,N_40455);
xnor U41670 (N_41670,N_40652,N_40517);
nor U41671 (N_41671,N_40651,N_40206);
and U41672 (N_41672,N_40015,N_40758);
and U41673 (N_41673,N_40579,N_40854);
or U41674 (N_41674,N_40694,N_40866);
nor U41675 (N_41675,N_40984,N_40276);
xnor U41676 (N_41676,N_40493,N_40580);
or U41677 (N_41677,N_40541,N_40930);
or U41678 (N_41678,N_40314,N_40834);
nor U41679 (N_41679,N_40583,N_40300);
nand U41680 (N_41680,N_40169,N_40970);
or U41681 (N_41681,N_40644,N_40288);
and U41682 (N_41682,N_40276,N_40662);
nor U41683 (N_41683,N_40899,N_40772);
nand U41684 (N_41684,N_40490,N_40379);
xor U41685 (N_41685,N_40430,N_40936);
nor U41686 (N_41686,N_40747,N_40749);
xor U41687 (N_41687,N_40916,N_40002);
xnor U41688 (N_41688,N_40548,N_40604);
xor U41689 (N_41689,N_40642,N_40987);
nand U41690 (N_41690,N_40910,N_40199);
and U41691 (N_41691,N_40206,N_40605);
xnor U41692 (N_41692,N_40433,N_40159);
nand U41693 (N_41693,N_40212,N_40703);
nand U41694 (N_41694,N_40332,N_40517);
nor U41695 (N_41695,N_40858,N_40125);
and U41696 (N_41696,N_40078,N_40919);
and U41697 (N_41697,N_40197,N_40328);
and U41698 (N_41698,N_40421,N_40002);
xor U41699 (N_41699,N_40639,N_40126);
or U41700 (N_41700,N_40610,N_40629);
nand U41701 (N_41701,N_40711,N_40382);
nand U41702 (N_41702,N_40155,N_40410);
nand U41703 (N_41703,N_40119,N_40464);
or U41704 (N_41704,N_40136,N_40089);
nand U41705 (N_41705,N_40580,N_40627);
and U41706 (N_41706,N_40405,N_40923);
and U41707 (N_41707,N_40664,N_40243);
and U41708 (N_41708,N_40064,N_40019);
and U41709 (N_41709,N_40666,N_40651);
nor U41710 (N_41710,N_40840,N_40210);
nor U41711 (N_41711,N_40038,N_40258);
nor U41712 (N_41712,N_40581,N_40821);
or U41713 (N_41713,N_40154,N_40985);
or U41714 (N_41714,N_40837,N_40329);
nor U41715 (N_41715,N_40046,N_40289);
or U41716 (N_41716,N_40979,N_40886);
and U41717 (N_41717,N_40163,N_40765);
and U41718 (N_41718,N_40369,N_40150);
xor U41719 (N_41719,N_40009,N_40322);
nand U41720 (N_41720,N_40817,N_40840);
nor U41721 (N_41721,N_40321,N_40859);
or U41722 (N_41722,N_40126,N_40356);
nor U41723 (N_41723,N_40530,N_40625);
or U41724 (N_41724,N_40892,N_40860);
and U41725 (N_41725,N_40452,N_40909);
or U41726 (N_41726,N_40431,N_40549);
nand U41727 (N_41727,N_40695,N_40829);
xor U41728 (N_41728,N_40067,N_40307);
xnor U41729 (N_41729,N_40921,N_40017);
or U41730 (N_41730,N_40679,N_40282);
nand U41731 (N_41731,N_40107,N_40659);
or U41732 (N_41732,N_40172,N_40246);
xnor U41733 (N_41733,N_40033,N_40144);
xnor U41734 (N_41734,N_40953,N_40949);
nor U41735 (N_41735,N_40903,N_40035);
or U41736 (N_41736,N_40609,N_40735);
nor U41737 (N_41737,N_40494,N_40938);
xnor U41738 (N_41738,N_40474,N_40637);
xnor U41739 (N_41739,N_40377,N_40865);
and U41740 (N_41740,N_40755,N_40359);
nor U41741 (N_41741,N_40073,N_40506);
xnor U41742 (N_41742,N_40240,N_40579);
nor U41743 (N_41743,N_40066,N_40828);
nor U41744 (N_41744,N_40226,N_40181);
or U41745 (N_41745,N_40083,N_40560);
nor U41746 (N_41746,N_40478,N_40187);
or U41747 (N_41747,N_40294,N_40288);
and U41748 (N_41748,N_40683,N_40570);
or U41749 (N_41749,N_40685,N_40893);
xnor U41750 (N_41750,N_40127,N_40881);
nand U41751 (N_41751,N_40681,N_40353);
nand U41752 (N_41752,N_40930,N_40583);
nand U41753 (N_41753,N_40903,N_40270);
and U41754 (N_41754,N_40292,N_40259);
nand U41755 (N_41755,N_40512,N_40081);
nand U41756 (N_41756,N_40471,N_40466);
and U41757 (N_41757,N_40687,N_40222);
nand U41758 (N_41758,N_40808,N_40698);
or U41759 (N_41759,N_40235,N_40428);
nand U41760 (N_41760,N_40815,N_40470);
nand U41761 (N_41761,N_40249,N_40323);
xnor U41762 (N_41762,N_40754,N_40950);
or U41763 (N_41763,N_40014,N_40805);
and U41764 (N_41764,N_40482,N_40738);
and U41765 (N_41765,N_40669,N_40728);
and U41766 (N_41766,N_40481,N_40253);
or U41767 (N_41767,N_40349,N_40530);
or U41768 (N_41768,N_40801,N_40410);
and U41769 (N_41769,N_40232,N_40967);
and U41770 (N_41770,N_40646,N_40826);
nor U41771 (N_41771,N_40366,N_40119);
nand U41772 (N_41772,N_40790,N_40508);
and U41773 (N_41773,N_40262,N_40025);
xnor U41774 (N_41774,N_40618,N_40419);
nor U41775 (N_41775,N_40675,N_40446);
and U41776 (N_41776,N_40195,N_40858);
nand U41777 (N_41777,N_40129,N_40886);
nand U41778 (N_41778,N_40505,N_40727);
and U41779 (N_41779,N_40725,N_40514);
xnor U41780 (N_41780,N_40211,N_40297);
or U41781 (N_41781,N_40373,N_40604);
nand U41782 (N_41782,N_40384,N_40669);
or U41783 (N_41783,N_40637,N_40616);
nand U41784 (N_41784,N_40909,N_40762);
nor U41785 (N_41785,N_40790,N_40985);
nor U41786 (N_41786,N_40105,N_40418);
or U41787 (N_41787,N_40118,N_40605);
xnor U41788 (N_41788,N_40304,N_40058);
or U41789 (N_41789,N_40497,N_40507);
nor U41790 (N_41790,N_40928,N_40870);
nor U41791 (N_41791,N_40186,N_40398);
nor U41792 (N_41792,N_40230,N_40018);
nand U41793 (N_41793,N_40465,N_40661);
nand U41794 (N_41794,N_40339,N_40527);
nand U41795 (N_41795,N_40781,N_40114);
and U41796 (N_41796,N_40934,N_40404);
nand U41797 (N_41797,N_40531,N_40805);
nand U41798 (N_41798,N_40941,N_40248);
nor U41799 (N_41799,N_40394,N_40032);
nor U41800 (N_41800,N_40966,N_40636);
xor U41801 (N_41801,N_40986,N_40936);
xnor U41802 (N_41802,N_40145,N_40768);
xnor U41803 (N_41803,N_40563,N_40017);
nor U41804 (N_41804,N_40081,N_40719);
nor U41805 (N_41805,N_40958,N_40950);
xnor U41806 (N_41806,N_40853,N_40518);
nor U41807 (N_41807,N_40176,N_40059);
nand U41808 (N_41808,N_40887,N_40033);
or U41809 (N_41809,N_40230,N_40937);
or U41810 (N_41810,N_40237,N_40903);
nor U41811 (N_41811,N_40294,N_40960);
and U41812 (N_41812,N_40930,N_40080);
and U41813 (N_41813,N_40397,N_40042);
or U41814 (N_41814,N_40899,N_40576);
and U41815 (N_41815,N_40176,N_40204);
nor U41816 (N_41816,N_40432,N_40744);
nor U41817 (N_41817,N_40876,N_40473);
or U41818 (N_41818,N_40871,N_40525);
nor U41819 (N_41819,N_40806,N_40571);
nor U41820 (N_41820,N_40813,N_40716);
nand U41821 (N_41821,N_40380,N_40089);
nor U41822 (N_41822,N_40402,N_40289);
or U41823 (N_41823,N_40398,N_40057);
and U41824 (N_41824,N_40916,N_40021);
nor U41825 (N_41825,N_40188,N_40455);
and U41826 (N_41826,N_40775,N_40584);
xnor U41827 (N_41827,N_40129,N_40375);
nor U41828 (N_41828,N_40371,N_40882);
or U41829 (N_41829,N_40975,N_40138);
nand U41830 (N_41830,N_40091,N_40376);
nand U41831 (N_41831,N_40077,N_40778);
nor U41832 (N_41832,N_40708,N_40998);
and U41833 (N_41833,N_40131,N_40953);
nand U41834 (N_41834,N_40505,N_40199);
xor U41835 (N_41835,N_40551,N_40498);
or U41836 (N_41836,N_40673,N_40617);
and U41837 (N_41837,N_40121,N_40361);
and U41838 (N_41838,N_40342,N_40507);
or U41839 (N_41839,N_40628,N_40624);
or U41840 (N_41840,N_40417,N_40739);
nor U41841 (N_41841,N_40116,N_40576);
nor U41842 (N_41842,N_40863,N_40937);
and U41843 (N_41843,N_40836,N_40985);
nor U41844 (N_41844,N_40021,N_40868);
nor U41845 (N_41845,N_40980,N_40223);
or U41846 (N_41846,N_40377,N_40927);
or U41847 (N_41847,N_40708,N_40773);
nor U41848 (N_41848,N_40723,N_40647);
xnor U41849 (N_41849,N_40106,N_40148);
nor U41850 (N_41850,N_40427,N_40466);
xnor U41851 (N_41851,N_40467,N_40220);
xnor U41852 (N_41852,N_40591,N_40582);
nand U41853 (N_41853,N_40448,N_40149);
or U41854 (N_41854,N_40161,N_40755);
and U41855 (N_41855,N_40047,N_40961);
or U41856 (N_41856,N_40664,N_40630);
nand U41857 (N_41857,N_40861,N_40269);
nor U41858 (N_41858,N_40798,N_40097);
xor U41859 (N_41859,N_40142,N_40893);
nand U41860 (N_41860,N_40960,N_40154);
nand U41861 (N_41861,N_40393,N_40559);
xnor U41862 (N_41862,N_40831,N_40298);
xnor U41863 (N_41863,N_40356,N_40167);
nand U41864 (N_41864,N_40481,N_40335);
xnor U41865 (N_41865,N_40921,N_40117);
or U41866 (N_41866,N_40760,N_40412);
xor U41867 (N_41867,N_40550,N_40119);
nor U41868 (N_41868,N_40436,N_40201);
xnor U41869 (N_41869,N_40272,N_40877);
xnor U41870 (N_41870,N_40708,N_40925);
xor U41871 (N_41871,N_40241,N_40067);
nor U41872 (N_41872,N_40679,N_40302);
or U41873 (N_41873,N_40670,N_40328);
or U41874 (N_41874,N_40590,N_40160);
or U41875 (N_41875,N_40987,N_40897);
and U41876 (N_41876,N_40128,N_40564);
and U41877 (N_41877,N_40584,N_40191);
nor U41878 (N_41878,N_40096,N_40924);
or U41879 (N_41879,N_40039,N_40047);
or U41880 (N_41880,N_40892,N_40568);
or U41881 (N_41881,N_40110,N_40274);
xor U41882 (N_41882,N_40806,N_40509);
nand U41883 (N_41883,N_40677,N_40649);
nand U41884 (N_41884,N_40521,N_40530);
xnor U41885 (N_41885,N_40772,N_40878);
or U41886 (N_41886,N_40208,N_40907);
nand U41887 (N_41887,N_40276,N_40632);
xnor U41888 (N_41888,N_40239,N_40958);
or U41889 (N_41889,N_40551,N_40645);
and U41890 (N_41890,N_40107,N_40904);
nor U41891 (N_41891,N_40220,N_40254);
or U41892 (N_41892,N_40257,N_40517);
xor U41893 (N_41893,N_40517,N_40968);
nand U41894 (N_41894,N_40505,N_40427);
nand U41895 (N_41895,N_40396,N_40713);
nand U41896 (N_41896,N_40806,N_40595);
nand U41897 (N_41897,N_40646,N_40018);
nor U41898 (N_41898,N_40695,N_40728);
and U41899 (N_41899,N_40866,N_40875);
xor U41900 (N_41900,N_40212,N_40091);
or U41901 (N_41901,N_40175,N_40197);
nor U41902 (N_41902,N_40259,N_40067);
or U41903 (N_41903,N_40970,N_40692);
xnor U41904 (N_41904,N_40567,N_40796);
and U41905 (N_41905,N_40937,N_40343);
xnor U41906 (N_41906,N_40382,N_40009);
nand U41907 (N_41907,N_40703,N_40320);
nand U41908 (N_41908,N_40847,N_40572);
and U41909 (N_41909,N_40283,N_40751);
xnor U41910 (N_41910,N_40446,N_40686);
xor U41911 (N_41911,N_40709,N_40275);
and U41912 (N_41912,N_40730,N_40545);
xnor U41913 (N_41913,N_40337,N_40700);
nand U41914 (N_41914,N_40398,N_40991);
nand U41915 (N_41915,N_40293,N_40502);
xnor U41916 (N_41916,N_40614,N_40869);
or U41917 (N_41917,N_40644,N_40535);
and U41918 (N_41918,N_40939,N_40021);
nand U41919 (N_41919,N_40673,N_40430);
nand U41920 (N_41920,N_40135,N_40989);
nand U41921 (N_41921,N_40775,N_40600);
nor U41922 (N_41922,N_40067,N_40007);
nor U41923 (N_41923,N_40517,N_40286);
or U41924 (N_41924,N_40378,N_40838);
nand U41925 (N_41925,N_40705,N_40756);
or U41926 (N_41926,N_40763,N_40521);
and U41927 (N_41927,N_40428,N_40572);
nor U41928 (N_41928,N_40345,N_40938);
nand U41929 (N_41929,N_40182,N_40118);
xnor U41930 (N_41930,N_40507,N_40091);
and U41931 (N_41931,N_40711,N_40043);
and U41932 (N_41932,N_40970,N_40450);
or U41933 (N_41933,N_40944,N_40729);
or U41934 (N_41934,N_40084,N_40542);
xnor U41935 (N_41935,N_40572,N_40815);
or U41936 (N_41936,N_40578,N_40648);
nand U41937 (N_41937,N_40611,N_40650);
nand U41938 (N_41938,N_40741,N_40526);
nor U41939 (N_41939,N_40853,N_40200);
or U41940 (N_41940,N_40888,N_40277);
xnor U41941 (N_41941,N_40103,N_40073);
nand U41942 (N_41942,N_40125,N_40363);
and U41943 (N_41943,N_40369,N_40769);
and U41944 (N_41944,N_40420,N_40884);
xnor U41945 (N_41945,N_40606,N_40474);
xnor U41946 (N_41946,N_40975,N_40962);
and U41947 (N_41947,N_40946,N_40395);
xor U41948 (N_41948,N_40050,N_40231);
nand U41949 (N_41949,N_40176,N_40679);
xnor U41950 (N_41950,N_40590,N_40354);
and U41951 (N_41951,N_40059,N_40473);
and U41952 (N_41952,N_40648,N_40757);
nand U41953 (N_41953,N_40152,N_40574);
nand U41954 (N_41954,N_40488,N_40341);
or U41955 (N_41955,N_40570,N_40038);
and U41956 (N_41956,N_40752,N_40670);
nor U41957 (N_41957,N_40492,N_40261);
xnor U41958 (N_41958,N_40557,N_40347);
nor U41959 (N_41959,N_40263,N_40801);
nand U41960 (N_41960,N_40513,N_40316);
and U41961 (N_41961,N_40106,N_40721);
nor U41962 (N_41962,N_40271,N_40539);
nor U41963 (N_41963,N_40365,N_40320);
xor U41964 (N_41964,N_40160,N_40794);
and U41965 (N_41965,N_40702,N_40985);
nor U41966 (N_41966,N_40701,N_40986);
nand U41967 (N_41967,N_40546,N_40622);
nor U41968 (N_41968,N_40979,N_40190);
and U41969 (N_41969,N_40108,N_40647);
nand U41970 (N_41970,N_40466,N_40221);
nor U41971 (N_41971,N_40036,N_40153);
and U41972 (N_41972,N_40491,N_40560);
nor U41973 (N_41973,N_40676,N_40246);
nand U41974 (N_41974,N_40273,N_40331);
and U41975 (N_41975,N_40757,N_40915);
and U41976 (N_41976,N_40909,N_40383);
nand U41977 (N_41977,N_40100,N_40509);
nand U41978 (N_41978,N_40850,N_40775);
nand U41979 (N_41979,N_40907,N_40594);
xnor U41980 (N_41980,N_40722,N_40734);
or U41981 (N_41981,N_40649,N_40553);
and U41982 (N_41982,N_40511,N_40445);
nand U41983 (N_41983,N_40979,N_40797);
and U41984 (N_41984,N_40148,N_40442);
or U41985 (N_41985,N_40880,N_40884);
nand U41986 (N_41986,N_40407,N_40270);
or U41987 (N_41987,N_40921,N_40496);
nand U41988 (N_41988,N_40566,N_40468);
nor U41989 (N_41989,N_40336,N_40566);
or U41990 (N_41990,N_40860,N_40910);
xnor U41991 (N_41991,N_40651,N_40272);
nor U41992 (N_41992,N_40968,N_40163);
nor U41993 (N_41993,N_40467,N_40717);
and U41994 (N_41994,N_40883,N_40374);
xnor U41995 (N_41995,N_40981,N_40769);
and U41996 (N_41996,N_40396,N_40282);
xnor U41997 (N_41997,N_40673,N_40345);
and U41998 (N_41998,N_40574,N_40729);
xnor U41999 (N_41999,N_40467,N_40948);
xor U42000 (N_42000,N_41315,N_41744);
and U42001 (N_42001,N_41137,N_41178);
nor U42002 (N_42002,N_41907,N_41390);
xor U42003 (N_42003,N_41291,N_41088);
and U42004 (N_42004,N_41680,N_41201);
xor U42005 (N_42005,N_41087,N_41504);
or U42006 (N_42006,N_41404,N_41584);
xnor U42007 (N_42007,N_41518,N_41117);
nand U42008 (N_42008,N_41287,N_41316);
nor U42009 (N_42009,N_41711,N_41054);
and U42010 (N_42010,N_41926,N_41600);
and U42011 (N_42011,N_41121,N_41144);
nor U42012 (N_42012,N_41927,N_41228);
xnor U42013 (N_42013,N_41164,N_41715);
and U42014 (N_42014,N_41020,N_41353);
xor U42015 (N_42015,N_41917,N_41326);
nor U42016 (N_42016,N_41629,N_41602);
and U42017 (N_42017,N_41055,N_41156);
xnor U42018 (N_42018,N_41888,N_41505);
nand U42019 (N_42019,N_41550,N_41231);
nor U42020 (N_42020,N_41666,N_41023);
or U42021 (N_42021,N_41298,N_41698);
nor U42022 (N_42022,N_41650,N_41471);
and U42023 (N_42023,N_41753,N_41241);
nand U42024 (N_42024,N_41421,N_41302);
and U42025 (N_42025,N_41370,N_41045);
or U42026 (N_42026,N_41850,N_41000);
xnor U42027 (N_42027,N_41092,N_41519);
nor U42028 (N_42028,N_41104,N_41660);
xor U42029 (N_42029,N_41940,N_41996);
xnor U42030 (N_42030,N_41070,N_41516);
nor U42031 (N_42031,N_41236,N_41759);
nand U42032 (N_42032,N_41362,N_41153);
nor U42033 (N_42033,N_41269,N_41186);
or U42034 (N_42034,N_41735,N_41638);
nor U42035 (N_42035,N_41237,N_41299);
xor U42036 (N_42036,N_41657,N_41882);
xnor U42037 (N_42037,N_41464,N_41717);
nand U42038 (N_42038,N_41322,N_41846);
or U42039 (N_42039,N_41414,N_41488);
or U42040 (N_42040,N_41774,N_41713);
nor U42041 (N_42041,N_41468,N_41154);
xnor U42042 (N_42042,N_41158,N_41565);
nand U42043 (N_42043,N_41296,N_41730);
xnor U42044 (N_42044,N_41871,N_41244);
nand U42045 (N_42045,N_41494,N_41791);
nor U42046 (N_42046,N_41247,N_41474);
and U42047 (N_42047,N_41423,N_41285);
nand U42048 (N_42048,N_41913,N_41551);
or U42049 (N_42049,N_41146,N_41443);
or U42050 (N_42050,N_41559,N_41956);
nor U42051 (N_42051,N_41470,N_41341);
or U42052 (N_42052,N_41479,N_41364);
nor U42053 (N_42053,N_41403,N_41331);
nor U42054 (N_42054,N_41668,N_41694);
or U42055 (N_42055,N_41541,N_41903);
nand U42056 (N_42056,N_41094,N_41763);
xnor U42057 (N_42057,N_41928,N_41425);
and U42058 (N_42058,N_41528,N_41978);
nand U42059 (N_42059,N_41891,N_41811);
xor U42060 (N_42060,N_41409,N_41383);
or U42061 (N_42061,N_41952,N_41567);
nor U42062 (N_42062,N_41695,N_41879);
nor U42063 (N_42063,N_41480,N_41832);
nor U42064 (N_42064,N_41789,N_41496);
nor U42065 (N_42065,N_41582,N_41204);
nor U42066 (N_42066,N_41843,N_41658);
nand U42067 (N_42067,N_41040,N_41663);
xor U42068 (N_42068,N_41161,N_41662);
and U42069 (N_42069,N_41063,N_41481);
nand U42070 (N_42070,N_41624,N_41887);
and U42071 (N_42071,N_41128,N_41416);
nand U42072 (N_42072,N_41466,N_41612);
and U42073 (N_42073,N_41642,N_41152);
xnor U42074 (N_42074,N_41323,N_41742);
nor U42075 (N_42075,N_41399,N_41263);
or U42076 (N_42076,N_41256,N_41609);
xnor U42077 (N_42077,N_41805,N_41084);
nand U42078 (N_42078,N_41223,N_41992);
xor U42079 (N_42079,N_41623,N_41982);
nor U42080 (N_42080,N_41413,N_41573);
or U42081 (N_42081,N_41706,N_41821);
nand U42082 (N_42082,N_41412,N_41794);
xnor U42083 (N_42083,N_41163,N_41841);
nor U42084 (N_42084,N_41188,N_41671);
and U42085 (N_42085,N_41553,N_41576);
nor U42086 (N_42086,N_41618,N_41656);
or U42087 (N_42087,N_41184,N_41283);
xor U42088 (N_42088,N_41393,N_41429);
and U42089 (N_42089,N_41268,N_41292);
nand U42090 (N_42090,N_41312,N_41770);
and U42091 (N_42091,N_41459,N_41886);
nor U42092 (N_42092,N_41809,N_41043);
xor U42093 (N_42093,N_41754,N_41649);
xnor U42094 (N_42094,N_41214,N_41745);
nor U42095 (N_42095,N_41066,N_41977);
and U42096 (N_42096,N_41572,N_41251);
or U42097 (N_42097,N_41571,N_41951);
nor U42098 (N_42098,N_41540,N_41093);
or U42099 (N_42099,N_41743,N_41615);
or U42100 (N_42100,N_41167,N_41611);
nor U42101 (N_42101,N_41816,N_41056);
xor U42102 (N_42102,N_41297,N_41246);
nand U42103 (N_42103,N_41890,N_41939);
nor U42104 (N_42104,N_41249,N_41591);
and U42105 (N_42105,N_41239,N_41218);
nor U42106 (N_42106,N_41342,N_41053);
or U42107 (N_42107,N_41385,N_41086);
or U42108 (N_42108,N_41257,N_41673);
nand U42109 (N_42109,N_41356,N_41529);
nand U42110 (N_42110,N_41527,N_41457);
or U42111 (N_42111,N_41508,N_41391);
and U42112 (N_42112,N_41448,N_41955);
and U42113 (N_42113,N_41039,N_41456);
xor U42114 (N_42114,N_41260,N_41530);
nor U42115 (N_42115,N_41495,N_41892);
nor U42116 (N_42116,N_41254,N_41098);
or U42117 (N_42117,N_41752,N_41445);
nand U42118 (N_42118,N_41057,N_41129);
xnor U42119 (N_42119,N_41687,N_41865);
xnor U42120 (N_42120,N_41532,N_41279);
xor U42121 (N_42121,N_41106,N_41818);
and U42122 (N_42122,N_41637,N_41845);
nand U42123 (N_42123,N_41909,N_41904);
nor U42124 (N_42124,N_41724,N_41029);
nor U42125 (N_42125,N_41962,N_41276);
or U42126 (N_42126,N_41136,N_41130);
nor U42127 (N_42127,N_41709,N_41503);
xnor U42128 (N_42128,N_41587,N_41669);
nand U42129 (N_42129,N_41595,N_41901);
or U42130 (N_42130,N_41248,N_41555);
xnor U42131 (N_42131,N_41065,N_41802);
and U42132 (N_42132,N_41242,N_41697);
or U42133 (N_42133,N_41451,N_41003);
nand U42134 (N_42134,N_41337,N_41132);
nor U42135 (N_42135,N_41621,N_41622);
xnor U42136 (N_42136,N_41286,N_41883);
nor U42137 (N_42137,N_41710,N_41936);
xor U42138 (N_42138,N_41240,N_41755);
nand U42139 (N_42139,N_41203,N_41083);
and U42140 (N_42140,N_41515,N_41741);
or U42141 (N_42141,N_41047,N_41217);
xnor U42142 (N_42142,N_41096,N_41995);
or U42143 (N_42143,N_41827,N_41513);
xor U42144 (N_42144,N_41235,N_41922);
xor U42145 (N_42145,N_41069,N_41406);
nor U42146 (N_42146,N_41112,N_41931);
nand U42147 (N_42147,N_41169,N_41213);
or U42148 (N_42148,N_41168,N_41542);
xnor U42149 (N_42149,N_41655,N_41375);
and U42150 (N_42150,N_41024,N_41386);
or U42151 (N_42151,N_41111,N_41114);
nand U42152 (N_42152,N_41199,N_41958);
nand U42153 (N_42153,N_41699,N_41351);
nor U42154 (N_42154,N_41665,N_41925);
nor U42155 (N_42155,N_41506,N_41945);
or U42156 (N_42156,N_41125,N_41373);
or U42157 (N_42157,N_41749,N_41826);
or U42158 (N_42158,N_41060,N_41659);
nor U42159 (N_42159,N_41967,N_41243);
and U42160 (N_42160,N_41603,N_41258);
or U42161 (N_42161,N_41420,N_41469);
nor U42162 (N_42162,N_41033,N_41634);
and U42163 (N_42163,N_41366,N_41233);
xor U42164 (N_42164,N_41601,N_41358);
and U42165 (N_42165,N_41580,N_41041);
xnor U42166 (N_42166,N_41549,N_41525);
nor U42167 (N_42167,N_41537,N_41177);
nor U42168 (N_42168,N_41570,N_41538);
xnor U42169 (N_42169,N_41097,N_41196);
xor U42170 (N_42170,N_41830,N_41889);
xor U42171 (N_42171,N_41905,N_41062);
xor U42172 (N_42172,N_41215,N_41746);
nor U42173 (N_42173,N_41368,N_41482);
nand U42174 (N_42174,N_41173,N_41856);
or U42175 (N_42175,N_41613,N_41971);
nor U42176 (N_42176,N_41651,N_41514);
and U42177 (N_42177,N_41190,N_41119);
and U42178 (N_42178,N_41371,N_41339);
nand U42179 (N_42179,N_41124,N_41782);
and U42180 (N_42180,N_41881,N_41498);
or U42181 (N_42181,N_41648,N_41295);
xnor U42182 (N_42182,N_41685,N_41716);
nor U42183 (N_42183,N_41738,N_41035);
nor U42184 (N_42184,N_41902,N_41736);
nand U42185 (N_42185,N_41878,N_41419);
nor U42186 (N_42186,N_41543,N_41150);
or U42187 (N_42187,N_41313,N_41009);
or U42188 (N_42188,N_41378,N_41873);
and U42189 (N_42189,N_41667,N_41628);
xor U42190 (N_42190,N_41289,N_41085);
nor U42191 (N_42191,N_41783,N_41645);
nor U42192 (N_42192,N_41729,N_41946);
or U42193 (N_42193,N_41400,N_41046);
or U42194 (N_42194,N_41325,N_41820);
xnor U42195 (N_42195,N_41044,N_41367);
and U42196 (N_42196,N_41489,N_41558);
or U42197 (N_42197,N_41290,N_41557);
xor U42198 (N_42198,N_41211,N_41510);
or U42199 (N_42199,N_41463,N_41344);
xnor U42200 (N_42200,N_41189,N_41690);
nor U42201 (N_42201,N_41853,N_41010);
nor U42202 (N_42202,N_41467,N_41885);
and U42203 (N_42203,N_41935,N_41308);
xnor U42204 (N_42204,N_41359,N_41625);
nor U42205 (N_42205,N_41038,N_41499);
or U42206 (N_42206,N_41760,N_41895);
xnor U42207 (N_42207,N_41930,N_41485);
nor U42208 (N_42208,N_41734,N_41021);
xor U42209 (N_42209,N_41472,N_41293);
xor U42210 (N_42210,N_41018,N_41548);
nor U42211 (N_42211,N_41208,N_41999);
nor U42212 (N_42212,N_41013,N_41221);
and U42213 (N_42213,N_41985,N_41216);
and U42214 (N_42214,N_41552,N_41401);
nand U42215 (N_42215,N_41860,N_41397);
nor U42216 (N_42216,N_41539,N_41327);
xnor U42217 (N_42217,N_41808,N_41116);
and U42218 (N_42218,N_41079,N_41027);
and U42219 (N_42219,N_41869,N_41959);
or U42220 (N_42220,N_41280,N_41972);
xor U42221 (N_42221,N_41226,N_41300);
xnor U42222 (N_42222,N_41197,N_41200);
or U42223 (N_42223,N_41693,N_41630);
nor U42224 (N_42224,N_41707,N_41501);
or U42225 (N_42225,N_41594,N_41672);
nand U42226 (N_42226,N_41340,N_41848);
nand U42227 (N_42227,N_41077,N_41444);
nor U42228 (N_42228,N_41354,N_41122);
xor U42229 (N_42229,N_41080,N_41034);
nor U42230 (N_42230,N_41531,N_41960);
nand U42231 (N_42231,N_41943,N_41449);
and U42232 (N_42232,N_41912,N_41365);
nand U42233 (N_42233,N_41910,N_41118);
or U42234 (N_42234,N_41181,N_41148);
or U42235 (N_42235,N_41294,N_41704);
nor U42236 (N_42236,N_41987,N_41113);
and U42237 (N_42237,N_41032,N_41149);
xnor U42238 (N_42238,N_41855,N_41437);
nor U42239 (N_42239,N_41861,N_41311);
nand U42240 (N_42240,N_41319,N_41983);
or U42241 (N_42241,N_41174,N_41374);
xor U42242 (N_42242,N_41078,N_41270);
nand U42243 (N_42243,N_41473,N_41792);
xnor U42244 (N_42244,N_41574,N_41719);
xnor U42245 (N_42245,N_41636,N_41785);
nand U42246 (N_42246,N_41031,N_41854);
or U42247 (N_42247,N_41398,N_41747);
xnor U42248 (N_42248,N_41970,N_41453);
nor U42249 (N_42249,N_41692,N_41639);
and U42250 (N_42250,N_41307,N_41844);
nand U42251 (N_42251,N_41825,N_41028);
nor U42252 (N_42252,N_41949,N_41387);
nand U42253 (N_42253,N_41646,N_41839);
nor U42254 (N_42254,N_41108,N_41721);
and U42255 (N_42255,N_41859,N_41547);
xor U42256 (N_42256,N_41415,N_41779);
nand U42257 (N_42257,N_41162,N_41918);
and U42258 (N_42258,N_41598,N_41974);
or U42259 (N_42259,N_41986,N_41012);
and U42260 (N_42260,N_41090,N_41071);
nand U42261 (N_42261,N_41633,N_41833);
nor U42262 (N_42262,N_41838,N_41522);
or U42263 (N_42263,N_41806,N_41914);
and U42264 (N_42264,N_41145,N_41817);
nor U42265 (N_42265,N_41554,N_41266);
nor U42266 (N_42266,N_41739,N_41324);
nand U42267 (N_42267,N_41059,N_41050);
nor U42268 (N_42268,N_41193,N_41352);
nand U42269 (N_42269,N_41762,N_41377);
nor U42270 (N_42270,N_41477,N_41212);
nor U42271 (N_42271,N_41617,N_41388);
nand U42272 (N_42272,N_41911,N_41487);
xnor U42273 (N_42273,N_41272,N_41253);
or U42274 (N_42274,N_41165,N_41329);
nor U42275 (N_42275,N_41123,N_41963);
or U42276 (N_42276,N_41596,N_41320);
and U42277 (N_42277,N_41544,N_41831);
nand U42278 (N_42278,N_41245,N_41684);
and U42279 (N_42279,N_41756,N_41566);
xor U42280 (N_42280,N_41402,N_41523);
and U42281 (N_42281,N_41932,N_41274);
or U42282 (N_42282,N_41748,N_41874);
and U42283 (N_42283,N_41674,N_41143);
xor U42284 (N_42284,N_41824,N_41305);
xor U42285 (N_42285,N_41728,N_41686);
or U42286 (N_42286,N_41796,N_41653);
and U42287 (N_42287,N_41751,N_41593);
xnor U42288 (N_42288,N_41703,N_41652);
xor U42289 (N_42289,N_41076,N_41176);
nand U42290 (N_42290,N_41333,N_41769);
and U42291 (N_42291,N_41369,N_41823);
xor U42292 (N_42292,N_41834,N_41405);
or U42293 (N_42293,N_41001,N_41900);
nand U42294 (N_42294,N_41647,N_41110);
nand U42295 (N_42295,N_41458,N_41768);
nor U42296 (N_42296,N_41207,N_41536);
and U42297 (N_42297,N_41640,N_41157);
and U42298 (N_42298,N_41915,N_41568);
and U42299 (N_42299,N_41195,N_41675);
and U42300 (N_42300,N_41438,N_41560);
or U42301 (N_42301,N_41379,N_41585);
nor U42302 (N_42302,N_41896,N_41075);
nor U42303 (N_42303,N_41643,N_41604);
nand U42304 (N_42304,N_41142,N_41361);
nand U42305 (N_42305,N_41546,N_41847);
or U42306 (N_42306,N_41586,N_41346);
nor U42307 (N_42307,N_41778,N_41726);
and U42308 (N_42308,N_41938,N_41064);
nand U42309 (N_42309,N_41897,N_41347);
nand U42310 (N_42310,N_41011,N_41250);
and U42311 (N_42311,N_41099,N_41599);
nor U42312 (N_42312,N_41863,N_41107);
xor U42313 (N_42313,N_41944,N_41840);
and U42314 (N_42314,N_41493,N_41284);
nand U42315 (N_42315,N_41301,N_41141);
and U42316 (N_42316,N_41082,N_41776);
xor U42317 (N_42317,N_41440,N_41229);
xnor U42318 (N_42318,N_41998,N_41517);
xnor U42319 (N_42319,N_41828,N_41973);
xnor U42320 (N_42320,N_41700,N_41407);
nor U42321 (N_42321,N_41991,N_41670);
and U42322 (N_42322,N_41589,N_41172);
nand U42323 (N_42323,N_41336,N_41455);
or U42324 (N_42324,N_41194,N_41048);
or U42325 (N_42325,N_41089,N_41431);
and U42326 (N_42326,N_41424,N_41357);
or U42327 (N_42327,N_41608,N_41417);
and U42328 (N_42328,N_41696,N_41575);
xnor U42329 (N_42329,N_41714,N_41348);
nand U42330 (N_42330,N_41921,N_41563);
xor U42331 (N_42331,N_41908,N_41758);
nand U42332 (N_42332,N_41678,N_41767);
nand U42333 (N_42333,N_41507,N_41220);
and U42334 (N_42334,N_41835,N_41275);
or U42335 (N_42335,N_41005,N_41095);
nor U42336 (N_42336,N_41264,N_41786);
nand U42337 (N_42337,N_41880,N_41372);
xor U42338 (N_42338,N_41868,N_41303);
nand U42339 (N_42339,N_41937,N_41851);
and U42340 (N_42340,N_41171,N_41984);
nor U42341 (N_42341,N_41109,N_41037);
nand U42342 (N_42342,N_41990,N_41712);
nor U42343 (N_42343,N_41395,N_41723);
and U42344 (N_42344,N_41446,N_41893);
or U42345 (N_42345,N_41780,N_41884);
and U42346 (N_42346,N_41569,N_41411);
or U42347 (N_42347,N_41583,N_41392);
nor U42348 (N_42348,N_41476,N_41968);
xor U42349 (N_42349,N_41988,N_41120);
and U42350 (N_42350,N_41965,N_41948);
and U42351 (N_42351,N_41454,N_41989);
or U42352 (N_42352,N_41829,N_41626);
and U42353 (N_42353,N_41836,N_41483);
xor U42354 (N_42354,N_41314,N_41842);
xnor U42355 (N_42355,N_41017,N_41006);
nand U42356 (N_42356,N_41664,N_41261);
and U42357 (N_42357,N_41015,N_41631);
nor U42358 (N_42358,N_41238,N_41681);
or U42359 (N_42359,N_41804,N_41961);
xor U42360 (N_42360,N_41427,N_41491);
nor U42361 (N_42361,N_41306,N_41389);
nand U42362 (N_42362,N_41100,N_41073);
xnor U42363 (N_42363,N_41036,N_41934);
nand U42364 (N_42364,N_41761,N_41206);
nor U42365 (N_42365,N_41661,N_41725);
nor U42366 (N_42366,N_41271,N_41981);
nor U42367 (N_42367,N_41798,N_41556);
and U42368 (N_42368,N_41452,N_41432);
and U42369 (N_42369,N_41533,N_41434);
nand U42370 (N_42370,N_41797,N_41318);
or U42371 (N_42371,N_41191,N_41590);
or U42372 (N_42372,N_41966,N_41183);
xor U42373 (N_42373,N_41450,N_41155);
nand U42374 (N_42374,N_41722,N_41210);
nand U42375 (N_42375,N_41683,N_41180);
and U42376 (N_42376,N_41439,N_41676);
nand U42377 (N_42377,N_41175,N_41976);
nand U42378 (N_42378,N_41534,N_41923);
and U42379 (N_42379,N_41074,N_41535);
xnor U42380 (N_42380,N_41964,N_41781);
and U42381 (N_42381,N_41511,N_41492);
nor U42382 (N_42382,N_41267,N_41230);
or U42383 (N_42383,N_41234,N_41765);
and U42384 (N_42384,N_41081,N_41870);
xnor U42385 (N_42385,N_41278,N_41102);
nor U42386 (N_42386,N_41335,N_41577);
xnor U42387 (N_42387,N_41281,N_41795);
xnor U42388 (N_42388,N_41360,N_41304);
and U42389 (N_42389,N_41330,N_41520);
and U42390 (N_42390,N_41764,N_41265);
nor U42391 (N_42391,N_41788,N_41138);
or U42392 (N_42392,N_41740,N_41259);
or U42393 (N_42393,N_41619,N_41521);
and U42394 (N_42394,N_41310,N_41866);
and U42395 (N_42395,N_41837,N_41898);
xnor U42396 (N_42396,N_41954,N_41334);
nor U42397 (N_42397,N_41159,N_41708);
or U42398 (N_42398,N_41126,N_41426);
nor U42399 (N_42399,N_41793,N_41442);
nor U42400 (N_42400,N_41408,N_41610);
nor U42401 (N_42401,N_41381,N_41564);
xnor U42402 (N_42402,N_41115,N_41933);
or U42403 (N_42403,N_41894,N_41607);
nand U42404 (N_42404,N_41997,N_41396);
or U42405 (N_42405,N_41701,N_41969);
or U42406 (N_42406,N_41497,N_41022);
or U42407 (N_42407,N_41091,N_41376);
and U42408 (N_42408,N_41813,N_41008);
or U42409 (N_42409,N_41579,N_41916);
xor U42410 (N_42410,N_41133,N_41775);
or U42411 (N_42411,N_41994,N_41321);
and U42412 (N_42412,N_41309,N_41140);
nor U42413 (N_42413,N_41677,N_41428);
xor U42414 (N_42414,N_41328,N_41441);
and U42415 (N_42415,N_41807,N_41049);
nor U42416 (N_42416,N_41799,N_41957);
xor U42417 (N_42417,N_41766,N_41151);
nand U42418 (N_42418,N_41597,N_41950);
and U42419 (N_42419,N_41877,N_41461);
xnor U42420 (N_42420,N_41147,N_41502);
xor U42421 (N_42421,N_41790,N_41410);
and U42422 (N_42422,N_41688,N_41273);
or U42423 (N_42423,N_41170,N_41475);
nor U42424 (N_42424,N_41447,N_41052);
and U42425 (N_42425,N_41876,N_41019);
xnor U42426 (N_42426,N_41350,N_41953);
or U42427 (N_42427,N_41002,N_41731);
and U42428 (N_42428,N_41864,N_41227);
or U42429 (N_42429,N_41772,N_41733);
xor U42430 (N_42430,N_41819,N_41067);
or U42431 (N_42431,N_41486,N_41562);
and U42432 (N_42432,N_41277,N_41219);
nor U42433 (N_42433,N_41222,N_41867);
and U42434 (N_42434,N_41592,N_41771);
or U42435 (N_42435,N_41422,N_41436);
nand U42436 (N_42436,N_41317,N_41578);
or U42437 (N_42437,N_41526,N_41803);
and U42438 (N_42438,N_41588,N_41872);
xor U42439 (N_42439,N_41465,N_41105);
and U42440 (N_42440,N_41166,N_41349);
xor U42441 (N_42441,N_41460,N_41288);
xnor U42442 (N_42442,N_41004,N_41332);
nor U42443 (N_42443,N_41691,N_41500);
and U42444 (N_42444,N_41906,N_41682);
nand U42445 (N_42445,N_41187,N_41490);
or U42446 (N_42446,N_41635,N_41430);
or U42447 (N_42447,N_41030,N_41042);
nor U42448 (N_42448,N_41689,N_41524);
nor U42449 (N_42449,N_41185,N_41620);
nor U42450 (N_42450,N_41561,N_41394);
nand U42451 (N_42451,N_41801,N_41727);
and U42452 (N_42452,N_41929,N_41614);
nand U42453 (N_42453,N_41192,N_41815);
nand U42454 (N_42454,N_41026,N_41947);
or U42455 (N_42455,N_41345,N_41462);
or U42456 (N_42456,N_41512,N_41435);
nor U42457 (N_42457,N_41224,N_41135);
nand U42458 (N_42458,N_41899,N_41545);
and U42459 (N_42459,N_41338,N_41072);
nand U42460 (N_42460,N_41737,N_41581);
or U42461 (N_42461,N_41255,N_41644);
and U42462 (N_42462,N_41380,N_41363);
xnor U42463 (N_42463,N_41384,N_41773);
or U42464 (N_42464,N_41732,N_41757);
nand U42465 (N_42465,N_41016,N_41993);
xnor U42466 (N_42466,N_41014,N_41810);
nor U42467 (N_42467,N_41857,N_41209);
and U42468 (N_42468,N_41205,N_41777);
nor U42469 (N_42469,N_41606,N_41919);
xnor U42470 (N_42470,N_41858,N_41252);
or U42471 (N_42471,N_41616,N_41979);
and U42472 (N_42472,N_41051,N_41509);
or U42473 (N_42473,N_41179,N_41980);
or U42474 (N_42474,N_41750,N_41182);
or U42475 (N_42475,N_41225,N_41852);
nand U42476 (N_42476,N_41679,N_41941);
or U42477 (N_42477,N_41705,N_41127);
or U42478 (N_42478,N_41814,N_41160);
nor U42479 (N_42479,N_41718,N_41924);
xnor U42480 (N_42480,N_41103,N_41382);
and U42481 (N_42481,N_41282,N_41920);
nand U42482 (N_42482,N_41942,N_41007);
nand U42483 (N_42483,N_41849,N_41641);
nand U42484 (N_42484,N_41632,N_41787);
nand U42485 (N_42485,N_41812,N_41068);
nor U42486 (N_42486,N_41605,N_41822);
nand U42487 (N_42487,N_41134,N_41862);
xor U42488 (N_42488,N_41433,N_41784);
or U42489 (N_42489,N_41702,N_41800);
and U42490 (N_42490,N_41025,N_41139);
nand U42491 (N_42491,N_41720,N_41131);
nor U42492 (N_42492,N_41484,N_41975);
and U42493 (N_42493,N_41355,N_41418);
xnor U42494 (N_42494,N_41058,N_41061);
nor U42495 (N_42495,N_41627,N_41654);
xor U42496 (N_42496,N_41262,N_41202);
nand U42497 (N_42497,N_41232,N_41101);
and U42498 (N_42498,N_41198,N_41343);
nor U42499 (N_42499,N_41875,N_41478);
and U42500 (N_42500,N_41337,N_41072);
nand U42501 (N_42501,N_41792,N_41071);
nor U42502 (N_42502,N_41953,N_41138);
and U42503 (N_42503,N_41119,N_41817);
nor U42504 (N_42504,N_41777,N_41644);
or U42505 (N_42505,N_41582,N_41091);
xnor U42506 (N_42506,N_41623,N_41779);
and U42507 (N_42507,N_41895,N_41666);
xnor U42508 (N_42508,N_41378,N_41509);
nand U42509 (N_42509,N_41251,N_41173);
or U42510 (N_42510,N_41969,N_41852);
nor U42511 (N_42511,N_41450,N_41511);
and U42512 (N_42512,N_41036,N_41771);
and U42513 (N_42513,N_41338,N_41165);
nand U42514 (N_42514,N_41090,N_41219);
and U42515 (N_42515,N_41716,N_41865);
xor U42516 (N_42516,N_41526,N_41718);
nand U42517 (N_42517,N_41841,N_41343);
nor U42518 (N_42518,N_41764,N_41301);
nand U42519 (N_42519,N_41143,N_41824);
nand U42520 (N_42520,N_41902,N_41358);
xnor U42521 (N_42521,N_41790,N_41262);
and U42522 (N_42522,N_41712,N_41043);
and U42523 (N_42523,N_41509,N_41769);
or U42524 (N_42524,N_41525,N_41935);
nor U42525 (N_42525,N_41553,N_41441);
or U42526 (N_42526,N_41639,N_41316);
xnor U42527 (N_42527,N_41319,N_41290);
or U42528 (N_42528,N_41925,N_41574);
nor U42529 (N_42529,N_41105,N_41351);
and U42530 (N_42530,N_41151,N_41640);
and U42531 (N_42531,N_41241,N_41221);
xor U42532 (N_42532,N_41467,N_41539);
or U42533 (N_42533,N_41787,N_41142);
nand U42534 (N_42534,N_41907,N_41389);
and U42535 (N_42535,N_41267,N_41795);
or U42536 (N_42536,N_41586,N_41787);
nand U42537 (N_42537,N_41166,N_41068);
xor U42538 (N_42538,N_41945,N_41568);
xnor U42539 (N_42539,N_41251,N_41644);
nor U42540 (N_42540,N_41798,N_41783);
or U42541 (N_42541,N_41681,N_41348);
or U42542 (N_42542,N_41581,N_41410);
nor U42543 (N_42543,N_41001,N_41321);
nor U42544 (N_42544,N_41231,N_41954);
nand U42545 (N_42545,N_41080,N_41883);
and U42546 (N_42546,N_41891,N_41968);
and U42547 (N_42547,N_41734,N_41951);
nand U42548 (N_42548,N_41518,N_41995);
and U42549 (N_42549,N_41242,N_41089);
nand U42550 (N_42550,N_41291,N_41053);
or U42551 (N_42551,N_41038,N_41136);
xor U42552 (N_42552,N_41621,N_41876);
nand U42553 (N_42553,N_41540,N_41817);
nor U42554 (N_42554,N_41707,N_41647);
xnor U42555 (N_42555,N_41188,N_41797);
or U42556 (N_42556,N_41024,N_41375);
xor U42557 (N_42557,N_41916,N_41358);
xor U42558 (N_42558,N_41979,N_41177);
or U42559 (N_42559,N_41288,N_41715);
xnor U42560 (N_42560,N_41341,N_41862);
or U42561 (N_42561,N_41565,N_41059);
xnor U42562 (N_42562,N_41607,N_41054);
and U42563 (N_42563,N_41895,N_41938);
and U42564 (N_42564,N_41011,N_41258);
and U42565 (N_42565,N_41155,N_41972);
nor U42566 (N_42566,N_41512,N_41495);
nor U42567 (N_42567,N_41958,N_41636);
xnor U42568 (N_42568,N_41981,N_41243);
xnor U42569 (N_42569,N_41161,N_41901);
and U42570 (N_42570,N_41563,N_41255);
xor U42571 (N_42571,N_41331,N_41734);
nor U42572 (N_42572,N_41686,N_41878);
nand U42573 (N_42573,N_41166,N_41861);
and U42574 (N_42574,N_41515,N_41751);
nor U42575 (N_42575,N_41467,N_41978);
or U42576 (N_42576,N_41432,N_41317);
nor U42577 (N_42577,N_41006,N_41810);
nand U42578 (N_42578,N_41030,N_41671);
and U42579 (N_42579,N_41061,N_41826);
nand U42580 (N_42580,N_41740,N_41147);
nor U42581 (N_42581,N_41320,N_41455);
and U42582 (N_42582,N_41893,N_41457);
xor U42583 (N_42583,N_41873,N_41950);
or U42584 (N_42584,N_41614,N_41265);
nor U42585 (N_42585,N_41976,N_41096);
and U42586 (N_42586,N_41541,N_41400);
or U42587 (N_42587,N_41242,N_41379);
and U42588 (N_42588,N_41536,N_41783);
or U42589 (N_42589,N_41296,N_41297);
or U42590 (N_42590,N_41983,N_41205);
and U42591 (N_42591,N_41592,N_41363);
nand U42592 (N_42592,N_41962,N_41076);
or U42593 (N_42593,N_41301,N_41847);
nor U42594 (N_42594,N_41950,N_41309);
or U42595 (N_42595,N_41229,N_41789);
and U42596 (N_42596,N_41857,N_41037);
and U42597 (N_42597,N_41952,N_41213);
and U42598 (N_42598,N_41515,N_41247);
or U42599 (N_42599,N_41480,N_41406);
nand U42600 (N_42600,N_41768,N_41559);
and U42601 (N_42601,N_41469,N_41172);
nor U42602 (N_42602,N_41990,N_41053);
nor U42603 (N_42603,N_41160,N_41812);
and U42604 (N_42604,N_41964,N_41883);
or U42605 (N_42605,N_41922,N_41813);
nand U42606 (N_42606,N_41016,N_41121);
and U42607 (N_42607,N_41616,N_41801);
or U42608 (N_42608,N_41856,N_41272);
nand U42609 (N_42609,N_41533,N_41321);
nor U42610 (N_42610,N_41719,N_41551);
or U42611 (N_42611,N_41028,N_41442);
nor U42612 (N_42612,N_41116,N_41520);
xnor U42613 (N_42613,N_41794,N_41464);
and U42614 (N_42614,N_41392,N_41034);
xnor U42615 (N_42615,N_41551,N_41414);
nor U42616 (N_42616,N_41343,N_41653);
xnor U42617 (N_42617,N_41340,N_41043);
or U42618 (N_42618,N_41740,N_41155);
nand U42619 (N_42619,N_41525,N_41817);
or U42620 (N_42620,N_41384,N_41705);
and U42621 (N_42621,N_41905,N_41119);
and U42622 (N_42622,N_41363,N_41150);
nand U42623 (N_42623,N_41133,N_41210);
nand U42624 (N_42624,N_41700,N_41643);
and U42625 (N_42625,N_41396,N_41183);
or U42626 (N_42626,N_41786,N_41538);
nor U42627 (N_42627,N_41689,N_41777);
nand U42628 (N_42628,N_41882,N_41950);
nor U42629 (N_42629,N_41804,N_41848);
xor U42630 (N_42630,N_41041,N_41187);
nand U42631 (N_42631,N_41348,N_41605);
or U42632 (N_42632,N_41758,N_41034);
or U42633 (N_42633,N_41997,N_41052);
or U42634 (N_42634,N_41793,N_41997);
nand U42635 (N_42635,N_41279,N_41560);
xor U42636 (N_42636,N_41295,N_41223);
and U42637 (N_42637,N_41525,N_41960);
nand U42638 (N_42638,N_41368,N_41018);
nor U42639 (N_42639,N_41250,N_41186);
nor U42640 (N_42640,N_41310,N_41750);
and U42641 (N_42641,N_41301,N_41775);
or U42642 (N_42642,N_41090,N_41211);
xnor U42643 (N_42643,N_41839,N_41118);
nand U42644 (N_42644,N_41129,N_41936);
and U42645 (N_42645,N_41306,N_41195);
nand U42646 (N_42646,N_41008,N_41531);
and U42647 (N_42647,N_41299,N_41932);
xnor U42648 (N_42648,N_41203,N_41096);
nor U42649 (N_42649,N_41634,N_41912);
xnor U42650 (N_42650,N_41145,N_41033);
and U42651 (N_42651,N_41763,N_41663);
xnor U42652 (N_42652,N_41729,N_41933);
nand U42653 (N_42653,N_41036,N_41406);
nand U42654 (N_42654,N_41353,N_41088);
nor U42655 (N_42655,N_41844,N_41358);
nand U42656 (N_42656,N_41343,N_41159);
nor U42657 (N_42657,N_41604,N_41582);
xor U42658 (N_42658,N_41098,N_41741);
or U42659 (N_42659,N_41145,N_41158);
or U42660 (N_42660,N_41612,N_41204);
nor U42661 (N_42661,N_41164,N_41441);
xor U42662 (N_42662,N_41316,N_41292);
and U42663 (N_42663,N_41542,N_41565);
nor U42664 (N_42664,N_41440,N_41678);
nand U42665 (N_42665,N_41136,N_41196);
and U42666 (N_42666,N_41623,N_41602);
nand U42667 (N_42667,N_41683,N_41763);
nor U42668 (N_42668,N_41274,N_41993);
nand U42669 (N_42669,N_41321,N_41641);
nor U42670 (N_42670,N_41646,N_41570);
and U42671 (N_42671,N_41397,N_41921);
nor U42672 (N_42672,N_41959,N_41439);
xnor U42673 (N_42673,N_41224,N_41342);
nor U42674 (N_42674,N_41025,N_41330);
xnor U42675 (N_42675,N_41752,N_41249);
nand U42676 (N_42676,N_41483,N_41214);
and U42677 (N_42677,N_41035,N_41412);
xor U42678 (N_42678,N_41670,N_41863);
or U42679 (N_42679,N_41739,N_41289);
and U42680 (N_42680,N_41259,N_41378);
nand U42681 (N_42681,N_41394,N_41865);
nor U42682 (N_42682,N_41292,N_41384);
or U42683 (N_42683,N_41304,N_41211);
nor U42684 (N_42684,N_41239,N_41698);
nor U42685 (N_42685,N_41555,N_41005);
xnor U42686 (N_42686,N_41262,N_41782);
nor U42687 (N_42687,N_41687,N_41390);
nand U42688 (N_42688,N_41217,N_41530);
or U42689 (N_42689,N_41814,N_41108);
and U42690 (N_42690,N_41385,N_41340);
xnor U42691 (N_42691,N_41191,N_41951);
nor U42692 (N_42692,N_41357,N_41503);
and U42693 (N_42693,N_41883,N_41659);
and U42694 (N_42694,N_41626,N_41886);
and U42695 (N_42695,N_41122,N_41424);
and U42696 (N_42696,N_41232,N_41703);
nor U42697 (N_42697,N_41624,N_41307);
nor U42698 (N_42698,N_41759,N_41148);
and U42699 (N_42699,N_41458,N_41311);
or U42700 (N_42700,N_41221,N_41169);
nand U42701 (N_42701,N_41213,N_41269);
and U42702 (N_42702,N_41013,N_41956);
or U42703 (N_42703,N_41619,N_41054);
or U42704 (N_42704,N_41761,N_41465);
nor U42705 (N_42705,N_41932,N_41296);
and U42706 (N_42706,N_41315,N_41183);
xor U42707 (N_42707,N_41363,N_41236);
or U42708 (N_42708,N_41384,N_41382);
nand U42709 (N_42709,N_41951,N_41111);
xnor U42710 (N_42710,N_41237,N_41171);
nand U42711 (N_42711,N_41210,N_41610);
xnor U42712 (N_42712,N_41902,N_41664);
nand U42713 (N_42713,N_41205,N_41510);
or U42714 (N_42714,N_41628,N_41882);
nand U42715 (N_42715,N_41129,N_41944);
nor U42716 (N_42716,N_41922,N_41116);
and U42717 (N_42717,N_41895,N_41221);
nand U42718 (N_42718,N_41443,N_41749);
and U42719 (N_42719,N_41956,N_41306);
and U42720 (N_42720,N_41697,N_41530);
nand U42721 (N_42721,N_41288,N_41692);
xor U42722 (N_42722,N_41224,N_41404);
and U42723 (N_42723,N_41226,N_41067);
or U42724 (N_42724,N_41406,N_41509);
and U42725 (N_42725,N_41795,N_41085);
and U42726 (N_42726,N_41468,N_41530);
and U42727 (N_42727,N_41421,N_41224);
xnor U42728 (N_42728,N_41158,N_41731);
xor U42729 (N_42729,N_41787,N_41375);
xnor U42730 (N_42730,N_41279,N_41695);
or U42731 (N_42731,N_41456,N_41035);
and U42732 (N_42732,N_41537,N_41022);
nand U42733 (N_42733,N_41699,N_41856);
xnor U42734 (N_42734,N_41926,N_41442);
nor U42735 (N_42735,N_41884,N_41307);
nor U42736 (N_42736,N_41125,N_41029);
xor U42737 (N_42737,N_41266,N_41968);
or U42738 (N_42738,N_41600,N_41797);
nand U42739 (N_42739,N_41773,N_41980);
nand U42740 (N_42740,N_41915,N_41195);
and U42741 (N_42741,N_41634,N_41746);
nand U42742 (N_42742,N_41521,N_41263);
and U42743 (N_42743,N_41382,N_41125);
and U42744 (N_42744,N_41513,N_41550);
or U42745 (N_42745,N_41561,N_41937);
nor U42746 (N_42746,N_41121,N_41801);
nor U42747 (N_42747,N_41043,N_41154);
or U42748 (N_42748,N_41512,N_41123);
xor U42749 (N_42749,N_41458,N_41847);
nor U42750 (N_42750,N_41349,N_41888);
and U42751 (N_42751,N_41282,N_41369);
and U42752 (N_42752,N_41661,N_41276);
nor U42753 (N_42753,N_41564,N_41790);
or U42754 (N_42754,N_41977,N_41894);
and U42755 (N_42755,N_41476,N_41865);
or U42756 (N_42756,N_41660,N_41117);
or U42757 (N_42757,N_41454,N_41541);
or U42758 (N_42758,N_41989,N_41958);
and U42759 (N_42759,N_41362,N_41253);
nand U42760 (N_42760,N_41487,N_41852);
nor U42761 (N_42761,N_41288,N_41746);
xnor U42762 (N_42762,N_41596,N_41775);
or U42763 (N_42763,N_41384,N_41597);
nand U42764 (N_42764,N_41585,N_41163);
and U42765 (N_42765,N_41406,N_41356);
xor U42766 (N_42766,N_41348,N_41461);
or U42767 (N_42767,N_41010,N_41499);
xnor U42768 (N_42768,N_41301,N_41499);
nand U42769 (N_42769,N_41803,N_41250);
nor U42770 (N_42770,N_41049,N_41523);
xnor U42771 (N_42771,N_41494,N_41113);
nor U42772 (N_42772,N_41350,N_41627);
xnor U42773 (N_42773,N_41282,N_41193);
nor U42774 (N_42774,N_41219,N_41694);
nand U42775 (N_42775,N_41450,N_41750);
or U42776 (N_42776,N_41370,N_41942);
nand U42777 (N_42777,N_41022,N_41449);
or U42778 (N_42778,N_41351,N_41942);
xnor U42779 (N_42779,N_41506,N_41042);
xnor U42780 (N_42780,N_41747,N_41828);
xor U42781 (N_42781,N_41975,N_41631);
or U42782 (N_42782,N_41923,N_41230);
or U42783 (N_42783,N_41505,N_41363);
and U42784 (N_42784,N_41315,N_41780);
and U42785 (N_42785,N_41599,N_41842);
and U42786 (N_42786,N_41905,N_41536);
xor U42787 (N_42787,N_41716,N_41220);
or U42788 (N_42788,N_41717,N_41853);
nor U42789 (N_42789,N_41147,N_41737);
nor U42790 (N_42790,N_41335,N_41101);
or U42791 (N_42791,N_41826,N_41322);
or U42792 (N_42792,N_41055,N_41006);
and U42793 (N_42793,N_41331,N_41722);
xnor U42794 (N_42794,N_41112,N_41355);
nor U42795 (N_42795,N_41606,N_41855);
nand U42796 (N_42796,N_41655,N_41874);
and U42797 (N_42797,N_41909,N_41688);
nor U42798 (N_42798,N_41805,N_41679);
xnor U42799 (N_42799,N_41730,N_41909);
and U42800 (N_42800,N_41937,N_41134);
or U42801 (N_42801,N_41810,N_41706);
or U42802 (N_42802,N_41257,N_41100);
nor U42803 (N_42803,N_41313,N_41585);
xor U42804 (N_42804,N_41769,N_41427);
nor U42805 (N_42805,N_41572,N_41957);
nor U42806 (N_42806,N_41868,N_41434);
nor U42807 (N_42807,N_41073,N_41150);
nand U42808 (N_42808,N_41554,N_41227);
nand U42809 (N_42809,N_41767,N_41604);
or U42810 (N_42810,N_41635,N_41632);
and U42811 (N_42811,N_41855,N_41600);
and U42812 (N_42812,N_41637,N_41336);
xor U42813 (N_42813,N_41040,N_41127);
and U42814 (N_42814,N_41057,N_41230);
or U42815 (N_42815,N_41256,N_41283);
nor U42816 (N_42816,N_41653,N_41600);
xor U42817 (N_42817,N_41793,N_41711);
nor U42818 (N_42818,N_41833,N_41488);
and U42819 (N_42819,N_41250,N_41401);
and U42820 (N_42820,N_41291,N_41179);
or U42821 (N_42821,N_41551,N_41821);
nor U42822 (N_42822,N_41677,N_41935);
and U42823 (N_42823,N_41546,N_41614);
nand U42824 (N_42824,N_41715,N_41307);
or U42825 (N_42825,N_41945,N_41065);
nor U42826 (N_42826,N_41268,N_41397);
and U42827 (N_42827,N_41687,N_41163);
or U42828 (N_42828,N_41296,N_41852);
xnor U42829 (N_42829,N_41291,N_41469);
nand U42830 (N_42830,N_41456,N_41429);
and U42831 (N_42831,N_41541,N_41007);
xor U42832 (N_42832,N_41515,N_41188);
nor U42833 (N_42833,N_41211,N_41763);
nand U42834 (N_42834,N_41874,N_41132);
nand U42835 (N_42835,N_41371,N_41721);
nor U42836 (N_42836,N_41263,N_41368);
or U42837 (N_42837,N_41887,N_41261);
xnor U42838 (N_42838,N_41706,N_41074);
xnor U42839 (N_42839,N_41863,N_41534);
nand U42840 (N_42840,N_41687,N_41419);
or U42841 (N_42841,N_41223,N_41312);
nor U42842 (N_42842,N_41058,N_41723);
xor U42843 (N_42843,N_41264,N_41881);
nor U42844 (N_42844,N_41292,N_41469);
nand U42845 (N_42845,N_41893,N_41233);
or U42846 (N_42846,N_41014,N_41312);
nor U42847 (N_42847,N_41567,N_41824);
and U42848 (N_42848,N_41293,N_41003);
and U42849 (N_42849,N_41124,N_41364);
xnor U42850 (N_42850,N_41259,N_41699);
xnor U42851 (N_42851,N_41613,N_41311);
and U42852 (N_42852,N_41053,N_41055);
xnor U42853 (N_42853,N_41859,N_41642);
or U42854 (N_42854,N_41503,N_41131);
nand U42855 (N_42855,N_41134,N_41275);
nor U42856 (N_42856,N_41137,N_41221);
or U42857 (N_42857,N_41609,N_41356);
xor U42858 (N_42858,N_41915,N_41940);
xor U42859 (N_42859,N_41019,N_41390);
nand U42860 (N_42860,N_41701,N_41436);
and U42861 (N_42861,N_41768,N_41732);
nor U42862 (N_42862,N_41484,N_41839);
nor U42863 (N_42863,N_41401,N_41514);
nand U42864 (N_42864,N_41541,N_41933);
nor U42865 (N_42865,N_41493,N_41176);
and U42866 (N_42866,N_41525,N_41507);
xor U42867 (N_42867,N_41705,N_41561);
and U42868 (N_42868,N_41414,N_41441);
or U42869 (N_42869,N_41959,N_41295);
or U42870 (N_42870,N_41658,N_41551);
nand U42871 (N_42871,N_41730,N_41829);
or U42872 (N_42872,N_41556,N_41447);
xnor U42873 (N_42873,N_41459,N_41639);
and U42874 (N_42874,N_41196,N_41252);
and U42875 (N_42875,N_41314,N_41179);
xnor U42876 (N_42876,N_41754,N_41675);
or U42877 (N_42877,N_41219,N_41315);
or U42878 (N_42878,N_41387,N_41130);
nand U42879 (N_42879,N_41887,N_41380);
nand U42880 (N_42880,N_41286,N_41276);
xnor U42881 (N_42881,N_41993,N_41148);
nand U42882 (N_42882,N_41162,N_41568);
and U42883 (N_42883,N_41733,N_41458);
nor U42884 (N_42884,N_41619,N_41182);
nor U42885 (N_42885,N_41285,N_41950);
xor U42886 (N_42886,N_41287,N_41955);
nand U42887 (N_42887,N_41316,N_41224);
and U42888 (N_42888,N_41004,N_41519);
or U42889 (N_42889,N_41472,N_41769);
nand U42890 (N_42890,N_41032,N_41884);
or U42891 (N_42891,N_41719,N_41155);
nand U42892 (N_42892,N_41827,N_41787);
and U42893 (N_42893,N_41098,N_41829);
and U42894 (N_42894,N_41134,N_41522);
xor U42895 (N_42895,N_41775,N_41132);
nor U42896 (N_42896,N_41382,N_41019);
nor U42897 (N_42897,N_41761,N_41714);
and U42898 (N_42898,N_41944,N_41038);
nor U42899 (N_42899,N_41398,N_41495);
nor U42900 (N_42900,N_41816,N_41431);
nor U42901 (N_42901,N_41228,N_41739);
nor U42902 (N_42902,N_41383,N_41672);
xor U42903 (N_42903,N_41946,N_41715);
or U42904 (N_42904,N_41179,N_41255);
nand U42905 (N_42905,N_41601,N_41375);
and U42906 (N_42906,N_41694,N_41764);
nor U42907 (N_42907,N_41171,N_41628);
or U42908 (N_42908,N_41065,N_41416);
or U42909 (N_42909,N_41745,N_41856);
and U42910 (N_42910,N_41355,N_41264);
nor U42911 (N_42911,N_41106,N_41908);
nand U42912 (N_42912,N_41472,N_41977);
nand U42913 (N_42913,N_41188,N_41984);
nand U42914 (N_42914,N_41702,N_41314);
nand U42915 (N_42915,N_41797,N_41424);
and U42916 (N_42916,N_41200,N_41569);
and U42917 (N_42917,N_41895,N_41012);
nor U42918 (N_42918,N_41826,N_41190);
xor U42919 (N_42919,N_41520,N_41019);
xor U42920 (N_42920,N_41474,N_41795);
or U42921 (N_42921,N_41033,N_41110);
nand U42922 (N_42922,N_41633,N_41685);
and U42923 (N_42923,N_41241,N_41954);
nor U42924 (N_42924,N_41798,N_41356);
xnor U42925 (N_42925,N_41729,N_41654);
or U42926 (N_42926,N_41067,N_41607);
xor U42927 (N_42927,N_41836,N_41882);
nor U42928 (N_42928,N_41533,N_41651);
nor U42929 (N_42929,N_41688,N_41090);
or U42930 (N_42930,N_41049,N_41405);
nor U42931 (N_42931,N_41207,N_41629);
nand U42932 (N_42932,N_41059,N_41698);
nor U42933 (N_42933,N_41765,N_41590);
nand U42934 (N_42934,N_41678,N_41900);
or U42935 (N_42935,N_41827,N_41502);
xnor U42936 (N_42936,N_41894,N_41726);
or U42937 (N_42937,N_41017,N_41020);
nand U42938 (N_42938,N_41146,N_41745);
nand U42939 (N_42939,N_41031,N_41094);
nand U42940 (N_42940,N_41455,N_41810);
xnor U42941 (N_42941,N_41054,N_41951);
nand U42942 (N_42942,N_41381,N_41086);
xor U42943 (N_42943,N_41352,N_41592);
nor U42944 (N_42944,N_41901,N_41896);
nand U42945 (N_42945,N_41882,N_41776);
or U42946 (N_42946,N_41975,N_41120);
or U42947 (N_42947,N_41589,N_41161);
and U42948 (N_42948,N_41051,N_41254);
nor U42949 (N_42949,N_41483,N_41778);
and U42950 (N_42950,N_41214,N_41809);
xor U42951 (N_42951,N_41381,N_41311);
and U42952 (N_42952,N_41022,N_41338);
xor U42953 (N_42953,N_41592,N_41690);
nor U42954 (N_42954,N_41671,N_41309);
or U42955 (N_42955,N_41015,N_41134);
or U42956 (N_42956,N_41411,N_41320);
nor U42957 (N_42957,N_41155,N_41920);
nand U42958 (N_42958,N_41328,N_41874);
nor U42959 (N_42959,N_41375,N_41945);
xor U42960 (N_42960,N_41217,N_41762);
or U42961 (N_42961,N_41636,N_41418);
nor U42962 (N_42962,N_41330,N_41346);
and U42963 (N_42963,N_41788,N_41075);
nand U42964 (N_42964,N_41416,N_41398);
and U42965 (N_42965,N_41131,N_41536);
xor U42966 (N_42966,N_41420,N_41041);
nand U42967 (N_42967,N_41240,N_41474);
xor U42968 (N_42968,N_41624,N_41168);
or U42969 (N_42969,N_41974,N_41831);
xnor U42970 (N_42970,N_41769,N_41475);
xor U42971 (N_42971,N_41152,N_41132);
and U42972 (N_42972,N_41262,N_41405);
nor U42973 (N_42973,N_41033,N_41479);
or U42974 (N_42974,N_41855,N_41889);
or U42975 (N_42975,N_41162,N_41887);
nor U42976 (N_42976,N_41233,N_41775);
nor U42977 (N_42977,N_41030,N_41788);
xnor U42978 (N_42978,N_41478,N_41515);
or U42979 (N_42979,N_41905,N_41112);
and U42980 (N_42980,N_41763,N_41186);
or U42981 (N_42981,N_41215,N_41541);
nand U42982 (N_42982,N_41842,N_41311);
nor U42983 (N_42983,N_41924,N_41233);
and U42984 (N_42984,N_41566,N_41690);
nor U42985 (N_42985,N_41232,N_41522);
and U42986 (N_42986,N_41407,N_41298);
and U42987 (N_42987,N_41971,N_41149);
and U42988 (N_42988,N_41028,N_41238);
xor U42989 (N_42989,N_41157,N_41415);
nor U42990 (N_42990,N_41946,N_41319);
and U42991 (N_42991,N_41347,N_41344);
nor U42992 (N_42992,N_41071,N_41166);
nor U42993 (N_42993,N_41353,N_41997);
xnor U42994 (N_42994,N_41722,N_41353);
or U42995 (N_42995,N_41446,N_41414);
nand U42996 (N_42996,N_41339,N_41529);
nor U42997 (N_42997,N_41717,N_41574);
xnor U42998 (N_42998,N_41362,N_41199);
or U42999 (N_42999,N_41400,N_41028);
nor U43000 (N_43000,N_42234,N_42772);
and U43001 (N_43001,N_42010,N_42823);
or U43002 (N_43002,N_42703,N_42609);
nor U43003 (N_43003,N_42247,N_42924);
nand U43004 (N_43004,N_42559,N_42921);
and U43005 (N_43005,N_42911,N_42412);
and U43006 (N_43006,N_42202,N_42811);
nand U43007 (N_43007,N_42518,N_42131);
nor U43008 (N_43008,N_42012,N_42089);
nor U43009 (N_43009,N_42099,N_42425);
nor U43010 (N_43010,N_42964,N_42153);
xor U43011 (N_43011,N_42834,N_42997);
xnor U43012 (N_43012,N_42747,N_42926);
xor U43013 (N_43013,N_42646,N_42375);
and U43014 (N_43014,N_42711,N_42126);
nor U43015 (N_43015,N_42593,N_42041);
xor U43016 (N_43016,N_42420,N_42750);
nor U43017 (N_43017,N_42098,N_42956);
xnor U43018 (N_43018,N_42249,N_42695);
and U43019 (N_43019,N_42394,N_42773);
and U43020 (N_43020,N_42105,N_42951);
nand U43021 (N_43021,N_42448,N_42108);
or U43022 (N_43022,N_42831,N_42349);
nand U43023 (N_43023,N_42584,N_42445);
nor U43024 (N_43024,N_42193,N_42026);
xnor U43025 (N_43025,N_42158,N_42875);
nor U43026 (N_43026,N_42553,N_42621);
or U43027 (N_43027,N_42838,N_42051);
or U43028 (N_43028,N_42683,N_42025);
nor U43029 (N_43029,N_42873,N_42432);
and U43030 (N_43030,N_42916,N_42931);
xnor U43031 (N_43031,N_42038,N_42169);
nor U43032 (N_43032,N_42639,N_42685);
nand U43033 (N_43033,N_42334,N_42179);
nand U43034 (N_43034,N_42952,N_42517);
nor U43035 (N_43035,N_42422,N_42242);
and U43036 (N_43036,N_42266,N_42653);
xor U43037 (N_43037,N_42635,N_42596);
and U43038 (N_43038,N_42801,N_42171);
nand U43039 (N_43039,N_42223,N_42970);
xnor U43040 (N_43040,N_42476,N_42315);
or U43041 (N_43041,N_42037,N_42787);
nand U43042 (N_43042,N_42427,N_42002);
nand U43043 (N_43043,N_42638,N_42577);
xor U43044 (N_43044,N_42728,N_42307);
and U43045 (N_43045,N_42554,N_42156);
nor U43046 (N_43046,N_42928,N_42339);
nand U43047 (N_43047,N_42570,N_42246);
and U43048 (N_43048,N_42740,N_42119);
or U43049 (N_43049,N_42059,N_42331);
nor U43050 (N_43050,N_42645,N_42742);
nor U43051 (N_43051,N_42228,N_42981);
and U43052 (N_43052,N_42846,N_42194);
nor U43053 (N_43053,N_42473,N_42729);
or U43054 (N_43054,N_42296,N_42879);
nor U43055 (N_43055,N_42201,N_42550);
nand U43056 (N_43056,N_42467,N_42456);
or U43057 (N_43057,N_42894,N_42352);
or U43058 (N_43058,N_42035,N_42631);
and U43059 (N_43059,N_42763,N_42492);
nor U43060 (N_43060,N_42810,N_42450);
or U43061 (N_43061,N_42177,N_42039);
and U43062 (N_43062,N_42960,N_42084);
xor U43063 (N_43063,N_42140,N_42583);
or U43064 (N_43064,N_42321,N_42691);
xor U43065 (N_43065,N_42187,N_42300);
xnor U43066 (N_43066,N_42664,N_42566);
or U43067 (N_43067,N_42154,N_42071);
or U43068 (N_43068,N_42805,N_42398);
nand U43069 (N_43069,N_42934,N_42819);
nor U43070 (N_43070,N_42723,N_42876);
and U43071 (N_43071,N_42627,N_42016);
and U43072 (N_43072,N_42735,N_42895);
nand U43073 (N_43073,N_42898,N_42047);
xnor U43074 (N_43074,N_42549,N_42245);
and U43075 (N_43075,N_42243,N_42438);
or U43076 (N_43076,N_42910,N_42330);
xnor U43077 (N_43077,N_42062,N_42044);
xor U43078 (N_43078,N_42994,N_42305);
and U43079 (N_43079,N_42824,N_42925);
xor U43080 (N_43080,N_42142,N_42258);
nor U43081 (N_43081,N_42930,N_42019);
or U43082 (N_43082,N_42213,N_42594);
and U43083 (N_43083,N_42097,N_42125);
xnor U43084 (N_43084,N_42340,N_42409);
or U43085 (N_43085,N_42066,N_42705);
and U43086 (N_43086,N_42919,N_42618);
nand U43087 (N_43087,N_42157,N_42985);
and U43088 (N_43088,N_42459,N_42168);
xor U43089 (N_43089,N_42807,N_42866);
or U43090 (N_43090,N_42795,N_42411);
or U43091 (N_43091,N_42122,N_42941);
nand U43092 (N_43092,N_42607,N_42480);
and U43093 (N_43093,N_42498,N_42058);
and U43094 (N_43094,N_42167,N_42030);
nor U43095 (N_43095,N_42999,N_42995);
xnor U43096 (N_43096,N_42046,N_42946);
or U43097 (N_43097,N_42830,N_42967);
xnor U43098 (N_43098,N_42588,N_42191);
and U43099 (N_43099,N_42651,N_42575);
nand U43100 (N_43100,N_42185,N_42990);
nand U43101 (N_43101,N_42354,N_42102);
nand U43102 (N_43102,N_42989,N_42786);
nor U43103 (N_43103,N_42617,N_42769);
nand U43104 (N_43104,N_42240,N_42762);
xnor U43105 (N_43105,N_42103,N_42181);
or U43106 (N_43106,N_42272,N_42504);
or U43107 (N_43107,N_42820,N_42494);
or U43108 (N_43108,N_42392,N_42915);
nor U43109 (N_43109,N_42225,N_42310);
nor U43110 (N_43110,N_42341,N_42903);
nand U43111 (N_43111,N_42332,N_42610);
and U43112 (N_43112,N_42260,N_42835);
nand U43113 (N_43113,N_42658,N_42690);
xor U43114 (N_43114,N_42731,N_42912);
or U43115 (N_43115,N_42464,N_42348);
xor U43116 (N_43116,N_42086,N_42509);
xnor U43117 (N_43117,N_42545,N_42702);
xor U43118 (N_43118,N_42317,N_42323);
and U43119 (N_43119,N_42748,N_42163);
xnor U43120 (N_43120,N_42863,N_42939);
xnor U43121 (N_43121,N_42676,N_42134);
xnor U43122 (N_43122,N_42056,N_42857);
or U43123 (N_43123,N_42528,N_42632);
and U43124 (N_43124,N_42320,N_42948);
nand U43125 (N_43125,N_42767,N_42722);
nor U43126 (N_43126,N_42120,N_42574);
or U43127 (N_43127,N_42628,N_42129);
and U43128 (N_43128,N_42136,N_42556);
and U43129 (N_43129,N_42783,N_42414);
and U43130 (N_43130,N_42677,N_42184);
nand U43131 (N_43131,N_42267,N_42401);
nand U43132 (N_43132,N_42378,N_42211);
or U43133 (N_43133,N_42203,N_42555);
or U43134 (N_43134,N_42406,N_42982);
nor U43135 (N_43135,N_42539,N_42849);
and U43136 (N_43136,N_42252,N_42165);
or U43137 (N_43137,N_42650,N_42151);
or U43138 (N_43138,N_42852,N_42904);
xor U43139 (N_43139,N_42707,N_42978);
or U43140 (N_43140,N_42075,N_42888);
nor U43141 (N_43141,N_42180,N_42660);
nor U43142 (N_43142,N_42034,N_42620);
or U43143 (N_43143,N_42347,N_42382);
xnor U43144 (N_43144,N_42780,N_42519);
and U43145 (N_43145,N_42132,N_42490);
nor U43146 (N_43146,N_42273,N_42150);
or U43147 (N_43147,N_42829,N_42839);
or U43148 (N_43148,N_42547,N_42405);
nor U43149 (N_43149,N_42410,N_42477);
and U43150 (N_43150,N_42280,N_42471);
nor U43151 (N_43151,N_42788,N_42614);
and U43152 (N_43152,N_42322,N_42031);
or U43153 (N_43153,N_42800,N_42430);
or U43154 (N_43154,N_42087,N_42155);
xnor U43155 (N_43155,N_42085,N_42095);
and U43156 (N_43156,N_42848,N_42993);
nor U43157 (N_43157,N_42011,N_42419);
nand U43158 (N_43158,N_42862,N_42061);
or U43159 (N_43159,N_42074,N_42815);
nand U43160 (N_43160,N_42488,N_42442);
nor U43161 (N_43161,N_42262,N_42753);
nor U43162 (N_43162,N_42461,N_42966);
nand U43163 (N_43163,N_42901,N_42673);
nor U43164 (N_43164,N_42072,N_42276);
and U43165 (N_43165,N_42256,N_42714);
nor U43166 (N_43166,N_42962,N_42591);
nand U43167 (N_43167,N_42732,N_42080);
and U43168 (N_43168,N_42804,N_42469);
or U43169 (N_43169,N_42853,N_42532);
nand U43170 (N_43170,N_42986,N_42586);
nor U43171 (N_43171,N_42661,N_42291);
or U43172 (N_43172,N_42444,N_42563);
nor U43173 (N_43173,N_42316,N_42486);
nor U43174 (N_43174,N_42268,N_42694);
nor U43175 (N_43175,N_42526,N_42230);
xor U43176 (N_43176,N_42980,N_42389);
nand U43177 (N_43177,N_42541,N_42437);
xor U43178 (N_43178,N_42634,N_42015);
nand U43179 (N_43179,N_42736,N_42782);
or U43180 (N_43180,N_42579,N_42938);
nand U43181 (N_43181,N_42250,N_42278);
nand U43182 (N_43182,N_42741,N_42647);
nand U43183 (N_43183,N_42612,N_42353);
nand U43184 (N_43184,N_42739,N_42395);
and U43185 (N_43185,N_42560,N_42914);
or U43186 (N_43186,N_42581,N_42452);
nand U43187 (N_43187,N_42943,N_42543);
or U43188 (N_43188,N_42351,N_42468);
or U43189 (N_43189,N_42188,N_42388);
or U43190 (N_43190,N_42417,N_42359);
xor U43191 (N_43191,N_42754,N_42657);
and U43192 (N_43192,N_42641,N_42544);
nor U43193 (N_43193,N_42149,N_42957);
and U43194 (N_43194,N_42623,N_42333);
or U43195 (N_43195,N_42124,N_42812);
or U43196 (N_43196,N_42073,N_42506);
and U43197 (N_43197,N_42053,N_42701);
and U43198 (N_43198,N_42209,N_42902);
or U43199 (N_43199,N_42858,N_42364);
and U43200 (N_43200,N_42048,N_42949);
nand U43201 (N_43201,N_42624,N_42215);
or U43202 (N_43202,N_42604,N_42060);
nand U43203 (N_43203,N_42152,N_42299);
nand U43204 (N_43204,N_42837,N_42988);
and U43205 (N_43205,N_42996,N_42176);
nor U43206 (N_43206,N_42619,N_42345);
and U43207 (N_43207,N_42128,N_42885);
nand U43208 (N_43208,N_42712,N_42537);
nor U43209 (N_43209,N_42953,N_42809);
xnor U43210 (N_43210,N_42717,N_42582);
xor U43211 (N_43211,N_42479,N_42766);
and U43212 (N_43212,N_42832,N_42697);
nor U43213 (N_43213,N_42318,N_42237);
xnor U43214 (N_43214,N_42141,N_42020);
xor U43215 (N_43215,N_42578,N_42045);
and U43216 (N_43216,N_42704,N_42992);
and U43217 (N_43217,N_42174,N_42599);
and U43218 (N_43218,N_42489,N_42285);
and U43219 (N_43219,N_42922,N_42502);
xnor U43220 (N_43220,N_42196,N_42874);
nor U43221 (N_43221,N_42238,N_42752);
and U43222 (N_43222,N_42336,N_42887);
nor U43223 (N_43223,N_42587,N_42861);
xnor U43224 (N_43224,N_42561,N_42446);
nor U43225 (N_43225,N_42022,N_42940);
and U43226 (N_43226,N_42231,N_42897);
nand U43227 (N_43227,N_42719,N_42173);
nor U43228 (N_43228,N_42972,N_42516);
and U43229 (N_43229,N_42841,N_42770);
xor U43230 (N_43230,N_42166,N_42598);
nor U43231 (N_43231,N_42615,N_42463);
xnor U43232 (N_43232,N_42212,N_42293);
nand U43233 (N_43233,N_42878,N_42495);
nor U43234 (N_43234,N_42205,N_42525);
xor U43235 (N_43235,N_42868,N_42112);
nor U43236 (N_43236,N_42738,N_42564);
or U43237 (N_43237,N_42458,N_42470);
xor U43238 (N_43238,N_42567,N_42844);
or U43239 (N_43239,N_42207,N_42600);
xor U43240 (N_43240,N_42626,N_42263);
and U43241 (N_43241,N_42021,N_42573);
and U43242 (N_43242,N_42913,N_42720);
and U43243 (N_43243,N_42816,N_42271);
or U43244 (N_43244,N_42253,N_42514);
xnor U43245 (N_43245,N_42050,N_42929);
xor U43246 (N_43246,N_42472,N_42808);
and U43247 (N_43247,N_42496,N_42313);
xor U43248 (N_43248,N_42281,N_42360);
nor U43249 (N_43249,N_42540,N_42096);
nor U43250 (N_43250,N_42255,N_42793);
or U43251 (N_43251,N_42342,N_42756);
nor U43252 (N_43252,N_42590,N_42029);
xor U43253 (N_43253,N_42920,N_42160);
nor U43254 (N_43254,N_42507,N_42670);
or U43255 (N_43255,N_42803,N_42523);
and U43256 (N_43256,N_42935,N_42308);
and U43257 (N_43257,N_42637,N_42482);
nand U43258 (N_43258,N_42379,N_42908);
or U43259 (N_43259,N_42259,N_42251);
and U43260 (N_43260,N_42533,N_42358);
nor U43261 (N_43261,N_42190,N_42216);
and U43262 (N_43262,N_42715,N_42270);
xor U43263 (N_43263,N_42441,N_42091);
and U43264 (N_43264,N_42484,N_42017);
or U43265 (N_43265,N_42552,N_42065);
nand U43266 (N_43266,N_42485,N_42478);
nand U43267 (N_43267,N_42568,N_42608);
nor U43268 (N_43268,N_42955,N_42674);
and U43269 (N_43269,N_42778,N_42297);
xor U43270 (N_43270,N_42971,N_42208);
xnor U43271 (N_43271,N_42290,N_42453);
and U43272 (N_43272,N_42546,N_42726);
and U43273 (N_43273,N_42000,N_42036);
or U43274 (N_43274,N_42696,N_42372);
and U43275 (N_43275,N_42603,N_42531);
or U43276 (N_43276,N_42135,N_42755);
or U43277 (N_43277,N_42402,N_42282);
xor U43278 (N_43278,N_42630,N_42344);
nor U43279 (N_43279,N_42433,N_42123);
nand U43280 (N_43280,N_42369,N_42497);
nand U43281 (N_43281,N_42973,N_42636);
nand U43282 (N_43282,N_42622,N_42279);
xnor U43283 (N_43283,N_42368,N_42900);
xnor U43284 (N_43284,N_42328,N_42693);
or U43285 (N_43285,N_42936,N_42192);
xnor U43286 (N_43286,N_42261,N_42881);
and U43287 (N_43287,N_42451,N_42447);
nor U43288 (N_43288,N_42233,N_42295);
nand U43289 (N_43289,N_42423,N_42367);
nand U43290 (N_43290,N_42889,N_42505);
and U43291 (N_43291,N_42148,N_42856);
nor U43292 (N_43292,N_42325,N_42004);
or U43293 (N_43293,N_42965,N_42092);
xnor U43294 (N_43294,N_42146,N_42277);
nor U43295 (N_43295,N_42662,N_42055);
xor U43296 (N_43296,N_42906,N_42286);
and U43297 (N_43297,N_42896,N_42408);
or U43298 (N_43298,N_42042,N_42927);
and U43299 (N_43299,N_42666,N_42241);
nor U43300 (N_43300,N_42975,N_42139);
xnor U43301 (N_43301,N_42730,N_42535);
or U43302 (N_43302,N_42580,N_42569);
or U43303 (N_43303,N_42681,N_42529);
or U43304 (N_43304,N_42845,N_42548);
and U43305 (N_43305,N_42520,N_42562);
xor U43306 (N_43306,N_42254,N_42595);
or U43307 (N_43307,N_42698,N_42117);
nand U43308 (N_43308,N_42558,N_42133);
nand U43309 (N_43309,N_42718,N_42799);
nor U43310 (N_43310,N_42457,N_42796);
and U43311 (N_43311,N_42186,N_42170);
nand U43312 (N_43312,N_42515,N_42081);
nor U43313 (N_43313,N_42983,N_42137);
or U43314 (N_43314,N_42028,N_42700);
nand U43315 (N_43315,N_42870,N_42284);
and U43316 (N_43316,N_42798,N_42138);
nor U43317 (N_43317,N_42393,N_42536);
and U43318 (N_43318,N_42654,N_42426);
or U43319 (N_43319,N_42043,N_42008);
and U43320 (N_43320,N_42880,N_42524);
xor U43321 (N_43321,N_42768,N_42629);
xor U43322 (N_43322,N_42391,N_42784);
nor U43323 (N_43323,N_42033,N_42797);
nand U43324 (N_43324,N_42269,N_42968);
xnor U43325 (N_43325,N_42049,N_42355);
nand U43326 (N_43326,N_42371,N_42932);
nand U43327 (N_43327,N_42454,N_42104);
nor U43328 (N_43328,N_42396,N_42842);
nand U43329 (N_43329,N_42481,N_42503);
nand U43330 (N_43330,N_42067,N_42984);
nor U43331 (N_43331,N_42460,N_42836);
and U43332 (N_43332,N_42465,N_42669);
and U43333 (N_43333,N_42298,N_42706);
xnor U43334 (N_43334,N_42283,N_42399);
or U43335 (N_43335,N_42172,N_42024);
nor U43336 (N_43336,N_42189,N_42501);
nor U43337 (N_43337,N_42439,N_42950);
and U43338 (N_43338,N_42671,N_42292);
or U43339 (N_43339,N_42064,N_42198);
and U43340 (N_43340,N_42377,N_42428);
nor U43341 (N_43341,N_42145,N_42387);
or U43342 (N_43342,N_42855,N_42642);
or U43343 (N_43343,N_42232,N_42449);
nand U43344 (N_43344,N_42821,N_42923);
or U43345 (N_43345,N_42527,N_42288);
nand U43346 (N_43346,N_42001,N_42571);
or U43347 (N_43347,N_42220,N_42306);
xnor U43348 (N_43348,N_42115,N_42365);
xnor U43349 (N_43349,N_42542,N_42942);
and U43350 (N_43350,N_42014,N_42329);
nor U43351 (N_43351,N_42850,N_42421);
xnor U43352 (N_43352,N_42871,N_42822);
and U43353 (N_43353,N_42937,N_42390);
nand U43354 (N_43354,N_42309,N_42958);
or U43355 (N_43355,N_42977,N_42551);
and U43356 (N_43356,N_42301,N_42483);
xor U43357 (N_43357,N_42302,N_42589);
xor U43358 (N_43358,N_42883,N_42840);
and U43359 (N_43359,N_42692,N_42403);
and U43360 (N_43360,N_42792,N_42493);
and U43361 (N_43361,N_42663,N_42147);
xor U43362 (N_43362,N_42775,N_42206);
xnor U43363 (N_43363,N_42969,N_42200);
xor U43364 (N_43364,N_42265,N_42040);
or U43365 (N_43365,N_42510,N_42774);
nand U43366 (N_43366,N_42443,N_42027);
or U43367 (N_43367,N_42431,N_42113);
nor U43368 (N_43368,N_42781,N_42385);
nand U43369 (N_43369,N_42491,N_42337);
nor U43370 (N_43370,N_42987,N_42751);
or U43371 (N_43371,N_42376,N_42708);
nor U43372 (N_43372,N_42689,N_42090);
or U43373 (N_43373,N_42789,N_42761);
nor U43374 (N_43374,N_42400,N_42161);
and U43375 (N_43375,N_42063,N_42164);
nand U43376 (N_43376,N_42759,N_42833);
nor U43377 (N_43377,N_42828,N_42397);
or U43378 (N_43378,N_42362,N_42776);
nor U43379 (N_43379,N_42366,N_42791);
and U43380 (N_43380,N_42311,N_42592);
xor U43381 (N_43381,N_42032,N_42765);
or U43382 (N_43382,N_42790,N_42854);
xnor U43383 (N_43383,N_42802,N_42304);
or U43384 (N_43384,N_42633,N_42415);
nand U43385 (N_43385,N_42144,N_42383);
xor U43386 (N_43386,N_42758,N_42917);
xor U43387 (N_43387,N_42236,N_42864);
xnor U43388 (N_43388,N_42865,N_42737);
and U43389 (N_43389,N_42979,N_42257);
or U43390 (N_43390,N_42734,N_42370);
or U43391 (N_43391,N_42724,N_42338);
nor U43392 (N_43392,N_42757,N_42576);
nor U43393 (N_43393,N_42974,N_42709);
nor U43394 (N_43394,N_42721,N_42944);
and U43395 (N_43395,N_42210,N_42006);
or U43396 (N_43396,N_42699,N_42991);
and U43397 (N_43397,N_42667,N_42054);
nand U43398 (N_43398,N_42162,N_42616);
and U43399 (N_43399,N_42440,N_42424);
and U43400 (N_43400,N_42127,N_42686);
xnor U43401 (N_43401,N_42688,N_42648);
nand U43402 (N_43402,N_42314,N_42649);
and U43403 (N_43403,N_42565,N_42764);
nor U43404 (N_43404,N_42182,N_42374);
nand U43405 (N_43405,N_42289,N_42204);
and U43406 (N_43406,N_42101,N_42687);
and U43407 (N_43407,N_42287,N_42106);
xor U43408 (N_43408,N_42511,N_42585);
and U43409 (N_43409,N_42214,N_42640);
xnor U43410 (N_43410,N_42843,N_42918);
or U43411 (N_43411,N_42892,N_42899);
or U43412 (N_43412,N_42665,N_42613);
nor U43413 (N_43413,N_42350,N_42818);
and U43414 (N_43414,N_42429,N_42221);
or U43415 (N_43415,N_42659,N_42785);
xor U43416 (N_43416,N_42672,N_42416);
xor U43417 (N_43417,N_42143,N_42678);
nor U43418 (N_43418,N_42384,N_42746);
nor U43419 (N_43419,N_42079,N_42572);
or U43420 (N_43420,N_42611,N_42418);
nand U43421 (N_43421,N_42771,N_42508);
nor U43422 (N_43422,N_42264,N_42407);
or U43423 (N_43423,N_42343,N_42682);
nand U43424 (N_43424,N_42197,N_42083);
nand U43425 (N_43425,N_42625,N_42710);
nor U43426 (N_43426,N_42357,N_42869);
or U43427 (N_43427,N_42294,N_42684);
xor U43428 (N_43428,N_42744,N_42813);
xor U43429 (N_43429,N_42005,N_42312);
nor U43430 (N_43430,N_42976,N_42827);
and U43431 (N_43431,N_42324,N_42078);
nand U43432 (N_43432,N_42436,N_42070);
xor U43433 (N_43433,N_42363,N_42111);
and U43434 (N_43434,N_42224,N_42057);
nor U43435 (N_43435,N_42413,N_42947);
nand U43436 (N_43436,N_42275,N_42199);
or U43437 (N_43437,N_42326,N_42118);
and U43438 (N_43438,N_42905,N_42606);
and U43439 (N_43439,N_42373,N_42239);
or U43440 (N_43440,N_42727,N_42093);
nand U43441 (N_43441,N_42859,N_42512);
xor U43442 (N_43442,N_42893,N_42244);
nand U43443 (N_43443,N_42130,N_42725);
or U43444 (N_43444,N_42779,N_42963);
or U43445 (N_43445,N_42013,N_42218);
nor U43446 (N_43446,N_42601,N_42745);
xor U43447 (N_43447,N_42749,N_42226);
xor U43448 (N_43448,N_42380,N_42882);
nand U43449 (N_43449,N_42023,N_42680);
nand U43450 (N_43450,N_42675,N_42222);
or U43451 (N_43451,N_42381,N_42175);
or U43452 (N_43452,N_42500,N_42094);
or U43453 (N_43453,N_42522,N_42886);
nor U43454 (N_43454,N_42159,N_42114);
or U43455 (N_43455,N_42814,N_42959);
or U43456 (N_43456,N_42088,N_42487);
nand U43457 (N_43457,N_42100,N_42743);
xnor U43458 (N_43458,N_42597,N_42217);
nor U43459 (N_43459,N_42656,N_42077);
or U43460 (N_43460,N_42655,N_42435);
or U43461 (N_43461,N_42327,N_42891);
or U43462 (N_43462,N_42933,N_42109);
nand U43463 (N_43463,N_42826,N_42361);
or U43464 (N_43464,N_42530,N_42499);
xnor U43465 (N_43465,N_42643,N_42319);
nand U43466 (N_43466,N_42068,N_42998);
or U43467 (N_43467,N_42884,N_42434);
and U43468 (N_43468,N_42817,N_42652);
nor U43469 (N_43469,N_42825,N_42521);
nand U43470 (N_43470,N_42235,N_42602);
or U43471 (N_43471,N_42195,N_42557);
nor U43472 (N_43472,N_42018,N_42605);
and U43473 (N_43473,N_42860,N_42116);
nand U43474 (N_43474,N_42248,N_42227);
and U43475 (N_43475,N_42847,N_42455);
nand U43476 (N_43476,N_42069,N_42777);
nand U43477 (N_43477,N_42121,N_42110);
nor U43478 (N_43478,N_42644,N_42475);
and U43479 (N_43479,N_42346,N_42534);
and U43480 (N_43480,N_42713,N_42386);
xor U43481 (N_43481,N_42462,N_42219);
nor U43482 (N_43482,N_42945,N_42303);
or U43483 (N_43483,N_42178,N_42076);
xnor U43484 (N_43484,N_42794,N_42474);
or U43485 (N_43485,N_42760,N_42716);
xor U43486 (N_43486,N_42867,N_42806);
nand U43487 (N_43487,N_42733,N_42909);
xor U43488 (N_43488,N_42183,N_42679);
xor U43489 (N_43489,N_42877,N_42404);
xor U43490 (N_43490,N_42356,N_42009);
xor U43491 (N_43491,N_42229,N_42513);
and U43492 (N_43492,N_42274,N_42954);
or U43493 (N_43493,N_42052,N_42851);
nor U43494 (N_43494,N_42007,N_42003);
nand U43495 (N_43495,N_42082,N_42466);
nand U43496 (N_43496,N_42961,N_42907);
nor U43497 (N_43497,N_42872,N_42107);
nand U43498 (N_43498,N_42335,N_42668);
nor U43499 (N_43499,N_42538,N_42890);
xor U43500 (N_43500,N_42539,N_42659);
and U43501 (N_43501,N_42932,N_42907);
and U43502 (N_43502,N_42807,N_42696);
and U43503 (N_43503,N_42364,N_42662);
nor U43504 (N_43504,N_42132,N_42476);
and U43505 (N_43505,N_42562,N_42583);
nor U43506 (N_43506,N_42367,N_42177);
nand U43507 (N_43507,N_42225,N_42840);
xor U43508 (N_43508,N_42413,N_42853);
xor U43509 (N_43509,N_42316,N_42867);
and U43510 (N_43510,N_42718,N_42236);
and U43511 (N_43511,N_42925,N_42270);
or U43512 (N_43512,N_42153,N_42303);
xnor U43513 (N_43513,N_42750,N_42786);
or U43514 (N_43514,N_42679,N_42665);
and U43515 (N_43515,N_42915,N_42823);
xor U43516 (N_43516,N_42453,N_42049);
or U43517 (N_43517,N_42770,N_42508);
and U43518 (N_43518,N_42714,N_42463);
or U43519 (N_43519,N_42250,N_42084);
or U43520 (N_43520,N_42943,N_42770);
nor U43521 (N_43521,N_42612,N_42821);
nor U43522 (N_43522,N_42520,N_42796);
or U43523 (N_43523,N_42060,N_42946);
nor U43524 (N_43524,N_42395,N_42574);
nor U43525 (N_43525,N_42393,N_42921);
nor U43526 (N_43526,N_42477,N_42155);
xnor U43527 (N_43527,N_42587,N_42916);
xnor U43528 (N_43528,N_42823,N_42015);
or U43529 (N_43529,N_42483,N_42867);
nor U43530 (N_43530,N_42828,N_42734);
xnor U43531 (N_43531,N_42587,N_42758);
nor U43532 (N_43532,N_42561,N_42229);
nor U43533 (N_43533,N_42582,N_42787);
xor U43534 (N_43534,N_42239,N_42001);
xor U43535 (N_43535,N_42479,N_42460);
and U43536 (N_43536,N_42887,N_42745);
or U43537 (N_43537,N_42662,N_42743);
and U43538 (N_43538,N_42856,N_42044);
nor U43539 (N_43539,N_42986,N_42420);
xnor U43540 (N_43540,N_42294,N_42043);
and U43541 (N_43541,N_42094,N_42197);
nor U43542 (N_43542,N_42143,N_42457);
and U43543 (N_43543,N_42525,N_42845);
nor U43544 (N_43544,N_42757,N_42040);
or U43545 (N_43545,N_42470,N_42750);
and U43546 (N_43546,N_42679,N_42601);
or U43547 (N_43547,N_42313,N_42733);
nor U43548 (N_43548,N_42211,N_42891);
nor U43549 (N_43549,N_42518,N_42351);
or U43550 (N_43550,N_42359,N_42749);
and U43551 (N_43551,N_42856,N_42037);
xor U43552 (N_43552,N_42272,N_42346);
xnor U43553 (N_43553,N_42671,N_42659);
and U43554 (N_43554,N_42644,N_42278);
and U43555 (N_43555,N_42696,N_42358);
xor U43556 (N_43556,N_42690,N_42547);
nand U43557 (N_43557,N_42761,N_42152);
nor U43558 (N_43558,N_42306,N_42674);
nor U43559 (N_43559,N_42643,N_42446);
and U43560 (N_43560,N_42205,N_42962);
and U43561 (N_43561,N_42894,N_42957);
xor U43562 (N_43562,N_42491,N_42611);
and U43563 (N_43563,N_42998,N_42016);
nand U43564 (N_43564,N_42570,N_42811);
nor U43565 (N_43565,N_42911,N_42020);
xnor U43566 (N_43566,N_42758,N_42719);
xor U43567 (N_43567,N_42587,N_42569);
xor U43568 (N_43568,N_42654,N_42607);
nor U43569 (N_43569,N_42663,N_42091);
nor U43570 (N_43570,N_42075,N_42228);
nor U43571 (N_43571,N_42677,N_42030);
nor U43572 (N_43572,N_42185,N_42059);
nand U43573 (N_43573,N_42073,N_42011);
nor U43574 (N_43574,N_42611,N_42449);
nand U43575 (N_43575,N_42278,N_42269);
xor U43576 (N_43576,N_42360,N_42548);
and U43577 (N_43577,N_42287,N_42507);
and U43578 (N_43578,N_42862,N_42304);
nor U43579 (N_43579,N_42211,N_42209);
or U43580 (N_43580,N_42881,N_42144);
nor U43581 (N_43581,N_42298,N_42217);
nand U43582 (N_43582,N_42115,N_42253);
nand U43583 (N_43583,N_42183,N_42322);
or U43584 (N_43584,N_42034,N_42130);
xnor U43585 (N_43585,N_42852,N_42930);
xor U43586 (N_43586,N_42879,N_42099);
and U43587 (N_43587,N_42937,N_42025);
nor U43588 (N_43588,N_42593,N_42431);
or U43589 (N_43589,N_42047,N_42466);
nor U43590 (N_43590,N_42344,N_42474);
and U43591 (N_43591,N_42686,N_42419);
nand U43592 (N_43592,N_42544,N_42946);
nor U43593 (N_43593,N_42817,N_42658);
or U43594 (N_43594,N_42672,N_42794);
or U43595 (N_43595,N_42259,N_42506);
or U43596 (N_43596,N_42090,N_42527);
xor U43597 (N_43597,N_42447,N_42273);
or U43598 (N_43598,N_42506,N_42251);
or U43599 (N_43599,N_42252,N_42568);
and U43600 (N_43600,N_42135,N_42027);
nor U43601 (N_43601,N_42599,N_42114);
nand U43602 (N_43602,N_42548,N_42988);
nand U43603 (N_43603,N_42008,N_42180);
and U43604 (N_43604,N_42956,N_42266);
nand U43605 (N_43605,N_42533,N_42297);
nor U43606 (N_43606,N_42210,N_42565);
xnor U43607 (N_43607,N_42630,N_42723);
xnor U43608 (N_43608,N_42767,N_42840);
nand U43609 (N_43609,N_42567,N_42340);
nand U43610 (N_43610,N_42751,N_42055);
nor U43611 (N_43611,N_42393,N_42696);
xor U43612 (N_43612,N_42110,N_42204);
xor U43613 (N_43613,N_42820,N_42911);
and U43614 (N_43614,N_42315,N_42825);
xor U43615 (N_43615,N_42819,N_42365);
and U43616 (N_43616,N_42014,N_42982);
xor U43617 (N_43617,N_42321,N_42830);
nand U43618 (N_43618,N_42769,N_42184);
nand U43619 (N_43619,N_42133,N_42104);
nand U43620 (N_43620,N_42349,N_42631);
and U43621 (N_43621,N_42047,N_42032);
nand U43622 (N_43622,N_42667,N_42763);
nand U43623 (N_43623,N_42033,N_42929);
xor U43624 (N_43624,N_42564,N_42584);
nand U43625 (N_43625,N_42645,N_42968);
and U43626 (N_43626,N_42468,N_42008);
nor U43627 (N_43627,N_42810,N_42455);
xor U43628 (N_43628,N_42255,N_42328);
xor U43629 (N_43629,N_42639,N_42584);
and U43630 (N_43630,N_42163,N_42144);
nor U43631 (N_43631,N_42973,N_42989);
or U43632 (N_43632,N_42230,N_42464);
nor U43633 (N_43633,N_42359,N_42696);
or U43634 (N_43634,N_42168,N_42050);
nand U43635 (N_43635,N_42714,N_42095);
nand U43636 (N_43636,N_42752,N_42129);
or U43637 (N_43637,N_42739,N_42093);
and U43638 (N_43638,N_42582,N_42743);
nor U43639 (N_43639,N_42549,N_42649);
xor U43640 (N_43640,N_42684,N_42614);
xor U43641 (N_43641,N_42399,N_42969);
or U43642 (N_43642,N_42314,N_42647);
or U43643 (N_43643,N_42648,N_42462);
xnor U43644 (N_43644,N_42353,N_42175);
or U43645 (N_43645,N_42088,N_42537);
nor U43646 (N_43646,N_42138,N_42942);
nor U43647 (N_43647,N_42866,N_42005);
xor U43648 (N_43648,N_42860,N_42662);
nor U43649 (N_43649,N_42585,N_42467);
nor U43650 (N_43650,N_42554,N_42307);
xor U43651 (N_43651,N_42777,N_42320);
xnor U43652 (N_43652,N_42971,N_42425);
or U43653 (N_43653,N_42995,N_42939);
nor U43654 (N_43654,N_42705,N_42442);
or U43655 (N_43655,N_42347,N_42637);
xor U43656 (N_43656,N_42547,N_42554);
or U43657 (N_43657,N_42354,N_42227);
or U43658 (N_43658,N_42808,N_42894);
xnor U43659 (N_43659,N_42756,N_42811);
and U43660 (N_43660,N_42296,N_42098);
and U43661 (N_43661,N_42450,N_42563);
xor U43662 (N_43662,N_42837,N_42941);
nor U43663 (N_43663,N_42692,N_42189);
and U43664 (N_43664,N_42494,N_42809);
or U43665 (N_43665,N_42318,N_42676);
nand U43666 (N_43666,N_42709,N_42786);
and U43667 (N_43667,N_42939,N_42778);
nor U43668 (N_43668,N_42244,N_42875);
and U43669 (N_43669,N_42284,N_42967);
xnor U43670 (N_43670,N_42137,N_42010);
nor U43671 (N_43671,N_42684,N_42538);
nand U43672 (N_43672,N_42414,N_42604);
and U43673 (N_43673,N_42467,N_42383);
and U43674 (N_43674,N_42726,N_42628);
xnor U43675 (N_43675,N_42428,N_42471);
nand U43676 (N_43676,N_42189,N_42412);
or U43677 (N_43677,N_42434,N_42630);
or U43678 (N_43678,N_42920,N_42906);
xnor U43679 (N_43679,N_42254,N_42630);
nand U43680 (N_43680,N_42807,N_42658);
nor U43681 (N_43681,N_42873,N_42483);
nand U43682 (N_43682,N_42735,N_42200);
nand U43683 (N_43683,N_42509,N_42682);
or U43684 (N_43684,N_42884,N_42615);
xnor U43685 (N_43685,N_42684,N_42493);
xor U43686 (N_43686,N_42976,N_42742);
and U43687 (N_43687,N_42763,N_42664);
and U43688 (N_43688,N_42497,N_42141);
nand U43689 (N_43689,N_42553,N_42243);
nand U43690 (N_43690,N_42266,N_42407);
nor U43691 (N_43691,N_42500,N_42499);
nor U43692 (N_43692,N_42757,N_42923);
nand U43693 (N_43693,N_42967,N_42879);
or U43694 (N_43694,N_42977,N_42597);
and U43695 (N_43695,N_42269,N_42351);
nor U43696 (N_43696,N_42577,N_42910);
nand U43697 (N_43697,N_42383,N_42292);
or U43698 (N_43698,N_42850,N_42380);
xnor U43699 (N_43699,N_42455,N_42987);
nand U43700 (N_43700,N_42416,N_42932);
nand U43701 (N_43701,N_42391,N_42708);
xnor U43702 (N_43702,N_42604,N_42127);
and U43703 (N_43703,N_42899,N_42310);
or U43704 (N_43704,N_42765,N_42086);
xnor U43705 (N_43705,N_42259,N_42072);
and U43706 (N_43706,N_42534,N_42749);
and U43707 (N_43707,N_42920,N_42631);
nand U43708 (N_43708,N_42900,N_42320);
or U43709 (N_43709,N_42974,N_42232);
or U43710 (N_43710,N_42190,N_42737);
or U43711 (N_43711,N_42304,N_42207);
xnor U43712 (N_43712,N_42630,N_42535);
xor U43713 (N_43713,N_42399,N_42741);
xnor U43714 (N_43714,N_42597,N_42599);
or U43715 (N_43715,N_42836,N_42341);
nand U43716 (N_43716,N_42188,N_42369);
xor U43717 (N_43717,N_42774,N_42265);
nor U43718 (N_43718,N_42593,N_42719);
or U43719 (N_43719,N_42200,N_42461);
nand U43720 (N_43720,N_42743,N_42402);
nor U43721 (N_43721,N_42696,N_42382);
nor U43722 (N_43722,N_42881,N_42964);
nand U43723 (N_43723,N_42398,N_42320);
xor U43724 (N_43724,N_42105,N_42492);
nand U43725 (N_43725,N_42442,N_42618);
nor U43726 (N_43726,N_42875,N_42441);
nand U43727 (N_43727,N_42490,N_42484);
nor U43728 (N_43728,N_42555,N_42757);
xor U43729 (N_43729,N_42089,N_42474);
nand U43730 (N_43730,N_42087,N_42946);
and U43731 (N_43731,N_42914,N_42911);
and U43732 (N_43732,N_42851,N_42105);
or U43733 (N_43733,N_42283,N_42437);
and U43734 (N_43734,N_42068,N_42393);
nor U43735 (N_43735,N_42651,N_42416);
xor U43736 (N_43736,N_42775,N_42754);
nor U43737 (N_43737,N_42324,N_42977);
xnor U43738 (N_43738,N_42302,N_42819);
or U43739 (N_43739,N_42314,N_42390);
xnor U43740 (N_43740,N_42380,N_42236);
nand U43741 (N_43741,N_42662,N_42554);
and U43742 (N_43742,N_42539,N_42280);
and U43743 (N_43743,N_42418,N_42529);
or U43744 (N_43744,N_42237,N_42827);
nand U43745 (N_43745,N_42425,N_42521);
nor U43746 (N_43746,N_42103,N_42235);
nor U43747 (N_43747,N_42629,N_42104);
or U43748 (N_43748,N_42875,N_42693);
nand U43749 (N_43749,N_42888,N_42556);
nor U43750 (N_43750,N_42717,N_42536);
or U43751 (N_43751,N_42244,N_42498);
nor U43752 (N_43752,N_42609,N_42080);
xor U43753 (N_43753,N_42626,N_42435);
or U43754 (N_43754,N_42404,N_42763);
nor U43755 (N_43755,N_42610,N_42396);
xnor U43756 (N_43756,N_42119,N_42742);
nand U43757 (N_43757,N_42678,N_42725);
nor U43758 (N_43758,N_42296,N_42999);
nor U43759 (N_43759,N_42224,N_42198);
nand U43760 (N_43760,N_42285,N_42817);
and U43761 (N_43761,N_42941,N_42670);
or U43762 (N_43762,N_42682,N_42002);
nor U43763 (N_43763,N_42546,N_42156);
and U43764 (N_43764,N_42824,N_42259);
or U43765 (N_43765,N_42335,N_42832);
nand U43766 (N_43766,N_42616,N_42852);
nand U43767 (N_43767,N_42620,N_42022);
nand U43768 (N_43768,N_42729,N_42053);
or U43769 (N_43769,N_42981,N_42091);
nor U43770 (N_43770,N_42407,N_42817);
and U43771 (N_43771,N_42067,N_42187);
and U43772 (N_43772,N_42709,N_42981);
and U43773 (N_43773,N_42205,N_42164);
xor U43774 (N_43774,N_42441,N_42209);
nor U43775 (N_43775,N_42099,N_42250);
or U43776 (N_43776,N_42748,N_42852);
xnor U43777 (N_43777,N_42594,N_42809);
nor U43778 (N_43778,N_42238,N_42746);
xnor U43779 (N_43779,N_42881,N_42632);
or U43780 (N_43780,N_42470,N_42087);
nand U43781 (N_43781,N_42394,N_42508);
nand U43782 (N_43782,N_42612,N_42288);
nand U43783 (N_43783,N_42177,N_42990);
nor U43784 (N_43784,N_42059,N_42010);
xnor U43785 (N_43785,N_42595,N_42144);
nor U43786 (N_43786,N_42379,N_42983);
xor U43787 (N_43787,N_42847,N_42713);
and U43788 (N_43788,N_42574,N_42164);
xor U43789 (N_43789,N_42071,N_42615);
xnor U43790 (N_43790,N_42454,N_42485);
and U43791 (N_43791,N_42040,N_42748);
nor U43792 (N_43792,N_42883,N_42495);
nand U43793 (N_43793,N_42966,N_42980);
and U43794 (N_43794,N_42348,N_42578);
xnor U43795 (N_43795,N_42433,N_42575);
xor U43796 (N_43796,N_42097,N_42982);
nor U43797 (N_43797,N_42156,N_42908);
nand U43798 (N_43798,N_42951,N_42409);
nor U43799 (N_43799,N_42623,N_42327);
xnor U43800 (N_43800,N_42495,N_42619);
nor U43801 (N_43801,N_42507,N_42042);
or U43802 (N_43802,N_42958,N_42738);
and U43803 (N_43803,N_42668,N_42967);
or U43804 (N_43804,N_42277,N_42298);
or U43805 (N_43805,N_42496,N_42472);
xor U43806 (N_43806,N_42197,N_42023);
or U43807 (N_43807,N_42011,N_42353);
nand U43808 (N_43808,N_42866,N_42521);
nand U43809 (N_43809,N_42879,N_42268);
and U43810 (N_43810,N_42517,N_42279);
or U43811 (N_43811,N_42286,N_42123);
xnor U43812 (N_43812,N_42327,N_42381);
nor U43813 (N_43813,N_42531,N_42798);
nor U43814 (N_43814,N_42509,N_42081);
or U43815 (N_43815,N_42257,N_42595);
nor U43816 (N_43816,N_42351,N_42427);
or U43817 (N_43817,N_42691,N_42228);
or U43818 (N_43818,N_42236,N_42351);
and U43819 (N_43819,N_42130,N_42976);
nor U43820 (N_43820,N_42075,N_42648);
nor U43821 (N_43821,N_42757,N_42789);
or U43822 (N_43822,N_42804,N_42656);
nor U43823 (N_43823,N_42509,N_42315);
nor U43824 (N_43824,N_42205,N_42654);
nor U43825 (N_43825,N_42391,N_42153);
xor U43826 (N_43826,N_42230,N_42125);
nor U43827 (N_43827,N_42872,N_42812);
nor U43828 (N_43828,N_42662,N_42302);
nor U43829 (N_43829,N_42879,N_42197);
xor U43830 (N_43830,N_42274,N_42814);
nor U43831 (N_43831,N_42736,N_42194);
nor U43832 (N_43832,N_42775,N_42847);
and U43833 (N_43833,N_42256,N_42546);
nand U43834 (N_43834,N_42107,N_42744);
nor U43835 (N_43835,N_42402,N_42549);
xor U43836 (N_43836,N_42932,N_42941);
xnor U43837 (N_43837,N_42043,N_42239);
or U43838 (N_43838,N_42074,N_42699);
and U43839 (N_43839,N_42748,N_42892);
or U43840 (N_43840,N_42168,N_42707);
xor U43841 (N_43841,N_42039,N_42788);
nand U43842 (N_43842,N_42006,N_42329);
nor U43843 (N_43843,N_42650,N_42622);
or U43844 (N_43844,N_42101,N_42142);
and U43845 (N_43845,N_42394,N_42535);
nor U43846 (N_43846,N_42737,N_42113);
or U43847 (N_43847,N_42652,N_42891);
nand U43848 (N_43848,N_42871,N_42708);
or U43849 (N_43849,N_42549,N_42729);
and U43850 (N_43850,N_42521,N_42506);
nor U43851 (N_43851,N_42966,N_42592);
or U43852 (N_43852,N_42255,N_42002);
nand U43853 (N_43853,N_42553,N_42374);
and U43854 (N_43854,N_42076,N_42921);
xor U43855 (N_43855,N_42704,N_42947);
and U43856 (N_43856,N_42383,N_42918);
nand U43857 (N_43857,N_42452,N_42140);
and U43858 (N_43858,N_42340,N_42225);
and U43859 (N_43859,N_42948,N_42934);
nor U43860 (N_43860,N_42016,N_42690);
xor U43861 (N_43861,N_42356,N_42580);
xnor U43862 (N_43862,N_42860,N_42696);
or U43863 (N_43863,N_42415,N_42314);
and U43864 (N_43864,N_42263,N_42679);
and U43865 (N_43865,N_42638,N_42575);
xnor U43866 (N_43866,N_42092,N_42602);
or U43867 (N_43867,N_42297,N_42751);
nand U43868 (N_43868,N_42149,N_42706);
or U43869 (N_43869,N_42516,N_42913);
or U43870 (N_43870,N_42936,N_42734);
xor U43871 (N_43871,N_42571,N_42753);
and U43872 (N_43872,N_42185,N_42330);
xor U43873 (N_43873,N_42464,N_42706);
xnor U43874 (N_43874,N_42845,N_42641);
or U43875 (N_43875,N_42718,N_42707);
nand U43876 (N_43876,N_42532,N_42079);
nor U43877 (N_43877,N_42104,N_42189);
or U43878 (N_43878,N_42283,N_42087);
or U43879 (N_43879,N_42600,N_42274);
xor U43880 (N_43880,N_42169,N_42633);
nor U43881 (N_43881,N_42834,N_42169);
nor U43882 (N_43882,N_42481,N_42836);
or U43883 (N_43883,N_42076,N_42662);
and U43884 (N_43884,N_42362,N_42113);
and U43885 (N_43885,N_42932,N_42048);
or U43886 (N_43886,N_42048,N_42032);
xnor U43887 (N_43887,N_42738,N_42775);
nor U43888 (N_43888,N_42395,N_42223);
nand U43889 (N_43889,N_42394,N_42250);
and U43890 (N_43890,N_42383,N_42595);
nand U43891 (N_43891,N_42509,N_42829);
and U43892 (N_43892,N_42687,N_42660);
nor U43893 (N_43893,N_42399,N_42143);
xnor U43894 (N_43894,N_42866,N_42532);
and U43895 (N_43895,N_42116,N_42290);
and U43896 (N_43896,N_42144,N_42031);
nor U43897 (N_43897,N_42742,N_42917);
xor U43898 (N_43898,N_42769,N_42470);
nor U43899 (N_43899,N_42193,N_42727);
nand U43900 (N_43900,N_42347,N_42231);
xnor U43901 (N_43901,N_42536,N_42615);
nor U43902 (N_43902,N_42598,N_42264);
and U43903 (N_43903,N_42839,N_42000);
nand U43904 (N_43904,N_42972,N_42628);
and U43905 (N_43905,N_42246,N_42735);
nor U43906 (N_43906,N_42661,N_42930);
xnor U43907 (N_43907,N_42469,N_42889);
nand U43908 (N_43908,N_42228,N_42450);
nor U43909 (N_43909,N_42214,N_42911);
nand U43910 (N_43910,N_42697,N_42948);
xor U43911 (N_43911,N_42072,N_42656);
or U43912 (N_43912,N_42736,N_42246);
or U43913 (N_43913,N_42391,N_42400);
and U43914 (N_43914,N_42173,N_42661);
and U43915 (N_43915,N_42756,N_42443);
xor U43916 (N_43916,N_42210,N_42962);
and U43917 (N_43917,N_42211,N_42138);
xor U43918 (N_43918,N_42264,N_42845);
xor U43919 (N_43919,N_42694,N_42600);
xor U43920 (N_43920,N_42477,N_42306);
nand U43921 (N_43921,N_42617,N_42599);
nor U43922 (N_43922,N_42798,N_42665);
nor U43923 (N_43923,N_42720,N_42786);
and U43924 (N_43924,N_42030,N_42850);
nor U43925 (N_43925,N_42002,N_42521);
nand U43926 (N_43926,N_42391,N_42254);
nor U43927 (N_43927,N_42753,N_42237);
or U43928 (N_43928,N_42843,N_42489);
xnor U43929 (N_43929,N_42226,N_42378);
nor U43930 (N_43930,N_42660,N_42278);
or U43931 (N_43931,N_42994,N_42017);
xnor U43932 (N_43932,N_42685,N_42631);
nor U43933 (N_43933,N_42667,N_42425);
nand U43934 (N_43934,N_42079,N_42693);
or U43935 (N_43935,N_42671,N_42807);
xor U43936 (N_43936,N_42810,N_42548);
xor U43937 (N_43937,N_42036,N_42523);
nor U43938 (N_43938,N_42547,N_42129);
and U43939 (N_43939,N_42485,N_42880);
or U43940 (N_43940,N_42282,N_42561);
nor U43941 (N_43941,N_42452,N_42216);
nor U43942 (N_43942,N_42195,N_42111);
nand U43943 (N_43943,N_42614,N_42450);
xor U43944 (N_43944,N_42370,N_42314);
xor U43945 (N_43945,N_42911,N_42127);
xor U43946 (N_43946,N_42220,N_42369);
nand U43947 (N_43947,N_42870,N_42071);
nand U43948 (N_43948,N_42331,N_42829);
or U43949 (N_43949,N_42345,N_42341);
or U43950 (N_43950,N_42529,N_42974);
and U43951 (N_43951,N_42210,N_42580);
and U43952 (N_43952,N_42715,N_42739);
nor U43953 (N_43953,N_42819,N_42191);
nand U43954 (N_43954,N_42204,N_42970);
xnor U43955 (N_43955,N_42625,N_42706);
nand U43956 (N_43956,N_42386,N_42264);
nor U43957 (N_43957,N_42757,N_42263);
or U43958 (N_43958,N_42963,N_42569);
or U43959 (N_43959,N_42099,N_42903);
nor U43960 (N_43960,N_42990,N_42425);
nor U43961 (N_43961,N_42376,N_42696);
nor U43962 (N_43962,N_42571,N_42126);
nand U43963 (N_43963,N_42322,N_42751);
or U43964 (N_43964,N_42993,N_42777);
xnor U43965 (N_43965,N_42658,N_42130);
and U43966 (N_43966,N_42782,N_42720);
nor U43967 (N_43967,N_42228,N_42159);
nand U43968 (N_43968,N_42696,N_42063);
xor U43969 (N_43969,N_42931,N_42565);
or U43970 (N_43970,N_42796,N_42563);
nor U43971 (N_43971,N_42153,N_42762);
and U43972 (N_43972,N_42713,N_42567);
xor U43973 (N_43973,N_42297,N_42469);
nand U43974 (N_43974,N_42558,N_42933);
nor U43975 (N_43975,N_42349,N_42250);
nand U43976 (N_43976,N_42149,N_42357);
nand U43977 (N_43977,N_42654,N_42155);
xnor U43978 (N_43978,N_42205,N_42262);
nand U43979 (N_43979,N_42412,N_42244);
xnor U43980 (N_43980,N_42405,N_42184);
nand U43981 (N_43981,N_42481,N_42311);
nor U43982 (N_43982,N_42139,N_42154);
or U43983 (N_43983,N_42537,N_42134);
and U43984 (N_43984,N_42443,N_42764);
nor U43985 (N_43985,N_42378,N_42167);
nor U43986 (N_43986,N_42012,N_42817);
nand U43987 (N_43987,N_42215,N_42574);
nor U43988 (N_43988,N_42465,N_42857);
and U43989 (N_43989,N_42903,N_42967);
or U43990 (N_43990,N_42912,N_42063);
nor U43991 (N_43991,N_42817,N_42225);
or U43992 (N_43992,N_42378,N_42466);
xnor U43993 (N_43993,N_42917,N_42422);
and U43994 (N_43994,N_42853,N_42976);
and U43995 (N_43995,N_42187,N_42523);
xor U43996 (N_43996,N_42740,N_42426);
xor U43997 (N_43997,N_42933,N_42310);
nand U43998 (N_43998,N_42077,N_42629);
or U43999 (N_43999,N_42953,N_42876);
nor U44000 (N_44000,N_43798,N_43180);
xor U44001 (N_44001,N_43689,N_43391);
or U44002 (N_44002,N_43264,N_43523);
or U44003 (N_44003,N_43290,N_43144);
and U44004 (N_44004,N_43673,N_43522);
xor U44005 (N_44005,N_43920,N_43303);
xnor U44006 (N_44006,N_43655,N_43637);
and U44007 (N_44007,N_43250,N_43823);
or U44008 (N_44008,N_43577,N_43829);
and U44009 (N_44009,N_43593,N_43441);
nor U44010 (N_44010,N_43267,N_43414);
and U44011 (N_44011,N_43618,N_43240);
nand U44012 (N_44012,N_43474,N_43625);
nand U44013 (N_44013,N_43682,N_43320);
nor U44014 (N_44014,N_43998,N_43179);
nor U44015 (N_44015,N_43480,N_43857);
nor U44016 (N_44016,N_43221,N_43862);
and U44017 (N_44017,N_43919,N_43098);
nand U44018 (N_44018,N_43923,N_43395);
and U44019 (N_44019,N_43960,N_43470);
nand U44020 (N_44020,N_43317,N_43888);
xor U44021 (N_44021,N_43776,N_43819);
nand U44022 (N_44022,N_43724,N_43357);
nor U44023 (N_44023,N_43204,N_43729);
and U44024 (N_44024,N_43217,N_43633);
and U44025 (N_44025,N_43503,N_43695);
nand U44026 (N_44026,N_43182,N_43068);
nor U44027 (N_44027,N_43559,N_43782);
nand U44028 (N_44028,N_43620,N_43773);
nor U44029 (N_44029,N_43984,N_43059);
and U44030 (N_44030,N_43659,N_43652);
and U44031 (N_44031,N_43093,N_43330);
and U44032 (N_44032,N_43425,N_43361);
nand U44033 (N_44033,N_43450,N_43260);
nor U44034 (N_44034,N_43460,N_43584);
or U44035 (N_44035,N_43585,N_43530);
and U44036 (N_44036,N_43266,N_43594);
nand U44037 (N_44037,N_43868,N_43427);
and U44038 (N_44038,N_43708,N_43821);
nand U44039 (N_44039,N_43948,N_43174);
and U44040 (N_44040,N_43797,N_43141);
or U44041 (N_44041,N_43884,N_43793);
nor U44042 (N_44042,N_43331,N_43915);
or U44043 (N_44043,N_43152,N_43022);
xnor U44044 (N_44044,N_43748,N_43513);
nand U44045 (N_44045,N_43945,N_43565);
nor U44046 (N_44046,N_43928,N_43683);
xnor U44047 (N_44047,N_43996,N_43483);
and U44048 (N_44048,N_43482,N_43670);
nand U44049 (N_44049,N_43115,N_43661);
nand U44050 (N_44050,N_43164,N_43281);
and U44051 (N_44051,N_43751,N_43101);
nand U44052 (N_44052,N_43185,N_43771);
xnor U44053 (N_44053,N_43785,N_43699);
or U44054 (N_44054,N_43551,N_43234);
xor U44055 (N_44055,N_43381,N_43018);
nand U44056 (N_44056,N_43490,N_43615);
xor U44057 (N_44057,N_43306,N_43844);
nand U44058 (N_44058,N_43858,N_43639);
nand U44059 (N_44059,N_43613,N_43826);
or U44060 (N_44060,N_43904,N_43006);
and U44061 (N_44061,N_43867,N_43027);
nand U44062 (N_44062,N_43273,N_43032);
and U44063 (N_44063,N_43953,N_43665);
nor U44064 (N_44064,N_43493,N_43009);
nor U44065 (N_44065,N_43869,N_43464);
nand U44066 (N_44066,N_43367,N_43050);
and U44067 (N_44067,N_43942,N_43225);
and U44068 (N_44068,N_43061,N_43031);
nor U44069 (N_44069,N_43548,N_43411);
nor U44070 (N_44070,N_43406,N_43456);
or U44071 (N_44071,N_43983,N_43758);
nor U44072 (N_44072,N_43759,N_43562);
and U44073 (N_44073,N_43828,N_43873);
xnor U44074 (N_44074,N_43910,N_43311);
nand U44075 (N_44075,N_43210,N_43728);
xnor U44076 (N_44076,N_43335,N_43448);
nor U44077 (N_44077,N_43872,N_43783);
nor U44078 (N_44078,N_43892,N_43726);
nand U44079 (N_44079,N_43796,N_43226);
nor U44080 (N_44080,N_43866,N_43712);
or U44081 (N_44081,N_43787,N_43012);
and U44082 (N_44082,N_43775,N_43128);
nand U44083 (N_44083,N_43140,N_43667);
nor U44084 (N_44084,N_43265,N_43014);
or U44085 (N_44085,N_43781,N_43791);
nand U44086 (N_44086,N_43081,N_43478);
or U44087 (N_44087,N_43889,N_43738);
or U44088 (N_44088,N_43696,N_43623);
or U44089 (N_44089,N_43853,N_43039);
nor U44090 (N_44090,N_43531,N_43519);
nand U44091 (N_44091,N_43930,N_43360);
nor U44092 (N_44092,N_43725,N_43774);
or U44093 (N_44093,N_43205,N_43851);
and U44094 (N_44094,N_43020,N_43354);
and U44095 (N_44095,N_43497,N_43291);
xnor U44096 (N_44096,N_43627,N_43046);
nand U44097 (N_44097,N_43878,N_43704);
xnor U44098 (N_44098,N_43003,N_43702);
and U44099 (N_44099,N_43143,N_43258);
and U44100 (N_44100,N_43526,N_43899);
xor U44101 (N_44101,N_43465,N_43447);
nor U44102 (N_44102,N_43309,N_43874);
and U44103 (N_44103,N_43811,N_43193);
xor U44104 (N_44104,N_43355,N_43803);
nor U44105 (N_44105,N_43084,N_43235);
or U44106 (N_44106,N_43590,N_43230);
and U44107 (N_44107,N_43149,N_43408);
and U44108 (N_44108,N_43897,N_43177);
nand U44109 (N_44109,N_43974,N_43108);
nor U44110 (N_44110,N_43206,N_43376);
nor U44111 (N_44111,N_43606,N_43938);
nor U44112 (N_44112,N_43799,N_43064);
and U44113 (N_44113,N_43589,N_43687);
xor U44114 (N_44114,N_43933,N_43778);
and U44115 (N_44115,N_43795,N_43552);
nand U44116 (N_44116,N_43214,N_43911);
or U44117 (N_44117,N_43901,N_43649);
or U44118 (N_44118,N_43534,N_43096);
xor U44119 (N_44119,N_43207,N_43476);
nand U44120 (N_44120,N_43788,N_43847);
nand U44121 (N_44121,N_43691,N_43527);
or U44122 (N_44122,N_43656,N_43895);
or U44123 (N_44123,N_43505,N_43834);
nor U44124 (N_44124,N_43040,N_43610);
or U44125 (N_44125,N_43780,N_43405);
and U44126 (N_44126,N_43626,N_43302);
and U44127 (N_44127,N_43727,N_43431);
and U44128 (N_44128,N_43877,N_43327);
xor U44129 (N_44129,N_43663,N_43069);
or U44130 (N_44130,N_43021,N_43364);
and U44131 (N_44131,N_43971,N_43338);
or U44132 (N_44132,N_43525,N_43843);
or U44133 (N_44133,N_43574,N_43734);
and U44134 (N_44134,N_43042,N_43351);
and U44135 (N_44135,N_43028,N_43047);
nand U44136 (N_44136,N_43218,N_43619);
and U44137 (N_44137,N_43103,N_43404);
nand U44138 (N_44138,N_43416,N_43166);
xnor U44139 (N_44139,N_43550,N_43010);
xor U44140 (N_44140,N_43669,N_43254);
nor U44141 (N_44141,N_43444,N_43510);
xnor U44142 (N_44142,N_43608,N_43628);
nand U44143 (N_44143,N_43840,N_43169);
xor U44144 (N_44144,N_43440,N_43388);
nand U44145 (N_44145,N_43817,N_43342);
and U44146 (N_44146,N_43555,N_43135);
xor U44147 (N_44147,N_43664,N_43162);
xor U44148 (N_44148,N_43657,N_43209);
and U44149 (N_44149,N_43413,N_43688);
or U44150 (N_44150,N_43442,N_43345);
nand U44151 (N_44151,N_43019,N_43779);
xnor U44152 (N_44152,N_43975,N_43638);
xor U44153 (N_44153,N_43126,N_43514);
or U44154 (N_44154,N_43242,N_43232);
or U44155 (N_44155,N_43592,N_43130);
or U44156 (N_44156,N_43245,N_43453);
xnor U44157 (N_44157,N_43644,N_43418);
and U44158 (N_44158,N_43350,N_43127);
xnor U44159 (N_44159,N_43706,N_43622);
and U44160 (N_44160,N_43479,N_43893);
xnor U44161 (N_44161,N_43386,N_43880);
nor U44162 (N_44162,N_43934,N_43715);
nor U44163 (N_44163,N_43473,N_43949);
nand U44164 (N_44164,N_43600,N_43832);
or U44165 (N_44165,N_43110,N_43927);
or U44166 (N_44166,N_43237,N_43253);
nor U44167 (N_44167,N_43255,N_43457);
or U44168 (N_44168,N_43885,N_43172);
nor U44169 (N_44169,N_43756,N_43407);
nand U44170 (N_44170,N_43336,N_43506);
nor U44171 (N_44171,N_43836,N_43362);
or U44172 (N_44172,N_43203,N_43583);
nand U44173 (N_44173,N_43859,N_43197);
nor U44174 (N_44174,N_43353,N_43684);
or U44175 (N_44175,N_43499,N_43641);
and U44176 (N_44176,N_43384,N_43681);
and U44177 (N_44177,N_43597,N_43060);
nor U44178 (N_44178,N_43539,N_43288);
and U44179 (N_44179,N_43990,N_43374);
nand U44180 (N_44180,N_43154,N_43153);
and U44181 (N_44181,N_43563,N_43117);
nand U44182 (N_44182,N_43243,N_43881);
nand U44183 (N_44183,N_43275,N_43257);
nand U44184 (N_44184,N_43321,N_43786);
xor U44185 (N_44185,N_43958,N_43168);
nor U44186 (N_44186,N_43557,N_43701);
nor U44187 (N_44187,N_43511,N_43766);
nand U44188 (N_44188,N_43090,N_43377);
xnor U44189 (N_44189,N_43845,N_43591);
nor U44190 (N_44190,N_43994,N_43297);
nand U44191 (N_44191,N_43274,N_43417);
nand U44192 (N_44192,N_43926,N_43807);
xor U44193 (N_44193,N_43790,N_43856);
and U44194 (N_44194,N_43211,N_43894);
or U44195 (N_44195,N_43538,N_43403);
nand U44196 (N_44196,N_43484,N_43215);
nor U44197 (N_44197,N_43650,N_43251);
nor U44198 (N_44198,N_43157,N_43635);
xnor U44199 (N_44199,N_43973,N_43269);
and U44200 (N_44200,N_43380,N_43515);
xor U44201 (N_44201,N_43762,N_43167);
or U44202 (N_44202,N_43842,N_43461);
xor U44203 (N_44203,N_43294,N_43272);
nor U44204 (N_44204,N_43744,N_43854);
and U44205 (N_44205,N_43993,N_43801);
or U44206 (N_44206,N_43908,N_43041);
xor U44207 (N_44207,N_43063,N_43770);
or U44208 (N_44208,N_43151,N_43914);
nor U44209 (N_44209,N_43287,N_43871);
or U44210 (N_44210,N_43703,N_43013);
xnor U44211 (N_44211,N_43825,N_43717);
nor U44212 (N_44212,N_43238,N_43936);
nor U44213 (N_44213,N_43337,N_43498);
xor U44214 (N_44214,N_43223,N_43423);
nor U44215 (N_44215,N_43079,N_43102);
and U44216 (N_44216,N_43595,N_43668);
nor U44217 (N_44217,N_43772,N_43433);
xor U44218 (N_44218,N_43653,N_43792);
xnor U44219 (N_44219,N_43816,N_43968);
and U44220 (N_44220,N_43752,N_43183);
and U44221 (N_44221,N_43753,N_43077);
nor U44222 (N_44222,N_43976,N_43198);
nand U44223 (N_44223,N_43768,N_43138);
xnor U44224 (N_44224,N_43369,N_43978);
or U44225 (N_44225,N_43654,N_43318);
nand U44226 (N_44226,N_43698,N_43158);
nand U44227 (N_44227,N_43742,N_43307);
and U44228 (N_44228,N_43091,N_43863);
xor U44229 (N_44229,N_43602,N_43429);
nor U44230 (N_44230,N_43679,N_43882);
nand U44231 (N_44231,N_43755,N_43319);
and U44232 (N_44232,N_43194,N_43105);
nand U44233 (N_44233,N_43849,N_43767);
or U44234 (N_44234,N_43937,N_43074);
nand U44235 (N_44235,N_43229,N_43095);
and U44236 (N_44236,N_43556,N_43282);
and U44237 (N_44237,N_43412,N_43283);
or U44238 (N_44238,N_43446,N_43463);
and U44239 (N_44239,N_43846,N_43390);
or U44240 (N_44240,N_43261,N_43067);
or U44241 (N_44241,N_43760,N_43458);
nand U44242 (N_44242,N_43344,N_43426);
nand U44243 (N_44243,N_43244,N_43542);
and U44244 (N_44244,N_43137,N_43436);
and U44245 (N_44245,N_43520,N_43705);
nor U44246 (N_44246,N_43045,N_43113);
and U44247 (N_44247,N_43213,N_43645);
xnor U44248 (N_44248,N_43420,N_43733);
and U44249 (N_44249,N_43969,N_43370);
nand U44250 (N_44250,N_43544,N_43747);
or U44251 (N_44251,N_43710,N_43268);
nor U44252 (N_44252,N_43488,N_43349);
or U44253 (N_44253,N_43509,N_43572);
xnor U44254 (N_44254,N_43718,N_43246);
or U44255 (N_44255,N_43106,N_43905);
xor U44256 (N_44256,N_43375,N_43954);
nand U44257 (N_44257,N_43611,N_43735);
or U44258 (N_44258,N_43459,N_43475);
nand U44259 (N_44259,N_43070,N_43328);
nor U44260 (N_44260,N_43629,N_43947);
or U44261 (N_44261,N_43578,N_43002);
xor U44262 (N_44262,N_43765,N_43648);
xor U44263 (N_44263,N_43502,N_43588);
xor U44264 (N_44264,N_43087,N_43686);
and U44265 (N_44265,N_43026,N_43902);
or U44266 (N_44266,N_43389,N_43746);
and U44267 (N_44267,N_43913,N_43017);
or U44268 (N_44268,N_43222,N_43850);
or U44269 (N_44269,N_43004,N_43721);
and U44270 (N_44270,N_43379,N_43270);
and U44271 (N_44271,N_43955,N_43449);
nand U44272 (N_44272,N_43672,N_43818);
and U44273 (N_44273,N_43887,N_43394);
xnor U44274 (N_44274,N_43604,N_43300);
or U44275 (N_44275,N_43991,N_43271);
and U44276 (N_44276,N_43815,N_43900);
xor U44277 (N_44277,N_43929,N_43324);
xor U44278 (N_44278,N_43575,N_43249);
and U44279 (N_44279,N_43359,N_43835);
and U44280 (N_44280,N_43005,N_43363);
nand U44281 (N_44281,N_43248,N_43398);
and U44282 (N_44282,N_43011,N_43500);
and U44283 (N_44283,N_43750,N_43912);
xor U44284 (N_44284,N_43956,N_43932);
xor U44285 (N_44285,N_43827,N_43219);
nand U44286 (N_44286,N_43924,N_43233);
nor U44287 (N_44287,N_43195,N_43481);
xnor U44288 (N_44288,N_43037,N_43739);
nand U44289 (N_44289,N_43580,N_43886);
or U44290 (N_44290,N_43546,N_43609);
and U44291 (N_44291,N_43421,N_43730);
or U44292 (N_44292,N_43935,N_43016);
nor U44293 (N_44293,N_43196,N_43316);
xor U44294 (N_44294,N_43333,N_43252);
or U44295 (N_44295,N_43651,N_43961);
nand U44296 (N_44296,N_43830,N_43891);
or U44297 (N_44297,N_43025,N_43468);
and U44298 (N_44298,N_43099,N_43477);
or U44299 (N_44299,N_43278,N_43997);
or U44300 (N_44300,N_43680,N_43368);
xor U44301 (N_44301,N_43434,N_43118);
or U44302 (N_44302,N_43295,N_43382);
and U44303 (N_44303,N_43631,N_43146);
xor U44304 (N_44304,N_43392,N_43241);
nor U44305 (N_44305,N_43305,N_43088);
nor U44306 (N_44306,N_43922,N_43100);
nand U44307 (N_44307,N_43008,N_43524);
and U44308 (N_44308,N_43860,N_43224);
and U44309 (N_44309,N_43634,N_43136);
nand U44310 (N_44310,N_43432,N_43000);
xor U44311 (N_44311,N_43171,N_43570);
and U44312 (N_44312,N_43455,N_43310);
nor U44313 (N_44313,N_43617,N_43612);
and U44314 (N_44314,N_43685,N_43055);
xor U44315 (N_44315,N_43848,N_43078);
nand U44316 (N_44316,N_43341,N_43616);
xnor U44317 (N_44317,N_43133,N_43097);
nand U44318 (N_44318,N_43443,N_43076);
or U44319 (N_44319,N_43831,N_43424);
nand U44320 (N_44320,N_43707,N_43841);
and U44321 (N_44321,N_43714,N_43540);
and U44322 (N_44322,N_43605,N_43709);
or U44323 (N_44323,N_43279,N_43116);
xnor U44324 (N_44324,N_43247,N_43800);
nand U44325 (N_44325,N_43190,N_43112);
and U44326 (N_44326,N_43082,N_43131);
and U44327 (N_44327,N_43228,N_43023);
xor U44328 (N_44328,N_43621,N_43549);
and U44329 (N_44329,N_43794,N_43532);
nand U44330 (N_44330,N_43950,N_43284);
xor U44331 (N_44331,N_43992,N_43155);
or U44332 (N_44332,N_43987,N_43208);
and U44333 (N_44333,N_43940,N_43967);
nor U44334 (N_44334,N_43723,N_43693);
nand U44335 (N_44335,N_43601,N_43537);
nand U44336 (N_44336,N_43038,N_43372);
xor U44337 (N_44337,N_43301,N_43065);
xnor U44338 (N_44338,N_43861,N_43554);
nand U44339 (N_44339,N_43262,N_43982);
or U44340 (N_44340,N_43371,N_43286);
xnor U44341 (N_44341,N_43276,N_43467);
nand U44342 (N_44342,N_43690,N_43256);
nand U44343 (N_44343,N_43259,N_43486);
nand U44344 (N_44344,N_43263,N_43086);
nand U44345 (N_44345,N_43543,N_43517);
or U44346 (N_44346,N_43957,N_43986);
and U44347 (N_44347,N_43397,N_43358);
and U44348 (N_44348,N_43339,N_43666);
or U44349 (N_44349,N_43757,N_43373);
and U44350 (N_44350,N_43365,N_43719);
nor U44351 (N_44351,N_43989,N_43876);
or U44352 (N_44352,N_43139,N_43917);
xor U44353 (N_44353,N_43521,N_43736);
and U44354 (N_44354,N_43569,N_43896);
nor U44355 (N_44355,N_43573,N_43784);
nand U44356 (N_44356,N_43007,N_43178);
or U44357 (N_44357,N_43504,N_43495);
and U44358 (N_44358,N_43553,N_43356);
nand U44359 (N_44359,N_43737,N_43864);
nand U44360 (N_44360,N_43428,N_43805);
nor U44361 (N_44361,N_43491,N_43348);
xor U44362 (N_44362,N_43277,N_43820);
and U44363 (N_44363,N_43722,N_43329);
nand U44364 (N_44364,N_43567,N_43471);
nor U44365 (N_44365,N_43492,N_43058);
and U44366 (N_44366,N_43676,N_43430);
nand U44367 (N_44367,N_43496,N_43184);
nand U44368 (N_44368,N_43163,N_43299);
nor U44369 (N_44369,N_43073,N_43325);
xnor U44370 (N_44370,N_43134,N_43870);
xnor U44371 (N_44371,N_43199,N_43660);
and U44372 (N_44372,N_43312,N_43813);
xnor U44373 (N_44373,N_43995,N_43966);
nand U44374 (N_44374,N_43528,N_43814);
xnor U44375 (N_44375,N_43646,N_43323);
nor U44376 (N_44376,N_43024,N_43985);
xor U44377 (N_44377,N_43720,N_43123);
or U44378 (N_44378,N_43466,N_43422);
xnor U44379 (N_44379,N_43603,N_43571);
nand U44380 (N_44380,N_43094,N_43700);
xnor U44381 (N_44381,N_43401,N_43396);
nor U44382 (N_44382,N_43125,N_43314);
and U44383 (N_44383,N_43564,N_43160);
nand U44384 (N_44384,N_43536,N_43907);
and U44385 (N_44385,N_43366,N_43107);
nor U44386 (N_44386,N_43962,N_43675);
and U44387 (N_44387,N_43545,N_43231);
xnor U44388 (N_44388,N_43822,N_43075);
nand U44389 (N_44389,N_43202,N_43315);
xnor U44390 (N_44390,N_43340,N_43121);
xnor U44391 (N_44391,N_43036,N_43711);
and U44392 (N_44392,N_43630,N_43713);
nand U44393 (N_44393,N_43963,N_43030);
or U44394 (N_44394,N_43547,N_43201);
nand U44395 (N_44395,N_43918,N_43582);
xor U44396 (N_44396,N_43965,N_43692);
nor U44397 (N_44397,N_43147,N_43501);
nand U44398 (N_44398,N_43313,N_43981);
nor U44399 (N_44399,N_43632,N_43001);
or U44400 (N_44400,N_43581,N_43409);
or U44401 (N_44401,N_43494,N_43150);
xnor U44402 (N_44402,N_43883,N_43764);
nand U44403 (N_44403,N_43561,N_43212);
xnor U44404 (N_44404,N_43142,N_43763);
nand U44405 (N_44405,N_43034,N_43640);
or U44406 (N_44406,N_43109,N_43393);
xnor U44407 (N_44407,N_43454,N_43120);
or U44408 (N_44408,N_43732,N_43906);
or U44409 (N_44409,N_43298,N_43879);
nand U44410 (N_44410,N_43740,N_43192);
nand U44411 (N_44411,N_43239,N_43541);
xnor U44412 (N_44412,N_43035,N_43293);
xnor U44413 (N_44413,N_43944,N_43508);
xnor U44414 (N_44414,N_43308,N_43469);
and U44415 (N_44415,N_43809,N_43529);
or U44416 (N_44416,N_43326,N_43216);
or U44417 (N_44417,N_43921,N_43598);
nor U44418 (N_44418,N_43343,N_43806);
or U44419 (N_44419,N_43435,N_43033);
nand U44420 (N_44420,N_43159,N_43062);
or U44421 (N_44421,N_43200,N_43769);
xor U44422 (N_44422,N_43674,N_43614);
nor U44423 (N_44423,N_43999,N_43236);
nor U44424 (N_44424,N_43485,N_43472);
or U44425 (N_44425,N_43964,N_43187);
and U44426 (N_44426,N_43643,N_43385);
xor U44427 (N_44427,N_43642,N_43439);
nor U44428 (N_44428,N_43898,N_43754);
nor U44429 (N_44429,N_43579,N_43399);
nor U44430 (N_44430,N_43015,N_43462);
nand U44431 (N_44431,N_43452,N_43925);
or U44432 (N_44432,N_43916,N_43951);
xor U44433 (N_44433,N_43083,N_43931);
xnor U44434 (N_44434,N_43292,N_43749);
nand U44435 (N_44435,N_43839,N_43952);
nand U44436 (N_44436,N_43186,N_43285);
xnor U44437 (N_44437,N_43568,N_43148);
xor U44438 (N_44438,N_43970,N_43587);
or U44439 (N_44439,N_43533,N_43662);
and U44440 (N_44440,N_43512,N_43437);
nor U44441 (N_44441,N_43636,N_43560);
nor U44442 (N_44442,N_43156,N_43596);
and U44443 (N_44443,N_43378,N_43658);
xor U44444 (N_44444,N_43535,N_43352);
and U44445 (N_44445,N_43808,N_43451);
and U44446 (N_44446,N_43056,N_43145);
xor U44447 (N_44447,N_43647,N_43049);
or U44448 (N_44448,N_43789,N_43052);
nand U44449 (N_44449,N_43119,N_43487);
xnor U44450 (N_44450,N_43387,N_43189);
and U44451 (N_44451,N_43875,N_43607);
nor U44452 (N_44452,N_43122,N_43802);
xnor U44453 (N_44453,N_43289,N_43838);
or U44454 (N_44454,N_43777,N_43518);
and U44455 (N_44455,N_43053,N_43132);
and U44456 (N_44456,N_43048,N_43029);
and U44457 (N_44457,N_43810,N_43445);
nor U44458 (N_44458,N_43220,N_43402);
and U44459 (N_44459,N_43066,N_43181);
nor U44460 (N_44460,N_43694,N_43833);
nand U44461 (N_44461,N_43939,N_43812);
and U44462 (N_44462,N_43716,N_43104);
or U44463 (N_44463,N_43347,N_43415);
nand U44464 (N_44464,N_43165,N_43980);
nand U44465 (N_44465,N_43979,N_43188);
and U44466 (N_44466,N_43671,N_43852);
nand U44467 (N_44467,N_43697,N_43054);
xor U44468 (N_44468,N_43678,N_43129);
or U44469 (N_44469,N_43988,N_43855);
nor U44470 (N_44470,N_43161,N_43890);
or U44471 (N_44471,N_43191,N_43332);
nor U44472 (N_44472,N_43280,N_43089);
xor U44473 (N_44473,N_43072,N_43400);
nand U44474 (N_44474,N_43304,N_43837);
nor U44475 (N_44475,N_43043,N_43346);
nor U44476 (N_44476,N_43176,N_43092);
nand U44477 (N_44477,N_43057,N_43946);
or U44478 (N_44478,N_43909,N_43175);
nand U44479 (N_44479,N_43438,N_43383);
nor U44480 (N_44480,N_43080,N_43865);
nor U44481 (N_44481,N_43824,N_43576);
and U44482 (N_44482,N_43745,N_43124);
nor U44483 (N_44483,N_43941,N_43111);
and U44484 (N_44484,N_43761,N_43558);
or U44485 (N_44485,N_43071,N_43903);
and U44486 (N_44486,N_43419,N_43051);
and U44487 (N_44487,N_43959,N_43977);
nand U44488 (N_44488,N_43943,N_43516);
nand U44489 (N_44489,N_43489,N_43804);
and U44490 (N_44490,N_43227,N_43599);
xor U44491 (N_44491,N_43731,N_43173);
nor U44492 (N_44492,N_43334,N_43507);
xor U44493 (N_44493,N_43085,N_43170);
xor U44494 (N_44494,N_43677,N_43741);
xor U44495 (N_44495,N_43044,N_43114);
nand U44496 (N_44496,N_43566,N_43743);
nor U44497 (N_44497,N_43624,N_43296);
xnor U44498 (N_44498,N_43410,N_43322);
nor U44499 (N_44499,N_43972,N_43586);
nand U44500 (N_44500,N_43744,N_43961);
xnor U44501 (N_44501,N_43343,N_43163);
xor U44502 (N_44502,N_43574,N_43713);
xnor U44503 (N_44503,N_43639,N_43314);
or U44504 (N_44504,N_43483,N_43395);
nand U44505 (N_44505,N_43339,N_43786);
or U44506 (N_44506,N_43998,N_43779);
xnor U44507 (N_44507,N_43086,N_43198);
xor U44508 (N_44508,N_43214,N_43800);
nor U44509 (N_44509,N_43171,N_43734);
or U44510 (N_44510,N_43299,N_43491);
nand U44511 (N_44511,N_43353,N_43018);
and U44512 (N_44512,N_43354,N_43460);
or U44513 (N_44513,N_43782,N_43141);
and U44514 (N_44514,N_43902,N_43204);
and U44515 (N_44515,N_43920,N_43133);
and U44516 (N_44516,N_43026,N_43826);
nand U44517 (N_44517,N_43624,N_43573);
or U44518 (N_44518,N_43607,N_43748);
or U44519 (N_44519,N_43073,N_43349);
or U44520 (N_44520,N_43227,N_43396);
and U44521 (N_44521,N_43996,N_43723);
or U44522 (N_44522,N_43904,N_43964);
nand U44523 (N_44523,N_43889,N_43090);
nor U44524 (N_44524,N_43076,N_43233);
or U44525 (N_44525,N_43138,N_43301);
nor U44526 (N_44526,N_43425,N_43325);
nor U44527 (N_44527,N_43747,N_43858);
nand U44528 (N_44528,N_43423,N_43893);
nor U44529 (N_44529,N_43862,N_43153);
or U44530 (N_44530,N_43725,N_43107);
or U44531 (N_44531,N_43240,N_43472);
and U44532 (N_44532,N_43533,N_43104);
or U44533 (N_44533,N_43608,N_43190);
and U44534 (N_44534,N_43907,N_43963);
nand U44535 (N_44535,N_43062,N_43507);
nor U44536 (N_44536,N_43804,N_43697);
and U44537 (N_44537,N_43523,N_43069);
nor U44538 (N_44538,N_43976,N_43431);
and U44539 (N_44539,N_43533,N_43780);
xnor U44540 (N_44540,N_43866,N_43614);
nor U44541 (N_44541,N_43228,N_43819);
and U44542 (N_44542,N_43849,N_43397);
and U44543 (N_44543,N_43110,N_43975);
nor U44544 (N_44544,N_43605,N_43985);
nand U44545 (N_44545,N_43627,N_43545);
or U44546 (N_44546,N_43061,N_43243);
and U44547 (N_44547,N_43577,N_43540);
nor U44548 (N_44548,N_43315,N_43761);
and U44549 (N_44549,N_43532,N_43091);
nor U44550 (N_44550,N_43542,N_43156);
nor U44551 (N_44551,N_43124,N_43030);
xnor U44552 (N_44552,N_43952,N_43245);
nand U44553 (N_44553,N_43855,N_43937);
or U44554 (N_44554,N_43014,N_43850);
and U44555 (N_44555,N_43418,N_43802);
xor U44556 (N_44556,N_43677,N_43642);
nand U44557 (N_44557,N_43705,N_43188);
nor U44558 (N_44558,N_43744,N_43571);
nand U44559 (N_44559,N_43308,N_43950);
xor U44560 (N_44560,N_43923,N_43009);
and U44561 (N_44561,N_43896,N_43292);
xor U44562 (N_44562,N_43411,N_43119);
nand U44563 (N_44563,N_43243,N_43322);
and U44564 (N_44564,N_43557,N_43743);
xor U44565 (N_44565,N_43033,N_43097);
or U44566 (N_44566,N_43828,N_43113);
and U44567 (N_44567,N_43400,N_43807);
nand U44568 (N_44568,N_43315,N_43865);
xor U44569 (N_44569,N_43974,N_43951);
and U44570 (N_44570,N_43680,N_43700);
or U44571 (N_44571,N_43173,N_43161);
nor U44572 (N_44572,N_43010,N_43156);
nand U44573 (N_44573,N_43274,N_43612);
and U44574 (N_44574,N_43879,N_43791);
nand U44575 (N_44575,N_43834,N_43165);
xor U44576 (N_44576,N_43516,N_43926);
nand U44577 (N_44577,N_43213,N_43139);
and U44578 (N_44578,N_43826,N_43473);
or U44579 (N_44579,N_43510,N_43132);
xor U44580 (N_44580,N_43339,N_43121);
nor U44581 (N_44581,N_43903,N_43252);
nand U44582 (N_44582,N_43340,N_43657);
nand U44583 (N_44583,N_43299,N_43882);
xnor U44584 (N_44584,N_43535,N_43515);
xor U44585 (N_44585,N_43817,N_43469);
xor U44586 (N_44586,N_43421,N_43133);
nor U44587 (N_44587,N_43122,N_43928);
or U44588 (N_44588,N_43381,N_43247);
and U44589 (N_44589,N_43105,N_43223);
xnor U44590 (N_44590,N_43123,N_43638);
nand U44591 (N_44591,N_43331,N_43261);
nor U44592 (N_44592,N_43038,N_43020);
nand U44593 (N_44593,N_43039,N_43467);
xnor U44594 (N_44594,N_43368,N_43117);
nor U44595 (N_44595,N_43250,N_43448);
nor U44596 (N_44596,N_43042,N_43066);
xor U44597 (N_44597,N_43733,N_43957);
and U44598 (N_44598,N_43434,N_43183);
nor U44599 (N_44599,N_43724,N_43602);
or U44600 (N_44600,N_43522,N_43775);
or U44601 (N_44601,N_43128,N_43542);
and U44602 (N_44602,N_43062,N_43746);
xnor U44603 (N_44603,N_43561,N_43096);
or U44604 (N_44604,N_43464,N_43654);
nor U44605 (N_44605,N_43688,N_43211);
xor U44606 (N_44606,N_43989,N_43402);
or U44607 (N_44607,N_43802,N_43850);
or U44608 (N_44608,N_43928,N_43116);
nand U44609 (N_44609,N_43507,N_43428);
nor U44610 (N_44610,N_43957,N_43370);
nand U44611 (N_44611,N_43767,N_43408);
nor U44612 (N_44612,N_43304,N_43282);
nor U44613 (N_44613,N_43139,N_43186);
nor U44614 (N_44614,N_43752,N_43282);
xor U44615 (N_44615,N_43123,N_43070);
nor U44616 (N_44616,N_43986,N_43987);
and U44617 (N_44617,N_43336,N_43773);
or U44618 (N_44618,N_43903,N_43189);
or U44619 (N_44619,N_43976,N_43900);
or U44620 (N_44620,N_43372,N_43110);
nor U44621 (N_44621,N_43763,N_43658);
nand U44622 (N_44622,N_43636,N_43476);
or U44623 (N_44623,N_43676,N_43413);
or U44624 (N_44624,N_43365,N_43592);
and U44625 (N_44625,N_43571,N_43535);
or U44626 (N_44626,N_43460,N_43537);
xnor U44627 (N_44627,N_43413,N_43523);
or U44628 (N_44628,N_43120,N_43759);
nand U44629 (N_44629,N_43838,N_43506);
or U44630 (N_44630,N_43270,N_43951);
or U44631 (N_44631,N_43713,N_43993);
nand U44632 (N_44632,N_43669,N_43570);
nand U44633 (N_44633,N_43208,N_43436);
or U44634 (N_44634,N_43437,N_43214);
or U44635 (N_44635,N_43995,N_43313);
nor U44636 (N_44636,N_43171,N_43097);
or U44637 (N_44637,N_43110,N_43654);
nor U44638 (N_44638,N_43089,N_43180);
and U44639 (N_44639,N_43554,N_43487);
xnor U44640 (N_44640,N_43767,N_43111);
and U44641 (N_44641,N_43096,N_43281);
or U44642 (N_44642,N_43499,N_43513);
and U44643 (N_44643,N_43297,N_43222);
nor U44644 (N_44644,N_43392,N_43568);
or U44645 (N_44645,N_43510,N_43823);
and U44646 (N_44646,N_43853,N_43693);
and U44647 (N_44647,N_43575,N_43354);
and U44648 (N_44648,N_43690,N_43722);
nand U44649 (N_44649,N_43455,N_43255);
nor U44650 (N_44650,N_43859,N_43833);
xor U44651 (N_44651,N_43870,N_43167);
or U44652 (N_44652,N_43039,N_43925);
xnor U44653 (N_44653,N_43062,N_43772);
nor U44654 (N_44654,N_43920,N_43342);
and U44655 (N_44655,N_43198,N_43140);
or U44656 (N_44656,N_43774,N_43646);
xor U44657 (N_44657,N_43468,N_43783);
xnor U44658 (N_44658,N_43662,N_43077);
xor U44659 (N_44659,N_43443,N_43452);
xor U44660 (N_44660,N_43577,N_43757);
or U44661 (N_44661,N_43420,N_43655);
or U44662 (N_44662,N_43599,N_43916);
and U44663 (N_44663,N_43125,N_43419);
nor U44664 (N_44664,N_43989,N_43913);
nand U44665 (N_44665,N_43192,N_43985);
nand U44666 (N_44666,N_43131,N_43445);
nand U44667 (N_44667,N_43242,N_43866);
nor U44668 (N_44668,N_43513,N_43573);
nand U44669 (N_44669,N_43516,N_43504);
or U44670 (N_44670,N_43421,N_43092);
xor U44671 (N_44671,N_43985,N_43987);
or U44672 (N_44672,N_43696,N_43085);
and U44673 (N_44673,N_43235,N_43588);
nand U44674 (N_44674,N_43560,N_43254);
nor U44675 (N_44675,N_43618,N_43610);
xor U44676 (N_44676,N_43033,N_43695);
nand U44677 (N_44677,N_43023,N_43846);
nor U44678 (N_44678,N_43251,N_43883);
xor U44679 (N_44679,N_43652,N_43079);
nand U44680 (N_44680,N_43734,N_43279);
or U44681 (N_44681,N_43225,N_43984);
nor U44682 (N_44682,N_43831,N_43390);
nor U44683 (N_44683,N_43567,N_43599);
and U44684 (N_44684,N_43652,N_43983);
and U44685 (N_44685,N_43103,N_43166);
or U44686 (N_44686,N_43584,N_43053);
or U44687 (N_44687,N_43012,N_43629);
nand U44688 (N_44688,N_43024,N_43797);
xor U44689 (N_44689,N_43884,N_43012);
or U44690 (N_44690,N_43169,N_43617);
and U44691 (N_44691,N_43201,N_43838);
xor U44692 (N_44692,N_43138,N_43150);
or U44693 (N_44693,N_43741,N_43728);
xor U44694 (N_44694,N_43312,N_43339);
xor U44695 (N_44695,N_43706,N_43256);
nand U44696 (N_44696,N_43690,N_43143);
and U44697 (N_44697,N_43428,N_43911);
nand U44698 (N_44698,N_43544,N_43620);
and U44699 (N_44699,N_43872,N_43934);
or U44700 (N_44700,N_43689,N_43787);
xnor U44701 (N_44701,N_43050,N_43292);
and U44702 (N_44702,N_43341,N_43461);
or U44703 (N_44703,N_43324,N_43486);
and U44704 (N_44704,N_43214,N_43072);
and U44705 (N_44705,N_43636,N_43894);
or U44706 (N_44706,N_43850,N_43268);
or U44707 (N_44707,N_43552,N_43368);
nand U44708 (N_44708,N_43033,N_43305);
nand U44709 (N_44709,N_43272,N_43621);
and U44710 (N_44710,N_43936,N_43472);
and U44711 (N_44711,N_43929,N_43170);
nor U44712 (N_44712,N_43644,N_43951);
xnor U44713 (N_44713,N_43573,N_43230);
xnor U44714 (N_44714,N_43803,N_43150);
xnor U44715 (N_44715,N_43751,N_43140);
nand U44716 (N_44716,N_43427,N_43885);
and U44717 (N_44717,N_43558,N_43967);
xnor U44718 (N_44718,N_43501,N_43260);
nand U44719 (N_44719,N_43801,N_43504);
nand U44720 (N_44720,N_43408,N_43394);
xnor U44721 (N_44721,N_43492,N_43645);
xor U44722 (N_44722,N_43476,N_43005);
xor U44723 (N_44723,N_43864,N_43223);
xor U44724 (N_44724,N_43394,N_43087);
or U44725 (N_44725,N_43577,N_43926);
nor U44726 (N_44726,N_43192,N_43313);
or U44727 (N_44727,N_43653,N_43363);
and U44728 (N_44728,N_43646,N_43096);
nor U44729 (N_44729,N_43906,N_43636);
nor U44730 (N_44730,N_43437,N_43952);
nand U44731 (N_44731,N_43133,N_43364);
nor U44732 (N_44732,N_43197,N_43508);
nand U44733 (N_44733,N_43150,N_43379);
or U44734 (N_44734,N_43628,N_43556);
nor U44735 (N_44735,N_43779,N_43657);
nor U44736 (N_44736,N_43085,N_43479);
xor U44737 (N_44737,N_43338,N_43019);
nor U44738 (N_44738,N_43717,N_43018);
or U44739 (N_44739,N_43312,N_43057);
or U44740 (N_44740,N_43042,N_43572);
xor U44741 (N_44741,N_43974,N_43357);
and U44742 (N_44742,N_43915,N_43276);
and U44743 (N_44743,N_43847,N_43513);
and U44744 (N_44744,N_43284,N_43379);
nand U44745 (N_44745,N_43740,N_43978);
nor U44746 (N_44746,N_43449,N_43278);
or U44747 (N_44747,N_43727,N_43740);
xor U44748 (N_44748,N_43000,N_43320);
and U44749 (N_44749,N_43837,N_43144);
xor U44750 (N_44750,N_43866,N_43941);
nor U44751 (N_44751,N_43998,N_43582);
nor U44752 (N_44752,N_43052,N_43004);
and U44753 (N_44753,N_43140,N_43396);
and U44754 (N_44754,N_43613,N_43947);
and U44755 (N_44755,N_43540,N_43394);
or U44756 (N_44756,N_43004,N_43787);
and U44757 (N_44757,N_43089,N_43034);
and U44758 (N_44758,N_43300,N_43454);
and U44759 (N_44759,N_43079,N_43760);
nor U44760 (N_44760,N_43751,N_43513);
and U44761 (N_44761,N_43543,N_43981);
or U44762 (N_44762,N_43314,N_43996);
and U44763 (N_44763,N_43464,N_43313);
nor U44764 (N_44764,N_43168,N_43403);
nand U44765 (N_44765,N_43122,N_43257);
or U44766 (N_44766,N_43460,N_43156);
and U44767 (N_44767,N_43121,N_43243);
and U44768 (N_44768,N_43349,N_43903);
or U44769 (N_44769,N_43204,N_43338);
and U44770 (N_44770,N_43147,N_43299);
nor U44771 (N_44771,N_43205,N_43709);
and U44772 (N_44772,N_43133,N_43008);
nand U44773 (N_44773,N_43138,N_43139);
and U44774 (N_44774,N_43500,N_43910);
nand U44775 (N_44775,N_43537,N_43626);
and U44776 (N_44776,N_43992,N_43909);
nor U44777 (N_44777,N_43947,N_43496);
xnor U44778 (N_44778,N_43266,N_43590);
nor U44779 (N_44779,N_43049,N_43175);
and U44780 (N_44780,N_43295,N_43461);
xor U44781 (N_44781,N_43073,N_43367);
and U44782 (N_44782,N_43235,N_43370);
nand U44783 (N_44783,N_43454,N_43597);
and U44784 (N_44784,N_43159,N_43971);
xor U44785 (N_44785,N_43077,N_43632);
nand U44786 (N_44786,N_43565,N_43140);
and U44787 (N_44787,N_43600,N_43744);
xor U44788 (N_44788,N_43898,N_43891);
and U44789 (N_44789,N_43652,N_43590);
xnor U44790 (N_44790,N_43298,N_43130);
nand U44791 (N_44791,N_43884,N_43680);
and U44792 (N_44792,N_43399,N_43227);
nand U44793 (N_44793,N_43948,N_43226);
or U44794 (N_44794,N_43013,N_43579);
nor U44795 (N_44795,N_43540,N_43411);
or U44796 (N_44796,N_43164,N_43174);
nand U44797 (N_44797,N_43131,N_43971);
xnor U44798 (N_44798,N_43095,N_43734);
and U44799 (N_44799,N_43310,N_43836);
nor U44800 (N_44800,N_43448,N_43098);
xor U44801 (N_44801,N_43900,N_43896);
xor U44802 (N_44802,N_43216,N_43626);
nand U44803 (N_44803,N_43934,N_43633);
and U44804 (N_44804,N_43434,N_43713);
xnor U44805 (N_44805,N_43277,N_43797);
or U44806 (N_44806,N_43450,N_43601);
or U44807 (N_44807,N_43311,N_43485);
and U44808 (N_44808,N_43053,N_43388);
xnor U44809 (N_44809,N_43913,N_43435);
or U44810 (N_44810,N_43180,N_43814);
nand U44811 (N_44811,N_43249,N_43083);
nand U44812 (N_44812,N_43776,N_43089);
xor U44813 (N_44813,N_43812,N_43112);
xor U44814 (N_44814,N_43609,N_43051);
xor U44815 (N_44815,N_43288,N_43371);
and U44816 (N_44816,N_43595,N_43149);
or U44817 (N_44817,N_43395,N_43231);
or U44818 (N_44818,N_43342,N_43437);
nand U44819 (N_44819,N_43108,N_43977);
nor U44820 (N_44820,N_43873,N_43256);
xor U44821 (N_44821,N_43068,N_43687);
nor U44822 (N_44822,N_43325,N_43708);
xor U44823 (N_44823,N_43035,N_43992);
or U44824 (N_44824,N_43149,N_43358);
nand U44825 (N_44825,N_43616,N_43469);
and U44826 (N_44826,N_43412,N_43755);
nand U44827 (N_44827,N_43673,N_43191);
nand U44828 (N_44828,N_43590,N_43737);
or U44829 (N_44829,N_43883,N_43364);
or U44830 (N_44830,N_43341,N_43635);
nand U44831 (N_44831,N_43819,N_43195);
nand U44832 (N_44832,N_43869,N_43765);
or U44833 (N_44833,N_43666,N_43580);
nor U44834 (N_44834,N_43919,N_43059);
xor U44835 (N_44835,N_43092,N_43667);
or U44836 (N_44836,N_43646,N_43425);
xor U44837 (N_44837,N_43164,N_43724);
and U44838 (N_44838,N_43606,N_43747);
nand U44839 (N_44839,N_43083,N_43006);
nor U44840 (N_44840,N_43856,N_43824);
xor U44841 (N_44841,N_43865,N_43996);
and U44842 (N_44842,N_43742,N_43387);
xor U44843 (N_44843,N_43596,N_43744);
xor U44844 (N_44844,N_43926,N_43056);
nand U44845 (N_44845,N_43548,N_43939);
and U44846 (N_44846,N_43198,N_43375);
xor U44847 (N_44847,N_43698,N_43340);
or U44848 (N_44848,N_43446,N_43997);
nand U44849 (N_44849,N_43389,N_43598);
or U44850 (N_44850,N_43496,N_43895);
nor U44851 (N_44851,N_43044,N_43098);
or U44852 (N_44852,N_43533,N_43096);
nand U44853 (N_44853,N_43658,N_43366);
nand U44854 (N_44854,N_43601,N_43206);
xnor U44855 (N_44855,N_43536,N_43308);
nand U44856 (N_44856,N_43544,N_43781);
nor U44857 (N_44857,N_43810,N_43051);
xnor U44858 (N_44858,N_43611,N_43948);
nor U44859 (N_44859,N_43351,N_43270);
xor U44860 (N_44860,N_43310,N_43038);
and U44861 (N_44861,N_43378,N_43602);
nor U44862 (N_44862,N_43421,N_43627);
nor U44863 (N_44863,N_43347,N_43298);
nand U44864 (N_44864,N_43982,N_43574);
nand U44865 (N_44865,N_43088,N_43371);
xnor U44866 (N_44866,N_43698,N_43436);
or U44867 (N_44867,N_43639,N_43798);
or U44868 (N_44868,N_43391,N_43439);
or U44869 (N_44869,N_43070,N_43026);
and U44870 (N_44870,N_43556,N_43320);
nor U44871 (N_44871,N_43899,N_43110);
xor U44872 (N_44872,N_43745,N_43024);
nand U44873 (N_44873,N_43586,N_43303);
xnor U44874 (N_44874,N_43586,N_43676);
nand U44875 (N_44875,N_43811,N_43183);
nand U44876 (N_44876,N_43522,N_43331);
xor U44877 (N_44877,N_43523,N_43780);
xor U44878 (N_44878,N_43916,N_43489);
nor U44879 (N_44879,N_43270,N_43979);
and U44880 (N_44880,N_43052,N_43374);
and U44881 (N_44881,N_43320,N_43976);
and U44882 (N_44882,N_43243,N_43312);
nor U44883 (N_44883,N_43239,N_43802);
nor U44884 (N_44884,N_43864,N_43398);
and U44885 (N_44885,N_43064,N_43228);
and U44886 (N_44886,N_43746,N_43769);
nand U44887 (N_44887,N_43187,N_43700);
xor U44888 (N_44888,N_43444,N_43469);
nand U44889 (N_44889,N_43256,N_43440);
xor U44890 (N_44890,N_43655,N_43932);
nand U44891 (N_44891,N_43717,N_43481);
or U44892 (N_44892,N_43488,N_43160);
nor U44893 (N_44893,N_43014,N_43784);
or U44894 (N_44894,N_43172,N_43820);
and U44895 (N_44895,N_43229,N_43380);
nand U44896 (N_44896,N_43217,N_43452);
nor U44897 (N_44897,N_43934,N_43564);
nand U44898 (N_44898,N_43260,N_43792);
nor U44899 (N_44899,N_43667,N_43115);
xnor U44900 (N_44900,N_43162,N_43510);
or U44901 (N_44901,N_43178,N_43191);
nand U44902 (N_44902,N_43266,N_43953);
or U44903 (N_44903,N_43508,N_43936);
xnor U44904 (N_44904,N_43652,N_43296);
nor U44905 (N_44905,N_43272,N_43835);
nand U44906 (N_44906,N_43515,N_43666);
nor U44907 (N_44907,N_43245,N_43630);
and U44908 (N_44908,N_43601,N_43984);
or U44909 (N_44909,N_43812,N_43833);
nand U44910 (N_44910,N_43136,N_43122);
and U44911 (N_44911,N_43661,N_43838);
and U44912 (N_44912,N_43669,N_43766);
nand U44913 (N_44913,N_43207,N_43340);
nand U44914 (N_44914,N_43617,N_43191);
or U44915 (N_44915,N_43438,N_43596);
nor U44916 (N_44916,N_43559,N_43154);
nand U44917 (N_44917,N_43377,N_43001);
nand U44918 (N_44918,N_43835,N_43083);
nor U44919 (N_44919,N_43227,N_43081);
nor U44920 (N_44920,N_43806,N_43349);
or U44921 (N_44921,N_43378,N_43111);
nor U44922 (N_44922,N_43307,N_43187);
nor U44923 (N_44923,N_43922,N_43420);
or U44924 (N_44924,N_43077,N_43989);
xnor U44925 (N_44925,N_43130,N_43855);
or U44926 (N_44926,N_43757,N_43975);
xnor U44927 (N_44927,N_43508,N_43877);
nand U44928 (N_44928,N_43696,N_43821);
xor U44929 (N_44929,N_43856,N_43322);
or U44930 (N_44930,N_43501,N_43757);
or U44931 (N_44931,N_43960,N_43842);
nor U44932 (N_44932,N_43783,N_43241);
xnor U44933 (N_44933,N_43159,N_43781);
and U44934 (N_44934,N_43285,N_43274);
xnor U44935 (N_44935,N_43544,N_43602);
and U44936 (N_44936,N_43360,N_43512);
nor U44937 (N_44937,N_43555,N_43515);
xnor U44938 (N_44938,N_43111,N_43895);
and U44939 (N_44939,N_43840,N_43149);
and U44940 (N_44940,N_43080,N_43317);
nor U44941 (N_44941,N_43249,N_43796);
xor U44942 (N_44942,N_43759,N_43518);
and U44943 (N_44943,N_43711,N_43254);
nor U44944 (N_44944,N_43580,N_43399);
xnor U44945 (N_44945,N_43338,N_43076);
xnor U44946 (N_44946,N_43632,N_43586);
nand U44947 (N_44947,N_43690,N_43650);
or U44948 (N_44948,N_43783,N_43437);
nor U44949 (N_44949,N_43843,N_43924);
nand U44950 (N_44950,N_43888,N_43119);
nand U44951 (N_44951,N_43628,N_43783);
or U44952 (N_44952,N_43336,N_43781);
or U44953 (N_44953,N_43626,N_43030);
nand U44954 (N_44954,N_43488,N_43771);
nor U44955 (N_44955,N_43407,N_43109);
nor U44956 (N_44956,N_43339,N_43056);
and U44957 (N_44957,N_43302,N_43129);
and U44958 (N_44958,N_43622,N_43579);
nand U44959 (N_44959,N_43061,N_43575);
nand U44960 (N_44960,N_43284,N_43938);
nor U44961 (N_44961,N_43200,N_43438);
and U44962 (N_44962,N_43424,N_43527);
or U44963 (N_44963,N_43235,N_43552);
nand U44964 (N_44964,N_43431,N_43928);
nand U44965 (N_44965,N_43527,N_43132);
nand U44966 (N_44966,N_43145,N_43651);
xnor U44967 (N_44967,N_43732,N_43495);
nor U44968 (N_44968,N_43314,N_43327);
nand U44969 (N_44969,N_43921,N_43323);
nand U44970 (N_44970,N_43214,N_43444);
nor U44971 (N_44971,N_43436,N_43635);
nor U44972 (N_44972,N_43490,N_43781);
and U44973 (N_44973,N_43671,N_43666);
nand U44974 (N_44974,N_43262,N_43300);
xor U44975 (N_44975,N_43154,N_43293);
xnor U44976 (N_44976,N_43374,N_43387);
or U44977 (N_44977,N_43244,N_43837);
nor U44978 (N_44978,N_43972,N_43114);
nor U44979 (N_44979,N_43319,N_43903);
nand U44980 (N_44980,N_43831,N_43913);
nor U44981 (N_44981,N_43516,N_43401);
nand U44982 (N_44982,N_43690,N_43762);
nor U44983 (N_44983,N_43880,N_43772);
or U44984 (N_44984,N_43178,N_43763);
nor U44985 (N_44985,N_43729,N_43736);
and U44986 (N_44986,N_43056,N_43193);
or U44987 (N_44987,N_43466,N_43608);
nor U44988 (N_44988,N_43053,N_43487);
nor U44989 (N_44989,N_43559,N_43940);
nor U44990 (N_44990,N_43575,N_43449);
or U44991 (N_44991,N_43996,N_43765);
nand U44992 (N_44992,N_43361,N_43111);
xnor U44993 (N_44993,N_43464,N_43200);
xnor U44994 (N_44994,N_43859,N_43326);
xor U44995 (N_44995,N_43151,N_43183);
xor U44996 (N_44996,N_43169,N_43692);
xnor U44997 (N_44997,N_43951,N_43276);
nand U44998 (N_44998,N_43249,N_43303);
or U44999 (N_44999,N_43373,N_43160);
xnor U45000 (N_45000,N_44161,N_44425);
xor U45001 (N_45001,N_44881,N_44244);
and U45002 (N_45002,N_44458,N_44112);
nor U45003 (N_45003,N_44405,N_44487);
and U45004 (N_45004,N_44948,N_44786);
nand U45005 (N_45005,N_44764,N_44566);
nor U45006 (N_45006,N_44263,N_44024);
nor U45007 (N_45007,N_44247,N_44351);
xor U45008 (N_45008,N_44571,N_44479);
nor U45009 (N_45009,N_44876,N_44751);
nor U45010 (N_45010,N_44445,N_44505);
and U45011 (N_45011,N_44086,N_44229);
or U45012 (N_45012,N_44653,N_44712);
xnor U45013 (N_45013,N_44152,N_44611);
nor U45014 (N_45014,N_44107,N_44612);
nand U45015 (N_45015,N_44676,N_44070);
nor U45016 (N_45016,N_44499,N_44727);
nor U45017 (N_45017,N_44713,N_44057);
nand U45018 (N_45018,N_44928,N_44327);
nand U45019 (N_45019,N_44300,N_44201);
nor U45020 (N_45020,N_44678,N_44624);
xor U45021 (N_45021,N_44944,N_44698);
nand U45022 (N_45022,N_44397,N_44210);
and U45023 (N_45023,N_44343,N_44549);
or U45024 (N_45024,N_44789,N_44480);
or U45025 (N_45025,N_44128,N_44004);
or U45026 (N_45026,N_44158,N_44124);
nand U45027 (N_45027,N_44842,N_44598);
nor U45028 (N_45028,N_44752,N_44440);
nor U45029 (N_45029,N_44335,N_44819);
nand U45030 (N_45030,N_44980,N_44531);
nor U45031 (N_45031,N_44707,N_44272);
nor U45032 (N_45032,N_44682,N_44400);
or U45033 (N_45033,N_44172,N_44448);
or U45034 (N_45034,N_44242,N_44204);
nand U45035 (N_45035,N_44364,N_44562);
or U45036 (N_45036,N_44492,N_44741);
and U45037 (N_45037,N_44062,N_44469);
xnor U45038 (N_45038,N_44625,N_44932);
and U45039 (N_45039,N_44567,N_44546);
nor U45040 (N_45040,N_44514,N_44910);
or U45041 (N_45041,N_44403,N_44260);
xnor U45042 (N_45042,N_44889,N_44494);
nor U45043 (N_45043,N_44563,N_44643);
or U45044 (N_45044,N_44040,N_44880);
nor U45045 (N_45045,N_44541,N_44329);
nand U45046 (N_45046,N_44601,N_44583);
or U45047 (N_45047,N_44388,N_44095);
and U45048 (N_45048,N_44166,N_44017);
nor U45049 (N_45049,N_44331,N_44780);
nand U45050 (N_45050,N_44305,N_44600);
and U45051 (N_45051,N_44162,N_44317);
or U45052 (N_45052,N_44042,N_44451);
xnor U45053 (N_45053,N_44279,N_44964);
nor U45054 (N_45054,N_44695,N_44486);
nand U45055 (N_45055,N_44491,N_44150);
nand U45056 (N_45056,N_44831,N_44389);
nand U45057 (N_45057,N_44907,N_44387);
nor U45058 (N_45058,N_44287,N_44737);
nor U45059 (N_45059,N_44079,N_44334);
nand U45060 (N_45060,N_44515,N_44614);
and U45061 (N_45061,N_44700,N_44168);
or U45062 (N_45062,N_44946,N_44560);
or U45063 (N_45063,N_44116,N_44374);
and U45064 (N_45064,N_44544,N_44794);
xor U45065 (N_45065,N_44885,N_44288);
and U45066 (N_45066,N_44209,N_44103);
nor U45067 (N_45067,N_44308,N_44901);
nor U45068 (N_45068,N_44963,N_44019);
and U45069 (N_45069,N_44465,N_44576);
nor U45070 (N_45070,N_44996,N_44188);
xnor U45071 (N_45071,N_44856,N_44132);
and U45072 (N_45072,N_44022,N_44319);
and U45073 (N_45073,N_44850,N_44268);
and U45074 (N_45074,N_44313,N_44981);
xnor U45075 (N_45075,N_44587,N_44151);
xor U45076 (N_45076,N_44453,N_44809);
and U45077 (N_45077,N_44130,N_44489);
or U45078 (N_45078,N_44767,N_44048);
nand U45079 (N_45079,N_44165,N_44519);
xnor U45080 (N_45080,N_44952,N_44140);
or U45081 (N_45081,N_44690,N_44344);
nand U45082 (N_45082,N_44868,N_44740);
xor U45083 (N_45083,N_44482,N_44959);
nor U45084 (N_45084,N_44258,N_44339);
and U45085 (N_45085,N_44854,N_44609);
or U45086 (N_45086,N_44729,N_44355);
nor U45087 (N_45087,N_44921,N_44264);
and U45088 (N_45088,N_44621,N_44187);
nor U45089 (N_45089,N_44592,N_44820);
nor U45090 (N_45090,N_44018,N_44096);
xor U45091 (N_45091,N_44315,N_44723);
xor U45092 (N_45092,N_44163,N_44449);
or U45093 (N_45093,N_44380,N_44495);
nor U45094 (N_45094,N_44628,N_44424);
and U45095 (N_45095,N_44270,N_44671);
nor U45096 (N_45096,N_44685,N_44147);
xor U45097 (N_45097,N_44537,N_44431);
nor U45098 (N_45098,N_44568,N_44212);
xnor U45099 (N_45099,N_44955,N_44659);
nor U45100 (N_45100,N_44362,N_44386);
or U45101 (N_45101,N_44186,N_44990);
xnor U45102 (N_45102,N_44021,N_44845);
nor U45103 (N_45103,N_44524,N_44573);
nor U45104 (N_45104,N_44904,N_44146);
xor U45105 (N_45105,N_44805,N_44254);
xor U45106 (N_45106,N_44010,N_44966);
nor U45107 (N_45107,N_44255,N_44784);
nor U45108 (N_45108,N_44135,N_44848);
or U45109 (N_45109,N_44199,N_44858);
xor U45110 (N_45110,N_44768,N_44131);
or U45111 (N_45111,N_44615,N_44454);
xor U45112 (N_45112,N_44687,N_44092);
or U45113 (N_45113,N_44450,N_44629);
and U45114 (N_45114,N_44940,N_44093);
or U45115 (N_45115,N_44087,N_44510);
and U45116 (N_45116,N_44657,N_44935);
xnor U45117 (N_45117,N_44861,N_44281);
and U45118 (N_45118,N_44617,N_44117);
xor U45119 (N_45119,N_44763,N_44719);
nor U45120 (N_45120,N_44137,N_44083);
nand U45121 (N_45121,N_44797,N_44363);
xnor U45122 (N_45122,N_44227,N_44637);
or U45123 (N_45123,N_44972,N_44641);
nand U45124 (N_45124,N_44872,N_44666);
nand U45125 (N_45125,N_44539,N_44304);
xor U45126 (N_45126,N_44520,N_44558);
or U45127 (N_45127,N_44839,N_44860);
or U45128 (N_45128,N_44989,N_44336);
nand U45129 (N_45129,N_44297,N_44938);
nor U45130 (N_45130,N_44826,N_44538);
xor U45131 (N_45131,N_44274,N_44230);
xor U45132 (N_45132,N_44542,N_44060);
or U45133 (N_45133,N_44728,N_44059);
nand U45134 (N_45134,N_44604,N_44123);
or U45135 (N_45135,N_44591,N_44547);
nand U45136 (N_45136,N_44138,N_44870);
or U45137 (N_45137,N_44957,N_44704);
nor U45138 (N_45138,N_44200,N_44613);
and U45139 (N_45139,N_44661,N_44973);
and U45140 (N_45140,N_44867,N_44250);
xor U45141 (N_45141,N_44159,N_44974);
nor U45142 (N_45142,N_44559,N_44055);
xor U45143 (N_45143,N_44912,N_44792);
nor U45144 (N_45144,N_44894,N_44762);
or U45145 (N_45145,N_44667,N_44085);
nor U45146 (N_45146,N_44370,N_44345);
nor U45147 (N_45147,N_44550,N_44597);
xnor U45148 (N_45148,N_44032,N_44090);
or U45149 (N_45149,N_44222,N_44808);
nand U45150 (N_45150,N_44824,N_44337);
or U45151 (N_45151,N_44954,N_44501);
or U45152 (N_45152,N_44841,N_44012);
or U45153 (N_45153,N_44652,N_44000);
nor U45154 (N_45154,N_44960,N_44474);
xnor U45155 (N_45155,N_44094,N_44978);
and U45156 (N_45156,N_44496,N_44065);
and U45157 (N_45157,N_44303,N_44468);
nor U45158 (N_45158,N_44338,N_44804);
or U45159 (N_45159,N_44582,N_44655);
or U45160 (N_45160,N_44787,N_44461);
and U45161 (N_45161,N_44895,N_44324);
and U45162 (N_45162,N_44711,N_44008);
nand U45163 (N_45163,N_44193,N_44239);
or U45164 (N_45164,N_44377,N_44834);
nand U45165 (N_45165,N_44790,N_44905);
nor U45166 (N_45166,N_44349,N_44234);
and U45167 (N_45167,N_44699,N_44314);
xnor U45168 (N_45168,N_44758,N_44523);
nor U45169 (N_45169,N_44354,N_44703);
nor U45170 (N_45170,N_44545,N_44476);
and U45171 (N_45171,N_44185,N_44577);
nand U45172 (N_45172,N_44005,N_44899);
xnor U45173 (N_45173,N_44077,N_44836);
and U45174 (N_45174,N_44580,N_44748);
nand U45175 (N_45175,N_44100,N_44962);
nand U45176 (N_45176,N_44033,N_44432);
nand U45177 (N_45177,N_44635,N_44992);
nor U45178 (N_45178,N_44738,N_44777);
nor U45179 (N_45179,N_44434,N_44988);
xor U45180 (N_45180,N_44656,N_44235);
xnor U45181 (N_45181,N_44673,N_44706);
nand U45182 (N_45182,N_44633,N_44067);
nor U45183 (N_45183,N_44717,N_44155);
xor U45184 (N_45184,N_44419,N_44616);
nor U45185 (N_45185,N_44183,N_44348);
xnor U45186 (N_45186,N_44759,N_44267);
and U45187 (N_45187,N_44099,N_44481);
xnor U45188 (N_45188,N_44731,N_44642);
nand U45189 (N_45189,N_44154,N_44463);
xor U45190 (N_45190,N_44669,N_44007);
nand U45191 (N_45191,N_44423,N_44284);
xnor U45192 (N_45192,N_44073,N_44755);
or U45193 (N_45193,N_44555,N_44645);
nand U45194 (N_45194,N_44498,N_44618);
or U45195 (N_45195,N_44392,N_44620);
xnor U45196 (N_45196,N_44192,N_44770);
and U45197 (N_45197,N_44754,N_44488);
xnor U45198 (N_45198,N_44879,N_44925);
xnor U45199 (N_45199,N_44599,N_44701);
or U45200 (N_45200,N_44252,N_44157);
xnor U45201 (N_45201,N_44502,N_44811);
xnor U45202 (N_45202,N_44565,N_44941);
xnor U45203 (N_45203,N_44142,N_44749);
and U45204 (N_45204,N_44716,N_44353);
xnor U45205 (N_45205,N_44529,N_44736);
and U45206 (N_45206,N_44467,N_44245);
xnor U45207 (N_45207,N_44833,N_44970);
nor U45208 (N_45208,N_44361,N_44821);
xnor U45209 (N_45209,N_44603,N_44002);
and U45210 (N_45210,N_44807,N_44174);
or U45211 (N_45211,N_44816,N_44511);
nor U45212 (N_45212,N_44779,N_44991);
xor U45213 (N_45213,N_44995,N_44898);
nand U45214 (N_45214,N_44735,N_44799);
nand U45215 (N_45215,N_44847,N_44822);
or U45216 (N_45216,N_44217,N_44875);
nor U45217 (N_45217,N_44223,N_44294);
and U45218 (N_45218,N_44051,N_44477);
or U45219 (N_45219,N_44893,N_44594);
and U45220 (N_45220,N_44081,N_44001);
nand U45221 (N_45221,N_44564,N_44459);
nor U45222 (N_45222,N_44182,N_44806);
xor U45223 (N_45223,N_44082,N_44038);
and U45224 (N_45224,N_44967,N_44983);
nor U45225 (N_45225,N_44115,N_44177);
and U45226 (N_45226,N_44730,N_44293);
nor U45227 (N_45227,N_44114,N_44072);
nor U45228 (N_45228,N_44061,N_44466);
and U45229 (N_45229,N_44026,N_44111);
xnor U45230 (N_45230,N_44902,N_44148);
nand U45231 (N_45231,N_44859,N_44049);
xor U45232 (N_45232,N_44009,N_44757);
or U45233 (N_45233,N_44526,N_44385);
and U45234 (N_45234,N_44307,N_44862);
and U45235 (N_45235,N_44760,N_44534);
nand U45236 (N_45236,N_44064,N_44918);
nand U45237 (N_45237,N_44634,N_44118);
or U45238 (N_45238,N_44674,N_44164);
nor U45239 (N_45239,N_44887,N_44993);
nand U45240 (N_45240,N_44586,N_44874);
nand U45241 (N_45241,N_44399,N_44034);
and U45242 (N_45242,N_44373,N_44369);
nand U45243 (N_45243,N_44382,N_44088);
or U45244 (N_45244,N_44979,N_44843);
and U45245 (N_45245,N_44406,N_44823);
nand U45246 (N_45246,N_44144,N_44427);
or U45247 (N_45247,N_44950,N_44470);
or U45248 (N_45248,N_44815,N_44548);
nor U45249 (N_45249,N_44922,N_44143);
xnor U45250 (N_45250,N_44483,N_44783);
and U45251 (N_45251,N_44202,N_44746);
xnor U45252 (N_45252,N_44189,N_44068);
nand U45253 (N_45253,N_44043,N_44953);
or U45254 (N_45254,N_44683,N_44198);
or U45255 (N_45255,N_44692,N_44984);
xnor U45256 (N_45256,N_44773,N_44825);
nand U45257 (N_45257,N_44769,N_44404);
or U45258 (N_45258,N_44251,N_44133);
nor U45259 (N_45259,N_44640,N_44551);
xor U45260 (N_45260,N_44662,N_44347);
nand U45261 (N_45261,N_44041,N_44851);
nand U45262 (N_45262,N_44460,N_44897);
xor U45263 (N_45263,N_44378,N_44688);
and U45264 (N_45264,N_44595,N_44302);
xor U45265 (N_45265,N_44054,N_44999);
xnor U45266 (N_45266,N_44679,N_44761);
nor U45267 (N_45267,N_44398,N_44195);
xnor U45268 (N_45268,N_44119,N_44422);
nand U45269 (N_45269,N_44827,N_44330);
nand U45270 (N_45270,N_44426,N_44947);
or U45271 (N_45271,N_44101,N_44771);
or U45272 (N_45272,N_44273,N_44225);
nand U45273 (N_45273,N_44853,N_44791);
or U45274 (N_45274,N_44718,N_44240);
or U45275 (N_45275,N_44462,N_44122);
xor U45276 (N_45276,N_44838,N_44788);
nor U45277 (N_45277,N_44015,N_44365);
nor U45278 (N_45278,N_44803,N_44610);
xor U45279 (N_45279,N_44917,N_44321);
nand U45280 (N_45280,N_44167,N_44722);
or U45281 (N_45281,N_44888,N_44141);
nor U45282 (N_45282,N_44360,N_44277);
or U45283 (N_45283,N_44710,N_44063);
nor U45284 (N_45284,N_44631,N_44873);
and U45285 (N_45285,N_44997,N_44923);
or U45286 (N_45286,N_44607,N_44105);
or U45287 (N_45287,N_44023,N_44934);
xnor U45288 (N_45288,N_44817,N_44914);
xor U45289 (N_45289,N_44578,N_44396);
or U45290 (N_45290,N_44249,N_44725);
nor U45291 (N_45291,N_44261,N_44197);
nor U45292 (N_45292,N_44056,N_44484);
or U45293 (N_45293,N_44664,N_44203);
or U45294 (N_45294,N_44689,N_44569);
nor U45295 (N_45295,N_44556,N_44646);
nor U45296 (N_45296,N_44557,N_44913);
xor U45297 (N_45297,N_44310,N_44175);
xor U45298 (N_45298,N_44686,N_44346);
nor U45299 (N_45299,N_44207,N_44437);
nand U45300 (N_45300,N_44025,N_44069);
nor U45301 (N_45301,N_44160,N_44194);
xor U45302 (N_45302,N_44464,N_44776);
or U45303 (N_45303,N_44016,N_44906);
nand U45304 (N_45304,N_44801,N_44285);
nand U45305 (N_45305,N_44774,N_44903);
and U45306 (N_45306,N_44781,N_44412);
or U45307 (N_45307,N_44052,N_44433);
xnor U45308 (N_45308,N_44106,N_44417);
or U45309 (N_45309,N_44246,N_44933);
and U45310 (N_45310,N_44213,N_44224);
xnor U45311 (N_45311,N_44253,N_44596);
nor U45312 (N_45312,N_44608,N_44532);
and U45313 (N_45313,N_44473,N_44226);
xor U45314 (N_45314,N_44184,N_44765);
xor U45315 (N_45315,N_44295,N_44920);
or U45316 (N_45316,N_44886,N_44572);
xor U45317 (N_45317,N_44512,N_44011);
nor U45318 (N_45318,N_44931,N_44503);
or U45319 (N_45319,N_44724,N_44593);
or U45320 (N_45320,N_44844,N_44058);
nand U45321 (N_45321,N_44371,N_44930);
and U45322 (N_45322,N_44402,N_44219);
nor U45323 (N_45323,N_44316,N_44878);
or U45324 (N_45324,N_44518,N_44084);
xnor U45325 (N_45325,N_44782,N_44332);
and U45326 (N_45326,N_44139,N_44756);
nor U45327 (N_45327,N_44733,N_44156);
or U45328 (N_45328,N_44527,N_44436);
nor U45329 (N_45329,N_44091,N_44421);
or U45330 (N_45330,N_44098,N_44446);
nand U45331 (N_45331,N_44985,N_44681);
and U45332 (N_45332,N_44649,N_44383);
nand U45333 (N_45333,N_44866,N_44630);
xor U45334 (N_45334,N_44720,N_44742);
and U45335 (N_45335,N_44283,N_44909);
or U45336 (N_45336,N_44376,N_44136);
nand U45337 (N_45337,N_44668,N_44452);
and U45338 (N_45338,N_44619,N_44180);
or U45339 (N_45339,N_44409,N_44663);
nor U45340 (N_45340,N_44588,N_44442);
xnor U45341 (N_45341,N_44029,N_44037);
and U45342 (N_45342,N_44220,N_44636);
and U45343 (N_45343,N_44290,N_44120);
nand U45344 (N_45344,N_44750,N_44228);
nand U45345 (N_45345,N_44949,N_44233);
xnor U45346 (N_45346,N_44726,N_44301);
or U45347 (N_45347,N_44916,N_44884);
nand U45348 (N_45348,N_44271,N_44044);
or U45349 (N_45349,N_44855,N_44456);
nand U45350 (N_45350,N_44053,N_44020);
and U45351 (N_45351,N_44795,N_44071);
xnor U45352 (N_45352,N_44214,N_44936);
nand U45353 (N_45353,N_44149,N_44863);
nand U45354 (N_45354,N_44248,N_44413);
nor U45355 (N_45355,N_44046,N_44677);
xnor U45356 (N_45356,N_44178,N_44575);
nor U45357 (N_45357,N_44318,N_44036);
nand U45358 (N_45358,N_44325,N_44030);
or U45359 (N_45359,N_44262,N_44408);
nor U45360 (N_45360,N_44181,N_44766);
nand U45361 (N_45361,N_44929,N_44455);
or U45362 (N_45362,N_44179,N_44420);
nor U45363 (N_45363,N_44753,N_44366);
or U45364 (N_45364,N_44394,N_44939);
nand U45365 (N_45365,N_44622,N_44145);
nor U45366 (N_45366,N_44775,N_44076);
xor U45367 (N_45367,N_44702,N_44384);
xor U45368 (N_45368,N_44237,N_44977);
and U45369 (N_45369,N_44987,N_44798);
xor U45370 (N_45370,N_44435,N_44943);
nor U45371 (N_45371,N_44444,N_44414);
xor U45372 (N_45372,N_44958,N_44418);
or U45373 (N_45373,N_44975,N_44439);
and U45374 (N_45374,N_44080,N_44299);
xnor U45375 (N_45375,N_44045,N_44238);
or U45376 (N_45376,N_44506,N_44994);
and U45377 (N_45377,N_44896,N_44109);
nor U45378 (N_45378,N_44956,N_44543);
or U45379 (N_45379,N_44243,N_44694);
and U45380 (N_45380,N_44734,N_44108);
and U45381 (N_45381,N_44328,N_44937);
nor U45382 (N_45382,N_44497,N_44153);
nor U45383 (N_45383,N_44323,N_44357);
nor U45384 (N_45384,N_44216,N_44047);
and U45385 (N_45385,N_44393,N_44276);
and U45386 (N_45386,N_44478,N_44513);
xor U45387 (N_45387,N_44554,N_44982);
nand U45388 (N_45388,N_44102,N_44951);
nor U45389 (N_45389,N_44129,N_44684);
and U45390 (N_45390,N_44078,N_44352);
nand U45391 (N_45391,N_44697,N_44428);
or U45392 (N_45392,N_44006,N_44340);
or U45393 (N_45393,N_44035,N_44648);
nand U45394 (N_45394,N_44693,N_44778);
or U45395 (N_45395,N_44410,N_44113);
or U45396 (N_45396,N_44915,N_44971);
xor U45397 (N_45397,N_44176,N_44533);
and U45398 (N_45398,N_44430,N_44840);
or U45399 (N_45399,N_44900,N_44127);
or U45400 (N_45400,N_44632,N_44945);
or U45401 (N_45401,N_44490,N_44375);
or U45402 (N_45402,N_44236,N_44522);
nand U45403 (N_45403,N_44257,N_44651);
or U45404 (N_45404,N_44475,N_44919);
nand U45405 (N_45405,N_44626,N_44832);
and U45406 (N_45406,N_44882,N_44368);
or U45407 (N_45407,N_44976,N_44221);
nor U45408 (N_45408,N_44606,N_44709);
xnor U45409 (N_45409,N_44411,N_44013);
nor U45410 (N_45410,N_44961,N_44416);
xnor U45411 (N_45411,N_44359,N_44282);
nor U45412 (N_45412,N_44849,N_44381);
xor U45413 (N_45413,N_44561,N_44259);
or U45414 (N_45414,N_44747,N_44097);
xnor U45415 (N_45415,N_44443,N_44828);
and U45416 (N_45416,N_44367,N_44715);
xor U45417 (N_45417,N_44802,N_44291);
xor U45418 (N_45418,N_44732,N_44066);
and U45419 (N_45419,N_44275,N_44877);
and U45420 (N_45420,N_44320,N_44472);
or U45421 (N_45421,N_44280,N_44846);
nor U45422 (N_45422,N_44891,N_44171);
or U45423 (N_45423,N_44438,N_44721);
nand U45424 (N_45424,N_44341,N_44675);
or U45425 (N_45425,N_44865,N_44027);
xor U45426 (N_45426,N_44342,N_44585);
nand U45427 (N_45427,N_44785,N_44638);
and U45428 (N_45428,N_44206,N_44517);
or U45429 (N_45429,N_44926,N_44714);
or U45430 (N_45430,N_44516,N_44772);
nor U45431 (N_45431,N_44391,N_44326);
or U45432 (N_45432,N_44218,N_44708);
and U45433 (N_45433,N_44289,N_44231);
xor U45434 (N_45434,N_44509,N_44508);
or U45435 (N_45435,N_44447,N_44208);
nor U45436 (N_45436,N_44627,N_44215);
nor U45437 (N_45437,N_44590,N_44521);
xor U45438 (N_45438,N_44528,N_44269);
or U45439 (N_45439,N_44670,N_44892);
or U45440 (N_45440,N_44191,N_44356);
or U45441 (N_45441,N_44837,N_44504);
xor U45442 (N_45442,N_44211,N_44278);
nand U45443 (N_45443,N_44390,N_44372);
nor U45444 (N_45444,N_44457,N_44969);
and U45445 (N_45445,N_44471,N_44170);
xor U45446 (N_45446,N_44535,N_44395);
or U45447 (N_45447,N_44232,N_44003);
or U45448 (N_45448,N_44286,N_44441);
and U45449 (N_45449,N_44241,N_44639);
xnor U45450 (N_45450,N_44089,N_44800);
and U45451 (N_45451,N_44818,N_44813);
xor U45452 (N_45452,N_44552,N_44744);
or U45453 (N_45453,N_44312,N_44500);
nor U45454 (N_45454,N_44190,N_44830);
or U45455 (N_45455,N_44968,N_44415);
nand U45456 (N_45456,N_44266,N_44796);
nor U45457 (N_45457,N_44650,N_44743);
nor U45458 (N_45458,N_44829,N_44265);
and U45459 (N_45459,N_44379,N_44986);
nor U45460 (N_45460,N_44574,N_44605);
or U45461 (N_45461,N_44965,N_44014);
and U45462 (N_45462,N_44835,N_44298);
or U45463 (N_45463,N_44814,N_44908);
xnor U45464 (N_45464,N_44584,N_44602);
or U45465 (N_45465,N_44536,N_44665);
or U45466 (N_45466,N_44104,N_44196);
nand U45467 (N_45467,N_44857,N_44696);
xor U45468 (N_45468,N_44306,N_44660);
nor U45469 (N_45469,N_44871,N_44942);
nand U45470 (N_45470,N_44869,N_44644);
or U45471 (N_45471,N_44296,N_44075);
xnor U45472 (N_45472,N_44169,N_44309);
or U45473 (N_45473,N_44173,N_44126);
nand U45474 (N_45474,N_44493,N_44256);
nand U45475 (N_45475,N_44553,N_44658);
and U45476 (N_45476,N_44031,N_44407);
and U45477 (N_45477,N_44647,N_44927);
or U45478 (N_45478,N_44121,N_44540);
xor U45479 (N_45479,N_44311,N_44134);
or U45480 (N_45480,N_44292,N_44205);
xor U45481 (N_45481,N_44333,N_44911);
and U45482 (N_45482,N_44864,N_44350);
nand U45483 (N_45483,N_44812,N_44623);
and U45484 (N_45484,N_44883,N_44570);
nand U45485 (N_45485,N_44589,N_44810);
and U45486 (N_45486,N_44485,N_44998);
nand U45487 (N_45487,N_44507,N_44525);
or U45488 (N_45488,N_44705,N_44890);
xnor U45489 (N_45489,N_44745,N_44793);
or U45490 (N_45490,N_44039,N_44672);
xor U45491 (N_45491,N_44924,N_44358);
or U45492 (N_45492,N_44429,N_44050);
nand U45493 (N_45493,N_44852,N_44654);
and U45494 (N_45494,N_44074,N_44691);
nand U45495 (N_45495,N_44579,N_44028);
and U45496 (N_45496,N_44125,N_44739);
or U45497 (N_45497,N_44581,N_44110);
or U45498 (N_45498,N_44680,N_44530);
nand U45499 (N_45499,N_44322,N_44401);
nand U45500 (N_45500,N_44148,N_44809);
and U45501 (N_45501,N_44147,N_44977);
or U45502 (N_45502,N_44352,N_44607);
nand U45503 (N_45503,N_44062,N_44539);
nand U45504 (N_45504,N_44179,N_44377);
nor U45505 (N_45505,N_44440,N_44412);
xor U45506 (N_45506,N_44082,N_44591);
nand U45507 (N_45507,N_44008,N_44092);
nor U45508 (N_45508,N_44190,N_44384);
nand U45509 (N_45509,N_44387,N_44014);
and U45510 (N_45510,N_44198,N_44018);
or U45511 (N_45511,N_44838,N_44230);
nor U45512 (N_45512,N_44618,N_44300);
nand U45513 (N_45513,N_44933,N_44572);
or U45514 (N_45514,N_44692,N_44138);
nand U45515 (N_45515,N_44980,N_44066);
nor U45516 (N_45516,N_44459,N_44087);
nand U45517 (N_45517,N_44627,N_44317);
and U45518 (N_45518,N_44860,N_44128);
xnor U45519 (N_45519,N_44074,N_44278);
or U45520 (N_45520,N_44673,N_44331);
nor U45521 (N_45521,N_44839,N_44192);
nand U45522 (N_45522,N_44848,N_44053);
nor U45523 (N_45523,N_44933,N_44032);
nand U45524 (N_45524,N_44205,N_44410);
nand U45525 (N_45525,N_44346,N_44054);
and U45526 (N_45526,N_44562,N_44242);
and U45527 (N_45527,N_44409,N_44792);
or U45528 (N_45528,N_44839,N_44008);
xnor U45529 (N_45529,N_44908,N_44793);
nand U45530 (N_45530,N_44114,N_44724);
nor U45531 (N_45531,N_44321,N_44529);
nor U45532 (N_45532,N_44816,N_44669);
or U45533 (N_45533,N_44766,N_44590);
or U45534 (N_45534,N_44072,N_44725);
nand U45535 (N_45535,N_44426,N_44224);
nor U45536 (N_45536,N_44581,N_44970);
nand U45537 (N_45537,N_44937,N_44589);
xnor U45538 (N_45538,N_44680,N_44415);
xnor U45539 (N_45539,N_44858,N_44890);
or U45540 (N_45540,N_44649,N_44158);
and U45541 (N_45541,N_44581,N_44615);
xor U45542 (N_45542,N_44975,N_44395);
and U45543 (N_45543,N_44563,N_44296);
xor U45544 (N_45544,N_44020,N_44332);
or U45545 (N_45545,N_44946,N_44642);
or U45546 (N_45546,N_44473,N_44200);
xor U45547 (N_45547,N_44371,N_44250);
nor U45548 (N_45548,N_44355,N_44052);
nand U45549 (N_45549,N_44151,N_44304);
nor U45550 (N_45550,N_44286,N_44106);
or U45551 (N_45551,N_44827,N_44548);
or U45552 (N_45552,N_44555,N_44444);
nor U45553 (N_45553,N_44792,N_44078);
nand U45554 (N_45554,N_44197,N_44205);
nand U45555 (N_45555,N_44999,N_44066);
nand U45556 (N_45556,N_44363,N_44924);
or U45557 (N_45557,N_44840,N_44392);
or U45558 (N_45558,N_44451,N_44327);
nand U45559 (N_45559,N_44397,N_44934);
nor U45560 (N_45560,N_44980,N_44550);
or U45561 (N_45561,N_44106,N_44891);
nand U45562 (N_45562,N_44092,N_44703);
nor U45563 (N_45563,N_44218,N_44330);
xor U45564 (N_45564,N_44602,N_44861);
nand U45565 (N_45565,N_44206,N_44992);
and U45566 (N_45566,N_44481,N_44932);
and U45567 (N_45567,N_44307,N_44879);
xnor U45568 (N_45568,N_44819,N_44245);
or U45569 (N_45569,N_44483,N_44020);
and U45570 (N_45570,N_44027,N_44586);
or U45571 (N_45571,N_44048,N_44530);
nand U45572 (N_45572,N_44227,N_44687);
xor U45573 (N_45573,N_44409,N_44847);
xor U45574 (N_45574,N_44437,N_44273);
and U45575 (N_45575,N_44926,N_44827);
or U45576 (N_45576,N_44769,N_44738);
nand U45577 (N_45577,N_44107,N_44141);
nor U45578 (N_45578,N_44618,N_44018);
nor U45579 (N_45579,N_44297,N_44107);
or U45580 (N_45580,N_44184,N_44983);
xor U45581 (N_45581,N_44928,N_44425);
nor U45582 (N_45582,N_44412,N_44490);
and U45583 (N_45583,N_44176,N_44166);
and U45584 (N_45584,N_44791,N_44305);
xnor U45585 (N_45585,N_44505,N_44509);
or U45586 (N_45586,N_44412,N_44409);
nor U45587 (N_45587,N_44449,N_44789);
or U45588 (N_45588,N_44152,N_44843);
xnor U45589 (N_45589,N_44756,N_44277);
or U45590 (N_45590,N_44320,N_44689);
nor U45591 (N_45591,N_44823,N_44027);
and U45592 (N_45592,N_44595,N_44316);
and U45593 (N_45593,N_44654,N_44837);
nor U45594 (N_45594,N_44424,N_44775);
nand U45595 (N_45595,N_44708,N_44681);
xor U45596 (N_45596,N_44599,N_44773);
and U45597 (N_45597,N_44176,N_44380);
and U45598 (N_45598,N_44123,N_44305);
xnor U45599 (N_45599,N_44090,N_44086);
nand U45600 (N_45600,N_44505,N_44969);
or U45601 (N_45601,N_44791,N_44481);
xnor U45602 (N_45602,N_44516,N_44115);
or U45603 (N_45603,N_44614,N_44323);
or U45604 (N_45604,N_44606,N_44398);
or U45605 (N_45605,N_44668,N_44683);
nor U45606 (N_45606,N_44866,N_44186);
nand U45607 (N_45607,N_44441,N_44814);
nand U45608 (N_45608,N_44823,N_44014);
nand U45609 (N_45609,N_44430,N_44196);
nand U45610 (N_45610,N_44907,N_44775);
and U45611 (N_45611,N_44074,N_44942);
nor U45612 (N_45612,N_44349,N_44148);
xor U45613 (N_45613,N_44202,N_44434);
nand U45614 (N_45614,N_44380,N_44938);
nand U45615 (N_45615,N_44154,N_44331);
or U45616 (N_45616,N_44212,N_44783);
and U45617 (N_45617,N_44043,N_44924);
xor U45618 (N_45618,N_44727,N_44126);
and U45619 (N_45619,N_44068,N_44095);
nor U45620 (N_45620,N_44929,N_44227);
or U45621 (N_45621,N_44171,N_44972);
nand U45622 (N_45622,N_44410,N_44952);
and U45623 (N_45623,N_44195,N_44479);
nor U45624 (N_45624,N_44929,N_44763);
nor U45625 (N_45625,N_44775,N_44874);
or U45626 (N_45626,N_44808,N_44638);
or U45627 (N_45627,N_44813,N_44627);
nand U45628 (N_45628,N_44266,N_44684);
xnor U45629 (N_45629,N_44496,N_44385);
xnor U45630 (N_45630,N_44078,N_44704);
nor U45631 (N_45631,N_44430,N_44230);
and U45632 (N_45632,N_44988,N_44528);
and U45633 (N_45633,N_44437,N_44333);
nand U45634 (N_45634,N_44178,N_44261);
nand U45635 (N_45635,N_44286,N_44449);
xnor U45636 (N_45636,N_44902,N_44423);
nor U45637 (N_45637,N_44032,N_44576);
nand U45638 (N_45638,N_44363,N_44131);
nor U45639 (N_45639,N_44312,N_44628);
nand U45640 (N_45640,N_44267,N_44623);
xnor U45641 (N_45641,N_44575,N_44339);
nor U45642 (N_45642,N_44801,N_44470);
or U45643 (N_45643,N_44512,N_44285);
nor U45644 (N_45644,N_44450,N_44588);
nor U45645 (N_45645,N_44662,N_44972);
and U45646 (N_45646,N_44955,N_44565);
nand U45647 (N_45647,N_44435,N_44209);
or U45648 (N_45648,N_44422,N_44220);
nand U45649 (N_45649,N_44103,N_44106);
or U45650 (N_45650,N_44887,N_44376);
nor U45651 (N_45651,N_44814,N_44412);
or U45652 (N_45652,N_44356,N_44069);
xnor U45653 (N_45653,N_44033,N_44656);
xor U45654 (N_45654,N_44379,N_44827);
or U45655 (N_45655,N_44635,N_44930);
xnor U45656 (N_45656,N_44779,N_44802);
nand U45657 (N_45657,N_44550,N_44780);
nor U45658 (N_45658,N_44218,N_44479);
and U45659 (N_45659,N_44807,N_44910);
nor U45660 (N_45660,N_44809,N_44267);
nor U45661 (N_45661,N_44948,N_44814);
or U45662 (N_45662,N_44336,N_44361);
or U45663 (N_45663,N_44371,N_44115);
xnor U45664 (N_45664,N_44053,N_44558);
or U45665 (N_45665,N_44527,N_44615);
or U45666 (N_45666,N_44239,N_44834);
xnor U45667 (N_45667,N_44280,N_44611);
or U45668 (N_45668,N_44906,N_44972);
xnor U45669 (N_45669,N_44807,N_44109);
xnor U45670 (N_45670,N_44948,N_44822);
or U45671 (N_45671,N_44367,N_44270);
nor U45672 (N_45672,N_44609,N_44618);
and U45673 (N_45673,N_44909,N_44790);
and U45674 (N_45674,N_44776,N_44593);
xor U45675 (N_45675,N_44417,N_44020);
or U45676 (N_45676,N_44492,N_44149);
xnor U45677 (N_45677,N_44621,N_44358);
nand U45678 (N_45678,N_44305,N_44909);
or U45679 (N_45679,N_44125,N_44975);
nor U45680 (N_45680,N_44356,N_44032);
nand U45681 (N_45681,N_44904,N_44753);
and U45682 (N_45682,N_44252,N_44731);
or U45683 (N_45683,N_44014,N_44296);
nor U45684 (N_45684,N_44223,N_44940);
xnor U45685 (N_45685,N_44535,N_44424);
or U45686 (N_45686,N_44191,N_44681);
nor U45687 (N_45687,N_44724,N_44651);
xor U45688 (N_45688,N_44808,N_44381);
and U45689 (N_45689,N_44147,N_44338);
nor U45690 (N_45690,N_44238,N_44390);
and U45691 (N_45691,N_44709,N_44836);
or U45692 (N_45692,N_44223,N_44376);
and U45693 (N_45693,N_44285,N_44386);
or U45694 (N_45694,N_44651,N_44977);
xnor U45695 (N_45695,N_44023,N_44206);
or U45696 (N_45696,N_44556,N_44091);
nand U45697 (N_45697,N_44430,N_44846);
or U45698 (N_45698,N_44640,N_44567);
or U45699 (N_45699,N_44580,N_44427);
nand U45700 (N_45700,N_44519,N_44760);
nand U45701 (N_45701,N_44098,N_44449);
nor U45702 (N_45702,N_44435,N_44592);
and U45703 (N_45703,N_44817,N_44527);
or U45704 (N_45704,N_44387,N_44481);
nor U45705 (N_45705,N_44275,N_44455);
and U45706 (N_45706,N_44722,N_44546);
nand U45707 (N_45707,N_44451,N_44436);
and U45708 (N_45708,N_44376,N_44044);
nand U45709 (N_45709,N_44260,N_44352);
and U45710 (N_45710,N_44525,N_44364);
xor U45711 (N_45711,N_44840,N_44198);
or U45712 (N_45712,N_44547,N_44223);
nand U45713 (N_45713,N_44780,N_44271);
and U45714 (N_45714,N_44343,N_44376);
and U45715 (N_45715,N_44472,N_44988);
nor U45716 (N_45716,N_44541,N_44325);
and U45717 (N_45717,N_44160,N_44782);
or U45718 (N_45718,N_44130,N_44424);
and U45719 (N_45719,N_44795,N_44557);
nor U45720 (N_45720,N_44571,N_44404);
nand U45721 (N_45721,N_44648,N_44739);
nor U45722 (N_45722,N_44286,N_44073);
and U45723 (N_45723,N_44514,N_44435);
and U45724 (N_45724,N_44010,N_44776);
or U45725 (N_45725,N_44939,N_44895);
nand U45726 (N_45726,N_44424,N_44592);
or U45727 (N_45727,N_44927,N_44690);
and U45728 (N_45728,N_44791,N_44013);
or U45729 (N_45729,N_44822,N_44846);
xnor U45730 (N_45730,N_44034,N_44287);
or U45731 (N_45731,N_44437,N_44752);
nor U45732 (N_45732,N_44389,N_44281);
or U45733 (N_45733,N_44234,N_44795);
xnor U45734 (N_45734,N_44055,N_44189);
xnor U45735 (N_45735,N_44417,N_44939);
nor U45736 (N_45736,N_44650,N_44145);
nor U45737 (N_45737,N_44721,N_44391);
or U45738 (N_45738,N_44052,N_44274);
or U45739 (N_45739,N_44348,N_44775);
nor U45740 (N_45740,N_44747,N_44665);
or U45741 (N_45741,N_44491,N_44949);
or U45742 (N_45742,N_44109,N_44492);
nand U45743 (N_45743,N_44433,N_44233);
or U45744 (N_45744,N_44530,N_44801);
xor U45745 (N_45745,N_44913,N_44698);
or U45746 (N_45746,N_44439,N_44267);
nor U45747 (N_45747,N_44818,N_44913);
nor U45748 (N_45748,N_44311,N_44416);
nor U45749 (N_45749,N_44188,N_44755);
and U45750 (N_45750,N_44912,N_44252);
and U45751 (N_45751,N_44076,N_44792);
or U45752 (N_45752,N_44832,N_44143);
nand U45753 (N_45753,N_44670,N_44099);
or U45754 (N_45754,N_44892,N_44317);
nor U45755 (N_45755,N_44720,N_44574);
nor U45756 (N_45756,N_44419,N_44954);
or U45757 (N_45757,N_44457,N_44523);
nor U45758 (N_45758,N_44035,N_44062);
or U45759 (N_45759,N_44724,N_44600);
nor U45760 (N_45760,N_44158,N_44201);
and U45761 (N_45761,N_44139,N_44742);
nor U45762 (N_45762,N_44544,N_44591);
and U45763 (N_45763,N_44111,N_44169);
nor U45764 (N_45764,N_44207,N_44291);
nor U45765 (N_45765,N_44667,N_44778);
or U45766 (N_45766,N_44357,N_44362);
or U45767 (N_45767,N_44723,N_44391);
and U45768 (N_45768,N_44172,N_44828);
nand U45769 (N_45769,N_44560,N_44066);
xor U45770 (N_45770,N_44076,N_44997);
nand U45771 (N_45771,N_44650,N_44771);
xnor U45772 (N_45772,N_44399,N_44424);
or U45773 (N_45773,N_44333,N_44509);
nor U45774 (N_45774,N_44303,N_44520);
nor U45775 (N_45775,N_44437,N_44851);
nand U45776 (N_45776,N_44839,N_44351);
nor U45777 (N_45777,N_44373,N_44786);
or U45778 (N_45778,N_44340,N_44176);
nor U45779 (N_45779,N_44008,N_44232);
nor U45780 (N_45780,N_44690,N_44360);
nand U45781 (N_45781,N_44326,N_44551);
and U45782 (N_45782,N_44208,N_44510);
xnor U45783 (N_45783,N_44647,N_44278);
nor U45784 (N_45784,N_44442,N_44999);
and U45785 (N_45785,N_44699,N_44658);
and U45786 (N_45786,N_44640,N_44041);
nand U45787 (N_45787,N_44728,N_44299);
or U45788 (N_45788,N_44123,N_44357);
nor U45789 (N_45789,N_44812,N_44322);
and U45790 (N_45790,N_44403,N_44535);
xor U45791 (N_45791,N_44159,N_44877);
nor U45792 (N_45792,N_44936,N_44793);
and U45793 (N_45793,N_44112,N_44065);
xor U45794 (N_45794,N_44999,N_44080);
nand U45795 (N_45795,N_44293,N_44888);
and U45796 (N_45796,N_44636,N_44128);
and U45797 (N_45797,N_44620,N_44618);
xor U45798 (N_45798,N_44837,N_44325);
xor U45799 (N_45799,N_44224,N_44110);
or U45800 (N_45800,N_44005,N_44653);
and U45801 (N_45801,N_44688,N_44041);
nand U45802 (N_45802,N_44023,N_44893);
nand U45803 (N_45803,N_44229,N_44772);
nor U45804 (N_45804,N_44352,N_44357);
nor U45805 (N_45805,N_44095,N_44628);
nor U45806 (N_45806,N_44271,N_44584);
and U45807 (N_45807,N_44828,N_44878);
xnor U45808 (N_45808,N_44908,N_44341);
nor U45809 (N_45809,N_44179,N_44899);
and U45810 (N_45810,N_44273,N_44412);
nand U45811 (N_45811,N_44333,N_44524);
xnor U45812 (N_45812,N_44611,N_44252);
xnor U45813 (N_45813,N_44321,N_44642);
or U45814 (N_45814,N_44440,N_44703);
nor U45815 (N_45815,N_44199,N_44966);
and U45816 (N_45816,N_44305,N_44516);
nand U45817 (N_45817,N_44615,N_44030);
nor U45818 (N_45818,N_44061,N_44029);
xnor U45819 (N_45819,N_44600,N_44887);
nor U45820 (N_45820,N_44468,N_44383);
xnor U45821 (N_45821,N_44639,N_44944);
xor U45822 (N_45822,N_44374,N_44200);
nor U45823 (N_45823,N_44339,N_44473);
or U45824 (N_45824,N_44697,N_44619);
xor U45825 (N_45825,N_44393,N_44081);
xor U45826 (N_45826,N_44445,N_44847);
and U45827 (N_45827,N_44588,N_44984);
nand U45828 (N_45828,N_44405,N_44281);
or U45829 (N_45829,N_44846,N_44964);
or U45830 (N_45830,N_44927,N_44305);
nand U45831 (N_45831,N_44764,N_44006);
nor U45832 (N_45832,N_44503,N_44030);
xnor U45833 (N_45833,N_44943,N_44503);
xor U45834 (N_45834,N_44898,N_44796);
nor U45835 (N_45835,N_44108,N_44225);
nor U45836 (N_45836,N_44526,N_44200);
and U45837 (N_45837,N_44136,N_44169);
and U45838 (N_45838,N_44201,N_44654);
and U45839 (N_45839,N_44848,N_44927);
nor U45840 (N_45840,N_44040,N_44331);
xor U45841 (N_45841,N_44026,N_44046);
or U45842 (N_45842,N_44716,N_44854);
nor U45843 (N_45843,N_44426,N_44341);
xor U45844 (N_45844,N_44543,N_44455);
nand U45845 (N_45845,N_44781,N_44349);
nor U45846 (N_45846,N_44585,N_44077);
nor U45847 (N_45847,N_44038,N_44930);
nand U45848 (N_45848,N_44089,N_44746);
and U45849 (N_45849,N_44978,N_44905);
nand U45850 (N_45850,N_44723,N_44456);
nand U45851 (N_45851,N_44646,N_44369);
xor U45852 (N_45852,N_44656,N_44539);
and U45853 (N_45853,N_44473,N_44819);
nand U45854 (N_45854,N_44598,N_44600);
nor U45855 (N_45855,N_44166,N_44662);
nor U45856 (N_45856,N_44563,N_44739);
nand U45857 (N_45857,N_44324,N_44517);
and U45858 (N_45858,N_44641,N_44275);
and U45859 (N_45859,N_44873,N_44289);
or U45860 (N_45860,N_44090,N_44917);
or U45861 (N_45861,N_44700,N_44195);
and U45862 (N_45862,N_44961,N_44619);
or U45863 (N_45863,N_44348,N_44634);
nand U45864 (N_45864,N_44145,N_44613);
nor U45865 (N_45865,N_44953,N_44991);
and U45866 (N_45866,N_44101,N_44897);
or U45867 (N_45867,N_44982,N_44148);
and U45868 (N_45868,N_44879,N_44106);
xnor U45869 (N_45869,N_44078,N_44596);
or U45870 (N_45870,N_44894,N_44260);
nand U45871 (N_45871,N_44316,N_44057);
and U45872 (N_45872,N_44697,N_44173);
or U45873 (N_45873,N_44539,N_44460);
nand U45874 (N_45874,N_44162,N_44363);
nor U45875 (N_45875,N_44209,N_44281);
or U45876 (N_45876,N_44606,N_44815);
nand U45877 (N_45877,N_44702,N_44389);
nand U45878 (N_45878,N_44907,N_44309);
nand U45879 (N_45879,N_44837,N_44124);
nand U45880 (N_45880,N_44869,N_44945);
nor U45881 (N_45881,N_44458,N_44133);
nand U45882 (N_45882,N_44701,N_44964);
nor U45883 (N_45883,N_44680,N_44770);
xnor U45884 (N_45884,N_44545,N_44634);
and U45885 (N_45885,N_44272,N_44571);
xnor U45886 (N_45886,N_44742,N_44258);
nand U45887 (N_45887,N_44960,N_44290);
or U45888 (N_45888,N_44421,N_44857);
xnor U45889 (N_45889,N_44535,N_44841);
xnor U45890 (N_45890,N_44017,N_44264);
nor U45891 (N_45891,N_44790,N_44926);
and U45892 (N_45892,N_44538,N_44728);
xnor U45893 (N_45893,N_44734,N_44500);
nor U45894 (N_45894,N_44318,N_44012);
and U45895 (N_45895,N_44964,N_44818);
nand U45896 (N_45896,N_44185,N_44581);
or U45897 (N_45897,N_44295,N_44701);
xor U45898 (N_45898,N_44837,N_44248);
or U45899 (N_45899,N_44482,N_44609);
or U45900 (N_45900,N_44368,N_44118);
and U45901 (N_45901,N_44666,N_44810);
and U45902 (N_45902,N_44573,N_44326);
nand U45903 (N_45903,N_44503,N_44046);
xor U45904 (N_45904,N_44909,N_44063);
nand U45905 (N_45905,N_44460,N_44853);
nand U45906 (N_45906,N_44893,N_44990);
xor U45907 (N_45907,N_44207,N_44967);
or U45908 (N_45908,N_44976,N_44224);
nand U45909 (N_45909,N_44748,N_44262);
or U45910 (N_45910,N_44836,N_44760);
xor U45911 (N_45911,N_44131,N_44853);
and U45912 (N_45912,N_44861,N_44633);
xnor U45913 (N_45913,N_44019,N_44923);
nor U45914 (N_45914,N_44554,N_44098);
xnor U45915 (N_45915,N_44518,N_44213);
nor U45916 (N_45916,N_44088,N_44945);
nand U45917 (N_45917,N_44139,N_44658);
and U45918 (N_45918,N_44035,N_44695);
or U45919 (N_45919,N_44740,N_44266);
xor U45920 (N_45920,N_44872,N_44477);
xor U45921 (N_45921,N_44473,N_44776);
or U45922 (N_45922,N_44409,N_44174);
nand U45923 (N_45923,N_44877,N_44293);
or U45924 (N_45924,N_44385,N_44054);
nor U45925 (N_45925,N_44411,N_44903);
or U45926 (N_45926,N_44397,N_44079);
nand U45927 (N_45927,N_44620,N_44962);
xnor U45928 (N_45928,N_44413,N_44338);
and U45929 (N_45929,N_44600,N_44492);
and U45930 (N_45930,N_44182,N_44702);
nand U45931 (N_45931,N_44667,N_44075);
xor U45932 (N_45932,N_44925,N_44466);
xnor U45933 (N_45933,N_44990,N_44224);
nand U45934 (N_45934,N_44015,N_44465);
nand U45935 (N_45935,N_44735,N_44436);
nand U45936 (N_45936,N_44866,N_44805);
or U45937 (N_45937,N_44437,N_44886);
and U45938 (N_45938,N_44924,N_44810);
and U45939 (N_45939,N_44633,N_44142);
and U45940 (N_45940,N_44690,N_44028);
or U45941 (N_45941,N_44015,N_44738);
nand U45942 (N_45942,N_44760,N_44135);
nand U45943 (N_45943,N_44282,N_44468);
nor U45944 (N_45944,N_44480,N_44436);
xnor U45945 (N_45945,N_44299,N_44290);
or U45946 (N_45946,N_44902,N_44598);
nand U45947 (N_45947,N_44017,N_44399);
or U45948 (N_45948,N_44653,N_44850);
nor U45949 (N_45949,N_44841,N_44580);
or U45950 (N_45950,N_44067,N_44350);
and U45951 (N_45951,N_44061,N_44641);
xor U45952 (N_45952,N_44521,N_44958);
and U45953 (N_45953,N_44865,N_44721);
or U45954 (N_45954,N_44468,N_44410);
xor U45955 (N_45955,N_44023,N_44833);
or U45956 (N_45956,N_44294,N_44959);
or U45957 (N_45957,N_44027,N_44325);
or U45958 (N_45958,N_44404,N_44060);
nor U45959 (N_45959,N_44470,N_44254);
nand U45960 (N_45960,N_44637,N_44927);
or U45961 (N_45961,N_44460,N_44432);
nor U45962 (N_45962,N_44143,N_44306);
or U45963 (N_45963,N_44760,N_44622);
xnor U45964 (N_45964,N_44414,N_44105);
nand U45965 (N_45965,N_44456,N_44858);
or U45966 (N_45966,N_44036,N_44264);
nor U45967 (N_45967,N_44824,N_44797);
and U45968 (N_45968,N_44086,N_44636);
or U45969 (N_45969,N_44806,N_44130);
xor U45970 (N_45970,N_44788,N_44830);
nand U45971 (N_45971,N_44801,N_44768);
nand U45972 (N_45972,N_44215,N_44380);
or U45973 (N_45973,N_44654,N_44727);
or U45974 (N_45974,N_44724,N_44094);
xnor U45975 (N_45975,N_44090,N_44033);
and U45976 (N_45976,N_44057,N_44044);
and U45977 (N_45977,N_44644,N_44202);
nand U45978 (N_45978,N_44764,N_44463);
nor U45979 (N_45979,N_44024,N_44387);
nor U45980 (N_45980,N_44470,N_44174);
or U45981 (N_45981,N_44493,N_44769);
or U45982 (N_45982,N_44720,N_44037);
nand U45983 (N_45983,N_44307,N_44173);
nand U45984 (N_45984,N_44617,N_44333);
xor U45985 (N_45985,N_44604,N_44692);
or U45986 (N_45986,N_44806,N_44415);
nand U45987 (N_45987,N_44251,N_44960);
or U45988 (N_45988,N_44762,N_44211);
nor U45989 (N_45989,N_44240,N_44453);
xnor U45990 (N_45990,N_44198,N_44731);
xor U45991 (N_45991,N_44119,N_44864);
nor U45992 (N_45992,N_44394,N_44378);
nor U45993 (N_45993,N_44197,N_44202);
nor U45994 (N_45994,N_44291,N_44316);
and U45995 (N_45995,N_44037,N_44129);
nand U45996 (N_45996,N_44247,N_44040);
nor U45997 (N_45997,N_44833,N_44653);
nand U45998 (N_45998,N_44331,N_44883);
and U45999 (N_45999,N_44736,N_44154);
and U46000 (N_46000,N_45790,N_45597);
xor U46001 (N_46001,N_45074,N_45512);
and U46002 (N_46002,N_45288,N_45735);
or U46003 (N_46003,N_45690,N_45822);
nand U46004 (N_46004,N_45547,N_45862);
and U46005 (N_46005,N_45410,N_45158);
xnor U46006 (N_46006,N_45255,N_45305);
or U46007 (N_46007,N_45326,N_45328);
nor U46008 (N_46008,N_45975,N_45230);
nor U46009 (N_46009,N_45083,N_45107);
or U46010 (N_46010,N_45519,N_45032);
xor U46011 (N_46011,N_45659,N_45495);
and U46012 (N_46012,N_45123,N_45800);
xor U46013 (N_46013,N_45769,N_45589);
nand U46014 (N_46014,N_45275,N_45139);
and U46015 (N_46015,N_45730,N_45660);
or U46016 (N_46016,N_45220,N_45142);
xor U46017 (N_46017,N_45842,N_45023);
nor U46018 (N_46018,N_45063,N_45049);
nand U46019 (N_46019,N_45093,N_45056);
nor U46020 (N_46020,N_45043,N_45183);
xor U46021 (N_46021,N_45670,N_45219);
nor U46022 (N_46022,N_45529,N_45084);
nand U46023 (N_46023,N_45118,N_45710);
nand U46024 (N_46024,N_45907,N_45443);
or U46025 (N_46025,N_45169,N_45454);
and U46026 (N_46026,N_45173,N_45828);
nand U46027 (N_46027,N_45613,N_45696);
nor U46028 (N_46028,N_45112,N_45198);
nand U46029 (N_46029,N_45532,N_45464);
and U46030 (N_46030,N_45188,N_45815);
or U46031 (N_46031,N_45967,N_45362);
and U46032 (N_46032,N_45944,N_45590);
nand U46033 (N_46033,N_45177,N_45037);
and U46034 (N_46034,N_45683,N_45436);
or U46035 (N_46035,N_45217,N_45915);
or U46036 (N_46036,N_45951,N_45916);
or U46037 (N_46037,N_45665,N_45076);
xor U46038 (N_46038,N_45736,N_45044);
and U46039 (N_46039,N_45920,N_45634);
or U46040 (N_46040,N_45026,N_45666);
nor U46041 (N_46041,N_45997,N_45749);
xnor U46042 (N_46042,N_45178,N_45005);
nand U46043 (N_46043,N_45854,N_45941);
xnor U46044 (N_46044,N_45126,N_45408);
and U46045 (N_46045,N_45880,N_45066);
or U46046 (N_46046,N_45896,N_45294);
nand U46047 (N_46047,N_45162,N_45671);
xor U46048 (N_46048,N_45085,N_45246);
nand U46049 (N_46049,N_45416,N_45164);
or U46050 (N_46050,N_45424,N_45349);
xnor U46051 (N_46051,N_45447,N_45639);
and U46052 (N_46052,N_45563,N_45306);
or U46053 (N_46053,N_45705,N_45000);
xor U46054 (N_46054,N_45797,N_45831);
or U46055 (N_46055,N_45558,N_45500);
nand U46056 (N_46056,N_45174,N_45546);
nor U46057 (N_46057,N_45817,N_45419);
and U46058 (N_46058,N_45475,N_45391);
nor U46059 (N_46059,N_45003,N_45324);
nand U46060 (N_46060,N_45273,N_45816);
nor U46061 (N_46061,N_45827,N_45763);
or U46062 (N_46062,N_45726,N_45157);
or U46063 (N_46063,N_45926,N_45439);
nor U46064 (N_46064,N_45276,N_45473);
and U46065 (N_46065,N_45082,N_45572);
nor U46066 (N_46066,N_45526,N_45140);
nor U46067 (N_46067,N_45366,N_45741);
or U46068 (N_46068,N_45132,N_45320);
nor U46069 (N_46069,N_45394,N_45938);
nand U46070 (N_46070,N_45646,N_45611);
nand U46071 (N_46071,N_45434,N_45963);
nor U46072 (N_46072,N_45562,N_45829);
xor U46073 (N_46073,N_45502,N_45090);
nor U46074 (N_46074,N_45861,N_45950);
and U46075 (N_46075,N_45773,N_45708);
and U46076 (N_46076,N_45048,N_45633);
nand U46077 (N_46077,N_45551,N_45190);
or U46078 (N_46078,N_45612,N_45755);
and U46079 (N_46079,N_45565,N_45717);
nor U46080 (N_46080,N_45588,N_45598);
and U46081 (N_46081,N_45307,N_45069);
and U46082 (N_46082,N_45898,N_45834);
xor U46083 (N_46083,N_45935,N_45490);
or U46084 (N_46084,N_45619,N_45878);
nor U46085 (N_46085,N_45549,N_45550);
xnor U46086 (N_46086,N_45095,N_45658);
and U46087 (N_46087,N_45218,N_45413);
or U46088 (N_46088,N_45728,N_45238);
nor U46089 (N_46089,N_45936,N_45160);
xor U46090 (N_46090,N_45046,N_45807);
nand U46091 (N_46091,N_45165,N_45061);
and U46092 (N_46092,N_45811,N_45144);
or U46093 (N_46093,N_45301,N_45461);
nor U46094 (N_46094,N_45882,N_45632);
nor U46095 (N_46095,N_45592,N_45538);
nor U46096 (N_46096,N_45647,N_45501);
or U46097 (N_46097,N_45575,N_45956);
xnor U46098 (N_46098,N_45333,N_45035);
and U46099 (N_46099,N_45561,N_45367);
nor U46100 (N_46100,N_45297,N_45930);
or U46101 (N_46101,N_45459,N_45928);
xnor U46102 (N_46102,N_45285,N_45693);
or U46103 (N_46103,N_45480,N_45688);
nand U46104 (N_46104,N_45743,N_45168);
or U46105 (N_46105,N_45020,N_45376);
or U46106 (N_46106,N_45681,N_45989);
or U46107 (N_46107,N_45718,N_45729);
nor U46108 (N_46108,N_45809,N_45591);
or U46109 (N_46109,N_45931,N_45466);
or U46110 (N_46110,N_45117,N_45796);
or U46111 (N_46111,N_45054,N_45483);
and U46112 (N_46112,N_45962,N_45282);
xnor U46113 (N_46113,N_45689,N_45787);
and U46114 (N_46114,N_45456,N_45848);
nand U46115 (N_46115,N_45389,N_45120);
nor U46116 (N_46116,N_45296,N_45175);
and U46117 (N_46117,N_45096,N_45953);
xor U46118 (N_46118,N_45396,N_45525);
xnor U46119 (N_46119,N_45996,N_45694);
or U46120 (N_46120,N_45616,N_45476);
xnor U46121 (N_46121,N_45628,N_45203);
and U46122 (N_46122,N_45109,N_45171);
and U46123 (N_46123,N_45040,N_45300);
nand U46124 (N_46124,N_45978,N_45406);
nand U46125 (N_46125,N_45852,N_45783);
or U46126 (N_46126,N_45554,N_45062);
or U46127 (N_46127,N_45824,N_45888);
nand U46128 (N_46128,N_45498,N_45627);
and U46129 (N_46129,N_45474,N_45445);
xnor U46130 (N_46130,N_45785,N_45341);
nand U46131 (N_46131,N_45031,N_45704);
and U46132 (N_46132,N_45847,N_45653);
xnor U46133 (N_46133,N_45594,N_45354);
xnor U46134 (N_46134,N_45489,N_45912);
or U46135 (N_46135,N_45645,N_45423);
xnor U46136 (N_46136,N_45004,N_45334);
nand U46137 (N_46137,N_45793,N_45499);
nand U46138 (N_46138,N_45957,N_45292);
nor U46139 (N_46139,N_45271,N_45511);
nor U46140 (N_46140,N_45640,N_45414);
and U46141 (N_46141,N_45135,N_45733);
nand U46142 (N_46142,N_45960,N_45313);
nand U46143 (N_46143,N_45648,N_45885);
xor U46144 (N_46144,N_45195,N_45053);
and U46145 (N_46145,N_45876,N_45421);
xor U46146 (N_46146,N_45161,N_45460);
or U46147 (N_46147,N_45223,N_45855);
xnor U46148 (N_46148,N_45317,N_45662);
nand U46149 (N_46149,N_45227,N_45411);
nand U46150 (N_46150,N_45578,N_45825);
nand U46151 (N_46151,N_45196,N_45780);
nor U46152 (N_46152,N_45014,N_45448);
nand U46153 (N_46153,N_45493,N_45969);
xnor U46154 (N_46154,N_45994,N_45116);
nor U46155 (N_46155,N_45266,N_45172);
and U46156 (N_46156,N_45064,N_45644);
nor U46157 (N_46157,N_45843,N_45030);
xor U46158 (N_46158,N_45853,N_45260);
xnor U46159 (N_46159,N_45510,N_45257);
and U46160 (N_46160,N_45622,N_45819);
nor U46161 (N_46161,N_45833,N_45587);
xor U46162 (N_46162,N_45965,N_45901);
nor U46163 (N_46163,N_45202,N_45373);
nor U46164 (N_46164,N_45954,N_45034);
or U46165 (N_46165,N_45678,N_45206);
and U46166 (N_46166,N_45702,N_45012);
or U46167 (N_46167,N_45740,N_45208);
nand U46168 (N_46168,N_45544,N_45103);
or U46169 (N_46169,N_45939,N_45539);
xor U46170 (N_46170,N_45264,N_45985);
nor U46171 (N_46171,N_45802,N_45570);
nand U46172 (N_46172,N_45451,N_45826);
xnor U46173 (N_46173,N_45184,N_45378);
xnor U46174 (N_46174,N_45309,N_45060);
nor U46175 (N_46175,N_45509,N_45075);
nor U46176 (N_46176,N_45959,N_45810);
xor U46177 (N_46177,N_45984,N_45929);
nand U46178 (N_46178,N_45318,N_45786);
nand U46179 (N_46179,N_45441,N_45747);
xor U46180 (N_46180,N_45642,N_45637);
nor U46181 (N_46181,N_45656,N_45618);
or U46182 (N_46182,N_45988,N_45152);
nand U46183 (N_46183,N_45993,N_45185);
xor U46184 (N_46184,N_45820,N_45222);
nor U46185 (N_46185,N_45527,N_45521);
or U46186 (N_46186,N_45721,N_45484);
nand U46187 (N_46187,N_45187,N_45105);
nor U46188 (N_46188,N_45018,N_45601);
nand U46189 (N_46189,N_45906,N_45463);
or U46190 (N_46190,N_45148,N_45114);
nor U46191 (N_46191,N_45359,N_45432);
nor U46192 (N_46192,N_45340,N_45478);
nor U46193 (N_46193,N_45002,N_45774);
nand U46194 (N_46194,N_45277,N_45290);
nor U46195 (N_46195,N_45345,N_45615);
and U46196 (N_46196,N_45207,N_45086);
and U46197 (N_46197,N_45189,N_45269);
nor U46198 (N_46198,N_45315,N_45390);
or U46199 (N_46199,N_45585,N_45111);
nor U46200 (N_46200,N_45039,N_45137);
or U46201 (N_46201,N_45823,N_45245);
or U46202 (N_46202,N_45009,N_45837);
nor U46203 (N_46203,N_45363,N_45050);
xnor U46204 (N_46204,N_45332,N_45055);
nand U46205 (N_46205,N_45404,N_45537);
nor U46206 (N_46206,N_45961,N_45518);
and U46207 (N_46207,N_45351,N_45194);
nor U46208 (N_46208,N_45635,N_45435);
and U46209 (N_46209,N_45933,N_45553);
and U46210 (N_46210,N_45347,N_45893);
nor U46211 (N_46211,N_45364,N_45361);
or U46212 (N_46212,N_45750,N_45279);
nor U46213 (N_46213,N_45709,N_45455);
and U46214 (N_46214,N_45609,N_45520);
or U46215 (N_46215,N_45052,N_45453);
nand U46216 (N_46216,N_45346,N_45143);
nand U46217 (N_46217,N_45712,N_45652);
and U46218 (N_46218,N_45580,N_45159);
xor U46219 (N_46219,N_45803,N_45754);
or U46220 (N_46220,N_45564,N_45059);
and U46221 (N_46221,N_45081,N_45226);
nand U46222 (N_46222,N_45507,N_45923);
and U46223 (N_46223,N_45851,N_45374);
nand U46224 (N_46224,N_45291,N_45779);
and U46225 (N_46225,N_45121,N_45504);
or U46226 (N_46226,N_45398,N_45886);
or U46227 (N_46227,N_45497,N_45182);
xor U46228 (N_46228,N_45119,N_45995);
nor U46229 (N_46229,N_45595,N_45088);
nand U46230 (N_46230,N_45732,N_45677);
nor U46231 (N_46231,N_45706,N_45968);
nor U46232 (N_46232,N_45267,N_45479);
and U46233 (N_46233,N_45765,N_45813);
nand U46234 (N_46234,N_45127,N_45180);
nand U46235 (N_46235,N_45228,N_45225);
nand U46236 (N_46236,N_45715,N_45981);
and U46237 (N_46237,N_45428,N_45600);
and U46238 (N_46238,N_45099,N_45673);
nand U46239 (N_46239,N_45940,N_45725);
or U46240 (N_46240,N_45734,N_45908);
xor U46241 (N_46241,N_45760,N_45496);
nand U46242 (N_46242,N_45372,N_45900);
nor U46243 (N_46243,N_45610,N_45723);
and U46244 (N_46244,N_45259,N_45442);
nor U46245 (N_46245,N_45982,N_45412);
xor U46246 (N_46246,N_45249,N_45714);
nand U46247 (N_46247,N_45231,N_45884);
nand U46248 (N_46248,N_45685,N_45946);
xnor U46249 (N_46249,N_45626,N_45883);
nand U46250 (N_46250,N_45097,N_45716);
and U46251 (N_46251,N_45859,N_45767);
nand U46252 (N_46252,N_45524,N_45641);
xor U46253 (N_46253,N_45649,N_45557);
nand U46254 (N_46254,N_45235,N_45329);
and U46255 (N_46255,N_45007,N_45452);
or U46256 (N_46256,N_45759,N_45293);
nand U46257 (N_46257,N_45087,N_45395);
xor U46258 (N_46258,N_45571,N_45166);
or U46259 (N_46259,N_45348,N_45323);
and U46260 (N_46260,N_45200,N_45025);
nand U46261 (N_46261,N_45910,N_45698);
xnor U46262 (N_46262,N_45402,N_45895);
xor U46263 (N_46263,N_45289,N_45427);
or U46264 (N_46264,N_45617,N_45192);
xnor U46265 (N_46265,N_45624,N_45661);
xor U46266 (N_46266,N_45552,N_45253);
or U46267 (N_46267,N_45927,N_45719);
and U46268 (N_46268,N_45322,N_45577);
xnor U46269 (N_46269,N_45979,N_45115);
xor U46270 (N_46270,N_45417,N_45457);
and U46271 (N_46271,N_45091,N_45836);
and U46272 (N_46272,N_45674,N_45687);
xor U46273 (N_46273,N_45942,N_45776);
xor U46274 (N_46274,N_45299,N_45835);
nor U46275 (N_46275,N_45806,N_45244);
and U46276 (N_46276,N_45338,N_45782);
and U46277 (N_46277,N_45711,N_45596);
xor U46278 (N_46278,N_45492,N_45679);
nor U46279 (N_46279,N_45124,N_45420);
nand U46280 (N_46280,N_45379,N_45657);
and U46281 (N_46281,N_45250,N_45021);
nand U46282 (N_46282,N_45605,N_45738);
nor U46283 (N_46283,N_45934,N_45327);
or U46284 (N_46284,N_45889,N_45278);
nand U46285 (N_46285,N_45757,N_45872);
and U46286 (N_46286,N_45943,N_45789);
nor U46287 (N_46287,N_45270,N_45205);
and U46288 (N_46288,N_45446,N_45958);
nand U46289 (N_46289,N_45151,N_45233);
nor U46290 (N_46290,N_45752,N_45625);
nor U46291 (N_46291,N_45422,N_45543);
xnor U46292 (N_46292,N_45080,N_45254);
and U46293 (N_46293,N_45703,N_45745);
nand U46294 (N_46294,N_45481,N_45176);
nor U46295 (N_46295,N_45153,N_45016);
or U46296 (N_46296,N_45795,N_45821);
xnor U46297 (N_46297,N_45232,N_45983);
or U46298 (N_46298,N_45899,N_45573);
or U46299 (N_46299,N_45316,N_45579);
nand U46300 (N_46300,N_45869,N_45990);
nand U46301 (N_46301,N_45211,N_45130);
xor U46302 (N_46302,N_45154,N_45098);
nand U46303 (N_46303,N_45970,N_45197);
and U46304 (N_46304,N_45506,N_45343);
and U46305 (N_46305,N_45686,N_45241);
nor U46306 (N_46306,N_45067,N_45638);
nand U46307 (N_46307,N_45672,N_45015);
xor U46308 (N_46308,N_45469,N_45545);
or U46309 (N_46309,N_45017,N_45891);
and U46310 (N_46310,N_45758,N_45280);
nand U46311 (N_46311,N_45472,N_45339);
nor U46312 (N_46312,N_45149,N_45071);
or U46313 (N_46313,N_45146,N_45494);
nor U46314 (N_46314,N_45914,N_45358);
and U46315 (N_46315,N_45314,N_45281);
nor U46316 (N_46316,N_45860,N_45801);
and U46317 (N_46317,N_45513,N_45430);
or U46318 (N_46318,N_45503,N_45304);
nand U46319 (N_46319,N_45337,N_45991);
xor U46320 (N_46320,N_45384,N_45488);
and U46321 (N_46321,N_45163,N_45385);
xor U46322 (N_46322,N_45866,N_45794);
and U46323 (N_46323,N_45251,N_45027);
nor U46324 (N_46324,N_45330,N_45470);
or U46325 (N_46325,N_45382,N_45193);
nand U46326 (N_46326,N_45237,N_45375);
and U46327 (N_46327,N_45636,N_45089);
xor U46328 (N_46328,N_45047,N_45136);
nand U46329 (N_46329,N_45778,N_45764);
xnor U46330 (N_46330,N_45236,N_45485);
or U46331 (N_46331,N_45058,N_45429);
or U46332 (N_46332,N_45234,N_45684);
nand U46333 (N_46333,N_45917,N_45409);
nand U46334 (N_46334,N_45849,N_45041);
nor U46335 (N_46335,N_45945,N_45310);
nor U46336 (N_46336,N_45630,N_45437);
or U46337 (N_46337,N_45042,N_45535);
nor U46338 (N_46338,N_45751,N_45101);
nand U46339 (N_46339,N_45283,N_45212);
nor U46340 (N_46340,N_45073,N_45643);
xor U46341 (N_46341,N_45312,N_45010);
nand U46342 (N_46342,N_45737,N_45365);
xor U46343 (N_46343,N_45937,N_45350);
nand U46344 (N_46344,N_45383,N_45971);
xnor U46345 (N_46345,N_45516,N_45788);
nor U46346 (N_46346,N_45077,N_45458);
nand U46347 (N_46347,N_45569,N_45070);
or U46348 (N_46348,N_45224,N_45426);
nand U46349 (N_46349,N_45584,N_45128);
nand U46350 (N_46350,N_45263,N_45675);
or U46351 (N_46351,N_45201,N_45331);
nand U46352 (N_46352,N_45792,N_45602);
and U46353 (N_46353,N_45746,N_45909);
nor U46354 (N_46354,N_45482,N_45287);
xor U46355 (N_46355,N_45804,N_45676);
nand U46356 (N_46356,N_45321,N_45522);
and U46357 (N_46357,N_45371,N_45808);
and U46358 (N_46358,N_45863,N_45134);
and U46359 (N_46359,N_45298,N_45770);
or U46360 (N_46360,N_45839,N_45431);
or U46361 (N_46361,N_45667,N_45742);
xnor U46362 (N_46362,N_45523,N_45336);
xnor U46363 (N_46363,N_45812,N_45799);
xnor U46364 (N_46364,N_45845,N_45925);
and U46365 (N_46365,N_45604,N_45621);
xnor U46366 (N_46366,N_45870,N_45556);
or U46367 (N_46367,N_45387,N_45664);
nor U46368 (N_46368,N_45311,N_45401);
nor U46369 (N_46369,N_45104,N_45548);
or U46370 (N_46370,N_45145,N_45583);
nand U46371 (N_46371,N_45724,N_45707);
nand U46372 (N_46372,N_45980,N_45045);
and U46373 (N_46373,N_45798,N_45850);
nand U46374 (N_46374,N_45840,N_45302);
and U46375 (N_46375,N_45620,N_45654);
nand U46376 (N_46376,N_45904,N_45964);
or U46377 (N_46377,N_45874,N_45335);
nand U46378 (N_46378,N_45036,N_45922);
nor U46379 (N_46379,N_45614,N_45897);
nor U46380 (N_46380,N_45303,N_45213);
or U46381 (N_46381,N_45533,N_45753);
and U46382 (N_46382,N_45932,N_45008);
or U46383 (N_46383,N_45695,N_45924);
nand U46384 (N_46384,N_45720,N_45381);
and U46385 (N_46385,N_45508,N_45186);
nand U46386 (N_46386,N_45541,N_45902);
xor U46387 (N_46387,N_45029,N_45239);
xnor U46388 (N_46388,N_45668,N_45542);
xnor U46389 (N_46389,N_45013,N_45100);
nor U46390 (N_46390,N_45057,N_45566);
nand U46391 (N_46391,N_45701,N_45540);
or U46392 (N_46392,N_45370,N_45155);
nor U46393 (N_46393,N_45272,N_45369);
and U46394 (N_46394,N_45599,N_45999);
nor U46395 (N_46395,N_45467,N_45739);
and U46396 (N_46396,N_45342,N_45353);
nor U46397 (N_46397,N_45477,N_45515);
and U46398 (N_46398,N_45766,N_45818);
nor U46399 (N_46399,N_45150,N_45356);
nand U46400 (N_46400,N_45857,N_45106);
nand U46401 (N_46401,N_45215,N_45700);
or U46402 (N_46402,N_45918,N_45992);
nand U46403 (N_46403,N_45903,N_45468);
or U46404 (N_46404,N_45775,N_45181);
nor U46405 (N_46405,N_45129,N_45777);
xnor U46406 (N_46406,N_45167,N_45352);
nor U46407 (N_46407,N_45407,N_45011);
or U46408 (N_46408,N_45781,N_45768);
nor U46409 (N_46409,N_45078,N_45948);
or U46410 (N_46410,N_45252,N_45449);
or U46411 (N_46411,N_45913,N_45325);
or U46412 (N_46412,N_45438,N_45517);
nor U46413 (N_46413,N_45905,N_45377);
xor U46414 (N_46414,N_45261,N_45240);
or U46415 (N_46415,N_45418,N_45110);
and U46416 (N_46416,N_45830,N_45051);
and U46417 (N_46417,N_45838,N_45380);
nand U46418 (N_46418,N_45505,N_45344);
or U46419 (N_46419,N_45415,N_45977);
or U46420 (N_46420,N_45268,N_45576);
and U46421 (N_46421,N_45444,N_45581);
and U46422 (N_46422,N_45919,N_45393);
nand U46423 (N_46423,N_45976,N_45761);
nor U46424 (N_46424,N_45868,N_45921);
xnor U46425 (N_46425,N_45947,N_45871);
or U46426 (N_46426,N_45388,N_45762);
and U46427 (N_46427,N_45890,N_45586);
nor U46428 (N_46428,N_45974,N_45873);
and U46429 (N_46429,N_45425,N_45141);
xor U46430 (N_46430,N_45791,N_45170);
or U46431 (N_46431,N_45308,N_45471);
nand U46432 (N_46432,N_45879,N_45727);
and U46433 (N_46433,N_45199,N_45006);
xnor U46434 (N_46434,N_45131,N_45846);
nor U46435 (N_46435,N_45844,N_45286);
and U46436 (N_46436,N_45399,N_45191);
xnor U46437 (N_46437,N_45368,N_45386);
and U46438 (N_46438,N_45400,N_45568);
and U46439 (N_46439,N_45772,N_45731);
nand U46440 (N_46440,N_45113,N_45072);
xor U46441 (N_46441,N_45360,N_45487);
nand U46442 (N_46442,N_45856,N_45748);
or U46443 (N_46443,N_45892,N_45911);
nand U46444 (N_46444,N_45065,N_45465);
nand U46445 (N_46445,N_45629,N_45582);
and U46446 (N_46446,N_45001,N_45651);
nor U46447 (N_46447,N_45247,N_45229);
and U46448 (N_46448,N_45295,N_45606);
and U46449 (N_46449,N_45603,N_45210);
or U46450 (N_46450,N_45209,N_45867);
xor U46451 (N_46451,N_45771,N_45022);
or U46452 (N_46452,N_45987,N_45691);
and U46453 (N_46453,N_45019,N_45125);
xor U46454 (N_46454,N_45722,N_45242);
and U46455 (N_46455,N_45881,N_45179);
nand U46456 (N_46456,N_45784,N_45530);
xnor U46457 (N_46457,N_45258,N_45875);
nor U46458 (N_46458,N_45559,N_45894);
nand U46459 (N_46459,N_45214,N_45607);
nand U46460 (N_46460,N_45440,N_45998);
nand U46461 (N_46461,N_45682,N_45284);
xor U46462 (N_46462,N_45669,N_45699);
and U46463 (N_46463,N_45555,N_45623);
xor U46464 (N_46464,N_45138,N_45887);
nand U46465 (N_46465,N_45534,N_45514);
or U46466 (N_46466,N_45248,N_45102);
or U46467 (N_46467,N_45262,N_45650);
nor U46468 (N_46468,N_45865,N_45528);
xnor U46469 (N_46469,N_45986,N_45567);
and U46470 (N_46470,N_45858,N_45486);
nor U46471 (N_46471,N_45133,N_45574);
nand U46472 (N_46472,N_45814,N_45216);
xor U46473 (N_46473,N_45274,N_45663);
nand U46474 (N_46474,N_45713,N_45243);
nor U46475 (N_46475,N_45955,N_45024);
xor U46476 (N_46476,N_45756,N_45038);
nor U46477 (N_46477,N_45952,N_45841);
xor U46478 (N_46478,N_45033,N_45122);
nand U46479 (N_46479,N_45744,N_45068);
nand U46480 (N_46480,N_45805,N_45433);
and U46481 (N_46481,N_45147,N_45973);
nor U46482 (N_46482,N_45462,N_45966);
nand U46483 (N_46483,N_45028,N_45405);
xor U46484 (N_46484,N_45319,N_45536);
xnor U46485 (N_46485,N_45832,N_45256);
nand U46486 (N_46486,N_45593,N_45655);
nand U46487 (N_46487,N_45491,N_45094);
or U46488 (N_46488,N_45949,N_45265);
nor U46489 (N_46489,N_45692,N_45156);
xor U46490 (N_46490,N_45972,N_45560);
or U46491 (N_46491,N_45877,N_45355);
and U46492 (N_46492,N_45221,N_45079);
nand U46493 (N_46493,N_45531,N_45092);
and U46494 (N_46494,N_45680,N_45864);
and U46495 (N_46495,N_45392,N_45631);
nor U46496 (N_46496,N_45608,N_45108);
xnor U46497 (N_46497,N_45403,N_45697);
nand U46498 (N_46498,N_45204,N_45357);
xor U46499 (N_46499,N_45397,N_45450);
or U46500 (N_46500,N_45414,N_45458);
xnor U46501 (N_46501,N_45748,N_45417);
or U46502 (N_46502,N_45893,N_45703);
nor U46503 (N_46503,N_45764,N_45097);
nor U46504 (N_46504,N_45253,N_45028);
nand U46505 (N_46505,N_45141,N_45880);
nand U46506 (N_46506,N_45317,N_45163);
xnor U46507 (N_46507,N_45701,N_45691);
and U46508 (N_46508,N_45959,N_45026);
and U46509 (N_46509,N_45889,N_45853);
xnor U46510 (N_46510,N_45521,N_45898);
xor U46511 (N_46511,N_45350,N_45913);
or U46512 (N_46512,N_45574,N_45324);
nand U46513 (N_46513,N_45669,N_45405);
or U46514 (N_46514,N_45337,N_45939);
and U46515 (N_46515,N_45884,N_45663);
nand U46516 (N_46516,N_45219,N_45498);
nand U46517 (N_46517,N_45181,N_45157);
xor U46518 (N_46518,N_45918,N_45930);
nor U46519 (N_46519,N_45804,N_45448);
and U46520 (N_46520,N_45946,N_45446);
nor U46521 (N_46521,N_45715,N_45176);
xnor U46522 (N_46522,N_45105,N_45361);
nor U46523 (N_46523,N_45259,N_45025);
xnor U46524 (N_46524,N_45720,N_45822);
or U46525 (N_46525,N_45442,N_45224);
or U46526 (N_46526,N_45021,N_45458);
nand U46527 (N_46527,N_45763,N_45132);
and U46528 (N_46528,N_45975,N_45922);
or U46529 (N_46529,N_45282,N_45287);
nand U46530 (N_46530,N_45638,N_45484);
xor U46531 (N_46531,N_45465,N_45849);
nand U46532 (N_46532,N_45234,N_45380);
xnor U46533 (N_46533,N_45768,N_45029);
or U46534 (N_46534,N_45154,N_45214);
xnor U46535 (N_46535,N_45870,N_45267);
or U46536 (N_46536,N_45954,N_45484);
and U46537 (N_46537,N_45861,N_45917);
and U46538 (N_46538,N_45025,N_45658);
or U46539 (N_46539,N_45931,N_45679);
xor U46540 (N_46540,N_45720,N_45159);
nor U46541 (N_46541,N_45322,N_45805);
nand U46542 (N_46542,N_45005,N_45265);
or U46543 (N_46543,N_45341,N_45606);
and U46544 (N_46544,N_45321,N_45451);
nand U46545 (N_46545,N_45791,N_45811);
or U46546 (N_46546,N_45300,N_45303);
xnor U46547 (N_46547,N_45547,N_45981);
nand U46548 (N_46548,N_45177,N_45415);
and U46549 (N_46549,N_45015,N_45581);
or U46550 (N_46550,N_45565,N_45619);
nand U46551 (N_46551,N_45043,N_45929);
and U46552 (N_46552,N_45011,N_45550);
xor U46553 (N_46553,N_45796,N_45509);
xor U46554 (N_46554,N_45864,N_45872);
nand U46555 (N_46555,N_45641,N_45025);
xor U46556 (N_46556,N_45572,N_45013);
nor U46557 (N_46557,N_45133,N_45922);
xnor U46558 (N_46558,N_45448,N_45598);
xnor U46559 (N_46559,N_45155,N_45804);
and U46560 (N_46560,N_45985,N_45583);
or U46561 (N_46561,N_45401,N_45728);
or U46562 (N_46562,N_45302,N_45225);
and U46563 (N_46563,N_45692,N_45430);
or U46564 (N_46564,N_45973,N_45245);
nand U46565 (N_46565,N_45445,N_45497);
xor U46566 (N_46566,N_45708,N_45092);
and U46567 (N_46567,N_45549,N_45044);
and U46568 (N_46568,N_45996,N_45486);
nor U46569 (N_46569,N_45127,N_45225);
nand U46570 (N_46570,N_45430,N_45015);
and U46571 (N_46571,N_45472,N_45436);
and U46572 (N_46572,N_45389,N_45744);
nor U46573 (N_46573,N_45898,N_45378);
and U46574 (N_46574,N_45148,N_45682);
nand U46575 (N_46575,N_45654,N_45259);
xnor U46576 (N_46576,N_45988,N_45770);
nor U46577 (N_46577,N_45039,N_45719);
or U46578 (N_46578,N_45532,N_45731);
nor U46579 (N_46579,N_45001,N_45790);
or U46580 (N_46580,N_45062,N_45671);
nand U46581 (N_46581,N_45017,N_45172);
nor U46582 (N_46582,N_45657,N_45236);
xnor U46583 (N_46583,N_45371,N_45897);
and U46584 (N_46584,N_45170,N_45571);
nor U46585 (N_46585,N_45359,N_45312);
nand U46586 (N_46586,N_45533,N_45025);
or U46587 (N_46587,N_45912,N_45917);
or U46588 (N_46588,N_45392,N_45151);
xnor U46589 (N_46589,N_45839,N_45264);
xnor U46590 (N_46590,N_45499,N_45494);
xor U46591 (N_46591,N_45476,N_45861);
nor U46592 (N_46592,N_45806,N_45258);
or U46593 (N_46593,N_45022,N_45170);
or U46594 (N_46594,N_45472,N_45069);
nor U46595 (N_46595,N_45920,N_45717);
nor U46596 (N_46596,N_45563,N_45185);
nand U46597 (N_46597,N_45869,N_45415);
and U46598 (N_46598,N_45654,N_45752);
xor U46599 (N_46599,N_45821,N_45387);
nor U46600 (N_46600,N_45604,N_45030);
or U46601 (N_46601,N_45124,N_45567);
xor U46602 (N_46602,N_45037,N_45052);
nand U46603 (N_46603,N_45606,N_45544);
nor U46604 (N_46604,N_45447,N_45977);
nand U46605 (N_46605,N_45490,N_45911);
xor U46606 (N_46606,N_45788,N_45938);
nand U46607 (N_46607,N_45488,N_45118);
nand U46608 (N_46608,N_45578,N_45604);
or U46609 (N_46609,N_45939,N_45463);
and U46610 (N_46610,N_45745,N_45746);
nand U46611 (N_46611,N_45949,N_45520);
nand U46612 (N_46612,N_45880,N_45566);
or U46613 (N_46613,N_45818,N_45626);
nor U46614 (N_46614,N_45956,N_45706);
xor U46615 (N_46615,N_45312,N_45252);
and U46616 (N_46616,N_45014,N_45999);
and U46617 (N_46617,N_45950,N_45023);
or U46618 (N_46618,N_45157,N_45943);
nand U46619 (N_46619,N_45278,N_45306);
nand U46620 (N_46620,N_45070,N_45064);
nand U46621 (N_46621,N_45776,N_45745);
or U46622 (N_46622,N_45713,N_45506);
nor U46623 (N_46623,N_45906,N_45633);
xnor U46624 (N_46624,N_45360,N_45580);
nor U46625 (N_46625,N_45091,N_45641);
nand U46626 (N_46626,N_45244,N_45315);
xor U46627 (N_46627,N_45217,N_45811);
or U46628 (N_46628,N_45692,N_45651);
xnor U46629 (N_46629,N_45241,N_45888);
xnor U46630 (N_46630,N_45670,N_45034);
nand U46631 (N_46631,N_45914,N_45905);
and U46632 (N_46632,N_45524,N_45301);
and U46633 (N_46633,N_45370,N_45916);
nor U46634 (N_46634,N_45515,N_45852);
nor U46635 (N_46635,N_45867,N_45679);
and U46636 (N_46636,N_45797,N_45525);
or U46637 (N_46637,N_45781,N_45004);
xor U46638 (N_46638,N_45560,N_45783);
nand U46639 (N_46639,N_45954,N_45996);
and U46640 (N_46640,N_45887,N_45419);
or U46641 (N_46641,N_45079,N_45451);
and U46642 (N_46642,N_45515,N_45849);
nand U46643 (N_46643,N_45141,N_45148);
nand U46644 (N_46644,N_45181,N_45603);
or U46645 (N_46645,N_45469,N_45622);
and U46646 (N_46646,N_45022,N_45070);
nand U46647 (N_46647,N_45106,N_45826);
nand U46648 (N_46648,N_45444,N_45808);
nor U46649 (N_46649,N_45828,N_45296);
nand U46650 (N_46650,N_45262,N_45539);
xor U46651 (N_46651,N_45055,N_45854);
nand U46652 (N_46652,N_45791,N_45486);
nand U46653 (N_46653,N_45875,N_45347);
or U46654 (N_46654,N_45394,N_45140);
nor U46655 (N_46655,N_45437,N_45101);
xnor U46656 (N_46656,N_45925,N_45390);
xnor U46657 (N_46657,N_45256,N_45759);
nand U46658 (N_46658,N_45317,N_45500);
nor U46659 (N_46659,N_45339,N_45816);
or U46660 (N_46660,N_45750,N_45351);
and U46661 (N_46661,N_45555,N_45968);
and U46662 (N_46662,N_45567,N_45053);
xnor U46663 (N_46663,N_45511,N_45156);
nor U46664 (N_46664,N_45284,N_45610);
and U46665 (N_46665,N_45621,N_45322);
nor U46666 (N_46666,N_45070,N_45938);
or U46667 (N_46667,N_45431,N_45350);
or U46668 (N_46668,N_45451,N_45447);
nand U46669 (N_46669,N_45522,N_45811);
and U46670 (N_46670,N_45755,N_45501);
or U46671 (N_46671,N_45851,N_45296);
nand U46672 (N_46672,N_45826,N_45355);
or U46673 (N_46673,N_45140,N_45393);
nand U46674 (N_46674,N_45723,N_45405);
and U46675 (N_46675,N_45354,N_45151);
nand U46676 (N_46676,N_45350,N_45970);
xor U46677 (N_46677,N_45220,N_45396);
nor U46678 (N_46678,N_45766,N_45027);
xor U46679 (N_46679,N_45750,N_45577);
nand U46680 (N_46680,N_45504,N_45484);
and U46681 (N_46681,N_45732,N_45000);
nor U46682 (N_46682,N_45568,N_45416);
nor U46683 (N_46683,N_45986,N_45926);
xnor U46684 (N_46684,N_45978,N_45197);
xnor U46685 (N_46685,N_45298,N_45584);
and U46686 (N_46686,N_45657,N_45967);
nor U46687 (N_46687,N_45373,N_45625);
nor U46688 (N_46688,N_45523,N_45942);
nand U46689 (N_46689,N_45545,N_45540);
nand U46690 (N_46690,N_45260,N_45710);
nand U46691 (N_46691,N_45043,N_45070);
xor U46692 (N_46692,N_45265,N_45856);
and U46693 (N_46693,N_45431,N_45847);
nand U46694 (N_46694,N_45294,N_45118);
xnor U46695 (N_46695,N_45533,N_45770);
and U46696 (N_46696,N_45080,N_45117);
and U46697 (N_46697,N_45924,N_45748);
and U46698 (N_46698,N_45869,N_45323);
and U46699 (N_46699,N_45737,N_45828);
xnor U46700 (N_46700,N_45032,N_45958);
xor U46701 (N_46701,N_45614,N_45257);
nand U46702 (N_46702,N_45550,N_45735);
xor U46703 (N_46703,N_45690,N_45009);
xor U46704 (N_46704,N_45103,N_45290);
nor U46705 (N_46705,N_45203,N_45373);
and U46706 (N_46706,N_45960,N_45053);
xor U46707 (N_46707,N_45712,N_45502);
xor U46708 (N_46708,N_45013,N_45944);
nor U46709 (N_46709,N_45560,N_45058);
xnor U46710 (N_46710,N_45687,N_45326);
xnor U46711 (N_46711,N_45828,N_45092);
nand U46712 (N_46712,N_45707,N_45246);
nand U46713 (N_46713,N_45043,N_45875);
and U46714 (N_46714,N_45061,N_45003);
nand U46715 (N_46715,N_45927,N_45870);
nor U46716 (N_46716,N_45291,N_45504);
nand U46717 (N_46717,N_45044,N_45190);
nand U46718 (N_46718,N_45682,N_45595);
xnor U46719 (N_46719,N_45001,N_45378);
or U46720 (N_46720,N_45461,N_45500);
and U46721 (N_46721,N_45489,N_45828);
or U46722 (N_46722,N_45549,N_45367);
and U46723 (N_46723,N_45022,N_45970);
and U46724 (N_46724,N_45993,N_45533);
nand U46725 (N_46725,N_45132,N_45530);
nor U46726 (N_46726,N_45175,N_45235);
xnor U46727 (N_46727,N_45948,N_45495);
nand U46728 (N_46728,N_45970,N_45868);
nor U46729 (N_46729,N_45437,N_45609);
xnor U46730 (N_46730,N_45934,N_45736);
and U46731 (N_46731,N_45612,N_45096);
nor U46732 (N_46732,N_45378,N_45963);
xor U46733 (N_46733,N_45287,N_45874);
xnor U46734 (N_46734,N_45758,N_45393);
nor U46735 (N_46735,N_45316,N_45014);
nand U46736 (N_46736,N_45832,N_45111);
and U46737 (N_46737,N_45757,N_45940);
xor U46738 (N_46738,N_45176,N_45460);
nand U46739 (N_46739,N_45912,N_45253);
or U46740 (N_46740,N_45228,N_45174);
nor U46741 (N_46741,N_45376,N_45194);
or U46742 (N_46742,N_45629,N_45934);
xor U46743 (N_46743,N_45184,N_45482);
and U46744 (N_46744,N_45475,N_45997);
or U46745 (N_46745,N_45738,N_45026);
or U46746 (N_46746,N_45830,N_45029);
xor U46747 (N_46747,N_45897,N_45615);
nor U46748 (N_46748,N_45358,N_45592);
xnor U46749 (N_46749,N_45623,N_45561);
xor U46750 (N_46750,N_45708,N_45260);
nand U46751 (N_46751,N_45367,N_45035);
nand U46752 (N_46752,N_45046,N_45927);
nand U46753 (N_46753,N_45024,N_45360);
or U46754 (N_46754,N_45621,N_45890);
nor U46755 (N_46755,N_45986,N_45495);
or U46756 (N_46756,N_45802,N_45660);
xnor U46757 (N_46757,N_45480,N_45737);
nand U46758 (N_46758,N_45663,N_45295);
xor U46759 (N_46759,N_45642,N_45175);
and U46760 (N_46760,N_45582,N_45859);
nor U46761 (N_46761,N_45257,N_45493);
nor U46762 (N_46762,N_45970,N_45643);
xor U46763 (N_46763,N_45220,N_45129);
nand U46764 (N_46764,N_45497,N_45074);
nand U46765 (N_46765,N_45023,N_45069);
xnor U46766 (N_46766,N_45071,N_45527);
or U46767 (N_46767,N_45272,N_45841);
or U46768 (N_46768,N_45567,N_45814);
nor U46769 (N_46769,N_45027,N_45790);
nor U46770 (N_46770,N_45721,N_45150);
nand U46771 (N_46771,N_45026,N_45237);
or U46772 (N_46772,N_45385,N_45047);
nand U46773 (N_46773,N_45840,N_45050);
xor U46774 (N_46774,N_45103,N_45819);
and U46775 (N_46775,N_45863,N_45986);
nor U46776 (N_46776,N_45814,N_45528);
xnor U46777 (N_46777,N_45615,N_45969);
nand U46778 (N_46778,N_45300,N_45245);
and U46779 (N_46779,N_45907,N_45363);
xnor U46780 (N_46780,N_45370,N_45807);
nor U46781 (N_46781,N_45948,N_45990);
xnor U46782 (N_46782,N_45978,N_45501);
nand U46783 (N_46783,N_45901,N_45646);
and U46784 (N_46784,N_45158,N_45757);
and U46785 (N_46785,N_45641,N_45209);
nor U46786 (N_46786,N_45864,N_45071);
nor U46787 (N_46787,N_45257,N_45494);
nand U46788 (N_46788,N_45523,N_45474);
and U46789 (N_46789,N_45778,N_45938);
or U46790 (N_46790,N_45237,N_45079);
or U46791 (N_46791,N_45616,N_45277);
and U46792 (N_46792,N_45115,N_45940);
and U46793 (N_46793,N_45712,N_45618);
nor U46794 (N_46794,N_45430,N_45045);
and U46795 (N_46795,N_45954,N_45636);
nand U46796 (N_46796,N_45472,N_45395);
xnor U46797 (N_46797,N_45152,N_45285);
or U46798 (N_46798,N_45923,N_45077);
xor U46799 (N_46799,N_45672,N_45943);
nand U46800 (N_46800,N_45191,N_45786);
xor U46801 (N_46801,N_45058,N_45084);
nor U46802 (N_46802,N_45870,N_45706);
xnor U46803 (N_46803,N_45936,N_45401);
nand U46804 (N_46804,N_45806,N_45570);
or U46805 (N_46805,N_45031,N_45351);
xor U46806 (N_46806,N_45045,N_45791);
nor U46807 (N_46807,N_45875,N_45511);
nand U46808 (N_46808,N_45891,N_45922);
nand U46809 (N_46809,N_45266,N_45050);
or U46810 (N_46810,N_45836,N_45803);
nor U46811 (N_46811,N_45560,N_45676);
nor U46812 (N_46812,N_45002,N_45823);
or U46813 (N_46813,N_45150,N_45423);
nand U46814 (N_46814,N_45029,N_45200);
and U46815 (N_46815,N_45070,N_45298);
nor U46816 (N_46816,N_45959,N_45069);
xor U46817 (N_46817,N_45520,N_45177);
and U46818 (N_46818,N_45267,N_45774);
nor U46819 (N_46819,N_45787,N_45426);
nor U46820 (N_46820,N_45902,N_45952);
nand U46821 (N_46821,N_45191,N_45364);
xnor U46822 (N_46822,N_45452,N_45037);
nand U46823 (N_46823,N_45532,N_45913);
nand U46824 (N_46824,N_45948,N_45119);
and U46825 (N_46825,N_45240,N_45836);
xnor U46826 (N_46826,N_45758,N_45714);
xnor U46827 (N_46827,N_45754,N_45221);
nand U46828 (N_46828,N_45946,N_45336);
xor U46829 (N_46829,N_45479,N_45894);
xnor U46830 (N_46830,N_45266,N_45193);
nor U46831 (N_46831,N_45798,N_45812);
xnor U46832 (N_46832,N_45329,N_45808);
nor U46833 (N_46833,N_45387,N_45673);
or U46834 (N_46834,N_45816,N_45622);
and U46835 (N_46835,N_45191,N_45304);
and U46836 (N_46836,N_45735,N_45484);
nand U46837 (N_46837,N_45854,N_45429);
nand U46838 (N_46838,N_45959,N_45597);
and U46839 (N_46839,N_45140,N_45888);
and U46840 (N_46840,N_45849,N_45114);
nor U46841 (N_46841,N_45792,N_45562);
xnor U46842 (N_46842,N_45848,N_45750);
and U46843 (N_46843,N_45461,N_45091);
xnor U46844 (N_46844,N_45914,N_45145);
nor U46845 (N_46845,N_45566,N_45620);
xnor U46846 (N_46846,N_45254,N_45164);
nor U46847 (N_46847,N_45602,N_45179);
and U46848 (N_46848,N_45788,N_45475);
nor U46849 (N_46849,N_45320,N_45321);
and U46850 (N_46850,N_45330,N_45172);
or U46851 (N_46851,N_45826,N_45905);
and U46852 (N_46852,N_45442,N_45214);
nand U46853 (N_46853,N_45392,N_45334);
nor U46854 (N_46854,N_45346,N_45367);
nand U46855 (N_46855,N_45265,N_45090);
or U46856 (N_46856,N_45755,N_45013);
and U46857 (N_46857,N_45487,N_45112);
or U46858 (N_46858,N_45889,N_45026);
nand U46859 (N_46859,N_45425,N_45752);
and U46860 (N_46860,N_45454,N_45725);
xor U46861 (N_46861,N_45288,N_45462);
or U46862 (N_46862,N_45203,N_45210);
and U46863 (N_46863,N_45790,N_45769);
nor U46864 (N_46864,N_45142,N_45294);
or U46865 (N_46865,N_45883,N_45356);
and U46866 (N_46866,N_45459,N_45702);
and U46867 (N_46867,N_45057,N_45879);
or U46868 (N_46868,N_45759,N_45371);
nor U46869 (N_46869,N_45206,N_45845);
and U46870 (N_46870,N_45128,N_45664);
nand U46871 (N_46871,N_45624,N_45294);
nand U46872 (N_46872,N_45976,N_45798);
and U46873 (N_46873,N_45227,N_45409);
xnor U46874 (N_46874,N_45266,N_45095);
nand U46875 (N_46875,N_45230,N_45420);
xor U46876 (N_46876,N_45824,N_45288);
xnor U46877 (N_46877,N_45388,N_45583);
xor U46878 (N_46878,N_45647,N_45265);
nor U46879 (N_46879,N_45530,N_45277);
nand U46880 (N_46880,N_45829,N_45221);
xor U46881 (N_46881,N_45873,N_45556);
and U46882 (N_46882,N_45461,N_45740);
nor U46883 (N_46883,N_45480,N_45519);
nand U46884 (N_46884,N_45584,N_45557);
nand U46885 (N_46885,N_45706,N_45465);
and U46886 (N_46886,N_45324,N_45177);
and U46887 (N_46887,N_45765,N_45503);
nand U46888 (N_46888,N_45303,N_45741);
nor U46889 (N_46889,N_45941,N_45229);
and U46890 (N_46890,N_45445,N_45653);
nor U46891 (N_46891,N_45946,N_45439);
nand U46892 (N_46892,N_45617,N_45342);
nor U46893 (N_46893,N_45399,N_45562);
nand U46894 (N_46894,N_45981,N_45691);
and U46895 (N_46895,N_45550,N_45677);
and U46896 (N_46896,N_45068,N_45310);
or U46897 (N_46897,N_45740,N_45809);
and U46898 (N_46898,N_45325,N_45544);
or U46899 (N_46899,N_45271,N_45325);
nand U46900 (N_46900,N_45516,N_45050);
nand U46901 (N_46901,N_45894,N_45209);
and U46902 (N_46902,N_45852,N_45428);
xor U46903 (N_46903,N_45832,N_45075);
or U46904 (N_46904,N_45663,N_45929);
or U46905 (N_46905,N_45853,N_45125);
nor U46906 (N_46906,N_45413,N_45023);
or U46907 (N_46907,N_45420,N_45883);
nand U46908 (N_46908,N_45242,N_45024);
or U46909 (N_46909,N_45091,N_45571);
and U46910 (N_46910,N_45172,N_45674);
xnor U46911 (N_46911,N_45942,N_45325);
nor U46912 (N_46912,N_45638,N_45184);
nand U46913 (N_46913,N_45513,N_45336);
or U46914 (N_46914,N_45897,N_45965);
and U46915 (N_46915,N_45191,N_45540);
nand U46916 (N_46916,N_45606,N_45563);
xnor U46917 (N_46917,N_45887,N_45123);
and U46918 (N_46918,N_45852,N_45578);
or U46919 (N_46919,N_45120,N_45836);
and U46920 (N_46920,N_45980,N_45593);
nor U46921 (N_46921,N_45819,N_45438);
xnor U46922 (N_46922,N_45843,N_45502);
xor U46923 (N_46923,N_45458,N_45567);
xor U46924 (N_46924,N_45589,N_45782);
nand U46925 (N_46925,N_45097,N_45571);
or U46926 (N_46926,N_45255,N_45761);
and U46927 (N_46927,N_45431,N_45750);
and U46928 (N_46928,N_45437,N_45148);
and U46929 (N_46929,N_45072,N_45992);
and U46930 (N_46930,N_45653,N_45475);
xnor U46931 (N_46931,N_45619,N_45064);
nand U46932 (N_46932,N_45878,N_45074);
nor U46933 (N_46933,N_45031,N_45940);
or U46934 (N_46934,N_45416,N_45316);
or U46935 (N_46935,N_45086,N_45976);
xor U46936 (N_46936,N_45012,N_45196);
or U46937 (N_46937,N_45848,N_45177);
or U46938 (N_46938,N_45551,N_45504);
nand U46939 (N_46939,N_45381,N_45881);
xnor U46940 (N_46940,N_45627,N_45586);
and U46941 (N_46941,N_45700,N_45327);
nand U46942 (N_46942,N_45399,N_45903);
and U46943 (N_46943,N_45227,N_45607);
nor U46944 (N_46944,N_45108,N_45269);
nor U46945 (N_46945,N_45763,N_45193);
nor U46946 (N_46946,N_45413,N_45198);
and U46947 (N_46947,N_45860,N_45927);
and U46948 (N_46948,N_45333,N_45426);
nand U46949 (N_46949,N_45946,N_45890);
or U46950 (N_46950,N_45073,N_45651);
xnor U46951 (N_46951,N_45697,N_45586);
and U46952 (N_46952,N_45487,N_45719);
and U46953 (N_46953,N_45572,N_45328);
or U46954 (N_46954,N_45827,N_45073);
nor U46955 (N_46955,N_45546,N_45001);
or U46956 (N_46956,N_45590,N_45692);
and U46957 (N_46957,N_45178,N_45889);
or U46958 (N_46958,N_45768,N_45722);
nor U46959 (N_46959,N_45372,N_45689);
xnor U46960 (N_46960,N_45883,N_45305);
nor U46961 (N_46961,N_45518,N_45440);
nor U46962 (N_46962,N_45776,N_45431);
nand U46963 (N_46963,N_45415,N_45787);
and U46964 (N_46964,N_45067,N_45269);
xnor U46965 (N_46965,N_45049,N_45344);
xor U46966 (N_46966,N_45007,N_45201);
and U46967 (N_46967,N_45942,N_45701);
nand U46968 (N_46968,N_45859,N_45694);
nand U46969 (N_46969,N_45671,N_45522);
nor U46970 (N_46970,N_45609,N_45841);
nand U46971 (N_46971,N_45704,N_45184);
nand U46972 (N_46972,N_45187,N_45649);
xnor U46973 (N_46973,N_45299,N_45746);
xor U46974 (N_46974,N_45384,N_45814);
nor U46975 (N_46975,N_45010,N_45989);
and U46976 (N_46976,N_45899,N_45216);
nand U46977 (N_46977,N_45956,N_45034);
or U46978 (N_46978,N_45097,N_45066);
or U46979 (N_46979,N_45085,N_45563);
and U46980 (N_46980,N_45870,N_45579);
and U46981 (N_46981,N_45919,N_45332);
nand U46982 (N_46982,N_45900,N_45234);
nor U46983 (N_46983,N_45025,N_45578);
nor U46984 (N_46984,N_45400,N_45705);
nor U46985 (N_46985,N_45028,N_45006);
nand U46986 (N_46986,N_45450,N_45027);
nand U46987 (N_46987,N_45945,N_45585);
or U46988 (N_46988,N_45239,N_45258);
nor U46989 (N_46989,N_45094,N_45164);
and U46990 (N_46990,N_45941,N_45265);
and U46991 (N_46991,N_45162,N_45526);
and U46992 (N_46992,N_45407,N_45040);
xnor U46993 (N_46993,N_45185,N_45289);
xnor U46994 (N_46994,N_45809,N_45393);
xor U46995 (N_46995,N_45146,N_45178);
nand U46996 (N_46996,N_45941,N_45683);
nor U46997 (N_46997,N_45095,N_45118);
or U46998 (N_46998,N_45437,N_45084);
and U46999 (N_46999,N_45130,N_45527);
xor U47000 (N_47000,N_46127,N_46037);
and U47001 (N_47001,N_46909,N_46378);
xnor U47002 (N_47002,N_46282,N_46947);
nor U47003 (N_47003,N_46849,N_46192);
xor U47004 (N_47004,N_46358,N_46995);
and U47005 (N_47005,N_46013,N_46865);
and U47006 (N_47006,N_46341,N_46689);
xor U47007 (N_47007,N_46837,N_46871);
xor U47008 (N_47008,N_46915,N_46548);
or U47009 (N_47009,N_46510,N_46039);
nor U47010 (N_47010,N_46890,N_46092);
nand U47011 (N_47011,N_46447,N_46119);
or U47012 (N_47012,N_46681,N_46607);
nand U47013 (N_47013,N_46894,N_46258);
nand U47014 (N_47014,N_46186,N_46695);
nand U47015 (N_47015,N_46091,N_46961);
nor U47016 (N_47016,N_46716,N_46924);
nor U47017 (N_47017,N_46266,N_46189);
nand U47018 (N_47018,N_46723,N_46169);
and U47019 (N_47019,N_46280,N_46868);
or U47020 (N_47020,N_46130,N_46353);
nand U47021 (N_47021,N_46674,N_46409);
xor U47022 (N_47022,N_46416,N_46797);
nand U47023 (N_47023,N_46066,N_46468);
nand U47024 (N_47024,N_46914,N_46584);
or U47025 (N_47025,N_46106,N_46232);
nand U47026 (N_47026,N_46509,N_46854);
xor U47027 (N_47027,N_46090,N_46290);
nor U47028 (N_47028,N_46940,N_46496);
nor U47029 (N_47029,N_46658,N_46850);
nand U47030 (N_47030,N_46948,N_46593);
nor U47031 (N_47031,N_46929,N_46205);
nand U47032 (N_47032,N_46034,N_46029);
nor U47033 (N_47033,N_46454,N_46880);
and U47034 (N_47034,N_46970,N_46113);
or U47035 (N_47035,N_46283,N_46394);
nand U47036 (N_47036,N_46807,N_46698);
nor U47037 (N_47037,N_46105,N_46984);
xor U47038 (N_47038,N_46620,N_46009);
xnor U47039 (N_47039,N_46370,N_46041);
nor U47040 (N_47040,N_46663,N_46457);
or U47041 (N_47041,N_46456,N_46706);
nor U47042 (N_47042,N_46533,N_46863);
nor U47043 (N_47043,N_46323,N_46964);
xor U47044 (N_47044,N_46212,N_46730);
nand U47045 (N_47045,N_46249,N_46881);
and U47046 (N_47046,N_46740,N_46616);
and U47047 (N_47047,N_46306,N_46256);
and U47048 (N_47048,N_46081,N_46200);
xnor U47049 (N_47049,N_46839,N_46634);
xnor U47050 (N_47050,N_46460,N_46823);
nor U47051 (N_47051,N_46263,N_46506);
and U47052 (N_47052,N_46810,N_46361);
or U47053 (N_47053,N_46571,N_46419);
nand U47054 (N_47054,N_46683,N_46500);
xor U47055 (N_47055,N_46042,N_46324);
and U47056 (N_47056,N_46618,N_46343);
xor U47057 (N_47057,N_46809,N_46694);
nor U47058 (N_47058,N_46910,N_46063);
and U47059 (N_47059,N_46768,N_46462);
or U47060 (N_47060,N_46545,N_46110);
and U47061 (N_47061,N_46675,N_46216);
or U47062 (N_47062,N_46491,N_46828);
nor U47063 (N_47063,N_46832,N_46313);
or U47064 (N_47064,N_46356,N_46421);
or U47065 (N_47065,N_46523,N_46776);
and U47066 (N_47066,N_46733,N_46629);
nor U47067 (N_47067,N_46762,N_46685);
or U47068 (N_47068,N_46008,N_46573);
nand U47069 (N_47069,N_46722,N_46067);
nor U47070 (N_47070,N_46404,N_46236);
and U47071 (N_47071,N_46728,N_46588);
nand U47072 (N_47072,N_46682,N_46650);
nor U47073 (N_47073,N_46911,N_46741);
nor U47074 (N_47074,N_46161,N_46412);
and U47075 (N_47075,N_46662,N_46250);
or U47076 (N_47076,N_46707,N_46426);
nor U47077 (N_47077,N_46575,N_46815);
and U47078 (N_47078,N_46763,N_46905);
nor U47079 (N_47079,N_46992,N_46112);
nand U47080 (N_47080,N_46570,N_46145);
nor U47081 (N_47081,N_46614,N_46641);
or U47082 (N_47082,N_46483,N_46163);
nand U47083 (N_47083,N_46852,N_46131);
and U47084 (N_47084,N_46949,N_46279);
nor U47085 (N_47085,N_46184,N_46851);
nor U47086 (N_47086,N_46516,N_46596);
or U47087 (N_47087,N_46595,N_46269);
or U47088 (N_47088,N_46450,N_46676);
or U47089 (N_47089,N_46494,N_46308);
nor U47090 (N_47090,N_46811,N_46726);
nor U47091 (N_47091,N_46490,N_46417);
or U47092 (N_47092,N_46051,N_46338);
xor U47093 (N_47093,N_46739,N_46679);
and U47094 (N_47094,N_46374,N_46011);
nor U47095 (N_47095,N_46297,N_46284);
xor U47096 (N_47096,N_46512,N_46959);
nor U47097 (N_47097,N_46774,N_46070);
and U47098 (N_47098,N_46691,N_46368);
xnor U47099 (N_47099,N_46633,N_46291);
and U47100 (N_47100,N_46973,N_46165);
or U47101 (N_47101,N_46055,N_46415);
or U47102 (N_47102,N_46845,N_46923);
and U47103 (N_47103,N_46143,N_46793);
and U47104 (N_47104,N_46974,N_46922);
and U47105 (N_47105,N_46759,N_46157);
nand U47106 (N_47106,N_46170,N_46213);
and U47107 (N_47107,N_46073,N_46962);
and U47108 (N_47108,N_46887,N_46862);
nand U47109 (N_47109,N_46628,N_46968);
nor U47110 (N_47110,N_46791,N_46393);
xor U47111 (N_47111,N_46238,N_46798);
or U47112 (N_47112,N_46861,N_46919);
and U47113 (N_47113,N_46336,N_46502);
nand U47114 (N_47114,N_46151,N_46064);
nor U47115 (N_47115,N_46321,N_46757);
and U47116 (N_47116,N_46908,N_46729);
xnor U47117 (N_47117,N_46830,N_46557);
nand U47118 (N_47118,N_46060,N_46826);
nor U47119 (N_47119,N_46111,N_46414);
xnor U47120 (N_47120,N_46221,N_46373);
xor U47121 (N_47121,N_46167,N_46482);
nand U47122 (N_47122,N_46268,N_46162);
and U47123 (N_47123,N_46299,N_46337);
nand U47124 (N_47124,N_46149,N_46672);
or U47125 (N_47125,N_46814,N_46437);
nor U47126 (N_47126,N_46044,N_46960);
or U47127 (N_47127,N_46208,N_46334);
nor U47128 (N_47128,N_46972,N_46779);
nand U47129 (N_47129,N_46943,N_46230);
nor U47130 (N_47130,N_46549,N_46996);
nand U47131 (N_47131,N_46859,N_46101);
nor U47132 (N_47132,N_46538,N_46524);
or U47133 (N_47133,N_46198,N_46848);
or U47134 (N_47134,N_46649,N_46591);
or U47135 (N_47135,N_46876,N_46339);
xor U47136 (N_47136,N_46952,N_46276);
nand U47137 (N_47137,N_46532,N_46428);
or U47138 (N_47138,N_46001,N_46470);
and U47139 (N_47139,N_46272,N_46875);
or U47140 (N_47140,N_46692,N_46701);
nand U47141 (N_47141,N_46069,N_46436);
xor U47142 (N_47142,N_46802,N_46185);
nor U47143 (N_47143,N_46085,N_46438);
nand U47144 (N_47144,N_46176,N_46277);
nor U47145 (N_47145,N_46049,N_46800);
or U47146 (N_47146,N_46246,N_46357);
nand U47147 (N_47147,N_46079,N_46093);
and U47148 (N_47148,N_46035,N_46535);
or U47149 (N_47149,N_46777,N_46829);
or U47150 (N_47150,N_46138,N_46316);
nor U47151 (N_47151,N_46076,N_46869);
nand U47152 (N_47152,N_46242,N_46062);
nor U47153 (N_47153,N_46918,N_46362);
nand U47154 (N_47154,N_46825,N_46420);
or U47155 (N_47155,N_46660,N_46801);
nor U47156 (N_47156,N_46898,N_46521);
xnor U47157 (N_47157,N_46214,N_46015);
nor U47158 (N_47158,N_46147,N_46432);
xor U47159 (N_47159,N_46177,N_46738);
nand U47160 (N_47160,N_46096,N_46963);
or U47161 (N_47161,N_46465,N_46006);
nand U47162 (N_47162,N_46030,N_46844);
nand U47163 (N_47163,N_46673,N_46471);
or U47164 (N_47164,N_46585,N_46582);
xor U47165 (N_47165,N_46813,N_46322);
and U47166 (N_47166,N_46708,N_46155);
xor U47167 (N_47167,N_46325,N_46354);
and U47168 (N_47168,N_46900,N_46474);
xnor U47169 (N_47169,N_46193,N_46109);
nor U47170 (N_47170,N_46997,N_46160);
or U47171 (N_47171,N_46648,N_46550);
nand U47172 (N_47172,N_46957,N_46427);
nor U47173 (N_47173,N_46363,N_46466);
and U47174 (N_47174,N_46921,N_46690);
nor U47175 (N_47175,N_46100,N_46259);
xnor U47176 (N_47176,N_46142,N_46241);
nand U47177 (N_47177,N_46889,N_46439);
nand U47178 (N_47178,N_46985,N_46603);
nand U47179 (N_47179,N_46396,N_46913);
nor U47180 (N_47180,N_46937,N_46377);
xor U47181 (N_47181,N_46054,N_46770);
nand U47182 (N_47182,N_46040,N_46950);
nor U47183 (N_47183,N_46072,N_46315);
and U47184 (N_47184,N_46194,N_46756);
nand U47185 (N_47185,N_46441,N_46806);
xnor U47186 (N_47186,N_46772,N_46651);
nand U47187 (N_47187,N_46349,N_46712);
or U47188 (N_47188,N_46834,N_46243);
nand U47189 (N_47189,N_46265,N_46418);
and U47190 (N_47190,N_46342,N_46817);
or U47191 (N_47191,N_46075,N_46017);
or U47192 (N_47192,N_46696,N_46047);
nor U47193 (N_47193,N_46643,N_46355);
and U47194 (N_47194,N_46812,N_46877);
xnor U47195 (N_47195,N_46391,N_46872);
and U47196 (N_47196,N_46540,N_46032);
nand U47197 (N_47197,N_46024,N_46107);
nor U47198 (N_47198,N_46711,N_46347);
nor U47199 (N_47199,N_46389,N_46804);
and U47200 (N_47200,N_46411,N_46498);
and U47201 (N_47201,N_46139,N_46977);
nor U47202 (N_47202,N_46794,N_46993);
xor U47203 (N_47203,N_46764,N_46710);
nor U47204 (N_47204,N_46602,N_46517);
xor U47205 (N_47205,N_46400,N_46114);
xnor U47206 (N_47206,N_46704,N_46352);
nor U47207 (N_47207,N_46320,N_46188);
or U47208 (N_47208,N_46061,N_46182);
and U47209 (N_47209,N_46560,N_46318);
nand U47210 (N_47210,N_46951,N_46164);
and U47211 (N_47211,N_46159,N_46892);
nor U47212 (N_47212,N_46860,N_46749);
nor U47213 (N_47213,N_46522,N_46744);
and U47214 (N_47214,N_46492,N_46223);
nand U47215 (N_47215,N_46592,N_46452);
xor U47216 (N_47216,N_46309,N_46270);
nand U47217 (N_47217,N_46327,N_46481);
nor U47218 (N_47218,N_46218,N_46990);
xnor U47219 (N_47219,N_46172,N_46754);
nor U47220 (N_47220,N_46399,N_46551);
nand U47221 (N_47221,N_46350,N_46191);
nand U47222 (N_47222,N_46818,N_46088);
and U47223 (N_47223,N_46286,N_46330);
or U47224 (N_47224,N_46897,N_46906);
nand U47225 (N_47225,N_46788,N_46783);
nor U47226 (N_47226,N_46244,N_46307);
nor U47227 (N_47227,N_46767,N_46464);
and U47228 (N_47228,N_46442,N_46511);
nor U47229 (N_47229,N_46004,N_46262);
xor U47230 (N_47230,N_46916,N_46359);
nand U47231 (N_47231,N_46513,N_46099);
nor U47232 (N_47232,N_46397,N_46632);
nor U47233 (N_47233,N_46742,N_46917);
or U47234 (N_47234,N_46469,N_46448);
and U47235 (N_47235,N_46821,N_46463);
xor U47236 (N_47236,N_46458,N_46273);
or U47237 (N_47237,N_46120,N_46606);
xnor U47238 (N_47238,N_46989,N_46669);
nand U47239 (N_47239,N_46022,N_46805);
and U47240 (N_47240,N_46048,N_46007);
xnor U47241 (N_47241,N_46652,N_46202);
xor U47242 (N_47242,N_46670,N_46928);
nor U47243 (N_47243,N_46058,N_46253);
nand U47244 (N_47244,N_46976,N_46478);
xor U47245 (N_47245,N_46116,N_46944);
nor U47246 (N_47246,N_46598,N_46537);
nor U47247 (N_47247,N_46904,N_46773);
nor U47248 (N_47248,N_46688,N_46424);
xor U47249 (N_47249,N_46687,N_46056);
nor U47250 (N_47250,N_46727,N_46750);
or U47251 (N_47251,N_46587,N_46667);
or U47252 (N_47252,N_46925,N_46453);
or U47253 (N_47253,N_46736,N_46899);
or U47254 (N_47254,N_46385,N_46274);
and U47255 (N_47255,N_46755,N_46140);
nand U47256 (N_47256,N_46835,N_46623);
and U47257 (N_47257,N_46576,N_46636);
xor U47258 (N_47258,N_46901,N_46975);
xor U47259 (N_47259,N_46311,N_46095);
and U47260 (N_47260,N_46920,N_46581);
or U47261 (N_47261,N_46534,N_46847);
nand U47262 (N_47262,N_46033,N_46748);
or U47263 (N_47263,N_46827,N_46611);
xnor U47264 (N_47264,N_46045,N_46833);
xor U47265 (N_47265,N_46732,N_46668);
nor U47266 (N_47266,N_46375,N_46195);
nor U47267 (N_47267,N_46831,N_46528);
nand U47268 (N_47268,N_46068,N_46403);
xor U47269 (N_47269,N_46994,N_46945);
or U47270 (N_47270,N_46933,N_46751);
xor U47271 (N_47271,N_46697,N_46637);
nor U47272 (N_47272,N_46659,N_46335);
or U47273 (N_47273,N_46747,N_46154);
or U47274 (N_47274,N_46087,N_46803);
nor U47275 (N_47275,N_46329,N_46175);
xnor U47276 (N_47276,N_46539,N_46724);
nor U47277 (N_47277,N_46866,N_46518);
nor U47278 (N_47278,N_46954,N_46501);
or U47279 (N_47279,N_46792,N_46050);
nand U47280 (N_47280,N_46519,N_46129);
and U47281 (N_47281,N_46879,N_46955);
or U47282 (N_47282,N_46365,N_46612);
and U47283 (N_47283,N_46884,N_46302);
or U47284 (N_47284,N_46656,N_46211);
or U47285 (N_47285,N_46778,N_46179);
or U47286 (N_47286,N_46010,N_46664);
nor U47287 (N_47287,N_46134,N_46326);
nand U47288 (N_47288,N_46445,N_46126);
nand U47289 (N_47289,N_46558,N_46398);
xnor U47290 (N_47290,N_46562,N_46758);
nand U47291 (N_47291,N_46719,N_46544);
and U47292 (N_47292,N_46451,N_46247);
nor U47293 (N_47293,N_46215,N_46018);
or U47294 (N_47294,N_46122,N_46261);
or U47295 (N_47295,N_46619,N_46016);
and U47296 (N_47296,N_46407,N_46383);
and U47297 (N_47297,N_46796,N_46264);
and U47298 (N_47298,N_46666,N_46245);
or U47299 (N_47299,N_46608,N_46965);
xnor U47300 (N_47300,N_46178,N_46405);
nand U47301 (N_47301,N_46577,N_46461);
and U47302 (N_47302,N_46431,N_46146);
xor U47303 (N_47303,N_46183,N_46328);
and U47304 (N_47304,N_46382,N_46480);
nand U47305 (N_47305,N_46319,N_46477);
nand U47306 (N_47306,N_46966,N_46639);
and U47307 (N_47307,N_46433,N_46625);
or U47308 (N_47308,N_46507,N_46304);
nor U47309 (N_47309,N_46765,N_46609);
or U47310 (N_47310,N_46379,N_46434);
xnor U47311 (N_47311,N_46021,N_46564);
nor U47312 (N_47312,N_46234,N_46958);
nand U47313 (N_47313,N_46305,N_46893);
xor U47314 (N_47314,N_46784,N_46731);
xor U47315 (N_47315,N_46144,N_46148);
or U47316 (N_47316,N_46569,N_46333);
nand U47317 (N_47317,N_46487,N_46734);
xnor U47318 (N_47318,N_46671,N_46858);
or U47319 (N_47319,N_46401,N_46753);
or U47320 (N_47320,N_46345,N_46028);
nand U47321 (N_47321,N_46310,N_46621);
and U47322 (N_47322,N_46019,N_46402);
nand U47323 (N_47323,N_46873,N_46430);
and U47324 (N_47324,N_46074,N_46484);
nor U47325 (N_47325,N_46372,N_46158);
and U47326 (N_47326,N_46298,N_46429);
nor U47327 (N_47327,N_46766,N_46714);
nor U47328 (N_47328,N_46240,N_46941);
xor U47329 (N_47329,N_46289,N_46455);
nor U47330 (N_47330,N_46390,N_46786);
nor U47331 (N_47331,N_46166,N_46281);
nand U47332 (N_47332,N_46853,N_46002);
or U47333 (N_47333,N_46499,N_46233);
and U47334 (N_47334,N_46980,N_46610);
nand U47335 (N_47335,N_46317,N_46220);
nand U47336 (N_47336,N_46926,N_46423);
and U47337 (N_47337,N_46953,N_46536);
nand U47338 (N_47338,N_46824,N_46991);
xor U47339 (N_47339,N_46857,N_46855);
nand U47340 (N_47340,N_46082,N_46312);
nor U47341 (N_47341,N_46137,N_46257);
and U47342 (N_47342,N_46787,N_46475);
nand U47343 (N_47343,N_46979,N_46617);
or U47344 (N_47344,N_46935,N_46206);
and U47345 (N_47345,N_46364,N_46392);
nand U47346 (N_47346,N_46999,N_46229);
and U47347 (N_47347,N_46907,N_46235);
xnor U47348 (N_47348,N_46117,N_46295);
or U47349 (N_47349,N_46680,N_46841);
and U47350 (N_47350,N_46231,N_46563);
or U47351 (N_47351,N_46485,N_46574);
and U47352 (N_47352,N_46566,N_46572);
nand U47353 (N_47353,N_46878,N_46026);
xor U47354 (N_47354,N_46971,N_46084);
xnor U47355 (N_47355,N_46267,N_46473);
xor U47356 (N_47356,N_46296,N_46406);
or U47357 (N_47357,N_46381,N_46956);
nand U47358 (N_47358,N_46912,N_46579);
nand U47359 (N_47359,N_46882,N_46775);
and U47360 (N_47360,N_46156,N_46555);
and U47361 (N_47361,N_46780,N_46699);
xor U47362 (N_47362,N_46553,N_46344);
and U47363 (N_47363,N_46526,N_46987);
and U47364 (N_47364,N_46440,N_46981);
nand U47365 (N_47365,N_46624,N_46816);
and U47366 (N_47366,N_46896,N_46104);
nor U47367 (N_47367,N_46644,N_46867);
xor U47368 (N_47368,N_46586,N_46038);
xor U47369 (N_47369,N_46790,N_46713);
xor U47370 (N_47370,N_46781,N_46927);
or U47371 (N_47371,N_46180,N_46479);
nand U47372 (N_47372,N_46376,N_46559);
and U47373 (N_47373,N_46053,N_46799);
nand U47374 (N_47374,N_46367,N_46525);
and U47375 (N_47375,N_46278,N_46141);
xor U47376 (N_47376,N_46599,N_46505);
or U47377 (N_47377,N_46174,N_46410);
or U47378 (N_47378,N_46546,N_46969);
or U47379 (N_47379,N_46888,N_46745);
and U47380 (N_47380,N_46702,N_46023);
xnor U47381 (N_47381,N_46568,N_46700);
and U47382 (N_47382,N_46102,N_46446);
nor U47383 (N_47383,N_46503,N_46275);
nand U47384 (N_47384,N_46657,N_46870);
and U47385 (N_47385,N_46046,N_46902);
xor U47386 (N_47386,N_46089,N_46635);
nor U47387 (N_47387,N_46005,N_46171);
xnor U47388 (N_47388,N_46360,N_46108);
nor U47389 (N_47389,N_46565,N_46583);
and U47390 (N_47390,N_46604,N_46486);
or U47391 (N_47391,N_46613,N_46939);
xnor U47392 (N_47392,N_46721,N_46371);
or U47393 (N_47393,N_46493,N_46590);
nor U47394 (N_47394,N_46210,N_46718);
nor U47395 (N_47395,N_46459,N_46932);
xnor U47396 (N_47396,N_46025,N_46287);
nand U47397 (N_47397,N_46541,N_46514);
or U47398 (N_47398,N_46133,N_46136);
xnor U47399 (N_47399,N_46207,N_46883);
nor U47400 (N_47400,N_46098,N_46886);
and U47401 (N_47401,N_46653,N_46237);
or U47402 (N_47402,N_46065,N_46665);
and U47403 (N_47403,N_46225,N_46654);
nor U47404 (N_47404,N_46217,N_46168);
nor U47405 (N_47405,N_46661,N_46201);
xor U47406 (N_47406,N_46934,N_46292);
or U47407 (N_47407,N_46626,N_46543);
nor U47408 (N_47408,N_46083,N_46260);
xnor U47409 (N_47409,N_46578,N_46303);
or U47410 (N_47410,N_46071,N_46150);
and U47411 (N_47411,N_46589,N_46931);
xor U47412 (N_47412,N_46597,N_46000);
xnor U47413 (N_47413,N_46746,N_46020);
nand U47414 (N_47414,N_46838,N_46331);
xnor U47415 (N_47415,N_46228,N_46594);
nand U47416 (N_47416,N_46715,N_46388);
xor U47417 (N_47417,N_46580,N_46631);
or U47418 (N_47418,N_46622,N_46895);
nor U47419 (N_47419,N_46836,N_46467);
nand U47420 (N_47420,N_46314,N_46422);
nor U47421 (N_47421,N_46226,N_46530);
and U47422 (N_47422,N_46782,N_46735);
and U47423 (N_47423,N_46605,N_46080);
nor U47424 (N_47424,N_46251,N_46743);
nor U47425 (N_47425,N_46301,N_46097);
xor U47426 (N_47426,N_46982,N_46248);
and U47427 (N_47427,N_46647,N_46115);
xnor U47428 (N_47428,N_46840,N_46488);
nor U47429 (N_47429,N_46425,N_46332);
nor U47430 (N_47430,N_46556,N_46197);
or U47431 (N_47431,N_46627,N_46891);
or U47432 (N_47432,N_46489,N_46630);
or U47433 (N_47433,N_46737,N_46036);
and U47434 (N_47434,N_46472,N_46938);
xor U47435 (N_47435,N_46476,N_46057);
or U47436 (N_47436,N_46703,N_46254);
nor U47437 (N_47437,N_46808,N_46785);
nor U47438 (N_47438,N_46520,N_46642);
and U47439 (N_47439,N_46340,N_46795);
and U47440 (N_47440,N_46094,N_46942);
nand U47441 (N_47441,N_46395,N_46190);
nor U47442 (N_47442,N_46567,N_46132);
nand U47443 (N_47443,N_46531,N_46408);
xnor U47444 (N_47444,N_46181,N_46936);
and U47445 (N_47445,N_46078,N_46027);
and U47446 (N_47446,N_46387,N_46227);
and U47447 (N_47447,N_46600,N_46615);
or U47448 (N_47448,N_46123,N_46843);
or U47449 (N_47449,N_46125,N_46118);
nand U47450 (N_47450,N_46173,N_46789);
and U47451 (N_47451,N_46252,N_46542);
nor U47452 (N_47452,N_46293,N_46384);
xor U47453 (N_47453,N_46444,N_46271);
nand U47454 (N_47454,N_46413,N_46885);
nor U47455 (N_47455,N_46443,N_46820);
nand U47456 (N_47456,N_46135,N_46705);
or U47457 (N_47457,N_46822,N_46012);
and U47458 (N_47458,N_46638,N_46645);
nand U47459 (N_47459,N_46846,N_46504);
and U47460 (N_47460,N_46864,N_46196);
nor U47461 (N_47461,N_46300,N_46014);
and U47462 (N_47462,N_46222,N_46720);
nand U47463 (N_47463,N_46003,N_46380);
nand U47464 (N_47464,N_46449,N_46219);
nor U47465 (N_47465,N_46204,N_46086);
nand U47466 (N_47466,N_46761,N_46752);
nand U47467 (N_47467,N_46967,N_46819);
nand U47468 (N_47468,N_46239,N_46121);
and U47469 (N_47469,N_46209,N_46874);
and U47470 (N_47470,N_46527,N_46495);
nand U47471 (N_47471,N_46348,N_46043);
nand U47472 (N_47472,N_46152,N_46717);
nand U47473 (N_47473,N_46077,N_46124);
xor U47474 (N_47474,N_46255,N_46725);
or U47475 (N_47475,N_46760,N_46986);
xor U47476 (N_47476,N_46856,N_46369);
xnor U47477 (N_47477,N_46294,N_46978);
nand U47478 (N_47478,N_46128,N_46655);
xnor U47479 (N_47479,N_46386,N_46351);
or U47480 (N_47480,N_46684,N_46946);
xnor U47481 (N_47481,N_46103,N_46677);
and U47482 (N_47482,N_46769,N_46285);
nor U47483 (N_47483,N_46435,N_46497);
nor U47484 (N_47484,N_46515,N_46224);
and U47485 (N_47485,N_46366,N_46988);
nand U47486 (N_47486,N_46554,N_46059);
or U47487 (N_47487,N_46693,N_46601);
nor U47488 (N_47488,N_46346,N_46529);
and U47489 (N_47489,N_46842,N_46199);
nor U47490 (N_47490,N_46187,N_46983);
nand U47491 (N_47491,N_46646,N_46678);
nor U47492 (N_47492,N_46552,N_46903);
and U47493 (N_47493,N_46709,N_46508);
xnor U47494 (N_47494,N_46561,N_46153);
or U47495 (N_47495,N_46771,N_46203);
nor U47496 (N_47496,N_46052,N_46031);
xnor U47497 (N_47497,N_46930,N_46288);
xnor U47498 (N_47498,N_46998,N_46640);
nor U47499 (N_47499,N_46686,N_46547);
and U47500 (N_47500,N_46038,N_46234);
or U47501 (N_47501,N_46342,N_46483);
xnor U47502 (N_47502,N_46588,N_46938);
and U47503 (N_47503,N_46246,N_46700);
and U47504 (N_47504,N_46668,N_46956);
xnor U47505 (N_47505,N_46727,N_46638);
and U47506 (N_47506,N_46989,N_46007);
or U47507 (N_47507,N_46574,N_46390);
xor U47508 (N_47508,N_46344,N_46908);
and U47509 (N_47509,N_46031,N_46330);
or U47510 (N_47510,N_46327,N_46602);
and U47511 (N_47511,N_46987,N_46444);
or U47512 (N_47512,N_46809,N_46441);
xnor U47513 (N_47513,N_46940,N_46734);
or U47514 (N_47514,N_46845,N_46045);
nor U47515 (N_47515,N_46539,N_46978);
or U47516 (N_47516,N_46403,N_46112);
xnor U47517 (N_47517,N_46435,N_46329);
nor U47518 (N_47518,N_46743,N_46581);
or U47519 (N_47519,N_46790,N_46600);
or U47520 (N_47520,N_46175,N_46472);
or U47521 (N_47521,N_46389,N_46543);
and U47522 (N_47522,N_46121,N_46959);
nand U47523 (N_47523,N_46874,N_46049);
nand U47524 (N_47524,N_46638,N_46364);
nand U47525 (N_47525,N_46132,N_46595);
nor U47526 (N_47526,N_46060,N_46886);
nand U47527 (N_47527,N_46320,N_46294);
nand U47528 (N_47528,N_46830,N_46428);
nand U47529 (N_47529,N_46586,N_46058);
nand U47530 (N_47530,N_46168,N_46190);
nor U47531 (N_47531,N_46214,N_46862);
xor U47532 (N_47532,N_46198,N_46698);
and U47533 (N_47533,N_46494,N_46014);
or U47534 (N_47534,N_46915,N_46308);
nor U47535 (N_47535,N_46812,N_46714);
and U47536 (N_47536,N_46983,N_46545);
nor U47537 (N_47537,N_46284,N_46761);
nor U47538 (N_47538,N_46990,N_46807);
or U47539 (N_47539,N_46790,N_46983);
nor U47540 (N_47540,N_46642,N_46933);
or U47541 (N_47541,N_46103,N_46230);
or U47542 (N_47542,N_46841,N_46562);
and U47543 (N_47543,N_46867,N_46061);
nor U47544 (N_47544,N_46540,N_46461);
xnor U47545 (N_47545,N_46025,N_46662);
xnor U47546 (N_47546,N_46113,N_46218);
nand U47547 (N_47547,N_46967,N_46546);
nor U47548 (N_47548,N_46292,N_46027);
nor U47549 (N_47549,N_46165,N_46220);
nand U47550 (N_47550,N_46693,N_46169);
and U47551 (N_47551,N_46611,N_46431);
or U47552 (N_47552,N_46160,N_46318);
xor U47553 (N_47553,N_46265,N_46676);
nand U47554 (N_47554,N_46513,N_46880);
xor U47555 (N_47555,N_46518,N_46043);
xnor U47556 (N_47556,N_46810,N_46834);
nor U47557 (N_47557,N_46631,N_46461);
nand U47558 (N_47558,N_46347,N_46909);
nor U47559 (N_47559,N_46146,N_46360);
xnor U47560 (N_47560,N_46911,N_46567);
or U47561 (N_47561,N_46082,N_46525);
nand U47562 (N_47562,N_46991,N_46590);
or U47563 (N_47563,N_46209,N_46936);
nor U47564 (N_47564,N_46757,N_46605);
and U47565 (N_47565,N_46723,N_46294);
xnor U47566 (N_47566,N_46988,N_46368);
and U47567 (N_47567,N_46125,N_46515);
nand U47568 (N_47568,N_46288,N_46299);
and U47569 (N_47569,N_46144,N_46455);
and U47570 (N_47570,N_46690,N_46548);
nand U47571 (N_47571,N_46034,N_46706);
nand U47572 (N_47572,N_46392,N_46445);
and U47573 (N_47573,N_46450,N_46551);
nor U47574 (N_47574,N_46325,N_46496);
xnor U47575 (N_47575,N_46589,N_46111);
or U47576 (N_47576,N_46524,N_46743);
nor U47577 (N_47577,N_46062,N_46517);
and U47578 (N_47578,N_46155,N_46136);
nor U47579 (N_47579,N_46810,N_46454);
or U47580 (N_47580,N_46498,N_46977);
xnor U47581 (N_47581,N_46082,N_46239);
nor U47582 (N_47582,N_46174,N_46635);
nor U47583 (N_47583,N_46604,N_46450);
or U47584 (N_47584,N_46562,N_46512);
nor U47585 (N_47585,N_46647,N_46744);
or U47586 (N_47586,N_46882,N_46069);
xnor U47587 (N_47587,N_46342,N_46946);
xor U47588 (N_47588,N_46082,N_46090);
xnor U47589 (N_47589,N_46203,N_46416);
and U47590 (N_47590,N_46280,N_46962);
nor U47591 (N_47591,N_46554,N_46402);
nand U47592 (N_47592,N_46141,N_46938);
and U47593 (N_47593,N_46556,N_46851);
nand U47594 (N_47594,N_46391,N_46845);
xor U47595 (N_47595,N_46160,N_46002);
nand U47596 (N_47596,N_46725,N_46280);
or U47597 (N_47597,N_46355,N_46522);
xnor U47598 (N_47598,N_46895,N_46617);
nand U47599 (N_47599,N_46923,N_46367);
nand U47600 (N_47600,N_46154,N_46063);
nand U47601 (N_47601,N_46239,N_46795);
or U47602 (N_47602,N_46895,N_46836);
or U47603 (N_47603,N_46434,N_46913);
or U47604 (N_47604,N_46864,N_46035);
nand U47605 (N_47605,N_46127,N_46733);
nand U47606 (N_47606,N_46222,N_46463);
xor U47607 (N_47607,N_46785,N_46257);
and U47608 (N_47608,N_46707,N_46230);
and U47609 (N_47609,N_46512,N_46659);
xnor U47610 (N_47610,N_46702,N_46525);
nand U47611 (N_47611,N_46732,N_46252);
or U47612 (N_47612,N_46327,N_46071);
or U47613 (N_47613,N_46078,N_46205);
xor U47614 (N_47614,N_46963,N_46836);
or U47615 (N_47615,N_46658,N_46608);
and U47616 (N_47616,N_46204,N_46274);
or U47617 (N_47617,N_46784,N_46677);
xor U47618 (N_47618,N_46505,N_46782);
xor U47619 (N_47619,N_46020,N_46583);
nor U47620 (N_47620,N_46954,N_46218);
nand U47621 (N_47621,N_46645,N_46109);
and U47622 (N_47622,N_46807,N_46485);
nor U47623 (N_47623,N_46463,N_46408);
nor U47624 (N_47624,N_46479,N_46875);
and U47625 (N_47625,N_46032,N_46436);
nand U47626 (N_47626,N_46737,N_46946);
nor U47627 (N_47627,N_46790,N_46049);
nor U47628 (N_47628,N_46044,N_46417);
nor U47629 (N_47629,N_46536,N_46684);
or U47630 (N_47630,N_46305,N_46890);
and U47631 (N_47631,N_46930,N_46138);
nand U47632 (N_47632,N_46823,N_46464);
or U47633 (N_47633,N_46712,N_46333);
or U47634 (N_47634,N_46109,N_46565);
xor U47635 (N_47635,N_46018,N_46200);
nor U47636 (N_47636,N_46749,N_46326);
or U47637 (N_47637,N_46131,N_46332);
and U47638 (N_47638,N_46840,N_46577);
or U47639 (N_47639,N_46780,N_46046);
and U47640 (N_47640,N_46128,N_46909);
nor U47641 (N_47641,N_46611,N_46493);
nand U47642 (N_47642,N_46839,N_46037);
nand U47643 (N_47643,N_46329,N_46622);
and U47644 (N_47644,N_46709,N_46357);
nor U47645 (N_47645,N_46175,N_46988);
or U47646 (N_47646,N_46116,N_46991);
or U47647 (N_47647,N_46433,N_46220);
xor U47648 (N_47648,N_46789,N_46865);
nand U47649 (N_47649,N_46836,N_46288);
nand U47650 (N_47650,N_46231,N_46071);
nor U47651 (N_47651,N_46040,N_46195);
or U47652 (N_47652,N_46881,N_46734);
and U47653 (N_47653,N_46140,N_46988);
or U47654 (N_47654,N_46620,N_46257);
nor U47655 (N_47655,N_46024,N_46109);
or U47656 (N_47656,N_46742,N_46121);
or U47657 (N_47657,N_46916,N_46582);
and U47658 (N_47658,N_46927,N_46468);
and U47659 (N_47659,N_46614,N_46128);
nor U47660 (N_47660,N_46537,N_46285);
or U47661 (N_47661,N_46905,N_46500);
or U47662 (N_47662,N_46839,N_46758);
and U47663 (N_47663,N_46577,N_46477);
and U47664 (N_47664,N_46288,N_46013);
xor U47665 (N_47665,N_46275,N_46339);
xnor U47666 (N_47666,N_46131,N_46602);
nor U47667 (N_47667,N_46899,N_46958);
and U47668 (N_47668,N_46529,N_46059);
nor U47669 (N_47669,N_46214,N_46360);
and U47670 (N_47670,N_46058,N_46162);
and U47671 (N_47671,N_46148,N_46896);
nand U47672 (N_47672,N_46258,N_46948);
nand U47673 (N_47673,N_46172,N_46430);
or U47674 (N_47674,N_46939,N_46072);
or U47675 (N_47675,N_46899,N_46760);
and U47676 (N_47676,N_46750,N_46329);
and U47677 (N_47677,N_46811,N_46384);
and U47678 (N_47678,N_46098,N_46685);
nand U47679 (N_47679,N_46945,N_46294);
xnor U47680 (N_47680,N_46430,N_46139);
or U47681 (N_47681,N_46922,N_46505);
nand U47682 (N_47682,N_46008,N_46646);
xnor U47683 (N_47683,N_46530,N_46241);
xnor U47684 (N_47684,N_46216,N_46698);
xnor U47685 (N_47685,N_46887,N_46615);
and U47686 (N_47686,N_46243,N_46202);
xor U47687 (N_47687,N_46909,N_46699);
and U47688 (N_47688,N_46916,N_46113);
nand U47689 (N_47689,N_46037,N_46045);
xor U47690 (N_47690,N_46088,N_46244);
nor U47691 (N_47691,N_46433,N_46120);
or U47692 (N_47692,N_46860,N_46431);
nand U47693 (N_47693,N_46809,N_46440);
nand U47694 (N_47694,N_46124,N_46622);
or U47695 (N_47695,N_46084,N_46552);
nor U47696 (N_47696,N_46650,N_46697);
and U47697 (N_47697,N_46355,N_46514);
and U47698 (N_47698,N_46099,N_46522);
nor U47699 (N_47699,N_46384,N_46578);
xnor U47700 (N_47700,N_46098,N_46966);
xor U47701 (N_47701,N_46312,N_46861);
nor U47702 (N_47702,N_46002,N_46132);
nor U47703 (N_47703,N_46725,N_46212);
nor U47704 (N_47704,N_46300,N_46673);
nand U47705 (N_47705,N_46163,N_46910);
nor U47706 (N_47706,N_46304,N_46045);
or U47707 (N_47707,N_46317,N_46920);
nor U47708 (N_47708,N_46859,N_46542);
nand U47709 (N_47709,N_46833,N_46542);
and U47710 (N_47710,N_46976,N_46057);
or U47711 (N_47711,N_46653,N_46663);
nand U47712 (N_47712,N_46162,N_46450);
or U47713 (N_47713,N_46956,N_46092);
and U47714 (N_47714,N_46268,N_46076);
nor U47715 (N_47715,N_46917,N_46606);
nand U47716 (N_47716,N_46585,N_46810);
nor U47717 (N_47717,N_46627,N_46742);
xnor U47718 (N_47718,N_46014,N_46068);
or U47719 (N_47719,N_46305,N_46635);
nor U47720 (N_47720,N_46110,N_46242);
nor U47721 (N_47721,N_46441,N_46290);
nor U47722 (N_47722,N_46787,N_46733);
or U47723 (N_47723,N_46817,N_46184);
and U47724 (N_47724,N_46345,N_46301);
nor U47725 (N_47725,N_46884,N_46694);
xnor U47726 (N_47726,N_46922,N_46830);
xor U47727 (N_47727,N_46701,N_46808);
nand U47728 (N_47728,N_46124,N_46884);
or U47729 (N_47729,N_46901,N_46028);
nor U47730 (N_47730,N_46293,N_46141);
xnor U47731 (N_47731,N_46774,N_46240);
xor U47732 (N_47732,N_46048,N_46630);
or U47733 (N_47733,N_46080,N_46328);
or U47734 (N_47734,N_46604,N_46232);
and U47735 (N_47735,N_46210,N_46317);
nor U47736 (N_47736,N_46996,N_46407);
xnor U47737 (N_47737,N_46531,N_46391);
and U47738 (N_47738,N_46902,N_46444);
nor U47739 (N_47739,N_46658,N_46840);
xor U47740 (N_47740,N_46467,N_46611);
xnor U47741 (N_47741,N_46517,N_46048);
or U47742 (N_47742,N_46794,N_46812);
nor U47743 (N_47743,N_46703,N_46546);
nand U47744 (N_47744,N_46505,N_46102);
nand U47745 (N_47745,N_46077,N_46818);
nand U47746 (N_47746,N_46486,N_46821);
and U47747 (N_47747,N_46649,N_46328);
xnor U47748 (N_47748,N_46702,N_46745);
nor U47749 (N_47749,N_46051,N_46300);
nand U47750 (N_47750,N_46272,N_46609);
nand U47751 (N_47751,N_46089,N_46143);
or U47752 (N_47752,N_46256,N_46964);
and U47753 (N_47753,N_46931,N_46156);
nand U47754 (N_47754,N_46543,N_46753);
or U47755 (N_47755,N_46067,N_46232);
and U47756 (N_47756,N_46395,N_46812);
and U47757 (N_47757,N_46313,N_46609);
and U47758 (N_47758,N_46278,N_46730);
xnor U47759 (N_47759,N_46850,N_46546);
nand U47760 (N_47760,N_46393,N_46554);
or U47761 (N_47761,N_46368,N_46820);
nor U47762 (N_47762,N_46012,N_46217);
or U47763 (N_47763,N_46178,N_46314);
nor U47764 (N_47764,N_46447,N_46706);
and U47765 (N_47765,N_46960,N_46647);
nand U47766 (N_47766,N_46745,N_46160);
xnor U47767 (N_47767,N_46953,N_46469);
nand U47768 (N_47768,N_46749,N_46136);
nand U47769 (N_47769,N_46381,N_46369);
and U47770 (N_47770,N_46217,N_46259);
and U47771 (N_47771,N_46081,N_46373);
xor U47772 (N_47772,N_46447,N_46214);
nor U47773 (N_47773,N_46972,N_46301);
nand U47774 (N_47774,N_46847,N_46080);
or U47775 (N_47775,N_46924,N_46388);
xnor U47776 (N_47776,N_46766,N_46651);
or U47777 (N_47777,N_46487,N_46575);
and U47778 (N_47778,N_46013,N_46224);
and U47779 (N_47779,N_46937,N_46206);
and U47780 (N_47780,N_46794,N_46244);
nor U47781 (N_47781,N_46554,N_46743);
or U47782 (N_47782,N_46775,N_46377);
nand U47783 (N_47783,N_46600,N_46539);
xor U47784 (N_47784,N_46372,N_46908);
nand U47785 (N_47785,N_46519,N_46833);
and U47786 (N_47786,N_46280,N_46816);
nor U47787 (N_47787,N_46473,N_46133);
xnor U47788 (N_47788,N_46708,N_46419);
nor U47789 (N_47789,N_46887,N_46195);
or U47790 (N_47790,N_46357,N_46369);
nor U47791 (N_47791,N_46733,N_46492);
nand U47792 (N_47792,N_46322,N_46724);
xnor U47793 (N_47793,N_46087,N_46116);
nand U47794 (N_47794,N_46395,N_46853);
and U47795 (N_47795,N_46041,N_46767);
xnor U47796 (N_47796,N_46200,N_46359);
xor U47797 (N_47797,N_46388,N_46446);
or U47798 (N_47798,N_46809,N_46822);
or U47799 (N_47799,N_46007,N_46408);
nor U47800 (N_47800,N_46117,N_46162);
nand U47801 (N_47801,N_46313,N_46627);
nand U47802 (N_47802,N_46739,N_46973);
or U47803 (N_47803,N_46017,N_46787);
nand U47804 (N_47804,N_46904,N_46548);
and U47805 (N_47805,N_46592,N_46690);
nand U47806 (N_47806,N_46770,N_46572);
and U47807 (N_47807,N_46573,N_46746);
and U47808 (N_47808,N_46700,N_46308);
and U47809 (N_47809,N_46585,N_46919);
nand U47810 (N_47810,N_46785,N_46212);
xnor U47811 (N_47811,N_46249,N_46045);
nand U47812 (N_47812,N_46601,N_46782);
and U47813 (N_47813,N_46715,N_46816);
or U47814 (N_47814,N_46885,N_46318);
nor U47815 (N_47815,N_46771,N_46327);
nor U47816 (N_47816,N_46935,N_46253);
xor U47817 (N_47817,N_46345,N_46654);
nor U47818 (N_47818,N_46102,N_46646);
xnor U47819 (N_47819,N_46968,N_46475);
nand U47820 (N_47820,N_46559,N_46783);
and U47821 (N_47821,N_46597,N_46585);
nand U47822 (N_47822,N_46913,N_46403);
or U47823 (N_47823,N_46213,N_46851);
or U47824 (N_47824,N_46878,N_46865);
nor U47825 (N_47825,N_46711,N_46889);
and U47826 (N_47826,N_46136,N_46564);
nor U47827 (N_47827,N_46428,N_46313);
xnor U47828 (N_47828,N_46762,N_46030);
xor U47829 (N_47829,N_46257,N_46416);
xnor U47830 (N_47830,N_46213,N_46169);
xnor U47831 (N_47831,N_46497,N_46246);
nor U47832 (N_47832,N_46199,N_46711);
and U47833 (N_47833,N_46726,N_46176);
nand U47834 (N_47834,N_46188,N_46608);
xnor U47835 (N_47835,N_46678,N_46265);
xor U47836 (N_47836,N_46548,N_46824);
nor U47837 (N_47837,N_46408,N_46353);
xnor U47838 (N_47838,N_46166,N_46520);
and U47839 (N_47839,N_46026,N_46250);
xnor U47840 (N_47840,N_46790,N_46353);
nand U47841 (N_47841,N_46422,N_46769);
or U47842 (N_47842,N_46561,N_46052);
xnor U47843 (N_47843,N_46655,N_46809);
nor U47844 (N_47844,N_46518,N_46383);
and U47845 (N_47845,N_46403,N_46604);
xor U47846 (N_47846,N_46898,N_46115);
xor U47847 (N_47847,N_46664,N_46505);
and U47848 (N_47848,N_46280,N_46414);
and U47849 (N_47849,N_46594,N_46968);
nor U47850 (N_47850,N_46983,N_46295);
or U47851 (N_47851,N_46443,N_46560);
xnor U47852 (N_47852,N_46913,N_46451);
or U47853 (N_47853,N_46158,N_46707);
and U47854 (N_47854,N_46357,N_46129);
or U47855 (N_47855,N_46230,N_46314);
nor U47856 (N_47856,N_46392,N_46709);
xnor U47857 (N_47857,N_46245,N_46634);
or U47858 (N_47858,N_46342,N_46621);
xnor U47859 (N_47859,N_46530,N_46975);
or U47860 (N_47860,N_46929,N_46338);
or U47861 (N_47861,N_46199,N_46680);
nand U47862 (N_47862,N_46191,N_46462);
and U47863 (N_47863,N_46295,N_46894);
nand U47864 (N_47864,N_46276,N_46153);
or U47865 (N_47865,N_46309,N_46516);
or U47866 (N_47866,N_46074,N_46663);
nand U47867 (N_47867,N_46672,N_46080);
or U47868 (N_47868,N_46095,N_46945);
or U47869 (N_47869,N_46010,N_46603);
or U47870 (N_47870,N_46751,N_46451);
xor U47871 (N_47871,N_46411,N_46702);
and U47872 (N_47872,N_46450,N_46369);
nor U47873 (N_47873,N_46657,N_46058);
or U47874 (N_47874,N_46256,N_46172);
nor U47875 (N_47875,N_46441,N_46137);
or U47876 (N_47876,N_46592,N_46968);
and U47877 (N_47877,N_46484,N_46697);
nor U47878 (N_47878,N_46410,N_46211);
xnor U47879 (N_47879,N_46172,N_46132);
and U47880 (N_47880,N_46617,N_46257);
xor U47881 (N_47881,N_46309,N_46078);
nor U47882 (N_47882,N_46077,N_46439);
xor U47883 (N_47883,N_46430,N_46634);
or U47884 (N_47884,N_46767,N_46829);
or U47885 (N_47885,N_46360,N_46810);
nor U47886 (N_47886,N_46531,N_46726);
and U47887 (N_47887,N_46872,N_46116);
nor U47888 (N_47888,N_46217,N_46296);
nor U47889 (N_47889,N_46718,N_46179);
xor U47890 (N_47890,N_46107,N_46232);
nor U47891 (N_47891,N_46407,N_46080);
xor U47892 (N_47892,N_46294,N_46840);
and U47893 (N_47893,N_46062,N_46539);
or U47894 (N_47894,N_46342,N_46855);
nor U47895 (N_47895,N_46413,N_46268);
and U47896 (N_47896,N_46856,N_46426);
nand U47897 (N_47897,N_46963,N_46837);
nor U47898 (N_47898,N_46724,N_46136);
and U47899 (N_47899,N_46380,N_46888);
nand U47900 (N_47900,N_46740,N_46381);
nor U47901 (N_47901,N_46453,N_46423);
nor U47902 (N_47902,N_46637,N_46519);
nor U47903 (N_47903,N_46035,N_46406);
or U47904 (N_47904,N_46608,N_46064);
xor U47905 (N_47905,N_46874,N_46713);
and U47906 (N_47906,N_46194,N_46929);
nor U47907 (N_47907,N_46960,N_46191);
and U47908 (N_47908,N_46012,N_46048);
nand U47909 (N_47909,N_46767,N_46119);
nand U47910 (N_47910,N_46802,N_46793);
xor U47911 (N_47911,N_46433,N_46016);
xor U47912 (N_47912,N_46463,N_46572);
nand U47913 (N_47913,N_46365,N_46966);
and U47914 (N_47914,N_46517,N_46974);
xor U47915 (N_47915,N_46390,N_46380);
nor U47916 (N_47916,N_46410,N_46191);
xnor U47917 (N_47917,N_46970,N_46541);
nand U47918 (N_47918,N_46784,N_46321);
xor U47919 (N_47919,N_46540,N_46390);
and U47920 (N_47920,N_46654,N_46846);
nor U47921 (N_47921,N_46902,N_46905);
xor U47922 (N_47922,N_46999,N_46858);
nor U47923 (N_47923,N_46873,N_46221);
nor U47924 (N_47924,N_46486,N_46550);
xor U47925 (N_47925,N_46043,N_46703);
and U47926 (N_47926,N_46020,N_46268);
and U47927 (N_47927,N_46776,N_46351);
nand U47928 (N_47928,N_46498,N_46991);
nand U47929 (N_47929,N_46812,N_46592);
nor U47930 (N_47930,N_46506,N_46483);
xnor U47931 (N_47931,N_46874,N_46978);
or U47932 (N_47932,N_46893,N_46615);
and U47933 (N_47933,N_46858,N_46326);
xor U47934 (N_47934,N_46896,N_46732);
nand U47935 (N_47935,N_46239,N_46550);
and U47936 (N_47936,N_46536,N_46146);
nand U47937 (N_47937,N_46965,N_46959);
xor U47938 (N_47938,N_46439,N_46923);
nor U47939 (N_47939,N_46365,N_46661);
nor U47940 (N_47940,N_46705,N_46719);
or U47941 (N_47941,N_46744,N_46835);
or U47942 (N_47942,N_46661,N_46835);
or U47943 (N_47943,N_46189,N_46183);
and U47944 (N_47944,N_46077,N_46628);
or U47945 (N_47945,N_46168,N_46420);
xnor U47946 (N_47946,N_46850,N_46315);
xnor U47947 (N_47947,N_46437,N_46112);
nand U47948 (N_47948,N_46131,N_46330);
nor U47949 (N_47949,N_46452,N_46476);
xnor U47950 (N_47950,N_46967,N_46960);
xor U47951 (N_47951,N_46843,N_46096);
xnor U47952 (N_47952,N_46137,N_46885);
or U47953 (N_47953,N_46740,N_46467);
and U47954 (N_47954,N_46080,N_46795);
nand U47955 (N_47955,N_46649,N_46924);
or U47956 (N_47956,N_46907,N_46369);
or U47957 (N_47957,N_46120,N_46438);
or U47958 (N_47958,N_46680,N_46097);
nand U47959 (N_47959,N_46448,N_46025);
xor U47960 (N_47960,N_46163,N_46177);
and U47961 (N_47961,N_46140,N_46178);
or U47962 (N_47962,N_46273,N_46509);
nor U47963 (N_47963,N_46414,N_46166);
xnor U47964 (N_47964,N_46667,N_46578);
nor U47965 (N_47965,N_46086,N_46362);
and U47966 (N_47966,N_46948,N_46188);
nor U47967 (N_47967,N_46718,N_46401);
xnor U47968 (N_47968,N_46293,N_46453);
xnor U47969 (N_47969,N_46164,N_46259);
or U47970 (N_47970,N_46212,N_46573);
and U47971 (N_47971,N_46569,N_46899);
or U47972 (N_47972,N_46666,N_46126);
nand U47973 (N_47973,N_46087,N_46932);
nand U47974 (N_47974,N_46177,N_46821);
or U47975 (N_47975,N_46989,N_46570);
or U47976 (N_47976,N_46038,N_46307);
or U47977 (N_47977,N_46064,N_46933);
xor U47978 (N_47978,N_46673,N_46467);
nor U47979 (N_47979,N_46859,N_46930);
nand U47980 (N_47980,N_46018,N_46330);
nand U47981 (N_47981,N_46079,N_46729);
and U47982 (N_47982,N_46300,N_46109);
and U47983 (N_47983,N_46252,N_46297);
or U47984 (N_47984,N_46393,N_46290);
nor U47985 (N_47985,N_46355,N_46180);
or U47986 (N_47986,N_46664,N_46033);
or U47987 (N_47987,N_46601,N_46462);
and U47988 (N_47988,N_46607,N_46017);
or U47989 (N_47989,N_46422,N_46638);
and U47990 (N_47990,N_46540,N_46981);
nand U47991 (N_47991,N_46686,N_46702);
and U47992 (N_47992,N_46503,N_46732);
nor U47993 (N_47993,N_46887,N_46244);
nand U47994 (N_47994,N_46260,N_46380);
and U47995 (N_47995,N_46341,N_46321);
xor U47996 (N_47996,N_46318,N_46484);
xor U47997 (N_47997,N_46802,N_46187);
xnor U47998 (N_47998,N_46386,N_46260);
and U47999 (N_47999,N_46352,N_46845);
nor U48000 (N_48000,N_47254,N_47091);
xor U48001 (N_48001,N_47675,N_47443);
and U48002 (N_48002,N_47304,N_47578);
nand U48003 (N_48003,N_47402,N_47914);
xor U48004 (N_48004,N_47556,N_47761);
and U48005 (N_48005,N_47856,N_47251);
nor U48006 (N_48006,N_47013,N_47234);
nor U48007 (N_48007,N_47472,N_47613);
nand U48008 (N_48008,N_47296,N_47282);
xor U48009 (N_48009,N_47899,N_47961);
nand U48010 (N_48010,N_47575,N_47098);
xor U48011 (N_48011,N_47804,N_47763);
and U48012 (N_48012,N_47186,N_47680);
or U48013 (N_48013,N_47765,N_47330);
or U48014 (N_48014,N_47464,N_47998);
and U48015 (N_48015,N_47805,N_47191);
and U48016 (N_48016,N_47302,N_47642);
and U48017 (N_48017,N_47696,N_47429);
nor U48018 (N_48018,N_47218,N_47999);
nand U48019 (N_48019,N_47517,N_47648);
or U48020 (N_48020,N_47983,N_47801);
nor U48021 (N_48021,N_47310,N_47023);
xor U48022 (N_48022,N_47984,N_47123);
and U48023 (N_48023,N_47551,N_47256);
xnor U48024 (N_48024,N_47930,N_47270);
and U48025 (N_48025,N_47986,N_47548);
or U48026 (N_48026,N_47352,N_47547);
nand U48027 (N_48027,N_47272,N_47668);
nor U48028 (N_48028,N_47824,N_47810);
nor U48029 (N_48029,N_47513,N_47058);
xor U48030 (N_48030,N_47397,N_47408);
or U48031 (N_48031,N_47629,N_47711);
or U48032 (N_48032,N_47424,N_47299);
nor U48033 (N_48033,N_47002,N_47284);
xnor U48034 (N_48034,N_47670,N_47661);
or U48035 (N_48035,N_47571,N_47677);
or U48036 (N_48036,N_47518,N_47647);
xnor U48037 (N_48037,N_47562,N_47393);
xor U48038 (N_48038,N_47250,N_47292);
xnor U48039 (N_48039,N_47275,N_47946);
and U48040 (N_48040,N_47932,N_47701);
and U48041 (N_48041,N_47372,N_47414);
nand U48042 (N_48042,N_47877,N_47707);
or U48043 (N_48043,N_47697,N_47830);
and U48044 (N_48044,N_47404,N_47364);
nand U48045 (N_48045,N_47271,N_47576);
and U48046 (N_48046,N_47175,N_47796);
xor U48047 (N_48047,N_47523,N_47622);
nor U48048 (N_48048,N_47970,N_47014);
or U48049 (N_48049,N_47850,N_47486);
xor U48050 (N_48050,N_47913,N_47164);
or U48051 (N_48051,N_47503,N_47423);
and U48052 (N_48052,N_47638,N_47832);
or U48053 (N_48053,N_47734,N_47106);
xor U48054 (N_48054,N_47311,N_47498);
nand U48055 (N_48055,N_47569,N_47315);
and U48056 (N_48056,N_47216,N_47005);
or U48057 (N_48057,N_47199,N_47229);
or U48058 (N_48058,N_47470,N_47589);
and U48059 (N_48059,N_47502,N_47236);
or U48060 (N_48060,N_47965,N_47545);
or U48061 (N_48061,N_47174,N_47268);
xor U48062 (N_48062,N_47626,N_47855);
nand U48063 (N_48063,N_47845,N_47185);
and U48064 (N_48064,N_47156,N_47620);
nor U48065 (N_48065,N_47957,N_47603);
xnor U48066 (N_48066,N_47431,N_47122);
and U48067 (N_48067,N_47510,N_47777);
nor U48068 (N_48068,N_47827,N_47025);
xnor U48069 (N_48069,N_47528,N_47361);
xor U48070 (N_48070,N_47066,N_47048);
and U48071 (N_48071,N_47289,N_47055);
nand U48072 (N_48072,N_47099,N_47690);
xor U48073 (N_48073,N_47771,N_47349);
and U48074 (N_48074,N_47394,N_47323);
nand U48075 (N_48075,N_47803,N_47053);
nor U48076 (N_48076,N_47729,N_47504);
nor U48077 (N_48077,N_47604,N_47587);
nor U48078 (N_48078,N_47076,N_47662);
xnor U48079 (N_48079,N_47125,N_47356);
nand U48080 (N_48080,N_47557,N_47406);
xor U48081 (N_48081,N_47415,N_47886);
and U48082 (N_48082,N_47499,N_47781);
nor U48083 (N_48083,N_47150,N_47410);
and U48084 (N_48084,N_47420,N_47463);
and U48085 (N_48085,N_47319,N_47445);
nor U48086 (N_48086,N_47501,N_47248);
xnor U48087 (N_48087,N_47317,N_47552);
xnor U48088 (N_48088,N_47522,N_47770);
and U48089 (N_48089,N_47829,N_47081);
nor U48090 (N_48090,N_47258,N_47934);
xor U48091 (N_48091,N_47067,N_47838);
nand U48092 (N_48092,N_47800,N_47221);
nand U48093 (N_48093,N_47573,N_47339);
nor U48094 (N_48094,N_47039,N_47274);
nor U48095 (N_48095,N_47792,N_47419);
and U48096 (N_48096,N_47943,N_47674);
or U48097 (N_48097,N_47795,N_47514);
or U48098 (N_48098,N_47778,N_47812);
nand U48099 (N_48099,N_47187,N_47568);
nand U48100 (N_48100,N_47911,N_47375);
nor U48101 (N_48101,N_47931,N_47779);
nand U48102 (N_48102,N_47612,N_47749);
nor U48103 (N_48103,N_47412,N_47997);
and U48104 (N_48104,N_47338,N_47045);
xnor U48105 (N_48105,N_47403,N_47480);
xor U48106 (N_48106,N_47793,N_47298);
nand U48107 (N_48107,N_47724,N_47471);
nor U48108 (N_48108,N_47136,N_47512);
and U48109 (N_48109,N_47667,N_47206);
and U48110 (N_48110,N_47259,N_47226);
and U48111 (N_48111,N_47698,N_47625);
nand U48112 (N_48112,N_47280,N_47909);
nor U48113 (N_48113,N_47484,N_47822);
nand U48114 (N_48114,N_47321,N_47482);
nor U48115 (N_48115,N_47332,N_47614);
or U48116 (N_48116,N_47828,N_47363);
nor U48117 (N_48117,N_47851,N_47900);
xor U48118 (N_48118,N_47083,N_47505);
nand U48119 (N_48119,N_47193,N_47333);
and U48120 (N_48120,N_47741,N_47813);
nand U48121 (N_48121,N_47168,N_47097);
or U48122 (N_48122,N_47586,N_47920);
nor U48123 (N_48123,N_47991,N_47712);
and U48124 (N_48124,N_47705,N_47555);
xor U48125 (N_48125,N_47543,N_47146);
nor U48126 (N_48126,N_47010,N_47689);
nand U48127 (N_48127,N_47788,N_47026);
or U48128 (N_48128,N_47672,N_47059);
and U48129 (N_48129,N_47879,N_47411);
and U48130 (N_48130,N_47633,N_47244);
nor U48131 (N_48131,N_47782,N_47452);
nand U48132 (N_48132,N_47540,N_47837);
or U48133 (N_48133,N_47354,N_47996);
xor U48134 (N_48134,N_47645,N_47541);
xor U48135 (N_48135,N_47024,N_47774);
nand U48136 (N_48136,N_47883,N_47987);
nor U48137 (N_48137,N_47173,N_47857);
nor U48138 (N_48138,N_47882,N_47331);
xnor U48139 (N_48139,N_47912,N_47316);
or U48140 (N_48140,N_47862,N_47885);
or U48141 (N_48141,N_47903,N_47184);
nor U48142 (N_48142,N_47069,N_47746);
nor U48143 (N_48143,N_47001,N_47153);
xor U48144 (N_48144,N_47038,N_47927);
nor U48145 (N_48145,N_47172,N_47699);
nor U48146 (N_48146,N_47073,N_47599);
nand U48147 (N_48147,N_47643,N_47385);
and U48148 (N_48148,N_47937,N_47151);
or U48149 (N_48149,N_47003,N_47861);
or U48150 (N_48150,N_47956,N_47806);
and U48151 (N_48151,N_47869,N_47748);
xnor U48152 (N_48152,N_47371,N_47736);
or U48153 (N_48153,N_47863,N_47119);
or U48154 (N_48154,N_47876,N_47112);
nor U48155 (N_48155,N_47659,N_47233);
nor U48156 (N_48156,N_47092,N_47581);
nand U48157 (N_48157,N_47080,N_47227);
xor U48158 (N_48158,N_47816,N_47181);
nand U48159 (N_48159,N_47290,N_47731);
or U48160 (N_48160,N_47866,N_47052);
nand U48161 (N_48161,N_47938,N_47031);
and U48162 (N_48162,N_47209,N_47117);
nor U48163 (N_48163,N_47834,N_47871);
or U48164 (N_48164,N_47017,N_47347);
xnor U48165 (N_48165,N_47606,N_47867);
and U48166 (N_48166,N_47190,N_47644);
and U48167 (N_48167,N_47084,N_47466);
nand U48168 (N_48168,N_47213,N_47751);
or U48169 (N_48169,N_47074,N_47183);
xor U48170 (N_48170,N_47362,N_47618);
nor U48171 (N_48171,N_47046,N_47716);
nand U48172 (N_48172,N_47988,N_47958);
and U48173 (N_48173,N_47760,N_47596);
nand U48174 (N_48174,N_47437,N_47809);
nor U48175 (N_48175,N_47020,N_47567);
xor U48176 (N_48176,N_47101,N_47343);
nand U48177 (N_48177,N_47239,N_47859);
xnor U48178 (N_48178,N_47341,N_47008);
or U48179 (N_48179,N_47088,N_47468);
nor U48180 (N_48180,N_47458,N_47844);
and U48181 (N_48181,N_47149,N_47278);
nand U48182 (N_48182,N_47497,N_47500);
nand U48183 (N_48183,N_47678,N_47494);
or U48184 (N_48184,N_47391,N_47245);
and U48185 (N_48185,N_47688,N_47337);
nor U48186 (N_48186,N_47665,N_47169);
xor U48187 (N_48187,N_47973,N_47444);
nand U48188 (N_48188,N_47605,N_47483);
or U48189 (N_48189,N_47742,N_47351);
nand U48190 (N_48190,N_47089,N_47840);
or U48191 (N_48191,N_47653,N_47893);
nor U48192 (N_48192,N_47496,N_47635);
nor U48193 (N_48193,N_47446,N_47491);
nor U48194 (N_48194,N_47728,N_47691);
nor U48195 (N_48195,N_47407,N_47891);
and U48196 (N_48196,N_47610,N_47959);
nor U48197 (N_48197,N_47950,N_47060);
xnor U48198 (N_48198,N_47880,N_47739);
nor U48199 (N_48199,N_47474,N_47888);
nand U48200 (N_48200,N_47579,N_47242);
nand U48201 (N_48201,N_47057,N_47945);
or U48202 (N_48202,N_47135,N_47454);
nor U48203 (N_48203,N_47560,N_47447);
or U48204 (N_48204,N_47919,N_47154);
or U48205 (N_48205,N_47232,N_47249);
nand U48206 (N_48206,N_47238,N_47582);
nor U48207 (N_48207,N_47884,N_47344);
and U48208 (N_48208,N_47720,N_47821);
nand U48209 (N_48209,N_47421,N_47157);
nor U48210 (N_48210,N_47260,N_47584);
or U48211 (N_48211,N_47846,N_47875);
nor U48212 (N_48212,N_47124,N_47949);
xnor U48213 (N_48213,N_47536,N_47892);
nand U48214 (N_48214,N_47217,N_47188);
or U48215 (N_48215,N_47116,N_47322);
nand U48216 (N_48216,N_47944,N_47353);
or U48217 (N_48217,N_47030,N_47598);
xor U48218 (N_48218,N_47980,N_47435);
nand U48219 (N_48219,N_47954,N_47147);
nor U48220 (N_48220,N_47365,N_47758);
or U48221 (N_48221,N_47107,N_47225);
and U48222 (N_48222,N_47974,N_47253);
or U48223 (N_48223,N_47926,N_47434);
nor U48224 (N_48224,N_47159,N_47416);
nand U48225 (N_48225,N_47607,N_47537);
or U48226 (N_48226,N_47901,N_47594);
nor U48227 (N_48227,N_47370,N_47422);
nor U48228 (N_48228,N_47704,N_47355);
or U48229 (N_48229,N_47049,N_47087);
or U48230 (N_48230,N_47526,N_47652);
nand U48231 (N_48231,N_47207,N_47897);
nor U48232 (N_48232,N_47525,N_47843);
nand U48233 (N_48233,N_47047,N_47636);
nor U48234 (N_48234,N_47747,N_47348);
or U48235 (N_48235,N_47395,N_47390);
nor U48236 (N_48236,N_47657,N_47405);
or U48237 (N_48237,N_47448,N_47947);
nor U48238 (N_48238,N_47865,N_47095);
xor U48239 (N_48239,N_47487,N_47671);
nand U48240 (N_48240,N_47007,N_47574);
xor U48241 (N_48241,N_47971,N_47791);
and U48242 (N_48242,N_47588,N_47917);
or U48243 (N_48243,N_47683,N_47179);
and U48244 (N_48244,N_47127,N_47538);
xor U48245 (N_48245,N_47440,N_47577);
xnor U48246 (N_48246,N_47787,N_47068);
or U48247 (N_48247,N_47294,N_47915);
nor U48248 (N_48248,N_47161,N_47759);
xnor U48249 (N_48249,N_47286,N_47195);
nand U48250 (N_48250,N_47709,N_47768);
nand U48251 (N_48251,N_47817,N_47703);
and U48252 (N_48252,N_47976,N_47539);
xor U48253 (N_48253,N_47121,N_47293);
and U48254 (N_48254,N_47281,N_47532);
nand U48255 (N_48255,N_47075,N_47379);
or U48256 (N_48256,N_47114,N_47040);
nor U48257 (N_48257,N_47750,N_47336);
or U48258 (N_48258,N_47602,N_47077);
or U48259 (N_48259,N_47212,N_47632);
nor U48260 (N_48260,N_47940,N_47328);
nand U48261 (N_48261,N_47243,N_47035);
xnor U48262 (N_48262,N_47790,N_47165);
xor U48263 (N_48263,N_47767,N_47962);
nor U48264 (N_48264,N_47094,N_47326);
or U48265 (N_48265,N_47283,N_47418);
nor U48266 (N_48266,N_47743,N_47327);
and U48267 (N_48267,N_47033,N_47490);
nand U48268 (N_48268,N_47554,N_47019);
nand U48269 (N_48269,N_47120,N_47318);
xnor U48270 (N_48270,N_47969,N_47433);
or U48271 (N_48271,N_47714,N_47324);
xnor U48272 (N_48272,N_47797,N_47194);
nor U48273 (N_48273,N_47717,N_47307);
nor U48274 (N_48274,N_47432,N_47627);
or U48275 (N_48275,N_47478,N_47475);
nor U48276 (N_48276,N_47687,N_47263);
and U48277 (N_48277,N_47651,N_47754);
xnor U48278 (N_48278,N_47182,N_47223);
xnor U48279 (N_48279,N_47219,N_47426);
nand U48280 (N_48280,N_47203,N_47167);
nand U48281 (N_48281,N_47802,N_47507);
and U48282 (N_48282,N_47710,N_47860);
and U48283 (N_48283,N_47684,N_47706);
and U48284 (N_48284,N_47065,N_47898);
and U48285 (N_48285,N_47142,N_47308);
nand U48286 (N_48286,N_47848,N_47438);
nor U48287 (N_48287,N_47872,N_47312);
nand U48288 (N_48288,N_47220,N_47392);
nand U48289 (N_48289,N_47692,N_47237);
nand U48290 (N_48290,N_47814,N_47138);
xor U48291 (N_48291,N_47616,N_47305);
nor U48292 (N_48292,N_47085,N_47745);
nand U48293 (N_48293,N_47807,N_47941);
and U48294 (N_48294,N_47388,N_47713);
nand U48295 (N_48295,N_47527,N_47935);
and U48296 (N_48296,N_47533,N_47939);
or U48297 (N_48297,N_47131,N_47495);
xor U48298 (N_48298,N_47744,N_47450);
and U48299 (N_48299,N_47902,N_47032);
nand U48300 (N_48300,N_47211,N_47108);
nand U48301 (N_48301,N_47439,N_47295);
nor U48302 (N_48302,N_47350,N_47204);
nor U48303 (N_48303,N_47277,N_47300);
xnor U48304 (N_48304,N_47320,N_47043);
xnor U48305 (N_48305,N_47104,N_47849);
xnor U48306 (N_48306,N_47925,N_47580);
or U48307 (N_48307,N_47600,N_47649);
and U48308 (N_48308,N_47905,N_47126);
nand U48309 (N_48309,N_47477,N_47978);
xnor U48310 (N_48310,N_47255,N_47853);
nor U48311 (N_48311,N_47544,N_47715);
nand U48312 (N_48312,N_47386,N_47951);
and U48313 (N_48313,N_47000,N_47210);
nand U48314 (N_48314,N_47521,N_47881);
or U48315 (N_48315,N_47178,N_47467);
nor U48316 (N_48316,N_47357,N_47384);
and U48317 (N_48317,N_47982,N_47064);
and U48318 (N_48318,N_47006,N_47921);
and U48319 (N_48319,N_47368,N_47459);
nand U48320 (N_48320,N_47011,N_47456);
xnor U48321 (N_48321,N_47655,N_47623);
or U48322 (N_48322,N_47966,N_47918);
or U48323 (N_48323,N_47550,N_47868);
or U48324 (N_48324,N_47342,N_47723);
xor U48325 (N_48325,N_47798,N_47534);
and U48326 (N_48326,N_47180,N_47485);
nand U48327 (N_48327,N_47819,N_47906);
xor U48328 (N_48328,N_47041,N_47208);
and U48329 (N_48329,N_47531,N_47037);
and U48330 (N_48330,N_47972,N_47702);
xnor U48331 (N_48331,N_47228,N_47593);
nand U48332 (N_48332,N_47409,N_47676);
nor U48333 (N_48333,N_47462,N_47725);
and U48334 (N_48334,N_47631,N_47874);
and U48335 (N_48335,N_47858,N_47093);
nand U48336 (N_48336,N_47383,N_47894);
nand U48337 (N_48337,N_47764,N_47994);
or U48338 (N_48338,N_47786,N_47162);
and U48339 (N_48339,N_47262,N_47451);
and U48340 (N_48340,N_47654,N_47028);
and U48341 (N_48341,N_47722,N_47340);
and U48342 (N_48342,N_47133,N_47910);
nand U48343 (N_48343,N_47492,N_47382);
nor U48344 (N_48344,N_47380,N_47646);
or U48345 (N_48345,N_47737,N_47481);
or U48346 (N_48346,N_47726,N_47685);
nor U48347 (N_48347,N_47285,N_47265);
nor U48348 (N_48348,N_47009,N_47663);
nand U48349 (N_48349,N_47542,N_47794);
and U48350 (N_48350,N_47297,N_47465);
or U48351 (N_48351,N_47682,N_47441);
nor U48352 (N_48352,N_47718,N_47109);
and U48353 (N_48353,N_47266,N_47100);
xnor U48354 (N_48354,N_47279,N_47034);
xnor U48355 (N_48355,N_47325,N_47158);
xnor U48356 (N_48356,N_47955,N_47303);
or U48357 (N_48357,N_47565,N_47854);
or U48358 (N_48358,N_47769,N_47110);
nor U48359 (N_48359,N_47137,N_47753);
or U48360 (N_48360,N_47953,N_47755);
and U48361 (N_48361,N_47784,N_47287);
nor U48362 (N_48362,N_47130,N_47942);
nand U48363 (N_48363,N_47072,N_47833);
xor U48364 (N_48364,N_47460,N_47735);
nor U48365 (N_48365,N_47373,N_47847);
or U48366 (N_48366,N_47924,N_47508);
and U48367 (N_48367,N_47170,N_47063);
and U48368 (N_48368,N_47314,N_47374);
nor U48369 (N_48369,N_47398,N_47608);
nor U48370 (N_48370,N_47177,N_47776);
nor U48371 (N_48371,N_47401,N_47358);
and U48372 (N_48372,N_47078,N_47042);
or U48373 (N_48373,N_47595,N_47660);
xnor U48374 (N_48374,N_47489,N_47928);
and U48375 (N_48375,N_47141,N_47870);
or U48376 (N_48376,N_47115,N_47772);
or U48377 (N_48377,N_47686,N_47476);
and U48378 (N_48378,N_47963,N_47591);
nand U48379 (N_48379,N_47430,N_47214);
and U48380 (N_48380,N_47695,N_47740);
and U48381 (N_48381,N_47570,N_47252);
or U48382 (N_48382,N_47873,N_47785);
or U48383 (N_48383,N_47139,N_47975);
nand U48384 (N_48384,N_47773,N_47818);
nor U48385 (N_48385,N_47442,N_47730);
and U48386 (N_48386,N_47733,N_47823);
nor U48387 (N_48387,N_47839,N_47634);
or U48388 (N_48388,N_47488,N_47479);
xnor U48389 (N_48389,N_47198,N_47896);
xnor U48390 (N_48390,N_47826,N_47396);
xor U48391 (N_48391,N_47916,N_47417);
nand U48392 (N_48392,N_47641,N_47990);
nor U48393 (N_48393,N_47143,N_47968);
nor U48394 (N_48394,N_47658,N_47639);
and U48395 (N_48395,N_47389,N_47656);
xnor U48396 (N_48396,N_47134,N_47205);
nand U48397 (N_48397,N_47148,N_47269);
and U48398 (N_48398,N_47449,N_47096);
and U48399 (N_48399,N_47062,N_47273);
nor U48400 (N_48400,N_47511,N_47852);
nand U48401 (N_48401,N_47050,N_47756);
nand U48402 (N_48402,N_47700,N_47335);
xnor U48403 (N_48403,N_47637,N_47140);
nor U48404 (N_48404,N_47789,N_47288);
and U48405 (N_48405,N_47673,N_47611);
and U48406 (N_48406,N_47309,N_47276);
or U48407 (N_48407,N_47895,N_47820);
nand U48408 (N_48408,N_47118,N_47246);
nand U48409 (N_48409,N_47473,N_47979);
and U48410 (N_48410,N_47530,N_47904);
and U48411 (N_48411,N_47235,N_47021);
nor U48412 (N_48412,N_47376,N_47952);
nand U48413 (N_48413,N_47329,N_47012);
nand U48414 (N_48414,N_47346,N_47546);
xnor U48415 (N_48415,N_47775,N_47400);
or U48416 (N_48416,N_47624,N_47842);
nor U48417 (N_48417,N_47360,N_47129);
xor U48418 (N_48418,N_47241,N_47176);
and U48419 (N_48419,N_47145,N_47630);
xor U48420 (N_48420,N_47313,N_47036);
or U48421 (N_48421,N_47985,N_47694);
or U48422 (N_48422,N_47301,N_47054);
and U48423 (N_48423,N_47381,N_47436);
and U48424 (N_48424,N_47202,N_47825);
and U48425 (N_48425,N_47615,N_47564);
and U48426 (N_48426,N_47732,N_47079);
nor U48427 (N_48427,N_47964,N_47132);
nand U48428 (N_48428,N_47061,N_47572);
or U48429 (N_48429,N_47808,N_47609);
and U48430 (N_48430,N_47948,N_47922);
nand U48431 (N_48431,N_47345,N_47506);
or U48432 (N_48432,N_47889,N_47166);
nor U48433 (N_48433,N_47493,N_47650);
xor U48434 (N_48434,N_47192,N_47359);
nand U48435 (N_48435,N_47619,N_47051);
xor U48436 (N_48436,N_47469,N_47590);
nand U48437 (N_48437,N_47831,N_47524);
xnor U48438 (N_48438,N_47836,N_47669);
nand U48439 (N_48439,N_47369,N_47908);
or U48440 (N_48440,N_47222,N_47334);
and U48441 (N_48441,N_47509,N_47783);
nor U48442 (N_48442,N_47907,N_47721);
nor U48443 (N_48443,N_47103,N_47887);
nor U48444 (N_48444,N_47936,N_47231);
nor U48445 (N_48445,N_47780,N_47261);
or U48446 (N_48446,N_47977,N_47247);
or U48447 (N_48447,N_47022,N_47144);
or U48448 (N_48448,N_47291,N_47549);
nand U48449 (N_48449,N_47617,N_47455);
nor U48450 (N_48450,N_47757,N_47535);
nand U48451 (N_48451,N_47558,N_47111);
or U48452 (N_48452,N_47993,N_47529);
xor U48453 (N_48453,N_47128,N_47841);
or U48454 (N_48454,N_47044,N_47923);
xnor U48455 (N_48455,N_47693,N_47240);
and U48456 (N_48456,N_47457,N_47727);
nor U48457 (N_48457,N_47864,N_47799);
nor U48458 (N_48458,N_47811,N_47519);
and U48459 (N_48459,N_47306,N_47082);
or U48460 (N_48460,N_47762,N_47428);
or U48461 (N_48461,N_47399,N_47163);
and U48462 (N_48462,N_47015,N_47461);
or U48463 (N_48463,N_47427,N_47230);
or U48464 (N_48464,N_47257,N_47664);
nand U48465 (N_48465,N_47520,N_47621);
xor U48466 (N_48466,N_47553,N_47835);
nor U48467 (N_48467,N_47981,N_47878);
and U48468 (N_48468,N_47515,N_47933);
nor U48469 (N_48469,N_47666,N_47267);
and U48470 (N_48470,N_47070,N_47592);
nor U48471 (N_48471,N_47413,N_47929);
xor U48472 (N_48472,N_47090,N_47601);
nor U48473 (N_48473,N_47171,N_47566);
or U48474 (N_48474,N_47102,N_47815);
nor U48475 (N_48475,N_47366,N_47640);
or U48476 (N_48476,N_47585,N_47583);
nand U48477 (N_48477,N_47152,N_47752);
xnor U48478 (N_48478,N_47377,N_47995);
or U48479 (N_48479,N_47113,N_47367);
nand U48480 (N_48480,N_47890,N_47197);
or U48481 (N_48481,N_47201,N_47027);
xor U48482 (N_48482,N_47004,N_47029);
nor U48483 (N_48483,N_47563,N_47597);
nor U48484 (N_48484,N_47453,N_47967);
or U48485 (N_48485,N_47378,N_47189);
nand U48486 (N_48486,N_47992,N_47679);
nand U48487 (N_48487,N_47708,N_47561);
xnor U48488 (N_48488,N_47155,N_47766);
or U48489 (N_48489,N_47071,N_47016);
xor U48490 (N_48490,N_47264,N_47086);
xor U48491 (N_48491,N_47387,N_47516);
nor U48492 (N_48492,N_47196,N_47425);
nor U48493 (N_48493,N_47224,N_47200);
xnor U48494 (N_48494,N_47628,N_47105);
nand U48495 (N_48495,N_47719,N_47559);
xnor U48496 (N_48496,N_47681,N_47018);
and U48497 (N_48497,N_47960,N_47056);
xnor U48498 (N_48498,N_47989,N_47160);
xnor U48499 (N_48499,N_47738,N_47215);
or U48500 (N_48500,N_47762,N_47605);
nor U48501 (N_48501,N_47606,N_47575);
nor U48502 (N_48502,N_47757,N_47172);
and U48503 (N_48503,N_47468,N_47471);
nand U48504 (N_48504,N_47617,N_47975);
or U48505 (N_48505,N_47654,N_47644);
nand U48506 (N_48506,N_47117,N_47413);
xnor U48507 (N_48507,N_47718,N_47942);
and U48508 (N_48508,N_47558,N_47971);
and U48509 (N_48509,N_47149,N_47622);
xor U48510 (N_48510,N_47291,N_47753);
nand U48511 (N_48511,N_47567,N_47733);
nor U48512 (N_48512,N_47957,N_47535);
nand U48513 (N_48513,N_47312,N_47155);
nand U48514 (N_48514,N_47694,N_47902);
and U48515 (N_48515,N_47663,N_47413);
nor U48516 (N_48516,N_47277,N_47901);
or U48517 (N_48517,N_47003,N_47910);
and U48518 (N_48518,N_47429,N_47139);
nor U48519 (N_48519,N_47545,N_47699);
xor U48520 (N_48520,N_47595,N_47158);
and U48521 (N_48521,N_47579,N_47787);
or U48522 (N_48522,N_47332,N_47633);
and U48523 (N_48523,N_47230,N_47126);
xor U48524 (N_48524,N_47433,N_47859);
nor U48525 (N_48525,N_47980,N_47998);
xnor U48526 (N_48526,N_47848,N_47606);
xor U48527 (N_48527,N_47688,N_47760);
or U48528 (N_48528,N_47587,N_47483);
nor U48529 (N_48529,N_47083,N_47899);
and U48530 (N_48530,N_47947,N_47658);
nand U48531 (N_48531,N_47597,N_47890);
or U48532 (N_48532,N_47540,N_47144);
or U48533 (N_48533,N_47688,N_47643);
xnor U48534 (N_48534,N_47413,N_47704);
and U48535 (N_48535,N_47003,N_47733);
nand U48536 (N_48536,N_47135,N_47905);
and U48537 (N_48537,N_47412,N_47223);
nand U48538 (N_48538,N_47392,N_47339);
xnor U48539 (N_48539,N_47134,N_47577);
xnor U48540 (N_48540,N_47590,N_47642);
nor U48541 (N_48541,N_47107,N_47426);
nand U48542 (N_48542,N_47672,N_47855);
nor U48543 (N_48543,N_47253,N_47159);
xor U48544 (N_48544,N_47860,N_47347);
and U48545 (N_48545,N_47691,N_47375);
nor U48546 (N_48546,N_47051,N_47848);
xnor U48547 (N_48547,N_47006,N_47100);
nor U48548 (N_48548,N_47378,N_47656);
nand U48549 (N_48549,N_47338,N_47894);
nor U48550 (N_48550,N_47222,N_47028);
or U48551 (N_48551,N_47929,N_47470);
and U48552 (N_48552,N_47710,N_47425);
nand U48553 (N_48553,N_47442,N_47299);
nor U48554 (N_48554,N_47599,N_47749);
xor U48555 (N_48555,N_47703,N_47901);
xor U48556 (N_48556,N_47022,N_47915);
xnor U48557 (N_48557,N_47953,N_47882);
and U48558 (N_48558,N_47251,N_47016);
or U48559 (N_48559,N_47184,N_47362);
xnor U48560 (N_48560,N_47262,N_47691);
nor U48561 (N_48561,N_47821,N_47628);
nor U48562 (N_48562,N_47392,N_47905);
and U48563 (N_48563,N_47589,N_47416);
xor U48564 (N_48564,N_47813,N_47370);
or U48565 (N_48565,N_47747,N_47844);
xnor U48566 (N_48566,N_47185,N_47919);
xnor U48567 (N_48567,N_47715,N_47983);
xor U48568 (N_48568,N_47325,N_47802);
xnor U48569 (N_48569,N_47992,N_47907);
and U48570 (N_48570,N_47167,N_47698);
or U48571 (N_48571,N_47214,N_47947);
xor U48572 (N_48572,N_47161,N_47381);
and U48573 (N_48573,N_47104,N_47938);
or U48574 (N_48574,N_47213,N_47977);
xor U48575 (N_48575,N_47103,N_47436);
and U48576 (N_48576,N_47515,N_47860);
nand U48577 (N_48577,N_47314,N_47699);
xnor U48578 (N_48578,N_47984,N_47036);
or U48579 (N_48579,N_47975,N_47575);
nor U48580 (N_48580,N_47116,N_47814);
and U48581 (N_48581,N_47207,N_47317);
nor U48582 (N_48582,N_47925,N_47744);
nor U48583 (N_48583,N_47191,N_47437);
xor U48584 (N_48584,N_47925,N_47194);
xnor U48585 (N_48585,N_47219,N_47735);
nand U48586 (N_48586,N_47434,N_47383);
or U48587 (N_48587,N_47808,N_47900);
nor U48588 (N_48588,N_47598,N_47547);
and U48589 (N_48589,N_47211,N_47293);
xor U48590 (N_48590,N_47059,N_47912);
nor U48591 (N_48591,N_47088,N_47679);
and U48592 (N_48592,N_47079,N_47181);
xor U48593 (N_48593,N_47385,N_47145);
nand U48594 (N_48594,N_47291,N_47367);
xor U48595 (N_48595,N_47570,N_47868);
and U48596 (N_48596,N_47569,N_47225);
xor U48597 (N_48597,N_47737,N_47023);
or U48598 (N_48598,N_47949,N_47583);
or U48599 (N_48599,N_47006,N_47103);
nand U48600 (N_48600,N_47206,N_47373);
and U48601 (N_48601,N_47854,N_47042);
nor U48602 (N_48602,N_47345,N_47430);
nand U48603 (N_48603,N_47900,N_47611);
and U48604 (N_48604,N_47784,N_47225);
xnor U48605 (N_48605,N_47409,N_47636);
nand U48606 (N_48606,N_47661,N_47911);
nand U48607 (N_48607,N_47418,N_47449);
xor U48608 (N_48608,N_47247,N_47075);
nand U48609 (N_48609,N_47409,N_47262);
nand U48610 (N_48610,N_47726,N_47082);
or U48611 (N_48611,N_47082,N_47811);
nor U48612 (N_48612,N_47247,N_47036);
nor U48613 (N_48613,N_47873,N_47420);
and U48614 (N_48614,N_47489,N_47977);
xor U48615 (N_48615,N_47726,N_47759);
nand U48616 (N_48616,N_47872,N_47112);
nor U48617 (N_48617,N_47996,N_47746);
nor U48618 (N_48618,N_47518,N_47778);
or U48619 (N_48619,N_47444,N_47330);
nor U48620 (N_48620,N_47155,N_47110);
xor U48621 (N_48621,N_47622,N_47987);
or U48622 (N_48622,N_47868,N_47870);
and U48623 (N_48623,N_47746,N_47207);
nand U48624 (N_48624,N_47338,N_47269);
nand U48625 (N_48625,N_47095,N_47968);
and U48626 (N_48626,N_47893,N_47338);
nand U48627 (N_48627,N_47617,N_47920);
nor U48628 (N_48628,N_47663,N_47247);
xor U48629 (N_48629,N_47223,N_47286);
nor U48630 (N_48630,N_47666,N_47064);
or U48631 (N_48631,N_47352,N_47305);
or U48632 (N_48632,N_47658,N_47900);
or U48633 (N_48633,N_47335,N_47375);
nand U48634 (N_48634,N_47192,N_47022);
nor U48635 (N_48635,N_47074,N_47033);
nand U48636 (N_48636,N_47835,N_47393);
nor U48637 (N_48637,N_47345,N_47902);
or U48638 (N_48638,N_47069,N_47082);
nand U48639 (N_48639,N_47093,N_47017);
nor U48640 (N_48640,N_47331,N_47673);
nor U48641 (N_48641,N_47831,N_47696);
or U48642 (N_48642,N_47463,N_47974);
and U48643 (N_48643,N_47792,N_47891);
nand U48644 (N_48644,N_47760,N_47050);
or U48645 (N_48645,N_47121,N_47148);
and U48646 (N_48646,N_47320,N_47270);
nor U48647 (N_48647,N_47312,N_47468);
xnor U48648 (N_48648,N_47112,N_47475);
and U48649 (N_48649,N_47982,N_47970);
or U48650 (N_48650,N_47426,N_47519);
xor U48651 (N_48651,N_47360,N_47588);
nor U48652 (N_48652,N_47447,N_47038);
xor U48653 (N_48653,N_47201,N_47342);
or U48654 (N_48654,N_47734,N_47927);
or U48655 (N_48655,N_47652,N_47145);
or U48656 (N_48656,N_47570,N_47123);
nand U48657 (N_48657,N_47881,N_47768);
nand U48658 (N_48658,N_47145,N_47075);
and U48659 (N_48659,N_47167,N_47149);
or U48660 (N_48660,N_47742,N_47790);
xnor U48661 (N_48661,N_47428,N_47872);
xnor U48662 (N_48662,N_47563,N_47283);
and U48663 (N_48663,N_47627,N_47929);
or U48664 (N_48664,N_47340,N_47048);
xor U48665 (N_48665,N_47805,N_47786);
xor U48666 (N_48666,N_47237,N_47362);
nor U48667 (N_48667,N_47820,N_47658);
and U48668 (N_48668,N_47338,N_47195);
or U48669 (N_48669,N_47078,N_47499);
or U48670 (N_48670,N_47977,N_47458);
and U48671 (N_48671,N_47327,N_47172);
nor U48672 (N_48672,N_47110,N_47456);
xor U48673 (N_48673,N_47814,N_47522);
nor U48674 (N_48674,N_47465,N_47909);
xnor U48675 (N_48675,N_47465,N_47522);
nand U48676 (N_48676,N_47190,N_47058);
nand U48677 (N_48677,N_47168,N_47127);
or U48678 (N_48678,N_47817,N_47785);
or U48679 (N_48679,N_47784,N_47357);
nor U48680 (N_48680,N_47956,N_47732);
nand U48681 (N_48681,N_47171,N_47157);
nor U48682 (N_48682,N_47553,N_47504);
nor U48683 (N_48683,N_47213,N_47394);
and U48684 (N_48684,N_47961,N_47724);
or U48685 (N_48685,N_47840,N_47731);
xor U48686 (N_48686,N_47750,N_47617);
nand U48687 (N_48687,N_47059,N_47357);
and U48688 (N_48688,N_47306,N_47302);
xnor U48689 (N_48689,N_47439,N_47778);
or U48690 (N_48690,N_47844,N_47909);
nand U48691 (N_48691,N_47730,N_47713);
or U48692 (N_48692,N_47132,N_47255);
and U48693 (N_48693,N_47329,N_47921);
xor U48694 (N_48694,N_47294,N_47828);
and U48695 (N_48695,N_47220,N_47228);
xnor U48696 (N_48696,N_47864,N_47296);
nor U48697 (N_48697,N_47249,N_47365);
nand U48698 (N_48698,N_47027,N_47204);
nand U48699 (N_48699,N_47298,N_47575);
and U48700 (N_48700,N_47732,N_47794);
and U48701 (N_48701,N_47694,N_47720);
or U48702 (N_48702,N_47377,N_47426);
xnor U48703 (N_48703,N_47643,N_47279);
xor U48704 (N_48704,N_47933,N_47880);
xor U48705 (N_48705,N_47393,N_47042);
and U48706 (N_48706,N_47497,N_47396);
and U48707 (N_48707,N_47004,N_47086);
or U48708 (N_48708,N_47377,N_47924);
xor U48709 (N_48709,N_47144,N_47749);
xor U48710 (N_48710,N_47627,N_47301);
nor U48711 (N_48711,N_47052,N_47267);
nand U48712 (N_48712,N_47916,N_47938);
nor U48713 (N_48713,N_47564,N_47900);
and U48714 (N_48714,N_47227,N_47549);
nand U48715 (N_48715,N_47631,N_47728);
nor U48716 (N_48716,N_47690,N_47419);
nand U48717 (N_48717,N_47394,N_47711);
nand U48718 (N_48718,N_47307,N_47830);
nor U48719 (N_48719,N_47882,N_47755);
nor U48720 (N_48720,N_47189,N_47381);
and U48721 (N_48721,N_47249,N_47604);
xor U48722 (N_48722,N_47805,N_47334);
nand U48723 (N_48723,N_47236,N_47916);
xor U48724 (N_48724,N_47740,N_47571);
xnor U48725 (N_48725,N_47740,N_47395);
or U48726 (N_48726,N_47082,N_47639);
nor U48727 (N_48727,N_47394,N_47866);
and U48728 (N_48728,N_47732,N_47331);
and U48729 (N_48729,N_47418,N_47147);
xnor U48730 (N_48730,N_47570,N_47626);
and U48731 (N_48731,N_47894,N_47189);
and U48732 (N_48732,N_47768,N_47593);
or U48733 (N_48733,N_47765,N_47399);
nand U48734 (N_48734,N_47752,N_47342);
nand U48735 (N_48735,N_47981,N_47448);
nor U48736 (N_48736,N_47300,N_47294);
xnor U48737 (N_48737,N_47489,N_47306);
and U48738 (N_48738,N_47226,N_47278);
and U48739 (N_48739,N_47613,N_47477);
and U48740 (N_48740,N_47159,N_47470);
nor U48741 (N_48741,N_47070,N_47321);
and U48742 (N_48742,N_47275,N_47664);
or U48743 (N_48743,N_47346,N_47019);
and U48744 (N_48744,N_47700,N_47038);
xnor U48745 (N_48745,N_47955,N_47266);
and U48746 (N_48746,N_47225,N_47558);
or U48747 (N_48747,N_47011,N_47735);
nand U48748 (N_48748,N_47021,N_47225);
xor U48749 (N_48749,N_47840,N_47118);
xor U48750 (N_48750,N_47582,N_47204);
xnor U48751 (N_48751,N_47510,N_47049);
and U48752 (N_48752,N_47080,N_47445);
and U48753 (N_48753,N_47792,N_47137);
nand U48754 (N_48754,N_47972,N_47759);
or U48755 (N_48755,N_47261,N_47334);
nand U48756 (N_48756,N_47055,N_47425);
nor U48757 (N_48757,N_47103,N_47797);
or U48758 (N_48758,N_47536,N_47341);
nand U48759 (N_48759,N_47552,N_47537);
nor U48760 (N_48760,N_47129,N_47877);
or U48761 (N_48761,N_47145,N_47859);
nor U48762 (N_48762,N_47598,N_47199);
nand U48763 (N_48763,N_47356,N_47809);
or U48764 (N_48764,N_47527,N_47044);
or U48765 (N_48765,N_47512,N_47440);
and U48766 (N_48766,N_47837,N_47128);
nand U48767 (N_48767,N_47475,N_47027);
and U48768 (N_48768,N_47046,N_47690);
xor U48769 (N_48769,N_47506,N_47220);
xor U48770 (N_48770,N_47522,N_47354);
nand U48771 (N_48771,N_47403,N_47048);
nand U48772 (N_48772,N_47262,N_47114);
nor U48773 (N_48773,N_47433,N_47850);
and U48774 (N_48774,N_47351,N_47234);
xor U48775 (N_48775,N_47913,N_47853);
or U48776 (N_48776,N_47992,N_47695);
nor U48777 (N_48777,N_47988,N_47400);
nor U48778 (N_48778,N_47985,N_47348);
nor U48779 (N_48779,N_47570,N_47488);
nand U48780 (N_48780,N_47998,N_47062);
or U48781 (N_48781,N_47444,N_47882);
nand U48782 (N_48782,N_47498,N_47536);
xnor U48783 (N_48783,N_47373,N_47733);
or U48784 (N_48784,N_47870,N_47413);
and U48785 (N_48785,N_47882,N_47333);
and U48786 (N_48786,N_47520,N_47680);
and U48787 (N_48787,N_47470,N_47016);
xor U48788 (N_48788,N_47718,N_47595);
nand U48789 (N_48789,N_47984,N_47003);
and U48790 (N_48790,N_47482,N_47095);
nor U48791 (N_48791,N_47440,N_47488);
xor U48792 (N_48792,N_47382,N_47821);
nand U48793 (N_48793,N_47236,N_47261);
nand U48794 (N_48794,N_47357,N_47029);
or U48795 (N_48795,N_47162,N_47964);
xor U48796 (N_48796,N_47282,N_47320);
and U48797 (N_48797,N_47802,N_47041);
or U48798 (N_48798,N_47702,N_47367);
xor U48799 (N_48799,N_47293,N_47426);
xnor U48800 (N_48800,N_47061,N_47900);
xnor U48801 (N_48801,N_47043,N_47704);
nor U48802 (N_48802,N_47326,N_47146);
nand U48803 (N_48803,N_47420,N_47069);
nor U48804 (N_48804,N_47169,N_47423);
or U48805 (N_48805,N_47586,N_47293);
nand U48806 (N_48806,N_47148,N_47115);
and U48807 (N_48807,N_47421,N_47467);
nand U48808 (N_48808,N_47607,N_47548);
nor U48809 (N_48809,N_47048,N_47448);
or U48810 (N_48810,N_47294,N_47526);
and U48811 (N_48811,N_47520,N_47800);
nand U48812 (N_48812,N_47131,N_47610);
xor U48813 (N_48813,N_47721,N_47414);
and U48814 (N_48814,N_47468,N_47863);
xnor U48815 (N_48815,N_47205,N_47907);
xnor U48816 (N_48816,N_47693,N_47815);
and U48817 (N_48817,N_47594,N_47445);
or U48818 (N_48818,N_47084,N_47606);
or U48819 (N_48819,N_47791,N_47026);
and U48820 (N_48820,N_47315,N_47400);
xnor U48821 (N_48821,N_47445,N_47075);
xnor U48822 (N_48822,N_47577,N_47404);
nor U48823 (N_48823,N_47338,N_47986);
and U48824 (N_48824,N_47170,N_47700);
nand U48825 (N_48825,N_47412,N_47161);
nor U48826 (N_48826,N_47853,N_47949);
nor U48827 (N_48827,N_47238,N_47018);
nor U48828 (N_48828,N_47847,N_47196);
xnor U48829 (N_48829,N_47938,N_47021);
or U48830 (N_48830,N_47127,N_47218);
xor U48831 (N_48831,N_47070,N_47275);
or U48832 (N_48832,N_47244,N_47130);
or U48833 (N_48833,N_47478,N_47592);
nand U48834 (N_48834,N_47892,N_47904);
or U48835 (N_48835,N_47714,N_47349);
or U48836 (N_48836,N_47496,N_47459);
and U48837 (N_48837,N_47895,N_47729);
nand U48838 (N_48838,N_47865,N_47237);
and U48839 (N_48839,N_47829,N_47284);
xor U48840 (N_48840,N_47754,N_47071);
or U48841 (N_48841,N_47946,N_47233);
xor U48842 (N_48842,N_47002,N_47581);
nand U48843 (N_48843,N_47827,N_47705);
or U48844 (N_48844,N_47428,N_47909);
and U48845 (N_48845,N_47723,N_47582);
or U48846 (N_48846,N_47040,N_47464);
and U48847 (N_48847,N_47894,N_47130);
or U48848 (N_48848,N_47319,N_47394);
xor U48849 (N_48849,N_47133,N_47459);
xnor U48850 (N_48850,N_47035,N_47544);
or U48851 (N_48851,N_47672,N_47787);
nand U48852 (N_48852,N_47523,N_47030);
xnor U48853 (N_48853,N_47863,N_47749);
nor U48854 (N_48854,N_47907,N_47581);
or U48855 (N_48855,N_47885,N_47985);
or U48856 (N_48856,N_47975,N_47236);
or U48857 (N_48857,N_47346,N_47341);
or U48858 (N_48858,N_47636,N_47607);
or U48859 (N_48859,N_47258,N_47337);
and U48860 (N_48860,N_47866,N_47522);
and U48861 (N_48861,N_47893,N_47234);
xnor U48862 (N_48862,N_47006,N_47430);
and U48863 (N_48863,N_47157,N_47947);
and U48864 (N_48864,N_47571,N_47226);
and U48865 (N_48865,N_47753,N_47129);
nor U48866 (N_48866,N_47908,N_47658);
nand U48867 (N_48867,N_47648,N_47541);
or U48868 (N_48868,N_47913,N_47784);
xor U48869 (N_48869,N_47610,N_47625);
and U48870 (N_48870,N_47453,N_47129);
nand U48871 (N_48871,N_47527,N_47163);
xnor U48872 (N_48872,N_47225,N_47934);
xor U48873 (N_48873,N_47255,N_47579);
or U48874 (N_48874,N_47185,N_47025);
xor U48875 (N_48875,N_47404,N_47497);
xor U48876 (N_48876,N_47849,N_47410);
nor U48877 (N_48877,N_47749,N_47454);
nand U48878 (N_48878,N_47755,N_47292);
or U48879 (N_48879,N_47101,N_47207);
or U48880 (N_48880,N_47748,N_47617);
and U48881 (N_48881,N_47171,N_47014);
and U48882 (N_48882,N_47621,N_47121);
xor U48883 (N_48883,N_47518,N_47621);
and U48884 (N_48884,N_47148,N_47108);
nand U48885 (N_48885,N_47726,N_47438);
xor U48886 (N_48886,N_47171,N_47013);
and U48887 (N_48887,N_47480,N_47725);
nor U48888 (N_48888,N_47532,N_47516);
nand U48889 (N_48889,N_47693,N_47502);
nor U48890 (N_48890,N_47158,N_47001);
xnor U48891 (N_48891,N_47348,N_47207);
nand U48892 (N_48892,N_47629,N_47103);
and U48893 (N_48893,N_47736,N_47209);
xor U48894 (N_48894,N_47996,N_47325);
nor U48895 (N_48895,N_47614,N_47732);
and U48896 (N_48896,N_47013,N_47012);
and U48897 (N_48897,N_47402,N_47860);
or U48898 (N_48898,N_47421,N_47540);
and U48899 (N_48899,N_47003,N_47031);
xor U48900 (N_48900,N_47165,N_47174);
xor U48901 (N_48901,N_47157,N_47680);
and U48902 (N_48902,N_47391,N_47401);
nand U48903 (N_48903,N_47076,N_47543);
nor U48904 (N_48904,N_47510,N_47819);
and U48905 (N_48905,N_47354,N_47557);
nand U48906 (N_48906,N_47082,N_47662);
nor U48907 (N_48907,N_47386,N_47910);
and U48908 (N_48908,N_47533,N_47986);
xor U48909 (N_48909,N_47485,N_47645);
xor U48910 (N_48910,N_47841,N_47659);
nor U48911 (N_48911,N_47960,N_47178);
and U48912 (N_48912,N_47177,N_47185);
nor U48913 (N_48913,N_47384,N_47611);
or U48914 (N_48914,N_47340,N_47453);
and U48915 (N_48915,N_47726,N_47974);
xnor U48916 (N_48916,N_47159,N_47739);
nand U48917 (N_48917,N_47074,N_47837);
nand U48918 (N_48918,N_47353,N_47037);
nor U48919 (N_48919,N_47433,N_47041);
nor U48920 (N_48920,N_47940,N_47132);
or U48921 (N_48921,N_47414,N_47565);
and U48922 (N_48922,N_47372,N_47463);
nor U48923 (N_48923,N_47101,N_47357);
or U48924 (N_48924,N_47133,N_47884);
or U48925 (N_48925,N_47038,N_47444);
nor U48926 (N_48926,N_47519,N_47389);
xnor U48927 (N_48927,N_47469,N_47706);
and U48928 (N_48928,N_47222,N_47830);
or U48929 (N_48929,N_47972,N_47543);
nor U48930 (N_48930,N_47545,N_47670);
nor U48931 (N_48931,N_47057,N_47718);
or U48932 (N_48932,N_47413,N_47772);
xor U48933 (N_48933,N_47377,N_47099);
nand U48934 (N_48934,N_47730,N_47646);
or U48935 (N_48935,N_47500,N_47550);
and U48936 (N_48936,N_47000,N_47776);
xnor U48937 (N_48937,N_47377,N_47298);
nand U48938 (N_48938,N_47701,N_47339);
or U48939 (N_48939,N_47058,N_47115);
and U48940 (N_48940,N_47884,N_47658);
and U48941 (N_48941,N_47342,N_47954);
and U48942 (N_48942,N_47557,N_47285);
nand U48943 (N_48943,N_47359,N_47065);
and U48944 (N_48944,N_47179,N_47119);
and U48945 (N_48945,N_47228,N_47047);
and U48946 (N_48946,N_47686,N_47767);
or U48947 (N_48947,N_47601,N_47614);
nor U48948 (N_48948,N_47963,N_47744);
nand U48949 (N_48949,N_47447,N_47650);
nor U48950 (N_48950,N_47889,N_47712);
or U48951 (N_48951,N_47941,N_47888);
nand U48952 (N_48952,N_47997,N_47186);
or U48953 (N_48953,N_47403,N_47472);
or U48954 (N_48954,N_47856,N_47911);
nor U48955 (N_48955,N_47293,N_47896);
xor U48956 (N_48956,N_47088,N_47408);
xnor U48957 (N_48957,N_47007,N_47329);
or U48958 (N_48958,N_47276,N_47722);
nand U48959 (N_48959,N_47811,N_47304);
nand U48960 (N_48960,N_47784,N_47345);
or U48961 (N_48961,N_47115,N_47880);
nand U48962 (N_48962,N_47830,N_47562);
and U48963 (N_48963,N_47083,N_47577);
or U48964 (N_48964,N_47729,N_47854);
and U48965 (N_48965,N_47370,N_47111);
xnor U48966 (N_48966,N_47942,N_47683);
nor U48967 (N_48967,N_47564,N_47312);
and U48968 (N_48968,N_47275,N_47926);
or U48969 (N_48969,N_47508,N_47700);
nand U48970 (N_48970,N_47663,N_47457);
and U48971 (N_48971,N_47550,N_47109);
and U48972 (N_48972,N_47804,N_47270);
nand U48973 (N_48973,N_47488,N_47131);
nor U48974 (N_48974,N_47689,N_47217);
or U48975 (N_48975,N_47682,N_47068);
and U48976 (N_48976,N_47623,N_47635);
nor U48977 (N_48977,N_47120,N_47602);
and U48978 (N_48978,N_47245,N_47413);
nand U48979 (N_48979,N_47900,N_47321);
nand U48980 (N_48980,N_47189,N_47056);
and U48981 (N_48981,N_47439,N_47000);
xnor U48982 (N_48982,N_47328,N_47338);
and U48983 (N_48983,N_47502,N_47300);
nand U48984 (N_48984,N_47930,N_47045);
and U48985 (N_48985,N_47344,N_47952);
and U48986 (N_48986,N_47277,N_47511);
xnor U48987 (N_48987,N_47036,N_47025);
xor U48988 (N_48988,N_47835,N_47200);
or U48989 (N_48989,N_47569,N_47250);
nand U48990 (N_48990,N_47361,N_47358);
xnor U48991 (N_48991,N_47893,N_47165);
xor U48992 (N_48992,N_47893,N_47230);
nand U48993 (N_48993,N_47655,N_47837);
nor U48994 (N_48994,N_47015,N_47617);
or U48995 (N_48995,N_47024,N_47568);
nand U48996 (N_48996,N_47925,N_47999);
xor U48997 (N_48997,N_47124,N_47574);
nor U48998 (N_48998,N_47654,N_47765);
xnor U48999 (N_48999,N_47938,N_47258);
or U49000 (N_49000,N_48941,N_48855);
nor U49001 (N_49001,N_48524,N_48622);
or U49002 (N_49002,N_48812,N_48271);
xor U49003 (N_49003,N_48245,N_48918);
nand U49004 (N_49004,N_48935,N_48386);
or U49005 (N_49005,N_48669,N_48710);
xor U49006 (N_49006,N_48639,N_48649);
and U49007 (N_49007,N_48690,N_48410);
nand U49008 (N_49008,N_48411,N_48704);
and U49009 (N_49009,N_48845,N_48232);
nand U49010 (N_49010,N_48928,N_48937);
xnor U49011 (N_49011,N_48351,N_48580);
or U49012 (N_49012,N_48289,N_48511);
and U49013 (N_49013,N_48480,N_48692);
nor U49014 (N_49014,N_48507,N_48071);
or U49015 (N_49015,N_48777,N_48129);
nor U49016 (N_49016,N_48005,N_48431);
nand U49017 (N_49017,N_48343,N_48719);
xnor U49018 (N_49018,N_48416,N_48050);
or U49019 (N_49019,N_48378,N_48568);
or U49020 (N_49020,N_48577,N_48659);
and U49021 (N_49021,N_48617,N_48678);
xor U49022 (N_49022,N_48303,N_48977);
nor U49023 (N_49023,N_48728,N_48015);
nor U49024 (N_49024,N_48479,N_48801);
and U49025 (N_49025,N_48607,N_48342);
xor U49026 (N_49026,N_48832,N_48175);
or U49027 (N_49027,N_48395,N_48672);
nor U49028 (N_49028,N_48074,N_48909);
nor U49029 (N_49029,N_48557,N_48247);
and U49030 (N_49030,N_48775,N_48367);
xor U49031 (N_49031,N_48644,N_48520);
xor U49032 (N_49032,N_48993,N_48985);
nand U49033 (N_49033,N_48847,N_48003);
or U49034 (N_49034,N_48357,N_48699);
nor U49035 (N_49035,N_48171,N_48798);
and U49036 (N_49036,N_48809,N_48348);
or U49037 (N_49037,N_48179,N_48078);
or U49038 (N_49038,N_48926,N_48360);
and U49039 (N_49039,N_48760,N_48340);
and U49040 (N_49040,N_48194,N_48666);
or U49041 (N_49041,N_48685,N_48133);
nor U49042 (N_49042,N_48455,N_48654);
and U49043 (N_49043,N_48599,N_48069);
nor U49044 (N_49044,N_48353,N_48093);
or U49045 (N_49045,N_48060,N_48402);
or U49046 (N_49046,N_48804,N_48439);
and U49047 (N_49047,N_48796,N_48778);
or U49048 (N_49048,N_48998,N_48330);
xnor U49049 (N_49049,N_48092,N_48125);
nand U49050 (N_49050,N_48508,N_48035);
nand U49051 (N_49051,N_48814,N_48504);
nor U49052 (N_49052,N_48304,N_48542);
or U49053 (N_49053,N_48314,N_48493);
and U49054 (N_49054,N_48359,N_48682);
nand U49055 (N_49055,N_48588,N_48866);
xnor U49056 (N_49056,N_48356,N_48612);
or U49057 (N_49057,N_48382,N_48581);
nand U49058 (N_49058,N_48959,N_48296);
nand U49059 (N_49059,N_48829,N_48602);
nor U49060 (N_49060,N_48957,N_48295);
nand U49061 (N_49061,N_48198,N_48141);
nand U49062 (N_49062,N_48980,N_48625);
or U49063 (N_49063,N_48843,N_48252);
and U49064 (N_49064,N_48932,N_48226);
and U49065 (N_49065,N_48254,N_48558);
or U49066 (N_49066,N_48893,N_48009);
nor U49067 (N_49067,N_48502,N_48063);
xnor U49068 (N_49068,N_48265,N_48564);
and U49069 (N_49069,N_48266,N_48865);
nand U49070 (N_49070,N_48901,N_48967);
xor U49071 (N_49071,N_48503,N_48774);
and U49072 (N_49072,N_48280,N_48551);
or U49073 (N_49073,N_48754,N_48421);
and U49074 (N_49074,N_48700,N_48428);
nor U49075 (N_49075,N_48461,N_48905);
xor U49076 (N_49076,N_48067,N_48910);
nand U49077 (N_49077,N_48301,N_48867);
nor U49078 (N_49078,N_48243,N_48627);
and U49079 (N_49079,N_48756,N_48995);
nand U49080 (N_49080,N_48338,N_48684);
xor U49081 (N_49081,N_48495,N_48800);
nor U49082 (N_49082,N_48374,N_48570);
nor U49083 (N_49083,N_48651,N_48675);
and U49084 (N_49084,N_48033,N_48234);
or U49085 (N_49085,N_48540,N_48268);
xor U49086 (N_49086,N_48592,N_48730);
nor U49087 (N_49087,N_48380,N_48201);
nor U49088 (N_49088,N_48242,N_48115);
or U49089 (N_49089,N_48769,N_48586);
and U49090 (N_49090,N_48354,N_48709);
or U49091 (N_49091,N_48992,N_48022);
nor U49092 (N_49092,N_48341,N_48991);
nor U49093 (N_49093,N_48292,N_48116);
nor U49094 (N_49094,N_48598,N_48166);
and U49095 (N_49095,N_48165,N_48827);
xor U49096 (N_49096,N_48447,N_48954);
or U49097 (N_49097,N_48857,N_48702);
and U49098 (N_49098,N_48097,N_48594);
nor U49099 (N_49099,N_48648,N_48290);
and U49100 (N_49100,N_48489,N_48002);
xnor U49101 (N_49101,N_48745,N_48830);
xnor U49102 (N_49102,N_48294,N_48876);
or U49103 (N_49103,N_48652,N_48427);
and U49104 (N_49104,N_48211,N_48562);
or U49105 (N_49105,N_48291,N_48048);
nand U49106 (N_49106,N_48761,N_48531);
and U49107 (N_49107,N_48687,N_48922);
xor U49108 (N_49108,N_48573,N_48988);
and U49109 (N_49109,N_48929,N_48544);
and U49110 (N_49110,N_48436,N_48975);
nor U49111 (N_49111,N_48401,N_48476);
nand U49112 (N_49112,N_48267,N_48256);
and U49113 (N_49113,N_48442,N_48080);
and U49114 (N_49114,N_48720,N_48591);
nor U49115 (N_49115,N_48786,N_48638);
nand U49116 (N_49116,N_48131,N_48117);
nand U49117 (N_49117,N_48323,N_48239);
and U49118 (N_49118,N_48384,N_48039);
nand U49119 (N_49119,N_48123,N_48169);
nor U49120 (N_49120,N_48947,N_48898);
nor U49121 (N_49121,N_48757,N_48258);
xnor U49122 (N_49122,N_48075,N_48674);
nand U49123 (N_49123,N_48608,N_48197);
nor U49124 (N_49124,N_48433,N_48499);
xor U49125 (N_49125,N_48471,N_48013);
nand U49126 (N_49126,N_48152,N_48882);
and U49127 (N_49127,N_48478,N_48144);
and U49128 (N_49128,N_48936,N_48206);
and U49129 (N_49129,N_48514,N_48065);
and U49130 (N_49130,N_48787,N_48895);
nor U49131 (N_49131,N_48244,N_48713);
or U49132 (N_49132,N_48210,N_48269);
xnor U49133 (N_49133,N_48309,N_48135);
and U49134 (N_49134,N_48264,N_48460);
and U49135 (N_49135,N_48387,N_48057);
xnor U49136 (N_49136,N_48438,N_48474);
xor U49137 (N_49137,N_48597,N_48444);
nor U49138 (N_49138,N_48885,N_48191);
nand U49139 (N_49139,N_48541,N_48956);
nor U49140 (N_49140,N_48276,N_48224);
xor U49141 (N_49141,N_48925,N_48731);
nor U49142 (N_49142,N_48958,N_48413);
or U49143 (N_49143,N_48660,N_48714);
xor U49144 (N_49144,N_48192,N_48556);
and U49145 (N_49145,N_48846,N_48613);
or U49146 (N_49146,N_48664,N_48740);
nand U49147 (N_49147,N_48099,N_48579);
nand U49148 (N_49148,N_48062,N_48717);
xnor U49149 (N_49149,N_48465,N_48743);
and U49150 (N_49150,N_48076,N_48393);
xor U49151 (N_49151,N_48528,N_48283);
and U49152 (N_49152,N_48631,N_48167);
xnor U49153 (N_49153,N_48213,N_48240);
nor U49154 (N_49154,N_48547,N_48772);
and U49155 (N_49155,N_48722,N_48320);
xnor U49156 (N_49156,N_48994,N_48082);
or U49157 (N_49157,N_48485,N_48420);
or U49158 (N_49158,N_48365,N_48228);
or U49159 (N_49159,N_48056,N_48459);
xnor U49160 (N_49160,N_48752,N_48792);
nor U49161 (N_49161,N_48180,N_48443);
nand U49162 (N_49162,N_48396,N_48931);
or U49163 (N_49163,N_48081,N_48263);
xor U49164 (N_49164,N_48456,N_48842);
nor U49165 (N_49165,N_48668,N_48146);
or U49166 (N_49166,N_48358,N_48202);
and U49167 (N_49167,N_48111,N_48369);
nor U49168 (N_49168,N_48043,N_48884);
or U49169 (N_49169,N_48878,N_48810);
xor U49170 (N_49170,N_48986,N_48151);
xnor U49171 (N_49171,N_48231,N_48744);
xnor U49172 (N_49172,N_48583,N_48864);
or U49173 (N_49173,N_48630,N_48571);
and U49174 (N_49174,N_48753,N_48596);
nor U49175 (N_49175,N_48697,N_48087);
nor U49176 (N_49176,N_48446,N_48698);
and U49177 (N_49177,N_48220,N_48188);
or U49178 (N_49178,N_48789,N_48559);
nor U49179 (N_49179,N_48399,N_48724);
and U49180 (N_49180,N_48324,N_48279);
and U49181 (N_49181,N_48694,N_48322);
and U49182 (N_49182,N_48046,N_48405);
or U49183 (N_49183,N_48620,N_48536);
xor U49184 (N_49184,N_48961,N_48712);
xor U49185 (N_49185,N_48634,N_48145);
and U49186 (N_49186,N_48124,N_48751);
and U49187 (N_49187,N_48575,N_48236);
and U49188 (N_49188,N_48275,N_48453);
nand U49189 (N_49189,N_48134,N_48705);
nand U49190 (N_49190,N_48066,N_48739);
and U49191 (N_49191,N_48737,N_48222);
or U49192 (N_49192,N_48091,N_48372);
nor U49193 (N_49193,N_48229,N_48887);
xnor U49194 (N_49194,N_48112,N_48762);
or U49195 (N_49195,N_48758,N_48020);
nand U49196 (N_49196,N_48333,N_48390);
or U49197 (N_49197,N_48138,N_48516);
nand U49198 (N_49198,N_48892,N_48451);
xnor U49199 (N_49199,N_48225,N_48526);
nor U49200 (N_49200,N_48635,N_48335);
nor U49201 (N_49201,N_48418,N_48938);
or U49202 (N_49202,N_48127,N_48679);
nand U49203 (N_49203,N_48477,N_48844);
or U49204 (N_49204,N_48982,N_48429);
xor U49205 (N_49205,N_48137,N_48454);
and U49206 (N_49206,N_48053,N_48595);
nand U49207 (N_49207,N_48587,N_48629);
and U49208 (N_49208,N_48107,N_48006);
nand U49209 (N_49209,N_48227,N_48337);
nand U49210 (N_49210,N_48084,N_48363);
or U49211 (N_49211,N_48951,N_48400);
xnor U49212 (N_49212,N_48773,N_48949);
nand U49213 (N_49213,N_48911,N_48072);
nor U49214 (N_49214,N_48077,N_48223);
nor U49215 (N_49215,N_48339,N_48716);
or U49216 (N_49216,N_48207,N_48718);
and U49217 (N_49217,N_48848,N_48912);
or U49218 (N_49218,N_48734,N_48904);
and U49219 (N_49219,N_48469,N_48199);
or U49220 (N_49220,N_48921,N_48549);
or U49221 (N_49221,N_48394,N_48726);
nor U49222 (N_49222,N_48492,N_48965);
and U49223 (N_49223,N_48670,N_48661);
xnor U49224 (N_49224,N_48894,N_48034);
and U49225 (N_49225,N_48457,N_48632);
and U49226 (N_49226,N_48671,N_48767);
and U49227 (N_49227,N_48611,N_48621);
xor U49228 (N_49228,N_48344,N_48979);
nor U49229 (N_49229,N_48467,N_48868);
or U49230 (N_49230,N_48852,N_48715);
and U49231 (N_49231,N_48486,N_48328);
and U49232 (N_49232,N_48253,N_48512);
nor U49233 (N_49233,N_48491,N_48601);
nand U49234 (N_49234,N_48021,N_48934);
xor U49235 (N_49235,N_48248,N_48302);
and U49236 (N_49236,N_48791,N_48689);
nand U49237 (N_49237,N_48037,N_48004);
and U49238 (N_49238,N_48858,N_48425);
nand U49239 (N_49239,N_48923,N_48184);
or U49240 (N_49240,N_48011,N_48623);
or U49241 (N_49241,N_48680,N_48768);
xnor U49242 (N_49242,N_48889,N_48437);
xnor U49243 (N_49243,N_48837,N_48899);
or U49244 (N_49244,N_48535,N_48217);
nor U49245 (N_49245,N_48733,N_48933);
xnor U49246 (N_49246,N_48582,N_48440);
xnor U49247 (N_49247,N_48441,N_48120);
xnor U49248 (N_49248,N_48423,N_48041);
xor U49249 (N_49249,N_48628,N_48736);
or U49250 (N_49250,N_48150,N_48040);
nand U49251 (N_49251,N_48347,N_48797);
nand U49252 (N_49252,N_48870,N_48162);
xor U49253 (N_49253,N_48088,N_48793);
or U49254 (N_49254,N_48070,N_48808);
xnor U49255 (N_49255,N_48908,N_48838);
nor U49256 (N_49256,N_48001,N_48505);
nand U49257 (N_49257,N_48497,N_48155);
nand U49258 (N_49258,N_48103,N_48158);
nor U49259 (N_49259,N_48388,N_48249);
xor U49260 (N_49260,N_48110,N_48560);
xnor U49261 (N_49261,N_48874,N_48350);
nand U49262 (N_49262,N_48398,N_48316);
or U49263 (N_49263,N_48108,N_48946);
or U49264 (N_49264,N_48185,N_48119);
xor U49265 (N_49265,N_48822,N_48310);
xor U49266 (N_49266,N_48696,N_48605);
and U49267 (N_49267,N_48308,N_48723);
nand U49268 (N_49268,N_48813,N_48686);
and U49269 (N_49269,N_48259,N_48101);
nand U49270 (N_49270,N_48907,N_48945);
xor U49271 (N_49271,N_48422,N_48010);
xnor U49272 (N_49272,N_48329,N_48098);
nor U49273 (N_49273,N_48089,N_48695);
or U49274 (N_49274,N_48811,N_48250);
or U49275 (N_49275,N_48881,N_48193);
xnor U49276 (N_49276,N_48000,N_48312);
xor U49277 (N_49277,N_48260,N_48869);
or U49278 (N_49278,N_48803,N_48321);
xnor U49279 (N_49279,N_48325,N_48548);
nor U49280 (N_49280,N_48653,N_48045);
xnor U49281 (N_49281,N_48955,N_48313);
nor U49282 (N_49282,N_48780,N_48770);
or U49283 (N_49283,N_48424,N_48142);
nor U49284 (N_49284,N_48470,N_48068);
or U49285 (N_49285,N_48539,N_48136);
and U49286 (N_49286,N_48408,N_48732);
nand U49287 (N_49287,N_48619,N_48121);
xnor U49288 (N_49288,N_48532,N_48017);
or U49289 (N_49289,N_48430,N_48606);
and U49290 (N_49290,N_48272,N_48159);
and U49291 (N_49291,N_48100,N_48873);
or U49292 (N_49292,N_48759,N_48805);
nor U49293 (N_49293,N_48029,N_48783);
nand U49294 (N_49294,N_48462,N_48891);
nor U49295 (N_49295,N_48102,N_48984);
nor U49296 (N_49296,N_48545,N_48799);
nand U49297 (N_49297,N_48174,N_48538);
and U49298 (N_49298,N_48331,N_48235);
xor U49299 (N_49299,N_48779,N_48498);
and U49300 (N_49300,N_48214,N_48044);
and U49301 (N_49301,N_48854,N_48432);
or U49302 (N_49302,N_48833,N_48915);
xor U49303 (N_49303,N_48600,N_48172);
and U49304 (N_49304,N_48434,N_48795);
xnor U49305 (N_49305,N_48880,N_48153);
and U49306 (N_49306,N_48083,N_48389);
or U49307 (N_49307,N_48860,N_48297);
and U49308 (N_49308,N_48412,N_48435);
nand U49309 (N_49309,N_48525,N_48018);
and U49310 (N_49310,N_48543,N_48897);
nand U49311 (N_49311,N_48284,N_48807);
and U49312 (N_49312,N_48989,N_48128);
nor U49313 (N_49313,N_48472,N_48085);
xor U49314 (N_49314,N_48515,N_48187);
and U49315 (N_49315,N_48130,N_48825);
or U49316 (N_49316,N_48618,N_48537);
nand U49317 (N_49317,N_48725,N_48708);
nand U49318 (N_49318,N_48007,N_48319);
nor U49319 (N_49319,N_48942,N_48997);
and U49320 (N_49320,N_48332,N_48143);
nor U49321 (N_49321,N_48445,N_48764);
or U49322 (N_49322,N_48299,N_48305);
nor U49323 (N_49323,N_48482,N_48836);
or U49324 (N_49324,N_48626,N_48765);
or U49325 (N_49325,N_48534,N_48823);
xor U49326 (N_49326,N_48966,N_48721);
nor U49327 (N_49327,N_48841,N_48746);
or U49328 (N_49328,N_48940,N_48230);
xnor U49329 (N_49329,N_48640,N_48061);
or U49330 (N_49330,N_48375,N_48939);
nor U49331 (N_49331,N_48978,N_48533);
and U49332 (N_49332,N_48204,N_48452);
or U49333 (N_49333,N_48327,N_48964);
or U49334 (N_49334,N_48963,N_48968);
or U49335 (N_49335,N_48181,N_48785);
or U49336 (N_49336,N_48913,N_48806);
xor U49337 (N_49337,N_48662,N_48590);
or U49338 (N_49338,N_48593,N_48711);
or U49339 (N_49339,N_48409,N_48106);
xor U49340 (N_49340,N_48962,N_48530);
xnor U49341 (N_49341,N_48983,N_48552);
and U49342 (N_49342,N_48036,N_48856);
or U49343 (N_49343,N_48886,N_48168);
and U49344 (N_49344,N_48771,N_48032);
or U49345 (N_49345,N_48277,N_48379);
nor U49346 (N_49346,N_48794,N_48016);
xnor U49347 (N_49347,N_48377,N_48049);
and U49348 (N_49348,N_48219,N_48604);
nand U49349 (N_49349,N_48614,N_48449);
nand U49350 (N_49350,N_48561,N_48642);
nand U49351 (N_49351,N_48368,N_48285);
nor U49352 (N_49352,N_48113,N_48944);
xor U49353 (N_49353,N_48090,N_48521);
or U49354 (N_49354,N_48902,N_48496);
and U49355 (N_49355,N_48750,N_48815);
nand U49356 (N_49356,N_48487,N_48987);
nand U49357 (N_49357,N_48518,N_48209);
nor U49358 (N_49358,N_48177,N_48972);
nor U49359 (N_49359,N_48336,N_48385);
or U49360 (N_49360,N_48318,N_48173);
or U49361 (N_49361,N_48615,N_48610);
nand U49362 (N_49362,N_48976,N_48567);
nor U49363 (N_49363,N_48414,N_48346);
nand U49364 (N_49364,N_48849,N_48157);
or U49365 (N_49365,N_48326,N_48999);
and U49366 (N_49366,N_48677,N_48246);
nand U49367 (N_49367,N_48840,N_48763);
nor U49368 (N_49368,N_48481,N_48555);
and U49369 (N_49369,N_48510,N_48052);
nor U49370 (N_49370,N_48834,N_48196);
or U49371 (N_49371,N_48650,N_48458);
nand U49372 (N_49372,N_48916,N_48371);
nor U49373 (N_49373,N_48450,N_48519);
or U49374 (N_49374,N_48546,N_48352);
nand U49375 (N_49375,N_48306,N_48943);
or U49376 (N_49376,N_48589,N_48051);
xor U49377 (N_49377,N_48633,N_48550);
nand U49378 (N_49378,N_48574,N_48397);
nor U49379 (N_49379,N_48208,N_48376);
and U49380 (N_49380,N_48156,N_48109);
nand U49381 (N_49381,N_48748,N_48563);
xnor U49382 (N_49382,N_48373,N_48673);
nand U49383 (N_49383,N_48784,N_48578);
or U49384 (N_49384,N_48883,N_48023);
and U49385 (N_49385,N_48417,N_48027);
xor U49386 (N_49386,N_48251,N_48257);
nor U49387 (N_49387,N_48233,N_48270);
nand U49388 (N_49388,N_48647,N_48665);
xor U49389 (N_49389,N_48079,N_48178);
or U49390 (N_49390,N_48426,N_48370);
or U49391 (N_49391,N_48790,N_48749);
nand U49392 (N_49392,N_48788,N_48237);
nand U49393 (N_49393,N_48362,N_48747);
nor U49394 (N_49394,N_48862,N_48676);
nand U49395 (N_49395,N_48114,N_48974);
and U49396 (N_49396,N_48616,N_48553);
xnor U49397 (N_49397,N_48042,N_48691);
nor U49398 (N_49398,N_48655,N_48960);
or U49399 (N_49399,N_48415,N_48667);
and U49400 (N_49400,N_48609,N_48293);
xor U49401 (N_49401,N_48569,N_48298);
and U49402 (N_49402,N_48490,N_48817);
nand U49403 (N_49403,N_48990,N_48139);
xor U49404 (N_49404,N_48215,N_48161);
or U49405 (N_49405,N_48973,N_48154);
nand U49406 (N_49406,N_48924,N_48658);
nand U49407 (N_49407,N_48241,N_48286);
xor U49408 (N_49408,N_48643,N_48906);
and U49409 (N_49409,N_48147,N_48930);
nand U49410 (N_49410,N_48028,N_48821);
or U49411 (N_49411,N_48996,N_48317);
nor U49412 (N_49412,N_48288,N_48073);
xnor U49413 (N_49413,N_48527,N_48058);
xor U49414 (N_49414,N_48900,N_48483);
nand U49415 (N_49415,N_48872,N_48917);
or U49416 (N_49416,N_48488,N_48261);
nand U49417 (N_49417,N_48701,N_48688);
or U49418 (N_49418,N_48681,N_48952);
nor U49419 (N_49419,N_48448,N_48646);
nand U49420 (N_49420,N_48981,N_48850);
nor U49421 (N_49421,N_48030,N_48703);
nor U49422 (N_49422,N_48741,N_48182);
nand U49423 (N_49423,N_48118,N_48064);
nor U49424 (N_49424,N_48802,N_48566);
nand U49425 (N_49425,N_48255,N_48024);
or U49426 (N_49426,N_48645,N_48683);
and U49427 (N_49427,N_48624,N_48054);
xor U49428 (N_49428,N_48176,N_48274);
and U49429 (N_49429,N_48839,N_48506);
and U49430 (N_49430,N_48663,N_48729);
nor U49431 (N_49431,N_48554,N_48950);
nor U49432 (N_49432,N_48104,N_48927);
or U49433 (N_49433,N_48742,N_48896);
nand U49434 (N_49434,N_48565,N_48781);
nand U49435 (N_49435,N_48381,N_48148);
nor U49436 (N_49436,N_48953,N_48766);
and U49437 (N_49437,N_48170,N_48183);
and U49438 (N_49438,N_48278,N_48826);
nor U49439 (N_49439,N_48853,N_48513);
and U49440 (N_49440,N_48824,N_48464);
or U49441 (N_49441,N_48888,N_48473);
and U49442 (N_49442,N_48149,N_48205);
nor U49443 (N_49443,N_48391,N_48273);
xor U49444 (N_49444,N_48238,N_48383);
or U49445 (N_49445,N_48816,N_48025);
nand U49446 (N_49446,N_48831,N_48311);
and U49447 (N_49447,N_48404,N_48871);
xnor U49448 (N_49448,N_48221,N_48186);
or U49449 (N_49449,N_48105,N_48637);
or U49450 (N_49450,N_48727,N_48877);
xnor U49451 (N_49451,N_48509,N_48484);
nand U49452 (N_49452,N_48095,N_48392);
xnor U49453 (N_49453,N_48307,N_48861);
xnor U49454 (N_49454,N_48190,N_48517);
nand U49455 (N_49455,N_48576,N_48863);
and U49456 (N_49456,N_48879,N_48407);
and U49457 (N_49457,N_48160,N_48755);
and U49458 (N_49458,N_48735,N_48406);
nand U49459 (N_49459,N_48026,N_48287);
nor U49460 (N_49460,N_48820,N_48463);
nand U49461 (N_49461,N_48361,N_48163);
and U49462 (N_49462,N_48212,N_48585);
and U49463 (N_49463,N_48315,N_48970);
and U49464 (N_49464,N_48403,N_48776);
or U49465 (N_49465,N_48059,N_48875);
nand U49466 (N_49466,N_48468,N_48008);
or U49467 (N_49467,N_48216,N_48890);
xor U49468 (N_49468,N_48707,N_48366);
or U49469 (N_49469,N_48218,N_48055);
or U49470 (N_49470,N_48038,N_48047);
or U49471 (N_49471,N_48195,N_48086);
or U49472 (N_49472,N_48818,N_48282);
nand U49473 (N_49473,N_48919,N_48693);
nor U49474 (N_49474,N_48364,N_48706);
or U49475 (N_49475,N_48969,N_48782);
and U49476 (N_49476,N_48122,N_48522);
nand U49477 (N_49477,N_48019,N_48657);
xor U49478 (N_49478,N_48971,N_48920);
nor U49479 (N_49479,N_48851,N_48132);
nand U49480 (N_49480,N_48014,N_48096);
nor U49481 (N_49481,N_48475,N_48012);
and U49482 (N_49482,N_48641,N_48164);
xnor U49483 (N_49483,N_48914,N_48345);
nand U49484 (N_49484,N_48334,N_48529);
and U49485 (N_49485,N_48189,N_48094);
xor U49486 (N_49486,N_48603,N_48523);
and U49487 (N_49487,N_48466,N_48828);
nand U49488 (N_49488,N_48738,N_48948);
xor U49489 (N_49489,N_48656,N_48419);
nor U49490 (N_49490,N_48819,N_48835);
and U49491 (N_49491,N_48859,N_48262);
or U49492 (N_49492,N_48355,N_48126);
and U49493 (N_49493,N_48203,N_48494);
nor U49494 (N_49494,N_48300,N_48636);
and U49495 (N_49495,N_48572,N_48031);
nor U49496 (N_49496,N_48903,N_48349);
nand U49497 (N_49497,N_48140,N_48501);
xor U49498 (N_49498,N_48281,N_48500);
or U49499 (N_49499,N_48584,N_48200);
nand U49500 (N_49500,N_48088,N_48126);
or U49501 (N_49501,N_48453,N_48666);
or U49502 (N_49502,N_48774,N_48317);
nor U49503 (N_49503,N_48080,N_48598);
nor U49504 (N_49504,N_48431,N_48501);
or U49505 (N_49505,N_48342,N_48609);
or U49506 (N_49506,N_48582,N_48390);
nor U49507 (N_49507,N_48132,N_48642);
nand U49508 (N_49508,N_48080,N_48949);
xor U49509 (N_49509,N_48846,N_48633);
nand U49510 (N_49510,N_48441,N_48882);
nand U49511 (N_49511,N_48686,N_48146);
nor U49512 (N_49512,N_48042,N_48372);
or U49513 (N_49513,N_48860,N_48671);
or U49514 (N_49514,N_48330,N_48678);
xnor U49515 (N_49515,N_48690,N_48898);
and U49516 (N_49516,N_48644,N_48634);
nor U49517 (N_49517,N_48063,N_48048);
xnor U49518 (N_49518,N_48722,N_48020);
or U49519 (N_49519,N_48677,N_48214);
nor U49520 (N_49520,N_48643,N_48540);
xor U49521 (N_49521,N_48639,N_48080);
nor U49522 (N_49522,N_48869,N_48067);
or U49523 (N_49523,N_48178,N_48453);
nor U49524 (N_49524,N_48238,N_48731);
and U49525 (N_49525,N_48035,N_48077);
and U49526 (N_49526,N_48343,N_48770);
nand U49527 (N_49527,N_48152,N_48224);
xnor U49528 (N_49528,N_48227,N_48438);
and U49529 (N_49529,N_48869,N_48020);
nor U49530 (N_49530,N_48978,N_48562);
nor U49531 (N_49531,N_48591,N_48815);
nor U49532 (N_49532,N_48704,N_48627);
nor U49533 (N_49533,N_48109,N_48968);
nor U49534 (N_49534,N_48794,N_48966);
nor U49535 (N_49535,N_48704,N_48087);
and U49536 (N_49536,N_48362,N_48880);
xnor U49537 (N_49537,N_48402,N_48775);
nor U49538 (N_49538,N_48712,N_48227);
nor U49539 (N_49539,N_48099,N_48429);
xor U49540 (N_49540,N_48649,N_48611);
and U49541 (N_49541,N_48885,N_48322);
xnor U49542 (N_49542,N_48070,N_48706);
xnor U49543 (N_49543,N_48233,N_48105);
nor U49544 (N_49544,N_48477,N_48355);
nor U49545 (N_49545,N_48771,N_48310);
nor U49546 (N_49546,N_48562,N_48663);
nor U49547 (N_49547,N_48321,N_48657);
nand U49548 (N_49548,N_48659,N_48911);
nor U49549 (N_49549,N_48081,N_48737);
or U49550 (N_49550,N_48940,N_48278);
xnor U49551 (N_49551,N_48918,N_48623);
and U49552 (N_49552,N_48762,N_48221);
and U49553 (N_49553,N_48642,N_48943);
xnor U49554 (N_49554,N_48376,N_48449);
nand U49555 (N_49555,N_48619,N_48535);
nand U49556 (N_49556,N_48790,N_48787);
nand U49557 (N_49557,N_48713,N_48504);
nand U49558 (N_49558,N_48331,N_48271);
or U49559 (N_49559,N_48303,N_48193);
xor U49560 (N_49560,N_48348,N_48319);
nor U49561 (N_49561,N_48507,N_48745);
nor U49562 (N_49562,N_48917,N_48044);
xor U49563 (N_49563,N_48817,N_48619);
or U49564 (N_49564,N_48652,N_48025);
and U49565 (N_49565,N_48107,N_48585);
nor U49566 (N_49566,N_48651,N_48807);
nor U49567 (N_49567,N_48714,N_48630);
nor U49568 (N_49568,N_48690,N_48849);
nor U49569 (N_49569,N_48812,N_48967);
or U49570 (N_49570,N_48746,N_48508);
or U49571 (N_49571,N_48537,N_48139);
xnor U49572 (N_49572,N_48935,N_48022);
xnor U49573 (N_49573,N_48583,N_48070);
nor U49574 (N_49574,N_48296,N_48277);
or U49575 (N_49575,N_48483,N_48669);
xnor U49576 (N_49576,N_48624,N_48136);
or U49577 (N_49577,N_48057,N_48190);
xnor U49578 (N_49578,N_48420,N_48718);
or U49579 (N_49579,N_48283,N_48228);
or U49580 (N_49580,N_48743,N_48563);
or U49581 (N_49581,N_48769,N_48416);
or U49582 (N_49582,N_48459,N_48356);
and U49583 (N_49583,N_48241,N_48926);
nor U49584 (N_49584,N_48665,N_48473);
nand U49585 (N_49585,N_48162,N_48422);
and U49586 (N_49586,N_48076,N_48985);
nand U49587 (N_49587,N_48825,N_48424);
nand U49588 (N_49588,N_48875,N_48590);
and U49589 (N_49589,N_48499,N_48014);
nor U49590 (N_49590,N_48042,N_48030);
or U49591 (N_49591,N_48449,N_48959);
xnor U49592 (N_49592,N_48424,N_48910);
nand U49593 (N_49593,N_48687,N_48433);
xor U49594 (N_49594,N_48587,N_48577);
nor U49595 (N_49595,N_48738,N_48511);
nand U49596 (N_49596,N_48969,N_48236);
and U49597 (N_49597,N_48001,N_48315);
or U49598 (N_49598,N_48358,N_48771);
nor U49599 (N_49599,N_48547,N_48490);
or U49600 (N_49600,N_48788,N_48877);
nand U49601 (N_49601,N_48874,N_48378);
xnor U49602 (N_49602,N_48116,N_48737);
or U49603 (N_49603,N_48756,N_48182);
and U49604 (N_49604,N_48580,N_48735);
and U49605 (N_49605,N_48964,N_48549);
nor U49606 (N_49606,N_48691,N_48110);
xor U49607 (N_49607,N_48008,N_48808);
nand U49608 (N_49608,N_48126,N_48157);
and U49609 (N_49609,N_48871,N_48092);
and U49610 (N_49610,N_48788,N_48201);
nand U49611 (N_49611,N_48938,N_48031);
and U49612 (N_49612,N_48014,N_48217);
nand U49613 (N_49613,N_48175,N_48614);
nor U49614 (N_49614,N_48346,N_48583);
xor U49615 (N_49615,N_48469,N_48254);
nand U49616 (N_49616,N_48575,N_48407);
or U49617 (N_49617,N_48207,N_48397);
or U49618 (N_49618,N_48683,N_48585);
xnor U49619 (N_49619,N_48839,N_48521);
xnor U49620 (N_49620,N_48433,N_48763);
or U49621 (N_49621,N_48163,N_48776);
and U49622 (N_49622,N_48021,N_48231);
nor U49623 (N_49623,N_48285,N_48554);
nor U49624 (N_49624,N_48488,N_48203);
xnor U49625 (N_49625,N_48212,N_48001);
nand U49626 (N_49626,N_48759,N_48274);
xor U49627 (N_49627,N_48023,N_48479);
nand U49628 (N_49628,N_48931,N_48407);
nand U49629 (N_49629,N_48513,N_48528);
and U49630 (N_49630,N_48722,N_48544);
nor U49631 (N_49631,N_48154,N_48576);
or U49632 (N_49632,N_48627,N_48960);
nor U49633 (N_49633,N_48722,N_48936);
xor U49634 (N_49634,N_48819,N_48533);
and U49635 (N_49635,N_48150,N_48015);
nand U49636 (N_49636,N_48214,N_48168);
or U49637 (N_49637,N_48711,N_48032);
and U49638 (N_49638,N_48006,N_48901);
nand U49639 (N_49639,N_48386,N_48002);
xor U49640 (N_49640,N_48898,N_48528);
xor U49641 (N_49641,N_48810,N_48307);
nand U49642 (N_49642,N_48461,N_48183);
and U49643 (N_49643,N_48813,N_48605);
and U49644 (N_49644,N_48577,N_48650);
nand U49645 (N_49645,N_48826,N_48612);
nor U49646 (N_49646,N_48164,N_48165);
nor U49647 (N_49647,N_48197,N_48026);
nand U49648 (N_49648,N_48824,N_48018);
nand U49649 (N_49649,N_48491,N_48216);
nor U49650 (N_49650,N_48174,N_48386);
xnor U49651 (N_49651,N_48902,N_48063);
nand U49652 (N_49652,N_48075,N_48553);
and U49653 (N_49653,N_48604,N_48400);
or U49654 (N_49654,N_48281,N_48356);
xnor U49655 (N_49655,N_48798,N_48955);
xor U49656 (N_49656,N_48922,N_48960);
xor U49657 (N_49657,N_48016,N_48172);
nand U49658 (N_49658,N_48539,N_48662);
and U49659 (N_49659,N_48101,N_48363);
nor U49660 (N_49660,N_48767,N_48390);
nor U49661 (N_49661,N_48414,N_48583);
nand U49662 (N_49662,N_48011,N_48885);
nor U49663 (N_49663,N_48738,N_48705);
nor U49664 (N_49664,N_48246,N_48916);
nor U49665 (N_49665,N_48576,N_48269);
nand U49666 (N_49666,N_48102,N_48241);
and U49667 (N_49667,N_48664,N_48191);
nand U49668 (N_49668,N_48046,N_48389);
nand U49669 (N_49669,N_48426,N_48199);
nand U49670 (N_49670,N_48118,N_48880);
and U49671 (N_49671,N_48184,N_48752);
xor U49672 (N_49672,N_48765,N_48692);
and U49673 (N_49673,N_48830,N_48924);
and U49674 (N_49674,N_48342,N_48442);
or U49675 (N_49675,N_48152,N_48421);
nor U49676 (N_49676,N_48573,N_48659);
nand U49677 (N_49677,N_48496,N_48653);
nand U49678 (N_49678,N_48758,N_48541);
nand U49679 (N_49679,N_48138,N_48097);
xor U49680 (N_49680,N_48204,N_48538);
nor U49681 (N_49681,N_48849,N_48325);
xor U49682 (N_49682,N_48393,N_48111);
and U49683 (N_49683,N_48967,N_48265);
and U49684 (N_49684,N_48770,N_48381);
nor U49685 (N_49685,N_48181,N_48172);
nor U49686 (N_49686,N_48935,N_48875);
and U49687 (N_49687,N_48033,N_48703);
nand U49688 (N_49688,N_48098,N_48953);
xor U49689 (N_49689,N_48234,N_48971);
nor U49690 (N_49690,N_48178,N_48437);
nor U49691 (N_49691,N_48056,N_48498);
xor U49692 (N_49692,N_48303,N_48135);
or U49693 (N_49693,N_48603,N_48579);
or U49694 (N_49694,N_48659,N_48330);
nand U49695 (N_49695,N_48489,N_48138);
nand U49696 (N_49696,N_48616,N_48254);
xor U49697 (N_49697,N_48388,N_48268);
xor U49698 (N_49698,N_48975,N_48804);
or U49699 (N_49699,N_48511,N_48347);
xor U49700 (N_49700,N_48051,N_48492);
nor U49701 (N_49701,N_48607,N_48460);
and U49702 (N_49702,N_48456,N_48531);
and U49703 (N_49703,N_48413,N_48035);
nor U49704 (N_49704,N_48513,N_48095);
or U49705 (N_49705,N_48728,N_48190);
xor U49706 (N_49706,N_48510,N_48144);
and U49707 (N_49707,N_48119,N_48784);
or U49708 (N_49708,N_48983,N_48937);
nand U49709 (N_49709,N_48467,N_48097);
or U49710 (N_49710,N_48403,N_48821);
or U49711 (N_49711,N_48074,N_48144);
and U49712 (N_49712,N_48019,N_48761);
nor U49713 (N_49713,N_48473,N_48191);
xnor U49714 (N_49714,N_48027,N_48026);
nand U49715 (N_49715,N_48643,N_48104);
nor U49716 (N_49716,N_48702,N_48683);
or U49717 (N_49717,N_48093,N_48427);
or U49718 (N_49718,N_48493,N_48059);
nand U49719 (N_49719,N_48596,N_48318);
nor U49720 (N_49720,N_48241,N_48036);
and U49721 (N_49721,N_48905,N_48817);
nor U49722 (N_49722,N_48448,N_48338);
or U49723 (N_49723,N_48862,N_48414);
nand U49724 (N_49724,N_48110,N_48530);
nand U49725 (N_49725,N_48221,N_48426);
and U49726 (N_49726,N_48896,N_48345);
nand U49727 (N_49727,N_48075,N_48376);
xor U49728 (N_49728,N_48260,N_48226);
or U49729 (N_49729,N_48222,N_48002);
or U49730 (N_49730,N_48722,N_48065);
nor U49731 (N_49731,N_48810,N_48020);
and U49732 (N_49732,N_48585,N_48870);
xnor U49733 (N_49733,N_48705,N_48746);
xnor U49734 (N_49734,N_48757,N_48895);
or U49735 (N_49735,N_48345,N_48492);
nor U49736 (N_49736,N_48635,N_48862);
and U49737 (N_49737,N_48724,N_48381);
xor U49738 (N_49738,N_48660,N_48876);
and U49739 (N_49739,N_48851,N_48774);
or U49740 (N_49740,N_48612,N_48360);
nor U49741 (N_49741,N_48420,N_48737);
or U49742 (N_49742,N_48858,N_48674);
xnor U49743 (N_49743,N_48407,N_48441);
or U49744 (N_49744,N_48052,N_48804);
xor U49745 (N_49745,N_48272,N_48117);
and U49746 (N_49746,N_48851,N_48109);
or U49747 (N_49747,N_48418,N_48575);
and U49748 (N_49748,N_48308,N_48096);
xnor U49749 (N_49749,N_48068,N_48425);
or U49750 (N_49750,N_48515,N_48100);
or U49751 (N_49751,N_48794,N_48895);
or U49752 (N_49752,N_48631,N_48749);
nor U49753 (N_49753,N_48565,N_48471);
nor U49754 (N_49754,N_48674,N_48848);
xor U49755 (N_49755,N_48714,N_48313);
and U49756 (N_49756,N_48901,N_48599);
or U49757 (N_49757,N_48204,N_48944);
xor U49758 (N_49758,N_48634,N_48935);
or U49759 (N_49759,N_48288,N_48563);
or U49760 (N_49760,N_48673,N_48271);
xnor U49761 (N_49761,N_48610,N_48227);
nor U49762 (N_49762,N_48081,N_48880);
nand U49763 (N_49763,N_48958,N_48437);
nand U49764 (N_49764,N_48483,N_48798);
nand U49765 (N_49765,N_48304,N_48692);
nand U49766 (N_49766,N_48500,N_48356);
and U49767 (N_49767,N_48401,N_48120);
nand U49768 (N_49768,N_48913,N_48761);
or U49769 (N_49769,N_48808,N_48799);
xor U49770 (N_49770,N_48326,N_48107);
or U49771 (N_49771,N_48271,N_48920);
nor U49772 (N_49772,N_48195,N_48151);
or U49773 (N_49773,N_48064,N_48706);
nor U49774 (N_49774,N_48294,N_48490);
and U49775 (N_49775,N_48555,N_48288);
xnor U49776 (N_49776,N_48370,N_48554);
nand U49777 (N_49777,N_48036,N_48207);
nor U49778 (N_49778,N_48526,N_48375);
xor U49779 (N_49779,N_48584,N_48013);
nor U49780 (N_49780,N_48180,N_48936);
and U49781 (N_49781,N_48886,N_48681);
or U49782 (N_49782,N_48252,N_48217);
or U49783 (N_49783,N_48875,N_48724);
nor U49784 (N_49784,N_48573,N_48321);
xor U49785 (N_49785,N_48424,N_48450);
nand U49786 (N_49786,N_48877,N_48025);
nand U49787 (N_49787,N_48230,N_48506);
nor U49788 (N_49788,N_48346,N_48730);
nand U49789 (N_49789,N_48946,N_48406);
xor U49790 (N_49790,N_48912,N_48647);
or U49791 (N_49791,N_48717,N_48683);
and U49792 (N_49792,N_48050,N_48810);
xnor U49793 (N_49793,N_48537,N_48574);
or U49794 (N_49794,N_48388,N_48332);
nand U49795 (N_49795,N_48327,N_48010);
nand U49796 (N_49796,N_48386,N_48920);
xor U49797 (N_49797,N_48954,N_48737);
xor U49798 (N_49798,N_48187,N_48833);
and U49799 (N_49799,N_48672,N_48382);
nand U49800 (N_49800,N_48567,N_48374);
nand U49801 (N_49801,N_48386,N_48721);
xor U49802 (N_49802,N_48780,N_48335);
nand U49803 (N_49803,N_48409,N_48964);
xor U49804 (N_49804,N_48197,N_48802);
or U49805 (N_49805,N_48028,N_48820);
or U49806 (N_49806,N_48008,N_48015);
or U49807 (N_49807,N_48216,N_48543);
xnor U49808 (N_49808,N_48074,N_48268);
nor U49809 (N_49809,N_48711,N_48199);
nand U49810 (N_49810,N_48634,N_48568);
and U49811 (N_49811,N_48569,N_48883);
or U49812 (N_49812,N_48461,N_48225);
or U49813 (N_49813,N_48051,N_48701);
xnor U49814 (N_49814,N_48765,N_48461);
and U49815 (N_49815,N_48893,N_48770);
xor U49816 (N_49816,N_48006,N_48678);
xnor U49817 (N_49817,N_48262,N_48659);
nand U49818 (N_49818,N_48377,N_48204);
nor U49819 (N_49819,N_48127,N_48964);
nor U49820 (N_49820,N_48532,N_48983);
nor U49821 (N_49821,N_48656,N_48205);
and U49822 (N_49822,N_48213,N_48191);
nand U49823 (N_49823,N_48837,N_48512);
xnor U49824 (N_49824,N_48736,N_48757);
nor U49825 (N_49825,N_48196,N_48533);
or U49826 (N_49826,N_48680,N_48734);
xnor U49827 (N_49827,N_48390,N_48500);
xor U49828 (N_49828,N_48317,N_48421);
and U49829 (N_49829,N_48199,N_48246);
nand U49830 (N_49830,N_48714,N_48189);
or U49831 (N_49831,N_48306,N_48052);
or U49832 (N_49832,N_48920,N_48904);
nand U49833 (N_49833,N_48850,N_48259);
or U49834 (N_49834,N_48792,N_48334);
or U49835 (N_49835,N_48143,N_48405);
nor U49836 (N_49836,N_48236,N_48211);
nand U49837 (N_49837,N_48884,N_48855);
or U49838 (N_49838,N_48848,N_48655);
and U49839 (N_49839,N_48011,N_48301);
xnor U49840 (N_49840,N_48502,N_48849);
nor U49841 (N_49841,N_48742,N_48783);
nand U49842 (N_49842,N_48588,N_48249);
or U49843 (N_49843,N_48802,N_48218);
nor U49844 (N_49844,N_48763,N_48204);
nand U49845 (N_49845,N_48420,N_48559);
and U49846 (N_49846,N_48347,N_48358);
nand U49847 (N_49847,N_48742,N_48013);
and U49848 (N_49848,N_48784,N_48833);
nand U49849 (N_49849,N_48717,N_48884);
xor U49850 (N_49850,N_48438,N_48563);
nor U49851 (N_49851,N_48675,N_48850);
xor U49852 (N_49852,N_48054,N_48485);
nor U49853 (N_49853,N_48078,N_48223);
or U49854 (N_49854,N_48201,N_48768);
xor U49855 (N_49855,N_48864,N_48968);
or U49856 (N_49856,N_48310,N_48791);
nor U49857 (N_49857,N_48566,N_48171);
and U49858 (N_49858,N_48212,N_48616);
xnor U49859 (N_49859,N_48404,N_48366);
nand U49860 (N_49860,N_48899,N_48589);
and U49861 (N_49861,N_48986,N_48213);
or U49862 (N_49862,N_48725,N_48770);
nor U49863 (N_49863,N_48077,N_48628);
or U49864 (N_49864,N_48126,N_48478);
or U49865 (N_49865,N_48636,N_48131);
and U49866 (N_49866,N_48463,N_48064);
nor U49867 (N_49867,N_48753,N_48720);
and U49868 (N_49868,N_48372,N_48480);
xor U49869 (N_49869,N_48154,N_48784);
or U49870 (N_49870,N_48232,N_48218);
nor U49871 (N_49871,N_48715,N_48053);
or U49872 (N_49872,N_48429,N_48165);
nand U49873 (N_49873,N_48241,N_48938);
or U49874 (N_49874,N_48667,N_48501);
or U49875 (N_49875,N_48165,N_48555);
nor U49876 (N_49876,N_48927,N_48838);
and U49877 (N_49877,N_48083,N_48597);
or U49878 (N_49878,N_48416,N_48571);
and U49879 (N_49879,N_48403,N_48293);
or U49880 (N_49880,N_48425,N_48819);
or U49881 (N_49881,N_48975,N_48244);
and U49882 (N_49882,N_48971,N_48539);
nor U49883 (N_49883,N_48340,N_48841);
or U49884 (N_49884,N_48505,N_48336);
and U49885 (N_49885,N_48278,N_48964);
xnor U49886 (N_49886,N_48630,N_48774);
or U49887 (N_49887,N_48719,N_48711);
and U49888 (N_49888,N_48492,N_48368);
nor U49889 (N_49889,N_48061,N_48458);
and U49890 (N_49890,N_48917,N_48296);
nand U49891 (N_49891,N_48585,N_48358);
and U49892 (N_49892,N_48099,N_48642);
xor U49893 (N_49893,N_48499,N_48911);
nand U49894 (N_49894,N_48317,N_48114);
or U49895 (N_49895,N_48046,N_48407);
nand U49896 (N_49896,N_48496,N_48969);
xor U49897 (N_49897,N_48357,N_48492);
nand U49898 (N_49898,N_48437,N_48792);
xor U49899 (N_49899,N_48312,N_48217);
xor U49900 (N_49900,N_48795,N_48394);
nand U49901 (N_49901,N_48227,N_48188);
nand U49902 (N_49902,N_48075,N_48095);
nand U49903 (N_49903,N_48082,N_48737);
and U49904 (N_49904,N_48853,N_48892);
nor U49905 (N_49905,N_48722,N_48874);
xnor U49906 (N_49906,N_48576,N_48097);
or U49907 (N_49907,N_48085,N_48562);
nand U49908 (N_49908,N_48031,N_48911);
nand U49909 (N_49909,N_48064,N_48302);
and U49910 (N_49910,N_48699,N_48306);
and U49911 (N_49911,N_48257,N_48124);
nand U49912 (N_49912,N_48520,N_48316);
xnor U49913 (N_49913,N_48391,N_48073);
xnor U49914 (N_49914,N_48424,N_48071);
xor U49915 (N_49915,N_48020,N_48267);
and U49916 (N_49916,N_48237,N_48801);
and U49917 (N_49917,N_48082,N_48157);
or U49918 (N_49918,N_48625,N_48705);
or U49919 (N_49919,N_48361,N_48517);
nor U49920 (N_49920,N_48149,N_48757);
xnor U49921 (N_49921,N_48439,N_48398);
nor U49922 (N_49922,N_48393,N_48326);
nor U49923 (N_49923,N_48834,N_48181);
xnor U49924 (N_49924,N_48351,N_48930);
xnor U49925 (N_49925,N_48204,N_48434);
nand U49926 (N_49926,N_48069,N_48429);
nand U49927 (N_49927,N_48676,N_48337);
and U49928 (N_49928,N_48705,N_48747);
and U49929 (N_49929,N_48710,N_48915);
nand U49930 (N_49930,N_48594,N_48278);
nor U49931 (N_49931,N_48772,N_48236);
nand U49932 (N_49932,N_48903,N_48256);
xor U49933 (N_49933,N_48854,N_48534);
or U49934 (N_49934,N_48111,N_48889);
or U49935 (N_49935,N_48126,N_48787);
and U49936 (N_49936,N_48268,N_48854);
xor U49937 (N_49937,N_48466,N_48341);
or U49938 (N_49938,N_48971,N_48793);
nor U49939 (N_49939,N_48150,N_48710);
or U49940 (N_49940,N_48119,N_48007);
nor U49941 (N_49941,N_48849,N_48480);
nand U49942 (N_49942,N_48589,N_48789);
nand U49943 (N_49943,N_48083,N_48032);
xor U49944 (N_49944,N_48504,N_48775);
nand U49945 (N_49945,N_48608,N_48774);
nor U49946 (N_49946,N_48506,N_48205);
xnor U49947 (N_49947,N_48722,N_48949);
xor U49948 (N_49948,N_48985,N_48016);
or U49949 (N_49949,N_48670,N_48663);
and U49950 (N_49950,N_48803,N_48881);
nand U49951 (N_49951,N_48614,N_48746);
or U49952 (N_49952,N_48094,N_48896);
or U49953 (N_49953,N_48321,N_48482);
nand U49954 (N_49954,N_48033,N_48136);
or U49955 (N_49955,N_48504,N_48684);
and U49956 (N_49956,N_48117,N_48473);
or U49957 (N_49957,N_48129,N_48040);
xor U49958 (N_49958,N_48009,N_48647);
or U49959 (N_49959,N_48057,N_48634);
nor U49960 (N_49960,N_48759,N_48557);
xor U49961 (N_49961,N_48896,N_48553);
nor U49962 (N_49962,N_48866,N_48582);
nand U49963 (N_49963,N_48462,N_48212);
nor U49964 (N_49964,N_48491,N_48797);
xor U49965 (N_49965,N_48591,N_48165);
or U49966 (N_49966,N_48111,N_48645);
xor U49967 (N_49967,N_48780,N_48490);
xor U49968 (N_49968,N_48549,N_48454);
xnor U49969 (N_49969,N_48653,N_48256);
nand U49970 (N_49970,N_48693,N_48479);
xor U49971 (N_49971,N_48887,N_48769);
nor U49972 (N_49972,N_48600,N_48743);
nor U49973 (N_49973,N_48643,N_48617);
nor U49974 (N_49974,N_48472,N_48749);
xnor U49975 (N_49975,N_48438,N_48616);
and U49976 (N_49976,N_48035,N_48187);
and U49977 (N_49977,N_48904,N_48867);
xor U49978 (N_49978,N_48777,N_48020);
and U49979 (N_49979,N_48778,N_48060);
or U49980 (N_49980,N_48962,N_48528);
or U49981 (N_49981,N_48124,N_48723);
nand U49982 (N_49982,N_48611,N_48093);
or U49983 (N_49983,N_48641,N_48540);
nor U49984 (N_49984,N_48523,N_48822);
nor U49985 (N_49985,N_48635,N_48642);
or U49986 (N_49986,N_48743,N_48595);
nand U49987 (N_49987,N_48898,N_48437);
nor U49988 (N_49988,N_48660,N_48793);
or U49989 (N_49989,N_48998,N_48762);
and U49990 (N_49990,N_48293,N_48907);
or U49991 (N_49991,N_48066,N_48479);
or U49992 (N_49992,N_48112,N_48326);
nor U49993 (N_49993,N_48367,N_48014);
xnor U49994 (N_49994,N_48220,N_48487);
and U49995 (N_49995,N_48755,N_48702);
nand U49996 (N_49996,N_48473,N_48984);
nand U49997 (N_49997,N_48519,N_48938);
nor U49998 (N_49998,N_48850,N_48876);
or U49999 (N_49999,N_48854,N_48906);
or UO_0 (O_0,N_49380,N_49755);
nand UO_1 (O_1,N_49310,N_49627);
nand UO_2 (O_2,N_49201,N_49996);
or UO_3 (O_3,N_49572,N_49948);
and UO_4 (O_4,N_49679,N_49391);
xor UO_5 (O_5,N_49161,N_49327);
or UO_6 (O_6,N_49997,N_49734);
or UO_7 (O_7,N_49731,N_49284);
nand UO_8 (O_8,N_49769,N_49180);
and UO_9 (O_9,N_49610,N_49272);
nor UO_10 (O_10,N_49780,N_49301);
nor UO_11 (O_11,N_49316,N_49534);
nand UO_12 (O_12,N_49902,N_49459);
or UO_13 (O_13,N_49417,N_49237);
nand UO_14 (O_14,N_49479,N_49430);
xor UO_15 (O_15,N_49596,N_49289);
or UO_16 (O_16,N_49219,N_49709);
xor UO_17 (O_17,N_49091,N_49633);
xor UO_18 (O_18,N_49052,N_49384);
nor UO_19 (O_19,N_49676,N_49949);
and UO_20 (O_20,N_49364,N_49764);
and UO_21 (O_21,N_49625,N_49507);
and UO_22 (O_22,N_49098,N_49589);
nand UO_23 (O_23,N_49887,N_49650);
nand UO_24 (O_24,N_49810,N_49136);
nor UO_25 (O_25,N_49279,N_49736);
and UO_26 (O_26,N_49646,N_49939);
nor UO_27 (O_27,N_49118,N_49290);
and UO_28 (O_28,N_49623,N_49457);
and UO_29 (O_29,N_49607,N_49154);
or UO_30 (O_30,N_49894,N_49465);
xnor UO_31 (O_31,N_49067,N_49250);
and UO_32 (O_32,N_49382,N_49271);
xor UO_33 (O_33,N_49409,N_49211);
or UO_34 (O_34,N_49852,N_49196);
nor UO_35 (O_35,N_49282,N_49673);
xnor UO_36 (O_36,N_49065,N_49022);
nand UO_37 (O_37,N_49719,N_49573);
nand UO_38 (O_38,N_49675,N_49372);
nand UO_39 (O_39,N_49790,N_49733);
nor UO_40 (O_40,N_49670,N_49492);
nor UO_41 (O_41,N_49622,N_49661);
nand UO_42 (O_42,N_49421,N_49545);
xor UO_43 (O_43,N_49376,N_49657);
and UO_44 (O_44,N_49975,N_49109);
and UO_45 (O_45,N_49268,N_49544);
xnor UO_46 (O_46,N_49163,N_49908);
xor UO_47 (O_47,N_49805,N_49885);
xnor UO_48 (O_48,N_49436,N_49818);
nor UO_49 (O_49,N_49016,N_49049);
xor UO_50 (O_50,N_49634,N_49449);
nor UO_51 (O_51,N_49744,N_49814);
nor UO_52 (O_52,N_49159,N_49139);
or UO_53 (O_53,N_49379,N_49728);
or UO_54 (O_54,N_49010,N_49796);
nor UO_55 (O_55,N_49555,N_49835);
xor UO_56 (O_56,N_49559,N_49832);
nand UO_57 (O_57,N_49145,N_49097);
and UO_58 (O_58,N_49432,N_49234);
nand UO_59 (O_59,N_49225,N_49073);
or UO_60 (O_60,N_49714,N_49864);
nand UO_61 (O_61,N_49438,N_49685);
or UO_62 (O_62,N_49226,N_49228);
nor UO_63 (O_63,N_49880,N_49392);
or UO_64 (O_64,N_49811,N_49355);
and UO_65 (O_65,N_49490,N_49952);
and UO_66 (O_66,N_49004,N_49577);
or UO_67 (O_67,N_49023,N_49322);
and UO_68 (O_68,N_49352,N_49450);
nor UO_69 (O_69,N_49717,N_49982);
xor UO_70 (O_70,N_49207,N_49765);
or UO_71 (O_71,N_49581,N_49215);
and UO_72 (O_72,N_49482,N_49970);
xor UO_73 (O_73,N_49303,N_49204);
nor UO_74 (O_74,N_49969,N_49149);
or UO_75 (O_75,N_49531,N_49822);
or UO_76 (O_76,N_49278,N_49587);
nor UO_77 (O_77,N_49339,N_49690);
nor UO_78 (O_78,N_49043,N_49433);
nand UO_79 (O_79,N_49486,N_49759);
or UO_80 (O_80,N_49963,N_49980);
nor UO_81 (O_81,N_49655,N_49312);
xnor UO_82 (O_82,N_49720,N_49954);
and UO_83 (O_83,N_49236,N_49048);
and UO_84 (O_84,N_49493,N_49513);
nor UO_85 (O_85,N_49924,N_49027);
and UO_86 (O_86,N_49659,N_49718);
xor UO_87 (O_87,N_49860,N_49212);
and UO_88 (O_88,N_49682,N_49746);
xor UO_89 (O_89,N_49406,N_49265);
and UO_90 (O_90,N_49653,N_49428);
nand UO_91 (O_91,N_49815,N_49509);
and UO_92 (O_92,N_49264,N_49414);
nand UO_93 (O_93,N_49754,N_49866);
nand UO_94 (O_94,N_49884,N_49134);
nor UO_95 (O_95,N_49167,N_49079);
nand UO_96 (O_96,N_49307,N_49407);
and UO_97 (O_97,N_49127,N_49514);
and UO_98 (O_98,N_49710,N_49671);
and UO_99 (O_99,N_49504,N_49546);
nor UO_100 (O_100,N_49605,N_49468);
xnor UO_101 (O_101,N_49617,N_49130);
or UO_102 (O_102,N_49213,N_49711);
nand UO_103 (O_103,N_49171,N_49469);
nand UO_104 (O_104,N_49491,N_49704);
or UO_105 (O_105,N_49242,N_49060);
xor UO_106 (O_106,N_49099,N_49606);
nand UO_107 (O_107,N_49697,N_49920);
nor UO_108 (O_108,N_49680,N_49967);
and UO_109 (O_109,N_49813,N_49828);
nor UO_110 (O_110,N_49648,N_49837);
or UO_111 (O_111,N_49886,N_49888);
nor UO_112 (O_112,N_49441,N_49463);
nand UO_113 (O_113,N_49988,N_49294);
and UO_114 (O_114,N_49921,N_49799);
or UO_115 (O_115,N_49732,N_49245);
nor UO_116 (O_116,N_49007,N_49834);
or UO_117 (O_117,N_49907,N_49055);
xnor UO_118 (O_118,N_49524,N_49229);
nand UO_119 (O_119,N_49692,N_49730);
or UO_120 (O_120,N_49873,N_49470);
and UO_121 (O_121,N_49683,N_49585);
nand UO_122 (O_122,N_49054,N_49342);
nand UO_123 (O_123,N_49235,N_49981);
nand UO_124 (O_124,N_49946,N_49713);
or UO_125 (O_125,N_49929,N_49926);
or UO_126 (O_126,N_49770,N_49418);
nand UO_127 (O_127,N_49898,N_49181);
xnor UO_128 (O_128,N_49398,N_49529);
xnor UO_129 (O_129,N_49508,N_49481);
and UO_130 (O_130,N_49602,N_49241);
and UO_131 (O_131,N_49269,N_49554);
xor UO_132 (O_132,N_49176,N_49495);
xor UO_133 (O_133,N_49341,N_49752);
and UO_134 (O_134,N_49773,N_49846);
or UO_135 (O_135,N_49345,N_49977);
nor UO_136 (O_136,N_49930,N_49938);
nor UO_137 (O_137,N_49120,N_49367);
or UO_138 (O_138,N_49257,N_49096);
or UO_139 (O_139,N_49922,N_49701);
nor UO_140 (O_140,N_49255,N_49893);
nor UO_141 (O_141,N_49574,N_49878);
nor UO_142 (O_142,N_49350,N_49360);
or UO_143 (O_143,N_49933,N_49896);
or UO_144 (O_144,N_49905,N_49590);
nand UO_145 (O_145,N_49941,N_49368);
and UO_146 (O_146,N_49777,N_49974);
nor UO_147 (O_147,N_49801,N_49044);
or UO_148 (O_148,N_49859,N_49900);
nor UO_149 (O_149,N_49081,N_49793);
and UO_150 (O_150,N_49137,N_49447);
xnor UO_151 (O_151,N_49369,N_49439);
nor UO_152 (O_152,N_49912,N_49336);
or UO_153 (O_153,N_49831,N_49408);
and UO_154 (O_154,N_49387,N_49442);
xnor UO_155 (O_155,N_49550,N_49543);
or UO_156 (O_156,N_49494,N_49522);
nand UO_157 (O_157,N_49142,N_49412);
or UO_158 (O_158,N_49259,N_49173);
nand UO_159 (O_159,N_49185,N_49735);
xnor UO_160 (O_160,N_49045,N_49128);
nor UO_161 (O_161,N_49666,N_49253);
xnor UO_162 (O_162,N_49512,N_49498);
and UO_163 (O_163,N_49454,N_49030);
and UO_164 (O_164,N_49363,N_49218);
nor UO_165 (O_165,N_49381,N_49869);
and UO_166 (O_166,N_49068,N_49784);
nor UO_167 (O_167,N_49458,N_49937);
xnor UO_168 (O_168,N_49779,N_49283);
nand UO_169 (O_169,N_49961,N_49162);
xnor UO_170 (O_170,N_49575,N_49089);
or UO_171 (O_171,N_49652,N_49419);
or UO_172 (O_172,N_49865,N_49936);
xor UO_173 (O_173,N_49103,N_49361);
or UO_174 (O_174,N_49612,N_49526);
or UO_175 (O_175,N_49778,N_49404);
nand UO_176 (O_176,N_49621,N_49170);
nor UO_177 (O_177,N_49989,N_49199);
nor UO_178 (O_178,N_49348,N_49667);
xnor UO_179 (O_179,N_49768,N_49193);
and UO_180 (O_180,N_49246,N_49824);
xor UO_181 (O_181,N_49791,N_49147);
and UO_182 (O_182,N_49940,N_49636);
nand UO_183 (O_183,N_49277,N_49110);
and UO_184 (O_184,N_49323,N_49783);
xor UO_185 (O_185,N_49040,N_49928);
and UO_186 (O_186,N_49474,N_49133);
nor UO_187 (O_187,N_49674,N_49453);
nor UO_188 (O_188,N_49399,N_49314);
xnor UO_189 (O_189,N_49809,N_49182);
and UO_190 (O_190,N_49725,N_49613);
and UO_191 (O_191,N_49897,N_49210);
and UO_192 (O_192,N_49415,N_49808);
xor UO_193 (O_193,N_49416,N_49955);
xor UO_194 (O_194,N_49155,N_49200);
xor UO_195 (O_195,N_49552,N_49321);
nand UO_196 (O_196,N_49035,N_49861);
or UO_197 (O_197,N_49797,N_49082);
nand UO_198 (O_198,N_49292,N_49645);
nor UO_199 (O_199,N_49743,N_49335);
and UO_200 (O_200,N_49538,N_49231);
or UO_201 (O_201,N_49338,N_49568);
or UO_202 (O_202,N_49413,N_49702);
nand UO_203 (O_203,N_49856,N_49817);
and UO_204 (O_204,N_49203,N_49121);
or UO_205 (O_205,N_49841,N_49558);
xnor UO_206 (O_206,N_49947,N_49086);
nor UO_207 (O_207,N_49388,N_49076);
or UO_208 (O_208,N_49169,N_49148);
nor UO_209 (O_209,N_49631,N_49224);
nor UO_210 (O_210,N_49001,N_49951);
or UO_211 (O_211,N_49911,N_49564);
and UO_212 (O_212,N_49340,N_49537);
and UO_213 (O_213,N_49140,N_49456);
nand UO_214 (O_214,N_49978,N_49757);
or UO_215 (O_215,N_49373,N_49243);
nor UO_216 (O_216,N_49638,N_49496);
or UO_217 (O_217,N_49729,N_49480);
xnor UO_218 (O_218,N_49998,N_49593);
xor UO_219 (O_219,N_49668,N_49117);
nor UO_220 (O_220,N_49346,N_49402);
nor UO_221 (O_221,N_49230,N_49895);
nor UO_222 (O_222,N_49037,N_49074);
xor UO_223 (O_223,N_49249,N_49254);
or UO_224 (O_224,N_49077,N_49582);
or UO_225 (O_225,N_49792,N_49324);
and UO_226 (O_226,N_49851,N_49694);
xnor UO_227 (O_227,N_49800,N_49319);
and UO_228 (O_228,N_49611,N_49516);
or UO_229 (O_229,N_49429,N_49700);
nand UO_230 (O_230,N_49113,N_49641);
or UO_231 (O_231,N_49256,N_49329);
nor UO_232 (O_232,N_49775,N_49706);
nor UO_233 (O_233,N_49431,N_49842);
or UO_234 (O_234,N_49542,N_49062);
nand UO_235 (O_235,N_49839,N_49644);
or UO_236 (O_236,N_49080,N_49325);
and UO_237 (O_237,N_49308,N_49616);
xnor UO_238 (O_238,N_49958,N_49475);
xnor UO_239 (O_239,N_49987,N_49553);
and UO_240 (O_240,N_49177,N_49530);
and UO_241 (O_241,N_49991,N_49070);
or UO_242 (O_242,N_49695,N_49000);
and UO_243 (O_243,N_49845,N_49385);
nand UO_244 (O_244,N_49354,N_49488);
xor UO_245 (O_245,N_49427,N_49571);
xnor UO_246 (O_246,N_49390,N_49515);
and UO_247 (O_247,N_49297,N_49789);
nand UO_248 (O_248,N_49464,N_49288);
xnor UO_249 (O_249,N_49807,N_49258);
nand UO_250 (O_250,N_49506,N_49262);
nor UO_251 (O_251,N_49051,N_49038);
or UO_252 (O_252,N_49748,N_49957);
xnor UO_253 (O_253,N_49665,N_49609);
or UO_254 (O_254,N_49707,N_49901);
or UO_255 (O_255,N_49794,N_49267);
or UO_256 (O_256,N_49643,N_49143);
xor UO_257 (O_257,N_49761,N_49150);
nand UO_258 (O_258,N_49604,N_49194);
nor UO_259 (O_259,N_49715,N_49471);
or UO_260 (O_260,N_49050,N_49642);
nor UO_261 (O_261,N_49510,N_49039);
or UO_262 (O_262,N_49280,N_49461);
or UO_263 (O_263,N_49699,N_49591);
xor UO_264 (O_264,N_49497,N_49078);
or UO_265 (O_265,N_49838,N_49222);
or UO_266 (O_266,N_49247,N_49124);
or UO_267 (O_267,N_49890,N_49615);
and UO_268 (O_268,N_49260,N_49628);
nand UO_269 (O_269,N_49108,N_49401);
xnor UO_270 (O_270,N_49477,N_49787);
and UO_271 (O_271,N_49011,N_49239);
nor UO_272 (O_272,N_49812,N_49141);
xnor UO_273 (O_273,N_49651,N_49012);
or UO_274 (O_274,N_49446,N_49105);
nor UO_275 (O_275,N_49750,N_49008);
and UO_276 (O_276,N_49904,N_49021);
nor UO_277 (O_277,N_49209,N_49122);
or UO_278 (O_278,N_49870,N_49330);
nand UO_279 (O_279,N_49383,N_49959);
and UO_280 (O_280,N_49548,N_49956);
or UO_281 (O_281,N_49934,N_49567);
nand UO_282 (O_282,N_49351,N_49501);
nand UO_283 (O_283,N_49662,N_49208);
or UO_284 (O_284,N_49462,N_49024);
or UO_285 (O_285,N_49036,N_49910);
and UO_286 (O_286,N_49296,N_49640);
xor UO_287 (O_287,N_49485,N_49273);
nand UO_288 (O_288,N_49397,N_49104);
and UO_289 (O_289,N_49649,N_49756);
nand UO_290 (O_290,N_49891,N_49523);
and UO_291 (O_291,N_49899,N_49374);
xor UO_292 (O_292,N_49976,N_49002);
or UO_293 (O_293,N_49825,N_49527);
and UO_294 (O_294,N_49424,N_49983);
or UO_295 (O_295,N_49119,N_49266);
xnor UO_296 (O_296,N_49708,N_49018);
nand UO_297 (O_297,N_49999,N_49326);
nor UO_298 (O_298,N_49608,N_49451);
and UO_299 (O_299,N_49563,N_49992);
or UO_300 (O_300,N_49460,N_49804);
nand UO_301 (O_301,N_49356,N_49315);
and UO_302 (O_302,N_49132,N_49619);
xnor UO_303 (O_303,N_49183,N_49723);
xor UO_304 (O_304,N_49802,N_49875);
xnor UO_305 (O_305,N_49214,N_49935);
or UO_306 (O_306,N_49738,N_49767);
and UO_307 (O_307,N_49047,N_49985);
nor UO_308 (O_308,N_49393,N_49663);
nand UO_309 (O_309,N_49931,N_49557);
or UO_310 (O_310,N_49320,N_49600);
nand UO_311 (O_311,N_49857,N_49740);
and UO_312 (O_312,N_49422,N_49854);
xor UO_313 (O_313,N_49549,N_49071);
or UO_314 (O_314,N_49853,N_49064);
nand UO_315 (O_315,N_49306,N_49305);
or UO_316 (O_316,N_49343,N_49276);
xnor UO_317 (O_317,N_49594,N_49503);
xnor UO_318 (O_318,N_49227,N_49069);
xnor UO_319 (O_319,N_49561,N_49090);
or UO_320 (O_320,N_49198,N_49906);
and UO_321 (O_321,N_49125,N_49112);
nor UO_322 (O_322,N_49876,N_49144);
and UO_323 (O_323,N_49165,N_49100);
or UO_324 (O_324,N_49129,N_49855);
and UO_325 (O_325,N_49932,N_49614);
xor UO_326 (O_326,N_49487,N_49620);
nor UO_327 (O_327,N_49032,N_49362);
nand UO_328 (O_328,N_49309,N_49295);
xor UO_329 (O_329,N_49116,N_49019);
nand UO_330 (O_330,N_49874,N_49909);
nand UO_331 (O_331,N_49088,N_49131);
xor UO_332 (O_332,N_49862,N_49584);
xnor UO_333 (O_333,N_49505,N_49009);
and UO_334 (O_334,N_49721,N_49377);
or UO_335 (O_335,N_49502,N_49601);
nand UO_336 (O_336,N_49889,N_49483);
nand UO_337 (O_337,N_49025,N_49058);
nor UO_338 (O_338,N_49848,N_49172);
nor UO_339 (O_339,N_49240,N_49261);
and UO_340 (O_340,N_49858,N_49703);
nor UO_341 (O_341,N_49688,N_49565);
xor UO_342 (O_342,N_49473,N_49164);
xor UO_343 (O_343,N_49686,N_49677);
nand UO_344 (O_344,N_49588,N_49195);
xor UO_345 (O_345,N_49101,N_49107);
nand UO_346 (O_346,N_49389,N_49629);
nor UO_347 (O_347,N_49344,N_49293);
and UO_348 (O_348,N_49484,N_49111);
or UO_349 (O_349,N_49892,N_49972);
nand UO_350 (O_350,N_49467,N_49034);
and UO_351 (O_351,N_49916,N_49075);
nor UO_352 (O_352,N_49434,N_49114);
nor UO_353 (O_353,N_49806,N_49445);
nor UO_354 (O_354,N_49925,N_49583);
nor UO_355 (O_355,N_49915,N_49191);
nor UO_356 (O_356,N_49973,N_49206);
nand UO_357 (O_357,N_49712,N_49375);
and UO_358 (O_358,N_49093,N_49664);
xnor UO_359 (O_359,N_49190,N_49106);
xnor UO_360 (O_360,N_49281,N_49452);
nor UO_361 (O_361,N_49216,N_49437);
or UO_362 (O_362,N_49592,N_49304);
and UO_363 (O_363,N_49849,N_49092);
nor UO_364 (O_364,N_49302,N_49877);
nor UO_365 (O_365,N_49238,N_49146);
and UO_366 (O_366,N_49472,N_49371);
nand UO_367 (O_367,N_49971,N_49626);
or UO_368 (O_368,N_49705,N_49400);
and UO_369 (O_369,N_49440,N_49739);
nor UO_370 (O_370,N_49576,N_49160);
nor UO_371 (O_371,N_49881,N_49006);
or UO_372 (O_372,N_49347,N_49722);
nand UO_373 (O_373,N_49580,N_49031);
nor UO_374 (O_374,N_49598,N_49727);
and UO_375 (O_375,N_49205,N_49681);
or UO_376 (O_376,N_49003,N_49630);
or UO_377 (O_377,N_49691,N_49994);
and UO_378 (O_378,N_49244,N_49370);
xor UO_379 (O_379,N_49313,N_49053);
nor UO_380 (O_380,N_49532,N_49639);
nor UO_381 (O_381,N_49152,N_49252);
nand UO_382 (O_382,N_49747,N_49328);
nor UO_383 (O_383,N_49556,N_49882);
or UO_384 (O_384,N_49560,N_49175);
or UO_385 (O_385,N_49521,N_49803);
or UO_386 (O_386,N_49923,N_49126);
nor UO_387 (O_387,N_49833,N_49063);
nor UO_388 (O_388,N_49156,N_49795);
xor UO_389 (O_389,N_49816,N_49918);
and UO_390 (O_390,N_49562,N_49840);
or UO_391 (O_391,N_49396,N_49566);
xor UO_392 (O_392,N_49540,N_49410);
or UO_393 (O_393,N_49046,N_49395);
or UO_394 (O_394,N_49760,N_49518);
xor UO_395 (O_395,N_49263,N_49829);
or UO_396 (O_396,N_49017,N_49174);
nand UO_397 (O_397,N_49300,N_49960);
nand UO_398 (O_398,N_49551,N_49569);
or UO_399 (O_399,N_49466,N_49741);
nor UO_400 (O_400,N_49693,N_49425);
and UO_401 (O_401,N_49353,N_49123);
and UO_402 (O_402,N_49084,N_49072);
nand UO_403 (O_403,N_49270,N_49570);
nor UO_404 (O_404,N_49758,N_49197);
nand UO_405 (O_405,N_49637,N_49157);
nor UO_406 (O_406,N_49285,N_49232);
and UO_407 (O_407,N_49299,N_49830);
nand UO_408 (O_408,N_49669,N_49448);
and UO_409 (O_409,N_49057,N_49943);
or UO_410 (O_410,N_49349,N_49083);
or UO_411 (O_411,N_49085,N_49950);
nor UO_412 (O_412,N_49333,N_49528);
nand UO_413 (O_413,N_49358,N_49188);
nor UO_414 (O_414,N_49726,N_49578);
or UO_415 (O_415,N_49026,N_49378);
xnor UO_416 (O_416,N_49318,N_49403);
xor UO_417 (O_417,N_49724,N_49595);
xnor UO_418 (O_418,N_49094,N_49095);
and UO_419 (O_419,N_49656,N_49586);
xor UO_420 (O_420,N_49995,N_49334);
nor UO_421 (O_421,N_49499,N_49944);
or UO_422 (O_422,N_49763,N_49455);
and UO_423 (O_423,N_49015,N_49984);
nand UO_424 (O_424,N_49635,N_49913);
nor UO_425 (O_425,N_49426,N_49771);
and UO_426 (O_426,N_49337,N_49056);
or UO_427 (O_427,N_49879,N_49766);
nor UO_428 (O_428,N_49696,N_49903);
or UO_429 (O_429,N_49749,N_49168);
nand UO_430 (O_430,N_49359,N_49444);
nand UO_431 (O_431,N_49966,N_49654);
nand UO_432 (O_432,N_49762,N_49192);
nand UO_433 (O_433,N_49115,N_49423);
nand UO_434 (O_434,N_49287,N_49624);
nand UO_435 (O_435,N_49579,N_49962);
xor UO_436 (O_436,N_49511,N_49689);
nand UO_437 (O_437,N_49500,N_49990);
and UO_438 (O_438,N_49737,N_49979);
and UO_439 (O_439,N_49151,N_49827);
and UO_440 (O_440,N_49914,N_49751);
nor UO_441 (O_441,N_49535,N_49883);
nand UO_442 (O_442,N_49217,N_49138);
nor UO_443 (O_443,N_49476,N_49774);
nand UO_444 (O_444,N_49435,N_49742);
nor UO_445 (O_445,N_49357,N_49520);
xor UO_446 (O_446,N_49823,N_49964);
nand UO_447 (O_447,N_49843,N_49184);
xor UO_448 (O_448,N_49221,N_49365);
or UO_449 (O_449,N_49153,N_49678);
or UO_450 (O_450,N_49863,N_49684);
nand UO_451 (O_451,N_49298,N_49785);
and UO_452 (O_452,N_49539,N_49993);
nor UO_453 (O_453,N_49716,N_49632);
nand UO_454 (O_454,N_49867,N_49618);
nor UO_455 (O_455,N_49223,N_49033);
xor UO_456 (O_456,N_49687,N_49519);
xor UO_457 (O_457,N_49411,N_49248);
and UO_458 (O_458,N_49847,N_49291);
nor UO_459 (O_459,N_49087,N_49821);
xnor UO_460 (O_460,N_49772,N_49233);
nor UO_461 (O_461,N_49917,N_49014);
or UO_462 (O_462,N_49541,N_49872);
nand UO_463 (O_463,N_49753,N_49919);
nor UO_464 (O_464,N_49061,N_49186);
or UO_465 (O_465,N_49332,N_49745);
nand UO_466 (O_466,N_49029,N_49536);
xnor UO_467 (O_467,N_49420,N_49776);
xor UO_468 (O_468,N_49819,N_49158);
or UO_469 (O_469,N_49286,N_49826);
and UO_470 (O_470,N_49603,N_49274);
or UO_471 (O_471,N_49311,N_49850);
nand UO_472 (O_472,N_49597,N_49331);
xor UO_473 (O_473,N_49028,N_49443);
and UO_474 (O_474,N_49945,N_49135);
nor UO_475 (O_475,N_49868,N_49178);
nor UO_476 (O_476,N_49366,N_49968);
nor UO_477 (O_477,N_49220,N_49042);
xnor UO_478 (O_478,N_49179,N_49489);
and UO_479 (O_479,N_49005,N_49478);
or UO_480 (O_480,N_49965,N_49647);
or UO_481 (O_481,N_49394,N_49942);
nand UO_482 (O_482,N_49525,N_49781);
xor UO_483 (O_483,N_49013,N_49698);
and UO_484 (O_484,N_49166,N_49820);
xor UO_485 (O_485,N_49547,N_49871);
nand UO_486 (O_486,N_49660,N_49202);
nor UO_487 (O_487,N_49275,N_49844);
xor UO_488 (O_488,N_49672,N_49405);
or UO_489 (O_489,N_49927,N_49066);
nand UO_490 (O_490,N_49788,N_49798);
nand UO_491 (O_491,N_49251,N_49517);
and UO_492 (O_492,N_49317,N_49386);
nand UO_493 (O_493,N_49599,N_49533);
nor UO_494 (O_494,N_49020,N_49953);
nand UO_495 (O_495,N_49986,N_49187);
and UO_496 (O_496,N_49786,N_49836);
or UO_497 (O_497,N_49102,N_49658);
nor UO_498 (O_498,N_49189,N_49059);
nand UO_499 (O_499,N_49041,N_49782);
nor UO_500 (O_500,N_49110,N_49300);
and UO_501 (O_501,N_49078,N_49988);
nand UO_502 (O_502,N_49001,N_49499);
xnor UO_503 (O_503,N_49356,N_49432);
nand UO_504 (O_504,N_49482,N_49531);
and UO_505 (O_505,N_49973,N_49944);
and UO_506 (O_506,N_49857,N_49449);
or UO_507 (O_507,N_49731,N_49131);
or UO_508 (O_508,N_49249,N_49751);
nand UO_509 (O_509,N_49525,N_49299);
nor UO_510 (O_510,N_49460,N_49721);
nor UO_511 (O_511,N_49126,N_49614);
or UO_512 (O_512,N_49951,N_49165);
xor UO_513 (O_513,N_49004,N_49684);
nand UO_514 (O_514,N_49892,N_49256);
and UO_515 (O_515,N_49249,N_49367);
and UO_516 (O_516,N_49253,N_49919);
and UO_517 (O_517,N_49280,N_49652);
xor UO_518 (O_518,N_49853,N_49244);
nor UO_519 (O_519,N_49520,N_49681);
xnor UO_520 (O_520,N_49949,N_49560);
or UO_521 (O_521,N_49645,N_49822);
or UO_522 (O_522,N_49040,N_49820);
or UO_523 (O_523,N_49737,N_49260);
and UO_524 (O_524,N_49634,N_49498);
or UO_525 (O_525,N_49858,N_49914);
or UO_526 (O_526,N_49344,N_49255);
nor UO_527 (O_527,N_49455,N_49423);
nor UO_528 (O_528,N_49372,N_49856);
or UO_529 (O_529,N_49504,N_49267);
or UO_530 (O_530,N_49566,N_49960);
nor UO_531 (O_531,N_49771,N_49774);
nor UO_532 (O_532,N_49581,N_49315);
nand UO_533 (O_533,N_49341,N_49092);
or UO_534 (O_534,N_49448,N_49138);
and UO_535 (O_535,N_49196,N_49759);
or UO_536 (O_536,N_49555,N_49836);
nor UO_537 (O_537,N_49678,N_49807);
nand UO_538 (O_538,N_49050,N_49410);
and UO_539 (O_539,N_49588,N_49534);
nand UO_540 (O_540,N_49949,N_49431);
nor UO_541 (O_541,N_49313,N_49728);
xnor UO_542 (O_542,N_49634,N_49299);
and UO_543 (O_543,N_49573,N_49842);
xor UO_544 (O_544,N_49602,N_49261);
xnor UO_545 (O_545,N_49599,N_49976);
or UO_546 (O_546,N_49591,N_49379);
or UO_547 (O_547,N_49695,N_49792);
or UO_548 (O_548,N_49068,N_49020);
or UO_549 (O_549,N_49507,N_49277);
or UO_550 (O_550,N_49813,N_49688);
and UO_551 (O_551,N_49113,N_49609);
xnor UO_552 (O_552,N_49400,N_49201);
or UO_553 (O_553,N_49111,N_49079);
or UO_554 (O_554,N_49280,N_49352);
nand UO_555 (O_555,N_49919,N_49716);
or UO_556 (O_556,N_49573,N_49297);
nand UO_557 (O_557,N_49825,N_49756);
nand UO_558 (O_558,N_49945,N_49820);
nor UO_559 (O_559,N_49550,N_49253);
nor UO_560 (O_560,N_49390,N_49624);
xnor UO_561 (O_561,N_49025,N_49032);
and UO_562 (O_562,N_49517,N_49278);
or UO_563 (O_563,N_49068,N_49803);
or UO_564 (O_564,N_49396,N_49092);
nand UO_565 (O_565,N_49235,N_49301);
nor UO_566 (O_566,N_49103,N_49283);
and UO_567 (O_567,N_49418,N_49365);
and UO_568 (O_568,N_49177,N_49244);
nand UO_569 (O_569,N_49735,N_49635);
or UO_570 (O_570,N_49914,N_49280);
xor UO_571 (O_571,N_49329,N_49926);
or UO_572 (O_572,N_49351,N_49710);
or UO_573 (O_573,N_49418,N_49140);
nor UO_574 (O_574,N_49419,N_49835);
nand UO_575 (O_575,N_49914,N_49893);
xor UO_576 (O_576,N_49790,N_49737);
xnor UO_577 (O_577,N_49364,N_49427);
xnor UO_578 (O_578,N_49290,N_49301);
nor UO_579 (O_579,N_49364,N_49812);
nand UO_580 (O_580,N_49063,N_49250);
or UO_581 (O_581,N_49162,N_49198);
or UO_582 (O_582,N_49313,N_49585);
nand UO_583 (O_583,N_49936,N_49960);
or UO_584 (O_584,N_49975,N_49075);
or UO_585 (O_585,N_49427,N_49673);
nor UO_586 (O_586,N_49949,N_49051);
nand UO_587 (O_587,N_49989,N_49256);
nor UO_588 (O_588,N_49172,N_49038);
and UO_589 (O_589,N_49417,N_49724);
or UO_590 (O_590,N_49026,N_49268);
nand UO_591 (O_591,N_49258,N_49924);
nor UO_592 (O_592,N_49599,N_49614);
nor UO_593 (O_593,N_49567,N_49349);
nand UO_594 (O_594,N_49033,N_49150);
nand UO_595 (O_595,N_49798,N_49649);
xnor UO_596 (O_596,N_49531,N_49006);
or UO_597 (O_597,N_49304,N_49657);
or UO_598 (O_598,N_49392,N_49866);
and UO_599 (O_599,N_49076,N_49517);
xnor UO_600 (O_600,N_49531,N_49120);
or UO_601 (O_601,N_49412,N_49023);
nor UO_602 (O_602,N_49633,N_49808);
or UO_603 (O_603,N_49520,N_49317);
nand UO_604 (O_604,N_49283,N_49335);
xor UO_605 (O_605,N_49094,N_49885);
xnor UO_606 (O_606,N_49262,N_49433);
or UO_607 (O_607,N_49225,N_49649);
nand UO_608 (O_608,N_49541,N_49802);
nand UO_609 (O_609,N_49364,N_49578);
or UO_610 (O_610,N_49337,N_49810);
nand UO_611 (O_611,N_49574,N_49796);
and UO_612 (O_612,N_49157,N_49645);
and UO_613 (O_613,N_49812,N_49802);
xnor UO_614 (O_614,N_49559,N_49782);
or UO_615 (O_615,N_49116,N_49858);
nor UO_616 (O_616,N_49157,N_49754);
nand UO_617 (O_617,N_49124,N_49185);
and UO_618 (O_618,N_49130,N_49373);
xnor UO_619 (O_619,N_49150,N_49726);
xor UO_620 (O_620,N_49727,N_49071);
xor UO_621 (O_621,N_49237,N_49885);
nand UO_622 (O_622,N_49516,N_49399);
nor UO_623 (O_623,N_49200,N_49439);
nor UO_624 (O_624,N_49909,N_49574);
and UO_625 (O_625,N_49573,N_49803);
xor UO_626 (O_626,N_49504,N_49950);
and UO_627 (O_627,N_49672,N_49889);
and UO_628 (O_628,N_49055,N_49894);
xnor UO_629 (O_629,N_49865,N_49329);
or UO_630 (O_630,N_49275,N_49355);
nor UO_631 (O_631,N_49269,N_49567);
xnor UO_632 (O_632,N_49383,N_49755);
or UO_633 (O_633,N_49018,N_49633);
or UO_634 (O_634,N_49463,N_49776);
xor UO_635 (O_635,N_49578,N_49566);
or UO_636 (O_636,N_49817,N_49344);
xor UO_637 (O_637,N_49627,N_49995);
nand UO_638 (O_638,N_49231,N_49414);
nor UO_639 (O_639,N_49329,N_49493);
xnor UO_640 (O_640,N_49320,N_49051);
xor UO_641 (O_641,N_49557,N_49542);
or UO_642 (O_642,N_49351,N_49880);
xnor UO_643 (O_643,N_49797,N_49180);
nand UO_644 (O_644,N_49364,N_49356);
nor UO_645 (O_645,N_49450,N_49752);
nand UO_646 (O_646,N_49898,N_49509);
xor UO_647 (O_647,N_49444,N_49997);
nor UO_648 (O_648,N_49855,N_49916);
nand UO_649 (O_649,N_49712,N_49077);
xnor UO_650 (O_650,N_49847,N_49086);
xor UO_651 (O_651,N_49231,N_49485);
nor UO_652 (O_652,N_49962,N_49509);
and UO_653 (O_653,N_49799,N_49778);
or UO_654 (O_654,N_49217,N_49024);
xor UO_655 (O_655,N_49486,N_49982);
and UO_656 (O_656,N_49053,N_49178);
or UO_657 (O_657,N_49669,N_49449);
xor UO_658 (O_658,N_49905,N_49198);
or UO_659 (O_659,N_49365,N_49532);
nor UO_660 (O_660,N_49964,N_49481);
nor UO_661 (O_661,N_49301,N_49824);
xor UO_662 (O_662,N_49559,N_49495);
nand UO_663 (O_663,N_49348,N_49507);
nor UO_664 (O_664,N_49975,N_49608);
and UO_665 (O_665,N_49008,N_49295);
xor UO_666 (O_666,N_49957,N_49819);
nor UO_667 (O_667,N_49074,N_49080);
or UO_668 (O_668,N_49770,N_49765);
nor UO_669 (O_669,N_49513,N_49096);
nand UO_670 (O_670,N_49103,N_49004);
xnor UO_671 (O_671,N_49690,N_49108);
nand UO_672 (O_672,N_49723,N_49090);
xnor UO_673 (O_673,N_49009,N_49384);
xnor UO_674 (O_674,N_49216,N_49953);
and UO_675 (O_675,N_49145,N_49066);
xnor UO_676 (O_676,N_49463,N_49963);
xnor UO_677 (O_677,N_49958,N_49037);
or UO_678 (O_678,N_49648,N_49054);
nor UO_679 (O_679,N_49799,N_49423);
xor UO_680 (O_680,N_49610,N_49116);
nor UO_681 (O_681,N_49732,N_49691);
or UO_682 (O_682,N_49898,N_49882);
nand UO_683 (O_683,N_49958,N_49439);
xor UO_684 (O_684,N_49868,N_49343);
nand UO_685 (O_685,N_49960,N_49740);
and UO_686 (O_686,N_49323,N_49977);
nor UO_687 (O_687,N_49209,N_49306);
and UO_688 (O_688,N_49205,N_49221);
nor UO_689 (O_689,N_49070,N_49900);
or UO_690 (O_690,N_49475,N_49262);
nor UO_691 (O_691,N_49048,N_49778);
and UO_692 (O_692,N_49042,N_49196);
and UO_693 (O_693,N_49396,N_49002);
nand UO_694 (O_694,N_49831,N_49748);
xor UO_695 (O_695,N_49379,N_49887);
or UO_696 (O_696,N_49316,N_49203);
or UO_697 (O_697,N_49157,N_49513);
nor UO_698 (O_698,N_49717,N_49370);
and UO_699 (O_699,N_49508,N_49825);
nor UO_700 (O_700,N_49576,N_49419);
or UO_701 (O_701,N_49925,N_49180);
and UO_702 (O_702,N_49304,N_49754);
xor UO_703 (O_703,N_49560,N_49400);
nor UO_704 (O_704,N_49566,N_49121);
nand UO_705 (O_705,N_49750,N_49958);
nor UO_706 (O_706,N_49634,N_49565);
nor UO_707 (O_707,N_49115,N_49050);
nor UO_708 (O_708,N_49612,N_49063);
and UO_709 (O_709,N_49933,N_49965);
nor UO_710 (O_710,N_49231,N_49521);
xnor UO_711 (O_711,N_49541,N_49480);
xor UO_712 (O_712,N_49375,N_49920);
or UO_713 (O_713,N_49589,N_49500);
xor UO_714 (O_714,N_49668,N_49957);
nor UO_715 (O_715,N_49729,N_49275);
and UO_716 (O_716,N_49120,N_49865);
nor UO_717 (O_717,N_49967,N_49614);
nor UO_718 (O_718,N_49575,N_49624);
nand UO_719 (O_719,N_49523,N_49044);
or UO_720 (O_720,N_49701,N_49026);
nor UO_721 (O_721,N_49895,N_49625);
nand UO_722 (O_722,N_49632,N_49767);
nor UO_723 (O_723,N_49047,N_49875);
or UO_724 (O_724,N_49224,N_49621);
and UO_725 (O_725,N_49971,N_49281);
nor UO_726 (O_726,N_49167,N_49071);
nor UO_727 (O_727,N_49819,N_49702);
and UO_728 (O_728,N_49937,N_49328);
nand UO_729 (O_729,N_49457,N_49513);
nor UO_730 (O_730,N_49941,N_49695);
or UO_731 (O_731,N_49247,N_49705);
nand UO_732 (O_732,N_49367,N_49150);
nor UO_733 (O_733,N_49528,N_49666);
nand UO_734 (O_734,N_49785,N_49063);
xor UO_735 (O_735,N_49249,N_49154);
or UO_736 (O_736,N_49486,N_49320);
or UO_737 (O_737,N_49134,N_49256);
xnor UO_738 (O_738,N_49921,N_49594);
xor UO_739 (O_739,N_49069,N_49281);
nand UO_740 (O_740,N_49282,N_49353);
nor UO_741 (O_741,N_49909,N_49196);
xnor UO_742 (O_742,N_49848,N_49560);
or UO_743 (O_743,N_49819,N_49263);
xor UO_744 (O_744,N_49472,N_49707);
or UO_745 (O_745,N_49920,N_49704);
xor UO_746 (O_746,N_49155,N_49549);
nor UO_747 (O_747,N_49955,N_49891);
or UO_748 (O_748,N_49179,N_49933);
xor UO_749 (O_749,N_49408,N_49680);
xor UO_750 (O_750,N_49919,N_49734);
xnor UO_751 (O_751,N_49145,N_49312);
nand UO_752 (O_752,N_49936,N_49896);
or UO_753 (O_753,N_49422,N_49098);
and UO_754 (O_754,N_49877,N_49142);
and UO_755 (O_755,N_49815,N_49344);
and UO_756 (O_756,N_49805,N_49197);
nand UO_757 (O_757,N_49322,N_49544);
xor UO_758 (O_758,N_49351,N_49381);
and UO_759 (O_759,N_49884,N_49801);
and UO_760 (O_760,N_49528,N_49795);
or UO_761 (O_761,N_49107,N_49972);
or UO_762 (O_762,N_49869,N_49265);
and UO_763 (O_763,N_49492,N_49429);
xnor UO_764 (O_764,N_49619,N_49191);
nand UO_765 (O_765,N_49321,N_49977);
or UO_766 (O_766,N_49431,N_49413);
or UO_767 (O_767,N_49845,N_49903);
nor UO_768 (O_768,N_49761,N_49358);
nand UO_769 (O_769,N_49976,N_49909);
xor UO_770 (O_770,N_49967,N_49734);
xor UO_771 (O_771,N_49664,N_49560);
xor UO_772 (O_772,N_49492,N_49389);
or UO_773 (O_773,N_49817,N_49655);
or UO_774 (O_774,N_49051,N_49974);
nand UO_775 (O_775,N_49167,N_49686);
or UO_776 (O_776,N_49475,N_49158);
and UO_777 (O_777,N_49543,N_49243);
or UO_778 (O_778,N_49843,N_49013);
nor UO_779 (O_779,N_49181,N_49900);
xnor UO_780 (O_780,N_49325,N_49103);
nor UO_781 (O_781,N_49458,N_49580);
nand UO_782 (O_782,N_49662,N_49089);
nor UO_783 (O_783,N_49268,N_49042);
and UO_784 (O_784,N_49695,N_49336);
and UO_785 (O_785,N_49895,N_49296);
nand UO_786 (O_786,N_49601,N_49569);
xor UO_787 (O_787,N_49370,N_49253);
nor UO_788 (O_788,N_49386,N_49053);
and UO_789 (O_789,N_49516,N_49621);
xor UO_790 (O_790,N_49976,N_49748);
nand UO_791 (O_791,N_49696,N_49246);
and UO_792 (O_792,N_49759,N_49691);
xor UO_793 (O_793,N_49755,N_49478);
nor UO_794 (O_794,N_49528,N_49547);
or UO_795 (O_795,N_49951,N_49469);
or UO_796 (O_796,N_49288,N_49252);
and UO_797 (O_797,N_49035,N_49804);
nand UO_798 (O_798,N_49764,N_49301);
or UO_799 (O_799,N_49380,N_49419);
or UO_800 (O_800,N_49736,N_49786);
xnor UO_801 (O_801,N_49478,N_49735);
or UO_802 (O_802,N_49126,N_49870);
nor UO_803 (O_803,N_49402,N_49760);
xnor UO_804 (O_804,N_49844,N_49034);
xor UO_805 (O_805,N_49403,N_49376);
nor UO_806 (O_806,N_49724,N_49233);
nand UO_807 (O_807,N_49952,N_49757);
nor UO_808 (O_808,N_49631,N_49171);
xor UO_809 (O_809,N_49125,N_49831);
xor UO_810 (O_810,N_49769,N_49001);
nand UO_811 (O_811,N_49519,N_49561);
or UO_812 (O_812,N_49006,N_49791);
nand UO_813 (O_813,N_49086,N_49304);
or UO_814 (O_814,N_49619,N_49489);
and UO_815 (O_815,N_49741,N_49598);
nand UO_816 (O_816,N_49915,N_49107);
nor UO_817 (O_817,N_49440,N_49782);
nor UO_818 (O_818,N_49508,N_49455);
nor UO_819 (O_819,N_49735,N_49579);
nor UO_820 (O_820,N_49342,N_49214);
nand UO_821 (O_821,N_49778,N_49464);
nand UO_822 (O_822,N_49058,N_49407);
and UO_823 (O_823,N_49140,N_49373);
nor UO_824 (O_824,N_49709,N_49454);
and UO_825 (O_825,N_49849,N_49356);
nand UO_826 (O_826,N_49468,N_49695);
and UO_827 (O_827,N_49045,N_49927);
xor UO_828 (O_828,N_49938,N_49654);
xor UO_829 (O_829,N_49764,N_49707);
and UO_830 (O_830,N_49410,N_49724);
nand UO_831 (O_831,N_49750,N_49034);
and UO_832 (O_832,N_49211,N_49445);
xor UO_833 (O_833,N_49620,N_49690);
or UO_834 (O_834,N_49009,N_49955);
nand UO_835 (O_835,N_49567,N_49853);
nor UO_836 (O_836,N_49952,N_49178);
and UO_837 (O_837,N_49969,N_49816);
nand UO_838 (O_838,N_49642,N_49920);
nor UO_839 (O_839,N_49513,N_49288);
nor UO_840 (O_840,N_49299,N_49446);
xnor UO_841 (O_841,N_49344,N_49451);
nor UO_842 (O_842,N_49651,N_49451);
or UO_843 (O_843,N_49885,N_49870);
or UO_844 (O_844,N_49711,N_49520);
nand UO_845 (O_845,N_49604,N_49280);
nand UO_846 (O_846,N_49867,N_49675);
or UO_847 (O_847,N_49369,N_49543);
xnor UO_848 (O_848,N_49167,N_49646);
and UO_849 (O_849,N_49825,N_49261);
nand UO_850 (O_850,N_49721,N_49599);
xnor UO_851 (O_851,N_49045,N_49314);
or UO_852 (O_852,N_49511,N_49204);
xor UO_853 (O_853,N_49422,N_49946);
nor UO_854 (O_854,N_49389,N_49254);
xnor UO_855 (O_855,N_49404,N_49498);
xor UO_856 (O_856,N_49732,N_49847);
xnor UO_857 (O_857,N_49486,N_49287);
and UO_858 (O_858,N_49614,N_49215);
nor UO_859 (O_859,N_49685,N_49004);
nand UO_860 (O_860,N_49025,N_49673);
and UO_861 (O_861,N_49405,N_49394);
nand UO_862 (O_862,N_49398,N_49562);
and UO_863 (O_863,N_49664,N_49347);
and UO_864 (O_864,N_49165,N_49734);
and UO_865 (O_865,N_49003,N_49511);
nand UO_866 (O_866,N_49067,N_49910);
xor UO_867 (O_867,N_49808,N_49070);
or UO_868 (O_868,N_49570,N_49819);
or UO_869 (O_869,N_49164,N_49195);
or UO_870 (O_870,N_49979,N_49061);
or UO_871 (O_871,N_49534,N_49777);
and UO_872 (O_872,N_49265,N_49572);
nand UO_873 (O_873,N_49599,N_49924);
xor UO_874 (O_874,N_49137,N_49321);
nand UO_875 (O_875,N_49141,N_49191);
or UO_876 (O_876,N_49649,N_49018);
nor UO_877 (O_877,N_49101,N_49935);
xor UO_878 (O_878,N_49475,N_49816);
nand UO_879 (O_879,N_49600,N_49034);
or UO_880 (O_880,N_49749,N_49100);
xor UO_881 (O_881,N_49630,N_49567);
nand UO_882 (O_882,N_49611,N_49392);
xor UO_883 (O_883,N_49916,N_49650);
nand UO_884 (O_884,N_49334,N_49212);
and UO_885 (O_885,N_49895,N_49349);
nand UO_886 (O_886,N_49648,N_49719);
xnor UO_887 (O_887,N_49715,N_49546);
nand UO_888 (O_888,N_49211,N_49308);
and UO_889 (O_889,N_49670,N_49310);
nand UO_890 (O_890,N_49335,N_49955);
nand UO_891 (O_891,N_49905,N_49862);
nor UO_892 (O_892,N_49791,N_49485);
and UO_893 (O_893,N_49498,N_49395);
nand UO_894 (O_894,N_49374,N_49452);
xor UO_895 (O_895,N_49960,N_49103);
nand UO_896 (O_896,N_49458,N_49839);
nand UO_897 (O_897,N_49199,N_49520);
nor UO_898 (O_898,N_49608,N_49858);
and UO_899 (O_899,N_49393,N_49962);
and UO_900 (O_900,N_49993,N_49880);
nand UO_901 (O_901,N_49485,N_49578);
nand UO_902 (O_902,N_49170,N_49640);
and UO_903 (O_903,N_49756,N_49872);
nand UO_904 (O_904,N_49233,N_49383);
and UO_905 (O_905,N_49467,N_49844);
nor UO_906 (O_906,N_49662,N_49314);
nor UO_907 (O_907,N_49637,N_49870);
nand UO_908 (O_908,N_49901,N_49413);
nor UO_909 (O_909,N_49769,N_49788);
nor UO_910 (O_910,N_49652,N_49838);
nand UO_911 (O_911,N_49895,N_49923);
and UO_912 (O_912,N_49142,N_49603);
nand UO_913 (O_913,N_49796,N_49138);
xor UO_914 (O_914,N_49109,N_49660);
xor UO_915 (O_915,N_49976,N_49339);
or UO_916 (O_916,N_49929,N_49525);
and UO_917 (O_917,N_49741,N_49397);
nor UO_918 (O_918,N_49804,N_49885);
nand UO_919 (O_919,N_49072,N_49458);
or UO_920 (O_920,N_49980,N_49643);
or UO_921 (O_921,N_49199,N_49351);
nor UO_922 (O_922,N_49104,N_49208);
xnor UO_923 (O_923,N_49353,N_49229);
and UO_924 (O_924,N_49830,N_49029);
nand UO_925 (O_925,N_49731,N_49857);
nor UO_926 (O_926,N_49195,N_49320);
nor UO_927 (O_927,N_49028,N_49116);
xor UO_928 (O_928,N_49768,N_49919);
xor UO_929 (O_929,N_49018,N_49878);
xnor UO_930 (O_930,N_49797,N_49351);
nand UO_931 (O_931,N_49846,N_49397);
and UO_932 (O_932,N_49901,N_49765);
nand UO_933 (O_933,N_49244,N_49277);
and UO_934 (O_934,N_49626,N_49519);
nor UO_935 (O_935,N_49542,N_49347);
nand UO_936 (O_936,N_49259,N_49376);
or UO_937 (O_937,N_49754,N_49383);
nand UO_938 (O_938,N_49135,N_49713);
and UO_939 (O_939,N_49089,N_49586);
nand UO_940 (O_940,N_49704,N_49404);
nand UO_941 (O_941,N_49350,N_49120);
xor UO_942 (O_942,N_49892,N_49430);
and UO_943 (O_943,N_49294,N_49101);
or UO_944 (O_944,N_49324,N_49791);
or UO_945 (O_945,N_49504,N_49555);
nor UO_946 (O_946,N_49936,N_49731);
xnor UO_947 (O_947,N_49184,N_49195);
or UO_948 (O_948,N_49172,N_49212);
nand UO_949 (O_949,N_49937,N_49715);
and UO_950 (O_950,N_49371,N_49925);
or UO_951 (O_951,N_49214,N_49398);
nand UO_952 (O_952,N_49056,N_49158);
and UO_953 (O_953,N_49125,N_49721);
or UO_954 (O_954,N_49237,N_49397);
or UO_955 (O_955,N_49372,N_49821);
xnor UO_956 (O_956,N_49922,N_49401);
and UO_957 (O_957,N_49196,N_49163);
nor UO_958 (O_958,N_49989,N_49135);
nand UO_959 (O_959,N_49993,N_49043);
nand UO_960 (O_960,N_49516,N_49820);
nand UO_961 (O_961,N_49379,N_49983);
xor UO_962 (O_962,N_49209,N_49918);
or UO_963 (O_963,N_49027,N_49828);
nand UO_964 (O_964,N_49194,N_49999);
nor UO_965 (O_965,N_49771,N_49735);
nor UO_966 (O_966,N_49617,N_49796);
nand UO_967 (O_967,N_49524,N_49206);
nor UO_968 (O_968,N_49263,N_49453);
xor UO_969 (O_969,N_49417,N_49024);
nor UO_970 (O_970,N_49344,N_49470);
or UO_971 (O_971,N_49770,N_49370);
nand UO_972 (O_972,N_49698,N_49201);
or UO_973 (O_973,N_49332,N_49033);
xnor UO_974 (O_974,N_49579,N_49617);
xor UO_975 (O_975,N_49237,N_49997);
nand UO_976 (O_976,N_49152,N_49902);
and UO_977 (O_977,N_49011,N_49309);
or UO_978 (O_978,N_49740,N_49305);
or UO_979 (O_979,N_49617,N_49700);
nand UO_980 (O_980,N_49278,N_49168);
xnor UO_981 (O_981,N_49474,N_49954);
nor UO_982 (O_982,N_49898,N_49377);
or UO_983 (O_983,N_49341,N_49007);
or UO_984 (O_984,N_49092,N_49718);
nor UO_985 (O_985,N_49809,N_49804);
xor UO_986 (O_986,N_49385,N_49470);
xnor UO_987 (O_987,N_49316,N_49369);
nand UO_988 (O_988,N_49798,N_49270);
or UO_989 (O_989,N_49129,N_49516);
nor UO_990 (O_990,N_49632,N_49701);
xor UO_991 (O_991,N_49527,N_49848);
or UO_992 (O_992,N_49668,N_49748);
xor UO_993 (O_993,N_49475,N_49488);
and UO_994 (O_994,N_49779,N_49832);
nand UO_995 (O_995,N_49822,N_49474);
and UO_996 (O_996,N_49916,N_49858);
xnor UO_997 (O_997,N_49804,N_49587);
xor UO_998 (O_998,N_49526,N_49715);
nor UO_999 (O_999,N_49148,N_49065);
nand UO_1000 (O_1000,N_49807,N_49907);
nand UO_1001 (O_1001,N_49063,N_49830);
xnor UO_1002 (O_1002,N_49168,N_49846);
or UO_1003 (O_1003,N_49783,N_49017);
nand UO_1004 (O_1004,N_49752,N_49204);
or UO_1005 (O_1005,N_49529,N_49608);
xnor UO_1006 (O_1006,N_49691,N_49972);
nor UO_1007 (O_1007,N_49917,N_49040);
xor UO_1008 (O_1008,N_49504,N_49999);
nand UO_1009 (O_1009,N_49838,N_49180);
nor UO_1010 (O_1010,N_49878,N_49861);
or UO_1011 (O_1011,N_49140,N_49506);
xnor UO_1012 (O_1012,N_49418,N_49372);
nand UO_1013 (O_1013,N_49812,N_49891);
nor UO_1014 (O_1014,N_49091,N_49208);
and UO_1015 (O_1015,N_49087,N_49072);
and UO_1016 (O_1016,N_49170,N_49928);
nor UO_1017 (O_1017,N_49771,N_49887);
xor UO_1018 (O_1018,N_49789,N_49091);
xnor UO_1019 (O_1019,N_49607,N_49595);
nor UO_1020 (O_1020,N_49477,N_49320);
and UO_1021 (O_1021,N_49203,N_49058);
xnor UO_1022 (O_1022,N_49901,N_49852);
xnor UO_1023 (O_1023,N_49350,N_49759);
nor UO_1024 (O_1024,N_49503,N_49613);
xnor UO_1025 (O_1025,N_49949,N_49230);
nor UO_1026 (O_1026,N_49948,N_49452);
xnor UO_1027 (O_1027,N_49170,N_49766);
nand UO_1028 (O_1028,N_49717,N_49251);
nand UO_1029 (O_1029,N_49923,N_49560);
nand UO_1030 (O_1030,N_49134,N_49872);
or UO_1031 (O_1031,N_49381,N_49870);
or UO_1032 (O_1032,N_49662,N_49962);
and UO_1033 (O_1033,N_49712,N_49818);
nor UO_1034 (O_1034,N_49839,N_49191);
and UO_1035 (O_1035,N_49440,N_49424);
xnor UO_1036 (O_1036,N_49402,N_49011);
and UO_1037 (O_1037,N_49107,N_49651);
nand UO_1038 (O_1038,N_49528,N_49557);
xor UO_1039 (O_1039,N_49716,N_49775);
and UO_1040 (O_1040,N_49448,N_49830);
xor UO_1041 (O_1041,N_49565,N_49352);
nand UO_1042 (O_1042,N_49434,N_49486);
or UO_1043 (O_1043,N_49038,N_49092);
or UO_1044 (O_1044,N_49746,N_49890);
xnor UO_1045 (O_1045,N_49001,N_49852);
nor UO_1046 (O_1046,N_49759,N_49242);
and UO_1047 (O_1047,N_49102,N_49474);
nand UO_1048 (O_1048,N_49359,N_49342);
or UO_1049 (O_1049,N_49698,N_49614);
nand UO_1050 (O_1050,N_49304,N_49089);
xor UO_1051 (O_1051,N_49477,N_49602);
nor UO_1052 (O_1052,N_49021,N_49544);
or UO_1053 (O_1053,N_49299,N_49395);
or UO_1054 (O_1054,N_49605,N_49895);
and UO_1055 (O_1055,N_49859,N_49333);
or UO_1056 (O_1056,N_49591,N_49214);
nor UO_1057 (O_1057,N_49530,N_49228);
nand UO_1058 (O_1058,N_49990,N_49456);
nand UO_1059 (O_1059,N_49639,N_49504);
or UO_1060 (O_1060,N_49007,N_49787);
nand UO_1061 (O_1061,N_49250,N_49695);
and UO_1062 (O_1062,N_49097,N_49709);
xor UO_1063 (O_1063,N_49596,N_49811);
nor UO_1064 (O_1064,N_49622,N_49740);
and UO_1065 (O_1065,N_49961,N_49790);
nor UO_1066 (O_1066,N_49006,N_49029);
nor UO_1067 (O_1067,N_49402,N_49107);
xor UO_1068 (O_1068,N_49983,N_49414);
nand UO_1069 (O_1069,N_49986,N_49013);
nand UO_1070 (O_1070,N_49407,N_49015);
or UO_1071 (O_1071,N_49355,N_49450);
nor UO_1072 (O_1072,N_49211,N_49400);
or UO_1073 (O_1073,N_49419,N_49103);
and UO_1074 (O_1074,N_49515,N_49756);
xor UO_1075 (O_1075,N_49545,N_49758);
or UO_1076 (O_1076,N_49547,N_49301);
nor UO_1077 (O_1077,N_49234,N_49561);
and UO_1078 (O_1078,N_49934,N_49852);
or UO_1079 (O_1079,N_49849,N_49113);
xor UO_1080 (O_1080,N_49389,N_49739);
or UO_1081 (O_1081,N_49007,N_49491);
or UO_1082 (O_1082,N_49530,N_49633);
nor UO_1083 (O_1083,N_49952,N_49702);
nand UO_1084 (O_1084,N_49286,N_49553);
and UO_1085 (O_1085,N_49610,N_49399);
xor UO_1086 (O_1086,N_49722,N_49267);
nand UO_1087 (O_1087,N_49170,N_49670);
or UO_1088 (O_1088,N_49931,N_49819);
nand UO_1089 (O_1089,N_49465,N_49215);
nor UO_1090 (O_1090,N_49380,N_49064);
nand UO_1091 (O_1091,N_49594,N_49211);
and UO_1092 (O_1092,N_49161,N_49166);
nor UO_1093 (O_1093,N_49401,N_49489);
nor UO_1094 (O_1094,N_49179,N_49343);
and UO_1095 (O_1095,N_49544,N_49616);
xnor UO_1096 (O_1096,N_49186,N_49782);
and UO_1097 (O_1097,N_49310,N_49805);
nor UO_1098 (O_1098,N_49202,N_49512);
nand UO_1099 (O_1099,N_49978,N_49784);
nand UO_1100 (O_1100,N_49201,N_49883);
nor UO_1101 (O_1101,N_49504,N_49191);
xnor UO_1102 (O_1102,N_49589,N_49025);
and UO_1103 (O_1103,N_49334,N_49168);
and UO_1104 (O_1104,N_49108,N_49380);
xor UO_1105 (O_1105,N_49134,N_49221);
nor UO_1106 (O_1106,N_49075,N_49892);
or UO_1107 (O_1107,N_49287,N_49661);
and UO_1108 (O_1108,N_49692,N_49413);
xnor UO_1109 (O_1109,N_49813,N_49018);
xnor UO_1110 (O_1110,N_49860,N_49616);
and UO_1111 (O_1111,N_49678,N_49087);
and UO_1112 (O_1112,N_49370,N_49919);
nor UO_1113 (O_1113,N_49115,N_49137);
or UO_1114 (O_1114,N_49303,N_49645);
and UO_1115 (O_1115,N_49332,N_49272);
or UO_1116 (O_1116,N_49182,N_49750);
or UO_1117 (O_1117,N_49846,N_49512);
nor UO_1118 (O_1118,N_49475,N_49661);
nand UO_1119 (O_1119,N_49143,N_49355);
and UO_1120 (O_1120,N_49927,N_49043);
and UO_1121 (O_1121,N_49493,N_49665);
or UO_1122 (O_1122,N_49809,N_49268);
nor UO_1123 (O_1123,N_49577,N_49293);
nand UO_1124 (O_1124,N_49198,N_49371);
nor UO_1125 (O_1125,N_49530,N_49096);
nand UO_1126 (O_1126,N_49274,N_49256);
xnor UO_1127 (O_1127,N_49434,N_49176);
and UO_1128 (O_1128,N_49898,N_49551);
xnor UO_1129 (O_1129,N_49584,N_49890);
xnor UO_1130 (O_1130,N_49969,N_49329);
nand UO_1131 (O_1131,N_49096,N_49377);
or UO_1132 (O_1132,N_49367,N_49771);
and UO_1133 (O_1133,N_49852,N_49375);
nor UO_1134 (O_1134,N_49503,N_49764);
or UO_1135 (O_1135,N_49720,N_49731);
or UO_1136 (O_1136,N_49933,N_49466);
nor UO_1137 (O_1137,N_49786,N_49759);
or UO_1138 (O_1138,N_49930,N_49824);
and UO_1139 (O_1139,N_49000,N_49400);
nor UO_1140 (O_1140,N_49044,N_49875);
and UO_1141 (O_1141,N_49035,N_49166);
nand UO_1142 (O_1142,N_49522,N_49713);
xor UO_1143 (O_1143,N_49855,N_49939);
nor UO_1144 (O_1144,N_49534,N_49596);
nor UO_1145 (O_1145,N_49001,N_49490);
xnor UO_1146 (O_1146,N_49856,N_49479);
nand UO_1147 (O_1147,N_49137,N_49687);
or UO_1148 (O_1148,N_49905,N_49279);
and UO_1149 (O_1149,N_49824,N_49254);
and UO_1150 (O_1150,N_49183,N_49436);
nand UO_1151 (O_1151,N_49717,N_49537);
nand UO_1152 (O_1152,N_49146,N_49940);
nand UO_1153 (O_1153,N_49052,N_49389);
nand UO_1154 (O_1154,N_49632,N_49638);
and UO_1155 (O_1155,N_49869,N_49422);
nand UO_1156 (O_1156,N_49240,N_49212);
xor UO_1157 (O_1157,N_49492,N_49120);
nor UO_1158 (O_1158,N_49930,N_49597);
xor UO_1159 (O_1159,N_49506,N_49389);
nand UO_1160 (O_1160,N_49854,N_49834);
or UO_1161 (O_1161,N_49243,N_49684);
and UO_1162 (O_1162,N_49364,N_49714);
and UO_1163 (O_1163,N_49077,N_49929);
nor UO_1164 (O_1164,N_49515,N_49590);
or UO_1165 (O_1165,N_49216,N_49022);
xnor UO_1166 (O_1166,N_49525,N_49738);
nand UO_1167 (O_1167,N_49936,N_49600);
nand UO_1168 (O_1168,N_49322,N_49130);
nand UO_1169 (O_1169,N_49168,N_49186);
or UO_1170 (O_1170,N_49129,N_49840);
xor UO_1171 (O_1171,N_49621,N_49807);
nor UO_1172 (O_1172,N_49976,N_49047);
nand UO_1173 (O_1173,N_49624,N_49392);
or UO_1174 (O_1174,N_49796,N_49088);
or UO_1175 (O_1175,N_49108,N_49591);
and UO_1176 (O_1176,N_49905,N_49788);
and UO_1177 (O_1177,N_49858,N_49558);
nand UO_1178 (O_1178,N_49800,N_49097);
or UO_1179 (O_1179,N_49835,N_49977);
nor UO_1180 (O_1180,N_49996,N_49639);
xor UO_1181 (O_1181,N_49864,N_49925);
nand UO_1182 (O_1182,N_49043,N_49258);
or UO_1183 (O_1183,N_49346,N_49102);
and UO_1184 (O_1184,N_49953,N_49438);
nor UO_1185 (O_1185,N_49376,N_49712);
nor UO_1186 (O_1186,N_49084,N_49897);
and UO_1187 (O_1187,N_49411,N_49793);
nand UO_1188 (O_1188,N_49107,N_49729);
nand UO_1189 (O_1189,N_49047,N_49597);
nor UO_1190 (O_1190,N_49494,N_49359);
nor UO_1191 (O_1191,N_49716,N_49446);
or UO_1192 (O_1192,N_49503,N_49397);
nor UO_1193 (O_1193,N_49380,N_49794);
and UO_1194 (O_1194,N_49188,N_49073);
and UO_1195 (O_1195,N_49042,N_49633);
and UO_1196 (O_1196,N_49404,N_49321);
nor UO_1197 (O_1197,N_49160,N_49215);
nand UO_1198 (O_1198,N_49004,N_49725);
or UO_1199 (O_1199,N_49305,N_49002);
nor UO_1200 (O_1200,N_49573,N_49710);
nand UO_1201 (O_1201,N_49801,N_49573);
nor UO_1202 (O_1202,N_49630,N_49215);
nand UO_1203 (O_1203,N_49641,N_49656);
nor UO_1204 (O_1204,N_49516,N_49500);
nand UO_1205 (O_1205,N_49801,N_49056);
xnor UO_1206 (O_1206,N_49120,N_49493);
nor UO_1207 (O_1207,N_49521,N_49533);
nor UO_1208 (O_1208,N_49385,N_49565);
nand UO_1209 (O_1209,N_49784,N_49175);
nand UO_1210 (O_1210,N_49010,N_49958);
nor UO_1211 (O_1211,N_49913,N_49033);
xor UO_1212 (O_1212,N_49845,N_49143);
xnor UO_1213 (O_1213,N_49120,N_49873);
nand UO_1214 (O_1214,N_49509,N_49181);
nand UO_1215 (O_1215,N_49911,N_49493);
and UO_1216 (O_1216,N_49210,N_49436);
and UO_1217 (O_1217,N_49339,N_49418);
or UO_1218 (O_1218,N_49058,N_49859);
or UO_1219 (O_1219,N_49206,N_49362);
nand UO_1220 (O_1220,N_49016,N_49408);
xor UO_1221 (O_1221,N_49889,N_49487);
or UO_1222 (O_1222,N_49327,N_49403);
nor UO_1223 (O_1223,N_49797,N_49980);
and UO_1224 (O_1224,N_49641,N_49999);
or UO_1225 (O_1225,N_49525,N_49308);
nand UO_1226 (O_1226,N_49869,N_49675);
xnor UO_1227 (O_1227,N_49906,N_49019);
or UO_1228 (O_1228,N_49875,N_49406);
or UO_1229 (O_1229,N_49957,N_49170);
xor UO_1230 (O_1230,N_49358,N_49665);
nand UO_1231 (O_1231,N_49983,N_49401);
nand UO_1232 (O_1232,N_49979,N_49556);
xnor UO_1233 (O_1233,N_49402,N_49672);
xnor UO_1234 (O_1234,N_49989,N_49435);
or UO_1235 (O_1235,N_49293,N_49410);
xor UO_1236 (O_1236,N_49419,N_49299);
nor UO_1237 (O_1237,N_49376,N_49865);
xor UO_1238 (O_1238,N_49410,N_49694);
and UO_1239 (O_1239,N_49031,N_49210);
or UO_1240 (O_1240,N_49195,N_49558);
or UO_1241 (O_1241,N_49486,N_49806);
and UO_1242 (O_1242,N_49325,N_49073);
and UO_1243 (O_1243,N_49550,N_49217);
and UO_1244 (O_1244,N_49194,N_49339);
and UO_1245 (O_1245,N_49740,N_49038);
or UO_1246 (O_1246,N_49457,N_49469);
nand UO_1247 (O_1247,N_49404,N_49020);
or UO_1248 (O_1248,N_49732,N_49712);
nand UO_1249 (O_1249,N_49543,N_49638);
nand UO_1250 (O_1250,N_49023,N_49429);
nor UO_1251 (O_1251,N_49150,N_49523);
xor UO_1252 (O_1252,N_49002,N_49079);
or UO_1253 (O_1253,N_49651,N_49971);
nand UO_1254 (O_1254,N_49592,N_49341);
nand UO_1255 (O_1255,N_49763,N_49947);
or UO_1256 (O_1256,N_49746,N_49598);
nor UO_1257 (O_1257,N_49754,N_49229);
nor UO_1258 (O_1258,N_49179,N_49900);
and UO_1259 (O_1259,N_49477,N_49524);
xnor UO_1260 (O_1260,N_49200,N_49419);
nand UO_1261 (O_1261,N_49068,N_49381);
or UO_1262 (O_1262,N_49610,N_49823);
and UO_1263 (O_1263,N_49749,N_49830);
or UO_1264 (O_1264,N_49792,N_49145);
or UO_1265 (O_1265,N_49992,N_49705);
or UO_1266 (O_1266,N_49829,N_49435);
or UO_1267 (O_1267,N_49948,N_49296);
nor UO_1268 (O_1268,N_49027,N_49026);
and UO_1269 (O_1269,N_49543,N_49186);
xnor UO_1270 (O_1270,N_49820,N_49506);
nand UO_1271 (O_1271,N_49102,N_49366);
xnor UO_1272 (O_1272,N_49348,N_49279);
nand UO_1273 (O_1273,N_49982,N_49151);
nor UO_1274 (O_1274,N_49986,N_49377);
and UO_1275 (O_1275,N_49952,N_49928);
nand UO_1276 (O_1276,N_49467,N_49979);
xnor UO_1277 (O_1277,N_49634,N_49382);
nand UO_1278 (O_1278,N_49860,N_49319);
nand UO_1279 (O_1279,N_49316,N_49555);
nand UO_1280 (O_1280,N_49321,N_49347);
or UO_1281 (O_1281,N_49701,N_49455);
or UO_1282 (O_1282,N_49930,N_49342);
nand UO_1283 (O_1283,N_49285,N_49329);
nand UO_1284 (O_1284,N_49546,N_49876);
xnor UO_1285 (O_1285,N_49677,N_49523);
nor UO_1286 (O_1286,N_49434,N_49545);
xor UO_1287 (O_1287,N_49633,N_49489);
xnor UO_1288 (O_1288,N_49895,N_49443);
and UO_1289 (O_1289,N_49611,N_49706);
nor UO_1290 (O_1290,N_49817,N_49313);
and UO_1291 (O_1291,N_49580,N_49778);
or UO_1292 (O_1292,N_49397,N_49209);
or UO_1293 (O_1293,N_49012,N_49725);
or UO_1294 (O_1294,N_49474,N_49695);
and UO_1295 (O_1295,N_49325,N_49821);
nor UO_1296 (O_1296,N_49988,N_49244);
nor UO_1297 (O_1297,N_49413,N_49924);
and UO_1298 (O_1298,N_49739,N_49213);
nand UO_1299 (O_1299,N_49975,N_49478);
nand UO_1300 (O_1300,N_49641,N_49133);
nand UO_1301 (O_1301,N_49768,N_49630);
xnor UO_1302 (O_1302,N_49955,N_49031);
nand UO_1303 (O_1303,N_49746,N_49587);
and UO_1304 (O_1304,N_49745,N_49916);
xor UO_1305 (O_1305,N_49543,N_49143);
nor UO_1306 (O_1306,N_49176,N_49481);
and UO_1307 (O_1307,N_49732,N_49108);
nor UO_1308 (O_1308,N_49001,N_49782);
and UO_1309 (O_1309,N_49120,N_49217);
or UO_1310 (O_1310,N_49241,N_49291);
xor UO_1311 (O_1311,N_49318,N_49014);
xnor UO_1312 (O_1312,N_49743,N_49620);
nor UO_1313 (O_1313,N_49312,N_49872);
or UO_1314 (O_1314,N_49364,N_49107);
xnor UO_1315 (O_1315,N_49416,N_49078);
xor UO_1316 (O_1316,N_49692,N_49004);
or UO_1317 (O_1317,N_49626,N_49254);
nand UO_1318 (O_1318,N_49620,N_49972);
and UO_1319 (O_1319,N_49424,N_49809);
nor UO_1320 (O_1320,N_49538,N_49094);
nor UO_1321 (O_1321,N_49330,N_49277);
nor UO_1322 (O_1322,N_49779,N_49409);
or UO_1323 (O_1323,N_49264,N_49779);
or UO_1324 (O_1324,N_49057,N_49186);
nor UO_1325 (O_1325,N_49914,N_49649);
xnor UO_1326 (O_1326,N_49284,N_49114);
nand UO_1327 (O_1327,N_49920,N_49451);
or UO_1328 (O_1328,N_49092,N_49472);
nand UO_1329 (O_1329,N_49930,N_49507);
or UO_1330 (O_1330,N_49846,N_49413);
xnor UO_1331 (O_1331,N_49912,N_49217);
or UO_1332 (O_1332,N_49293,N_49423);
or UO_1333 (O_1333,N_49674,N_49025);
or UO_1334 (O_1334,N_49340,N_49295);
nor UO_1335 (O_1335,N_49500,N_49961);
xor UO_1336 (O_1336,N_49023,N_49216);
xnor UO_1337 (O_1337,N_49935,N_49636);
or UO_1338 (O_1338,N_49329,N_49975);
and UO_1339 (O_1339,N_49830,N_49657);
xor UO_1340 (O_1340,N_49227,N_49522);
and UO_1341 (O_1341,N_49323,N_49004);
nand UO_1342 (O_1342,N_49440,N_49155);
and UO_1343 (O_1343,N_49426,N_49612);
nand UO_1344 (O_1344,N_49091,N_49007);
nand UO_1345 (O_1345,N_49105,N_49056);
or UO_1346 (O_1346,N_49768,N_49430);
nor UO_1347 (O_1347,N_49358,N_49743);
or UO_1348 (O_1348,N_49280,N_49224);
nor UO_1349 (O_1349,N_49390,N_49382);
or UO_1350 (O_1350,N_49968,N_49756);
and UO_1351 (O_1351,N_49578,N_49562);
nand UO_1352 (O_1352,N_49093,N_49595);
nand UO_1353 (O_1353,N_49703,N_49498);
xor UO_1354 (O_1354,N_49413,N_49004);
or UO_1355 (O_1355,N_49758,N_49167);
and UO_1356 (O_1356,N_49208,N_49990);
or UO_1357 (O_1357,N_49745,N_49712);
xnor UO_1358 (O_1358,N_49852,N_49302);
and UO_1359 (O_1359,N_49771,N_49488);
and UO_1360 (O_1360,N_49705,N_49969);
and UO_1361 (O_1361,N_49409,N_49394);
or UO_1362 (O_1362,N_49750,N_49835);
nand UO_1363 (O_1363,N_49302,N_49675);
nand UO_1364 (O_1364,N_49434,N_49819);
xor UO_1365 (O_1365,N_49479,N_49412);
nor UO_1366 (O_1366,N_49325,N_49713);
xnor UO_1367 (O_1367,N_49806,N_49736);
nand UO_1368 (O_1368,N_49725,N_49285);
xnor UO_1369 (O_1369,N_49451,N_49661);
nor UO_1370 (O_1370,N_49461,N_49255);
and UO_1371 (O_1371,N_49638,N_49121);
xor UO_1372 (O_1372,N_49905,N_49779);
and UO_1373 (O_1373,N_49062,N_49082);
xor UO_1374 (O_1374,N_49840,N_49080);
nor UO_1375 (O_1375,N_49117,N_49418);
nor UO_1376 (O_1376,N_49827,N_49961);
or UO_1377 (O_1377,N_49402,N_49216);
or UO_1378 (O_1378,N_49775,N_49634);
or UO_1379 (O_1379,N_49799,N_49093);
nor UO_1380 (O_1380,N_49129,N_49759);
or UO_1381 (O_1381,N_49226,N_49053);
xnor UO_1382 (O_1382,N_49115,N_49138);
xnor UO_1383 (O_1383,N_49624,N_49539);
xnor UO_1384 (O_1384,N_49605,N_49268);
and UO_1385 (O_1385,N_49607,N_49605);
nand UO_1386 (O_1386,N_49467,N_49625);
nor UO_1387 (O_1387,N_49167,N_49941);
and UO_1388 (O_1388,N_49131,N_49473);
nand UO_1389 (O_1389,N_49531,N_49929);
nand UO_1390 (O_1390,N_49021,N_49431);
nor UO_1391 (O_1391,N_49388,N_49393);
xnor UO_1392 (O_1392,N_49421,N_49088);
nand UO_1393 (O_1393,N_49391,N_49181);
nand UO_1394 (O_1394,N_49713,N_49192);
xnor UO_1395 (O_1395,N_49358,N_49448);
xor UO_1396 (O_1396,N_49012,N_49360);
or UO_1397 (O_1397,N_49366,N_49077);
xor UO_1398 (O_1398,N_49941,N_49006);
nor UO_1399 (O_1399,N_49892,N_49475);
xnor UO_1400 (O_1400,N_49377,N_49318);
nand UO_1401 (O_1401,N_49275,N_49030);
nor UO_1402 (O_1402,N_49978,N_49212);
nand UO_1403 (O_1403,N_49656,N_49223);
and UO_1404 (O_1404,N_49791,N_49044);
xor UO_1405 (O_1405,N_49259,N_49231);
nor UO_1406 (O_1406,N_49769,N_49449);
nor UO_1407 (O_1407,N_49675,N_49270);
xnor UO_1408 (O_1408,N_49099,N_49284);
nand UO_1409 (O_1409,N_49636,N_49447);
and UO_1410 (O_1410,N_49999,N_49330);
xnor UO_1411 (O_1411,N_49490,N_49954);
nand UO_1412 (O_1412,N_49547,N_49164);
nand UO_1413 (O_1413,N_49262,N_49751);
or UO_1414 (O_1414,N_49630,N_49037);
xor UO_1415 (O_1415,N_49934,N_49915);
or UO_1416 (O_1416,N_49349,N_49445);
xnor UO_1417 (O_1417,N_49434,N_49192);
nor UO_1418 (O_1418,N_49607,N_49287);
nor UO_1419 (O_1419,N_49001,N_49458);
nand UO_1420 (O_1420,N_49125,N_49890);
xnor UO_1421 (O_1421,N_49163,N_49317);
or UO_1422 (O_1422,N_49098,N_49184);
nor UO_1423 (O_1423,N_49653,N_49403);
nand UO_1424 (O_1424,N_49411,N_49195);
nor UO_1425 (O_1425,N_49802,N_49962);
xnor UO_1426 (O_1426,N_49795,N_49564);
nor UO_1427 (O_1427,N_49420,N_49603);
nand UO_1428 (O_1428,N_49401,N_49669);
nor UO_1429 (O_1429,N_49028,N_49654);
xor UO_1430 (O_1430,N_49710,N_49667);
nor UO_1431 (O_1431,N_49998,N_49328);
nand UO_1432 (O_1432,N_49902,N_49814);
nor UO_1433 (O_1433,N_49443,N_49266);
or UO_1434 (O_1434,N_49036,N_49843);
or UO_1435 (O_1435,N_49759,N_49697);
nor UO_1436 (O_1436,N_49136,N_49793);
xnor UO_1437 (O_1437,N_49061,N_49248);
and UO_1438 (O_1438,N_49611,N_49388);
nand UO_1439 (O_1439,N_49510,N_49691);
or UO_1440 (O_1440,N_49893,N_49545);
nand UO_1441 (O_1441,N_49474,N_49772);
and UO_1442 (O_1442,N_49241,N_49741);
nor UO_1443 (O_1443,N_49614,N_49008);
and UO_1444 (O_1444,N_49090,N_49514);
nor UO_1445 (O_1445,N_49224,N_49924);
nand UO_1446 (O_1446,N_49136,N_49898);
nand UO_1447 (O_1447,N_49591,N_49470);
or UO_1448 (O_1448,N_49169,N_49760);
nand UO_1449 (O_1449,N_49988,N_49199);
nor UO_1450 (O_1450,N_49225,N_49455);
and UO_1451 (O_1451,N_49531,N_49445);
and UO_1452 (O_1452,N_49014,N_49158);
or UO_1453 (O_1453,N_49329,N_49781);
nand UO_1454 (O_1454,N_49343,N_49938);
xnor UO_1455 (O_1455,N_49634,N_49689);
nand UO_1456 (O_1456,N_49980,N_49823);
xor UO_1457 (O_1457,N_49612,N_49125);
or UO_1458 (O_1458,N_49162,N_49971);
or UO_1459 (O_1459,N_49132,N_49957);
nand UO_1460 (O_1460,N_49072,N_49437);
and UO_1461 (O_1461,N_49226,N_49338);
or UO_1462 (O_1462,N_49382,N_49235);
and UO_1463 (O_1463,N_49056,N_49214);
xor UO_1464 (O_1464,N_49076,N_49370);
or UO_1465 (O_1465,N_49611,N_49068);
nand UO_1466 (O_1466,N_49297,N_49076);
and UO_1467 (O_1467,N_49069,N_49768);
or UO_1468 (O_1468,N_49791,N_49511);
and UO_1469 (O_1469,N_49676,N_49312);
nor UO_1470 (O_1470,N_49709,N_49826);
and UO_1471 (O_1471,N_49824,N_49636);
xor UO_1472 (O_1472,N_49082,N_49557);
nor UO_1473 (O_1473,N_49149,N_49663);
xnor UO_1474 (O_1474,N_49185,N_49893);
nor UO_1475 (O_1475,N_49495,N_49197);
or UO_1476 (O_1476,N_49051,N_49909);
nor UO_1477 (O_1477,N_49582,N_49308);
or UO_1478 (O_1478,N_49160,N_49238);
or UO_1479 (O_1479,N_49990,N_49348);
and UO_1480 (O_1480,N_49702,N_49066);
and UO_1481 (O_1481,N_49282,N_49406);
nor UO_1482 (O_1482,N_49297,N_49784);
nand UO_1483 (O_1483,N_49218,N_49000);
nand UO_1484 (O_1484,N_49456,N_49783);
xor UO_1485 (O_1485,N_49024,N_49272);
and UO_1486 (O_1486,N_49012,N_49457);
or UO_1487 (O_1487,N_49952,N_49376);
xor UO_1488 (O_1488,N_49494,N_49634);
nor UO_1489 (O_1489,N_49322,N_49234);
or UO_1490 (O_1490,N_49660,N_49712);
and UO_1491 (O_1491,N_49929,N_49176);
nand UO_1492 (O_1492,N_49997,N_49675);
and UO_1493 (O_1493,N_49557,N_49451);
nor UO_1494 (O_1494,N_49079,N_49404);
xnor UO_1495 (O_1495,N_49569,N_49187);
and UO_1496 (O_1496,N_49394,N_49454);
and UO_1497 (O_1497,N_49584,N_49985);
or UO_1498 (O_1498,N_49208,N_49360);
nand UO_1499 (O_1499,N_49679,N_49964);
xnor UO_1500 (O_1500,N_49332,N_49525);
nor UO_1501 (O_1501,N_49574,N_49129);
nand UO_1502 (O_1502,N_49404,N_49844);
or UO_1503 (O_1503,N_49449,N_49799);
nand UO_1504 (O_1504,N_49087,N_49698);
xor UO_1505 (O_1505,N_49194,N_49078);
nand UO_1506 (O_1506,N_49201,N_49704);
or UO_1507 (O_1507,N_49301,N_49288);
and UO_1508 (O_1508,N_49804,N_49435);
nor UO_1509 (O_1509,N_49154,N_49425);
or UO_1510 (O_1510,N_49169,N_49632);
and UO_1511 (O_1511,N_49958,N_49267);
or UO_1512 (O_1512,N_49472,N_49918);
nor UO_1513 (O_1513,N_49627,N_49168);
or UO_1514 (O_1514,N_49818,N_49449);
or UO_1515 (O_1515,N_49755,N_49761);
nand UO_1516 (O_1516,N_49731,N_49040);
xor UO_1517 (O_1517,N_49516,N_49582);
and UO_1518 (O_1518,N_49197,N_49672);
and UO_1519 (O_1519,N_49487,N_49851);
xnor UO_1520 (O_1520,N_49446,N_49854);
xor UO_1521 (O_1521,N_49453,N_49966);
xnor UO_1522 (O_1522,N_49425,N_49175);
nor UO_1523 (O_1523,N_49222,N_49336);
nor UO_1524 (O_1524,N_49745,N_49398);
nand UO_1525 (O_1525,N_49191,N_49176);
xnor UO_1526 (O_1526,N_49433,N_49082);
and UO_1527 (O_1527,N_49901,N_49609);
and UO_1528 (O_1528,N_49076,N_49758);
nor UO_1529 (O_1529,N_49353,N_49743);
or UO_1530 (O_1530,N_49752,N_49591);
nand UO_1531 (O_1531,N_49898,N_49582);
or UO_1532 (O_1532,N_49397,N_49556);
and UO_1533 (O_1533,N_49988,N_49829);
nand UO_1534 (O_1534,N_49149,N_49440);
nor UO_1535 (O_1535,N_49771,N_49997);
and UO_1536 (O_1536,N_49291,N_49574);
and UO_1537 (O_1537,N_49659,N_49530);
xor UO_1538 (O_1538,N_49234,N_49550);
xor UO_1539 (O_1539,N_49832,N_49720);
or UO_1540 (O_1540,N_49022,N_49544);
nand UO_1541 (O_1541,N_49186,N_49705);
xnor UO_1542 (O_1542,N_49945,N_49763);
nand UO_1543 (O_1543,N_49659,N_49732);
nor UO_1544 (O_1544,N_49993,N_49144);
xnor UO_1545 (O_1545,N_49551,N_49225);
and UO_1546 (O_1546,N_49995,N_49347);
or UO_1547 (O_1547,N_49033,N_49052);
nor UO_1548 (O_1548,N_49702,N_49452);
nand UO_1549 (O_1549,N_49907,N_49164);
nand UO_1550 (O_1550,N_49796,N_49034);
nand UO_1551 (O_1551,N_49016,N_49099);
nand UO_1552 (O_1552,N_49192,N_49707);
nand UO_1553 (O_1553,N_49499,N_49985);
xor UO_1554 (O_1554,N_49362,N_49651);
nand UO_1555 (O_1555,N_49965,N_49435);
or UO_1556 (O_1556,N_49145,N_49431);
xnor UO_1557 (O_1557,N_49471,N_49603);
nor UO_1558 (O_1558,N_49791,N_49780);
nand UO_1559 (O_1559,N_49379,N_49731);
nand UO_1560 (O_1560,N_49469,N_49359);
and UO_1561 (O_1561,N_49321,N_49086);
nor UO_1562 (O_1562,N_49693,N_49564);
or UO_1563 (O_1563,N_49452,N_49522);
and UO_1564 (O_1564,N_49355,N_49765);
nor UO_1565 (O_1565,N_49388,N_49520);
nor UO_1566 (O_1566,N_49052,N_49161);
and UO_1567 (O_1567,N_49003,N_49966);
or UO_1568 (O_1568,N_49250,N_49991);
and UO_1569 (O_1569,N_49356,N_49748);
or UO_1570 (O_1570,N_49537,N_49127);
nand UO_1571 (O_1571,N_49523,N_49907);
nand UO_1572 (O_1572,N_49102,N_49229);
nand UO_1573 (O_1573,N_49697,N_49342);
or UO_1574 (O_1574,N_49427,N_49879);
nand UO_1575 (O_1575,N_49256,N_49008);
nand UO_1576 (O_1576,N_49303,N_49372);
xor UO_1577 (O_1577,N_49805,N_49769);
and UO_1578 (O_1578,N_49573,N_49654);
nand UO_1579 (O_1579,N_49784,N_49391);
or UO_1580 (O_1580,N_49079,N_49127);
and UO_1581 (O_1581,N_49216,N_49276);
nor UO_1582 (O_1582,N_49660,N_49755);
nor UO_1583 (O_1583,N_49471,N_49406);
and UO_1584 (O_1584,N_49917,N_49371);
xnor UO_1585 (O_1585,N_49085,N_49502);
nor UO_1586 (O_1586,N_49905,N_49922);
xor UO_1587 (O_1587,N_49056,N_49931);
and UO_1588 (O_1588,N_49925,N_49801);
nor UO_1589 (O_1589,N_49412,N_49708);
or UO_1590 (O_1590,N_49758,N_49902);
nand UO_1591 (O_1591,N_49870,N_49704);
nor UO_1592 (O_1592,N_49515,N_49930);
nor UO_1593 (O_1593,N_49536,N_49416);
nor UO_1594 (O_1594,N_49914,N_49068);
nand UO_1595 (O_1595,N_49251,N_49616);
nand UO_1596 (O_1596,N_49080,N_49515);
xor UO_1597 (O_1597,N_49401,N_49362);
nand UO_1598 (O_1598,N_49927,N_49875);
nand UO_1599 (O_1599,N_49742,N_49601);
or UO_1600 (O_1600,N_49437,N_49006);
xnor UO_1601 (O_1601,N_49898,N_49276);
nand UO_1602 (O_1602,N_49918,N_49407);
or UO_1603 (O_1603,N_49131,N_49559);
or UO_1604 (O_1604,N_49804,N_49028);
nor UO_1605 (O_1605,N_49234,N_49673);
or UO_1606 (O_1606,N_49842,N_49483);
and UO_1607 (O_1607,N_49807,N_49587);
and UO_1608 (O_1608,N_49417,N_49217);
xnor UO_1609 (O_1609,N_49898,N_49474);
nand UO_1610 (O_1610,N_49488,N_49888);
and UO_1611 (O_1611,N_49104,N_49641);
nand UO_1612 (O_1612,N_49910,N_49972);
nand UO_1613 (O_1613,N_49340,N_49410);
nand UO_1614 (O_1614,N_49325,N_49917);
xor UO_1615 (O_1615,N_49688,N_49764);
or UO_1616 (O_1616,N_49363,N_49847);
nand UO_1617 (O_1617,N_49237,N_49382);
nor UO_1618 (O_1618,N_49602,N_49004);
or UO_1619 (O_1619,N_49967,N_49433);
and UO_1620 (O_1620,N_49417,N_49794);
and UO_1621 (O_1621,N_49934,N_49417);
or UO_1622 (O_1622,N_49861,N_49117);
xnor UO_1623 (O_1623,N_49610,N_49779);
and UO_1624 (O_1624,N_49388,N_49290);
and UO_1625 (O_1625,N_49516,N_49960);
or UO_1626 (O_1626,N_49498,N_49889);
nor UO_1627 (O_1627,N_49762,N_49919);
or UO_1628 (O_1628,N_49375,N_49606);
xor UO_1629 (O_1629,N_49700,N_49725);
nand UO_1630 (O_1630,N_49230,N_49041);
nor UO_1631 (O_1631,N_49047,N_49815);
and UO_1632 (O_1632,N_49370,N_49214);
or UO_1633 (O_1633,N_49165,N_49163);
or UO_1634 (O_1634,N_49650,N_49483);
nor UO_1635 (O_1635,N_49262,N_49952);
or UO_1636 (O_1636,N_49978,N_49595);
and UO_1637 (O_1637,N_49640,N_49757);
nor UO_1638 (O_1638,N_49999,N_49157);
nor UO_1639 (O_1639,N_49114,N_49704);
or UO_1640 (O_1640,N_49787,N_49739);
nor UO_1641 (O_1641,N_49399,N_49975);
nand UO_1642 (O_1642,N_49507,N_49110);
xnor UO_1643 (O_1643,N_49450,N_49708);
nor UO_1644 (O_1644,N_49134,N_49361);
and UO_1645 (O_1645,N_49538,N_49841);
xor UO_1646 (O_1646,N_49109,N_49213);
xor UO_1647 (O_1647,N_49651,N_49848);
and UO_1648 (O_1648,N_49460,N_49872);
and UO_1649 (O_1649,N_49669,N_49966);
nand UO_1650 (O_1650,N_49264,N_49552);
xor UO_1651 (O_1651,N_49739,N_49584);
nand UO_1652 (O_1652,N_49819,N_49645);
and UO_1653 (O_1653,N_49216,N_49514);
or UO_1654 (O_1654,N_49318,N_49899);
nor UO_1655 (O_1655,N_49490,N_49857);
nand UO_1656 (O_1656,N_49624,N_49241);
or UO_1657 (O_1657,N_49776,N_49430);
and UO_1658 (O_1658,N_49159,N_49863);
or UO_1659 (O_1659,N_49570,N_49476);
xor UO_1660 (O_1660,N_49009,N_49237);
nor UO_1661 (O_1661,N_49271,N_49787);
or UO_1662 (O_1662,N_49204,N_49870);
xnor UO_1663 (O_1663,N_49482,N_49794);
nand UO_1664 (O_1664,N_49111,N_49049);
and UO_1665 (O_1665,N_49056,N_49250);
or UO_1666 (O_1666,N_49285,N_49164);
and UO_1667 (O_1667,N_49724,N_49513);
and UO_1668 (O_1668,N_49830,N_49301);
nor UO_1669 (O_1669,N_49563,N_49857);
xor UO_1670 (O_1670,N_49076,N_49987);
or UO_1671 (O_1671,N_49161,N_49624);
nand UO_1672 (O_1672,N_49432,N_49170);
nor UO_1673 (O_1673,N_49427,N_49061);
or UO_1674 (O_1674,N_49187,N_49761);
or UO_1675 (O_1675,N_49550,N_49527);
xor UO_1676 (O_1676,N_49912,N_49524);
xnor UO_1677 (O_1677,N_49269,N_49210);
and UO_1678 (O_1678,N_49263,N_49425);
nor UO_1679 (O_1679,N_49417,N_49961);
xnor UO_1680 (O_1680,N_49439,N_49722);
or UO_1681 (O_1681,N_49121,N_49587);
nor UO_1682 (O_1682,N_49996,N_49910);
and UO_1683 (O_1683,N_49799,N_49820);
xnor UO_1684 (O_1684,N_49413,N_49087);
xnor UO_1685 (O_1685,N_49072,N_49556);
nor UO_1686 (O_1686,N_49570,N_49548);
nor UO_1687 (O_1687,N_49559,N_49430);
and UO_1688 (O_1688,N_49423,N_49539);
xnor UO_1689 (O_1689,N_49561,N_49598);
or UO_1690 (O_1690,N_49781,N_49741);
and UO_1691 (O_1691,N_49767,N_49260);
or UO_1692 (O_1692,N_49635,N_49165);
xnor UO_1693 (O_1693,N_49112,N_49814);
nor UO_1694 (O_1694,N_49238,N_49006);
or UO_1695 (O_1695,N_49543,N_49851);
and UO_1696 (O_1696,N_49535,N_49658);
or UO_1697 (O_1697,N_49073,N_49521);
nand UO_1698 (O_1698,N_49780,N_49612);
xor UO_1699 (O_1699,N_49660,N_49268);
or UO_1700 (O_1700,N_49214,N_49712);
nor UO_1701 (O_1701,N_49196,N_49723);
or UO_1702 (O_1702,N_49947,N_49806);
or UO_1703 (O_1703,N_49783,N_49634);
or UO_1704 (O_1704,N_49784,N_49143);
and UO_1705 (O_1705,N_49436,N_49385);
xnor UO_1706 (O_1706,N_49788,N_49997);
xnor UO_1707 (O_1707,N_49824,N_49843);
xor UO_1708 (O_1708,N_49760,N_49866);
xor UO_1709 (O_1709,N_49160,N_49359);
nand UO_1710 (O_1710,N_49372,N_49279);
or UO_1711 (O_1711,N_49094,N_49461);
nor UO_1712 (O_1712,N_49766,N_49308);
and UO_1713 (O_1713,N_49711,N_49965);
or UO_1714 (O_1714,N_49480,N_49129);
and UO_1715 (O_1715,N_49596,N_49988);
nor UO_1716 (O_1716,N_49375,N_49003);
or UO_1717 (O_1717,N_49547,N_49679);
or UO_1718 (O_1718,N_49460,N_49626);
nand UO_1719 (O_1719,N_49633,N_49270);
nor UO_1720 (O_1720,N_49079,N_49616);
and UO_1721 (O_1721,N_49447,N_49301);
and UO_1722 (O_1722,N_49078,N_49569);
xnor UO_1723 (O_1723,N_49412,N_49544);
xnor UO_1724 (O_1724,N_49660,N_49742);
nand UO_1725 (O_1725,N_49963,N_49633);
xor UO_1726 (O_1726,N_49150,N_49435);
nand UO_1727 (O_1727,N_49780,N_49393);
nand UO_1728 (O_1728,N_49469,N_49139);
or UO_1729 (O_1729,N_49664,N_49903);
xnor UO_1730 (O_1730,N_49148,N_49386);
or UO_1731 (O_1731,N_49735,N_49970);
nand UO_1732 (O_1732,N_49975,N_49024);
or UO_1733 (O_1733,N_49848,N_49642);
and UO_1734 (O_1734,N_49733,N_49392);
nand UO_1735 (O_1735,N_49528,N_49854);
and UO_1736 (O_1736,N_49851,N_49314);
xnor UO_1737 (O_1737,N_49478,N_49036);
nand UO_1738 (O_1738,N_49441,N_49382);
or UO_1739 (O_1739,N_49068,N_49649);
xnor UO_1740 (O_1740,N_49199,N_49536);
or UO_1741 (O_1741,N_49331,N_49131);
and UO_1742 (O_1742,N_49539,N_49654);
and UO_1743 (O_1743,N_49918,N_49828);
or UO_1744 (O_1744,N_49988,N_49049);
xor UO_1745 (O_1745,N_49353,N_49184);
nor UO_1746 (O_1746,N_49297,N_49402);
xor UO_1747 (O_1747,N_49200,N_49232);
and UO_1748 (O_1748,N_49214,N_49355);
and UO_1749 (O_1749,N_49659,N_49267);
nor UO_1750 (O_1750,N_49875,N_49403);
xnor UO_1751 (O_1751,N_49444,N_49139);
xor UO_1752 (O_1752,N_49721,N_49993);
nor UO_1753 (O_1753,N_49165,N_49234);
xnor UO_1754 (O_1754,N_49044,N_49150);
and UO_1755 (O_1755,N_49050,N_49383);
and UO_1756 (O_1756,N_49792,N_49415);
xnor UO_1757 (O_1757,N_49975,N_49342);
nand UO_1758 (O_1758,N_49501,N_49011);
nand UO_1759 (O_1759,N_49572,N_49337);
or UO_1760 (O_1760,N_49320,N_49607);
xor UO_1761 (O_1761,N_49034,N_49381);
or UO_1762 (O_1762,N_49539,N_49988);
or UO_1763 (O_1763,N_49940,N_49758);
and UO_1764 (O_1764,N_49557,N_49032);
and UO_1765 (O_1765,N_49920,N_49123);
nand UO_1766 (O_1766,N_49502,N_49675);
nand UO_1767 (O_1767,N_49960,N_49696);
xnor UO_1768 (O_1768,N_49305,N_49564);
nand UO_1769 (O_1769,N_49309,N_49339);
nand UO_1770 (O_1770,N_49876,N_49228);
or UO_1771 (O_1771,N_49431,N_49765);
xnor UO_1772 (O_1772,N_49561,N_49802);
or UO_1773 (O_1773,N_49949,N_49404);
and UO_1774 (O_1774,N_49728,N_49984);
or UO_1775 (O_1775,N_49717,N_49607);
or UO_1776 (O_1776,N_49814,N_49809);
nand UO_1777 (O_1777,N_49998,N_49032);
or UO_1778 (O_1778,N_49804,N_49397);
nand UO_1779 (O_1779,N_49250,N_49674);
nand UO_1780 (O_1780,N_49559,N_49599);
nor UO_1781 (O_1781,N_49688,N_49282);
nand UO_1782 (O_1782,N_49941,N_49802);
nand UO_1783 (O_1783,N_49193,N_49095);
nor UO_1784 (O_1784,N_49797,N_49504);
nor UO_1785 (O_1785,N_49522,N_49493);
nor UO_1786 (O_1786,N_49748,N_49442);
nor UO_1787 (O_1787,N_49377,N_49611);
nor UO_1788 (O_1788,N_49757,N_49017);
nand UO_1789 (O_1789,N_49409,N_49222);
or UO_1790 (O_1790,N_49885,N_49462);
xor UO_1791 (O_1791,N_49343,N_49116);
xor UO_1792 (O_1792,N_49099,N_49724);
xor UO_1793 (O_1793,N_49478,N_49178);
nor UO_1794 (O_1794,N_49277,N_49317);
nand UO_1795 (O_1795,N_49723,N_49678);
and UO_1796 (O_1796,N_49894,N_49732);
and UO_1797 (O_1797,N_49225,N_49328);
nor UO_1798 (O_1798,N_49519,N_49982);
or UO_1799 (O_1799,N_49896,N_49215);
nand UO_1800 (O_1800,N_49249,N_49520);
xor UO_1801 (O_1801,N_49401,N_49269);
nor UO_1802 (O_1802,N_49075,N_49069);
and UO_1803 (O_1803,N_49015,N_49142);
nor UO_1804 (O_1804,N_49435,N_49354);
xnor UO_1805 (O_1805,N_49088,N_49863);
nand UO_1806 (O_1806,N_49548,N_49327);
or UO_1807 (O_1807,N_49657,N_49677);
or UO_1808 (O_1808,N_49286,N_49199);
nor UO_1809 (O_1809,N_49915,N_49213);
and UO_1810 (O_1810,N_49110,N_49940);
or UO_1811 (O_1811,N_49869,N_49000);
or UO_1812 (O_1812,N_49191,N_49643);
nor UO_1813 (O_1813,N_49371,N_49260);
nor UO_1814 (O_1814,N_49815,N_49716);
xor UO_1815 (O_1815,N_49117,N_49486);
nand UO_1816 (O_1816,N_49546,N_49454);
or UO_1817 (O_1817,N_49865,N_49743);
xor UO_1818 (O_1818,N_49938,N_49270);
and UO_1819 (O_1819,N_49820,N_49311);
xnor UO_1820 (O_1820,N_49084,N_49703);
nor UO_1821 (O_1821,N_49003,N_49929);
xor UO_1822 (O_1822,N_49802,N_49279);
or UO_1823 (O_1823,N_49280,N_49138);
xnor UO_1824 (O_1824,N_49006,N_49499);
xor UO_1825 (O_1825,N_49429,N_49003);
xnor UO_1826 (O_1826,N_49424,N_49202);
and UO_1827 (O_1827,N_49190,N_49925);
nand UO_1828 (O_1828,N_49868,N_49618);
and UO_1829 (O_1829,N_49032,N_49194);
xor UO_1830 (O_1830,N_49345,N_49107);
or UO_1831 (O_1831,N_49698,N_49105);
nor UO_1832 (O_1832,N_49028,N_49949);
or UO_1833 (O_1833,N_49813,N_49611);
nand UO_1834 (O_1834,N_49566,N_49453);
nand UO_1835 (O_1835,N_49629,N_49126);
and UO_1836 (O_1836,N_49231,N_49234);
xnor UO_1837 (O_1837,N_49774,N_49452);
or UO_1838 (O_1838,N_49197,N_49628);
xnor UO_1839 (O_1839,N_49877,N_49244);
and UO_1840 (O_1840,N_49486,N_49229);
and UO_1841 (O_1841,N_49834,N_49744);
nand UO_1842 (O_1842,N_49581,N_49537);
nand UO_1843 (O_1843,N_49165,N_49670);
or UO_1844 (O_1844,N_49325,N_49440);
nor UO_1845 (O_1845,N_49954,N_49276);
nor UO_1846 (O_1846,N_49744,N_49037);
xnor UO_1847 (O_1847,N_49387,N_49220);
and UO_1848 (O_1848,N_49959,N_49629);
nor UO_1849 (O_1849,N_49629,N_49702);
xnor UO_1850 (O_1850,N_49826,N_49993);
or UO_1851 (O_1851,N_49026,N_49134);
or UO_1852 (O_1852,N_49256,N_49635);
or UO_1853 (O_1853,N_49815,N_49825);
xnor UO_1854 (O_1854,N_49463,N_49020);
xnor UO_1855 (O_1855,N_49526,N_49080);
nor UO_1856 (O_1856,N_49133,N_49227);
and UO_1857 (O_1857,N_49854,N_49182);
nor UO_1858 (O_1858,N_49876,N_49855);
nand UO_1859 (O_1859,N_49512,N_49431);
or UO_1860 (O_1860,N_49310,N_49375);
and UO_1861 (O_1861,N_49359,N_49238);
and UO_1862 (O_1862,N_49201,N_49299);
and UO_1863 (O_1863,N_49523,N_49804);
or UO_1864 (O_1864,N_49771,N_49229);
nand UO_1865 (O_1865,N_49458,N_49408);
xnor UO_1866 (O_1866,N_49594,N_49302);
nand UO_1867 (O_1867,N_49375,N_49005);
nand UO_1868 (O_1868,N_49345,N_49192);
nand UO_1869 (O_1869,N_49942,N_49824);
xnor UO_1870 (O_1870,N_49412,N_49556);
nand UO_1871 (O_1871,N_49584,N_49428);
xor UO_1872 (O_1872,N_49474,N_49150);
nand UO_1873 (O_1873,N_49894,N_49446);
xnor UO_1874 (O_1874,N_49280,N_49526);
xor UO_1875 (O_1875,N_49827,N_49303);
nand UO_1876 (O_1876,N_49720,N_49696);
nand UO_1877 (O_1877,N_49718,N_49385);
or UO_1878 (O_1878,N_49353,N_49051);
nand UO_1879 (O_1879,N_49573,N_49372);
or UO_1880 (O_1880,N_49099,N_49153);
nor UO_1881 (O_1881,N_49004,N_49846);
nor UO_1882 (O_1882,N_49658,N_49485);
or UO_1883 (O_1883,N_49801,N_49101);
nor UO_1884 (O_1884,N_49129,N_49538);
nor UO_1885 (O_1885,N_49298,N_49472);
and UO_1886 (O_1886,N_49879,N_49272);
or UO_1887 (O_1887,N_49984,N_49892);
nor UO_1888 (O_1888,N_49936,N_49577);
nand UO_1889 (O_1889,N_49663,N_49791);
or UO_1890 (O_1890,N_49680,N_49419);
xnor UO_1891 (O_1891,N_49849,N_49069);
nand UO_1892 (O_1892,N_49033,N_49700);
nor UO_1893 (O_1893,N_49653,N_49010);
xor UO_1894 (O_1894,N_49450,N_49634);
xor UO_1895 (O_1895,N_49214,N_49797);
or UO_1896 (O_1896,N_49918,N_49449);
nand UO_1897 (O_1897,N_49884,N_49031);
xor UO_1898 (O_1898,N_49682,N_49869);
nor UO_1899 (O_1899,N_49923,N_49026);
nand UO_1900 (O_1900,N_49026,N_49825);
nand UO_1901 (O_1901,N_49165,N_49397);
nor UO_1902 (O_1902,N_49088,N_49733);
and UO_1903 (O_1903,N_49612,N_49773);
nor UO_1904 (O_1904,N_49869,N_49450);
nand UO_1905 (O_1905,N_49253,N_49254);
nor UO_1906 (O_1906,N_49202,N_49198);
nand UO_1907 (O_1907,N_49285,N_49431);
and UO_1908 (O_1908,N_49228,N_49907);
nand UO_1909 (O_1909,N_49985,N_49573);
and UO_1910 (O_1910,N_49058,N_49008);
xor UO_1911 (O_1911,N_49549,N_49623);
and UO_1912 (O_1912,N_49612,N_49718);
and UO_1913 (O_1913,N_49127,N_49541);
nand UO_1914 (O_1914,N_49656,N_49540);
or UO_1915 (O_1915,N_49652,N_49065);
and UO_1916 (O_1916,N_49913,N_49110);
nor UO_1917 (O_1917,N_49448,N_49544);
and UO_1918 (O_1918,N_49355,N_49820);
nand UO_1919 (O_1919,N_49961,N_49004);
and UO_1920 (O_1920,N_49155,N_49952);
nand UO_1921 (O_1921,N_49740,N_49686);
nand UO_1922 (O_1922,N_49808,N_49708);
and UO_1923 (O_1923,N_49814,N_49522);
xor UO_1924 (O_1924,N_49032,N_49120);
nor UO_1925 (O_1925,N_49652,N_49966);
nand UO_1926 (O_1926,N_49062,N_49796);
xnor UO_1927 (O_1927,N_49491,N_49690);
xor UO_1928 (O_1928,N_49176,N_49375);
or UO_1929 (O_1929,N_49643,N_49177);
xor UO_1930 (O_1930,N_49774,N_49489);
nand UO_1931 (O_1931,N_49949,N_49752);
nor UO_1932 (O_1932,N_49307,N_49639);
nand UO_1933 (O_1933,N_49555,N_49394);
nand UO_1934 (O_1934,N_49649,N_49286);
and UO_1935 (O_1935,N_49719,N_49288);
and UO_1936 (O_1936,N_49360,N_49747);
and UO_1937 (O_1937,N_49967,N_49955);
and UO_1938 (O_1938,N_49269,N_49850);
or UO_1939 (O_1939,N_49849,N_49363);
nand UO_1940 (O_1940,N_49811,N_49496);
nor UO_1941 (O_1941,N_49229,N_49026);
and UO_1942 (O_1942,N_49727,N_49025);
nand UO_1943 (O_1943,N_49457,N_49014);
xor UO_1944 (O_1944,N_49707,N_49446);
nand UO_1945 (O_1945,N_49471,N_49533);
nand UO_1946 (O_1946,N_49119,N_49389);
or UO_1947 (O_1947,N_49883,N_49647);
and UO_1948 (O_1948,N_49805,N_49355);
nand UO_1949 (O_1949,N_49332,N_49221);
or UO_1950 (O_1950,N_49146,N_49819);
nor UO_1951 (O_1951,N_49712,N_49626);
or UO_1952 (O_1952,N_49964,N_49022);
and UO_1953 (O_1953,N_49393,N_49623);
or UO_1954 (O_1954,N_49084,N_49722);
xnor UO_1955 (O_1955,N_49856,N_49310);
nand UO_1956 (O_1956,N_49912,N_49137);
xor UO_1957 (O_1957,N_49748,N_49062);
nor UO_1958 (O_1958,N_49402,N_49401);
or UO_1959 (O_1959,N_49705,N_49034);
xnor UO_1960 (O_1960,N_49312,N_49101);
or UO_1961 (O_1961,N_49784,N_49716);
and UO_1962 (O_1962,N_49352,N_49097);
or UO_1963 (O_1963,N_49618,N_49265);
xnor UO_1964 (O_1964,N_49292,N_49447);
nor UO_1965 (O_1965,N_49420,N_49587);
nand UO_1966 (O_1966,N_49695,N_49007);
nand UO_1967 (O_1967,N_49060,N_49025);
or UO_1968 (O_1968,N_49784,N_49474);
xnor UO_1969 (O_1969,N_49376,N_49990);
and UO_1970 (O_1970,N_49469,N_49118);
nor UO_1971 (O_1971,N_49511,N_49258);
or UO_1972 (O_1972,N_49384,N_49743);
nor UO_1973 (O_1973,N_49760,N_49418);
nor UO_1974 (O_1974,N_49798,N_49430);
nand UO_1975 (O_1975,N_49205,N_49240);
and UO_1976 (O_1976,N_49661,N_49942);
or UO_1977 (O_1977,N_49498,N_49305);
xor UO_1978 (O_1978,N_49331,N_49451);
or UO_1979 (O_1979,N_49890,N_49768);
nand UO_1980 (O_1980,N_49718,N_49324);
xor UO_1981 (O_1981,N_49365,N_49439);
and UO_1982 (O_1982,N_49662,N_49905);
xor UO_1983 (O_1983,N_49650,N_49911);
nor UO_1984 (O_1984,N_49090,N_49534);
nor UO_1985 (O_1985,N_49124,N_49014);
and UO_1986 (O_1986,N_49997,N_49959);
nand UO_1987 (O_1987,N_49959,N_49666);
nand UO_1988 (O_1988,N_49670,N_49936);
xnor UO_1989 (O_1989,N_49766,N_49966);
or UO_1990 (O_1990,N_49147,N_49249);
xnor UO_1991 (O_1991,N_49525,N_49474);
nand UO_1992 (O_1992,N_49389,N_49926);
and UO_1993 (O_1993,N_49269,N_49579);
nor UO_1994 (O_1994,N_49633,N_49103);
or UO_1995 (O_1995,N_49591,N_49887);
or UO_1996 (O_1996,N_49710,N_49070);
xnor UO_1997 (O_1997,N_49286,N_49039);
or UO_1998 (O_1998,N_49281,N_49768);
nor UO_1999 (O_1999,N_49948,N_49638);
nand UO_2000 (O_2000,N_49920,N_49061);
xor UO_2001 (O_2001,N_49894,N_49820);
and UO_2002 (O_2002,N_49454,N_49873);
xnor UO_2003 (O_2003,N_49027,N_49456);
xnor UO_2004 (O_2004,N_49014,N_49863);
or UO_2005 (O_2005,N_49506,N_49088);
xnor UO_2006 (O_2006,N_49288,N_49404);
or UO_2007 (O_2007,N_49940,N_49515);
nand UO_2008 (O_2008,N_49070,N_49463);
xnor UO_2009 (O_2009,N_49676,N_49746);
nand UO_2010 (O_2010,N_49504,N_49556);
or UO_2011 (O_2011,N_49381,N_49610);
nor UO_2012 (O_2012,N_49822,N_49721);
or UO_2013 (O_2013,N_49773,N_49112);
nand UO_2014 (O_2014,N_49703,N_49880);
and UO_2015 (O_2015,N_49766,N_49860);
xor UO_2016 (O_2016,N_49983,N_49125);
and UO_2017 (O_2017,N_49711,N_49845);
xor UO_2018 (O_2018,N_49493,N_49850);
or UO_2019 (O_2019,N_49048,N_49699);
and UO_2020 (O_2020,N_49353,N_49612);
xor UO_2021 (O_2021,N_49376,N_49859);
or UO_2022 (O_2022,N_49951,N_49660);
nor UO_2023 (O_2023,N_49489,N_49332);
or UO_2024 (O_2024,N_49540,N_49698);
xor UO_2025 (O_2025,N_49724,N_49335);
nor UO_2026 (O_2026,N_49283,N_49519);
and UO_2027 (O_2027,N_49421,N_49132);
or UO_2028 (O_2028,N_49644,N_49198);
or UO_2029 (O_2029,N_49727,N_49511);
xnor UO_2030 (O_2030,N_49131,N_49887);
nor UO_2031 (O_2031,N_49878,N_49732);
and UO_2032 (O_2032,N_49300,N_49817);
nand UO_2033 (O_2033,N_49362,N_49760);
or UO_2034 (O_2034,N_49735,N_49247);
nand UO_2035 (O_2035,N_49354,N_49151);
and UO_2036 (O_2036,N_49866,N_49112);
or UO_2037 (O_2037,N_49093,N_49958);
and UO_2038 (O_2038,N_49642,N_49944);
nand UO_2039 (O_2039,N_49749,N_49849);
nor UO_2040 (O_2040,N_49058,N_49894);
nand UO_2041 (O_2041,N_49915,N_49872);
nand UO_2042 (O_2042,N_49519,N_49342);
nand UO_2043 (O_2043,N_49545,N_49586);
and UO_2044 (O_2044,N_49634,N_49492);
xnor UO_2045 (O_2045,N_49550,N_49757);
and UO_2046 (O_2046,N_49527,N_49147);
xnor UO_2047 (O_2047,N_49692,N_49850);
nand UO_2048 (O_2048,N_49791,N_49624);
and UO_2049 (O_2049,N_49369,N_49088);
or UO_2050 (O_2050,N_49411,N_49827);
nor UO_2051 (O_2051,N_49931,N_49016);
nor UO_2052 (O_2052,N_49924,N_49237);
nand UO_2053 (O_2053,N_49301,N_49667);
xor UO_2054 (O_2054,N_49597,N_49594);
or UO_2055 (O_2055,N_49774,N_49941);
or UO_2056 (O_2056,N_49576,N_49953);
and UO_2057 (O_2057,N_49957,N_49778);
xor UO_2058 (O_2058,N_49290,N_49280);
and UO_2059 (O_2059,N_49684,N_49699);
and UO_2060 (O_2060,N_49621,N_49962);
nor UO_2061 (O_2061,N_49835,N_49299);
nand UO_2062 (O_2062,N_49555,N_49567);
xnor UO_2063 (O_2063,N_49649,N_49987);
nor UO_2064 (O_2064,N_49422,N_49281);
xor UO_2065 (O_2065,N_49753,N_49740);
or UO_2066 (O_2066,N_49714,N_49062);
or UO_2067 (O_2067,N_49355,N_49823);
or UO_2068 (O_2068,N_49295,N_49684);
xnor UO_2069 (O_2069,N_49099,N_49559);
nor UO_2070 (O_2070,N_49727,N_49514);
xnor UO_2071 (O_2071,N_49013,N_49099);
nand UO_2072 (O_2072,N_49281,N_49538);
nand UO_2073 (O_2073,N_49478,N_49219);
and UO_2074 (O_2074,N_49726,N_49143);
nand UO_2075 (O_2075,N_49480,N_49155);
and UO_2076 (O_2076,N_49422,N_49008);
nand UO_2077 (O_2077,N_49503,N_49146);
or UO_2078 (O_2078,N_49876,N_49320);
and UO_2079 (O_2079,N_49992,N_49896);
xor UO_2080 (O_2080,N_49909,N_49926);
nor UO_2081 (O_2081,N_49675,N_49016);
nor UO_2082 (O_2082,N_49135,N_49668);
nand UO_2083 (O_2083,N_49751,N_49231);
nor UO_2084 (O_2084,N_49505,N_49622);
nand UO_2085 (O_2085,N_49247,N_49628);
and UO_2086 (O_2086,N_49079,N_49691);
nand UO_2087 (O_2087,N_49462,N_49096);
nor UO_2088 (O_2088,N_49725,N_49745);
nor UO_2089 (O_2089,N_49233,N_49765);
and UO_2090 (O_2090,N_49829,N_49083);
nor UO_2091 (O_2091,N_49446,N_49941);
nor UO_2092 (O_2092,N_49312,N_49450);
nand UO_2093 (O_2093,N_49429,N_49763);
nor UO_2094 (O_2094,N_49421,N_49430);
or UO_2095 (O_2095,N_49038,N_49785);
and UO_2096 (O_2096,N_49128,N_49302);
nand UO_2097 (O_2097,N_49147,N_49294);
xnor UO_2098 (O_2098,N_49927,N_49824);
and UO_2099 (O_2099,N_49414,N_49542);
nand UO_2100 (O_2100,N_49932,N_49214);
nand UO_2101 (O_2101,N_49287,N_49573);
nand UO_2102 (O_2102,N_49171,N_49470);
and UO_2103 (O_2103,N_49624,N_49227);
nand UO_2104 (O_2104,N_49694,N_49343);
nand UO_2105 (O_2105,N_49927,N_49412);
and UO_2106 (O_2106,N_49618,N_49786);
xnor UO_2107 (O_2107,N_49788,N_49576);
xnor UO_2108 (O_2108,N_49808,N_49669);
nor UO_2109 (O_2109,N_49982,N_49190);
xor UO_2110 (O_2110,N_49268,N_49069);
nor UO_2111 (O_2111,N_49329,N_49773);
or UO_2112 (O_2112,N_49879,N_49649);
xnor UO_2113 (O_2113,N_49736,N_49694);
and UO_2114 (O_2114,N_49770,N_49618);
nand UO_2115 (O_2115,N_49315,N_49733);
nor UO_2116 (O_2116,N_49207,N_49438);
nor UO_2117 (O_2117,N_49379,N_49974);
and UO_2118 (O_2118,N_49004,N_49098);
and UO_2119 (O_2119,N_49836,N_49936);
xor UO_2120 (O_2120,N_49991,N_49015);
xor UO_2121 (O_2121,N_49838,N_49034);
and UO_2122 (O_2122,N_49025,N_49179);
nand UO_2123 (O_2123,N_49760,N_49974);
xor UO_2124 (O_2124,N_49402,N_49286);
nor UO_2125 (O_2125,N_49260,N_49321);
and UO_2126 (O_2126,N_49995,N_49409);
and UO_2127 (O_2127,N_49483,N_49062);
nand UO_2128 (O_2128,N_49584,N_49550);
xor UO_2129 (O_2129,N_49707,N_49967);
nand UO_2130 (O_2130,N_49951,N_49754);
xor UO_2131 (O_2131,N_49218,N_49470);
nand UO_2132 (O_2132,N_49045,N_49770);
nor UO_2133 (O_2133,N_49116,N_49806);
xnor UO_2134 (O_2134,N_49059,N_49335);
or UO_2135 (O_2135,N_49785,N_49504);
nor UO_2136 (O_2136,N_49680,N_49481);
and UO_2137 (O_2137,N_49045,N_49063);
or UO_2138 (O_2138,N_49617,N_49031);
nor UO_2139 (O_2139,N_49950,N_49537);
nand UO_2140 (O_2140,N_49680,N_49673);
or UO_2141 (O_2141,N_49433,N_49801);
nor UO_2142 (O_2142,N_49173,N_49301);
and UO_2143 (O_2143,N_49733,N_49691);
nand UO_2144 (O_2144,N_49691,N_49173);
and UO_2145 (O_2145,N_49018,N_49987);
nor UO_2146 (O_2146,N_49650,N_49320);
nor UO_2147 (O_2147,N_49455,N_49390);
or UO_2148 (O_2148,N_49895,N_49209);
nor UO_2149 (O_2149,N_49725,N_49825);
and UO_2150 (O_2150,N_49447,N_49223);
nand UO_2151 (O_2151,N_49378,N_49890);
nor UO_2152 (O_2152,N_49667,N_49452);
nand UO_2153 (O_2153,N_49901,N_49114);
nand UO_2154 (O_2154,N_49006,N_49005);
xor UO_2155 (O_2155,N_49053,N_49441);
nand UO_2156 (O_2156,N_49110,N_49328);
xnor UO_2157 (O_2157,N_49904,N_49385);
nor UO_2158 (O_2158,N_49935,N_49142);
and UO_2159 (O_2159,N_49840,N_49585);
or UO_2160 (O_2160,N_49361,N_49241);
xnor UO_2161 (O_2161,N_49113,N_49986);
or UO_2162 (O_2162,N_49236,N_49708);
xor UO_2163 (O_2163,N_49302,N_49766);
and UO_2164 (O_2164,N_49390,N_49364);
xor UO_2165 (O_2165,N_49576,N_49037);
nand UO_2166 (O_2166,N_49819,N_49782);
xnor UO_2167 (O_2167,N_49490,N_49572);
nor UO_2168 (O_2168,N_49204,N_49323);
xnor UO_2169 (O_2169,N_49871,N_49544);
and UO_2170 (O_2170,N_49977,N_49155);
nor UO_2171 (O_2171,N_49267,N_49157);
nor UO_2172 (O_2172,N_49806,N_49937);
and UO_2173 (O_2173,N_49761,N_49645);
nand UO_2174 (O_2174,N_49836,N_49409);
xor UO_2175 (O_2175,N_49018,N_49399);
nand UO_2176 (O_2176,N_49966,N_49569);
or UO_2177 (O_2177,N_49913,N_49513);
and UO_2178 (O_2178,N_49740,N_49818);
or UO_2179 (O_2179,N_49807,N_49264);
nor UO_2180 (O_2180,N_49702,N_49766);
nand UO_2181 (O_2181,N_49417,N_49584);
or UO_2182 (O_2182,N_49518,N_49375);
or UO_2183 (O_2183,N_49664,N_49094);
nand UO_2184 (O_2184,N_49103,N_49775);
and UO_2185 (O_2185,N_49361,N_49686);
and UO_2186 (O_2186,N_49538,N_49224);
xnor UO_2187 (O_2187,N_49927,N_49973);
and UO_2188 (O_2188,N_49586,N_49551);
nand UO_2189 (O_2189,N_49359,N_49384);
or UO_2190 (O_2190,N_49877,N_49932);
xor UO_2191 (O_2191,N_49755,N_49368);
and UO_2192 (O_2192,N_49211,N_49582);
xnor UO_2193 (O_2193,N_49239,N_49456);
or UO_2194 (O_2194,N_49730,N_49060);
or UO_2195 (O_2195,N_49205,N_49881);
nor UO_2196 (O_2196,N_49641,N_49907);
nor UO_2197 (O_2197,N_49205,N_49047);
xnor UO_2198 (O_2198,N_49928,N_49523);
nor UO_2199 (O_2199,N_49493,N_49214);
xnor UO_2200 (O_2200,N_49864,N_49280);
and UO_2201 (O_2201,N_49376,N_49313);
and UO_2202 (O_2202,N_49562,N_49301);
and UO_2203 (O_2203,N_49435,N_49526);
xnor UO_2204 (O_2204,N_49980,N_49327);
xnor UO_2205 (O_2205,N_49224,N_49707);
nand UO_2206 (O_2206,N_49799,N_49132);
xnor UO_2207 (O_2207,N_49528,N_49871);
nand UO_2208 (O_2208,N_49475,N_49205);
nand UO_2209 (O_2209,N_49072,N_49499);
xnor UO_2210 (O_2210,N_49131,N_49432);
nand UO_2211 (O_2211,N_49902,N_49589);
and UO_2212 (O_2212,N_49313,N_49701);
nand UO_2213 (O_2213,N_49620,N_49187);
nand UO_2214 (O_2214,N_49028,N_49764);
and UO_2215 (O_2215,N_49491,N_49923);
nor UO_2216 (O_2216,N_49377,N_49472);
nor UO_2217 (O_2217,N_49936,N_49081);
xor UO_2218 (O_2218,N_49768,N_49623);
xnor UO_2219 (O_2219,N_49319,N_49113);
or UO_2220 (O_2220,N_49602,N_49773);
xor UO_2221 (O_2221,N_49016,N_49701);
nand UO_2222 (O_2222,N_49755,N_49426);
nor UO_2223 (O_2223,N_49938,N_49801);
and UO_2224 (O_2224,N_49454,N_49551);
or UO_2225 (O_2225,N_49537,N_49440);
nor UO_2226 (O_2226,N_49620,N_49175);
xor UO_2227 (O_2227,N_49964,N_49241);
nand UO_2228 (O_2228,N_49477,N_49833);
nor UO_2229 (O_2229,N_49547,N_49747);
nor UO_2230 (O_2230,N_49885,N_49504);
nand UO_2231 (O_2231,N_49610,N_49368);
or UO_2232 (O_2232,N_49573,N_49429);
nand UO_2233 (O_2233,N_49782,N_49199);
or UO_2234 (O_2234,N_49067,N_49439);
nor UO_2235 (O_2235,N_49804,N_49196);
or UO_2236 (O_2236,N_49528,N_49841);
and UO_2237 (O_2237,N_49465,N_49577);
xnor UO_2238 (O_2238,N_49842,N_49131);
xor UO_2239 (O_2239,N_49182,N_49428);
nor UO_2240 (O_2240,N_49611,N_49167);
nand UO_2241 (O_2241,N_49626,N_49237);
or UO_2242 (O_2242,N_49536,N_49902);
xor UO_2243 (O_2243,N_49577,N_49529);
xor UO_2244 (O_2244,N_49530,N_49461);
and UO_2245 (O_2245,N_49369,N_49697);
and UO_2246 (O_2246,N_49699,N_49468);
xnor UO_2247 (O_2247,N_49154,N_49213);
or UO_2248 (O_2248,N_49556,N_49332);
or UO_2249 (O_2249,N_49624,N_49671);
nor UO_2250 (O_2250,N_49723,N_49325);
or UO_2251 (O_2251,N_49545,N_49716);
nand UO_2252 (O_2252,N_49856,N_49021);
and UO_2253 (O_2253,N_49594,N_49813);
nand UO_2254 (O_2254,N_49529,N_49104);
xnor UO_2255 (O_2255,N_49542,N_49439);
nor UO_2256 (O_2256,N_49199,N_49454);
and UO_2257 (O_2257,N_49707,N_49943);
nor UO_2258 (O_2258,N_49290,N_49733);
nand UO_2259 (O_2259,N_49194,N_49200);
nor UO_2260 (O_2260,N_49980,N_49375);
nor UO_2261 (O_2261,N_49694,N_49504);
nor UO_2262 (O_2262,N_49525,N_49846);
and UO_2263 (O_2263,N_49207,N_49126);
and UO_2264 (O_2264,N_49730,N_49916);
and UO_2265 (O_2265,N_49078,N_49242);
xor UO_2266 (O_2266,N_49166,N_49450);
nand UO_2267 (O_2267,N_49027,N_49174);
or UO_2268 (O_2268,N_49629,N_49762);
nand UO_2269 (O_2269,N_49477,N_49538);
nand UO_2270 (O_2270,N_49281,N_49929);
nor UO_2271 (O_2271,N_49635,N_49065);
nor UO_2272 (O_2272,N_49763,N_49059);
or UO_2273 (O_2273,N_49181,N_49970);
and UO_2274 (O_2274,N_49416,N_49099);
or UO_2275 (O_2275,N_49630,N_49277);
nand UO_2276 (O_2276,N_49061,N_49426);
nand UO_2277 (O_2277,N_49423,N_49665);
xor UO_2278 (O_2278,N_49281,N_49295);
and UO_2279 (O_2279,N_49211,N_49210);
and UO_2280 (O_2280,N_49366,N_49384);
xnor UO_2281 (O_2281,N_49348,N_49301);
nor UO_2282 (O_2282,N_49621,N_49759);
or UO_2283 (O_2283,N_49864,N_49119);
nand UO_2284 (O_2284,N_49514,N_49403);
or UO_2285 (O_2285,N_49251,N_49974);
nor UO_2286 (O_2286,N_49765,N_49906);
nor UO_2287 (O_2287,N_49874,N_49662);
xnor UO_2288 (O_2288,N_49987,N_49053);
and UO_2289 (O_2289,N_49896,N_49801);
and UO_2290 (O_2290,N_49835,N_49857);
and UO_2291 (O_2291,N_49491,N_49273);
nor UO_2292 (O_2292,N_49764,N_49983);
or UO_2293 (O_2293,N_49803,N_49868);
or UO_2294 (O_2294,N_49852,N_49074);
and UO_2295 (O_2295,N_49630,N_49411);
nor UO_2296 (O_2296,N_49520,N_49891);
and UO_2297 (O_2297,N_49434,N_49974);
and UO_2298 (O_2298,N_49001,N_49049);
and UO_2299 (O_2299,N_49970,N_49589);
or UO_2300 (O_2300,N_49645,N_49666);
xor UO_2301 (O_2301,N_49863,N_49700);
nand UO_2302 (O_2302,N_49962,N_49453);
nor UO_2303 (O_2303,N_49194,N_49888);
nor UO_2304 (O_2304,N_49597,N_49704);
or UO_2305 (O_2305,N_49279,N_49704);
and UO_2306 (O_2306,N_49950,N_49837);
or UO_2307 (O_2307,N_49067,N_49083);
and UO_2308 (O_2308,N_49746,N_49850);
or UO_2309 (O_2309,N_49301,N_49161);
xnor UO_2310 (O_2310,N_49284,N_49707);
xor UO_2311 (O_2311,N_49814,N_49363);
nand UO_2312 (O_2312,N_49212,N_49300);
nand UO_2313 (O_2313,N_49294,N_49208);
and UO_2314 (O_2314,N_49048,N_49581);
nor UO_2315 (O_2315,N_49612,N_49306);
xor UO_2316 (O_2316,N_49654,N_49695);
and UO_2317 (O_2317,N_49752,N_49104);
nor UO_2318 (O_2318,N_49779,N_49493);
nor UO_2319 (O_2319,N_49434,N_49189);
nand UO_2320 (O_2320,N_49602,N_49524);
nand UO_2321 (O_2321,N_49003,N_49049);
and UO_2322 (O_2322,N_49257,N_49778);
or UO_2323 (O_2323,N_49591,N_49365);
and UO_2324 (O_2324,N_49247,N_49606);
xor UO_2325 (O_2325,N_49691,N_49472);
xnor UO_2326 (O_2326,N_49275,N_49319);
and UO_2327 (O_2327,N_49185,N_49045);
xor UO_2328 (O_2328,N_49417,N_49013);
nor UO_2329 (O_2329,N_49861,N_49580);
xnor UO_2330 (O_2330,N_49714,N_49485);
or UO_2331 (O_2331,N_49709,N_49927);
nand UO_2332 (O_2332,N_49884,N_49775);
nand UO_2333 (O_2333,N_49770,N_49108);
and UO_2334 (O_2334,N_49158,N_49738);
or UO_2335 (O_2335,N_49463,N_49537);
and UO_2336 (O_2336,N_49996,N_49927);
xnor UO_2337 (O_2337,N_49668,N_49890);
or UO_2338 (O_2338,N_49186,N_49166);
xor UO_2339 (O_2339,N_49121,N_49632);
xnor UO_2340 (O_2340,N_49208,N_49522);
or UO_2341 (O_2341,N_49976,N_49063);
and UO_2342 (O_2342,N_49069,N_49900);
xor UO_2343 (O_2343,N_49865,N_49660);
xnor UO_2344 (O_2344,N_49760,N_49562);
and UO_2345 (O_2345,N_49855,N_49084);
xnor UO_2346 (O_2346,N_49959,N_49252);
and UO_2347 (O_2347,N_49629,N_49157);
or UO_2348 (O_2348,N_49779,N_49006);
xor UO_2349 (O_2349,N_49652,N_49211);
xor UO_2350 (O_2350,N_49519,N_49044);
xor UO_2351 (O_2351,N_49943,N_49739);
or UO_2352 (O_2352,N_49173,N_49425);
xnor UO_2353 (O_2353,N_49420,N_49418);
nor UO_2354 (O_2354,N_49008,N_49862);
xor UO_2355 (O_2355,N_49596,N_49532);
nand UO_2356 (O_2356,N_49996,N_49263);
xnor UO_2357 (O_2357,N_49864,N_49293);
nor UO_2358 (O_2358,N_49943,N_49364);
or UO_2359 (O_2359,N_49982,N_49762);
and UO_2360 (O_2360,N_49103,N_49780);
and UO_2361 (O_2361,N_49693,N_49007);
and UO_2362 (O_2362,N_49582,N_49643);
and UO_2363 (O_2363,N_49007,N_49233);
xor UO_2364 (O_2364,N_49715,N_49423);
and UO_2365 (O_2365,N_49421,N_49288);
and UO_2366 (O_2366,N_49398,N_49196);
or UO_2367 (O_2367,N_49241,N_49938);
nor UO_2368 (O_2368,N_49702,N_49659);
nor UO_2369 (O_2369,N_49344,N_49208);
nor UO_2370 (O_2370,N_49483,N_49241);
xnor UO_2371 (O_2371,N_49263,N_49740);
and UO_2372 (O_2372,N_49982,N_49069);
nand UO_2373 (O_2373,N_49976,N_49430);
or UO_2374 (O_2374,N_49721,N_49064);
and UO_2375 (O_2375,N_49478,N_49206);
nor UO_2376 (O_2376,N_49003,N_49247);
nand UO_2377 (O_2377,N_49931,N_49540);
or UO_2378 (O_2378,N_49278,N_49197);
nor UO_2379 (O_2379,N_49612,N_49866);
and UO_2380 (O_2380,N_49936,N_49257);
and UO_2381 (O_2381,N_49251,N_49380);
and UO_2382 (O_2382,N_49155,N_49705);
and UO_2383 (O_2383,N_49141,N_49309);
xor UO_2384 (O_2384,N_49829,N_49979);
or UO_2385 (O_2385,N_49319,N_49697);
xnor UO_2386 (O_2386,N_49765,N_49269);
and UO_2387 (O_2387,N_49052,N_49036);
nand UO_2388 (O_2388,N_49971,N_49932);
or UO_2389 (O_2389,N_49227,N_49611);
or UO_2390 (O_2390,N_49355,N_49803);
nand UO_2391 (O_2391,N_49637,N_49405);
nor UO_2392 (O_2392,N_49198,N_49370);
or UO_2393 (O_2393,N_49533,N_49208);
and UO_2394 (O_2394,N_49468,N_49832);
or UO_2395 (O_2395,N_49102,N_49660);
nor UO_2396 (O_2396,N_49387,N_49963);
xor UO_2397 (O_2397,N_49647,N_49963);
and UO_2398 (O_2398,N_49042,N_49592);
nor UO_2399 (O_2399,N_49407,N_49103);
nand UO_2400 (O_2400,N_49629,N_49801);
nand UO_2401 (O_2401,N_49278,N_49003);
or UO_2402 (O_2402,N_49037,N_49586);
xnor UO_2403 (O_2403,N_49336,N_49153);
nand UO_2404 (O_2404,N_49428,N_49843);
nand UO_2405 (O_2405,N_49773,N_49755);
nor UO_2406 (O_2406,N_49419,N_49046);
xor UO_2407 (O_2407,N_49874,N_49324);
xor UO_2408 (O_2408,N_49723,N_49549);
xnor UO_2409 (O_2409,N_49112,N_49895);
or UO_2410 (O_2410,N_49771,N_49658);
nor UO_2411 (O_2411,N_49220,N_49413);
or UO_2412 (O_2412,N_49783,N_49051);
nor UO_2413 (O_2413,N_49784,N_49425);
nor UO_2414 (O_2414,N_49115,N_49999);
xnor UO_2415 (O_2415,N_49855,N_49606);
or UO_2416 (O_2416,N_49008,N_49833);
nor UO_2417 (O_2417,N_49915,N_49893);
nand UO_2418 (O_2418,N_49044,N_49518);
nor UO_2419 (O_2419,N_49150,N_49817);
nand UO_2420 (O_2420,N_49077,N_49206);
nor UO_2421 (O_2421,N_49300,N_49314);
or UO_2422 (O_2422,N_49423,N_49413);
and UO_2423 (O_2423,N_49749,N_49857);
nor UO_2424 (O_2424,N_49227,N_49200);
nor UO_2425 (O_2425,N_49124,N_49500);
nor UO_2426 (O_2426,N_49248,N_49046);
nand UO_2427 (O_2427,N_49403,N_49916);
and UO_2428 (O_2428,N_49864,N_49961);
nor UO_2429 (O_2429,N_49642,N_49902);
nand UO_2430 (O_2430,N_49941,N_49197);
xor UO_2431 (O_2431,N_49110,N_49606);
nor UO_2432 (O_2432,N_49085,N_49842);
or UO_2433 (O_2433,N_49080,N_49841);
and UO_2434 (O_2434,N_49967,N_49345);
and UO_2435 (O_2435,N_49323,N_49949);
xnor UO_2436 (O_2436,N_49979,N_49660);
nand UO_2437 (O_2437,N_49844,N_49324);
nand UO_2438 (O_2438,N_49409,N_49823);
and UO_2439 (O_2439,N_49173,N_49556);
or UO_2440 (O_2440,N_49337,N_49529);
or UO_2441 (O_2441,N_49355,N_49398);
and UO_2442 (O_2442,N_49719,N_49877);
xnor UO_2443 (O_2443,N_49057,N_49430);
nand UO_2444 (O_2444,N_49623,N_49104);
and UO_2445 (O_2445,N_49277,N_49273);
nor UO_2446 (O_2446,N_49851,N_49209);
and UO_2447 (O_2447,N_49194,N_49099);
nand UO_2448 (O_2448,N_49224,N_49717);
nor UO_2449 (O_2449,N_49001,N_49179);
and UO_2450 (O_2450,N_49773,N_49687);
xor UO_2451 (O_2451,N_49534,N_49266);
and UO_2452 (O_2452,N_49949,N_49979);
xor UO_2453 (O_2453,N_49173,N_49015);
and UO_2454 (O_2454,N_49958,N_49559);
nor UO_2455 (O_2455,N_49218,N_49124);
xor UO_2456 (O_2456,N_49232,N_49943);
or UO_2457 (O_2457,N_49887,N_49021);
or UO_2458 (O_2458,N_49088,N_49321);
and UO_2459 (O_2459,N_49982,N_49562);
xnor UO_2460 (O_2460,N_49039,N_49803);
nor UO_2461 (O_2461,N_49525,N_49754);
and UO_2462 (O_2462,N_49144,N_49249);
xnor UO_2463 (O_2463,N_49455,N_49457);
nand UO_2464 (O_2464,N_49326,N_49983);
xor UO_2465 (O_2465,N_49116,N_49504);
xnor UO_2466 (O_2466,N_49907,N_49297);
nor UO_2467 (O_2467,N_49145,N_49547);
and UO_2468 (O_2468,N_49163,N_49264);
xnor UO_2469 (O_2469,N_49947,N_49108);
or UO_2470 (O_2470,N_49202,N_49361);
xnor UO_2471 (O_2471,N_49684,N_49969);
and UO_2472 (O_2472,N_49591,N_49520);
nand UO_2473 (O_2473,N_49612,N_49668);
nand UO_2474 (O_2474,N_49017,N_49527);
nor UO_2475 (O_2475,N_49456,N_49170);
or UO_2476 (O_2476,N_49178,N_49350);
xor UO_2477 (O_2477,N_49589,N_49922);
nand UO_2478 (O_2478,N_49838,N_49114);
or UO_2479 (O_2479,N_49325,N_49248);
or UO_2480 (O_2480,N_49718,N_49714);
xor UO_2481 (O_2481,N_49123,N_49554);
xor UO_2482 (O_2482,N_49573,N_49414);
or UO_2483 (O_2483,N_49529,N_49796);
xor UO_2484 (O_2484,N_49315,N_49457);
nor UO_2485 (O_2485,N_49272,N_49704);
and UO_2486 (O_2486,N_49082,N_49639);
or UO_2487 (O_2487,N_49492,N_49767);
nor UO_2488 (O_2488,N_49119,N_49049);
and UO_2489 (O_2489,N_49129,N_49743);
xor UO_2490 (O_2490,N_49162,N_49660);
and UO_2491 (O_2491,N_49477,N_49079);
nand UO_2492 (O_2492,N_49294,N_49563);
nand UO_2493 (O_2493,N_49881,N_49534);
or UO_2494 (O_2494,N_49955,N_49347);
or UO_2495 (O_2495,N_49497,N_49253);
or UO_2496 (O_2496,N_49053,N_49445);
nand UO_2497 (O_2497,N_49932,N_49797);
or UO_2498 (O_2498,N_49505,N_49605);
nor UO_2499 (O_2499,N_49811,N_49931);
xnor UO_2500 (O_2500,N_49176,N_49678);
and UO_2501 (O_2501,N_49555,N_49479);
nand UO_2502 (O_2502,N_49889,N_49285);
xnor UO_2503 (O_2503,N_49692,N_49528);
nor UO_2504 (O_2504,N_49246,N_49581);
xor UO_2505 (O_2505,N_49821,N_49017);
and UO_2506 (O_2506,N_49701,N_49792);
xnor UO_2507 (O_2507,N_49094,N_49202);
and UO_2508 (O_2508,N_49893,N_49332);
xor UO_2509 (O_2509,N_49179,N_49077);
xor UO_2510 (O_2510,N_49192,N_49171);
nor UO_2511 (O_2511,N_49079,N_49472);
nand UO_2512 (O_2512,N_49342,N_49217);
and UO_2513 (O_2513,N_49866,N_49706);
and UO_2514 (O_2514,N_49139,N_49850);
or UO_2515 (O_2515,N_49919,N_49650);
and UO_2516 (O_2516,N_49174,N_49086);
nand UO_2517 (O_2517,N_49509,N_49156);
xnor UO_2518 (O_2518,N_49481,N_49669);
xnor UO_2519 (O_2519,N_49436,N_49734);
xnor UO_2520 (O_2520,N_49738,N_49704);
xnor UO_2521 (O_2521,N_49593,N_49493);
nand UO_2522 (O_2522,N_49275,N_49916);
and UO_2523 (O_2523,N_49593,N_49717);
nor UO_2524 (O_2524,N_49971,N_49018);
nand UO_2525 (O_2525,N_49093,N_49843);
xnor UO_2526 (O_2526,N_49454,N_49849);
and UO_2527 (O_2527,N_49505,N_49423);
or UO_2528 (O_2528,N_49249,N_49442);
xnor UO_2529 (O_2529,N_49039,N_49912);
xnor UO_2530 (O_2530,N_49118,N_49971);
nand UO_2531 (O_2531,N_49467,N_49995);
nand UO_2532 (O_2532,N_49310,N_49819);
and UO_2533 (O_2533,N_49389,N_49426);
or UO_2534 (O_2534,N_49082,N_49318);
xor UO_2535 (O_2535,N_49841,N_49708);
xor UO_2536 (O_2536,N_49078,N_49856);
nand UO_2537 (O_2537,N_49871,N_49910);
and UO_2538 (O_2538,N_49850,N_49739);
xnor UO_2539 (O_2539,N_49706,N_49310);
or UO_2540 (O_2540,N_49811,N_49696);
nand UO_2541 (O_2541,N_49716,N_49968);
nor UO_2542 (O_2542,N_49416,N_49861);
or UO_2543 (O_2543,N_49613,N_49155);
xnor UO_2544 (O_2544,N_49646,N_49423);
nor UO_2545 (O_2545,N_49618,N_49095);
or UO_2546 (O_2546,N_49728,N_49706);
or UO_2547 (O_2547,N_49764,N_49334);
and UO_2548 (O_2548,N_49156,N_49654);
and UO_2549 (O_2549,N_49050,N_49077);
xnor UO_2550 (O_2550,N_49772,N_49034);
nand UO_2551 (O_2551,N_49062,N_49884);
xor UO_2552 (O_2552,N_49933,N_49747);
nor UO_2553 (O_2553,N_49636,N_49932);
or UO_2554 (O_2554,N_49819,N_49517);
nor UO_2555 (O_2555,N_49321,N_49381);
nand UO_2556 (O_2556,N_49759,N_49198);
nand UO_2557 (O_2557,N_49279,N_49443);
and UO_2558 (O_2558,N_49220,N_49068);
xnor UO_2559 (O_2559,N_49682,N_49119);
nand UO_2560 (O_2560,N_49362,N_49167);
xnor UO_2561 (O_2561,N_49057,N_49407);
and UO_2562 (O_2562,N_49624,N_49376);
or UO_2563 (O_2563,N_49264,N_49150);
and UO_2564 (O_2564,N_49184,N_49351);
or UO_2565 (O_2565,N_49759,N_49197);
or UO_2566 (O_2566,N_49357,N_49102);
and UO_2567 (O_2567,N_49150,N_49457);
nor UO_2568 (O_2568,N_49816,N_49374);
and UO_2569 (O_2569,N_49011,N_49785);
nand UO_2570 (O_2570,N_49354,N_49366);
nor UO_2571 (O_2571,N_49351,N_49731);
and UO_2572 (O_2572,N_49341,N_49747);
nor UO_2573 (O_2573,N_49619,N_49109);
or UO_2574 (O_2574,N_49150,N_49986);
nor UO_2575 (O_2575,N_49375,N_49178);
and UO_2576 (O_2576,N_49798,N_49361);
nand UO_2577 (O_2577,N_49524,N_49799);
nand UO_2578 (O_2578,N_49581,N_49748);
nor UO_2579 (O_2579,N_49697,N_49368);
or UO_2580 (O_2580,N_49060,N_49214);
or UO_2581 (O_2581,N_49200,N_49590);
xor UO_2582 (O_2582,N_49307,N_49477);
or UO_2583 (O_2583,N_49354,N_49323);
and UO_2584 (O_2584,N_49939,N_49602);
and UO_2585 (O_2585,N_49695,N_49614);
and UO_2586 (O_2586,N_49802,N_49935);
or UO_2587 (O_2587,N_49113,N_49862);
nor UO_2588 (O_2588,N_49292,N_49371);
xnor UO_2589 (O_2589,N_49326,N_49216);
or UO_2590 (O_2590,N_49962,N_49370);
nor UO_2591 (O_2591,N_49622,N_49083);
or UO_2592 (O_2592,N_49726,N_49757);
nor UO_2593 (O_2593,N_49857,N_49800);
and UO_2594 (O_2594,N_49508,N_49447);
nor UO_2595 (O_2595,N_49362,N_49422);
xnor UO_2596 (O_2596,N_49727,N_49828);
xor UO_2597 (O_2597,N_49554,N_49156);
xnor UO_2598 (O_2598,N_49125,N_49608);
xnor UO_2599 (O_2599,N_49211,N_49057);
or UO_2600 (O_2600,N_49426,N_49413);
nor UO_2601 (O_2601,N_49266,N_49662);
and UO_2602 (O_2602,N_49226,N_49130);
nor UO_2603 (O_2603,N_49994,N_49204);
nor UO_2604 (O_2604,N_49670,N_49653);
nor UO_2605 (O_2605,N_49445,N_49888);
and UO_2606 (O_2606,N_49222,N_49358);
or UO_2607 (O_2607,N_49755,N_49898);
or UO_2608 (O_2608,N_49455,N_49437);
xnor UO_2609 (O_2609,N_49559,N_49030);
nor UO_2610 (O_2610,N_49681,N_49636);
nor UO_2611 (O_2611,N_49399,N_49441);
or UO_2612 (O_2612,N_49039,N_49644);
or UO_2613 (O_2613,N_49178,N_49482);
nand UO_2614 (O_2614,N_49342,N_49014);
xor UO_2615 (O_2615,N_49000,N_49299);
or UO_2616 (O_2616,N_49681,N_49647);
nand UO_2617 (O_2617,N_49407,N_49050);
nand UO_2618 (O_2618,N_49619,N_49677);
or UO_2619 (O_2619,N_49088,N_49766);
nor UO_2620 (O_2620,N_49491,N_49305);
xor UO_2621 (O_2621,N_49353,N_49469);
and UO_2622 (O_2622,N_49952,N_49809);
nand UO_2623 (O_2623,N_49297,N_49764);
or UO_2624 (O_2624,N_49253,N_49624);
or UO_2625 (O_2625,N_49115,N_49146);
and UO_2626 (O_2626,N_49815,N_49399);
nor UO_2627 (O_2627,N_49143,N_49626);
nor UO_2628 (O_2628,N_49758,N_49862);
and UO_2629 (O_2629,N_49156,N_49613);
or UO_2630 (O_2630,N_49800,N_49761);
nand UO_2631 (O_2631,N_49636,N_49897);
nor UO_2632 (O_2632,N_49614,N_49409);
or UO_2633 (O_2633,N_49918,N_49221);
nand UO_2634 (O_2634,N_49913,N_49288);
xor UO_2635 (O_2635,N_49728,N_49508);
nor UO_2636 (O_2636,N_49997,N_49155);
nand UO_2637 (O_2637,N_49764,N_49966);
nor UO_2638 (O_2638,N_49593,N_49605);
or UO_2639 (O_2639,N_49803,N_49027);
nand UO_2640 (O_2640,N_49795,N_49277);
xor UO_2641 (O_2641,N_49607,N_49876);
nor UO_2642 (O_2642,N_49055,N_49468);
xnor UO_2643 (O_2643,N_49685,N_49350);
or UO_2644 (O_2644,N_49935,N_49638);
nor UO_2645 (O_2645,N_49407,N_49623);
nand UO_2646 (O_2646,N_49940,N_49362);
or UO_2647 (O_2647,N_49704,N_49083);
nand UO_2648 (O_2648,N_49318,N_49855);
nor UO_2649 (O_2649,N_49433,N_49302);
or UO_2650 (O_2650,N_49793,N_49570);
or UO_2651 (O_2651,N_49695,N_49531);
nand UO_2652 (O_2652,N_49664,N_49958);
or UO_2653 (O_2653,N_49035,N_49262);
nand UO_2654 (O_2654,N_49361,N_49780);
nor UO_2655 (O_2655,N_49502,N_49993);
and UO_2656 (O_2656,N_49770,N_49193);
or UO_2657 (O_2657,N_49215,N_49696);
nand UO_2658 (O_2658,N_49359,N_49080);
nand UO_2659 (O_2659,N_49250,N_49376);
xor UO_2660 (O_2660,N_49175,N_49373);
and UO_2661 (O_2661,N_49807,N_49469);
nor UO_2662 (O_2662,N_49966,N_49357);
nor UO_2663 (O_2663,N_49803,N_49840);
nand UO_2664 (O_2664,N_49367,N_49434);
nor UO_2665 (O_2665,N_49591,N_49291);
xor UO_2666 (O_2666,N_49659,N_49071);
or UO_2667 (O_2667,N_49679,N_49640);
nand UO_2668 (O_2668,N_49365,N_49337);
and UO_2669 (O_2669,N_49081,N_49534);
xnor UO_2670 (O_2670,N_49595,N_49234);
or UO_2671 (O_2671,N_49787,N_49815);
xnor UO_2672 (O_2672,N_49277,N_49468);
and UO_2673 (O_2673,N_49504,N_49108);
nor UO_2674 (O_2674,N_49966,N_49137);
and UO_2675 (O_2675,N_49551,N_49179);
and UO_2676 (O_2676,N_49628,N_49416);
xor UO_2677 (O_2677,N_49120,N_49304);
nor UO_2678 (O_2678,N_49750,N_49138);
and UO_2679 (O_2679,N_49690,N_49914);
and UO_2680 (O_2680,N_49019,N_49773);
and UO_2681 (O_2681,N_49821,N_49297);
nor UO_2682 (O_2682,N_49807,N_49689);
xor UO_2683 (O_2683,N_49434,N_49762);
xnor UO_2684 (O_2684,N_49853,N_49645);
nand UO_2685 (O_2685,N_49594,N_49509);
nor UO_2686 (O_2686,N_49691,N_49022);
nand UO_2687 (O_2687,N_49938,N_49203);
nor UO_2688 (O_2688,N_49879,N_49518);
nor UO_2689 (O_2689,N_49244,N_49155);
and UO_2690 (O_2690,N_49193,N_49620);
or UO_2691 (O_2691,N_49115,N_49812);
xor UO_2692 (O_2692,N_49847,N_49484);
xnor UO_2693 (O_2693,N_49591,N_49035);
nor UO_2694 (O_2694,N_49763,N_49854);
nor UO_2695 (O_2695,N_49933,N_49218);
or UO_2696 (O_2696,N_49721,N_49922);
xor UO_2697 (O_2697,N_49457,N_49796);
or UO_2698 (O_2698,N_49803,N_49405);
nand UO_2699 (O_2699,N_49735,N_49685);
xnor UO_2700 (O_2700,N_49754,N_49864);
nor UO_2701 (O_2701,N_49987,N_49119);
xnor UO_2702 (O_2702,N_49562,N_49853);
nand UO_2703 (O_2703,N_49947,N_49779);
xor UO_2704 (O_2704,N_49501,N_49262);
nand UO_2705 (O_2705,N_49869,N_49907);
nand UO_2706 (O_2706,N_49061,N_49538);
nand UO_2707 (O_2707,N_49272,N_49378);
and UO_2708 (O_2708,N_49235,N_49253);
nor UO_2709 (O_2709,N_49121,N_49341);
and UO_2710 (O_2710,N_49679,N_49888);
xnor UO_2711 (O_2711,N_49440,N_49763);
nand UO_2712 (O_2712,N_49443,N_49802);
nand UO_2713 (O_2713,N_49356,N_49006);
and UO_2714 (O_2714,N_49709,N_49956);
or UO_2715 (O_2715,N_49227,N_49326);
or UO_2716 (O_2716,N_49139,N_49762);
nand UO_2717 (O_2717,N_49293,N_49159);
nor UO_2718 (O_2718,N_49757,N_49066);
and UO_2719 (O_2719,N_49441,N_49514);
nor UO_2720 (O_2720,N_49316,N_49022);
and UO_2721 (O_2721,N_49891,N_49659);
and UO_2722 (O_2722,N_49135,N_49488);
xor UO_2723 (O_2723,N_49634,N_49139);
nand UO_2724 (O_2724,N_49878,N_49877);
or UO_2725 (O_2725,N_49472,N_49759);
or UO_2726 (O_2726,N_49879,N_49918);
or UO_2727 (O_2727,N_49854,N_49932);
xor UO_2728 (O_2728,N_49724,N_49242);
and UO_2729 (O_2729,N_49465,N_49124);
nor UO_2730 (O_2730,N_49084,N_49475);
or UO_2731 (O_2731,N_49312,N_49931);
xor UO_2732 (O_2732,N_49458,N_49527);
or UO_2733 (O_2733,N_49182,N_49342);
or UO_2734 (O_2734,N_49986,N_49944);
nand UO_2735 (O_2735,N_49718,N_49090);
nand UO_2736 (O_2736,N_49041,N_49401);
nor UO_2737 (O_2737,N_49134,N_49000);
xor UO_2738 (O_2738,N_49123,N_49835);
or UO_2739 (O_2739,N_49562,N_49805);
xnor UO_2740 (O_2740,N_49327,N_49137);
and UO_2741 (O_2741,N_49817,N_49896);
or UO_2742 (O_2742,N_49549,N_49286);
nand UO_2743 (O_2743,N_49386,N_49683);
or UO_2744 (O_2744,N_49499,N_49377);
nand UO_2745 (O_2745,N_49755,N_49328);
and UO_2746 (O_2746,N_49929,N_49121);
nor UO_2747 (O_2747,N_49033,N_49904);
nor UO_2748 (O_2748,N_49380,N_49984);
nor UO_2749 (O_2749,N_49405,N_49382);
and UO_2750 (O_2750,N_49668,N_49186);
nand UO_2751 (O_2751,N_49332,N_49981);
nand UO_2752 (O_2752,N_49649,N_49094);
nor UO_2753 (O_2753,N_49344,N_49987);
nand UO_2754 (O_2754,N_49123,N_49418);
or UO_2755 (O_2755,N_49418,N_49298);
nor UO_2756 (O_2756,N_49677,N_49837);
nor UO_2757 (O_2757,N_49288,N_49110);
nor UO_2758 (O_2758,N_49659,N_49652);
xor UO_2759 (O_2759,N_49630,N_49549);
and UO_2760 (O_2760,N_49173,N_49841);
nand UO_2761 (O_2761,N_49554,N_49126);
nand UO_2762 (O_2762,N_49204,N_49366);
and UO_2763 (O_2763,N_49164,N_49459);
nor UO_2764 (O_2764,N_49175,N_49023);
nor UO_2765 (O_2765,N_49323,N_49111);
xnor UO_2766 (O_2766,N_49004,N_49104);
xnor UO_2767 (O_2767,N_49409,N_49502);
nand UO_2768 (O_2768,N_49324,N_49205);
and UO_2769 (O_2769,N_49453,N_49973);
or UO_2770 (O_2770,N_49695,N_49093);
and UO_2771 (O_2771,N_49945,N_49619);
xnor UO_2772 (O_2772,N_49993,N_49862);
xnor UO_2773 (O_2773,N_49741,N_49960);
or UO_2774 (O_2774,N_49251,N_49752);
and UO_2775 (O_2775,N_49182,N_49460);
nor UO_2776 (O_2776,N_49638,N_49787);
nand UO_2777 (O_2777,N_49825,N_49136);
or UO_2778 (O_2778,N_49670,N_49226);
and UO_2779 (O_2779,N_49485,N_49792);
xor UO_2780 (O_2780,N_49421,N_49659);
and UO_2781 (O_2781,N_49954,N_49850);
nor UO_2782 (O_2782,N_49823,N_49591);
xnor UO_2783 (O_2783,N_49889,N_49306);
or UO_2784 (O_2784,N_49723,N_49505);
or UO_2785 (O_2785,N_49632,N_49949);
and UO_2786 (O_2786,N_49823,N_49810);
nand UO_2787 (O_2787,N_49331,N_49109);
nand UO_2788 (O_2788,N_49603,N_49095);
nand UO_2789 (O_2789,N_49673,N_49987);
or UO_2790 (O_2790,N_49546,N_49195);
or UO_2791 (O_2791,N_49157,N_49508);
xnor UO_2792 (O_2792,N_49958,N_49049);
or UO_2793 (O_2793,N_49709,N_49499);
xnor UO_2794 (O_2794,N_49669,N_49728);
xor UO_2795 (O_2795,N_49412,N_49043);
and UO_2796 (O_2796,N_49101,N_49765);
nor UO_2797 (O_2797,N_49594,N_49042);
nor UO_2798 (O_2798,N_49047,N_49463);
or UO_2799 (O_2799,N_49746,N_49245);
or UO_2800 (O_2800,N_49528,N_49818);
nand UO_2801 (O_2801,N_49570,N_49015);
nand UO_2802 (O_2802,N_49368,N_49048);
xnor UO_2803 (O_2803,N_49678,N_49128);
and UO_2804 (O_2804,N_49520,N_49615);
and UO_2805 (O_2805,N_49251,N_49930);
nor UO_2806 (O_2806,N_49374,N_49162);
xnor UO_2807 (O_2807,N_49990,N_49505);
nor UO_2808 (O_2808,N_49092,N_49207);
or UO_2809 (O_2809,N_49266,N_49408);
nand UO_2810 (O_2810,N_49587,N_49453);
nand UO_2811 (O_2811,N_49992,N_49479);
or UO_2812 (O_2812,N_49209,N_49504);
and UO_2813 (O_2813,N_49622,N_49286);
nor UO_2814 (O_2814,N_49577,N_49975);
nor UO_2815 (O_2815,N_49737,N_49640);
nor UO_2816 (O_2816,N_49027,N_49024);
nor UO_2817 (O_2817,N_49325,N_49805);
nand UO_2818 (O_2818,N_49747,N_49718);
xor UO_2819 (O_2819,N_49817,N_49023);
nor UO_2820 (O_2820,N_49241,N_49550);
and UO_2821 (O_2821,N_49565,N_49337);
nor UO_2822 (O_2822,N_49726,N_49034);
xor UO_2823 (O_2823,N_49846,N_49966);
or UO_2824 (O_2824,N_49607,N_49452);
nor UO_2825 (O_2825,N_49275,N_49199);
or UO_2826 (O_2826,N_49875,N_49053);
and UO_2827 (O_2827,N_49202,N_49986);
or UO_2828 (O_2828,N_49833,N_49128);
nor UO_2829 (O_2829,N_49005,N_49536);
xnor UO_2830 (O_2830,N_49645,N_49643);
nand UO_2831 (O_2831,N_49489,N_49078);
xor UO_2832 (O_2832,N_49672,N_49136);
nor UO_2833 (O_2833,N_49517,N_49631);
nor UO_2834 (O_2834,N_49172,N_49445);
or UO_2835 (O_2835,N_49219,N_49442);
nand UO_2836 (O_2836,N_49653,N_49956);
and UO_2837 (O_2837,N_49448,N_49890);
nor UO_2838 (O_2838,N_49725,N_49491);
or UO_2839 (O_2839,N_49684,N_49744);
nor UO_2840 (O_2840,N_49435,N_49517);
and UO_2841 (O_2841,N_49910,N_49943);
xnor UO_2842 (O_2842,N_49265,N_49029);
xor UO_2843 (O_2843,N_49890,N_49123);
xor UO_2844 (O_2844,N_49141,N_49477);
nand UO_2845 (O_2845,N_49473,N_49821);
or UO_2846 (O_2846,N_49495,N_49822);
nand UO_2847 (O_2847,N_49453,N_49999);
and UO_2848 (O_2848,N_49054,N_49368);
nor UO_2849 (O_2849,N_49425,N_49496);
nand UO_2850 (O_2850,N_49688,N_49305);
nor UO_2851 (O_2851,N_49733,N_49363);
xor UO_2852 (O_2852,N_49104,N_49111);
xnor UO_2853 (O_2853,N_49604,N_49982);
nand UO_2854 (O_2854,N_49914,N_49277);
nand UO_2855 (O_2855,N_49739,N_49979);
or UO_2856 (O_2856,N_49484,N_49190);
or UO_2857 (O_2857,N_49198,N_49489);
xnor UO_2858 (O_2858,N_49135,N_49518);
and UO_2859 (O_2859,N_49265,N_49882);
nor UO_2860 (O_2860,N_49800,N_49314);
nor UO_2861 (O_2861,N_49388,N_49267);
xor UO_2862 (O_2862,N_49289,N_49367);
nor UO_2863 (O_2863,N_49169,N_49391);
nand UO_2864 (O_2864,N_49280,N_49356);
nor UO_2865 (O_2865,N_49907,N_49384);
nor UO_2866 (O_2866,N_49504,N_49856);
nand UO_2867 (O_2867,N_49489,N_49171);
nand UO_2868 (O_2868,N_49587,N_49977);
or UO_2869 (O_2869,N_49706,N_49432);
nor UO_2870 (O_2870,N_49435,N_49906);
nor UO_2871 (O_2871,N_49843,N_49047);
or UO_2872 (O_2872,N_49641,N_49971);
or UO_2873 (O_2873,N_49062,N_49636);
or UO_2874 (O_2874,N_49789,N_49740);
and UO_2875 (O_2875,N_49553,N_49434);
nand UO_2876 (O_2876,N_49386,N_49631);
nand UO_2877 (O_2877,N_49262,N_49430);
nand UO_2878 (O_2878,N_49628,N_49695);
nor UO_2879 (O_2879,N_49642,N_49414);
nor UO_2880 (O_2880,N_49474,N_49778);
nand UO_2881 (O_2881,N_49188,N_49151);
xnor UO_2882 (O_2882,N_49156,N_49197);
or UO_2883 (O_2883,N_49413,N_49345);
xor UO_2884 (O_2884,N_49566,N_49708);
nand UO_2885 (O_2885,N_49913,N_49849);
nor UO_2886 (O_2886,N_49620,N_49659);
nand UO_2887 (O_2887,N_49845,N_49809);
nand UO_2888 (O_2888,N_49565,N_49693);
nand UO_2889 (O_2889,N_49230,N_49566);
and UO_2890 (O_2890,N_49311,N_49966);
and UO_2891 (O_2891,N_49376,N_49443);
and UO_2892 (O_2892,N_49951,N_49408);
nor UO_2893 (O_2893,N_49824,N_49517);
or UO_2894 (O_2894,N_49719,N_49474);
or UO_2895 (O_2895,N_49783,N_49082);
or UO_2896 (O_2896,N_49367,N_49659);
or UO_2897 (O_2897,N_49704,N_49403);
nand UO_2898 (O_2898,N_49315,N_49483);
nor UO_2899 (O_2899,N_49463,N_49261);
xnor UO_2900 (O_2900,N_49625,N_49608);
or UO_2901 (O_2901,N_49892,N_49709);
nor UO_2902 (O_2902,N_49019,N_49108);
or UO_2903 (O_2903,N_49801,N_49960);
xnor UO_2904 (O_2904,N_49491,N_49669);
nand UO_2905 (O_2905,N_49140,N_49443);
nand UO_2906 (O_2906,N_49496,N_49011);
nand UO_2907 (O_2907,N_49663,N_49069);
nor UO_2908 (O_2908,N_49471,N_49261);
nor UO_2909 (O_2909,N_49132,N_49233);
and UO_2910 (O_2910,N_49276,N_49416);
or UO_2911 (O_2911,N_49748,N_49642);
or UO_2912 (O_2912,N_49747,N_49876);
xor UO_2913 (O_2913,N_49811,N_49569);
and UO_2914 (O_2914,N_49136,N_49077);
xnor UO_2915 (O_2915,N_49630,N_49324);
xor UO_2916 (O_2916,N_49133,N_49131);
and UO_2917 (O_2917,N_49423,N_49100);
nand UO_2918 (O_2918,N_49983,N_49909);
nor UO_2919 (O_2919,N_49877,N_49379);
nor UO_2920 (O_2920,N_49257,N_49786);
xor UO_2921 (O_2921,N_49427,N_49589);
and UO_2922 (O_2922,N_49937,N_49196);
nor UO_2923 (O_2923,N_49777,N_49048);
and UO_2924 (O_2924,N_49109,N_49286);
xor UO_2925 (O_2925,N_49741,N_49407);
xnor UO_2926 (O_2926,N_49716,N_49249);
or UO_2927 (O_2927,N_49933,N_49897);
or UO_2928 (O_2928,N_49564,N_49845);
nor UO_2929 (O_2929,N_49306,N_49156);
xnor UO_2930 (O_2930,N_49132,N_49901);
and UO_2931 (O_2931,N_49149,N_49376);
or UO_2932 (O_2932,N_49413,N_49037);
nand UO_2933 (O_2933,N_49150,N_49765);
xnor UO_2934 (O_2934,N_49700,N_49164);
nand UO_2935 (O_2935,N_49042,N_49664);
nor UO_2936 (O_2936,N_49862,N_49110);
and UO_2937 (O_2937,N_49870,N_49998);
xor UO_2938 (O_2938,N_49272,N_49305);
nand UO_2939 (O_2939,N_49652,N_49288);
or UO_2940 (O_2940,N_49786,N_49161);
and UO_2941 (O_2941,N_49656,N_49236);
and UO_2942 (O_2942,N_49652,N_49443);
and UO_2943 (O_2943,N_49582,N_49682);
xnor UO_2944 (O_2944,N_49742,N_49777);
nor UO_2945 (O_2945,N_49903,N_49433);
nand UO_2946 (O_2946,N_49460,N_49713);
and UO_2947 (O_2947,N_49764,N_49144);
nor UO_2948 (O_2948,N_49182,N_49461);
and UO_2949 (O_2949,N_49632,N_49229);
xor UO_2950 (O_2950,N_49411,N_49186);
nand UO_2951 (O_2951,N_49631,N_49062);
xnor UO_2952 (O_2952,N_49820,N_49972);
and UO_2953 (O_2953,N_49515,N_49669);
or UO_2954 (O_2954,N_49489,N_49415);
and UO_2955 (O_2955,N_49678,N_49493);
and UO_2956 (O_2956,N_49216,N_49252);
xor UO_2957 (O_2957,N_49107,N_49944);
and UO_2958 (O_2958,N_49497,N_49952);
and UO_2959 (O_2959,N_49237,N_49848);
nor UO_2960 (O_2960,N_49025,N_49884);
nor UO_2961 (O_2961,N_49059,N_49925);
and UO_2962 (O_2962,N_49727,N_49686);
nand UO_2963 (O_2963,N_49248,N_49216);
nor UO_2964 (O_2964,N_49127,N_49886);
or UO_2965 (O_2965,N_49733,N_49182);
nor UO_2966 (O_2966,N_49487,N_49011);
nand UO_2967 (O_2967,N_49666,N_49488);
xor UO_2968 (O_2968,N_49701,N_49177);
nor UO_2969 (O_2969,N_49882,N_49327);
and UO_2970 (O_2970,N_49219,N_49678);
xor UO_2971 (O_2971,N_49699,N_49240);
xnor UO_2972 (O_2972,N_49454,N_49035);
xnor UO_2973 (O_2973,N_49770,N_49768);
xor UO_2974 (O_2974,N_49597,N_49657);
xnor UO_2975 (O_2975,N_49757,N_49665);
nand UO_2976 (O_2976,N_49237,N_49989);
nor UO_2977 (O_2977,N_49608,N_49496);
xor UO_2978 (O_2978,N_49344,N_49225);
xnor UO_2979 (O_2979,N_49452,N_49210);
nand UO_2980 (O_2980,N_49151,N_49687);
nand UO_2981 (O_2981,N_49354,N_49876);
nand UO_2982 (O_2982,N_49038,N_49171);
nor UO_2983 (O_2983,N_49419,N_49694);
or UO_2984 (O_2984,N_49545,N_49950);
nand UO_2985 (O_2985,N_49976,N_49276);
nor UO_2986 (O_2986,N_49856,N_49986);
nand UO_2987 (O_2987,N_49759,N_49967);
xor UO_2988 (O_2988,N_49340,N_49798);
xnor UO_2989 (O_2989,N_49282,N_49415);
or UO_2990 (O_2990,N_49777,N_49994);
nor UO_2991 (O_2991,N_49996,N_49463);
nor UO_2992 (O_2992,N_49221,N_49330);
and UO_2993 (O_2993,N_49250,N_49490);
nor UO_2994 (O_2994,N_49184,N_49333);
and UO_2995 (O_2995,N_49694,N_49190);
nand UO_2996 (O_2996,N_49369,N_49413);
or UO_2997 (O_2997,N_49583,N_49565);
and UO_2998 (O_2998,N_49325,N_49565);
and UO_2999 (O_2999,N_49942,N_49288);
or UO_3000 (O_3000,N_49611,N_49287);
nand UO_3001 (O_3001,N_49179,N_49481);
and UO_3002 (O_3002,N_49289,N_49973);
and UO_3003 (O_3003,N_49646,N_49635);
and UO_3004 (O_3004,N_49457,N_49200);
nor UO_3005 (O_3005,N_49465,N_49261);
nand UO_3006 (O_3006,N_49521,N_49957);
nor UO_3007 (O_3007,N_49313,N_49878);
nor UO_3008 (O_3008,N_49086,N_49886);
and UO_3009 (O_3009,N_49309,N_49491);
and UO_3010 (O_3010,N_49706,N_49096);
xnor UO_3011 (O_3011,N_49177,N_49221);
nor UO_3012 (O_3012,N_49933,N_49682);
or UO_3013 (O_3013,N_49499,N_49717);
nand UO_3014 (O_3014,N_49796,N_49875);
or UO_3015 (O_3015,N_49999,N_49395);
xnor UO_3016 (O_3016,N_49750,N_49356);
nand UO_3017 (O_3017,N_49349,N_49448);
or UO_3018 (O_3018,N_49777,N_49979);
and UO_3019 (O_3019,N_49741,N_49989);
nand UO_3020 (O_3020,N_49088,N_49611);
or UO_3021 (O_3021,N_49495,N_49712);
nand UO_3022 (O_3022,N_49106,N_49926);
or UO_3023 (O_3023,N_49153,N_49260);
and UO_3024 (O_3024,N_49694,N_49255);
or UO_3025 (O_3025,N_49456,N_49873);
and UO_3026 (O_3026,N_49911,N_49515);
nand UO_3027 (O_3027,N_49104,N_49909);
xor UO_3028 (O_3028,N_49142,N_49982);
nor UO_3029 (O_3029,N_49706,N_49809);
nand UO_3030 (O_3030,N_49522,N_49166);
or UO_3031 (O_3031,N_49691,N_49938);
or UO_3032 (O_3032,N_49913,N_49050);
or UO_3033 (O_3033,N_49403,N_49454);
and UO_3034 (O_3034,N_49381,N_49096);
nand UO_3035 (O_3035,N_49156,N_49047);
nand UO_3036 (O_3036,N_49770,N_49491);
and UO_3037 (O_3037,N_49504,N_49723);
xor UO_3038 (O_3038,N_49266,N_49677);
nand UO_3039 (O_3039,N_49298,N_49872);
or UO_3040 (O_3040,N_49785,N_49981);
nand UO_3041 (O_3041,N_49805,N_49220);
and UO_3042 (O_3042,N_49663,N_49326);
xor UO_3043 (O_3043,N_49100,N_49765);
nand UO_3044 (O_3044,N_49638,N_49455);
and UO_3045 (O_3045,N_49099,N_49316);
nor UO_3046 (O_3046,N_49600,N_49770);
nand UO_3047 (O_3047,N_49560,N_49719);
xor UO_3048 (O_3048,N_49053,N_49742);
nor UO_3049 (O_3049,N_49667,N_49922);
nor UO_3050 (O_3050,N_49861,N_49010);
xnor UO_3051 (O_3051,N_49856,N_49418);
nor UO_3052 (O_3052,N_49083,N_49679);
nand UO_3053 (O_3053,N_49052,N_49203);
nand UO_3054 (O_3054,N_49280,N_49514);
or UO_3055 (O_3055,N_49873,N_49091);
nand UO_3056 (O_3056,N_49469,N_49871);
and UO_3057 (O_3057,N_49686,N_49159);
nand UO_3058 (O_3058,N_49878,N_49299);
nor UO_3059 (O_3059,N_49818,N_49982);
nand UO_3060 (O_3060,N_49288,N_49079);
nor UO_3061 (O_3061,N_49725,N_49132);
and UO_3062 (O_3062,N_49657,N_49218);
xnor UO_3063 (O_3063,N_49801,N_49970);
or UO_3064 (O_3064,N_49981,N_49167);
xnor UO_3065 (O_3065,N_49899,N_49430);
or UO_3066 (O_3066,N_49996,N_49977);
nor UO_3067 (O_3067,N_49718,N_49047);
nor UO_3068 (O_3068,N_49362,N_49393);
xnor UO_3069 (O_3069,N_49777,N_49525);
xor UO_3070 (O_3070,N_49809,N_49343);
or UO_3071 (O_3071,N_49295,N_49467);
nor UO_3072 (O_3072,N_49825,N_49524);
nor UO_3073 (O_3073,N_49598,N_49395);
and UO_3074 (O_3074,N_49180,N_49015);
nor UO_3075 (O_3075,N_49818,N_49610);
or UO_3076 (O_3076,N_49628,N_49732);
or UO_3077 (O_3077,N_49282,N_49028);
nor UO_3078 (O_3078,N_49116,N_49139);
and UO_3079 (O_3079,N_49432,N_49561);
nor UO_3080 (O_3080,N_49447,N_49793);
xor UO_3081 (O_3081,N_49920,N_49526);
nor UO_3082 (O_3082,N_49371,N_49815);
nand UO_3083 (O_3083,N_49855,N_49396);
xor UO_3084 (O_3084,N_49648,N_49458);
xor UO_3085 (O_3085,N_49073,N_49062);
xnor UO_3086 (O_3086,N_49576,N_49398);
or UO_3087 (O_3087,N_49153,N_49472);
and UO_3088 (O_3088,N_49111,N_49002);
xor UO_3089 (O_3089,N_49606,N_49237);
or UO_3090 (O_3090,N_49454,N_49068);
nand UO_3091 (O_3091,N_49285,N_49585);
xnor UO_3092 (O_3092,N_49851,N_49817);
and UO_3093 (O_3093,N_49601,N_49469);
nand UO_3094 (O_3094,N_49182,N_49582);
nor UO_3095 (O_3095,N_49600,N_49450);
or UO_3096 (O_3096,N_49621,N_49851);
and UO_3097 (O_3097,N_49881,N_49309);
nand UO_3098 (O_3098,N_49884,N_49805);
or UO_3099 (O_3099,N_49846,N_49742);
nand UO_3100 (O_3100,N_49707,N_49787);
xnor UO_3101 (O_3101,N_49661,N_49641);
nor UO_3102 (O_3102,N_49959,N_49389);
or UO_3103 (O_3103,N_49976,N_49014);
xnor UO_3104 (O_3104,N_49486,N_49822);
xnor UO_3105 (O_3105,N_49998,N_49338);
or UO_3106 (O_3106,N_49863,N_49892);
or UO_3107 (O_3107,N_49938,N_49965);
and UO_3108 (O_3108,N_49086,N_49263);
or UO_3109 (O_3109,N_49190,N_49053);
nand UO_3110 (O_3110,N_49461,N_49644);
and UO_3111 (O_3111,N_49624,N_49683);
nor UO_3112 (O_3112,N_49007,N_49716);
nand UO_3113 (O_3113,N_49251,N_49185);
nor UO_3114 (O_3114,N_49495,N_49785);
or UO_3115 (O_3115,N_49801,N_49665);
and UO_3116 (O_3116,N_49629,N_49961);
and UO_3117 (O_3117,N_49206,N_49967);
or UO_3118 (O_3118,N_49217,N_49595);
or UO_3119 (O_3119,N_49553,N_49379);
or UO_3120 (O_3120,N_49737,N_49797);
nand UO_3121 (O_3121,N_49822,N_49869);
nand UO_3122 (O_3122,N_49728,N_49572);
xor UO_3123 (O_3123,N_49257,N_49132);
nor UO_3124 (O_3124,N_49460,N_49706);
xnor UO_3125 (O_3125,N_49702,N_49549);
nor UO_3126 (O_3126,N_49968,N_49894);
xnor UO_3127 (O_3127,N_49896,N_49630);
and UO_3128 (O_3128,N_49013,N_49517);
and UO_3129 (O_3129,N_49991,N_49184);
or UO_3130 (O_3130,N_49404,N_49523);
xnor UO_3131 (O_3131,N_49316,N_49717);
or UO_3132 (O_3132,N_49384,N_49678);
or UO_3133 (O_3133,N_49168,N_49977);
nor UO_3134 (O_3134,N_49543,N_49481);
xnor UO_3135 (O_3135,N_49126,N_49797);
or UO_3136 (O_3136,N_49044,N_49685);
xor UO_3137 (O_3137,N_49272,N_49349);
xor UO_3138 (O_3138,N_49973,N_49057);
or UO_3139 (O_3139,N_49381,N_49000);
or UO_3140 (O_3140,N_49726,N_49229);
xor UO_3141 (O_3141,N_49645,N_49207);
nand UO_3142 (O_3142,N_49816,N_49801);
nor UO_3143 (O_3143,N_49762,N_49562);
nand UO_3144 (O_3144,N_49358,N_49259);
xor UO_3145 (O_3145,N_49386,N_49690);
and UO_3146 (O_3146,N_49336,N_49802);
nand UO_3147 (O_3147,N_49656,N_49801);
or UO_3148 (O_3148,N_49881,N_49968);
xnor UO_3149 (O_3149,N_49873,N_49544);
nand UO_3150 (O_3150,N_49081,N_49270);
xnor UO_3151 (O_3151,N_49091,N_49829);
or UO_3152 (O_3152,N_49764,N_49244);
nand UO_3153 (O_3153,N_49701,N_49161);
nor UO_3154 (O_3154,N_49328,N_49778);
nand UO_3155 (O_3155,N_49394,N_49300);
xnor UO_3156 (O_3156,N_49326,N_49366);
xnor UO_3157 (O_3157,N_49507,N_49011);
nor UO_3158 (O_3158,N_49854,N_49611);
and UO_3159 (O_3159,N_49515,N_49073);
nand UO_3160 (O_3160,N_49572,N_49899);
xor UO_3161 (O_3161,N_49016,N_49192);
or UO_3162 (O_3162,N_49791,N_49004);
or UO_3163 (O_3163,N_49554,N_49712);
nor UO_3164 (O_3164,N_49073,N_49986);
xor UO_3165 (O_3165,N_49639,N_49173);
nand UO_3166 (O_3166,N_49525,N_49034);
nand UO_3167 (O_3167,N_49055,N_49123);
nand UO_3168 (O_3168,N_49646,N_49751);
xor UO_3169 (O_3169,N_49022,N_49304);
xnor UO_3170 (O_3170,N_49906,N_49526);
xnor UO_3171 (O_3171,N_49693,N_49069);
xor UO_3172 (O_3172,N_49582,N_49537);
nor UO_3173 (O_3173,N_49493,N_49652);
xor UO_3174 (O_3174,N_49109,N_49950);
and UO_3175 (O_3175,N_49105,N_49542);
nand UO_3176 (O_3176,N_49677,N_49988);
and UO_3177 (O_3177,N_49579,N_49681);
and UO_3178 (O_3178,N_49386,N_49739);
nand UO_3179 (O_3179,N_49975,N_49725);
or UO_3180 (O_3180,N_49071,N_49468);
nand UO_3181 (O_3181,N_49062,N_49763);
nand UO_3182 (O_3182,N_49670,N_49935);
nand UO_3183 (O_3183,N_49359,N_49431);
nand UO_3184 (O_3184,N_49509,N_49943);
nand UO_3185 (O_3185,N_49284,N_49273);
nor UO_3186 (O_3186,N_49122,N_49667);
or UO_3187 (O_3187,N_49784,N_49339);
nor UO_3188 (O_3188,N_49288,N_49297);
nor UO_3189 (O_3189,N_49028,N_49664);
nand UO_3190 (O_3190,N_49122,N_49262);
nand UO_3191 (O_3191,N_49048,N_49426);
and UO_3192 (O_3192,N_49941,N_49656);
xor UO_3193 (O_3193,N_49465,N_49975);
xnor UO_3194 (O_3194,N_49951,N_49338);
nor UO_3195 (O_3195,N_49869,N_49927);
nand UO_3196 (O_3196,N_49571,N_49840);
nand UO_3197 (O_3197,N_49063,N_49761);
or UO_3198 (O_3198,N_49775,N_49326);
nand UO_3199 (O_3199,N_49517,N_49483);
xnor UO_3200 (O_3200,N_49047,N_49726);
nor UO_3201 (O_3201,N_49414,N_49458);
nor UO_3202 (O_3202,N_49524,N_49892);
xor UO_3203 (O_3203,N_49956,N_49488);
xnor UO_3204 (O_3204,N_49464,N_49512);
and UO_3205 (O_3205,N_49621,N_49534);
nand UO_3206 (O_3206,N_49532,N_49366);
nand UO_3207 (O_3207,N_49980,N_49623);
nand UO_3208 (O_3208,N_49029,N_49907);
nand UO_3209 (O_3209,N_49959,N_49564);
nand UO_3210 (O_3210,N_49486,N_49633);
and UO_3211 (O_3211,N_49013,N_49481);
and UO_3212 (O_3212,N_49181,N_49563);
or UO_3213 (O_3213,N_49797,N_49108);
nand UO_3214 (O_3214,N_49158,N_49173);
nor UO_3215 (O_3215,N_49703,N_49231);
xor UO_3216 (O_3216,N_49371,N_49615);
xor UO_3217 (O_3217,N_49311,N_49733);
or UO_3218 (O_3218,N_49728,N_49504);
nor UO_3219 (O_3219,N_49504,N_49911);
and UO_3220 (O_3220,N_49346,N_49629);
nand UO_3221 (O_3221,N_49433,N_49562);
nand UO_3222 (O_3222,N_49785,N_49181);
or UO_3223 (O_3223,N_49628,N_49417);
nor UO_3224 (O_3224,N_49195,N_49281);
or UO_3225 (O_3225,N_49414,N_49307);
xor UO_3226 (O_3226,N_49111,N_49558);
xor UO_3227 (O_3227,N_49565,N_49331);
and UO_3228 (O_3228,N_49238,N_49407);
xnor UO_3229 (O_3229,N_49109,N_49283);
nand UO_3230 (O_3230,N_49274,N_49149);
nand UO_3231 (O_3231,N_49976,N_49803);
nand UO_3232 (O_3232,N_49547,N_49632);
nand UO_3233 (O_3233,N_49062,N_49003);
and UO_3234 (O_3234,N_49843,N_49989);
and UO_3235 (O_3235,N_49322,N_49078);
nand UO_3236 (O_3236,N_49048,N_49344);
xor UO_3237 (O_3237,N_49627,N_49341);
xnor UO_3238 (O_3238,N_49339,N_49106);
and UO_3239 (O_3239,N_49847,N_49583);
xor UO_3240 (O_3240,N_49532,N_49867);
nor UO_3241 (O_3241,N_49168,N_49090);
and UO_3242 (O_3242,N_49190,N_49378);
nand UO_3243 (O_3243,N_49890,N_49687);
xor UO_3244 (O_3244,N_49863,N_49633);
nor UO_3245 (O_3245,N_49196,N_49880);
or UO_3246 (O_3246,N_49100,N_49452);
and UO_3247 (O_3247,N_49548,N_49585);
or UO_3248 (O_3248,N_49165,N_49787);
or UO_3249 (O_3249,N_49392,N_49691);
xor UO_3250 (O_3250,N_49244,N_49267);
xor UO_3251 (O_3251,N_49364,N_49562);
and UO_3252 (O_3252,N_49225,N_49994);
nand UO_3253 (O_3253,N_49474,N_49904);
and UO_3254 (O_3254,N_49025,N_49299);
or UO_3255 (O_3255,N_49992,N_49458);
and UO_3256 (O_3256,N_49362,N_49381);
and UO_3257 (O_3257,N_49930,N_49733);
or UO_3258 (O_3258,N_49619,N_49507);
nand UO_3259 (O_3259,N_49731,N_49383);
or UO_3260 (O_3260,N_49471,N_49106);
and UO_3261 (O_3261,N_49380,N_49982);
xnor UO_3262 (O_3262,N_49871,N_49848);
and UO_3263 (O_3263,N_49374,N_49466);
xor UO_3264 (O_3264,N_49051,N_49934);
nand UO_3265 (O_3265,N_49790,N_49648);
nor UO_3266 (O_3266,N_49611,N_49590);
and UO_3267 (O_3267,N_49800,N_49677);
or UO_3268 (O_3268,N_49965,N_49264);
xnor UO_3269 (O_3269,N_49920,N_49948);
or UO_3270 (O_3270,N_49318,N_49342);
or UO_3271 (O_3271,N_49925,N_49800);
xor UO_3272 (O_3272,N_49919,N_49951);
xnor UO_3273 (O_3273,N_49050,N_49768);
xnor UO_3274 (O_3274,N_49387,N_49629);
nor UO_3275 (O_3275,N_49825,N_49760);
nand UO_3276 (O_3276,N_49000,N_49508);
xor UO_3277 (O_3277,N_49473,N_49139);
xor UO_3278 (O_3278,N_49473,N_49221);
nand UO_3279 (O_3279,N_49502,N_49127);
nor UO_3280 (O_3280,N_49294,N_49884);
or UO_3281 (O_3281,N_49399,N_49263);
nor UO_3282 (O_3282,N_49619,N_49703);
nand UO_3283 (O_3283,N_49634,N_49803);
nor UO_3284 (O_3284,N_49736,N_49900);
and UO_3285 (O_3285,N_49585,N_49354);
xnor UO_3286 (O_3286,N_49169,N_49283);
or UO_3287 (O_3287,N_49298,N_49765);
and UO_3288 (O_3288,N_49496,N_49351);
nor UO_3289 (O_3289,N_49428,N_49062);
xor UO_3290 (O_3290,N_49807,N_49822);
nand UO_3291 (O_3291,N_49897,N_49499);
and UO_3292 (O_3292,N_49926,N_49835);
nand UO_3293 (O_3293,N_49618,N_49003);
and UO_3294 (O_3294,N_49201,N_49995);
nor UO_3295 (O_3295,N_49544,N_49622);
and UO_3296 (O_3296,N_49568,N_49192);
nand UO_3297 (O_3297,N_49974,N_49297);
and UO_3298 (O_3298,N_49922,N_49364);
nor UO_3299 (O_3299,N_49779,N_49740);
nand UO_3300 (O_3300,N_49183,N_49642);
and UO_3301 (O_3301,N_49892,N_49807);
nor UO_3302 (O_3302,N_49372,N_49184);
nor UO_3303 (O_3303,N_49855,N_49289);
xnor UO_3304 (O_3304,N_49629,N_49293);
and UO_3305 (O_3305,N_49102,N_49534);
nor UO_3306 (O_3306,N_49799,N_49286);
nor UO_3307 (O_3307,N_49351,N_49343);
xor UO_3308 (O_3308,N_49330,N_49249);
or UO_3309 (O_3309,N_49274,N_49383);
and UO_3310 (O_3310,N_49575,N_49439);
nor UO_3311 (O_3311,N_49260,N_49287);
and UO_3312 (O_3312,N_49738,N_49961);
xor UO_3313 (O_3313,N_49780,N_49539);
and UO_3314 (O_3314,N_49146,N_49603);
nand UO_3315 (O_3315,N_49103,N_49391);
xnor UO_3316 (O_3316,N_49033,N_49777);
or UO_3317 (O_3317,N_49962,N_49079);
nor UO_3318 (O_3318,N_49876,N_49656);
xor UO_3319 (O_3319,N_49950,N_49006);
and UO_3320 (O_3320,N_49541,N_49390);
nand UO_3321 (O_3321,N_49157,N_49126);
nor UO_3322 (O_3322,N_49494,N_49055);
nor UO_3323 (O_3323,N_49601,N_49568);
xor UO_3324 (O_3324,N_49753,N_49906);
nand UO_3325 (O_3325,N_49540,N_49726);
xor UO_3326 (O_3326,N_49320,N_49633);
nor UO_3327 (O_3327,N_49329,N_49211);
and UO_3328 (O_3328,N_49134,N_49555);
or UO_3329 (O_3329,N_49761,N_49953);
or UO_3330 (O_3330,N_49906,N_49230);
xor UO_3331 (O_3331,N_49018,N_49219);
and UO_3332 (O_3332,N_49349,N_49124);
nand UO_3333 (O_3333,N_49919,N_49154);
and UO_3334 (O_3334,N_49410,N_49390);
xnor UO_3335 (O_3335,N_49683,N_49295);
or UO_3336 (O_3336,N_49950,N_49214);
and UO_3337 (O_3337,N_49805,N_49547);
nand UO_3338 (O_3338,N_49643,N_49698);
and UO_3339 (O_3339,N_49198,N_49445);
and UO_3340 (O_3340,N_49892,N_49344);
and UO_3341 (O_3341,N_49045,N_49113);
nand UO_3342 (O_3342,N_49847,N_49004);
nand UO_3343 (O_3343,N_49333,N_49524);
xnor UO_3344 (O_3344,N_49193,N_49177);
nand UO_3345 (O_3345,N_49187,N_49879);
nand UO_3346 (O_3346,N_49209,N_49024);
and UO_3347 (O_3347,N_49715,N_49838);
and UO_3348 (O_3348,N_49396,N_49475);
xor UO_3349 (O_3349,N_49705,N_49777);
nand UO_3350 (O_3350,N_49811,N_49223);
or UO_3351 (O_3351,N_49788,N_49621);
and UO_3352 (O_3352,N_49483,N_49843);
or UO_3353 (O_3353,N_49408,N_49454);
nor UO_3354 (O_3354,N_49172,N_49738);
xnor UO_3355 (O_3355,N_49421,N_49782);
nand UO_3356 (O_3356,N_49804,N_49206);
and UO_3357 (O_3357,N_49759,N_49884);
and UO_3358 (O_3358,N_49315,N_49931);
xnor UO_3359 (O_3359,N_49980,N_49332);
nand UO_3360 (O_3360,N_49340,N_49406);
nand UO_3361 (O_3361,N_49280,N_49993);
nor UO_3362 (O_3362,N_49185,N_49022);
nor UO_3363 (O_3363,N_49123,N_49048);
nand UO_3364 (O_3364,N_49897,N_49865);
and UO_3365 (O_3365,N_49761,N_49446);
nor UO_3366 (O_3366,N_49048,N_49100);
xnor UO_3367 (O_3367,N_49714,N_49679);
xor UO_3368 (O_3368,N_49091,N_49701);
nor UO_3369 (O_3369,N_49719,N_49387);
or UO_3370 (O_3370,N_49746,N_49352);
xnor UO_3371 (O_3371,N_49988,N_49023);
xnor UO_3372 (O_3372,N_49779,N_49952);
and UO_3373 (O_3373,N_49670,N_49560);
nand UO_3374 (O_3374,N_49437,N_49857);
xor UO_3375 (O_3375,N_49802,N_49649);
nand UO_3376 (O_3376,N_49395,N_49758);
or UO_3377 (O_3377,N_49561,N_49553);
nor UO_3378 (O_3378,N_49885,N_49622);
nor UO_3379 (O_3379,N_49685,N_49543);
xnor UO_3380 (O_3380,N_49249,N_49431);
nand UO_3381 (O_3381,N_49425,N_49332);
nand UO_3382 (O_3382,N_49297,N_49696);
nand UO_3383 (O_3383,N_49789,N_49819);
and UO_3384 (O_3384,N_49212,N_49356);
and UO_3385 (O_3385,N_49346,N_49560);
and UO_3386 (O_3386,N_49728,N_49901);
nand UO_3387 (O_3387,N_49462,N_49280);
nor UO_3388 (O_3388,N_49083,N_49865);
or UO_3389 (O_3389,N_49627,N_49358);
xnor UO_3390 (O_3390,N_49577,N_49765);
or UO_3391 (O_3391,N_49180,N_49635);
xnor UO_3392 (O_3392,N_49630,N_49434);
and UO_3393 (O_3393,N_49273,N_49383);
nand UO_3394 (O_3394,N_49955,N_49144);
nand UO_3395 (O_3395,N_49954,N_49645);
nor UO_3396 (O_3396,N_49690,N_49888);
xnor UO_3397 (O_3397,N_49971,N_49035);
xor UO_3398 (O_3398,N_49708,N_49667);
nand UO_3399 (O_3399,N_49688,N_49489);
or UO_3400 (O_3400,N_49920,N_49277);
and UO_3401 (O_3401,N_49544,N_49719);
or UO_3402 (O_3402,N_49088,N_49731);
and UO_3403 (O_3403,N_49419,N_49270);
nand UO_3404 (O_3404,N_49918,N_49087);
and UO_3405 (O_3405,N_49918,N_49151);
or UO_3406 (O_3406,N_49939,N_49365);
and UO_3407 (O_3407,N_49540,N_49687);
nand UO_3408 (O_3408,N_49858,N_49861);
or UO_3409 (O_3409,N_49358,N_49546);
nand UO_3410 (O_3410,N_49900,N_49642);
nor UO_3411 (O_3411,N_49275,N_49246);
and UO_3412 (O_3412,N_49717,N_49893);
and UO_3413 (O_3413,N_49937,N_49614);
nand UO_3414 (O_3414,N_49942,N_49656);
xor UO_3415 (O_3415,N_49256,N_49520);
xnor UO_3416 (O_3416,N_49861,N_49715);
and UO_3417 (O_3417,N_49978,N_49742);
nand UO_3418 (O_3418,N_49387,N_49620);
nor UO_3419 (O_3419,N_49150,N_49910);
or UO_3420 (O_3420,N_49969,N_49817);
or UO_3421 (O_3421,N_49116,N_49206);
and UO_3422 (O_3422,N_49595,N_49219);
or UO_3423 (O_3423,N_49959,N_49068);
xnor UO_3424 (O_3424,N_49845,N_49357);
nor UO_3425 (O_3425,N_49572,N_49433);
and UO_3426 (O_3426,N_49709,N_49525);
or UO_3427 (O_3427,N_49249,N_49207);
xnor UO_3428 (O_3428,N_49688,N_49812);
or UO_3429 (O_3429,N_49251,N_49366);
or UO_3430 (O_3430,N_49329,N_49207);
nor UO_3431 (O_3431,N_49799,N_49026);
xor UO_3432 (O_3432,N_49216,N_49732);
nand UO_3433 (O_3433,N_49757,N_49648);
nand UO_3434 (O_3434,N_49825,N_49217);
and UO_3435 (O_3435,N_49608,N_49150);
nand UO_3436 (O_3436,N_49837,N_49037);
xor UO_3437 (O_3437,N_49604,N_49644);
nor UO_3438 (O_3438,N_49923,N_49245);
nand UO_3439 (O_3439,N_49592,N_49800);
nand UO_3440 (O_3440,N_49198,N_49659);
and UO_3441 (O_3441,N_49168,N_49525);
and UO_3442 (O_3442,N_49645,N_49512);
nand UO_3443 (O_3443,N_49935,N_49840);
xnor UO_3444 (O_3444,N_49565,N_49078);
or UO_3445 (O_3445,N_49248,N_49261);
and UO_3446 (O_3446,N_49812,N_49532);
and UO_3447 (O_3447,N_49907,N_49895);
nand UO_3448 (O_3448,N_49946,N_49415);
nand UO_3449 (O_3449,N_49695,N_49696);
nand UO_3450 (O_3450,N_49153,N_49736);
nand UO_3451 (O_3451,N_49752,N_49658);
nor UO_3452 (O_3452,N_49150,N_49396);
xnor UO_3453 (O_3453,N_49779,N_49625);
nand UO_3454 (O_3454,N_49431,N_49981);
and UO_3455 (O_3455,N_49457,N_49551);
or UO_3456 (O_3456,N_49374,N_49131);
xor UO_3457 (O_3457,N_49331,N_49365);
xnor UO_3458 (O_3458,N_49837,N_49688);
xor UO_3459 (O_3459,N_49266,N_49228);
nand UO_3460 (O_3460,N_49410,N_49954);
nand UO_3461 (O_3461,N_49152,N_49132);
nand UO_3462 (O_3462,N_49542,N_49852);
nand UO_3463 (O_3463,N_49266,N_49298);
xor UO_3464 (O_3464,N_49271,N_49595);
or UO_3465 (O_3465,N_49859,N_49731);
nor UO_3466 (O_3466,N_49957,N_49187);
or UO_3467 (O_3467,N_49709,N_49682);
xor UO_3468 (O_3468,N_49406,N_49024);
and UO_3469 (O_3469,N_49723,N_49031);
nor UO_3470 (O_3470,N_49275,N_49812);
and UO_3471 (O_3471,N_49323,N_49587);
nor UO_3472 (O_3472,N_49560,N_49231);
xnor UO_3473 (O_3473,N_49567,N_49474);
or UO_3474 (O_3474,N_49825,N_49456);
xnor UO_3475 (O_3475,N_49137,N_49977);
and UO_3476 (O_3476,N_49756,N_49889);
and UO_3477 (O_3477,N_49535,N_49821);
nor UO_3478 (O_3478,N_49507,N_49192);
nand UO_3479 (O_3479,N_49922,N_49515);
nor UO_3480 (O_3480,N_49108,N_49987);
nand UO_3481 (O_3481,N_49039,N_49037);
or UO_3482 (O_3482,N_49294,N_49610);
nor UO_3483 (O_3483,N_49490,N_49500);
xor UO_3484 (O_3484,N_49966,N_49801);
and UO_3485 (O_3485,N_49782,N_49396);
nand UO_3486 (O_3486,N_49118,N_49713);
nor UO_3487 (O_3487,N_49082,N_49792);
nor UO_3488 (O_3488,N_49048,N_49695);
and UO_3489 (O_3489,N_49095,N_49274);
nand UO_3490 (O_3490,N_49519,N_49369);
and UO_3491 (O_3491,N_49645,N_49299);
nand UO_3492 (O_3492,N_49215,N_49286);
or UO_3493 (O_3493,N_49124,N_49446);
and UO_3494 (O_3494,N_49498,N_49004);
or UO_3495 (O_3495,N_49976,N_49058);
nand UO_3496 (O_3496,N_49697,N_49560);
or UO_3497 (O_3497,N_49832,N_49366);
and UO_3498 (O_3498,N_49883,N_49836);
nand UO_3499 (O_3499,N_49525,N_49538);
or UO_3500 (O_3500,N_49105,N_49327);
nand UO_3501 (O_3501,N_49992,N_49258);
and UO_3502 (O_3502,N_49131,N_49246);
or UO_3503 (O_3503,N_49881,N_49402);
and UO_3504 (O_3504,N_49469,N_49240);
xor UO_3505 (O_3505,N_49286,N_49290);
and UO_3506 (O_3506,N_49747,N_49874);
nor UO_3507 (O_3507,N_49552,N_49356);
xnor UO_3508 (O_3508,N_49870,N_49322);
or UO_3509 (O_3509,N_49418,N_49642);
or UO_3510 (O_3510,N_49791,N_49092);
and UO_3511 (O_3511,N_49581,N_49946);
xnor UO_3512 (O_3512,N_49548,N_49386);
xor UO_3513 (O_3513,N_49705,N_49111);
nor UO_3514 (O_3514,N_49694,N_49177);
xor UO_3515 (O_3515,N_49615,N_49446);
xor UO_3516 (O_3516,N_49991,N_49977);
nor UO_3517 (O_3517,N_49598,N_49176);
or UO_3518 (O_3518,N_49601,N_49309);
or UO_3519 (O_3519,N_49378,N_49237);
or UO_3520 (O_3520,N_49671,N_49141);
xnor UO_3521 (O_3521,N_49731,N_49072);
xnor UO_3522 (O_3522,N_49944,N_49712);
xnor UO_3523 (O_3523,N_49560,N_49269);
nand UO_3524 (O_3524,N_49387,N_49377);
and UO_3525 (O_3525,N_49532,N_49560);
nor UO_3526 (O_3526,N_49819,N_49553);
nand UO_3527 (O_3527,N_49346,N_49958);
or UO_3528 (O_3528,N_49592,N_49622);
and UO_3529 (O_3529,N_49680,N_49429);
or UO_3530 (O_3530,N_49326,N_49019);
nor UO_3531 (O_3531,N_49794,N_49032);
or UO_3532 (O_3532,N_49817,N_49746);
nor UO_3533 (O_3533,N_49249,N_49382);
or UO_3534 (O_3534,N_49437,N_49542);
and UO_3535 (O_3535,N_49059,N_49504);
or UO_3536 (O_3536,N_49146,N_49742);
nand UO_3537 (O_3537,N_49408,N_49642);
xor UO_3538 (O_3538,N_49772,N_49370);
nor UO_3539 (O_3539,N_49661,N_49214);
xnor UO_3540 (O_3540,N_49104,N_49146);
or UO_3541 (O_3541,N_49243,N_49414);
or UO_3542 (O_3542,N_49867,N_49023);
and UO_3543 (O_3543,N_49736,N_49510);
nor UO_3544 (O_3544,N_49756,N_49004);
xor UO_3545 (O_3545,N_49483,N_49430);
and UO_3546 (O_3546,N_49182,N_49172);
or UO_3547 (O_3547,N_49810,N_49316);
nand UO_3548 (O_3548,N_49693,N_49882);
nor UO_3549 (O_3549,N_49367,N_49354);
xor UO_3550 (O_3550,N_49542,N_49865);
and UO_3551 (O_3551,N_49435,N_49057);
xnor UO_3552 (O_3552,N_49190,N_49640);
nor UO_3553 (O_3553,N_49230,N_49394);
or UO_3554 (O_3554,N_49267,N_49961);
xnor UO_3555 (O_3555,N_49691,N_49872);
and UO_3556 (O_3556,N_49429,N_49801);
nand UO_3557 (O_3557,N_49382,N_49606);
nor UO_3558 (O_3558,N_49126,N_49757);
nor UO_3559 (O_3559,N_49881,N_49202);
or UO_3560 (O_3560,N_49500,N_49706);
nand UO_3561 (O_3561,N_49739,N_49633);
or UO_3562 (O_3562,N_49645,N_49454);
or UO_3563 (O_3563,N_49737,N_49509);
nor UO_3564 (O_3564,N_49418,N_49056);
nand UO_3565 (O_3565,N_49613,N_49297);
nand UO_3566 (O_3566,N_49904,N_49694);
nor UO_3567 (O_3567,N_49561,N_49219);
nand UO_3568 (O_3568,N_49607,N_49401);
nor UO_3569 (O_3569,N_49149,N_49377);
nand UO_3570 (O_3570,N_49723,N_49878);
nand UO_3571 (O_3571,N_49974,N_49072);
and UO_3572 (O_3572,N_49500,N_49473);
nor UO_3573 (O_3573,N_49974,N_49388);
or UO_3574 (O_3574,N_49294,N_49674);
xnor UO_3575 (O_3575,N_49989,N_49059);
nand UO_3576 (O_3576,N_49947,N_49961);
or UO_3577 (O_3577,N_49283,N_49515);
nand UO_3578 (O_3578,N_49533,N_49319);
nand UO_3579 (O_3579,N_49716,N_49157);
nand UO_3580 (O_3580,N_49341,N_49346);
or UO_3581 (O_3581,N_49629,N_49252);
or UO_3582 (O_3582,N_49442,N_49015);
nand UO_3583 (O_3583,N_49368,N_49382);
nand UO_3584 (O_3584,N_49492,N_49860);
or UO_3585 (O_3585,N_49897,N_49620);
or UO_3586 (O_3586,N_49454,N_49202);
nand UO_3587 (O_3587,N_49966,N_49745);
and UO_3588 (O_3588,N_49566,N_49236);
nand UO_3589 (O_3589,N_49720,N_49122);
nand UO_3590 (O_3590,N_49304,N_49202);
xnor UO_3591 (O_3591,N_49189,N_49126);
and UO_3592 (O_3592,N_49939,N_49402);
nand UO_3593 (O_3593,N_49705,N_49594);
nand UO_3594 (O_3594,N_49896,N_49438);
and UO_3595 (O_3595,N_49527,N_49035);
nor UO_3596 (O_3596,N_49043,N_49315);
nor UO_3597 (O_3597,N_49374,N_49616);
nand UO_3598 (O_3598,N_49900,N_49794);
and UO_3599 (O_3599,N_49426,N_49931);
nand UO_3600 (O_3600,N_49887,N_49234);
nand UO_3601 (O_3601,N_49134,N_49581);
nand UO_3602 (O_3602,N_49428,N_49797);
nand UO_3603 (O_3603,N_49746,N_49074);
nor UO_3604 (O_3604,N_49051,N_49655);
or UO_3605 (O_3605,N_49657,N_49333);
nor UO_3606 (O_3606,N_49601,N_49222);
and UO_3607 (O_3607,N_49584,N_49480);
nand UO_3608 (O_3608,N_49692,N_49556);
nand UO_3609 (O_3609,N_49353,N_49476);
or UO_3610 (O_3610,N_49010,N_49084);
nor UO_3611 (O_3611,N_49852,N_49379);
xor UO_3612 (O_3612,N_49314,N_49184);
nor UO_3613 (O_3613,N_49973,N_49601);
xor UO_3614 (O_3614,N_49485,N_49698);
and UO_3615 (O_3615,N_49906,N_49320);
nand UO_3616 (O_3616,N_49567,N_49318);
xor UO_3617 (O_3617,N_49657,N_49788);
and UO_3618 (O_3618,N_49913,N_49803);
xor UO_3619 (O_3619,N_49249,N_49497);
or UO_3620 (O_3620,N_49754,N_49295);
or UO_3621 (O_3621,N_49476,N_49838);
nor UO_3622 (O_3622,N_49700,N_49001);
or UO_3623 (O_3623,N_49711,N_49743);
nand UO_3624 (O_3624,N_49892,N_49816);
and UO_3625 (O_3625,N_49243,N_49229);
nand UO_3626 (O_3626,N_49626,N_49939);
or UO_3627 (O_3627,N_49292,N_49642);
xor UO_3628 (O_3628,N_49671,N_49831);
nor UO_3629 (O_3629,N_49795,N_49684);
nand UO_3630 (O_3630,N_49819,N_49107);
nor UO_3631 (O_3631,N_49802,N_49367);
xor UO_3632 (O_3632,N_49572,N_49412);
nor UO_3633 (O_3633,N_49077,N_49918);
nor UO_3634 (O_3634,N_49254,N_49931);
and UO_3635 (O_3635,N_49393,N_49221);
and UO_3636 (O_3636,N_49169,N_49020);
nand UO_3637 (O_3637,N_49654,N_49215);
and UO_3638 (O_3638,N_49694,N_49596);
nor UO_3639 (O_3639,N_49551,N_49477);
and UO_3640 (O_3640,N_49503,N_49175);
nor UO_3641 (O_3641,N_49443,N_49111);
xor UO_3642 (O_3642,N_49713,N_49454);
or UO_3643 (O_3643,N_49014,N_49316);
nand UO_3644 (O_3644,N_49598,N_49565);
nor UO_3645 (O_3645,N_49368,N_49544);
nand UO_3646 (O_3646,N_49329,N_49096);
nand UO_3647 (O_3647,N_49252,N_49121);
and UO_3648 (O_3648,N_49627,N_49989);
and UO_3649 (O_3649,N_49812,N_49664);
nor UO_3650 (O_3650,N_49133,N_49188);
and UO_3651 (O_3651,N_49783,N_49332);
xnor UO_3652 (O_3652,N_49422,N_49928);
nor UO_3653 (O_3653,N_49554,N_49787);
and UO_3654 (O_3654,N_49265,N_49360);
nor UO_3655 (O_3655,N_49616,N_49703);
or UO_3656 (O_3656,N_49020,N_49305);
nand UO_3657 (O_3657,N_49723,N_49616);
and UO_3658 (O_3658,N_49826,N_49387);
nand UO_3659 (O_3659,N_49632,N_49288);
or UO_3660 (O_3660,N_49633,N_49161);
nand UO_3661 (O_3661,N_49510,N_49451);
and UO_3662 (O_3662,N_49738,N_49753);
nor UO_3663 (O_3663,N_49619,N_49669);
nor UO_3664 (O_3664,N_49173,N_49462);
nand UO_3665 (O_3665,N_49413,N_49463);
xor UO_3666 (O_3666,N_49550,N_49029);
nand UO_3667 (O_3667,N_49288,N_49134);
nand UO_3668 (O_3668,N_49958,N_49537);
and UO_3669 (O_3669,N_49033,N_49144);
nand UO_3670 (O_3670,N_49969,N_49215);
nand UO_3671 (O_3671,N_49972,N_49188);
xnor UO_3672 (O_3672,N_49872,N_49741);
xnor UO_3673 (O_3673,N_49380,N_49211);
nor UO_3674 (O_3674,N_49139,N_49972);
nor UO_3675 (O_3675,N_49721,N_49481);
and UO_3676 (O_3676,N_49752,N_49670);
nand UO_3677 (O_3677,N_49048,N_49968);
xnor UO_3678 (O_3678,N_49381,N_49792);
xor UO_3679 (O_3679,N_49433,N_49694);
or UO_3680 (O_3680,N_49969,N_49627);
or UO_3681 (O_3681,N_49153,N_49935);
and UO_3682 (O_3682,N_49440,N_49644);
xnor UO_3683 (O_3683,N_49984,N_49652);
nand UO_3684 (O_3684,N_49852,N_49844);
nand UO_3685 (O_3685,N_49968,N_49803);
or UO_3686 (O_3686,N_49910,N_49384);
xnor UO_3687 (O_3687,N_49935,N_49850);
nor UO_3688 (O_3688,N_49864,N_49164);
nor UO_3689 (O_3689,N_49417,N_49427);
nor UO_3690 (O_3690,N_49985,N_49842);
or UO_3691 (O_3691,N_49817,N_49421);
nor UO_3692 (O_3692,N_49041,N_49576);
xor UO_3693 (O_3693,N_49820,N_49791);
xnor UO_3694 (O_3694,N_49430,N_49915);
and UO_3695 (O_3695,N_49957,N_49659);
xor UO_3696 (O_3696,N_49129,N_49765);
xor UO_3697 (O_3697,N_49579,N_49472);
and UO_3698 (O_3698,N_49381,N_49657);
nand UO_3699 (O_3699,N_49417,N_49823);
or UO_3700 (O_3700,N_49663,N_49509);
xor UO_3701 (O_3701,N_49582,N_49810);
nand UO_3702 (O_3702,N_49993,N_49045);
nand UO_3703 (O_3703,N_49382,N_49389);
nand UO_3704 (O_3704,N_49868,N_49124);
nand UO_3705 (O_3705,N_49550,N_49827);
nand UO_3706 (O_3706,N_49247,N_49408);
or UO_3707 (O_3707,N_49814,N_49895);
nor UO_3708 (O_3708,N_49855,N_49641);
xor UO_3709 (O_3709,N_49323,N_49592);
and UO_3710 (O_3710,N_49264,N_49235);
or UO_3711 (O_3711,N_49860,N_49559);
and UO_3712 (O_3712,N_49503,N_49061);
nand UO_3713 (O_3713,N_49521,N_49419);
xor UO_3714 (O_3714,N_49887,N_49642);
xnor UO_3715 (O_3715,N_49758,N_49049);
nor UO_3716 (O_3716,N_49104,N_49548);
or UO_3717 (O_3717,N_49879,N_49343);
nand UO_3718 (O_3718,N_49035,N_49968);
or UO_3719 (O_3719,N_49712,N_49532);
nor UO_3720 (O_3720,N_49508,N_49647);
nand UO_3721 (O_3721,N_49359,N_49830);
or UO_3722 (O_3722,N_49983,N_49543);
and UO_3723 (O_3723,N_49854,N_49388);
xor UO_3724 (O_3724,N_49019,N_49053);
or UO_3725 (O_3725,N_49784,N_49723);
nor UO_3726 (O_3726,N_49411,N_49314);
nand UO_3727 (O_3727,N_49171,N_49188);
or UO_3728 (O_3728,N_49471,N_49956);
xnor UO_3729 (O_3729,N_49250,N_49114);
and UO_3730 (O_3730,N_49557,N_49429);
or UO_3731 (O_3731,N_49263,N_49952);
nor UO_3732 (O_3732,N_49338,N_49066);
xor UO_3733 (O_3733,N_49000,N_49905);
nand UO_3734 (O_3734,N_49211,N_49885);
and UO_3735 (O_3735,N_49955,N_49180);
nand UO_3736 (O_3736,N_49357,N_49140);
or UO_3737 (O_3737,N_49355,N_49953);
nor UO_3738 (O_3738,N_49142,N_49280);
xor UO_3739 (O_3739,N_49242,N_49573);
xnor UO_3740 (O_3740,N_49893,N_49887);
or UO_3741 (O_3741,N_49869,N_49875);
nand UO_3742 (O_3742,N_49972,N_49304);
and UO_3743 (O_3743,N_49451,N_49570);
and UO_3744 (O_3744,N_49643,N_49750);
nor UO_3745 (O_3745,N_49820,N_49144);
nand UO_3746 (O_3746,N_49971,N_49213);
nor UO_3747 (O_3747,N_49419,N_49912);
xor UO_3748 (O_3748,N_49780,N_49739);
nand UO_3749 (O_3749,N_49645,N_49614);
xor UO_3750 (O_3750,N_49570,N_49005);
nor UO_3751 (O_3751,N_49241,N_49343);
nand UO_3752 (O_3752,N_49591,N_49807);
nor UO_3753 (O_3753,N_49383,N_49077);
nand UO_3754 (O_3754,N_49868,N_49798);
or UO_3755 (O_3755,N_49574,N_49133);
or UO_3756 (O_3756,N_49417,N_49735);
nor UO_3757 (O_3757,N_49039,N_49500);
nor UO_3758 (O_3758,N_49659,N_49503);
nand UO_3759 (O_3759,N_49509,N_49456);
nand UO_3760 (O_3760,N_49703,N_49183);
or UO_3761 (O_3761,N_49083,N_49478);
xor UO_3762 (O_3762,N_49380,N_49546);
nor UO_3763 (O_3763,N_49857,N_49910);
and UO_3764 (O_3764,N_49856,N_49562);
nand UO_3765 (O_3765,N_49280,N_49748);
or UO_3766 (O_3766,N_49864,N_49895);
xor UO_3767 (O_3767,N_49553,N_49018);
or UO_3768 (O_3768,N_49074,N_49197);
and UO_3769 (O_3769,N_49966,N_49503);
nand UO_3770 (O_3770,N_49437,N_49846);
or UO_3771 (O_3771,N_49557,N_49929);
nor UO_3772 (O_3772,N_49261,N_49988);
xor UO_3773 (O_3773,N_49242,N_49337);
nor UO_3774 (O_3774,N_49316,N_49795);
or UO_3775 (O_3775,N_49620,N_49588);
nor UO_3776 (O_3776,N_49942,N_49246);
or UO_3777 (O_3777,N_49018,N_49416);
or UO_3778 (O_3778,N_49880,N_49654);
nand UO_3779 (O_3779,N_49420,N_49233);
xnor UO_3780 (O_3780,N_49684,N_49101);
xor UO_3781 (O_3781,N_49750,N_49063);
nand UO_3782 (O_3782,N_49935,N_49700);
or UO_3783 (O_3783,N_49726,N_49426);
xnor UO_3784 (O_3784,N_49923,N_49805);
xnor UO_3785 (O_3785,N_49073,N_49223);
or UO_3786 (O_3786,N_49238,N_49318);
and UO_3787 (O_3787,N_49253,N_49386);
xor UO_3788 (O_3788,N_49640,N_49085);
nand UO_3789 (O_3789,N_49079,N_49512);
nor UO_3790 (O_3790,N_49576,N_49736);
xor UO_3791 (O_3791,N_49309,N_49782);
and UO_3792 (O_3792,N_49731,N_49812);
and UO_3793 (O_3793,N_49032,N_49897);
nor UO_3794 (O_3794,N_49860,N_49200);
xor UO_3795 (O_3795,N_49060,N_49297);
xnor UO_3796 (O_3796,N_49250,N_49840);
and UO_3797 (O_3797,N_49266,N_49350);
or UO_3798 (O_3798,N_49195,N_49417);
or UO_3799 (O_3799,N_49218,N_49804);
xor UO_3800 (O_3800,N_49480,N_49623);
or UO_3801 (O_3801,N_49942,N_49843);
nor UO_3802 (O_3802,N_49682,N_49468);
nand UO_3803 (O_3803,N_49566,N_49722);
or UO_3804 (O_3804,N_49412,N_49754);
nand UO_3805 (O_3805,N_49908,N_49019);
nand UO_3806 (O_3806,N_49760,N_49134);
xnor UO_3807 (O_3807,N_49256,N_49073);
nand UO_3808 (O_3808,N_49380,N_49900);
or UO_3809 (O_3809,N_49700,N_49151);
xnor UO_3810 (O_3810,N_49792,N_49659);
xnor UO_3811 (O_3811,N_49538,N_49213);
and UO_3812 (O_3812,N_49361,N_49730);
and UO_3813 (O_3813,N_49619,N_49087);
nand UO_3814 (O_3814,N_49218,N_49785);
or UO_3815 (O_3815,N_49604,N_49726);
and UO_3816 (O_3816,N_49689,N_49910);
nor UO_3817 (O_3817,N_49633,N_49838);
xnor UO_3818 (O_3818,N_49481,N_49343);
or UO_3819 (O_3819,N_49461,N_49640);
nand UO_3820 (O_3820,N_49683,N_49275);
xor UO_3821 (O_3821,N_49269,N_49548);
and UO_3822 (O_3822,N_49477,N_49157);
nand UO_3823 (O_3823,N_49190,N_49842);
nand UO_3824 (O_3824,N_49419,N_49144);
or UO_3825 (O_3825,N_49040,N_49088);
nand UO_3826 (O_3826,N_49547,N_49241);
nand UO_3827 (O_3827,N_49791,N_49007);
nand UO_3828 (O_3828,N_49078,N_49238);
nor UO_3829 (O_3829,N_49892,N_49449);
xnor UO_3830 (O_3830,N_49700,N_49334);
and UO_3831 (O_3831,N_49346,N_49137);
and UO_3832 (O_3832,N_49317,N_49883);
xor UO_3833 (O_3833,N_49938,N_49620);
xnor UO_3834 (O_3834,N_49648,N_49079);
and UO_3835 (O_3835,N_49330,N_49025);
and UO_3836 (O_3836,N_49839,N_49936);
xor UO_3837 (O_3837,N_49230,N_49715);
xnor UO_3838 (O_3838,N_49149,N_49000);
nor UO_3839 (O_3839,N_49029,N_49131);
xnor UO_3840 (O_3840,N_49199,N_49533);
or UO_3841 (O_3841,N_49234,N_49079);
xnor UO_3842 (O_3842,N_49328,N_49158);
and UO_3843 (O_3843,N_49411,N_49218);
xnor UO_3844 (O_3844,N_49575,N_49829);
xor UO_3845 (O_3845,N_49808,N_49622);
nand UO_3846 (O_3846,N_49577,N_49612);
nor UO_3847 (O_3847,N_49233,N_49642);
nand UO_3848 (O_3848,N_49699,N_49351);
and UO_3849 (O_3849,N_49293,N_49287);
xnor UO_3850 (O_3850,N_49854,N_49337);
or UO_3851 (O_3851,N_49818,N_49738);
xnor UO_3852 (O_3852,N_49053,N_49377);
nand UO_3853 (O_3853,N_49064,N_49780);
nor UO_3854 (O_3854,N_49490,N_49916);
or UO_3855 (O_3855,N_49150,N_49470);
xor UO_3856 (O_3856,N_49315,N_49032);
xor UO_3857 (O_3857,N_49418,N_49722);
nor UO_3858 (O_3858,N_49919,N_49052);
nand UO_3859 (O_3859,N_49585,N_49696);
or UO_3860 (O_3860,N_49729,N_49635);
and UO_3861 (O_3861,N_49783,N_49485);
nand UO_3862 (O_3862,N_49670,N_49410);
and UO_3863 (O_3863,N_49345,N_49239);
nand UO_3864 (O_3864,N_49424,N_49236);
and UO_3865 (O_3865,N_49046,N_49120);
or UO_3866 (O_3866,N_49884,N_49873);
nand UO_3867 (O_3867,N_49220,N_49450);
nor UO_3868 (O_3868,N_49412,N_49946);
and UO_3869 (O_3869,N_49760,N_49261);
nand UO_3870 (O_3870,N_49465,N_49161);
or UO_3871 (O_3871,N_49454,N_49080);
and UO_3872 (O_3872,N_49186,N_49760);
and UO_3873 (O_3873,N_49231,N_49817);
and UO_3874 (O_3874,N_49940,N_49838);
xnor UO_3875 (O_3875,N_49464,N_49638);
xor UO_3876 (O_3876,N_49215,N_49725);
or UO_3877 (O_3877,N_49525,N_49364);
and UO_3878 (O_3878,N_49252,N_49594);
xnor UO_3879 (O_3879,N_49884,N_49700);
nand UO_3880 (O_3880,N_49997,N_49840);
and UO_3881 (O_3881,N_49107,N_49267);
and UO_3882 (O_3882,N_49666,N_49056);
nor UO_3883 (O_3883,N_49185,N_49338);
nand UO_3884 (O_3884,N_49025,N_49442);
nor UO_3885 (O_3885,N_49058,N_49839);
xor UO_3886 (O_3886,N_49935,N_49258);
nand UO_3887 (O_3887,N_49867,N_49024);
nand UO_3888 (O_3888,N_49192,N_49388);
or UO_3889 (O_3889,N_49534,N_49146);
nand UO_3890 (O_3890,N_49613,N_49953);
nand UO_3891 (O_3891,N_49593,N_49040);
and UO_3892 (O_3892,N_49021,N_49435);
nand UO_3893 (O_3893,N_49207,N_49683);
nor UO_3894 (O_3894,N_49386,N_49746);
or UO_3895 (O_3895,N_49153,N_49000);
or UO_3896 (O_3896,N_49086,N_49491);
nand UO_3897 (O_3897,N_49563,N_49859);
nand UO_3898 (O_3898,N_49586,N_49600);
nand UO_3899 (O_3899,N_49806,N_49821);
nand UO_3900 (O_3900,N_49355,N_49737);
and UO_3901 (O_3901,N_49320,N_49933);
xor UO_3902 (O_3902,N_49630,N_49596);
xnor UO_3903 (O_3903,N_49024,N_49480);
xnor UO_3904 (O_3904,N_49015,N_49200);
nor UO_3905 (O_3905,N_49961,N_49703);
nand UO_3906 (O_3906,N_49564,N_49707);
xnor UO_3907 (O_3907,N_49221,N_49964);
and UO_3908 (O_3908,N_49019,N_49686);
nor UO_3909 (O_3909,N_49477,N_49160);
and UO_3910 (O_3910,N_49383,N_49573);
xnor UO_3911 (O_3911,N_49246,N_49658);
or UO_3912 (O_3912,N_49978,N_49287);
or UO_3913 (O_3913,N_49902,N_49120);
nand UO_3914 (O_3914,N_49140,N_49613);
or UO_3915 (O_3915,N_49385,N_49703);
xor UO_3916 (O_3916,N_49587,N_49871);
and UO_3917 (O_3917,N_49289,N_49908);
or UO_3918 (O_3918,N_49992,N_49080);
and UO_3919 (O_3919,N_49249,N_49600);
or UO_3920 (O_3920,N_49951,N_49298);
nor UO_3921 (O_3921,N_49142,N_49336);
nand UO_3922 (O_3922,N_49352,N_49060);
xor UO_3923 (O_3923,N_49384,N_49107);
or UO_3924 (O_3924,N_49875,N_49522);
and UO_3925 (O_3925,N_49881,N_49812);
nor UO_3926 (O_3926,N_49526,N_49360);
nand UO_3927 (O_3927,N_49709,N_49668);
nor UO_3928 (O_3928,N_49154,N_49996);
nor UO_3929 (O_3929,N_49255,N_49732);
or UO_3930 (O_3930,N_49062,N_49352);
xor UO_3931 (O_3931,N_49471,N_49091);
nor UO_3932 (O_3932,N_49504,N_49057);
nor UO_3933 (O_3933,N_49998,N_49601);
xnor UO_3934 (O_3934,N_49954,N_49874);
nand UO_3935 (O_3935,N_49169,N_49513);
xnor UO_3936 (O_3936,N_49515,N_49031);
nand UO_3937 (O_3937,N_49840,N_49957);
nand UO_3938 (O_3938,N_49416,N_49409);
nand UO_3939 (O_3939,N_49485,N_49891);
or UO_3940 (O_3940,N_49009,N_49725);
nor UO_3941 (O_3941,N_49636,N_49873);
or UO_3942 (O_3942,N_49210,N_49003);
nand UO_3943 (O_3943,N_49336,N_49132);
nand UO_3944 (O_3944,N_49279,N_49784);
nand UO_3945 (O_3945,N_49466,N_49498);
and UO_3946 (O_3946,N_49563,N_49504);
nor UO_3947 (O_3947,N_49568,N_49547);
nand UO_3948 (O_3948,N_49609,N_49481);
xor UO_3949 (O_3949,N_49489,N_49866);
nor UO_3950 (O_3950,N_49262,N_49963);
or UO_3951 (O_3951,N_49696,N_49088);
nor UO_3952 (O_3952,N_49727,N_49760);
or UO_3953 (O_3953,N_49647,N_49027);
nor UO_3954 (O_3954,N_49058,N_49262);
nor UO_3955 (O_3955,N_49089,N_49432);
nand UO_3956 (O_3956,N_49690,N_49972);
nor UO_3957 (O_3957,N_49614,N_49380);
or UO_3958 (O_3958,N_49630,N_49200);
or UO_3959 (O_3959,N_49768,N_49512);
and UO_3960 (O_3960,N_49364,N_49560);
or UO_3961 (O_3961,N_49809,N_49736);
nand UO_3962 (O_3962,N_49694,N_49319);
and UO_3963 (O_3963,N_49454,N_49419);
and UO_3964 (O_3964,N_49581,N_49460);
nor UO_3965 (O_3965,N_49222,N_49730);
and UO_3966 (O_3966,N_49507,N_49771);
nand UO_3967 (O_3967,N_49203,N_49398);
xnor UO_3968 (O_3968,N_49393,N_49987);
or UO_3969 (O_3969,N_49230,N_49691);
and UO_3970 (O_3970,N_49218,N_49432);
and UO_3971 (O_3971,N_49520,N_49145);
xor UO_3972 (O_3972,N_49052,N_49221);
and UO_3973 (O_3973,N_49884,N_49128);
and UO_3974 (O_3974,N_49987,N_49504);
nand UO_3975 (O_3975,N_49135,N_49872);
and UO_3976 (O_3976,N_49735,N_49126);
or UO_3977 (O_3977,N_49378,N_49951);
nand UO_3978 (O_3978,N_49098,N_49496);
or UO_3979 (O_3979,N_49181,N_49270);
xor UO_3980 (O_3980,N_49357,N_49041);
nand UO_3981 (O_3981,N_49077,N_49536);
xnor UO_3982 (O_3982,N_49706,N_49051);
and UO_3983 (O_3983,N_49837,N_49844);
or UO_3984 (O_3984,N_49412,N_49311);
xor UO_3985 (O_3985,N_49221,N_49528);
and UO_3986 (O_3986,N_49070,N_49084);
or UO_3987 (O_3987,N_49483,N_49606);
xor UO_3988 (O_3988,N_49527,N_49118);
nor UO_3989 (O_3989,N_49549,N_49836);
and UO_3990 (O_3990,N_49600,N_49930);
nor UO_3991 (O_3991,N_49645,N_49816);
nand UO_3992 (O_3992,N_49450,N_49629);
and UO_3993 (O_3993,N_49319,N_49395);
xor UO_3994 (O_3994,N_49141,N_49050);
or UO_3995 (O_3995,N_49446,N_49143);
and UO_3996 (O_3996,N_49003,N_49610);
nand UO_3997 (O_3997,N_49980,N_49571);
nor UO_3998 (O_3998,N_49018,N_49348);
and UO_3999 (O_3999,N_49928,N_49283);
nor UO_4000 (O_4000,N_49605,N_49375);
nand UO_4001 (O_4001,N_49396,N_49499);
xor UO_4002 (O_4002,N_49203,N_49023);
and UO_4003 (O_4003,N_49884,N_49627);
xnor UO_4004 (O_4004,N_49233,N_49941);
nor UO_4005 (O_4005,N_49325,N_49796);
or UO_4006 (O_4006,N_49850,N_49691);
nor UO_4007 (O_4007,N_49143,N_49108);
and UO_4008 (O_4008,N_49039,N_49417);
and UO_4009 (O_4009,N_49890,N_49623);
or UO_4010 (O_4010,N_49375,N_49929);
nand UO_4011 (O_4011,N_49303,N_49464);
nor UO_4012 (O_4012,N_49780,N_49220);
nor UO_4013 (O_4013,N_49002,N_49048);
xor UO_4014 (O_4014,N_49716,N_49995);
or UO_4015 (O_4015,N_49231,N_49186);
nand UO_4016 (O_4016,N_49219,N_49294);
nand UO_4017 (O_4017,N_49044,N_49824);
and UO_4018 (O_4018,N_49572,N_49636);
nor UO_4019 (O_4019,N_49733,N_49131);
xnor UO_4020 (O_4020,N_49245,N_49466);
or UO_4021 (O_4021,N_49490,N_49742);
or UO_4022 (O_4022,N_49439,N_49676);
nor UO_4023 (O_4023,N_49129,N_49590);
xnor UO_4024 (O_4024,N_49501,N_49839);
xor UO_4025 (O_4025,N_49142,N_49532);
nand UO_4026 (O_4026,N_49309,N_49112);
xor UO_4027 (O_4027,N_49559,N_49823);
nor UO_4028 (O_4028,N_49650,N_49352);
xor UO_4029 (O_4029,N_49635,N_49374);
or UO_4030 (O_4030,N_49150,N_49851);
nand UO_4031 (O_4031,N_49313,N_49828);
nand UO_4032 (O_4032,N_49032,N_49292);
or UO_4033 (O_4033,N_49779,N_49480);
xnor UO_4034 (O_4034,N_49947,N_49921);
nand UO_4035 (O_4035,N_49492,N_49907);
nand UO_4036 (O_4036,N_49304,N_49333);
nor UO_4037 (O_4037,N_49020,N_49746);
nand UO_4038 (O_4038,N_49343,N_49637);
and UO_4039 (O_4039,N_49792,N_49586);
xnor UO_4040 (O_4040,N_49292,N_49921);
or UO_4041 (O_4041,N_49609,N_49916);
xnor UO_4042 (O_4042,N_49422,N_49353);
or UO_4043 (O_4043,N_49757,N_49476);
or UO_4044 (O_4044,N_49669,N_49468);
and UO_4045 (O_4045,N_49506,N_49690);
xnor UO_4046 (O_4046,N_49418,N_49187);
nor UO_4047 (O_4047,N_49634,N_49614);
xor UO_4048 (O_4048,N_49167,N_49678);
and UO_4049 (O_4049,N_49443,N_49286);
xnor UO_4050 (O_4050,N_49010,N_49570);
nor UO_4051 (O_4051,N_49740,N_49402);
nor UO_4052 (O_4052,N_49996,N_49302);
nor UO_4053 (O_4053,N_49246,N_49475);
or UO_4054 (O_4054,N_49863,N_49216);
nor UO_4055 (O_4055,N_49592,N_49920);
or UO_4056 (O_4056,N_49317,N_49394);
nand UO_4057 (O_4057,N_49283,N_49332);
and UO_4058 (O_4058,N_49136,N_49427);
xnor UO_4059 (O_4059,N_49969,N_49948);
nand UO_4060 (O_4060,N_49624,N_49936);
or UO_4061 (O_4061,N_49803,N_49594);
or UO_4062 (O_4062,N_49230,N_49990);
nand UO_4063 (O_4063,N_49899,N_49235);
nand UO_4064 (O_4064,N_49861,N_49772);
xor UO_4065 (O_4065,N_49572,N_49354);
xnor UO_4066 (O_4066,N_49332,N_49602);
and UO_4067 (O_4067,N_49315,N_49194);
and UO_4068 (O_4068,N_49003,N_49041);
xnor UO_4069 (O_4069,N_49900,N_49229);
and UO_4070 (O_4070,N_49548,N_49949);
nand UO_4071 (O_4071,N_49334,N_49141);
xnor UO_4072 (O_4072,N_49524,N_49298);
and UO_4073 (O_4073,N_49744,N_49197);
or UO_4074 (O_4074,N_49711,N_49572);
xor UO_4075 (O_4075,N_49858,N_49375);
nand UO_4076 (O_4076,N_49461,N_49469);
nand UO_4077 (O_4077,N_49797,N_49560);
xnor UO_4078 (O_4078,N_49867,N_49481);
nand UO_4079 (O_4079,N_49906,N_49292);
nor UO_4080 (O_4080,N_49036,N_49054);
and UO_4081 (O_4081,N_49374,N_49103);
nand UO_4082 (O_4082,N_49042,N_49948);
nor UO_4083 (O_4083,N_49277,N_49714);
nor UO_4084 (O_4084,N_49817,N_49053);
or UO_4085 (O_4085,N_49336,N_49426);
nor UO_4086 (O_4086,N_49265,N_49342);
xor UO_4087 (O_4087,N_49150,N_49266);
xnor UO_4088 (O_4088,N_49809,N_49399);
or UO_4089 (O_4089,N_49432,N_49530);
nor UO_4090 (O_4090,N_49671,N_49711);
xor UO_4091 (O_4091,N_49532,N_49290);
and UO_4092 (O_4092,N_49963,N_49661);
nand UO_4093 (O_4093,N_49992,N_49348);
and UO_4094 (O_4094,N_49316,N_49239);
nor UO_4095 (O_4095,N_49794,N_49940);
xnor UO_4096 (O_4096,N_49175,N_49386);
nand UO_4097 (O_4097,N_49848,N_49498);
and UO_4098 (O_4098,N_49553,N_49773);
nor UO_4099 (O_4099,N_49234,N_49359);
xnor UO_4100 (O_4100,N_49267,N_49596);
nor UO_4101 (O_4101,N_49450,N_49019);
nor UO_4102 (O_4102,N_49597,N_49596);
or UO_4103 (O_4103,N_49188,N_49663);
nor UO_4104 (O_4104,N_49646,N_49218);
nand UO_4105 (O_4105,N_49839,N_49960);
or UO_4106 (O_4106,N_49854,N_49417);
nor UO_4107 (O_4107,N_49748,N_49979);
nor UO_4108 (O_4108,N_49284,N_49460);
xor UO_4109 (O_4109,N_49281,N_49910);
and UO_4110 (O_4110,N_49129,N_49994);
nor UO_4111 (O_4111,N_49074,N_49317);
nand UO_4112 (O_4112,N_49814,N_49820);
nor UO_4113 (O_4113,N_49101,N_49685);
xor UO_4114 (O_4114,N_49907,N_49841);
or UO_4115 (O_4115,N_49946,N_49683);
xor UO_4116 (O_4116,N_49797,N_49111);
and UO_4117 (O_4117,N_49906,N_49717);
and UO_4118 (O_4118,N_49957,N_49148);
and UO_4119 (O_4119,N_49160,N_49964);
or UO_4120 (O_4120,N_49925,N_49575);
or UO_4121 (O_4121,N_49880,N_49460);
or UO_4122 (O_4122,N_49711,N_49086);
or UO_4123 (O_4123,N_49551,N_49238);
nor UO_4124 (O_4124,N_49442,N_49512);
xor UO_4125 (O_4125,N_49625,N_49599);
and UO_4126 (O_4126,N_49593,N_49185);
xor UO_4127 (O_4127,N_49011,N_49064);
xor UO_4128 (O_4128,N_49787,N_49291);
nand UO_4129 (O_4129,N_49210,N_49484);
nand UO_4130 (O_4130,N_49269,N_49518);
or UO_4131 (O_4131,N_49771,N_49639);
and UO_4132 (O_4132,N_49469,N_49890);
nor UO_4133 (O_4133,N_49548,N_49927);
and UO_4134 (O_4134,N_49942,N_49138);
and UO_4135 (O_4135,N_49492,N_49618);
nand UO_4136 (O_4136,N_49272,N_49938);
and UO_4137 (O_4137,N_49540,N_49598);
nand UO_4138 (O_4138,N_49642,N_49444);
or UO_4139 (O_4139,N_49662,N_49496);
and UO_4140 (O_4140,N_49757,N_49172);
nand UO_4141 (O_4141,N_49531,N_49116);
or UO_4142 (O_4142,N_49661,N_49729);
nand UO_4143 (O_4143,N_49247,N_49364);
nand UO_4144 (O_4144,N_49180,N_49145);
or UO_4145 (O_4145,N_49471,N_49431);
xnor UO_4146 (O_4146,N_49859,N_49392);
xnor UO_4147 (O_4147,N_49892,N_49743);
xnor UO_4148 (O_4148,N_49253,N_49781);
and UO_4149 (O_4149,N_49876,N_49370);
nor UO_4150 (O_4150,N_49713,N_49559);
and UO_4151 (O_4151,N_49000,N_49143);
nor UO_4152 (O_4152,N_49068,N_49390);
and UO_4153 (O_4153,N_49142,N_49259);
and UO_4154 (O_4154,N_49655,N_49889);
xnor UO_4155 (O_4155,N_49481,N_49727);
xnor UO_4156 (O_4156,N_49436,N_49832);
or UO_4157 (O_4157,N_49544,N_49638);
nor UO_4158 (O_4158,N_49764,N_49739);
and UO_4159 (O_4159,N_49907,N_49697);
or UO_4160 (O_4160,N_49535,N_49694);
nor UO_4161 (O_4161,N_49279,N_49700);
nand UO_4162 (O_4162,N_49555,N_49446);
nand UO_4163 (O_4163,N_49787,N_49010);
xor UO_4164 (O_4164,N_49543,N_49743);
or UO_4165 (O_4165,N_49549,N_49559);
or UO_4166 (O_4166,N_49547,N_49777);
nor UO_4167 (O_4167,N_49356,N_49585);
nand UO_4168 (O_4168,N_49138,N_49067);
or UO_4169 (O_4169,N_49061,N_49486);
xnor UO_4170 (O_4170,N_49225,N_49375);
and UO_4171 (O_4171,N_49754,N_49477);
nor UO_4172 (O_4172,N_49479,N_49395);
nand UO_4173 (O_4173,N_49419,N_49987);
and UO_4174 (O_4174,N_49386,N_49536);
and UO_4175 (O_4175,N_49465,N_49524);
xor UO_4176 (O_4176,N_49084,N_49686);
nor UO_4177 (O_4177,N_49826,N_49049);
and UO_4178 (O_4178,N_49541,N_49140);
or UO_4179 (O_4179,N_49497,N_49734);
or UO_4180 (O_4180,N_49672,N_49615);
nand UO_4181 (O_4181,N_49050,N_49710);
or UO_4182 (O_4182,N_49251,N_49076);
nor UO_4183 (O_4183,N_49486,N_49695);
xnor UO_4184 (O_4184,N_49624,N_49090);
xnor UO_4185 (O_4185,N_49283,N_49878);
xnor UO_4186 (O_4186,N_49819,N_49413);
xnor UO_4187 (O_4187,N_49416,N_49346);
xor UO_4188 (O_4188,N_49895,N_49198);
and UO_4189 (O_4189,N_49323,N_49719);
or UO_4190 (O_4190,N_49971,N_49642);
or UO_4191 (O_4191,N_49523,N_49743);
or UO_4192 (O_4192,N_49366,N_49828);
nor UO_4193 (O_4193,N_49286,N_49709);
or UO_4194 (O_4194,N_49537,N_49414);
and UO_4195 (O_4195,N_49206,N_49844);
and UO_4196 (O_4196,N_49379,N_49802);
nor UO_4197 (O_4197,N_49005,N_49841);
nor UO_4198 (O_4198,N_49671,N_49051);
nor UO_4199 (O_4199,N_49617,N_49099);
nand UO_4200 (O_4200,N_49416,N_49108);
nor UO_4201 (O_4201,N_49436,N_49820);
and UO_4202 (O_4202,N_49581,N_49099);
nand UO_4203 (O_4203,N_49649,N_49281);
and UO_4204 (O_4204,N_49697,N_49126);
or UO_4205 (O_4205,N_49218,N_49704);
xor UO_4206 (O_4206,N_49309,N_49727);
nor UO_4207 (O_4207,N_49266,N_49922);
and UO_4208 (O_4208,N_49359,N_49573);
nor UO_4209 (O_4209,N_49999,N_49580);
or UO_4210 (O_4210,N_49116,N_49089);
xnor UO_4211 (O_4211,N_49985,N_49890);
nand UO_4212 (O_4212,N_49411,N_49950);
and UO_4213 (O_4213,N_49103,N_49016);
nand UO_4214 (O_4214,N_49709,N_49721);
and UO_4215 (O_4215,N_49867,N_49254);
and UO_4216 (O_4216,N_49993,N_49386);
nand UO_4217 (O_4217,N_49244,N_49319);
nand UO_4218 (O_4218,N_49257,N_49895);
and UO_4219 (O_4219,N_49997,N_49516);
nor UO_4220 (O_4220,N_49956,N_49856);
nor UO_4221 (O_4221,N_49277,N_49323);
or UO_4222 (O_4222,N_49329,N_49135);
nand UO_4223 (O_4223,N_49970,N_49197);
nand UO_4224 (O_4224,N_49268,N_49725);
or UO_4225 (O_4225,N_49012,N_49224);
nor UO_4226 (O_4226,N_49048,N_49153);
and UO_4227 (O_4227,N_49367,N_49355);
nor UO_4228 (O_4228,N_49849,N_49155);
nand UO_4229 (O_4229,N_49160,N_49021);
nand UO_4230 (O_4230,N_49278,N_49173);
or UO_4231 (O_4231,N_49182,N_49796);
and UO_4232 (O_4232,N_49111,N_49234);
nor UO_4233 (O_4233,N_49918,N_49644);
nand UO_4234 (O_4234,N_49494,N_49278);
nor UO_4235 (O_4235,N_49967,N_49136);
xnor UO_4236 (O_4236,N_49683,N_49625);
xor UO_4237 (O_4237,N_49162,N_49286);
nand UO_4238 (O_4238,N_49785,N_49392);
nand UO_4239 (O_4239,N_49431,N_49067);
xor UO_4240 (O_4240,N_49871,N_49887);
and UO_4241 (O_4241,N_49497,N_49063);
nand UO_4242 (O_4242,N_49500,N_49579);
nor UO_4243 (O_4243,N_49744,N_49864);
xor UO_4244 (O_4244,N_49323,N_49618);
and UO_4245 (O_4245,N_49203,N_49945);
nand UO_4246 (O_4246,N_49689,N_49095);
xnor UO_4247 (O_4247,N_49909,N_49309);
nor UO_4248 (O_4248,N_49449,N_49804);
xnor UO_4249 (O_4249,N_49342,N_49872);
or UO_4250 (O_4250,N_49901,N_49030);
nand UO_4251 (O_4251,N_49799,N_49942);
xnor UO_4252 (O_4252,N_49466,N_49194);
nor UO_4253 (O_4253,N_49109,N_49146);
nor UO_4254 (O_4254,N_49009,N_49203);
xor UO_4255 (O_4255,N_49455,N_49194);
and UO_4256 (O_4256,N_49373,N_49060);
nor UO_4257 (O_4257,N_49310,N_49535);
xor UO_4258 (O_4258,N_49437,N_49077);
xnor UO_4259 (O_4259,N_49719,N_49361);
nand UO_4260 (O_4260,N_49737,N_49913);
nor UO_4261 (O_4261,N_49016,N_49969);
or UO_4262 (O_4262,N_49859,N_49515);
or UO_4263 (O_4263,N_49787,N_49134);
nor UO_4264 (O_4264,N_49386,N_49842);
nand UO_4265 (O_4265,N_49395,N_49415);
or UO_4266 (O_4266,N_49914,N_49355);
nand UO_4267 (O_4267,N_49138,N_49284);
or UO_4268 (O_4268,N_49540,N_49593);
or UO_4269 (O_4269,N_49325,N_49625);
xnor UO_4270 (O_4270,N_49167,N_49561);
or UO_4271 (O_4271,N_49672,N_49238);
nand UO_4272 (O_4272,N_49513,N_49788);
and UO_4273 (O_4273,N_49641,N_49522);
nand UO_4274 (O_4274,N_49863,N_49091);
nor UO_4275 (O_4275,N_49840,N_49561);
or UO_4276 (O_4276,N_49451,N_49125);
and UO_4277 (O_4277,N_49647,N_49840);
nand UO_4278 (O_4278,N_49558,N_49843);
xnor UO_4279 (O_4279,N_49443,N_49112);
nor UO_4280 (O_4280,N_49858,N_49632);
or UO_4281 (O_4281,N_49791,N_49335);
nor UO_4282 (O_4282,N_49806,N_49612);
nor UO_4283 (O_4283,N_49748,N_49810);
xnor UO_4284 (O_4284,N_49008,N_49370);
xnor UO_4285 (O_4285,N_49457,N_49997);
nand UO_4286 (O_4286,N_49168,N_49895);
and UO_4287 (O_4287,N_49385,N_49831);
xnor UO_4288 (O_4288,N_49620,N_49673);
or UO_4289 (O_4289,N_49942,N_49565);
xnor UO_4290 (O_4290,N_49398,N_49026);
and UO_4291 (O_4291,N_49869,N_49768);
xor UO_4292 (O_4292,N_49413,N_49896);
nand UO_4293 (O_4293,N_49607,N_49066);
or UO_4294 (O_4294,N_49764,N_49322);
nor UO_4295 (O_4295,N_49876,N_49997);
nor UO_4296 (O_4296,N_49376,N_49257);
xor UO_4297 (O_4297,N_49287,N_49938);
and UO_4298 (O_4298,N_49010,N_49692);
xnor UO_4299 (O_4299,N_49511,N_49097);
xor UO_4300 (O_4300,N_49624,N_49697);
xnor UO_4301 (O_4301,N_49577,N_49269);
nand UO_4302 (O_4302,N_49529,N_49736);
or UO_4303 (O_4303,N_49554,N_49164);
or UO_4304 (O_4304,N_49955,N_49563);
nor UO_4305 (O_4305,N_49783,N_49392);
xor UO_4306 (O_4306,N_49351,N_49151);
or UO_4307 (O_4307,N_49304,N_49851);
or UO_4308 (O_4308,N_49216,N_49735);
or UO_4309 (O_4309,N_49916,N_49386);
xnor UO_4310 (O_4310,N_49736,N_49416);
or UO_4311 (O_4311,N_49932,N_49689);
nand UO_4312 (O_4312,N_49439,N_49918);
nor UO_4313 (O_4313,N_49877,N_49077);
xnor UO_4314 (O_4314,N_49994,N_49764);
nor UO_4315 (O_4315,N_49156,N_49602);
xor UO_4316 (O_4316,N_49187,N_49333);
xor UO_4317 (O_4317,N_49566,N_49913);
nor UO_4318 (O_4318,N_49699,N_49901);
nor UO_4319 (O_4319,N_49529,N_49734);
nand UO_4320 (O_4320,N_49425,N_49635);
xor UO_4321 (O_4321,N_49841,N_49715);
and UO_4322 (O_4322,N_49970,N_49041);
nor UO_4323 (O_4323,N_49667,N_49049);
or UO_4324 (O_4324,N_49160,N_49114);
nor UO_4325 (O_4325,N_49044,N_49979);
xnor UO_4326 (O_4326,N_49196,N_49992);
or UO_4327 (O_4327,N_49278,N_49174);
or UO_4328 (O_4328,N_49884,N_49576);
xor UO_4329 (O_4329,N_49103,N_49679);
nand UO_4330 (O_4330,N_49589,N_49565);
or UO_4331 (O_4331,N_49822,N_49688);
xor UO_4332 (O_4332,N_49092,N_49907);
and UO_4333 (O_4333,N_49658,N_49519);
nand UO_4334 (O_4334,N_49942,N_49886);
or UO_4335 (O_4335,N_49936,N_49580);
xnor UO_4336 (O_4336,N_49155,N_49189);
or UO_4337 (O_4337,N_49184,N_49554);
or UO_4338 (O_4338,N_49248,N_49890);
nand UO_4339 (O_4339,N_49650,N_49791);
or UO_4340 (O_4340,N_49000,N_49196);
xnor UO_4341 (O_4341,N_49461,N_49206);
xor UO_4342 (O_4342,N_49316,N_49301);
nand UO_4343 (O_4343,N_49039,N_49506);
nor UO_4344 (O_4344,N_49169,N_49216);
nor UO_4345 (O_4345,N_49433,N_49500);
or UO_4346 (O_4346,N_49849,N_49455);
nand UO_4347 (O_4347,N_49253,N_49883);
or UO_4348 (O_4348,N_49271,N_49747);
and UO_4349 (O_4349,N_49715,N_49309);
xnor UO_4350 (O_4350,N_49342,N_49915);
and UO_4351 (O_4351,N_49008,N_49227);
nor UO_4352 (O_4352,N_49040,N_49199);
nor UO_4353 (O_4353,N_49483,N_49446);
or UO_4354 (O_4354,N_49758,N_49514);
nand UO_4355 (O_4355,N_49643,N_49099);
xnor UO_4356 (O_4356,N_49318,N_49568);
xor UO_4357 (O_4357,N_49283,N_49665);
xor UO_4358 (O_4358,N_49713,N_49201);
nand UO_4359 (O_4359,N_49656,N_49498);
and UO_4360 (O_4360,N_49560,N_49606);
nand UO_4361 (O_4361,N_49961,N_49003);
nor UO_4362 (O_4362,N_49414,N_49909);
nor UO_4363 (O_4363,N_49053,N_49034);
and UO_4364 (O_4364,N_49269,N_49377);
xor UO_4365 (O_4365,N_49211,N_49526);
xnor UO_4366 (O_4366,N_49881,N_49510);
nand UO_4367 (O_4367,N_49372,N_49989);
and UO_4368 (O_4368,N_49455,N_49037);
xor UO_4369 (O_4369,N_49703,N_49431);
and UO_4370 (O_4370,N_49894,N_49723);
nand UO_4371 (O_4371,N_49192,N_49398);
nor UO_4372 (O_4372,N_49773,N_49404);
nand UO_4373 (O_4373,N_49468,N_49210);
xor UO_4374 (O_4374,N_49258,N_49060);
nor UO_4375 (O_4375,N_49633,N_49133);
and UO_4376 (O_4376,N_49218,N_49648);
nor UO_4377 (O_4377,N_49932,N_49694);
nor UO_4378 (O_4378,N_49364,N_49366);
nand UO_4379 (O_4379,N_49053,N_49673);
xor UO_4380 (O_4380,N_49915,N_49008);
nand UO_4381 (O_4381,N_49020,N_49298);
nand UO_4382 (O_4382,N_49177,N_49971);
and UO_4383 (O_4383,N_49205,N_49517);
nor UO_4384 (O_4384,N_49503,N_49473);
and UO_4385 (O_4385,N_49945,N_49435);
or UO_4386 (O_4386,N_49111,N_49726);
and UO_4387 (O_4387,N_49649,N_49742);
xnor UO_4388 (O_4388,N_49932,N_49385);
xor UO_4389 (O_4389,N_49388,N_49234);
and UO_4390 (O_4390,N_49636,N_49292);
nor UO_4391 (O_4391,N_49553,N_49346);
nor UO_4392 (O_4392,N_49004,N_49939);
or UO_4393 (O_4393,N_49507,N_49038);
or UO_4394 (O_4394,N_49831,N_49252);
or UO_4395 (O_4395,N_49189,N_49730);
xor UO_4396 (O_4396,N_49878,N_49024);
and UO_4397 (O_4397,N_49127,N_49461);
nand UO_4398 (O_4398,N_49964,N_49926);
nand UO_4399 (O_4399,N_49207,N_49795);
or UO_4400 (O_4400,N_49412,N_49603);
nand UO_4401 (O_4401,N_49032,N_49647);
xor UO_4402 (O_4402,N_49512,N_49618);
nor UO_4403 (O_4403,N_49795,N_49331);
or UO_4404 (O_4404,N_49725,N_49671);
or UO_4405 (O_4405,N_49446,N_49723);
or UO_4406 (O_4406,N_49375,N_49417);
and UO_4407 (O_4407,N_49378,N_49532);
nand UO_4408 (O_4408,N_49203,N_49423);
and UO_4409 (O_4409,N_49728,N_49850);
or UO_4410 (O_4410,N_49571,N_49278);
xor UO_4411 (O_4411,N_49716,N_49988);
nand UO_4412 (O_4412,N_49872,N_49826);
nand UO_4413 (O_4413,N_49725,N_49632);
xor UO_4414 (O_4414,N_49442,N_49607);
nand UO_4415 (O_4415,N_49347,N_49858);
nand UO_4416 (O_4416,N_49663,N_49015);
and UO_4417 (O_4417,N_49997,N_49678);
nand UO_4418 (O_4418,N_49730,N_49555);
nor UO_4419 (O_4419,N_49841,N_49656);
and UO_4420 (O_4420,N_49622,N_49848);
xnor UO_4421 (O_4421,N_49256,N_49727);
and UO_4422 (O_4422,N_49973,N_49067);
nand UO_4423 (O_4423,N_49956,N_49555);
nor UO_4424 (O_4424,N_49584,N_49924);
nor UO_4425 (O_4425,N_49808,N_49321);
nor UO_4426 (O_4426,N_49046,N_49669);
or UO_4427 (O_4427,N_49709,N_49406);
nor UO_4428 (O_4428,N_49703,N_49438);
or UO_4429 (O_4429,N_49248,N_49096);
nor UO_4430 (O_4430,N_49218,N_49146);
nor UO_4431 (O_4431,N_49719,N_49277);
or UO_4432 (O_4432,N_49149,N_49853);
nand UO_4433 (O_4433,N_49579,N_49418);
nor UO_4434 (O_4434,N_49269,N_49851);
and UO_4435 (O_4435,N_49592,N_49766);
and UO_4436 (O_4436,N_49074,N_49040);
or UO_4437 (O_4437,N_49334,N_49052);
nand UO_4438 (O_4438,N_49251,N_49254);
nor UO_4439 (O_4439,N_49496,N_49355);
or UO_4440 (O_4440,N_49851,N_49811);
and UO_4441 (O_4441,N_49753,N_49423);
xor UO_4442 (O_4442,N_49941,N_49783);
nand UO_4443 (O_4443,N_49349,N_49037);
nand UO_4444 (O_4444,N_49272,N_49501);
nor UO_4445 (O_4445,N_49621,N_49479);
and UO_4446 (O_4446,N_49511,N_49786);
and UO_4447 (O_4447,N_49390,N_49738);
nor UO_4448 (O_4448,N_49695,N_49488);
and UO_4449 (O_4449,N_49965,N_49217);
nor UO_4450 (O_4450,N_49399,N_49492);
or UO_4451 (O_4451,N_49086,N_49867);
xnor UO_4452 (O_4452,N_49191,N_49982);
xnor UO_4453 (O_4453,N_49820,N_49871);
or UO_4454 (O_4454,N_49223,N_49691);
nor UO_4455 (O_4455,N_49879,N_49043);
nor UO_4456 (O_4456,N_49828,N_49153);
nor UO_4457 (O_4457,N_49826,N_49967);
and UO_4458 (O_4458,N_49552,N_49817);
xor UO_4459 (O_4459,N_49957,N_49612);
or UO_4460 (O_4460,N_49129,N_49022);
xor UO_4461 (O_4461,N_49706,N_49437);
nand UO_4462 (O_4462,N_49466,N_49630);
nand UO_4463 (O_4463,N_49312,N_49561);
xor UO_4464 (O_4464,N_49902,N_49101);
or UO_4465 (O_4465,N_49269,N_49037);
nor UO_4466 (O_4466,N_49298,N_49584);
nor UO_4467 (O_4467,N_49672,N_49613);
nand UO_4468 (O_4468,N_49688,N_49099);
and UO_4469 (O_4469,N_49568,N_49282);
xnor UO_4470 (O_4470,N_49302,N_49854);
nand UO_4471 (O_4471,N_49037,N_49650);
nand UO_4472 (O_4472,N_49895,N_49730);
xor UO_4473 (O_4473,N_49197,N_49874);
nor UO_4474 (O_4474,N_49979,N_49824);
and UO_4475 (O_4475,N_49501,N_49507);
xor UO_4476 (O_4476,N_49599,N_49250);
and UO_4477 (O_4477,N_49531,N_49350);
xnor UO_4478 (O_4478,N_49477,N_49572);
or UO_4479 (O_4479,N_49287,N_49347);
xnor UO_4480 (O_4480,N_49356,N_49916);
xnor UO_4481 (O_4481,N_49256,N_49806);
and UO_4482 (O_4482,N_49132,N_49835);
nor UO_4483 (O_4483,N_49544,N_49228);
nand UO_4484 (O_4484,N_49221,N_49532);
xnor UO_4485 (O_4485,N_49868,N_49213);
and UO_4486 (O_4486,N_49133,N_49062);
and UO_4487 (O_4487,N_49780,N_49367);
and UO_4488 (O_4488,N_49807,N_49133);
or UO_4489 (O_4489,N_49053,N_49203);
nor UO_4490 (O_4490,N_49941,N_49908);
or UO_4491 (O_4491,N_49706,N_49647);
nand UO_4492 (O_4492,N_49429,N_49840);
nand UO_4493 (O_4493,N_49384,N_49154);
nor UO_4494 (O_4494,N_49943,N_49502);
xnor UO_4495 (O_4495,N_49697,N_49091);
nor UO_4496 (O_4496,N_49240,N_49925);
nand UO_4497 (O_4497,N_49859,N_49231);
and UO_4498 (O_4498,N_49595,N_49797);
xnor UO_4499 (O_4499,N_49515,N_49089);
nand UO_4500 (O_4500,N_49111,N_49069);
nor UO_4501 (O_4501,N_49549,N_49863);
and UO_4502 (O_4502,N_49544,N_49274);
or UO_4503 (O_4503,N_49449,N_49435);
or UO_4504 (O_4504,N_49792,N_49949);
xor UO_4505 (O_4505,N_49416,N_49774);
and UO_4506 (O_4506,N_49311,N_49121);
xor UO_4507 (O_4507,N_49503,N_49283);
and UO_4508 (O_4508,N_49821,N_49970);
nand UO_4509 (O_4509,N_49338,N_49264);
or UO_4510 (O_4510,N_49929,N_49028);
or UO_4511 (O_4511,N_49644,N_49636);
nand UO_4512 (O_4512,N_49194,N_49566);
and UO_4513 (O_4513,N_49695,N_49142);
or UO_4514 (O_4514,N_49973,N_49665);
nand UO_4515 (O_4515,N_49384,N_49762);
xnor UO_4516 (O_4516,N_49371,N_49398);
nor UO_4517 (O_4517,N_49678,N_49458);
xnor UO_4518 (O_4518,N_49270,N_49092);
nand UO_4519 (O_4519,N_49249,N_49561);
nor UO_4520 (O_4520,N_49544,N_49106);
and UO_4521 (O_4521,N_49944,N_49335);
and UO_4522 (O_4522,N_49209,N_49561);
nand UO_4523 (O_4523,N_49219,N_49165);
nand UO_4524 (O_4524,N_49900,N_49212);
and UO_4525 (O_4525,N_49645,N_49090);
nor UO_4526 (O_4526,N_49884,N_49861);
or UO_4527 (O_4527,N_49376,N_49497);
nand UO_4528 (O_4528,N_49293,N_49799);
xor UO_4529 (O_4529,N_49471,N_49540);
or UO_4530 (O_4530,N_49891,N_49054);
nor UO_4531 (O_4531,N_49964,N_49398);
or UO_4532 (O_4532,N_49927,N_49932);
and UO_4533 (O_4533,N_49482,N_49762);
nand UO_4534 (O_4534,N_49275,N_49627);
xor UO_4535 (O_4535,N_49171,N_49379);
or UO_4536 (O_4536,N_49323,N_49830);
nand UO_4537 (O_4537,N_49809,N_49253);
or UO_4538 (O_4538,N_49613,N_49385);
nand UO_4539 (O_4539,N_49884,N_49101);
and UO_4540 (O_4540,N_49020,N_49520);
nor UO_4541 (O_4541,N_49278,N_49695);
xor UO_4542 (O_4542,N_49741,N_49585);
nand UO_4543 (O_4543,N_49348,N_49009);
nor UO_4544 (O_4544,N_49186,N_49886);
xor UO_4545 (O_4545,N_49906,N_49148);
nand UO_4546 (O_4546,N_49808,N_49998);
nand UO_4547 (O_4547,N_49429,N_49936);
xnor UO_4548 (O_4548,N_49014,N_49602);
nor UO_4549 (O_4549,N_49132,N_49766);
and UO_4550 (O_4550,N_49588,N_49652);
nand UO_4551 (O_4551,N_49074,N_49188);
or UO_4552 (O_4552,N_49185,N_49561);
nor UO_4553 (O_4553,N_49774,N_49153);
nor UO_4554 (O_4554,N_49049,N_49130);
nand UO_4555 (O_4555,N_49659,N_49448);
xnor UO_4556 (O_4556,N_49265,N_49380);
and UO_4557 (O_4557,N_49833,N_49818);
xnor UO_4558 (O_4558,N_49765,N_49820);
nand UO_4559 (O_4559,N_49479,N_49160);
and UO_4560 (O_4560,N_49774,N_49545);
nor UO_4561 (O_4561,N_49378,N_49596);
nor UO_4562 (O_4562,N_49585,N_49565);
and UO_4563 (O_4563,N_49952,N_49138);
nor UO_4564 (O_4564,N_49212,N_49421);
nand UO_4565 (O_4565,N_49514,N_49667);
or UO_4566 (O_4566,N_49514,N_49018);
or UO_4567 (O_4567,N_49723,N_49876);
or UO_4568 (O_4568,N_49127,N_49129);
nor UO_4569 (O_4569,N_49183,N_49216);
or UO_4570 (O_4570,N_49611,N_49395);
or UO_4571 (O_4571,N_49995,N_49516);
or UO_4572 (O_4572,N_49507,N_49614);
or UO_4573 (O_4573,N_49934,N_49768);
nor UO_4574 (O_4574,N_49907,N_49626);
nand UO_4575 (O_4575,N_49378,N_49585);
nand UO_4576 (O_4576,N_49961,N_49875);
and UO_4577 (O_4577,N_49316,N_49197);
xor UO_4578 (O_4578,N_49710,N_49228);
nand UO_4579 (O_4579,N_49588,N_49527);
or UO_4580 (O_4580,N_49144,N_49637);
or UO_4581 (O_4581,N_49652,N_49409);
xnor UO_4582 (O_4582,N_49023,N_49408);
or UO_4583 (O_4583,N_49031,N_49049);
and UO_4584 (O_4584,N_49431,N_49366);
and UO_4585 (O_4585,N_49881,N_49572);
and UO_4586 (O_4586,N_49187,N_49974);
nor UO_4587 (O_4587,N_49192,N_49767);
and UO_4588 (O_4588,N_49105,N_49434);
and UO_4589 (O_4589,N_49777,N_49094);
xnor UO_4590 (O_4590,N_49131,N_49423);
xnor UO_4591 (O_4591,N_49237,N_49912);
nor UO_4592 (O_4592,N_49251,N_49444);
or UO_4593 (O_4593,N_49860,N_49752);
nor UO_4594 (O_4594,N_49834,N_49438);
nor UO_4595 (O_4595,N_49092,N_49219);
xnor UO_4596 (O_4596,N_49156,N_49811);
nand UO_4597 (O_4597,N_49765,N_49087);
and UO_4598 (O_4598,N_49897,N_49214);
and UO_4599 (O_4599,N_49236,N_49341);
nor UO_4600 (O_4600,N_49651,N_49075);
xnor UO_4601 (O_4601,N_49091,N_49194);
xor UO_4602 (O_4602,N_49271,N_49549);
and UO_4603 (O_4603,N_49284,N_49445);
xor UO_4604 (O_4604,N_49127,N_49439);
or UO_4605 (O_4605,N_49999,N_49246);
nand UO_4606 (O_4606,N_49723,N_49341);
xor UO_4607 (O_4607,N_49232,N_49218);
xor UO_4608 (O_4608,N_49922,N_49960);
or UO_4609 (O_4609,N_49952,N_49544);
nand UO_4610 (O_4610,N_49871,N_49385);
nor UO_4611 (O_4611,N_49577,N_49050);
nor UO_4612 (O_4612,N_49165,N_49930);
nand UO_4613 (O_4613,N_49196,N_49674);
and UO_4614 (O_4614,N_49254,N_49873);
or UO_4615 (O_4615,N_49644,N_49809);
xor UO_4616 (O_4616,N_49053,N_49762);
or UO_4617 (O_4617,N_49826,N_49926);
and UO_4618 (O_4618,N_49836,N_49720);
and UO_4619 (O_4619,N_49428,N_49989);
nand UO_4620 (O_4620,N_49513,N_49075);
nand UO_4621 (O_4621,N_49249,N_49110);
nand UO_4622 (O_4622,N_49162,N_49418);
xnor UO_4623 (O_4623,N_49558,N_49740);
and UO_4624 (O_4624,N_49272,N_49841);
xnor UO_4625 (O_4625,N_49635,N_49915);
or UO_4626 (O_4626,N_49797,N_49992);
nor UO_4627 (O_4627,N_49043,N_49241);
nand UO_4628 (O_4628,N_49637,N_49941);
nor UO_4629 (O_4629,N_49204,N_49382);
and UO_4630 (O_4630,N_49566,N_49313);
nor UO_4631 (O_4631,N_49850,N_49062);
xnor UO_4632 (O_4632,N_49411,N_49125);
nor UO_4633 (O_4633,N_49174,N_49010);
xor UO_4634 (O_4634,N_49463,N_49695);
or UO_4635 (O_4635,N_49234,N_49334);
nand UO_4636 (O_4636,N_49921,N_49653);
and UO_4637 (O_4637,N_49961,N_49941);
nor UO_4638 (O_4638,N_49901,N_49491);
and UO_4639 (O_4639,N_49539,N_49060);
nand UO_4640 (O_4640,N_49722,N_49665);
nor UO_4641 (O_4641,N_49984,N_49651);
or UO_4642 (O_4642,N_49464,N_49781);
nor UO_4643 (O_4643,N_49291,N_49025);
or UO_4644 (O_4644,N_49640,N_49914);
and UO_4645 (O_4645,N_49591,N_49979);
or UO_4646 (O_4646,N_49319,N_49827);
and UO_4647 (O_4647,N_49396,N_49327);
nor UO_4648 (O_4648,N_49769,N_49445);
and UO_4649 (O_4649,N_49195,N_49755);
and UO_4650 (O_4650,N_49474,N_49821);
or UO_4651 (O_4651,N_49518,N_49356);
and UO_4652 (O_4652,N_49078,N_49705);
or UO_4653 (O_4653,N_49098,N_49567);
xnor UO_4654 (O_4654,N_49967,N_49772);
xnor UO_4655 (O_4655,N_49872,N_49890);
nand UO_4656 (O_4656,N_49636,N_49041);
or UO_4657 (O_4657,N_49400,N_49962);
xor UO_4658 (O_4658,N_49995,N_49677);
nand UO_4659 (O_4659,N_49024,N_49501);
and UO_4660 (O_4660,N_49255,N_49405);
or UO_4661 (O_4661,N_49392,N_49213);
xnor UO_4662 (O_4662,N_49905,N_49674);
nor UO_4663 (O_4663,N_49770,N_49684);
nor UO_4664 (O_4664,N_49589,N_49883);
or UO_4665 (O_4665,N_49705,N_49446);
and UO_4666 (O_4666,N_49511,N_49400);
xnor UO_4667 (O_4667,N_49385,N_49435);
or UO_4668 (O_4668,N_49813,N_49854);
nor UO_4669 (O_4669,N_49048,N_49180);
xor UO_4670 (O_4670,N_49536,N_49862);
nor UO_4671 (O_4671,N_49482,N_49101);
nand UO_4672 (O_4672,N_49294,N_49905);
and UO_4673 (O_4673,N_49508,N_49777);
nor UO_4674 (O_4674,N_49014,N_49132);
nor UO_4675 (O_4675,N_49320,N_49420);
nand UO_4676 (O_4676,N_49070,N_49872);
xnor UO_4677 (O_4677,N_49086,N_49026);
or UO_4678 (O_4678,N_49264,N_49320);
or UO_4679 (O_4679,N_49056,N_49382);
or UO_4680 (O_4680,N_49642,N_49149);
or UO_4681 (O_4681,N_49809,N_49653);
or UO_4682 (O_4682,N_49354,N_49211);
and UO_4683 (O_4683,N_49734,N_49667);
nor UO_4684 (O_4684,N_49369,N_49319);
or UO_4685 (O_4685,N_49455,N_49930);
xor UO_4686 (O_4686,N_49089,N_49639);
and UO_4687 (O_4687,N_49726,N_49180);
and UO_4688 (O_4688,N_49448,N_49901);
nor UO_4689 (O_4689,N_49622,N_49942);
nor UO_4690 (O_4690,N_49900,N_49569);
or UO_4691 (O_4691,N_49756,N_49021);
nand UO_4692 (O_4692,N_49387,N_49526);
nor UO_4693 (O_4693,N_49747,N_49073);
xor UO_4694 (O_4694,N_49033,N_49084);
nor UO_4695 (O_4695,N_49374,N_49312);
or UO_4696 (O_4696,N_49503,N_49015);
xnor UO_4697 (O_4697,N_49897,N_49086);
or UO_4698 (O_4698,N_49600,N_49993);
nand UO_4699 (O_4699,N_49429,N_49272);
nor UO_4700 (O_4700,N_49012,N_49427);
and UO_4701 (O_4701,N_49938,N_49189);
nand UO_4702 (O_4702,N_49550,N_49935);
nand UO_4703 (O_4703,N_49494,N_49652);
and UO_4704 (O_4704,N_49317,N_49443);
nand UO_4705 (O_4705,N_49406,N_49873);
nor UO_4706 (O_4706,N_49436,N_49058);
or UO_4707 (O_4707,N_49799,N_49584);
xnor UO_4708 (O_4708,N_49680,N_49812);
nor UO_4709 (O_4709,N_49769,N_49429);
or UO_4710 (O_4710,N_49754,N_49550);
xor UO_4711 (O_4711,N_49485,N_49633);
and UO_4712 (O_4712,N_49096,N_49716);
or UO_4713 (O_4713,N_49927,N_49723);
or UO_4714 (O_4714,N_49954,N_49941);
nand UO_4715 (O_4715,N_49151,N_49276);
nor UO_4716 (O_4716,N_49159,N_49516);
nor UO_4717 (O_4717,N_49192,N_49440);
or UO_4718 (O_4718,N_49863,N_49442);
nand UO_4719 (O_4719,N_49579,N_49635);
or UO_4720 (O_4720,N_49960,N_49884);
and UO_4721 (O_4721,N_49247,N_49525);
and UO_4722 (O_4722,N_49026,N_49516);
xnor UO_4723 (O_4723,N_49597,N_49656);
nor UO_4724 (O_4724,N_49986,N_49793);
or UO_4725 (O_4725,N_49749,N_49859);
and UO_4726 (O_4726,N_49572,N_49860);
nor UO_4727 (O_4727,N_49381,N_49272);
xnor UO_4728 (O_4728,N_49677,N_49907);
nand UO_4729 (O_4729,N_49878,N_49268);
nor UO_4730 (O_4730,N_49702,N_49147);
nor UO_4731 (O_4731,N_49931,N_49665);
nor UO_4732 (O_4732,N_49684,N_49104);
nand UO_4733 (O_4733,N_49324,N_49913);
nor UO_4734 (O_4734,N_49419,N_49989);
nand UO_4735 (O_4735,N_49616,N_49939);
xor UO_4736 (O_4736,N_49595,N_49845);
or UO_4737 (O_4737,N_49655,N_49180);
xnor UO_4738 (O_4738,N_49575,N_49266);
or UO_4739 (O_4739,N_49333,N_49598);
nor UO_4740 (O_4740,N_49008,N_49682);
or UO_4741 (O_4741,N_49683,N_49413);
nand UO_4742 (O_4742,N_49025,N_49572);
or UO_4743 (O_4743,N_49655,N_49834);
and UO_4744 (O_4744,N_49871,N_49408);
nand UO_4745 (O_4745,N_49696,N_49933);
or UO_4746 (O_4746,N_49773,N_49114);
xnor UO_4747 (O_4747,N_49031,N_49489);
or UO_4748 (O_4748,N_49228,N_49208);
xnor UO_4749 (O_4749,N_49094,N_49048);
xnor UO_4750 (O_4750,N_49550,N_49993);
and UO_4751 (O_4751,N_49236,N_49748);
or UO_4752 (O_4752,N_49790,N_49401);
nand UO_4753 (O_4753,N_49400,N_49520);
or UO_4754 (O_4754,N_49767,N_49866);
nor UO_4755 (O_4755,N_49526,N_49422);
nor UO_4756 (O_4756,N_49392,N_49600);
nor UO_4757 (O_4757,N_49198,N_49127);
xor UO_4758 (O_4758,N_49201,N_49072);
xnor UO_4759 (O_4759,N_49715,N_49437);
and UO_4760 (O_4760,N_49624,N_49984);
nor UO_4761 (O_4761,N_49132,N_49175);
nand UO_4762 (O_4762,N_49759,N_49690);
nor UO_4763 (O_4763,N_49294,N_49324);
nor UO_4764 (O_4764,N_49428,N_49003);
xor UO_4765 (O_4765,N_49864,N_49765);
nand UO_4766 (O_4766,N_49650,N_49295);
nor UO_4767 (O_4767,N_49950,N_49602);
or UO_4768 (O_4768,N_49474,N_49057);
nand UO_4769 (O_4769,N_49938,N_49517);
or UO_4770 (O_4770,N_49394,N_49419);
xnor UO_4771 (O_4771,N_49174,N_49356);
xor UO_4772 (O_4772,N_49802,N_49976);
xor UO_4773 (O_4773,N_49423,N_49742);
xnor UO_4774 (O_4774,N_49156,N_49316);
or UO_4775 (O_4775,N_49734,N_49770);
nand UO_4776 (O_4776,N_49785,N_49594);
or UO_4777 (O_4777,N_49606,N_49533);
xnor UO_4778 (O_4778,N_49606,N_49302);
nand UO_4779 (O_4779,N_49741,N_49330);
nor UO_4780 (O_4780,N_49719,N_49734);
nor UO_4781 (O_4781,N_49503,N_49542);
nand UO_4782 (O_4782,N_49762,N_49310);
nor UO_4783 (O_4783,N_49370,N_49148);
or UO_4784 (O_4784,N_49325,N_49102);
and UO_4785 (O_4785,N_49665,N_49098);
and UO_4786 (O_4786,N_49267,N_49164);
nand UO_4787 (O_4787,N_49397,N_49916);
xor UO_4788 (O_4788,N_49387,N_49176);
nor UO_4789 (O_4789,N_49133,N_49575);
xnor UO_4790 (O_4790,N_49364,N_49569);
or UO_4791 (O_4791,N_49989,N_49167);
and UO_4792 (O_4792,N_49731,N_49049);
or UO_4793 (O_4793,N_49016,N_49065);
nor UO_4794 (O_4794,N_49219,N_49243);
nor UO_4795 (O_4795,N_49105,N_49728);
nor UO_4796 (O_4796,N_49894,N_49512);
and UO_4797 (O_4797,N_49342,N_49954);
xor UO_4798 (O_4798,N_49851,N_49711);
nor UO_4799 (O_4799,N_49008,N_49910);
nand UO_4800 (O_4800,N_49224,N_49178);
nor UO_4801 (O_4801,N_49931,N_49438);
nand UO_4802 (O_4802,N_49493,N_49153);
or UO_4803 (O_4803,N_49367,N_49155);
or UO_4804 (O_4804,N_49750,N_49080);
or UO_4805 (O_4805,N_49403,N_49915);
or UO_4806 (O_4806,N_49961,N_49590);
nor UO_4807 (O_4807,N_49037,N_49052);
and UO_4808 (O_4808,N_49076,N_49523);
nor UO_4809 (O_4809,N_49102,N_49113);
nand UO_4810 (O_4810,N_49801,N_49124);
nand UO_4811 (O_4811,N_49442,N_49244);
or UO_4812 (O_4812,N_49741,N_49009);
nand UO_4813 (O_4813,N_49386,N_49803);
or UO_4814 (O_4814,N_49120,N_49651);
nor UO_4815 (O_4815,N_49184,N_49969);
nand UO_4816 (O_4816,N_49222,N_49874);
nor UO_4817 (O_4817,N_49650,N_49095);
nor UO_4818 (O_4818,N_49466,N_49680);
or UO_4819 (O_4819,N_49937,N_49779);
and UO_4820 (O_4820,N_49339,N_49613);
or UO_4821 (O_4821,N_49653,N_49936);
nor UO_4822 (O_4822,N_49894,N_49543);
and UO_4823 (O_4823,N_49806,N_49092);
or UO_4824 (O_4824,N_49416,N_49054);
nor UO_4825 (O_4825,N_49820,N_49029);
and UO_4826 (O_4826,N_49411,N_49974);
xor UO_4827 (O_4827,N_49850,N_49252);
nand UO_4828 (O_4828,N_49455,N_49143);
and UO_4829 (O_4829,N_49594,N_49374);
nor UO_4830 (O_4830,N_49733,N_49127);
and UO_4831 (O_4831,N_49460,N_49592);
nor UO_4832 (O_4832,N_49943,N_49258);
nand UO_4833 (O_4833,N_49252,N_49890);
and UO_4834 (O_4834,N_49799,N_49681);
xor UO_4835 (O_4835,N_49832,N_49838);
nand UO_4836 (O_4836,N_49197,N_49176);
nand UO_4837 (O_4837,N_49129,N_49034);
and UO_4838 (O_4838,N_49437,N_49522);
and UO_4839 (O_4839,N_49163,N_49702);
xnor UO_4840 (O_4840,N_49542,N_49602);
xor UO_4841 (O_4841,N_49513,N_49135);
nor UO_4842 (O_4842,N_49588,N_49876);
xnor UO_4843 (O_4843,N_49050,N_49680);
nand UO_4844 (O_4844,N_49610,N_49721);
xor UO_4845 (O_4845,N_49832,N_49102);
and UO_4846 (O_4846,N_49037,N_49421);
xor UO_4847 (O_4847,N_49363,N_49157);
and UO_4848 (O_4848,N_49875,N_49541);
nor UO_4849 (O_4849,N_49471,N_49901);
and UO_4850 (O_4850,N_49004,N_49516);
nor UO_4851 (O_4851,N_49571,N_49499);
or UO_4852 (O_4852,N_49412,N_49411);
and UO_4853 (O_4853,N_49602,N_49783);
or UO_4854 (O_4854,N_49396,N_49128);
nand UO_4855 (O_4855,N_49420,N_49716);
nor UO_4856 (O_4856,N_49935,N_49128);
or UO_4857 (O_4857,N_49071,N_49864);
nand UO_4858 (O_4858,N_49334,N_49958);
nand UO_4859 (O_4859,N_49535,N_49098);
nor UO_4860 (O_4860,N_49639,N_49444);
xnor UO_4861 (O_4861,N_49682,N_49215);
and UO_4862 (O_4862,N_49412,N_49807);
nand UO_4863 (O_4863,N_49560,N_49379);
nor UO_4864 (O_4864,N_49745,N_49840);
xnor UO_4865 (O_4865,N_49950,N_49502);
nand UO_4866 (O_4866,N_49176,N_49663);
nor UO_4867 (O_4867,N_49682,N_49303);
or UO_4868 (O_4868,N_49210,N_49985);
or UO_4869 (O_4869,N_49544,N_49456);
and UO_4870 (O_4870,N_49566,N_49972);
or UO_4871 (O_4871,N_49178,N_49778);
and UO_4872 (O_4872,N_49359,N_49190);
xor UO_4873 (O_4873,N_49770,N_49946);
xor UO_4874 (O_4874,N_49950,N_49724);
nand UO_4875 (O_4875,N_49928,N_49348);
and UO_4876 (O_4876,N_49396,N_49669);
xnor UO_4877 (O_4877,N_49532,N_49609);
or UO_4878 (O_4878,N_49739,N_49878);
xnor UO_4879 (O_4879,N_49920,N_49555);
nand UO_4880 (O_4880,N_49829,N_49029);
and UO_4881 (O_4881,N_49981,N_49312);
nor UO_4882 (O_4882,N_49595,N_49429);
and UO_4883 (O_4883,N_49641,N_49010);
or UO_4884 (O_4884,N_49829,N_49010);
nor UO_4885 (O_4885,N_49239,N_49391);
and UO_4886 (O_4886,N_49577,N_49171);
nand UO_4887 (O_4887,N_49260,N_49676);
xor UO_4888 (O_4888,N_49277,N_49573);
or UO_4889 (O_4889,N_49053,N_49788);
nand UO_4890 (O_4890,N_49916,N_49130);
or UO_4891 (O_4891,N_49770,N_49397);
and UO_4892 (O_4892,N_49281,N_49170);
nor UO_4893 (O_4893,N_49296,N_49753);
or UO_4894 (O_4894,N_49862,N_49538);
nor UO_4895 (O_4895,N_49511,N_49293);
nor UO_4896 (O_4896,N_49295,N_49968);
xnor UO_4897 (O_4897,N_49520,N_49457);
nand UO_4898 (O_4898,N_49843,N_49403);
or UO_4899 (O_4899,N_49812,N_49290);
and UO_4900 (O_4900,N_49340,N_49947);
nor UO_4901 (O_4901,N_49291,N_49185);
or UO_4902 (O_4902,N_49744,N_49141);
nor UO_4903 (O_4903,N_49969,N_49350);
nor UO_4904 (O_4904,N_49895,N_49108);
nand UO_4905 (O_4905,N_49978,N_49755);
and UO_4906 (O_4906,N_49366,N_49690);
xor UO_4907 (O_4907,N_49559,N_49194);
xor UO_4908 (O_4908,N_49820,N_49825);
or UO_4909 (O_4909,N_49597,N_49000);
or UO_4910 (O_4910,N_49789,N_49047);
nand UO_4911 (O_4911,N_49671,N_49403);
and UO_4912 (O_4912,N_49385,N_49316);
xor UO_4913 (O_4913,N_49518,N_49367);
or UO_4914 (O_4914,N_49671,N_49778);
nand UO_4915 (O_4915,N_49826,N_49028);
nor UO_4916 (O_4916,N_49055,N_49703);
and UO_4917 (O_4917,N_49350,N_49040);
or UO_4918 (O_4918,N_49020,N_49905);
nor UO_4919 (O_4919,N_49075,N_49070);
nand UO_4920 (O_4920,N_49540,N_49230);
and UO_4921 (O_4921,N_49148,N_49085);
or UO_4922 (O_4922,N_49097,N_49345);
nand UO_4923 (O_4923,N_49300,N_49722);
nor UO_4924 (O_4924,N_49969,N_49608);
and UO_4925 (O_4925,N_49116,N_49569);
or UO_4926 (O_4926,N_49205,N_49248);
and UO_4927 (O_4927,N_49646,N_49776);
or UO_4928 (O_4928,N_49357,N_49983);
nor UO_4929 (O_4929,N_49452,N_49246);
xnor UO_4930 (O_4930,N_49374,N_49326);
nand UO_4931 (O_4931,N_49343,N_49317);
xnor UO_4932 (O_4932,N_49689,N_49482);
nor UO_4933 (O_4933,N_49906,N_49338);
nor UO_4934 (O_4934,N_49552,N_49947);
and UO_4935 (O_4935,N_49909,N_49919);
xor UO_4936 (O_4936,N_49551,N_49154);
xor UO_4937 (O_4937,N_49139,N_49842);
and UO_4938 (O_4938,N_49611,N_49510);
nor UO_4939 (O_4939,N_49809,N_49354);
nor UO_4940 (O_4940,N_49210,N_49196);
and UO_4941 (O_4941,N_49723,N_49290);
nor UO_4942 (O_4942,N_49947,N_49177);
nand UO_4943 (O_4943,N_49264,N_49041);
nand UO_4944 (O_4944,N_49783,N_49360);
xnor UO_4945 (O_4945,N_49069,N_49383);
and UO_4946 (O_4946,N_49102,N_49526);
xor UO_4947 (O_4947,N_49704,N_49652);
nand UO_4948 (O_4948,N_49249,N_49601);
or UO_4949 (O_4949,N_49554,N_49957);
and UO_4950 (O_4950,N_49306,N_49003);
and UO_4951 (O_4951,N_49859,N_49466);
nor UO_4952 (O_4952,N_49654,N_49636);
or UO_4953 (O_4953,N_49296,N_49463);
or UO_4954 (O_4954,N_49328,N_49402);
and UO_4955 (O_4955,N_49653,N_49935);
xor UO_4956 (O_4956,N_49296,N_49645);
and UO_4957 (O_4957,N_49304,N_49880);
nand UO_4958 (O_4958,N_49287,N_49672);
nor UO_4959 (O_4959,N_49965,N_49048);
xor UO_4960 (O_4960,N_49586,N_49483);
nand UO_4961 (O_4961,N_49289,N_49050);
or UO_4962 (O_4962,N_49341,N_49114);
nor UO_4963 (O_4963,N_49058,N_49748);
xnor UO_4964 (O_4964,N_49702,N_49317);
or UO_4965 (O_4965,N_49349,N_49135);
nand UO_4966 (O_4966,N_49390,N_49616);
and UO_4967 (O_4967,N_49733,N_49273);
and UO_4968 (O_4968,N_49768,N_49245);
xor UO_4969 (O_4969,N_49535,N_49234);
and UO_4970 (O_4970,N_49491,N_49924);
and UO_4971 (O_4971,N_49043,N_49806);
xor UO_4972 (O_4972,N_49490,N_49324);
nand UO_4973 (O_4973,N_49098,N_49350);
or UO_4974 (O_4974,N_49837,N_49903);
or UO_4975 (O_4975,N_49849,N_49043);
nand UO_4976 (O_4976,N_49794,N_49157);
or UO_4977 (O_4977,N_49068,N_49407);
or UO_4978 (O_4978,N_49555,N_49934);
nand UO_4979 (O_4979,N_49595,N_49642);
and UO_4980 (O_4980,N_49545,N_49366);
or UO_4981 (O_4981,N_49190,N_49014);
xor UO_4982 (O_4982,N_49221,N_49839);
and UO_4983 (O_4983,N_49479,N_49652);
or UO_4984 (O_4984,N_49833,N_49769);
nor UO_4985 (O_4985,N_49500,N_49601);
or UO_4986 (O_4986,N_49004,N_49726);
nor UO_4987 (O_4987,N_49875,N_49570);
or UO_4988 (O_4988,N_49997,N_49248);
or UO_4989 (O_4989,N_49431,N_49940);
or UO_4990 (O_4990,N_49128,N_49344);
nor UO_4991 (O_4991,N_49371,N_49901);
nand UO_4992 (O_4992,N_49296,N_49740);
and UO_4993 (O_4993,N_49293,N_49671);
or UO_4994 (O_4994,N_49747,N_49673);
or UO_4995 (O_4995,N_49104,N_49884);
nor UO_4996 (O_4996,N_49812,N_49625);
nand UO_4997 (O_4997,N_49667,N_49015);
nand UO_4998 (O_4998,N_49557,N_49177);
and UO_4999 (O_4999,N_49780,N_49590);
endmodule