module basic_500_3000_500_60_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_467,In_46);
or U1 (N_1,In_18,In_168);
or U2 (N_2,In_268,In_227);
nor U3 (N_3,In_371,In_197);
nor U4 (N_4,In_409,In_278);
or U5 (N_5,In_426,In_362);
nor U6 (N_6,In_211,In_58);
nand U7 (N_7,In_230,In_115);
nand U8 (N_8,In_482,In_298);
nor U9 (N_9,In_402,In_427);
nor U10 (N_10,In_484,In_249);
nand U11 (N_11,In_349,In_246);
nand U12 (N_12,In_290,In_345);
nand U13 (N_13,In_254,In_135);
nand U14 (N_14,In_55,In_233);
xor U15 (N_15,In_244,In_70);
and U16 (N_16,In_223,In_174);
nand U17 (N_17,In_54,In_151);
and U18 (N_18,In_203,In_65);
and U19 (N_19,In_215,In_108);
or U20 (N_20,In_36,In_71);
nor U21 (N_21,In_98,In_103);
nor U22 (N_22,In_380,In_430);
nor U23 (N_23,In_106,In_454);
or U24 (N_24,In_433,In_165);
or U25 (N_25,In_314,In_95);
nor U26 (N_26,In_339,In_253);
nor U27 (N_27,In_384,In_358);
or U28 (N_28,In_125,In_16);
nor U29 (N_29,In_325,In_446);
nor U30 (N_30,In_444,In_264);
nor U31 (N_31,In_60,In_202);
or U32 (N_32,In_256,In_379);
and U33 (N_33,In_69,In_159);
or U34 (N_34,In_225,In_76);
xor U35 (N_35,In_81,In_485);
or U36 (N_36,In_85,In_285);
nand U37 (N_37,In_294,In_99);
nor U38 (N_38,In_305,In_483);
xnor U39 (N_39,In_259,In_421);
and U40 (N_40,In_293,In_473);
and U41 (N_41,In_178,In_89);
xor U42 (N_42,In_82,In_496);
or U43 (N_43,In_251,In_329);
or U44 (N_44,In_411,In_383);
xor U45 (N_45,In_406,In_222);
nor U46 (N_46,In_318,In_456);
and U47 (N_47,In_149,In_338);
nor U48 (N_48,In_10,In_272);
nor U49 (N_49,In_389,In_42);
xnor U50 (N_50,N_33,In_27);
xor U51 (N_51,N_43,In_187);
xnor U52 (N_52,In_438,In_492);
and U53 (N_53,In_398,In_351);
and U54 (N_54,In_455,In_327);
nand U55 (N_55,In_226,In_330);
nor U56 (N_56,In_377,In_57);
nand U57 (N_57,In_333,In_397);
xnor U58 (N_58,In_413,In_453);
xor U59 (N_59,In_401,In_376);
and U60 (N_60,In_364,In_231);
xor U61 (N_61,N_0,In_143);
nand U62 (N_62,In_90,In_140);
or U63 (N_63,In_50,In_498);
nand U64 (N_64,In_241,In_214);
nand U65 (N_65,In_212,In_119);
nand U66 (N_66,N_12,In_417);
nor U67 (N_67,N_41,In_188);
nor U68 (N_68,In_0,In_334);
and U69 (N_69,In_367,In_445);
or U70 (N_70,In_410,In_229);
nor U71 (N_71,In_471,In_260);
or U72 (N_72,In_129,In_435);
nand U73 (N_73,In_171,In_127);
nand U74 (N_74,In_163,N_34);
and U75 (N_75,In_240,In_350);
nor U76 (N_76,In_20,In_283);
nand U77 (N_77,In_110,In_30);
nor U78 (N_78,In_133,In_64);
and U79 (N_79,In_354,In_469);
nor U80 (N_80,In_310,In_80);
xnor U81 (N_81,In_346,In_21);
nor U82 (N_82,In_247,In_180);
xnor U83 (N_83,In_437,In_109);
xor U84 (N_84,In_185,N_11);
nor U85 (N_85,In_478,In_400);
or U86 (N_86,In_287,In_275);
nor U87 (N_87,In_365,In_201);
nor U88 (N_88,In_276,In_196);
xor U89 (N_89,In_475,In_424);
nor U90 (N_90,N_16,In_447);
nor U91 (N_91,N_39,In_153);
nand U92 (N_92,In_8,In_48);
nor U93 (N_93,In_493,In_368);
and U94 (N_94,In_189,In_167);
nand U95 (N_95,In_279,In_175);
or U96 (N_96,In_378,In_432);
nor U97 (N_97,In_466,In_138);
or U98 (N_98,In_270,N_28);
xor U99 (N_99,In_176,In_45);
or U100 (N_100,In_407,In_479);
nor U101 (N_101,In_359,In_495);
nor U102 (N_102,In_184,In_232);
xor U103 (N_103,In_273,In_173);
nand U104 (N_104,In_146,In_78);
and U105 (N_105,In_489,N_57);
or U106 (N_106,In_117,In_261);
nand U107 (N_107,In_102,In_113);
nand U108 (N_108,In_487,In_343);
nand U109 (N_109,In_316,In_341);
nor U110 (N_110,N_74,In_24);
and U111 (N_111,In_136,In_199);
and U112 (N_112,In_418,In_392);
nor U113 (N_113,N_92,N_4);
nor U114 (N_114,N_98,In_262);
nand U115 (N_115,N_21,N_54);
nor U116 (N_116,In_147,N_42);
or U117 (N_117,In_28,In_114);
xor U118 (N_118,In_460,In_208);
nor U119 (N_119,In_66,In_356);
and U120 (N_120,In_281,In_62);
nor U121 (N_121,N_58,N_87);
nand U122 (N_122,In_289,In_37);
and U123 (N_123,In_11,In_152);
nor U124 (N_124,In_449,In_388);
xnor U125 (N_125,N_86,In_156);
xnor U126 (N_126,In_158,N_14);
nor U127 (N_127,In_292,N_67);
nor U128 (N_128,N_65,In_322);
xnor U129 (N_129,N_22,N_94);
or U130 (N_130,In_239,In_468);
nand U131 (N_131,In_150,In_266);
nor U132 (N_132,In_463,In_331);
nand U133 (N_133,In_32,In_205);
xnor U134 (N_134,N_13,In_404);
or U135 (N_135,In_284,In_451);
xor U136 (N_136,In_206,In_19);
xor U137 (N_137,In_224,In_181);
and U138 (N_138,N_10,In_480);
and U139 (N_139,In_179,In_481);
and U140 (N_140,In_172,In_461);
and U141 (N_141,N_46,In_161);
xor U142 (N_142,In_491,N_83);
or U143 (N_143,In_399,In_248);
xnor U144 (N_144,In_269,In_169);
nand U145 (N_145,In_123,In_235);
xnor U146 (N_146,In_182,In_228);
or U147 (N_147,In_450,In_302);
or U148 (N_148,In_43,In_440);
or U149 (N_149,In_155,In_100);
xor U150 (N_150,N_64,In_328);
nor U151 (N_151,N_37,In_470);
xnor U152 (N_152,In_47,In_191);
nor U153 (N_153,In_164,N_111);
and U154 (N_154,In_116,N_107);
or U155 (N_155,In_41,N_131);
xnor U156 (N_156,N_32,In_296);
or U157 (N_157,N_101,N_133);
and U158 (N_158,In_9,In_6);
nor U159 (N_159,In_216,N_7);
nor U160 (N_160,In_312,In_295);
nand U161 (N_161,In_44,In_309);
nand U162 (N_162,In_342,In_49);
xnor U163 (N_163,N_82,In_23);
nor U164 (N_164,N_6,In_112);
or U165 (N_165,N_124,In_29);
nor U166 (N_166,In_474,N_104);
xnor U167 (N_167,In_218,N_26);
or U168 (N_168,In_236,N_109);
xnor U169 (N_169,N_3,In_393);
nor U170 (N_170,In_434,In_59);
nand U171 (N_171,N_146,N_2);
xnor U172 (N_172,In_405,N_25);
or U173 (N_173,In_441,In_183);
and U174 (N_174,N_113,In_67);
xnor U175 (N_175,N_19,In_361);
nand U176 (N_176,In_458,N_1);
nor U177 (N_177,In_360,In_38);
nand U178 (N_178,N_102,N_72);
nor U179 (N_179,In_303,In_439);
nand U180 (N_180,In_395,In_87);
or U181 (N_181,In_263,In_154);
and U182 (N_182,N_126,N_15);
nand U183 (N_183,In_210,N_29);
nor U184 (N_184,In_15,N_8);
nand U185 (N_185,N_45,In_436);
nand U186 (N_186,N_53,In_301);
or U187 (N_187,N_52,N_9);
and U188 (N_188,In_490,N_123);
nand U189 (N_189,N_59,N_80);
or U190 (N_190,In_237,In_375);
xnor U191 (N_191,In_477,In_258);
nand U192 (N_192,N_47,N_103);
or U193 (N_193,N_75,N_30);
xnor U194 (N_194,In_332,In_372);
or U195 (N_195,In_355,In_93);
and U196 (N_196,In_282,N_129);
nor U197 (N_197,In_14,In_363);
xor U198 (N_198,In_190,N_130);
or U199 (N_199,In_141,In_22);
or U200 (N_200,In_428,N_157);
nand U201 (N_201,N_68,N_17);
xor U202 (N_202,N_145,N_181);
nand U203 (N_203,N_55,In_51);
nor U204 (N_204,In_326,In_366);
or U205 (N_205,In_142,In_344);
nor U206 (N_206,In_170,In_234);
nand U207 (N_207,N_132,In_61);
nor U208 (N_208,N_118,In_52);
nor U209 (N_209,In_442,N_24);
nand U210 (N_210,In_34,In_2);
or U211 (N_211,In_308,In_1);
xor U212 (N_212,N_66,In_373);
nand U213 (N_213,In_452,N_106);
nand U214 (N_214,In_72,In_12);
and U215 (N_215,In_17,N_151);
and U216 (N_216,In_194,N_140);
nand U217 (N_217,In_465,In_416);
and U218 (N_218,N_27,In_391);
nor U219 (N_219,N_90,N_147);
nor U220 (N_220,In_297,In_369);
xor U221 (N_221,In_3,In_299);
or U222 (N_222,N_172,In_157);
nor U223 (N_223,In_288,In_131);
xor U224 (N_224,In_120,N_71);
nand U225 (N_225,In_457,In_101);
xor U226 (N_226,N_164,N_125);
or U227 (N_227,N_186,In_243);
xor U228 (N_228,N_179,In_403);
xor U229 (N_229,In_464,In_300);
nor U230 (N_230,In_74,In_84);
nor U231 (N_231,In_267,In_423);
xor U232 (N_232,In_381,In_387);
nor U233 (N_233,N_49,In_459);
or U234 (N_234,In_385,In_193);
xnor U235 (N_235,In_472,In_238);
xor U236 (N_236,In_271,N_170);
xnor U237 (N_237,In_40,In_104);
and U238 (N_238,N_38,In_422);
nand U239 (N_239,In_35,In_166);
xnor U240 (N_240,In_386,In_75);
nand U241 (N_241,N_160,N_141);
and U242 (N_242,N_128,N_73);
and U243 (N_243,N_194,In_192);
nor U244 (N_244,In_139,N_117);
xor U245 (N_245,N_110,In_353);
xnor U246 (N_246,N_174,In_494);
nand U247 (N_247,N_173,N_79);
and U248 (N_248,N_163,In_111);
xnor U249 (N_249,N_198,N_171);
nor U250 (N_250,N_142,In_77);
xor U251 (N_251,N_50,N_161);
or U252 (N_252,N_76,N_234);
xor U253 (N_253,In_390,In_336);
xor U254 (N_254,N_200,N_216);
nor U255 (N_255,N_223,N_96);
nor U256 (N_256,In_221,N_213);
nor U257 (N_257,N_138,In_476);
nand U258 (N_258,In_408,N_215);
nand U259 (N_259,In_242,N_247);
nor U260 (N_260,In_220,N_120);
nand U261 (N_261,In_317,N_97);
nor U262 (N_262,N_116,In_219);
xor U263 (N_263,In_306,In_107);
and U264 (N_264,N_187,N_212);
and U265 (N_265,In_352,N_167);
nor U266 (N_266,In_429,In_39);
or U267 (N_267,N_180,N_226);
xor U268 (N_268,N_136,In_337);
or U269 (N_269,N_23,N_122);
nor U270 (N_270,In_83,In_448);
xnor U271 (N_271,In_324,In_134);
nor U272 (N_272,N_139,N_183);
nand U273 (N_273,In_394,N_100);
and U274 (N_274,N_228,N_168);
and U275 (N_275,N_78,In_96);
nand U276 (N_276,In_488,N_189);
nor U277 (N_277,N_222,N_202);
or U278 (N_278,In_320,In_5);
xnor U279 (N_279,N_177,N_56);
nor U280 (N_280,N_203,In_497);
or U281 (N_281,In_4,In_291);
nand U282 (N_282,In_86,N_91);
nand U283 (N_283,In_304,N_81);
or U284 (N_284,In_431,In_124);
xnor U285 (N_285,N_235,In_132);
xnor U286 (N_286,In_412,In_53);
xnor U287 (N_287,N_143,N_159);
nand U288 (N_288,In_414,In_91);
xnor U289 (N_289,In_121,In_186);
nand U290 (N_290,N_89,In_321);
nor U291 (N_291,In_462,N_63);
and U292 (N_292,In_177,N_84);
nor U293 (N_293,N_238,In_209);
nand U294 (N_294,In_213,In_348);
nor U295 (N_295,N_150,N_184);
nor U296 (N_296,N_119,In_323);
xnor U297 (N_297,In_122,In_56);
or U298 (N_298,In_347,N_229);
or U299 (N_299,N_208,N_246);
nor U300 (N_300,N_299,In_319);
or U301 (N_301,In_374,N_219);
or U302 (N_302,N_288,N_191);
xnor U303 (N_303,N_236,N_210);
nand U304 (N_304,N_273,In_33);
nor U305 (N_305,In_137,N_61);
or U306 (N_306,N_99,In_357);
and U307 (N_307,N_195,N_35);
or U308 (N_308,N_220,N_248);
nor U309 (N_309,N_295,N_62);
nand U310 (N_310,N_232,N_256);
and U311 (N_311,N_190,N_214);
xnor U312 (N_312,In_92,N_257);
or U313 (N_313,In_396,N_217);
and U314 (N_314,In_257,N_281);
xnor U315 (N_315,In_130,In_144);
nor U316 (N_316,N_60,In_68);
nand U317 (N_317,N_261,In_420);
xnor U318 (N_318,N_70,N_114);
nand U319 (N_319,N_249,N_40);
xor U320 (N_320,N_206,N_196);
and U321 (N_321,N_268,N_277);
xnor U322 (N_322,N_199,N_121);
nor U323 (N_323,N_127,N_95);
nor U324 (N_324,N_278,N_108);
xor U325 (N_325,N_156,N_294);
nor U326 (N_326,N_204,N_243);
xor U327 (N_327,In_198,In_13);
nor U328 (N_328,In_26,N_239);
or U329 (N_329,N_5,N_272);
or U330 (N_330,In_145,N_251);
nand U331 (N_331,N_263,N_225);
nand U332 (N_332,In_88,In_97);
xnor U333 (N_333,In_162,N_169);
nand U334 (N_334,N_152,N_276);
and U335 (N_335,N_205,N_296);
nand U336 (N_336,N_105,In_160);
and U337 (N_337,N_292,N_193);
xor U338 (N_338,N_258,N_197);
and U339 (N_339,N_218,In_105);
xor U340 (N_340,N_44,N_137);
xnor U341 (N_341,N_224,N_290);
and U342 (N_342,In_217,N_282);
or U343 (N_343,N_69,N_231);
and U344 (N_344,N_245,In_382);
xnor U345 (N_345,In_207,N_221);
xnor U346 (N_346,In_252,N_227);
and U347 (N_347,In_200,N_176);
and U348 (N_348,N_253,In_148);
nor U349 (N_349,In_94,In_204);
and U350 (N_350,N_343,In_79);
xor U351 (N_351,N_300,N_303);
nor U352 (N_352,N_148,N_155);
or U353 (N_353,N_338,N_211);
nor U354 (N_354,N_201,In_73);
nand U355 (N_355,N_149,In_274);
xnor U356 (N_356,N_285,N_349);
and U357 (N_357,N_88,N_339);
nand U358 (N_358,N_342,In_335);
or U359 (N_359,N_310,In_443);
or U360 (N_360,In_250,N_18);
nand U361 (N_361,N_334,N_271);
xnor U362 (N_362,N_270,N_316);
and U363 (N_363,N_77,N_269);
or U364 (N_364,N_240,N_185);
nor U365 (N_365,N_250,N_298);
and U366 (N_366,N_301,N_237);
nor U367 (N_367,N_337,N_207);
and U368 (N_368,N_158,N_329);
nand U369 (N_369,N_259,N_304);
and U370 (N_370,N_115,N_244);
and U371 (N_371,N_154,In_315);
and U372 (N_372,N_311,N_209);
nor U373 (N_373,N_188,In_311);
or U374 (N_374,N_112,In_286);
and U375 (N_375,N_335,N_284);
and U376 (N_376,N_330,N_312);
nor U377 (N_377,N_51,N_320);
or U378 (N_378,N_346,N_252);
or U379 (N_379,N_315,N_340);
nand U380 (N_380,N_241,In_340);
xnor U381 (N_381,N_242,N_192);
or U382 (N_382,N_318,N_233);
and U383 (N_383,N_280,N_323);
or U384 (N_384,N_289,N_230);
nand U385 (N_385,N_260,N_341);
and U386 (N_386,N_336,N_321);
or U387 (N_387,N_331,N_165);
nand U388 (N_388,N_264,N_162);
or U389 (N_389,N_178,N_166);
or U390 (N_390,N_347,N_314);
and U391 (N_391,N_326,N_283);
or U392 (N_392,N_266,In_265);
xnor U393 (N_393,N_287,N_291);
xnor U394 (N_394,N_274,N_307);
and U395 (N_395,N_313,N_348);
nand U396 (N_396,In_7,N_267);
and U397 (N_397,N_322,In_255);
nand U398 (N_398,N_345,N_262);
xor U399 (N_399,N_93,In_415);
nor U400 (N_400,In_499,N_395);
or U401 (N_401,In_486,N_293);
nand U402 (N_402,N_352,N_355);
xnor U403 (N_403,N_286,N_332);
or U404 (N_404,N_302,In_31);
and U405 (N_405,N_305,N_350);
nand U406 (N_406,N_358,N_297);
nor U407 (N_407,N_374,N_375);
nor U408 (N_408,N_344,In_63);
and U409 (N_409,In_280,In_245);
xor U410 (N_410,N_381,In_313);
nand U411 (N_411,N_380,N_365);
nor U412 (N_412,N_353,N_319);
or U413 (N_413,N_379,N_328);
or U414 (N_414,N_324,N_327);
nor U415 (N_415,N_372,N_386);
nor U416 (N_416,N_254,N_309);
nor U417 (N_417,N_399,N_134);
nand U418 (N_418,N_370,N_388);
nor U419 (N_419,N_351,In_277);
nand U420 (N_420,N_362,N_396);
nand U421 (N_421,N_275,N_391);
and U422 (N_422,N_363,N_361);
xnor U423 (N_423,N_36,N_398);
nand U424 (N_424,N_367,In_307);
or U425 (N_425,In_25,N_85);
nor U426 (N_426,N_333,N_317);
xor U427 (N_427,N_359,N_382);
xnor U428 (N_428,N_376,N_366);
or U429 (N_429,N_378,N_389);
or U430 (N_430,N_279,N_306);
or U431 (N_431,N_387,N_182);
or U432 (N_432,N_357,N_255);
and U433 (N_433,N_356,N_371);
or U434 (N_434,N_392,N_265);
or U435 (N_435,N_377,N_369);
or U436 (N_436,In_195,N_153);
nor U437 (N_437,N_325,N_394);
nand U438 (N_438,N_393,N_397);
nand U439 (N_439,N_373,N_384);
and U440 (N_440,In_118,N_383);
xnor U441 (N_441,N_360,N_364);
nand U442 (N_442,N_175,N_20);
nor U443 (N_443,N_354,In_419);
nor U444 (N_444,N_390,In_128);
or U445 (N_445,N_308,N_31);
nor U446 (N_446,N_368,N_135);
and U447 (N_447,In_425,N_48);
or U448 (N_448,N_385,In_370);
and U449 (N_449,In_126,N_144);
nor U450 (N_450,N_419,N_402);
xnor U451 (N_451,N_449,N_437);
nor U452 (N_452,N_431,N_416);
nand U453 (N_453,N_426,N_424);
nand U454 (N_454,N_429,N_432);
or U455 (N_455,N_444,N_406);
xnor U456 (N_456,N_407,N_410);
xor U457 (N_457,N_411,N_448);
nand U458 (N_458,N_433,N_420);
nand U459 (N_459,N_403,N_442);
and U460 (N_460,N_436,N_417);
and U461 (N_461,N_408,N_443);
nor U462 (N_462,N_434,N_441);
nand U463 (N_463,N_421,N_405);
or U464 (N_464,N_423,N_414);
and U465 (N_465,N_425,N_447);
or U466 (N_466,N_422,N_439);
nor U467 (N_467,N_401,N_446);
nor U468 (N_468,N_435,N_412);
nor U469 (N_469,N_400,N_428);
nand U470 (N_470,N_415,N_438);
nor U471 (N_471,N_404,N_418);
and U472 (N_472,N_440,N_427);
and U473 (N_473,N_430,N_445);
and U474 (N_474,N_413,N_409);
nor U475 (N_475,N_447,N_423);
nand U476 (N_476,N_430,N_443);
and U477 (N_477,N_445,N_413);
nor U478 (N_478,N_444,N_430);
nand U479 (N_479,N_412,N_420);
nand U480 (N_480,N_442,N_414);
or U481 (N_481,N_419,N_429);
xnor U482 (N_482,N_434,N_410);
and U483 (N_483,N_413,N_414);
nand U484 (N_484,N_423,N_420);
xnor U485 (N_485,N_449,N_439);
nand U486 (N_486,N_429,N_408);
or U487 (N_487,N_434,N_447);
and U488 (N_488,N_448,N_410);
or U489 (N_489,N_407,N_420);
xnor U490 (N_490,N_432,N_437);
nand U491 (N_491,N_404,N_439);
nand U492 (N_492,N_413,N_402);
nand U493 (N_493,N_440,N_437);
xor U494 (N_494,N_402,N_448);
nor U495 (N_495,N_448,N_404);
or U496 (N_496,N_422,N_416);
or U497 (N_497,N_408,N_445);
nand U498 (N_498,N_424,N_411);
xnor U499 (N_499,N_444,N_413);
nand U500 (N_500,N_458,N_492);
and U501 (N_501,N_491,N_457);
or U502 (N_502,N_464,N_483);
and U503 (N_503,N_471,N_467);
xor U504 (N_504,N_473,N_460);
and U505 (N_505,N_454,N_486);
nand U506 (N_506,N_462,N_477);
or U507 (N_507,N_498,N_488);
and U508 (N_508,N_485,N_472);
nand U509 (N_509,N_499,N_461);
and U510 (N_510,N_465,N_455);
and U511 (N_511,N_468,N_475);
and U512 (N_512,N_453,N_451);
xnor U513 (N_513,N_470,N_495);
xor U514 (N_514,N_489,N_493);
nor U515 (N_515,N_466,N_494);
and U516 (N_516,N_496,N_481);
or U517 (N_517,N_490,N_484);
nand U518 (N_518,N_450,N_469);
and U519 (N_519,N_487,N_463);
or U520 (N_520,N_474,N_452);
or U521 (N_521,N_497,N_476);
or U522 (N_522,N_480,N_482);
and U523 (N_523,N_459,N_456);
nand U524 (N_524,N_478,N_479);
nand U525 (N_525,N_458,N_450);
nor U526 (N_526,N_487,N_499);
xor U527 (N_527,N_458,N_481);
nand U528 (N_528,N_455,N_491);
nand U529 (N_529,N_495,N_491);
xnor U530 (N_530,N_454,N_460);
and U531 (N_531,N_450,N_480);
or U532 (N_532,N_483,N_457);
and U533 (N_533,N_494,N_482);
xor U534 (N_534,N_494,N_495);
or U535 (N_535,N_464,N_451);
nor U536 (N_536,N_476,N_474);
and U537 (N_537,N_489,N_476);
nor U538 (N_538,N_464,N_472);
and U539 (N_539,N_464,N_498);
and U540 (N_540,N_494,N_453);
xnor U541 (N_541,N_460,N_472);
or U542 (N_542,N_482,N_497);
nand U543 (N_543,N_453,N_450);
nor U544 (N_544,N_495,N_498);
and U545 (N_545,N_455,N_471);
nand U546 (N_546,N_450,N_491);
and U547 (N_547,N_498,N_457);
nor U548 (N_548,N_471,N_498);
and U549 (N_549,N_465,N_457);
nor U550 (N_550,N_515,N_532);
nor U551 (N_551,N_524,N_518);
nand U552 (N_552,N_533,N_508);
or U553 (N_553,N_537,N_547);
or U554 (N_554,N_522,N_531);
xnor U555 (N_555,N_542,N_516);
xor U556 (N_556,N_513,N_506);
and U557 (N_557,N_528,N_535);
and U558 (N_558,N_534,N_526);
and U559 (N_559,N_539,N_507);
nor U560 (N_560,N_503,N_511);
or U561 (N_561,N_525,N_521);
nand U562 (N_562,N_500,N_504);
nand U563 (N_563,N_548,N_546);
nor U564 (N_564,N_529,N_519);
nor U565 (N_565,N_505,N_514);
nor U566 (N_566,N_538,N_543);
nor U567 (N_567,N_540,N_527);
xor U568 (N_568,N_523,N_501);
and U569 (N_569,N_545,N_541);
nand U570 (N_570,N_509,N_549);
nor U571 (N_571,N_544,N_536);
nor U572 (N_572,N_502,N_517);
nor U573 (N_573,N_512,N_510);
xor U574 (N_574,N_520,N_530);
and U575 (N_575,N_511,N_537);
and U576 (N_576,N_529,N_501);
or U577 (N_577,N_508,N_524);
and U578 (N_578,N_528,N_503);
or U579 (N_579,N_505,N_500);
xor U580 (N_580,N_535,N_529);
and U581 (N_581,N_545,N_509);
nand U582 (N_582,N_506,N_538);
xor U583 (N_583,N_504,N_541);
xnor U584 (N_584,N_533,N_500);
xor U585 (N_585,N_500,N_518);
nor U586 (N_586,N_545,N_523);
xnor U587 (N_587,N_540,N_547);
and U588 (N_588,N_522,N_513);
nor U589 (N_589,N_527,N_535);
nor U590 (N_590,N_537,N_505);
or U591 (N_591,N_543,N_542);
or U592 (N_592,N_506,N_518);
xnor U593 (N_593,N_518,N_505);
nor U594 (N_594,N_500,N_541);
xor U595 (N_595,N_507,N_501);
and U596 (N_596,N_514,N_502);
xnor U597 (N_597,N_544,N_548);
nor U598 (N_598,N_506,N_526);
xor U599 (N_599,N_533,N_544);
or U600 (N_600,N_590,N_572);
nor U601 (N_601,N_558,N_582);
and U602 (N_602,N_596,N_592);
and U603 (N_603,N_593,N_570);
and U604 (N_604,N_561,N_556);
and U605 (N_605,N_599,N_575);
and U606 (N_606,N_580,N_559);
nor U607 (N_607,N_579,N_567);
xnor U608 (N_608,N_568,N_552);
nor U609 (N_609,N_589,N_585);
and U610 (N_610,N_550,N_574);
and U611 (N_611,N_553,N_562);
or U612 (N_612,N_598,N_577);
xor U613 (N_613,N_566,N_578);
or U614 (N_614,N_594,N_595);
nor U615 (N_615,N_555,N_581);
xor U616 (N_616,N_573,N_565);
xor U617 (N_617,N_587,N_564);
nor U618 (N_618,N_588,N_551);
or U619 (N_619,N_597,N_576);
nand U620 (N_620,N_554,N_571);
and U621 (N_621,N_563,N_569);
xnor U622 (N_622,N_583,N_560);
nand U623 (N_623,N_557,N_591);
xnor U624 (N_624,N_586,N_584);
xor U625 (N_625,N_556,N_552);
and U626 (N_626,N_582,N_597);
xnor U627 (N_627,N_570,N_565);
and U628 (N_628,N_582,N_591);
and U629 (N_629,N_558,N_557);
nor U630 (N_630,N_570,N_566);
or U631 (N_631,N_563,N_559);
nand U632 (N_632,N_572,N_565);
nor U633 (N_633,N_575,N_568);
or U634 (N_634,N_568,N_586);
nor U635 (N_635,N_566,N_583);
nand U636 (N_636,N_587,N_586);
xor U637 (N_637,N_579,N_583);
xnor U638 (N_638,N_563,N_554);
and U639 (N_639,N_569,N_574);
nand U640 (N_640,N_597,N_566);
nand U641 (N_641,N_577,N_555);
or U642 (N_642,N_590,N_565);
xor U643 (N_643,N_557,N_575);
or U644 (N_644,N_584,N_590);
nand U645 (N_645,N_575,N_588);
nor U646 (N_646,N_590,N_579);
or U647 (N_647,N_591,N_555);
nand U648 (N_648,N_563,N_594);
nor U649 (N_649,N_576,N_579);
or U650 (N_650,N_603,N_614);
nand U651 (N_651,N_637,N_630);
nand U652 (N_652,N_600,N_621);
xor U653 (N_653,N_606,N_647);
nor U654 (N_654,N_645,N_623);
and U655 (N_655,N_602,N_615);
and U656 (N_656,N_636,N_611);
and U657 (N_657,N_638,N_620);
nor U658 (N_658,N_622,N_642);
nor U659 (N_659,N_634,N_607);
and U660 (N_660,N_619,N_627);
xor U661 (N_661,N_646,N_643);
xnor U662 (N_662,N_628,N_639);
and U663 (N_663,N_635,N_604);
or U664 (N_664,N_631,N_616);
and U665 (N_665,N_626,N_632);
and U666 (N_666,N_601,N_625);
nand U667 (N_667,N_617,N_612);
nand U668 (N_668,N_648,N_609);
or U669 (N_669,N_610,N_629);
or U670 (N_670,N_640,N_644);
nor U671 (N_671,N_641,N_608);
and U672 (N_672,N_624,N_649);
nor U673 (N_673,N_605,N_613);
and U674 (N_674,N_618,N_633);
nor U675 (N_675,N_615,N_649);
or U676 (N_676,N_631,N_622);
nor U677 (N_677,N_620,N_600);
or U678 (N_678,N_607,N_647);
nand U679 (N_679,N_603,N_622);
and U680 (N_680,N_614,N_647);
nor U681 (N_681,N_632,N_610);
or U682 (N_682,N_623,N_617);
and U683 (N_683,N_600,N_602);
nor U684 (N_684,N_621,N_622);
xor U685 (N_685,N_610,N_624);
nor U686 (N_686,N_626,N_614);
xor U687 (N_687,N_627,N_617);
nand U688 (N_688,N_643,N_616);
and U689 (N_689,N_640,N_645);
xnor U690 (N_690,N_639,N_623);
nor U691 (N_691,N_644,N_603);
or U692 (N_692,N_635,N_611);
or U693 (N_693,N_642,N_617);
and U694 (N_694,N_632,N_605);
xnor U695 (N_695,N_644,N_632);
and U696 (N_696,N_631,N_623);
nand U697 (N_697,N_629,N_643);
or U698 (N_698,N_600,N_603);
and U699 (N_699,N_649,N_637);
nor U700 (N_700,N_675,N_653);
or U701 (N_701,N_684,N_664);
or U702 (N_702,N_656,N_696);
nor U703 (N_703,N_665,N_682);
nand U704 (N_704,N_662,N_667);
and U705 (N_705,N_660,N_690);
nand U706 (N_706,N_657,N_670);
and U707 (N_707,N_677,N_680);
nand U708 (N_708,N_683,N_699);
nand U709 (N_709,N_695,N_658);
nand U710 (N_710,N_651,N_687);
xnor U711 (N_711,N_688,N_697);
or U712 (N_712,N_693,N_654);
nand U713 (N_713,N_650,N_698);
xor U714 (N_714,N_661,N_659);
xnor U715 (N_715,N_686,N_694);
nand U716 (N_716,N_679,N_666);
nand U717 (N_717,N_685,N_671);
or U718 (N_718,N_681,N_678);
and U719 (N_719,N_691,N_669);
and U720 (N_720,N_663,N_674);
and U721 (N_721,N_676,N_652);
nor U722 (N_722,N_668,N_689);
or U723 (N_723,N_673,N_672);
or U724 (N_724,N_655,N_692);
or U725 (N_725,N_673,N_663);
or U726 (N_726,N_679,N_652);
and U727 (N_727,N_662,N_665);
nand U728 (N_728,N_663,N_651);
xnor U729 (N_729,N_670,N_688);
or U730 (N_730,N_672,N_697);
nand U731 (N_731,N_659,N_658);
nand U732 (N_732,N_692,N_695);
xor U733 (N_733,N_659,N_696);
nand U734 (N_734,N_674,N_666);
or U735 (N_735,N_687,N_660);
xnor U736 (N_736,N_683,N_655);
xnor U737 (N_737,N_661,N_696);
xnor U738 (N_738,N_662,N_672);
nor U739 (N_739,N_688,N_662);
nor U740 (N_740,N_682,N_668);
and U741 (N_741,N_672,N_689);
nand U742 (N_742,N_690,N_685);
nand U743 (N_743,N_696,N_679);
nand U744 (N_744,N_651,N_654);
or U745 (N_745,N_680,N_699);
xor U746 (N_746,N_650,N_661);
xnor U747 (N_747,N_686,N_691);
or U748 (N_748,N_680,N_656);
or U749 (N_749,N_664,N_679);
and U750 (N_750,N_702,N_748);
and U751 (N_751,N_734,N_724);
xor U752 (N_752,N_736,N_729);
xnor U753 (N_753,N_722,N_708);
xor U754 (N_754,N_705,N_726);
and U755 (N_755,N_712,N_747);
nand U756 (N_756,N_711,N_707);
nor U757 (N_757,N_703,N_740);
nand U758 (N_758,N_706,N_719);
or U759 (N_759,N_717,N_723);
nor U760 (N_760,N_700,N_728);
nand U761 (N_761,N_720,N_738);
nand U762 (N_762,N_730,N_721);
nor U763 (N_763,N_727,N_716);
or U764 (N_764,N_732,N_709);
xor U765 (N_765,N_746,N_743);
or U766 (N_766,N_739,N_701);
and U767 (N_767,N_735,N_749);
and U768 (N_768,N_744,N_737);
or U769 (N_769,N_741,N_742);
nand U770 (N_770,N_710,N_725);
or U771 (N_771,N_715,N_713);
and U772 (N_772,N_704,N_718);
nor U773 (N_773,N_745,N_714);
xnor U774 (N_774,N_733,N_731);
or U775 (N_775,N_709,N_746);
xor U776 (N_776,N_725,N_740);
xnor U777 (N_777,N_738,N_725);
nand U778 (N_778,N_718,N_724);
xnor U779 (N_779,N_747,N_736);
xor U780 (N_780,N_733,N_728);
nor U781 (N_781,N_728,N_724);
xnor U782 (N_782,N_749,N_747);
and U783 (N_783,N_715,N_709);
nand U784 (N_784,N_730,N_709);
nand U785 (N_785,N_736,N_741);
or U786 (N_786,N_729,N_733);
and U787 (N_787,N_715,N_745);
nor U788 (N_788,N_720,N_731);
nand U789 (N_789,N_749,N_714);
xor U790 (N_790,N_719,N_713);
nor U791 (N_791,N_720,N_705);
and U792 (N_792,N_734,N_715);
nand U793 (N_793,N_747,N_730);
and U794 (N_794,N_735,N_741);
and U795 (N_795,N_743,N_740);
or U796 (N_796,N_730,N_716);
nand U797 (N_797,N_704,N_702);
nand U798 (N_798,N_720,N_718);
or U799 (N_799,N_734,N_701);
or U800 (N_800,N_757,N_768);
nand U801 (N_801,N_789,N_761);
and U802 (N_802,N_773,N_770);
and U803 (N_803,N_762,N_790);
xnor U804 (N_804,N_799,N_755);
and U805 (N_805,N_798,N_785);
xor U806 (N_806,N_781,N_780);
nor U807 (N_807,N_796,N_766);
or U808 (N_808,N_776,N_797);
nor U809 (N_809,N_791,N_779);
and U810 (N_810,N_777,N_784);
or U811 (N_811,N_758,N_795);
and U812 (N_812,N_759,N_771);
and U813 (N_813,N_769,N_752);
nor U814 (N_814,N_787,N_778);
xnor U815 (N_815,N_764,N_786);
and U816 (N_816,N_760,N_774);
and U817 (N_817,N_794,N_775);
nand U818 (N_818,N_751,N_753);
nor U819 (N_819,N_754,N_782);
and U820 (N_820,N_765,N_792);
or U821 (N_821,N_783,N_788);
nor U822 (N_822,N_750,N_763);
or U823 (N_823,N_793,N_756);
xnor U824 (N_824,N_772,N_767);
xor U825 (N_825,N_753,N_760);
nand U826 (N_826,N_774,N_767);
or U827 (N_827,N_793,N_784);
and U828 (N_828,N_785,N_760);
nand U829 (N_829,N_797,N_787);
nand U830 (N_830,N_759,N_777);
nand U831 (N_831,N_783,N_784);
nand U832 (N_832,N_750,N_753);
xor U833 (N_833,N_780,N_764);
or U834 (N_834,N_768,N_779);
nand U835 (N_835,N_765,N_796);
xor U836 (N_836,N_757,N_775);
nor U837 (N_837,N_773,N_760);
xor U838 (N_838,N_787,N_779);
xnor U839 (N_839,N_755,N_792);
and U840 (N_840,N_780,N_752);
or U841 (N_841,N_768,N_791);
and U842 (N_842,N_758,N_756);
and U843 (N_843,N_756,N_767);
xor U844 (N_844,N_795,N_755);
nand U845 (N_845,N_761,N_779);
or U846 (N_846,N_757,N_797);
xor U847 (N_847,N_762,N_792);
and U848 (N_848,N_752,N_754);
nor U849 (N_849,N_755,N_761);
xor U850 (N_850,N_820,N_808);
nor U851 (N_851,N_836,N_842);
and U852 (N_852,N_817,N_800);
nand U853 (N_853,N_844,N_812);
nand U854 (N_854,N_829,N_834);
and U855 (N_855,N_809,N_827);
nand U856 (N_856,N_815,N_801);
or U857 (N_857,N_822,N_841);
or U858 (N_858,N_824,N_849);
nand U859 (N_859,N_843,N_818);
or U860 (N_860,N_840,N_806);
or U861 (N_861,N_833,N_832);
nand U862 (N_862,N_811,N_813);
and U863 (N_863,N_803,N_831);
nor U864 (N_864,N_839,N_802);
nand U865 (N_865,N_823,N_814);
nand U866 (N_866,N_825,N_847);
xnor U867 (N_867,N_805,N_804);
nand U868 (N_868,N_846,N_845);
and U869 (N_869,N_826,N_835);
or U870 (N_870,N_838,N_810);
xnor U871 (N_871,N_830,N_807);
nand U872 (N_872,N_837,N_821);
nor U873 (N_873,N_816,N_819);
nor U874 (N_874,N_828,N_848);
or U875 (N_875,N_801,N_845);
and U876 (N_876,N_803,N_818);
xnor U877 (N_877,N_813,N_804);
and U878 (N_878,N_823,N_842);
nor U879 (N_879,N_804,N_841);
nor U880 (N_880,N_849,N_836);
xor U881 (N_881,N_834,N_809);
xor U882 (N_882,N_809,N_802);
nand U883 (N_883,N_812,N_822);
nand U884 (N_884,N_835,N_806);
nor U885 (N_885,N_805,N_812);
nand U886 (N_886,N_826,N_825);
and U887 (N_887,N_809,N_801);
or U888 (N_888,N_831,N_811);
nand U889 (N_889,N_805,N_836);
nor U890 (N_890,N_815,N_811);
and U891 (N_891,N_808,N_828);
nor U892 (N_892,N_800,N_838);
xor U893 (N_893,N_815,N_828);
or U894 (N_894,N_806,N_849);
xor U895 (N_895,N_804,N_838);
nand U896 (N_896,N_822,N_827);
nor U897 (N_897,N_848,N_835);
and U898 (N_898,N_819,N_847);
xnor U899 (N_899,N_849,N_820);
xnor U900 (N_900,N_885,N_886);
or U901 (N_901,N_864,N_873);
nand U902 (N_902,N_859,N_854);
or U903 (N_903,N_897,N_855);
or U904 (N_904,N_861,N_894);
and U905 (N_905,N_860,N_881);
or U906 (N_906,N_888,N_876);
or U907 (N_907,N_892,N_879);
or U908 (N_908,N_878,N_874);
xor U909 (N_909,N_856,N_890);
xor U910 (N_910,N_862,N_899);
or U911 (N_911,N_865,N_895);
nand U912 (N_912,N_870,N_868);
and U913 (N_913,N_867,N_850);
nor U914 (N_914,N_863,N_884);
nor U915 (N_915,N_893,N_882);
nand U916 (N_916,N_853,N_896);
xnor U917 (N_917,N_875,N_887);
nand U918 (N_918,N_871,N_880);
nor U919 (N_919,N_883,N_858);
or U920 (N_920,N_898,N_889);
nand U921 (N_921,N_852,N_869);
nand U922 (N_922,N_891,N_857);
nand U923 (N_923,N_872,N_851);
and U924 (N_924,N_866,N_877);
nor U925 (N_925,N_890,N_886);
nand U926 (N_926,N_875,N_871);
xnor U927 (N_927,N_880,N_864);
or U928 (N_928,N_896,N_857);
nor U929 (N_929,N_887,N_877);
or U930 (N_930,N_873,N_888);
and U931 (N_931,N_896,N_860);
and U932 (N_932,N_850,N_862);
or U933 (N_933,N_897,N_852);
nor U934 (N_934,N_871,N_893);
or U935 (N_935,N_888,N_889);
nor U936 (N_936,N_857,N_864);
and U937 (N_937,N_892,N_885);
nand U938 (N_938,N_887,N_891);
nor U939 (N_939,N_893,N_857);
or U940 (N_940,N_893,N_861);
nor U941 (N_941,N_875,N_892);
or U942 (N_942,N_857,N_875);
nand U943 (N_943,N_893,N_872);
nor U944 (N_944,N_887,N_864);
or U945 (N_945,N_890,N_887);
nor U946 (N_946,N_876,N_887);
xor U947 (N_947,N_855,N_862);
nor U948 (N_948,N_870,N_863);
and U949 (N_949,N_886,N_883);
and U950 (N_950,N_903,N_938);
nand U951 (N_951,N_906,N_912);
nand U952 (N_952,N_918,N_908);
and U953 (N_953,N_928,N_932);
nand U954 (N_954,N_943,N_923);
xnor U955 (N_955,N_921,N_916);
nor U956 (N_956,N_900,N_904);
or U957 (N_957,N_933,N_945);
nand U958 (N_958,N_937,N_939);
or U959 (N_959,N_946,N_941);
nand U960 (N_960,N_917,N_927);
and U961 (N_961,N_944,N_909);
xnor U962 (N_962,N_926,N_915);
nand U963 (N_963,N_920,N_949);
nand U964 (N_964,N_924,N_919);
or U965 (N_965,N_930,N_910);
and U966 (N_966,N_901,N_911);
nand U967 (N_967,N_922,N_914);
xnor U968 (N_968,N_934,N_907);
nand U969 (N_969,N_913,N_925);
nor U970 (N_970,N_936,N_929);
and U971 (N_971,N_902,N_931);
nor U972 (N_972,N_940,N_935);
and U973 (N_973,N_948,N_942);
or U974 (N_974,N_947,N_905);
or U975 (N_975,N_933,N_907);
nand U976 (N_976,N_910,N_948);
xnor U977 (N_977,N_905,N_904);
nand U978 (N_978,N_926,N_941);
nor U979 (N_979,N_907,N_911);
nor U980 (N_980,N_921,N_915);
nand U981 (N_981,N_933,N_931);
or U982 (N_982,N_902,N_901);
nor U983 (N_983,N_946,N_938);
or U984 (N_984,N_918,N_937);
nor U985 (N_985,N_931,N_925);
nand U986 (N_986,N_923,N_912);
or U987 (N_987,N_903,N_917);
or U988 (N_988,N_938,N_932);
nor U989 (N_989,N_909,N_936);
xnor U990 (N_990,N_901,N_943);
nor U991 (N_991,N_940,N_921);
nor U992 (N_992,N_916,N_929);
nand U993 (N_993,N_941,N_917);
and U994 (N_994,N_938,N_936);
and U995 (N_995,N_927,N_914);
nor U996 (N_996,N_909,N_919);
and U997 (N_997,N_912,N_933);
nor U998 (N_998,N_926,N_916);
and U999 (N_999,N_913,N_930);
nor U1000 (N_1000,N_966,N_964);
nand U1001 (N_1001,N_952,N_967);
nor U1002 (N_1002,N_965,N_982);
nand U1003 (N_1003,N_986,N_991);
or U1004 (N_1004,N_997,N_980);
or U1005 (N_1005,N_978,N_989);
nand U1006 (N_1006,N_976,N_993);
nor U1007 (N_1007,N_971,N_995);
nand U1008 (N_1008,N_984,N_994);
or U1009 (N_1009,N_990,N_960);
and U1010 (N_1010,N_958,N_973);
and U1011 (N_1011,N_968,N_981);
xor U1012 (N_1012,N_954,N_963);
or U1013 (N_1013,N_987,N_974);
nand U1014 (N_1014,N_969,N_950);
nand U1015 (N_1015,N_996,N_970);
xnor U1016 (N_1016,N_961,N_999);
and U1017 (N_1017,N_953,N_951);
nand U1018 (N_1018,N_957,N_983);
or U1019 (N_1019,N_972,N_955);
or U1020 (N_1020,N_988,N_998);
nor U1021 (N_1021,N_975,N_985);
or U1022 (N_1022,N_979,N_977);
and U1023 (N_1023,N_962,N_992);
nand U1024 (N_1024,N_959,N_956);
xnor U1025 (N_1025,N_985,N_967);
or U1026 (N_1026,N_955,N_956);
or U1027 (N_1027,N_959,N_966);
nand U1028 (N_1028,N_993,N_973);
and U1029 (N_1029,N_961,N_962);
and U1030 (N_1030,N_978,N_971);
nand U1031 (N_1031,N_958,N_962);
nand U1032 (N_1032,N_994,N_952);
or U1033 (N_1033,N_995,N_961);
xor U1034 (N_1034,N_979,N_997);
nor U1035 (N_1035,N_968,N_950);
and U1036 (N_1036,N_982,N_967);
and U1037 (N_1037,N_955,N_996);
or U1038 (N_1038,N_974,N_996);
nand U1039 (N_1039,N_958,N_954);
xnor U1040 (N_1040,N_960,N_981);
or U1041 (N_1041,N_979,N_961);
and U1042 (N_1042,N_981,N_999);
or U1043 (N_1043,N_955,N_979);
nand U1044 (N_1044,N_979,N_980);
nor U1045 (N_1045,N_966,N_974);
or U1046 (N_1046,N_969,N_967);
and U1047 (N_1047,N_974,N_992);
nor U1048 (N_1048,N_966,N_969);
nand U1049 (N_1049,N_974,N_957);
and U1050 (N_1050,N_1046,N_1009);
or U1051 (N_1051,N_1031,N_1048);
nand U1052 (N_1052,N_1001,N_1002);
nor U1053 (N_1053,N_1013,N_1000);
and U1054 (N_1054,N_1043,N_1014);
nor U1055 (N_1055,N_1030,N_1036);
or U1056 (N_1056,N_1015,N_1028);
or U1057 (N_1057,N_1049,N_1025);
or U1058 (N_1058,N_1003,N_1022);
or U1059 (N_1059,N_1007,N_1020);
xor U1060 (N_1060,N_1044,N_1012);
nor U1061 (N_1061,N_1029,N_1033);
xor U1062 (N_1062,N_1041,N_1018);
or U1063 (N_1063,N_1017,N_1024);
or U1064 (N_1064,N_1034,N_1016);
xnor U1065 (N_1065,N_1032,N_1004);
xor U1066 (N_1066,N_1008,N_1010);
or U1067 (N_1067,N_1035,N_1021);
nand U1068 (N_1068,N_1005,N_1026);
nor U1069 (N_1069,N_1045,N_1042);
xnor U1070 (N_1070,N_1037,N_1047);
nor U1071 (N_1071,N_1038,N_1011);
and U1072 (N_1072,N_1006,N_1040);
nor U1073 (N_1073,N_1023,N_1019);
nor U1074 (N_1074,N_1027,N_1039);
nor U1075 (N_1075,N_1008,N_1003);
nor U1076 (N_1076,N_1043,N_1000);
and U1077 (N_1077,N_1045,N_1017);
nand U1078 (N_1078,N_1046,N_1020);
nor U1079 (N_1079,N_1000,N_1020);
nor U1080 (N_1080,N_1018,N_1044);
nor U1081 (N_1081,N_1046,N_1023);
or U1082 (N_1082,N_1021,N_1032);
xnor U1083 (N_1083,N_1004,N_1002);
nor U1084 (N_1084,N_1005,N_1011);
xnor U1085 (N_1085,N_1017,N_1008);
nor U1086 (N_1086,N_1008,N_1024);
or U1087 (N_1087,N_1048,N_1003);
or U1088 (N_1088,N_1020,N_1024);
xor U1089 (N_1089,N_1013,N_1040);
nor U1090 (N_1090,N_1016,N_1048);
nor U1091 (N_1091,N_1039,N_1014);
nand U1092 (N_1092,N_1025,N_1032);
nand U1093 (N_1093,N_1028,N_1001);
nor U1094 (N_1094,N_1040,N_1020);
and U1095 (N_1095,N_1009,N_1044);
xnor U1096 (N_1096,N_1001,N_1014);
and U1097 (N_1097,N_1000,N_1048);
nand U1098 (N_1098,N_1032,N_1036);
and U1099 (N_1099,N_1028,N_1044);
nor U1100 (N_1100,N_1056,N_1097);
and U1101 (N_1101,N_1069,N_1078);
nand U1102 (N_1102,N_1085,N_1055);
xnor U1103 (N_1103,N_1072,N_1095);
and U1104 (N_1104,N_1073,N_1079);
and U1105 (N_1105,N_1092,N_1080);
or U1106 (N_1106,N_1087,N_1057);
xnor U1107 (N_1107,N_1068,N_1058);
or U1108 (N_1108,N_1070,N_1086);
and U1109 (N_1109,N_1083,N_1094);
xnor U1110 (N_1110,N_1088,N_1065);
xor U1111 (N_1111,N_1059,N_1099);
or U1112 (N_1112,N_1051,N_1053);
or U1113 (N_1113,N_1089,N_1077);
or U1114 (N_1114,N_1090,N_1067);
xnor U1115 (N_1115,N_1096,N_1052);
nor U1116 (N_1116,N_1098,N_1054);
and U1117 (N_1117,N_1064,N_1062);
or U1118 (N_1118,N_1066,N_1076);
and U1119 (N_1119,N_1082,N_1074);
xor U1120 (N_1120,N_1071,N_1075);
and U1121 (N_1121,N_1091,N_1063);
and U1122 (N_1122,N_1061,N_1081);
nand U1123 (N_1123,N_1050,N_1060);
xnor U1124 (N_1124,N_1093,N_1084);
or U1125 (N_1125,N_1051,N_1094);
nor U1126 (N_1126,N_1082,N_1089);
xor U1127 (N_1127,N_1075,N_1054);
or U1128 (N_1128,N_1053,N_1050);
or U1129 (N_1129,N_1062,N_1051);
nand U1130 (N_1130,N_1060,N_1065);
or U1131 (N_1131,N_1055,N_1069);
nand U1132 (N_1132,N_1051,N_1093);
and U1133 (N_1133,N_1056,N_1065);
nor U1134 (N_1134,N_1054,N_1079);
or U1135 (N_1135,N_1068,N_1089);
or U1136 (N_1136,N_1099,N_1078);
or U1137 (N_1137,N_1069,N_1090);
xnor U1138 (N_1138,N_1075,N_1050);
nand U1139 (N_1139,N_1066,N_1075);
xor U1140 (N_1140,N_1082,N_1054);
nand U1141 (N_1141,N_1074,N_1083);
and U1142 (N_1142,N_1064,N_1096);
and U1143 (N_1143,N_1097,N_1088);
or U1144 (N_1144,N_1072,N_1051);
or U1145 (N_1145,N_1071,N_1090);
xor U1146 (N_1146,N_1055,N_1091);
nor U1147 (N_1147,N_1054,N_1057);
xor U1148 (N_1148,N_1075,N_1068);
xor U1149 (N_1149,N_1081,N_1090);
nor U1150 (N_1150,N_1112,N_1143);
and U1151 (N_1151,N_1100,N_1113);
xnor U1152 (N_1152,N_1125,N_1122);
nand U1153 (N_1153,N_1146,N_1129);
xnor U1154 (N_1154,N_1141,N_1106);
nor U1155 (N_1155,N_1119,N_1111);
and U1156 (N_1156,N_1115,N_1108);
or U1157 (N_1157,N_1131,N_1117);
or U1158 (N_1158,N_1149,N_1105);
or U1159 (N_1159,N_1127,N_1139);
nor U1160 (N_1160,N_1107,N_1135);
and U1161 (N_1161,N_1132,N_1101);
xor U1162 (N_1162,N_1110,N_1134);
or U1163 (N_1163,N_1102,N_1137);
nand U1164 (N_1164,N_1140,N_1121);
xor U1165 (N_1165,N_1120,N_1104);
nor U1166 (N_1166,N_1145,N_1124);
or U1167 (N_1167,N_1133,N_1118);
nor U1168 (N_1168,N_1142,N_1116);
xnor U1169 (N_1169,N_1103,N_1138);
or U1170 (N_1170,N_1109,N_1144);
nand U1171 (N_1171,N_1147,N_1128);
and U1172 (N_1172,N_1126,N_1148);
or U1173 (N_1173,N_1114,N_1123);
or U1174 (N_1174,N_1130,N_1136);
nor U1175 (N_1175,N_1137,N_1118);
and U1176 (N_1176,N_1126,N_1128);
or U1177 (N_1177,N_1102,N_1127);
nor U1178 (N_1178,N_1115,N_1116);
xnor U1179 (N_1179,N_1115,N_1112);
or U1180 (N_1180,N_1101,N_1119);
nand U1181 (N_1181,N_1146,N_1105);
or U1182 (N_1182,N_1144,N_1117);
and U1183 (N_1183,N_1102,N_1111);
xnor U1184 (N_1184,N_1118,N_1140);
nand U1185 (N_1185,N_1146,N_1118);
or U1186 (N_1186,N_1124,N_1141);
nand U1187 (N_1187,N_1139,N_1126);
and U1188 (N_1188,N_1115,N_1104);
nand U1189 (N_1189,N_1121,N_1113);
and U1190 (N_1190,N_1124,N_1101);
or U1191 (N_1191,N_1133,N_1107);
xor U1192 (N_1192,N_1111,N_1101);
nor U1193 (N_1193,N_1123,N_1149);
xor U1194 (N_1194,N_1139,N_1106);
nand U1195 (N_1195,N_1101,N_1114);
nor U1196 (N_1196,N_1113,N_1108);
and U1197 (N_1197,N_1102,N_1103);
or U1198 (N_1198,N_1130,N_1147);
or U1199 (N_1199,N_1126,N_1133);
or U1200 (N_1200,N_1195,N_1164);
nand U1201 (N_1201,N_1162,N_1196);
xnor U1202 (N_1202,N_1189,N_1185);
nor U1203 (N_1203,N_1152,N_1187);
xnor U1204 (N_1204,N_1151,N_1150);
or U1205 (N_1205,N_1161,N_1153);
or U1206 (N_1206,N_1165,N_1188);
nor U1207 (N_1207,N_1182,N_1176);
or U1208 (N_1208,N_1194,N_1179);
or U1209 (N_1209,N_1170,N_1178);
xor U1210 (N_1210,N_1175,N_1180);
or U1211 (N_1211,N_1193,N_1168);
nand U1212 (N_1212,N_1177,N_1163);
nand U1213 (N_1213,N_1156,N_1154);
and U1214 (N_1214,N_1171,N_1167);
nand U1215 (N_1215,N_1158,N_1166);
xnor U1216 (N_1216,N_1181,N_1183);
nor U1217 (N_1217,N_1155,N_1157);
nor U1218 (N_1218,N_1198,N_1191);
nor U1219 (N_1219,N_1190,N_1186);
and U1220 (N_1220,N_1174,N_1173);
or U1221 (N_1221,N_1197,N_1169);
nor U1222 (N_1222,N_1199,N_1159);
nand U1223 (N_1223,N_1160,N_1172);
nand U1224 (N_1224,N_1184,N_1192);
nor U1225 (N_1225,N_1198,N_1182);
or U1226 (N_1226,N_1192,N_1162);
or U1227 (N_1227,N_1187,N_1182);
nand U1228 (N_1228,N_1171,N_1195);
nand U1229 (N_1229,N_1195,N_1180);
xnor U1230 (N_1230,N_1177,N_1181);
xnor U1231 (N_1231,N_1170,N_1163);
xnor U1232 (N_1232,N_1187,N_1150);
nor U1233 (N_1233,N_1178,N_1176);
nand U1234 (N_1234,N_1186,N_1171);
nand U1235 (N_1235,N_1162,N_1187);
nor U1236 (N_1236,N_1161,N_1181);
and U1237 (N_1237,N_1194,N_1171);
and U1238 (N_1238,N_1191,N_1153);
xor U1239 (N_1239,N_1172,N_1180);
and U1240 (N_1240,N_1150,N_1162);
and U1241 (N_1241,N_1183,N_1151);
or U1242 (N_1242,N_1157,N_1152);
and U1243 (N_1243,N_1173,N_1160);
nand U1244 (N_1244,N_1179,N_1167);
or U1245 (N_1245,N_1174,N_1194);
and U1246 (N_1246,N_1196,N_1190);
nor U1247 (N_1247,N_1155,N_1193);
nor U1248 (N_1248,N_1181,N_1160);
nand U1249 (N_1249,N_1168,N_1177);
xnor U1250 (N_1250,N_1247,N_1217);
or U1251 (N_1251,N_1235,N_1210);
xor U1252 (N_1252,N_1228,N_1214);
and U1253 (N_1253,N_1222,N_1221);
and U1254 (N_1254,N_1225,N_1245);
nor U1255 (N_1255,N_1213,N_1241);
and U1256 (N_1256,N_1238,N_1203);
xnor U1257 (N_1257,N_1209,N_1248);
or U1258 (N_1258,N_1232,N_1233);
nand U1259 (N_1259,N_1246,N_1223);
xor U1260 (N_1260,N_1237,N_1242);
nor U1261 (N_1261,N_1229,N_1211);
nand U1262 (N_1262,N_1236,N_1201);
nand U1263 (N_1263,N_1207,N_1219);
or U1264 (N_1264,N_1206,N_1230);
or U1265 (N_1265,N_1215,N_1200);
xor U1266 (N_1266,N_1249,N_1204);
or U1267 (N_1267,N_1202,N_1220);
xor U1268 (N_1268,N_1216,N_1243);
nor U1269 (N_1269,N_1226,N_1218);
xor U1270 (N_1270,N_1205,N_1231);
or U1271 (N_1271,N_1224,N_1239);
and U1272 (N_1272,N_1208,N_1227);
xnor U1273 (N_1273,N_1212,N_1240);
nor U1274 (N_1274,N_1244,N_1234);
xor U1275 (N_1275,N_1232,N_1237);
xnor U1276 (N_1276,N_1235,N_1232);
nand U1277 (N_1277,N_1231,N_1203);
nand U1278 (N_1278,N_1225,N_1218);
xor U1279 (N_1279,N_1247,N_1243);
nand U1280 (N_1280,N_1208,N_1228);
or U1281 (N_1281,N_1240,N_1205);
or U1282 (N_1282,N_1232,N_1215);
or U1283 (N_1283,N_1219,N_1213);
nand U1284 (N_1284,N_1240,N_1235);
nand U1285 (N_1285,N_1244,N_1220);
nor U1286 (N_1286,N_1244,N_1219);
xor U1287 (N_1287,N_1200,N_1229);
or U1288 (N_1288,N_1241,N_1201);
or U1289 (N_1289,N_1238,N_1212);
or U1290 (N_1290,N_1205,N_1224);
xor U1291 (N_1291,N_1224,N_1220);
nand U1292 (N_1292,N_1226,N_1208);
nand U1293 (N_1293,N_1205,N_1222);
nand U1294 (N_1294,N_1225,N_1236);
xor U1295 (N_1295,N_1244,N_1204);
and U1296 (N_1296,N_1230,N_1235);
or U1297 (N_1297,N_1211,N_1226);
or U1298 (N_1298,N_1245,N_1227);
nand U1299 (N_1299,N_1227,N_1201);
xor U1300 (N_1300,N_1283,N_1281);
nand U1301 (N_1301,N_1273,N_1263);
nor U1302 (N_1302,N_1274,N_1286);
nor U1303 (N_1303,N_1250,N_1282);
nor U1304 (N_1304,N_1255,N_1284);
xnor U1305 (N_1305,N_1289,N_1295);
or U1306 (N_1306,N_1292,N_1251);
xnor U1307 (N_1307,N_1285,N_1265);
and U1308 (N_1308,N_1287,N_1293);
nor U1309 (N_1309,N_1260,N_1298);
nor U1310 (N_1310,N_1267,N_1268);
nor U1311 (N_1311,N_1253,N_1252);
nand U1312 (N_1312,N_1299,N_1280);
nand U1313 (N_1313,N_1279,N_1276);
and U1314 (N_1314,N_1294,N_1254);
xor U1315 (N_1315,N_1261,N_1264);
or U1316 (N_1316,N_1266,N_1259);
nor U1317 (N_1317,N_1258,N_1256);
nor U1318 (N_1318,N_1262,N_1257);
nand U1319 (N_1319,N_1272,N_1278);
xor U1320 (N_1320,N_1296,N_1275);
or U1321 (N_1321,N_1277,N_1271);
nor U1322 (N_1322,N_1290,N_1270);
nand U1323 (N_1323,N_1269,N_1291);
nand U1324 (N_1324,N_1288,N_1297);
and U1325 (N_1325,N_1258,N_1294);
nand U1326 (N_1326,N_1280,N_1251);
nor U1327 (N_1327,N_1258,N_1270);
or U1328 (N_1328,N_1276,N_1263);
nand U1329 (N_1329,N_1260,N_1285);
nor U1330 (N_1330,N_1287,N_1281);
nand U1331 (N_1331,N_1250,N_1273);
and U1332 (N_1332,N_1277,N_1293);
nor U1333 (N_1333,N_1260,N_1251);
xnor U1334 (N_1334,N_1276,N_1297);
or U1335 (N_1335,N_1275,N_1254);
nor U1336 (N_1336,N_1259,N_1263);
nor U1337 (N_1337,N_1255,N_1278);
and U1338 (N_1338,N_1273,N_1260);
or U1339 (N_1339,N_1292,N_1288);
and U1340 (N_1340,N_1269,N_1265);
or U1341 (N_1341,N_1269,N_1258);
or U1342 (N_1342,N_1281,N_1282);
or U1343 (N_1343,N_1282,N_1280);
xor U1344 (N_1344,N_1272,N_1290);
or U1345 (N_1345,N_1263,N_1262);
or U1346 (N_1346,N_1298,N_1261);
or U1347 (N_1347,N_1290,N_1279);
xnor U1348 (N_1348,N_1255,N_1280);
and U1349 (N_1349,N_1269,N_1272);
or U1350 (N_1350,N_1309,N_1307);
nor U1351 (N_1351,N_1308,N_1336);
and U1352 (N_1352,N_1326,N_1338);
nor U1353 (N_1353,N_1328,N_1315);
and U1354 (N_1354,N_1304,N_1322);
nand U1355 (N_1355,N_1323,N_1327);
nor U1356 (N_1356,N_1337,N_1306);
nor U1357 (N_1357,N_1346,N_1302);
or U1358 (N_1358,N_1335,N_1342);
or U1359 (N_1359,N_1324,N_1340);
and U1360 (N_1360,N_1344,N_1318);
or U1361 (N_1361,N_1314,N_1341);
and U1362 (N_1362,N_1305,N_1339);
and U1363 (N_1363,N_1331,N_1329);
xnor U1364 (N_1364,N_1347,N_1345);
nor U1365 (N_1365,N_1300,N_1348);
and U1366 (N_1366,N_1310,N_1332);
and U1367 (N_1367,N_1349,N_1311);
nand U1368 (N_1368,N_1319,N_1303);
xor U1369 (N_1369,N_1330,N_1321);
or U1370 (N_1370,N_1320,N_1316);
nor U1371 (N_1371,N_1301,N_1312);
and U1372 (N_1372,N_1317,N_1325);
nand U1373 (N_1373,N_1334,N_1343);
or U1374 (N_1374,N_1313,N_1333);
xnor U1375 (N_1375,N_1310,N_1321);
nand U1376 (N_1376,N_1307,N_1328);
nor U1377 (N_1377,N_1330,N_1335);
nor U1378 (N_1378,N_1337,N_1328);
xnor U1379 (N_1379,N_1326,N_1322);
and U1380 (N_1380,N_1305,N_1317);
or U1381 (N_1381,N_1311,N_1346);
xor U1382 (N_1382,N_1344,N_1348);
nand U1383 (N_1383,N_1301,N_1309);
and U1384 (N_1384,N_1300,N_1313);
and U1385 (N_1385,N_1321,N_1339);
xnor U1386 (N_1386,N_1346,N_1338);
xnor U1387 (N_1387,N_1319,N_1315);
xor U1388 (N_1388,N_1340,N_1347);
xor U1389 (N_1389,N_1315,N_1302);
or U1390 (N_1390,N_1348,N_1341);
nor U1391 (N_1391,N_1322,N_1318);
nand U1392 (N_1392,N_1311,N_1329);
nor U1393 (N_1393,N_1300,N_1344);
nand U1394 (N_1394,N_1302,N_1311);
nor U1395 (N_1395,N_1338,N_1349);
nand U1396 (N_1396,N_1329,N_1330);
and U1397 (N_1397,N_1345,N_1318);
nand U1398 (N_1398,N_1328,N_1324);
nor U1399 (N_1399,N_1340,N_1311);
nand U1400 (N_1400,N_1367,N_1353);
and U1401 (N_1401,N_1381,N_1385);
xor U1402 (N_1402,N_1392,N_1356);
nor U1403 (N_1403,N_1386,N_1388);
nand U1404 (N_1404,N_1384,N_1372);
nand U1405 (N_1405,N_1359,N_1371);
nor U1406 (N_1406,N_1365,N_1389);
nor U1407 (N_1407,N_1379,N_1382);
and U1408 (N_1408,N_1374,N_1364);
and U1409 (N_1409,N_1395,N_1361);
or U1410 (N_1410,N_1396,N_1375);
nand U1411 (N_1411,N_1377,N_1355);
or U1412 (N_1412,N_1391,N_1383);
and U1413 (N_1413,N_1360,N_1390);
xnor U1414 (N_1414,N_1368,N_1393);
xor U1415 (N_1415,N_1354,N_1399);
nor U1416 (N_1416,N_1397,N_1358);
or U1417 (N_1417,N_1369,N_1376);
nand U1418 (N_1418,N_1378,N_1370);
nor U1419 (N_1419,N_1351,N_1352);
xnor U1420 (N_1420,N_1373,N_1350);
xor U1421 (N_1421,N_1394,N_1366);
and U1422 (N_1422,N_1362,N_1398);
nor U1423 (N_1423,N_1357,N_1380);
xor U1424 (N_1424,N_1363,N_1387);
xnor U1425 (N_1425,N_1382,N_1364);
nand U1426 (N_1426,N_1359,N_1361);
and U1427 (N_1427,N_1357,N_1396);
xor U1428 (N_1428,N_1388,N_1359);
or U1429 (N_1429,N_1387,N_1362);
nand U1430 (N_1430,N_1364,N_1368);
nand U1431 (N_1431,N_1372,N_1390);
nand U1432 (N_1432,N_1370,N_1354);
or U1433 (N_1433,N_1356,N_1388);
xor U1434 (N_1434,N_1370,N_1382);
and U1435 (N_1435,N_1362,N_1382);
nor U1436 (N_1436,N_1383,N_1350);
nor U1437 (N_1437,N_1371,N_1398);
and U1438 (N_1438,N_1382,N_1374);
xnor U1439 (N_1439,N_1370,N_1361);
and U1440 (N_1440,N_1357,N_1390);
and U1441 (N_1441,N_1386,N_1398);
xnor U1442 (N_1442,N_1387,N_1359);
xnor U1443 (N_1443,N_1396,N_1350);
or U1444 (N_1444,N_1366,N_1376);
xnor U1445 (N_1445,N_1367,N_1393);
and U1446 (N_1446,N_1393,N_1374);
xor U1447 (N_1447,N_1370,N_1368);
nor U1448 (N_1448,N_1352,N_1378);
and U1449 (N_1449,N_1372,N_1399);
xor U1450 (N_1450,N_1400,N_1421);
and U1451 (N_1451,N_1431,N_1430);
or U1452 (N_1452,N_1419,N_1446);
and U1453 (N_1453,N_1425,N_1428);
nor U1454 (N_1454,N_1444,N_1412);
nand U1455 (N_1455,N_1404,N_1437);
or U1456 (N_1456,N_1438,N_1447);
and U1457 (N_1457,N_1426,N_1435);
xor U1458 (N_1458,N_1449,N_1427);
nor U1459 (N_1459,N_1429,N_1411);
or U1460 (N_1460,N_1413,N_1434);
and U1461 (N_1461,N_1403,N_1416);
or U1462 (N_1462,N_1443,N_1424);
nor U1463 (N_1463,N_1405,N_1408);
nor U1464 (N_1464,N_1415,N_1433);
or U1465 (N_1465,N_1439,N_1402);
nand U1466 (N_1466,N_1406,N_1445);
nor U1467 (N_1467,N_1414,N_1422);
nor U1468 (N_1468,N_1417,N_1441);
xnor U1469 (N_1469,N_1410,N_1423);
nor U1470 (N_1470,N_1440,N_1432);
or U1471 (N_1471,N_1448,N_1407);
or U1472 (N_1472,N_1436,N_1409);
xnor U1473 (N_1473,N_1420,N_1418);
nand U1474 (N_1474,N_1442,N_1401);
nor U1475 (N_1475,N_1409,N_1406);
nand U1476 (N_1476,N_1444,N_1443);
xor U1477 (N_1477,N_1447,N_1417);
xor U1478 (N_1478,N_1415,N_1423);
nand U1479 (N_1479,N_1432,N_1435);
nor U1480 (N_1480,N_1424,N_1423);
xnor U1481 (N_1481,N_1425,N_1422);
or U1482 (N_1482,N_1432,N_1416);
and U1483 (N_1483,N_1425,N_1439);
or U1484 (N_1484,N_1411,N_1424);
or U1485 (N_1485,N_1443,N_1448);
xor U1486 (N_1486,N_1413,N_1409);
xor U1487 (N_1487,N_1432,N_1409);
and U1488 (N_1488,N_1410,N_1416);
and U1489 (N_1489,N_1444,N_1402);
or U1490 (N_1490,N_1425,N_1405);
or U1491 (N_1491,N_1446,N_1408);
xnor U1492 (N_1492,N_1406,N_1440);
and U1493 (N_1493,N_1429,N_1438);
or U1494 (N_1494,N_1449,N_1418);
or U1495 (N_1495,N_1437,N_1420);
nor U1496 (N_1496,N_1448,N_1414);
nand U1497 (N_1497,N_1434,N_1427);
nand U1498 (N_1498,N_1443,N_1434);
nand U1499 (N_1499,N_1432,N_1417);
nand U1500 (N_1500,N_1453,N_1454);
and U1501 (N_1501,N_1459,N_1473);
and U1502 (N_1502,N_1487,N_1468);
and U1503 (N_1503,N_1463,N_1480);
nor U1504 (N_1504,N_1460,N_1474);
xnor U1505 (N_1505,N_1451,N_1450);
or U1506 (N_1506,N_1458,N_1464);
xor U1507 (N_1507,N_1475,N_1483);
xor U1508 (N_1508,N_1497,N_1491);
nor U1509 (N_1509,N_1461,N_1485);
and U1510 (N_1510,N_1469,N_1457);
nand U1511 (N_1511,N_1479,N_1496);
xor U1512 (N_1512,N_1478,N_1456);
nand U1513 (N_1513,N_1495,N_1494);
and U1514 (N_1514,N_1492,N_1467);
nand U1515 (N_1515,N_1455,N_1486);
nand U1516 (N_1516,N_1471,N_1493);
xor U1517 (N_1517,N_1465,N_1477);
and U1518 (N_1518,N_1489,N_1466);
nand U1519 (N_1519,N_1476,N_1488);
nand U1520 (N_1520,N_1462,N_1490);
nand U1521 (N_1521,N_1470,N_1452);
nor U1522 (N_1522,N_1484,N_1499);
xnor U1523 (N_1523,N_1482,N_1481);
nand U1524 (N_1524,N_1472,N_1498);
xnor U1525 (N_1525,N_1452,N_1465);
and U1526 (N_1526,N_1461,N_1492);
xnor U1527 (N_1527,N_1456,N_1482);
or U1528 (N_1528,N_1477,N_1451);
nand U1529 (N_1529,N_1491,N_1464);
and U1530 (N_1530,N_1458,N_1473);
nor U1531 (N_1531,N_1473,N_1499);
xor U1532 (N_1532,N_1488,N_1495);
nor U1533 (N_1533,N_1473,N_1475);
xnor U1534 (N_1534,N_1484,N_1492);
and U1535 (N_1535,N_1469,N_1459);
nor U1536 (N_1536,N_1483,N_1460);
and U1537 (N_1537,N_1496,N_1481);
nand U1538 (N_1538,N_1497,N_1489);
nand U1539 (N_1539,N_1455,N_1475);
nor U1540 (N_1540,N_1455,N_1456);
and U1541 (N_1541,N_1479,N_1474);
nand U1542 (N_1542,N_1497,N_1456);
xnor U1543 (N_1543,N_1460,N_1465);
nor U1544 (N_1544,N_1469,N_1477);
nor U1545 (N_1545,N_1452,N_1479);
nand U1546 (N_1546,N_1478,N_1465);
nor U1547 (N_1547,N_1455,N_1464);
and U1548 (N_1548,N_1498,N_1490);
or U1549 (N_1549,N_1495,N_1472);
nand U1550 (N_1550,N_1518,N_1517);
or U1551 (N_1551,N_1538,N_1541);
nor U1552 (N_1552,N_1545,N_1532);
or U1553 (N_1553,N_1505,N_1534);
nor U1554 (N_1554,N_1525,N_1531);
or U1555 (N_1555,N_1522,N_1503);
or U1556 (N_1556,N_1520,N_1539);
or U1557 (N_1557,N_1542,N_1516);
nand U1558 (N_1558,N_1509,N_1537);
or U1559 (N_1559,N_1543,N_1527);
nand U1560 (N_1560,N_1502,N_1535);
xnor U1561 (N_1561,N_1501,N_1519);
nand U1562 (N_1562,N_1547,N_1530);
xnor U1563 (N_1563,N_1524,N_1526);
or U1564 (N_1564,N_1515,N_1546);
nor U1565 (N_1565,N_1513,N_1504);
and U1566 (N_1566,N_1544,N_1528);
and U1567 (N_1567,N_1549,N_1506);
nand U1568 (N_1568,N_1514,N_1529);
and U1569 (N_1569,N_1521,N_1540);
xor U1570 (N_1570,N_1511,N_1510);
and U1571 (N_1571,N_1523,N_1500);
and U1572 (N_1572,N_1548,N_1507);
and U1573 (N_1573,N_1512,N_1508);
and U1574 (N_1574,N_1536,N_1533);
nor U1575 (N_1575,N_1509,N_1521);
or U1576 (N_1576,N_1522,N_1514);
nor U1577 (N_1577,N_1546,N_1521);
nor U1578 (N_1578,N_1512,N_1500);
nand U1579 (N_1579,N_1510,N_1547);
xnor U1580 (N_1580,N_1533,N_1505);
nand U1581 (N_1581,N_1522,N_1510);
or U1582 (N_1582,N_1525,N_1537);
nor U1583 (N_1583,N_1544,N_1546);
or U1584 (N_1584,N_1543,N_1547);
or U1585 (N_1585,N_1537,N_1517);
xnor U1586 (N_1586,N_1512,N_1531);
xnor U1587 (N_1587,N_1537,N_1508);
and U1588 (N_1588,N_1549,N_1532);
nor U1589 (N_1589,N_1508,N_1528);
and U1590 (N_1590,N_1504,N_1506);
and U1591 (N_1591,N_1545,N_1502);
xnor U1592 (N_1592,N_1527,N_1528);
and U1593 (N_1593,N_1510,N_1533);
or U1594 (N_1594,N_1526,N_1525);
xor U1595 (N_1595,N_1529,N_1548);
xnor U1596 (N_1596,N_1524,N_1549);
nand U1597 (N_1597,N_1540,N_1505);
or U1598 (N_1598,N_1513,N_1528);
nand U1599 (N_1599,N_1541,N_1526);
and U1600 (N_1600,N_1567,N_1597);
or U1601 (N_1601,N_1553,N_1585);
nand U1602 (N_1602,N_1581,N_1565);
xnor U1603 (N_1603,N_1576,N_1561);
nand U1604 (N_1604,N_1575,N_1552);
or U1605 (N_1605,N_1595,N_1559);
or U1606 (N_1606,N_1558,N_1584);
or U1607 (N_1607,N_1599,N_1564);
or U1608 (N_1608,N_1568,N_1587);
nand U1609 (N_1609,N_1582,N_1580);
xnor U1610 (N_1610,N_1573,N_1569);
or U1611 (N_1611,N_1556,N_1586);
nor U1612 (N_1612,N_1570,N_1562);
xnor U1613 (N_1613,N_1557,N_1593);
or U1614 (N_1614,N_1590,N_1594);
nor U1615 (N_1615,N_1554,N_1572);
xor U1616 (N_1616,N_1578,N_1579);
xnor U1617 (N_1617,N_1588,N_1574);
nor U1618 (N_1618,N_1551,N_1583);
xnor U1619 (N_1619,N_1577,N_1592);
nor U1620 (N_1620,N_1566,N_1598);
nand U1621 (N_1621,N_1591,N_1555);
or U1622 (N_1622,N_1589,N_1563);
nor U1623 (N_1623,N_1596,N_1550);
nand U1624 (N_1624,N_1571,N_1560);
or U1625 (N_1625,N_1599,N_1573);
and U1626 (N_1626,N_1588,N_1560);
nor U1627 (N_1627,N_1594,N_1585);
and U1628 (N_1628,N_1594,N_1568);
and U1629 (N_1629,N_1582,N_1550);
nor U1630 (N_1630,N_1569,N_1598);
and U1631 (N_1631,N_1568,N_1567);
nor U1632 (N_1632,N_1580,N_1572);
nand U1633 (N_1633,N_1574,N_1595);
and U1634 (N_1634,N_1574,N_1585);
nand U1635 (N_1635,N_1577,N_1568);
xnor U1636 (N_1636,N_1560,N_1585);
and U1637 (N_1637,N_1573,N_1557);
xnor U1638 (N_1638,N_1567,N_1592);
nor U1639 (N_1639,N_1598,N_1550);
nor U1640 (N_1640,N_1564,N_1597);
nor U1641 (N_1641,N_1567,N_1550);
and U1642 (N_1642,N_1596,N_1575);
nor U1643 (N_1643,N_1580,N_1579);
or U1644 (N_1644,N_1592,N_1590);
nor U1645 (N_1645,N_1559,N_1560);
or U1646 (N_1646,N_1596,N_1592);
nand U1647 (N_1647,N_1556,N_1561);
and U1648 (N_1648,N_1578,N_1550);
xor U1649 (N_1649,N_1599,N_1588);
xnor U1650 (N_1650,N_1646,N_1621);
nor U1651 (N_1651,N_1634,N_1632);
and U1652 (N_1652,N_1609,N_1644);
xor U1653 (N_1653,N_1619,N_1612);
nor U1654 (N_1654,N_1615,N_1633);
or U1655 (N_1655,N_1629,N_1608);
or U1656 (N_1656,N_1642,N_1626);
xnor U1657 (N_1657,N_1622,N_1648);
nand U1658 (N_1658,N_1649,N_1643);
nand U1659 (N_1659,N_1617,N_1627);
nand U1660 (N_1660,N_1625,N_1631);
nand U1661 (N_1661,N_1607,N_1616);
nor U1662 (N_1662,N_1604,N_1623);
xor U1663 (N_1663,N_1645,N_1640);
nand U1664 (N_1664,N_1624,N_1635);
nor U1665 (N_1665,N_1613,N_1647);
nor U1666 (N_1666,N_1620,N_1606);
and U1667 (N_1667,N_1600,N_1636);
xor U1668 (N_1668,N_1618,N_1639);
and U1669 (N_1669,N_1638,N_1610);
nor U1670 (N_1670,N_1601,N_1603);
and U1671 (N_1671,N_1605,N_1602);
nor U1672 (N_1672,N_1637,N_1641);
and U1673 (N_1673,N_1614,N_1630);
nand U1674 (N_1674,N_1628,N_1611);
nand U1675 (N_1675,N_1624,N_1615);
xor U1676 (N_1676,N_1602,N_1612);
or U1677 (N_1677,N_1614,N_1648);
and U1678 (N_1678,N_1601,N_1607);
nand U1679 (N_1679,N_1637,N_1633);
nand U1680 (N_1680,N_1638,N_1615);
or U1681 (N_1681,N_1634,N_1602);
nand U1682 (N_1682,N_1628,N_1637);
nand U1683 (N_1683,N_1629,N_1606);
and U1684 (N_1684,N_1630,N_1634);
xnor U1685 (N_1685,N_1618,N_1608);
xnor U1686 (N_1686,N_1617,N_1637);
and U1687 (N_1687,N_1638,N_1619);
or U1688 (N_1688,N_1623,N_1626);
nand U1689 (N_1689,N_1643,N_1603);
and U1690 (N_1690,N_1627,N_1644);
xor U1691 (N_1691,N_1628,N_1622);
and U1692 (N_1692,N_1600,N_1605);
or U1693 (N_1693,N_1614,N_1600);
xor U1694 (N_1694,N_1605,N_1622);
nand U1695 (N_1695,N_1638,N_1601);
or U1696 (N_1696,N_1617,N_1642);
nand U1697 (N_1697,N_1634,N_1617);
xor U1698 (N_1698,N_1614,N_1604);
and U1699 (N_1699,N_1610,N_1648);
or U1700 (N_1700,N_1696,N_1680);
nor U1701 (N_1701,N_1691,N_1652);
or U1702 (N_1702,N_1670,N_1684);
xor U1703 (N_1703,N_1651,N_1663);
xor U1704 (N_1704,N_1672,N_1673);
or U1705 (N_1705,N_1662,N_1678);
and U1706 (N_1706,N_1679,N_1661);
nor U1707 (N_1707,N_1695,N_1676);
and U1708 (N_1708,N_1658,N_1683);
nor U1709 (N_1709,N_1653,N_1688);
or U1710 (N_1710,N_1674,N_1693);
nand U1711 (N_1711,N_1655,N_1685);
and U1712 (N_1712,N_1671,N_1666);
nand U1713 (N_1713,N_1694,N_1664);
and U1714 (N_1714,N_1660,N_1682);
xor U1715 (N_1715,N_1698,N_1687);
or U1716 (N_1716,N_1686,N_1692);
nor U1717 (N_1717,N_1668,N_1689);
or U1718 (N_1718,N_1657,N_1669);
nor U1719 (N_1719,N_1699,N_1677);
nor U1720 (N_1720,N_1681,N_1667);
or U1721 (N_1721,N_1675,N_1650);
or U1722 (N_1722,N_1665,N_1659);
nor U1723 (N_1723,N_1654,N_1690);
or U1724 (N_1724,N_1656,N_1697);
nand U1725 (N_1725,N_1665,N_1668);
nor U1726 (N_1726,N_1651,N_1660);
or U1727 (N_1727,N_1662,N_1699);
and U1728 (N_1728,N_1691,N_1663);
or U1729 (N_1729,N_1661,N_1662);
nor U1730 (N_1730,N_1668,N_1657);
or U1731 (N_1731,N_1677,N_1694);
or U1732 (N_1732,N_1653,N_1672);
nor U1733 (N_1733,N_1667,N_1671);
xnor U1734 (N_1734,N_1653,N_1660);
and U1735 (N_1735,N_1690,N_1692);
nand U1736 (N_1736,N_1697,N_1665);
xor U1737 (N_1737,N_1691,N_1662);
nor U1738 (N_1738,N_1685,N_1656);
nor U1739 (N_1739,N_1672,N_1651);
xor U1740 (N_1740,N_1650,N_1655);
nor U1741 (N_1741,N_1673,N_1677);
nor U1742 (N_1742,N_1653,N_1689);
xor U1743 (N_1743,N_1683,N_1699);
or U1744 (N_1744,N_1670,N_1663);
or U1745 (N_1745,N_1697,N_1650);
xor U1746 (N_1746,N_1651,N_1650);
nand U1747 (N_1747,N_1695,N_1675);
xnor U1748 (N_1748,N_1674,N_1667);
and U1749 (N_1749,N_1672,N_1692);
and U1750 (N_1750,N_1713,N_1730);
nand U1751 (N_1751,N_1705,N_1729);
nand U1752 (N_1752,N_1738,N_1710);
or U1753 (N_1753,N_1727,N_1743);
xor U1754 (N_1754,N_1715,N_1740);
or U1755 (N_1755,N_1701,N_1732);
and U1756 (N_1756,N_1726,N_1724);
nand U1757 (N_1757,N_1736,N_1745);
and U1758 (N_1758,N_1739,N_1748);
xnor U1759 (N_1759,N_1714,N_1728);
or U1760 (N_1760,N_1703,N_1747);
and U1761 (N_1761,N_1711,N_1721);
nand U1762 (N_1762,N_1731,N_1704);
or U1763 (N_1763,N_1702,N_1706);
and U1764 (N_1764,N_1733,N_1725);
xor U1765 (N_1765,N_1719,N_1707);
nor U1766 (N_1766,N_1749,N_1723);
or U1767 (N_1767,N_1744,N_1700);
and U1768 (N_1768,N_1712,N_1737);
xnor U1769 (N_1769,N_1709,N_1720);
xnor U1770 (N_1770,N_1708,N_1722);
nor U1771 (N_1771,N_1716,N_1717);
and U1772 (N_1772,N_1741,N_1735);
nand U1773 (N_1773,N_1734,N_1718);
xnor U1774 (N_1774,N_1742,N_1746);
nand U1775 (N_1775,N_1715,N_1729);
and U1776 (N_1776,N_1701,N_1733);
and U1777 (N_1777,N_1707,N_1730);
nand U1778 (N_1778,N_1724,N_1722);
nand U1779 (N_1779,N_1724,N_1734);
or U1780 (N_1780,N_1717,N_1707);
nand U1781 (N_1781,N_1736,N_1705);
nand U1782 (N_1782,N_1723,N_1742);
xor U1783 (N_1783,N_1743,N_1710);
xnor U1784 (N_1784,N_1734,N_1710);
xor U1785 (N_1785,N_1739,N_1737);
and U1786 (N_1786,N_1731,N_1705);
and U1787 (N_1787,N_1744,N_1723);
or U1788 (N_1788,N_1708,N_1737);
xnor U1789 (N_1789,N_1736,N_1729);
nand U1790 (N_1790,N_1710,N_1727);
and U1791 (N_1791,N_1734,N_1729);
nor U1792 (N_1792,N_1707,N_1731);
nand U1793 (N_1793,N_1749,N_1713);
or U1794 (N_1794,N_1719,N_1734);
or U1795 (N_1795,N_1705,N_1742);
and U1796 (N_1796,N_1705,N_1733);
nor U1797 (N_1797,N_1726,N_1713);
nand U1798 (N_1798,N_1700,N_1747);
xnor U1799 (N_1799,N_1712,N_1717);
and U1800 (N_1800,N_1793,N_1757);
or U1801 (N_1801,N_1781,N_1767);
or U1802 (N_1802,N_1797,N_1766);
or U1803 (N_1803,N_1795,N_1768);
or U1804 (N_1804,N_1774,N_1796);
or U1805 (N_1805,N_1765,N_1783);
xnor U1806 (N_1806,N_1763,N_1778);
nand U1807 (N_1807,N_1780,N_1787);
nor U1808 (N_1808,N_1786,N_1798);
xnor U1809 (N_1809,N_1760,N_1782);
xnor U1810 (N_1810,N_1751,N_1775);
nor U1811 (N_1811,N_1758,N_1771);
and U1812 (N_1812,N_1791,N_1772);
xnor U1813 (N_1813,N_1794,N_1759);
nand U1814 (N_1814,N_1769,N_1789);
and U1815 (N_1815,N_1761,N_1784);
or U1816 (N_1816,N_1755,N_1788);
or U1817 (N_1817,N_1776,N_1790);
and U1818 (N_1818,N_1753,N_1799);
nor U1819 (N_1819,N_1764,N_1756);
xnor U1820 (N_1820,N_1792,N_1785);
and U1821 (N_1821,N_1754,N_1750);
nand U1822 (N_1822,N_1773,N_1752);
nand U1823 (N_1823,N_1777,N_1770);
and U1824 (N_1824,N_1779,N_1762);
and U1825 (N_1825,N_1794,N_1788);
nand U1826 (N_1826,N_1768,N_1785);
nand U1827 (N_1827,N_1792,N_1768);
or U1828 (N_1828,N_1799,N_1766);
or U1829 (N_1829,N_1799,N_1763);
and U1830 (N_1830,N_1793,N_1799);
xnor U1831 (N_1831,N_1783,N_1796);
nor U1832 (N_1832,N_1793,N_1780);
and U1833 (N_1833,N_1790,N_1795);
nand U1834 (N_1834,N_1758,N_1785);
xnor U1835 (N_1835,N_1760,N_1797);
nand U1836 (N_1836,N_1771,N_1772);
and U1837 (N_1837,N_1780,N_1755);
xnor U1838 (N_1838,N_1758,N_1787);
or U1839 (N_1839,N_1763,N_1791);
xor U1840 (N_1840,N_1760,N_1766);
nor U1841 (N_1841,N_1773,N_1772);
and U1842 (N_1842,N_1756,N_1754);
and U1843 (N_1843,N_1791,N_1787);
and U1844 (N_1844,N_1785,N_1797);
and U1845 (N_1845,N_1769,N_1771);
or U1846 (N_1846,N_1763,N_1756);
nand U1847 (N_1847,N_1768,N_1754);
and U1848 (N_1848,N_1776,N_1797);
and U1849 (N_1849,N_1777,N_1756);
xor U1850 (N_1850,N_1808,N_1836);
xor U1851 (N_1851,N_1827,N_1820);
and U1852 (N_1852,N_1841,N_1837);
xor U1853 (N_1853,N_1840,N_1844);
nand U1854 (N_1854,N_1845,N_1833);
xor U1855 (N_1855,N_1810,N_1839);
and U1856 (N_1856,N_1848,N_1821);
nand U1857 (N_1857,N_1814,N_1843);
nand U1858 (N_1858,N_1838,N_1805);
and U1859 (N_1859,N_1812,N_1803);
and U1860 (N_1860,N_1816,N_1807);
xor U1861 (N_1861,N_1823,N_1835);
and U1862 (N_1862,N_1811,N_1828);
nor U1863 (N_1863,N_1802,N_1831);
nor U1864 (N_1864,N_1815,N_1822);
xor U1865 (N_1865,N_1846,N_1829);
or U1866 (N_1866,N_1819,N_1813);
nand U1867 (N_1867,N_1826,N_1800);
xor U1868 (N_1868,N_1806,N_1824);
xnor U1869 (N_1869,N_1801,N_1817);
and U1870 (N_1870,N_1804,N_1818);
nor U1871 (N_1871,N_1830,N_1834);
nor U1872 (N_1872,N_1847,N_1832);
nand U1873 (N_1873,N_1809,N_1849);
and U1874 (N_1874,N_1842,N_1825);
nand U1875 (N_1875,N_1833,N_1827);
or U1876 (N_1876,N_1845,N_1805);
xor U1877 (N_1877,N_1843,N_1812);
and U1878 (N_1878,N_1828,N_1808);
nand U1879 (N_1879,N_1842,N_1841);
xor U1880 (N_1880,N_1801,N_1808);
nor U1881 (N_1881,N_1816,N_1830);
nand U1882 (N_1882,N_1814,N_1848);
or U1883 (N_1883,N_1806,N_1825);
or U1884 (N_1884,N_1847,N_1808);
xnor U1885 (N_1885,N_1806,N_1821);
xor U1886 (N_1886,N_1835,N_1810);
nand U1887 (N_1887,N_1806,N_1847);
nand U1888 (N_1888,N_1811,N_1824);
and U1889 (N_1889,N_1843,N_1816);
and U1890 (N_1890,N_1836,N_1846);
nand U1891 (N_1891,N_1823,N_1810);
and U1892 (N_1892,N_1812,N_1841);
nor U1893 (N_1893,N_1833,N_1808);
nor U1894 (N_1894,N_1844,N_1841);
xnor U1895 (N_1895,N_1815,N_1825);
nor U1896 (N_1896,N_1811,N_1849);
nor U1897 (N_1897,N_1802,N_1842);
nand U1898 (N_1898,N_1819,N_1843);
xnor U1899 (N_1899,N_1825,N_1839);
and U1900 (N_1900,N_1889,N_1872);
nor U1901 (N_1901,N_1857,N_1896);
or U1902 (N_1902,N_1874,N_1886);
and U1903 (N_1903,N_1852,N_1862);
or U1904 (N_1904,N_1894,N_1882);
nor U1905 (N_1905,N_1885,N_1863);
or U1906 (N_1906,N_1895,N_1856);
nand U1907 (N_1907,N_1854,N_1853);
or U1908 (N_1908,N_1884,N_1851);
nor U1909 (N_1909,N_1887,N_1861);
nand U1910 (N_1910,N_1873,N_1883);
or U1911 (N_1911,N_1891,N_1855);
nor U1912 (N_1912,N_1878,N_1850);
or U1913 (N_1913,N_1897,N_1877);
or U1914 (N_1914,N_1865,N_1888);
xor U1915 (N_1915,N_1869,N_1871);
xor U1916 (N_1916,N_1881,N_1893);
nor U1917 (N_1917,N_1858,N_1875);
xor U1918 (N_1918,N_1864,N_1859);
nand U1919 (N_1919,N_1870,N_1879);
nor U1920 (N_1920,N_1866,N_1867);
xnor U1921 (N_1921,N_1892,N_1860);
nor U1922 (N_1922,N_1890,N_1898);
nor U1923 (N_1923,N_1868,N_1876);
or U1924 (N_1924,N_1899,N_1880);
xor U1925 (N_1925,N_1883,N_1858);
or U1926 (N_1926,N_1853,N_1897);
or U1927 (N_1927,N_1865,N_1893);
nand U1928 (N_1928,N_1881,N_1876);
or U1929 (N_1929,N_1856,N_1850);
nor U1930 (N_1930,N_1891,N_1850);
or U1931 (N_1931,N_1867,N_1854);
or U1932 (N_1932,N_1883,N_1855);
and U1933 (N_1933,N_1882,N_1877);
or U1934 (N_1934,N_1853,N_1861);
nand U1935 (N_1935,N_1896,N_1873);
nand U1936 (N_1936,N_1874,N_1872);
nor U1937 (N_1937,N_1868,N_1850);
or U1938 (N_1938,N_1877,N_1853);
xnor U1939 (N_1939,N_1851,N_1850);
or U1940 (N_1940,N_1880,N_1866);
and U1941 (N_1941,N_1885,N_1861);
nor U1942 (N_1942,N_1889,N_1861);
nor U1943 (N_1943,N_1871,N_1895);
and U1944 (N_1944,N_1878,N_1873);
and U1945 (N_1945,N_1869,N_1889);
nor U1946 (N_1946,N_1856,N_1871);
xnor U1947 (N_1947,N_1870,N_1863);
or U1948 (N_1948,N_1894,N_1888);
and U1949 (N_1949,N_1883,N_1862);
nand U1950 (N_1950,N_1902,N_1911);
nor U1951 (N_1951,N_1935,N_1926);
or U1952 (N_1952,N_1936,N_1920);
and U1953 (N_1953,N_1913,N_1947);
or U1954 (N_1954,N_1908,N_1918);
xor U1955 (N_1955,N_1919,N_1939);
and U1956 (N_1956,N_1941,N_1938);
or U1957 (N_1957,N_1949,N_1937);
and U1958 (N_1958,N_1930,N_1910);
and U1959 (N_1959,N_1931,N_1907);
xor U1960 (N_1960,N_1933,N_1915);
or U1961 (N_1961,N_1916,N_1901);
nor U1962 (N_1962,N_1924,N_1943);
nand U1963 (N_1963,N_1905,N_1940);
nor U1964 (N_1964,N_1925,N_1900);
nor U1965 (N_1965,N_1914,N_1922);
nand U1966 (N_1966,N_1917,N_1934);
or U1967 (N_1967,N_1904,N_1944);
or U1968 (N_1968,N_1946,N_1903);
nand U1969 (N_1969,N_1942,N_1928);
nand U1970 (N_1970,N_1945,N_1927);
and U1971 (N_1971,N_1923,N_1932);
or U1972 (N_1972,N_1909,N_1929);
xnor U1973 (N_1973,N_1906,N_1912);
or U1974 (N_1974,N_1948,N_1921);
and U1975 (N_1975,N_1915,N_1943);
and U1976 (N_1976,N_1920,N_1939);
and U1977 (N_1977,N_1930,N_1943);
or U1978 (N_1978,N_1937,N_1917);
xnor U1979 (N_1979,N_1927,N_1916);
or U1980 (N_1980,N_1904,N_1918);
nand U1981 (N_1981,N_1931,N_1925);
and U1982 (N_1982,N_1925,N_1901);
nor U1983 (N_1983,N_1901,N_1911);
and U1984 (N_1984,N_1934,N_1903);
or U1985 (N_1985,N_1930,N_1914);
nor U1986 (N_1986,N_1927,N_1912);
nand U1987 (N_1987,N_1912,N_1918);
and U1988 (N_1988,N_1911,N_1946);
xnor U1989 (N_1989,N_1919,N_1912);
xor U1990 (N_1990,N_1931,N_1928);
or U1991 (N_1991,N_1926,N_1947);
or U1992 (N_1992,N_1906,N_1907);
and U1993 (N_1993,N_1936,N_1913);
xor U1994 (N_1994,N_1928,N_1910);
nand U1995 (N_1995,N_1926,N_1932);
nand U1996 (N_1996,N_1932,N_1901);
and U1997 (N_1997,N_1939,N_1943);
xor U1998 (N_1998,N_1926,N_1936);
or U1999 (N_1999,N_1923,N_1903);
nand U2000 (N_2000,N_1976,N_1960);
nand U2001 (N_2001,N_1974,N_1996);
nand U2002 (N_2002,N_1969,N_1997);
nand U2003 (N_2003,N_1972,N_1952);
nand U2004 (N_2004,N_1970,N_1994);
xnor U2005 (N_2005,N_1962,N_1993);
or U2006 (N_2006,N_1951,N_1954);
and U2007 (N_2007,N_1963,N_1959);
and U2008 (N_2008,N_1983,N_1967);
nor U2009 (N_2009,N_1985,N_1984);
nand U2010 (N_2010,N_1968,N_1957);
and U2011 (N_2011,N_1979,N_1980);
or U2012 (N_2012,N_1955,N_1953);
or U2013 (N_2013,N_1989,N_1998);
or U2014 (N_2014,N_1977,N_1995);
xor U2015 (N_2015,N_1965,N_1956);
and U2016 (N_2016,N_1950,N_1975);
or U2017 (N_2017,N_1991,N_1986);
or U2018 (N_2018,N_1992,N_1973);
nor U2019 (N_2019,N_1990,N_1961);
nor U2020 (N_2020,N_1987,N_1958);
xor U2021 (N_2021,N_1964,N_1988);
nor U2022 (N_2022,N_1981,N_1978);
or U2023 (N_2023,N_1966,N_1971);
or U2024 (N_2024,N_1982,N_1999);
and U2025 (N_2025,N_1982,N_1981);
xor U2026 (N_2026,N_1989,N_1981);
xnor U2027 (N_2027,N_1951,N_1965);
nor U2028 (N_2028,N_1994,N_1977);
or U2029 (N_2029,N_1957,N_1998);
nand U2030 (N_2030,N_1996,N_1976);
xnor U2031 (N_2031,N_1957,N_1982);
nand U2032 (N_2032,N_1950,N_1998);
xnor U2033 (N_2033,N_1967,N_1954);
nor U2034 (N_2034,N_1969,N_1980);
and U2035 (N_2035,N_1987,N_1995);
or U2036 (N_2036,N_1986,N_1964);
nand U2037 (N_2037,N_1962,N_1958);
and U2038 (N_2038,N_1993,N_1951);
nor U2039 (N_2039,N_1974,N_1950);
nor U2040 (N_2040,N_1974,N_1992);
or U2041 (N_2041,N_1961,N_1965);
or U2042 (N_2042,N_1969,N_1973);
nor U2043 (N_2043,N_1980,N_1962);
xor U2044 (N_2044,N_1974,N_1959);
nor U2045 (N_2045,N_1985,N_1956);
nand U2046 (N_2046,N_1997,N_1990);
and U2047 (N_2047,N_1956,N_1986);
nand U2048 (N_2048,N_1984,N_1974);
nor U2049 (N_2049,N_1959,N_1960);
and U2050 (N_2050,N_2028,N_2004);
nor U2051 (N_2051,N_2047,N_2038);
nand U2052 (N_2052,N_2040,N_2029);
nand U2053 (N_2053,N_2044,N_2016);
and U2054 (N_2054,N_2042,N_2003);
nor U2055 (N_2055,N_2014,N_2033);
and U2056 (N_2056,N_2011,N_2012);
nand U2057 (N_2057,N_2043,N_2030);
and U2058 (N_2058,N_2005,N_2045);
or U2059 (N_2059,N_2036,N_2041);
or U2060 (N_2060,N_2001,N_2024);
or U2061 (N_2061,N_2009,N_2027);
and U2062 (N_2062,N_2032,N_2013);
nor U2063 (N_2063,N_2048,N_2022);
or U2064 (N_2064,N_2020,N_2018);
or U2065 (N_2065,N_2000,N_2031);
nand U2066 (N_2066,N_2025,N_2046);
nand U2067 (N_2067,N_2006,N_2010);
and U2068 (N_2068,N_2002,N_2019);
nor U2069 (N_2069,N_2026,N_2015);
xnor U2070 (N_2070,N_2023,N_2049);
nand U2071 (N_2071,N_2007,N_2008);
nand U2072 (N_2072,N_2037,N_2035);
or U2073 (N_2073,N_2021,N_2039);
or U2074 (N_2074,N_2034,N_2017);
and U2075 (N_2075,N_2011,N_2010);
nand U2076 (N_2076,N_2025,N_2030);
and U2077 (N_2077,N_2014,N_2020);
and U2078 (N_2078,N_2018,N_2047);
and U2079 (N_2079,N_2034,N_2021);
nand U2080 (N_2080,N_2018,N_2011);
and U2081 (N_2081,N_2027,N_2005);
or U2082 (N_2082,N_2031,N_2025);
nand U2083 (N_2083,N_2038,N_2008);
and U2084 (N_2084,N_2025,N_2033);
or U2085 (N_2085,N_2024,N_2010);
and U2086 (N_2086,N_2003,N_2021);
nand U2087 (N_2087,N_2000,N_2037);
or U2088 (N_2088,N_2035,N_2032);
and U2089 (N_2089,N_2033,N_2013);
nand U2090 (N_2090,N_2021,N_2005);
and U2091 (N_2091,N_2044,N_2020);
xor U2092 (N_2092,N_2032,N_2031);
xnor U2093 (N_2093,N_2044,N_2049);
or U2094 (N_2094,N_2009,N_2006);
nand U2095 (N_2095,N_2025,N_2024);
or U2096 (N_2096,N_2044,N_2000);
nor U2097 (N_2097,N_2017,N_2048);
nand U2098 (N_2098,N_2018,N_2032);
nand U2099 (N_2099,N_2009,N_2015);
or U2100 (N_2100,N_2099,N_2058);
and U2101 (N_2101,N_2071,N_2074);
or U2102 (N_2102,N_2061,N_2070);
and U2103 (N_2103,N_2089,N_2097);
nor U2104 (N_2104,N_2073,N_2092);
nor U2105 (N_2105,N_2095,N_2065);
or U2106 (N_2106,N_2067,N_2093);
or U2107 (N_2107,N_2091,N_2051);
xor U2108 (N_2108,N_2098,N_2054);
nand U2109 (N_2109,N_2060,N_2080);
nand U2110 (N_2110,N_2055,N_2081);
xor U2111 (N_2111,N_2086,N_2079);
and U2112 (N_2112,N_2076,N_2077);
xor U2113 (N_2113,N_2087,N_2057);
nor U2114 (N_2114,N_2063,N_2053);
nand U2115 (N_2115,N_2088,N_2075);
nand U2116 (N_2116,N_2072,N_2078);
nand U2117 (N_2117,N_2069,N_2068);
or U2118 (N_2118,N_2052,N_2064);
nand U2119 (N_2119,N_2066,N_2096);
nand U2120 (N_2120,N_2059,N_2062);
and U2121 (N_2121,N_2083,N_2050);
nor U2122 (N_2122,N_2084,N_2082);
xor U2123 (N_2123,N_2094,N_2056);
nor U2124 (N_2124,N_2085,N_2090);
and U2125 (N_2125,N_2068,N_2092);
and U2126 (N_2126,N_2070,N_2071);
nand U2127 (N_2127,N_2099,N_2055);
nand U2128 (N_2128,N_2059,N_2065);
or U2129 (N_2129,N_2085,N_2067);
or U2130 (N_2130,N_2082,N_2079);
xor U2131 (N_2131,N_2089,N_2059);
nor U2132 (N_2132,N_2061,N_2079);
nor U2133 (N_2133,N_2072,N_2095);
xor U2134 (N_2134,N_2091,N_2061);
or U2135 (N_2135,N_2077,N_2053);
and U2136 (N_2136,N_2097,N_2075);
and U2137 (N_2137,N_2054,N_2073);
and U2138 (N_2138,N_2077,N_2086);
nor U2139 (N_2139,N_2086,N_2060);
xnor U2140 (N_2140,N_2061,N_2064);
xnor U2141 (N_2141,N_2091,N_2062);
nand U2142 (N_2142,N_2086,N_2093);
or U2143 (N_2143,N_2078,N_2064);
and U2144 (N_2144,N_2090,N_2071);
xor U2145 (N_2145,N_2085,N_2053);
nand U2146 (N_2146,N_2058,N_2097);
xor U2147 (N_2147,N_2069,N_2062);
nand U2148 (N_2148,N_2068,N_2083);
and U2149 (N_2149,N_2079,N_2062);
nand U2150 (N_2150,N_2134,N_2131);
and U2151 (N_2151,N_2141,N_2146);
nor U2152 (N_2152,N_2118,N_2102);
nor U2153 (N_2153,N_2137,N_2100);
or U2154 (N_2154,N_2140,N_2109);
xnor U2155 (N_2155,N_2135,N_2120);
or U2156 (N_2156,N_2123,N_2121);
nand U2157 (N_2157,N_2117,N_2130);
or U2158 (N_2158,N_2113,N_2139);
xnor U2159 (N_2159,N_2126,N_2144);
or U2160 (N_2160,N_2129,N_2116);
and U2161 (N_2161,N_2125,N_2115);
nand U2162 (N_2162,N_2149,N_2127);
xor U2163 (N_2163,N_2145,N_2114);
and U2164 (N_2164,N_2138,N_2104);
xor U2165 (N_2165,N_2107,N_2101);
nor U2166 (N_2166,N_2105,N_2112);
xor U2167 (N_2167,N_2122,N_2132);
or U2168 (N_2168,N_2124,N_2106);
nand U2169 (N_2169,N_2128,N_2142);
nor U2170 (N_2170,N_2110,N_2136);
nor U2171 (N_2171,N_2111,N_2103);
and U2172 (N_2172,N_2143,N_2148);
xnor U2173 (N_2173,N_2108,N_2119);
nor U2174 (N_2174,N_2147,N_2133);
xor U2175 (N_2175,N_2144,N_2139);
xnor U2176 (N_2176,N_2122,N_2115);
and U2177 (N_2177,N_2133,N_2135);
xor U2178 (N_2178,N_2114,N_2132);
or U2179 (N_2179,N_2147,N_2132);
nor U2180 (N_2180,N_2133,N_2145);
and U2181 (N_2181,N_2140,N_2139);
xor U2182 (N_2182,N_2148,N_2116);
or U2183 (N_2183,N_2103,N_2107);
xor U2184 (N_2184,N_2136,N_2141);
and U2185 (N_2185,N_2118,N_2135);
nand U2186 (N_2186,N_2111,N_2139);
and U2187 (N_2187,N_2124,N_2145);
nor U2188 (N_2188,N_2100,N_2125);
xnor U2189 (N_2189,N_2129,N_2112);
nor U2190 (N_2190,N_2101,N_2148);
xor U2191 (N_2191,N_2130,N_2139);
xnor U2192 (N_2192,N_2148,N_2117);
xor U2193 (N_2193,N_2109,N_2110);
and U2194 (N_2194,N_2117,N_2143);
xor U2195 (N_2195,N_2109,N_2119);
and U2196 (N_2196,N_2123,N_2127);
nor U2197 (N_2197,N_2100,N_2131);
or U2198 (N_2198,N_2140,N_2145);
nor U2199 (N_2199,N_2100,N_2149);
xor U2200 (N_2200,N_2188,N_2167);
or U2201 (N_2201,N_2160,N_2186);
nand U2202 (N_2202,N_2197,N_2159);
nand U2203 (N_2203,N_2196,N_2182);
xnor U2204 (N_2204,N_2175,N_2179);
and U2205 (N_2205,N_2195,N_2185);
or U2206 (N_2206,N_2183,N_2194);
or U2207 (N_2207,N_2199,N_2169);
nor U2208 (N_2208,N_2154,N_2192);
nor U2209 (N_2209,N_2178,N_2176);
nor U2210 (N_2210,N_2180,N_2158);
nand U2211 (N_2211,N_2171,N_2153);
nor U2212 (N_2212,N_2155,N_2198);
nor U2213 (N_2213,N_2156,N_2177);
nand U2214 (N_2214,N_2184,N_2170);
or U2215 (N_2215,N_2157,N_2152);
xor U2216 (N_2216,N_2165,N_2173);
nand U2217 (N_2217,N_2174,N_2181);
and U2218 (N_2218,N_2151,N_2162);
and U2219 (N_2219,N_2168,N_2172);
nor U2220 (N_2220,N_2189,N_2187);
nor U2221 (N_2221,N_2150,N_2191);
or U2222 (N_2222,N_2161,N_2193);
xnor U2223 (N_2223,N_2164,N_2190);
nor U2224 (N_2224,N_2163,N_2166);
nand U2225 (N_2225,N_2154,N_2166);
or U2226 (N_2226,N_2180,N_2182);
or U2227 (N_2227,N_2153,N_2158);
and U2228 (N_2228,N_2179,N_2176);
and U2229 (N_2229,N_2184,N_2189);
nand U2230 (N_2230,N_2187,N_2177);
or U2231 (N_2231,N_2189,N_2164);
or U2232 (N_2232,N_2176,N_2150);
nand U2233 (N_2233,N_2151,N_2188);
xor U2234 (N_2234,N_2150,N_2186);
and U2235 (N_2235,N_2171,N_2197);
nand U2236 (N_2236,N_2150,N_2163);
nor U2237 (N_2237,N_2160,N_2176);
or U2238 (N_2238,N_2175,N_2190);
xnor U2239 (N_2239,N_2172,N_2153);
and U2240 (N_2240,N_2162,N_2190);
xor U2241 (N_2241,N_2180,N_2193);
or U2242 (N_2242,N_2158,N_2187);
nor U2243 (N_2243,N_2194,N_2197);
and U2244 (N_2244,N_2194,N_2195);
xor U2245 (N_2245,N_2183,N_2168);
xnor U2246 (N_2246,N_2155,N_2182);
or U2247 (N_2247,N_2186,N_2154);
or U2248 (N_2248,N_2171,N_2181);
and U2249 (N_2249,N_2185,N_2165);
and U2250 (N_2250,N_2205,N_2240);
and U2251 (N_2251,N_2203,N_2206);
xnor U2252 (N_2252,N_2226,N_2204);
xor U2253 (N_2253,N_2228,N_2210);
xnor U2254 (N_2254,N_2233,N_2201);
or U2255 (N_2255,N_2237,N_2220);
xor U2256 (N_2256,N_2217,N_2238);
xor U2257 (N_2257,N_2249,N_2239);
xor U2258 (N_2258,N_2216,N_2219);
xor U2259 (N_2259,N_2246,N_2208);
nor U2260 (N_2260,N_2213,N_2229);
or U2261 (N_2261,N_2242,N_2248);
or U2262 (N_2262,N_2214,N_2243);
nand U2263 (N_2263,N_2245,N_2211);
xnor U2264 (N_2264,N_2224,N_2218);
xor U2265 (N_2265,N_2227,N_2207);
nand U2266 (N_2266,N_2232,N_2231);
xnor U2267 (N_2267,N_2241,N_2236);
nand U2268 (N_2268,N_2221,N_2222);
nand U2269 (N_2269,N_2200,N_2215);
nor U2270 (N_2270,N_2234,N_2212);
xnor U2271 (N_2271,N_2225,N_2209);
xor U2272 (N_2272,N_2244,N_2230);
or U2273 (N_2273,N_2223,N_2247);
xor U2274 (N_2274,N_2202,N_2235);
and U2275 (N_2275,N_2244,N_2207);
and U2276 (N_2276,N_2240,N_2244);
nor U2277 (N_2277,N_2212,N_2200);
xor U2278 (N_2278,N_2201,N_2212);
or U2279 (N_2279,N_2205,N_2216);
or U2280 (N_2280,N_2209,N_2226);
and U2281 (N_2281,N_2233,N_2228);
and U2282 (N_2282,N_2207,N_2208);
or U2283 (N_2283,N_2232,N_2248);
nand U2284 (N_2284,N_2242,N_2239);
xnor U2285 (N_2285,N_2243,N_2221);
nand U2286 (N_2286,N_2211,N_2242);
xnor U2287 (N_2287,N_2216,N_2234);
or U2288 (N_2288,N_2226,N_2238);
xor U2289 (N_2289,N_2235,N_2212);
or U2290 (N_2290,N_2239,N_2240);
xor U2291 (N_2291,N_2242,N_2216);
or U2292 (N_2292,N_2206,N_2244);
xor U2293 (N_2293,N_2230,N_2219);
nand U2294 (N_2294,N_2236,N_2223);
xor U2295 (N_2295,N_2229,N_2215);
nor U2296 (N_2296,N_2222,N_2230);
nor U2297 (N_2297,N_2221,N_2204);
nor U2298 (N_2298,N_2229,N_2245);
or U2299 (N_2299,N_2231,N_2234);
nor U2300 (N_2300,N_2270,N_2269);
xor U2301 (N_2301,N_2254,N_2260);
xor U2302 (N_2302,N_2288,N_2251);
nor U2303 (N_2303,N_2298,N_2273);
nand U2304 (N_2304,N_2255,N_2265);
or U2305 (N_2305,N_2295,N_2293);
nor U2306 (N_2306,N_2287,N_2271);
xor U2307 (N_2307,N_2258,N_2268);
nand U2308 (N_2308,N_2284,N_2257);
or U2309 (N_2309,N_2252,N_2296);
or U2310 (N_2310,N_2275,N_2256);
nor U2311 (N_2311,N_2274,N_2263);
nand U2312 (N_2312,N_2282,N_2292);
and U2313 (N_2313,N_2262,N_2290);
and U2314 (N_2314,N_2285,N_2281);
nor U2315 (N_2315,N_2276,N_2286);
nor U2316 (N_2316,N_2259,N_2277);
and U2317 (N_2317,N_2261,N_2278);
xor U2318 (N_2318,N_2297,N_2294);
or U2319 (N_2319,N_2267,N_2291);
nand U2320 (N_2320,N_2272,N_2289);
or U2321 (N_2321,N_2299,N_2280);
and U2322 (N_2322,N_2283,N_2266);
xor U2323 (N_2323,N_2253,N_2250);
nor U2324 (N_2324,N_2279,N_2264);
nand U2325 (N_2325,N_2298,N_2287);
nor U2326 (N_2326,N_2267,N_2266);
or U2327 (N_2327,N_2299,N_2254);
xnor U2328 (N_2328,N_2270,N_2261);
nor U2329 (N_2329,N_2262,N_2292);
nand U2330 (N_2330,N_2271,N_2256);
and U2331 (N_2331,N_2280,N_2274);
nand U2332 (N_2332,N_2284,N_2251);
and U2333 (N_2333,N_2256,N_2288);
nor U2334 (N_2334,N_2284,N_2277);
nor U2335 (N_2335,N_2262,N_2288);
or U2336 (N_2336,N_2276,N_2281);
or U2337 (N_2337,N_2259,N_2250);
or U2338 (N_2338,N_2258,N_2278);
or U2339 (N_2339,N_2286,N_2265);
or U2340 (N_2340,N_2297,N_2266);
nor U2341 (N_2341,N_2297,N_2271);
nand U2342 (N_2342,N_2259,N_2264);
or U2343 (N_2343,N_2262,N_2255);
nand U2344 (N_2344,N_2284,N_2287);
nor U2345 (N_2345,N_2292,N_2260);
nor U2346 (N_2346,N_2292,N_2275);
nor U2347 (N_2347,N_2289,N_2285);
xor U2348 (N_2348,N_2255,N_2251);
xnor U2349 (N_2349,N_2268,N_2291);
nor U2350 (N_2350,N_2332,N_2323);
and U2351 (N_2351,N_2326,N_2345);
nor U2352 (N_2352,N_2311,N_2308);
nand U2353 (N_2353,N_2331,N_2337);
nand U2354 (N_2354,N_2307,N_2320);
nor U2355 (N_2355,N_2306,N_2341);
xor U2356 (N_2356,N_2338,N_2333);
and U2357 (N_2357,N_2328,N_2340);
nand U2358 (N_2358,N_2330,N_2304);
nor U2359 (N_2359,N_2339,N_2313);
nor U2360 (N_2360,N_2301,N_2334);
and U2361 (N_2361,N_2315,N_2336);
nor U2362 (N_2362,N_2342,N_2344);
nor U2363 (N_2363,N_2329,N_2312);
nand U2364 (N_2364,N_2302,N_2325);
nor U2365 (N_2365,N_2314,N_2316);
nand U2366 (N_2366,N_2343,N_2305);
nor U2367 (N_2367,N_2335,N_2327);
xnor U2368 (N_2368,N_2321,N_2309);
and U2369 (N_2369,N_2319,N_2310);
nand U2370 (N_2370,N_2303,N_2324);
nor U2371 (N_2371,N_2348,N_2322);
xor U2372 (N_2372,N_2300,N_2346);
and U2373 (N_2373,N_2318,N_2317);
or U2374 (N_2374,N_2347,N_2349);
and U2375 (N_2375,N_2336,N_2344);
nand U2376 (N_2376,N_2325,N_2304);
and U2377 (N_2377,N_2328,N_2338);
and U2378 (N_2378,N_2333,N_2342);
or U2379 (N_2379,N_2308,N_2346);
xnor U2380 (N_2380,N_2308,N_2335);
nor U2381 (N_2381,N_2331,N_2301);
nor U2382 (N_2382,N_2348,N_2314);
nand U2383 (N_2383,N_2342,N_2312);
xor U2384 (N_2384,N_2340,N_2345);
xor U2385 (N_2385,N_2332,N_2316);
nor U2386 (N_2386,N_2307,N_2339);
nand U2387 (N_2387,N_2303,N_2332);
and U2388 (N_2388,N_2315,N_2301);
and U2389 (N_2389,N_2320,N_2334);
nand U2390 (N_2390,N_2300,N_2319);
xnor U2391 (N_2391,N_2349,N_2322);
and U2392 (N_2392,N_2305,N_2302);
or U2393 (N_2393,N_2321,N_2334);
nand U2394 (N_2394,N_2339,N_2342);
or U2395 (N_2395,N_2338,N_2348);
xor U2396 (N_2396,N_2349,N_2345);
xnor U2397 (N_2397,N_2316,N_2307);
xnor U2398 (N_2398,N_2348,N_2336);
and U2399 (N_2399,N_2300,N_2337);
and U2400 (N_2400,N_2390,N_2355);
xnor U2401 (N_2401,N_2386,N_2398);
nor U2402 (N_2402,N_2366,N_2375);
xor U2403 (N_2403,N_2397,N_2367);
or U2404 (N_2404,N_2351,N_2363);
or U2405 (N_2405,N_2352,N_2357);
xnor U2406 (N_2406,N_2395,N_2396);
and U2407 (N_2407,N_2361,N_2371);
or U2408 (N_2408,N_2377,N_2394);
nand U2409 (N_2409,N_2381,N_2372);
and U2410 (N_2410,N_2391,N_2376);
xnor U2411 (N_2411,N_2393,N_2399);
nor U2412 (N_2412,N_2359,N_2385);
nor U2413 (N_2413,N_2392,N_2382);
nand U2414 (N_2414,N_2360,N_2373);
and U2415 (N_2415,N_2353,N_2365);
nand U2416 (N_2416,N_2378,N_2380);
and U2417 (N_2417,N_2356,N_2369);
or U2418 (N_2418,N_2368,N_2358);
nor U2419 (N_2419,N_2383,N_2379);
or U2420 (N_2420,N_2374,N_2389);
nor U2421 (N_2421,N_2354,N_2364);
or U2422 (N_2422,N_2370,N_2384);
nor U2423 (N_2423,N_2388,N_2387);
or U2424 (N_2424,N_2362,N_2350);
and U2425 (N_2425,N_2388,N_2381);
xor U2426 (N_2426,N_2387,N_2381);
or U2427 (N_2427,N_2359,N_2391);
xor U2428 (N_2428,N_2382,N_2352);
nand U2429 (N_2429,N_2370,N_2399);
nor U2430 (N_2430,N_2386,N_2368);
and U2431 (N_2431,N_2372,N_2355);
and U2432 (N_2432,N_2360,N_2387);
xnor U2433 (N_2433,N_2398,N_2353);
and U2434 (N_2434,N_2392,N_2385);
nand U2435 (N_2435,N_2387,N_2366);
or U2436 (N_2436,N_2350,N_2364);
nand U2437 (N_2437,N_2382,N_2381);
nand U2438 (N_2438,N_2361,N_2382);
nand U2439 (N_2439,N_2378,N_2387);
xnor U2440 (N_2440,N_2399,N_2390);
nor U2441 (N_2441,N_2397,N_2359);
nand U2442 (N_2442,N_2378,N_2363);
or U2443 (N_2443,N_2385,N_2398);
and U2444 (N_2444,N_2375,N_2352);
xor U2445 (N_2445,N_2356,N_2376);
nor U2446 (N_2446,N_2377,N_2393);
and U2447 (N_2447,N_2377,N_2378);
nor U2448 (N_2448,N_2385,N_2354);
or U2449 (N_2449,N_2355,N_2359);
nand U2450 (N_2450,N_2435,N_2411);
nor U2451 (N_2451,N_2404,N_2414);
or U2452 (N_2452,N_2442,N_2418);
nor U2453 (N_2453,N_2432,N_2410);
or U2454 (N_2454,N_2447,N_2402);
nor U2455 (N_2455,N_2401,N_2416);
nor U2456 (N_2456,N_2425,N_2406);
or U2457 (N_2457,N_2429,N_2422);
nor U2458 (N_2458,N_2400,N_2420);
and U2459 (N_2459,N_2415,N_2412);
or U2460 (N_2460,N_2436,N_2444);
xnor U2461 (N_2461,N_2424,N_2441);
and U2462 (N_2462,N_2409,N_2434);
or U2463 (N_2463,N_2413,N_2439);
nor U2464 (N_2464,N_2430,N_2408);
nand U2465 (N_2465,N_2438,N_2437);
and U2466 (N_2466,N_2443,N_2433);
xor U2467 (N_2467,N_2440,N_2431);
nor U2468 (N_2468,N_2421,N_2405);
nor U2469 (N_2469,N_2449,N_2419);
or U2470 (N_2470,N_2448,N_2423);
xnor U2471 (N_2471,N_2417,N_2426);
nor U2472 (N_2472,N_2403,N_2445);
nor U2473 (N_2473,N_2428,N_2427);
and U2474 (N_2474,N_2446,N_2407);
xor U2475 (N_2475,N_2437,N_2409);
or U2476 (N_2476,N_2430,N_2437);
xnor U2477 (N_2477,N_2428,N_2435);
xnor U2478 (N_2478,N_2421,N_2446);
nor U2479 (N_2479,N_2410,N_2404);
nand U2480 (N_2480,N_2417,N_2416);
xnor U2481 (N_2481,N_2444,N_2433);
xor U2482 (N_2482,N_2432,N_2417);
and U2483 (N_2483,N_2419,N_2427);
or U2484 (N_2484,N_2440,N_2407);
nor U2485 (N_2485,N_2400,N_2440);
or U2486 (N_2486,N_2437,N_2420);
nor U2487 (N_2487,N_2403,N_2435);
xnor U2488 (N_2488,N_2426,N_2424);
nand U2489 (N_2489,N_2434,N_2428);
or U2490 (N_2490,N_2402,N_2434);
and U2491 (N_2491,N_2403,N_2430);
and U2492 (N_2492,N_2431,N_2444);
nor U2493 (N_2493,N_2424,N_2433);
nand U2494 (N_2494,N_2415,N_2409);
or U2495 (N_2495,N_2431,N_2426);
and U2496 (N_2496,N_2444,N_2414);
or U2497 (N_2497,N_2406,N_2434);
xnor U2498 (N_2498,N_2449,N_2403);
or U2499 (N_2499,N_2445,N_2434);
nor U2500 (N_2500,N_2497,N_2457);
or U2501 (N_2501,N_2492,N_2478);
xnor U2502 (N_2502,N_2488,N_2468);
and U2503 (N_2503,N_2477,N_2473);
or U2504 (N_2504,N_2481,N_2465);
nor U2505 (N_2505,N_2487,N_2451);
xor U2506 (N_2506,N_2460,N_2459);
and U2507 (N_2507,N_2479,N_2476);
nand U2508 (N_2508,N_2455,N_2496);
and U2509 (N_2509,N_2470,N_2498);
nor U2510 (N_2510,N_2483,N_2464);
and U2511 (N_2511,N_2461,N_2485);
nor U2512 (N_2512,N_2489,N_2466);
xor U2513 (N_2513,N_2475,N_2458);
nand U2514 (N_2514,N_2486,N_2450);
nor U2515 (N_2515,N_2472,N_2499);
or U2516 (N_2516,N_2467,N_2491);
and U2517 (N_2517,N_2480,N_2453);
nor U2518 (N_2518,N_2452,N_2469);
xor U2519 (N_2519,N_2462,N_2463);
or U2520 (N_2520,N_2482,N_2474);
and U2521 (N_2521,N_2493,N_2456);
nand U2522 (N_2522,N_2484,N_2495);
and U2523 (N_2523,N_2494,N_2471);
or U2524 (N_2524,N_2490,N_2454);
nand U2525 (N_2525,N_2474,N_2450);
nand U2526 (N_2526,N_2480,N_2488);
and U2527 (N_2527,N_2495,N_2490);
nand U2528 (N_2528,N_2468,N_2485);
and U2529 (N_2529,N_2490,N_2480);
xnor U2530 (N_2530,N_2458,N_2495);
or U2531 (N_2531,N_2472,N_2495);
nand U2532 (N_2532,N_2472,N_2496);
nand U2533 (N_2533,N_2478,N_2472);
nand U2534 (N_2534,N_2480,N_2461);
xnor U2535 (N_2535,N_2470,N_2469);
nand U2536 (N_2536,N_2481,N_2478);
or U2537 (N_2537,N_2499,N_2467);
xor U2538 (N_2538,N_2465,N_2492);
nor U2539 (N_2539,N_2474,N_2498);
xnor U2540 (N_2540,N_2469,N_2462);
xnor U2541 (N_2541,N_2489,N_2459);
nand U2542 (N_2542,N_2467,N_2497);
nand U2543 (N_2543,N_2459,N_2496);
or U2544 (N_2544,N_2494,N_2474);
nand U2545 (N_2545,N_2452,N_2459);
nor U2546 (N_2546,N_2462,N_2468);
nor U2547 (N_2547,N_2487,N_2490);
nand U2548 (N_2548,N_2459,N_2492);
or U2549 (N_2549,N_2455,N_2490);
and U2550 (N_2550,N_2525,N_2514);
and U2551 (N_2551,N_2509,N_2549);
and U2552 (N_2552,N_2540,N_2532);
xor U2553 (N_2553,N_2542,N_2505);
nand U2554 (N_2554,N_2512,N_2543);
nor U2555 (N_2555,N_2526,N_2506);
and U2556 (N_2556,N_2528,N_2518);
and U2557 (N_2557,N_2502,N_2517);
or U2558 (N_2558,N_2508,N_2511);
or U2559 (N_2559,N_2521,N_2527);
nor U2560 (N_2560,N_2546,N_2544);
xnor U2561 (N_2561,N_2524,N_2538);
and U2562 (N_2562,N_2513,N_2536);
nor U2563 (N_2563,N_2522,N_2523);
nor U2564 (N_2564,N_2504,N_2501);
or U2565 (N_2565,N_2520,N_2530);
nor U2566 (N_2566,N_2500,N_2535);
nor U2567 (N_2567,N_2545,N_2519);
and U2568 (N_2568,N_2548,N_2547);
and U2569 (N_2569,N_2539,N_2503);
or U2570 (N_2570,N_2537,N_2534);
xor U2571 (N_2571,N_2510,N_2515);
or U2572 (N_2572,N_2533,N_2529);
nand U2573 (N_2573,N_2531,N_2507);
nor U2574 (N_2574,N_2516,N_2541);
xor U2575 (N_2575,N_2545,N_2501);
xnor U2576 (N_2576,N_2507,N_2524);
or U2577 (N_2577,N_2516,N_2535);
nand U2578 (N_2578,N_2531,N_2530);
xnor U2579 (N_2579,N_2515,N_2514);
nor U2580 (N_2580,N_2528,N_2531);
or U2581 (N_2581,N_2549,N_2510);
xnor U2582 (N_2582,N_2540,N_2502);
nand U2583 (N_2583,N_2519,N_2510);
nand U2584 (N_2584,N_2507,N_2516);
and U2585 (N_2585,N_2521,N_2516);
xor U2586 (N_2586,N_2532,N_2518);
xnor U2587 (N_2587,N_2549,N_2543);
nand U2588 (N_2588,N_2546,N_2511);
and U2589 (N_2589,N_2502,N_2549);
nand U2590 (N_2590,N_2517,N_2523);
or U2591 (N_2591,N_2517,N_2547);
xor U2592 (N_2592,N_2531,N_2538);
nor U2593 (N_2593,N_2532,N_2527);
xor U2594 (N_2594,N_2534,N_2513);
xnor U2595 (N_2595,N_2529,N_2500);
xnor U2596 (N_2596,N_2502,N_2542);
nor U2597 (N_2597,N_2527,N_2526);
or U2598 (N_2598,N_2514,N_2519);
xor U2599 (N_2599,N_2523,N_2504);
and U2600 (N_2600,N_2581,N_2599);
nand U2601 (N_2601,N_2563,N_2576);
nand U2602 (N_2602,N_2556,N_2596);
nand U2603 (N_2603,N_2590,N_2550);
xor U2604 (N_2604,N_2594,N_2572);
or U2605 (N_2605,N_2568,N_2559);
nor U2606 (N_2606,N_2570,N_2565);
and U2607 (N_2607,N_2573,N_2589);
nor U2608 (N_2608,N_2579,N_2561);
nor U2609 (N_2609,N_2562,N_2582);
xnor U2610 (N_2610,N_2558,N_2587);
nor U2611 (N_2611,N_2592,N_2567);
nand U2612 (N_2612,N_2571,N_2598);
or U2613 (N_2613,N_2580,N_2553);
xor U2614 (N_2614,N_2552,N_2595);
or U2615 (N_2615,N_2583,N_2585);
and U2616 (N_2616,N_2597,N_2578);
nand U2617 (N_2617,N_2564,N_2560);
or U2618 (N_2618,N_2555,N_2569);
or U2619 (N_2619,N_2566,N_2586);
xor U2620 (N_2620,N_2584,N_2575);
xor U2621 (N_2621,N_2588,N_2551);
and U2622 (N_2622,N_2574,N_2591);
or U2623 (N_2623,N_2557,N_2554);
nor U2624 (N_2624,N_2577,N_2593);
xor U2625 (N_2625,N_2554,N_2591);
nor U2626 (N_2626,N_2583,N_2581);
or U2627 (N_2627,N_2597,N_2595);
xnor U2628 (N_2628,N_2593,N_2569);
xor U2629 (N_2629,N_2582,N_2563);
and U2630 (N_2630,N_2550,N_2553);
or U2631 (N_2631,N_2567,N_2579);
xnor U2632 (N_2632,N_2578,N_2558);
or U2633 (N_2633,N_2563,N_2583);
nand U2634 (N_2634,N_2562,N_2566);
xor U2635 (N_2635,N_2587,N_2571);
and U2636 (N_2636,N_2577,N_2595);
xor U2637 (N_2637,N_2597,N_2550);
or U2638 (N_2638,N_2553,N_2573);
nand U2639 (N_2639,N_2570,N_2571);
nor U2640 (N_2640,N_2561,N_2556);
and U2641 (N_2641,N_2586,N_2551);
nor U2642 (N_2642,N_2577,N_2554);
nor U2643 (N_2643,N_2588,N_2594);
xor U2644 (N_2644,N_2573,N_2563);
or U2645 (N_2645,N_2595,N_2580);
nand U2646 (N_2646,N_2579,N_2569);
and U2647 (N_2647,N_2563,N_2597);
nand U2648 (N_2648,N_2560,N_2570);
xnor U2649 (N_2649,N_2577,N_2570);
and U2650 (N_2650,N_2634,N_2621);
xnor U2651 (N_2651,N_2600,N_2626);
and U2652 (N_2652,N_2613,N_2615);
nand U2653 (N_2653,N_2644,N_2605);
nor U2654 (N_2654,N_2633,N_2627);
and U2655 (N_2655,N_2628,N_2620);
or U2656 (N_2656,N_2622,N_2645);
nor U2657 (N_2657,N_2614,N_2639);
or U2658 (N_2658,N_2643,N_2625);
and U2659 (N_2659,N_2648,N_2630);
and U2660 (N_2660,N_2611,N_2631);
xor U2661 (N_2661,N_2608,N_2623);
nand U2662 (N_2662,N_2601,N_2604);
xnor U2663 (N_2663,N_2636,N_2629);
nor U2664 (N_2664,N_2603,N_2640);
and U2665 (N_2665,N_2624,N_2619);
or U2666 (N_2666,N_2606,N_2638);
nor U2667 (N_2667,N_2618,N_2609);
xor U2668 (N_2668,N_2632,N_2647);
xor U2669 (N_2669,N_2635,N_2612);
or U2670 (N_2670,N_2637,N_2642);
xnor U2671 (N_2671,N_2610,N_2646);
or U2672 (N_2672,N_2641,N_2616);
or U2673 (N_2673,N_2607,N_2649);
nor U2674 (N_2674,N_2602,N_2617);
nor U2675 (N_2675,N_2615,N_2622);
and U2676 (N_2676,N_2631,N_2610);
and U2677 (N_2677,N_2647,N_2602);
xor U2678 (N_2678,N_2618,N_2631);
and U2679 (N_2679,N_2625,N_2612);
or U2680 (N_2680,N_2628,N_2623);
or U2681 (N_2681,N_2615,N_2638);
xnor U2682 (N_2682,N_2611,N_2612);
nor U2683 (N_2683,N_2619,N_2602);
or U2684 (N_2684,N_2628,N_2617);
nor U2685 (N_2685,N_2627,N_2625);
and U2686 (N_2686,N_2640,N_2645);
nor U2687 (N_2687,N_2600,N_2614);
nor U2688 (N_2688,N_2649,N_2644);
and U2689 (N_2689,N_2616,N_2632);
and U2690 (N_2690,N_2643,N_2604);
xor U2691 (N_2691,N_2615,N_2643);
xor U2692 (N_2692,N_2618,N_2605);
nor U2693 (N_2693,N_2640,N_2604);
or U2694 (N_2694,N_2648,N_2649);
nand U2695 (N_2695,N_2623,N_2638);
nor U2696 (N_2696,N_2617,N_2609);
nand U2697 (N_2697,N_2611,N_2648);
xor U2698 (N_2698,N_2636,N_2602);
nand U2699 (N_2699,N_2634,N_2605);
and U2700 (N_2700,N_2679,N_2692);
and U2701 (N_2701,N_2691,N_2681);
nand U2702 (N_2702,N_2658,N_2680);
or U2703 (N_2703,N_2674,N_2678);
or U2704 (N_2704,N_2694,N_2677);
nand U2705 (N_2705,N_2651,N_2667);
nor U2706 (N_2706,N_2661,N_2682);
xor U2707 (N_2707,N_2695,N_2662);
nor U2708 (N_2708,N_2656,N_2676);
xor U2709 (N_2709,N_2650,N_2697);
nand U2710 (N_2710,N_2660,N_2670);
xnor U2711 (N_2711,N_2687,N_2665);
or U2712 (N_2712,N_2653,N_2689);
nand U2713 (N_2713,N_2671,N_2699);
nand U2714 (N_2714,N_2672,N_2686);
nand U2715 (N_2715,N_2663,N_2654);
nand U2716 (N_2716,N_2688,N_2657);
nor U2717 (N_2717,N_2652,N_2693);
or U2718 (N_2718,N_2675,N_2685);
or U2719 (N_2719,N_2690,N_2669);
xnor U2720 (N_2720,N_2666,N_2664);
nand U2721 (N_2721,N_2655,N_2673);
xnor U2722 (N_2722,N_2683,N_2684);
xor U2723 (N_2723,N_2668,N_2696);
nor U2724 (N_2724,N_2698,N_2659);
xnor U2725 (N_2725,N_2682,N_2662);
or U2726 (N_2726,N_2655,N_2658);
or U2727 (N_2727,N_2662,N_2680);
nand U2728 (N_2728,N_2699,N_2660);
nor U2729 (N_2729,N_2652,N_2697);
and U2730 (N_2730,N_2689,N_2662);
nor U2731 (N_2731,N_2661,N_2694);
nand U2732 (N_2732,N_2660,N_2654);
nand U2733 (N_2733,N_2695,N_2653);
nand U2734 (N_2734,N_2671,N_2665);
nor U2735 (N_2735,N_2690,N_2676);
nand U2736 (N_2736,N_2688,N_2660);
and U2737 (N_2737,N_2693,N_2684);
or U2738 (N_2738,N_2677,N_2664);
and U2739 (N_2739,N_2650,N_2656);
or U2740 (N_2740,N_2687,N_2667);
or U2741 (N_2741,N_2689,N_2655);
nor U2742 (N_2742,N_2680,N_2678);
xnor U2743 (N_2743,N_2694,N_2688);
or U2744 (N_2744,N_2657,N_2696);
nand U2745 (N_2745,N_2657,N_2654);
nor U2746 (N_2746,N_2696,N_2652);
xnor U2747 (N_2747,N_2673,N_2680);
nand U2748 (N_2748,N_2676,N_2651);
xnor U2749 (N_2749,N_2694,N_2696);
xnor U2750 (N_2750,N_2739,N_2729);
and U2751 (N_2751,N_2748,N_2738);
and U2752 (N_2752,N_2718,N_2720);
xor U2753 (N_2753,N_2703,N_2712);
nor U2754 (N_2754,N_2743,N_2741);
or U2755 (N_2755,N_2745,N_2746);
xor U2756 (N_2756,N_2731,N_2747);
or U2757 (N_2757,N_2709,N_2735);
nor U2758 (N_2758,N_2730,N_2706);
nand U2759 (N_2759,N_2732,N_2726);
xor U2760 (N_2760,N_2713,N_2724);
or U2761 (N_2761,N_2711,N_2704);
or U2762 (N_2762,N_2727,N_2702);
and U2763 (N_2763,N_2723,N_2719);
and U2764 (N_2764,N_2700,N_2722);
nor U2765 (N_2765,N_2725,N_2749);
nand U2766 (N_2766,N_2708,N_2734);
or U2767 (N_2767,N_2716,N_2721);
nor U2768 (N_2768,N_2733,N_2710);
xor U2769 (N_2769,N_2707,N_2715);
or U2770 (N_2770,N_2744,N_2736);
xnor U2771 (N_2771,N_2701,N_2742);
nand U2772 (N_2772,N_2728,N_2714);
and U2773 (N_2773,N_2737,N_2705);
nor U2774 (N_2774,N_2740,N_2717);
xor U2775 (N_2775,N_2715,N_2702);
xnor U2776 (N_2776,N_2737,N_2710);
or U2777 (N_2777,N_2743,N_2736);
xor U2778 (N_2778,N_2709,N_2733);
nand U2779 (N_2779,N_2736,N_2710);
nand U2780 (N_2780,N_2742,N_2746);
nand U2781 (N_2781,N_2727,N_2747);
xnor U2782 (N_2782,N_2725,N_2714);
xor U2783 (N_2783,N_2741,N_2711);
xnor U2784 (N_2784,N_2748,N_2703);
and U2785 (N_2785,N_2702,N_2738);
xnor U2786 (N_2786,N_2727,N_2742);
nand U2787 (N_2787,N_2744,N_2741);
nand U2788 (N_2788,N_2732,N_2718);
xnor U2789 (N_2789,N_2738,N_2716);
nand U2790 (N_2790,N_2726,N_2740);
or U2791 (N_2791,N_2730,N_2746);
xor U2792 (N_2792,N_2723,N_2727);
nor U2793 (N_2793,N_2702,N_2737);
xor U2794 (N_2794,N_2719,N_2712);
or U2795 (N_2795,N_2719,N_2738);
and U2796 (N_2796,N_2709,N_2700);
or U2797 (N_2797,N_2737,N_2715);
or U2798 (N_2798,N_2719,N_2740);
and U2799 (N_2799,N_2719,N_2705);
or U2800 (N_2800,N_2769,N_2766);
or U2801 (N_2801,N_2772,N_2798);
and U2802 (N_2802,N_2760,N_2768);
nor U2803 (N_2803,N_2771,N_2751);
xor U2804 (N_2804,N_2762,N_2759);
xnor U2805 (N_2805,N_2757,N_2750);
nand U2806 (N_2806,N_2775,N_2786);
nor U2807 (N_2807,N_2752,N_2784);
and U2808 (N_2808,N_2774,N_2793);
and U2809 (N_2809,N_2767,N_2797);
nand U2810 (N_2810,N_2770,N_2778);
and U2811 (N_2811,N_2783,N_2794);
and U2812 (N_2812,N_2792,N_2779);
xor U2813 (N_2813,N_2788,N_2763);
xnor U2814 (N_2814,N_2755,N_2753);
or U2815 (N_2815,N_2789,N_2777);
nand U2816 (N_2816,N_2796,N_2758);
nor U2817 (N_2817,N_2787,N_2754);
nor U2818 (N_2818,N_2782,N_2785);
nor U2819 (N_2819,N_2756,N_2791);
xor U2820 (N_2820,N_2780,N_2765);
or U2821 (N_2821,N_2799,N_2781);
and U2822 (N_2822,N_2776,N_2773);
and U2823 (N_2823,N_2795,N_2790);
nor U2824 (N_2824,N_2764,N_2761);
xnor U2825 (N_2825,N_2772,N_2756);
or U2826 (N_2826,N_2754,N_2768);
nor U2827 (N_2827,N_2776,N_2787);
nor U2828 (N_2828,N_2785,N_2770);
and U2829 (N_2829,N_2756,N_2777);
xnor U2830 (N_2830,N_2788,N_2774);
and U2831 (N_2831,N_2792,N_2778);
xnor U2832 (N_2832,N_2794,N_2776);
nand U2833 (N_2833,N_2750,N_2798);
nand U2834 (N_2834,N_2760,N_2754);
and U2835 (N_2835,N_2776,N_2795);
nor U2836 (N_2836,N_2754,N_2795);
nand U2837 (N_2837,N_2786,N_2777);
or U2838 (N_2838,N_2768,N_2764);
or U2839 (N_2839,N_2792,N_2787);
xnor U2840 (N_2840,N_2769,N_2764);
xor U2841 (N_2841,N_2772,N_2789);
or U2842 (N_2842,N_2794,N_2750);
or U2843 (N_2843,N_2797,N_2786);
and U2844 (N_2844,N_2760,N_2766);
or U2845 (N_2845,N_2781,N_2798);
nand U2846 (N_2846,N_2751,N_2775);
nand U2847 (N_2847,N_2786,N_2791);
and U2848 (N_2848,N_2754,N_2755);
nand U2849 (N_2849,N_2774,N_2779);
xor U2850 (N_2850,N_2842,N_2832);
nand U2851 (N_2851,N_2824,N_2804);
nand U2852 (N_2852,N_2800,N_2814);
nor U2853 (N_2853,N_2802,N_2835);
nand U2854 (N_2854,N_2806,N_2840);
and U2855 (N_2855,N_2803,N_2833);
nand U2856 (N_2856,N_2834,N_2817);
or U2857 (N_2857,N_2809,N_2807);
xnor U2858 (N_2858,N_2845,N_2811);
nor U2859 (N_2859,N_2808,N_2820);
nand U2860 (N_2860,N_2836,N_2813);
or U2861 (N_2861,N_2847,N_2827);
nand U2862 (N_2862,N_2829,N_2819);
and U2863 (N_2863,N_2805,N_2841);
nand U2864 (N_2864,N_2801,N_2822);
or U2865 (N_2865,N_2831,N_2826);
or U2866 (N_2866,N_2818,N_2812);
and U2867 (N_2867,N_2816,N_2823);
or U2868 (N_2868,N_2843,N_2828);
xnor U2869 (N_2869,N_2821,N_2825);
and U2870 (N_2870,N_2837,N_2849);
or U2871 (N_2871,N_2839,N_2846);
or U2872 (N_2872,N_2848,N_2830);
or U2873 (N_2873,N_2844,N_2838);
or U2874 (N_2874,N_2810,N_2815);
nor U2875 (N_2875,N_2804,N_2810);
nor U2876 (N_2876,N_2846,N_2819);
and U2877 (N_2877,N_2812,N_2800);
nand U2878 (N_2878,N_2822,N_2840);
or U2879 (N_2879,N_2809,N_2846);
nor U2880 (N_2880,N_2849,N_2828);
and U2881 (N_2881,N_2819,N_2806);
nand U2882 (N_2882,N_2807,N_2813);
xnor U2883 (N_2883,N_2824,N_2803);
or U2884 (N_2884,N_2834,N_2835);
nand U2885 (N_2885,N_2846,N_2811);
xnor U2886 (N_2886,N_2812,N_2814);
nor U2887 (N_2887,N_2814,N_2815);
and U2888 (N_2888,N_2830,N_2824);
or U2889 (N_2889,N_2811,N_2849);
nand U2890 (N_2890,N_2832,N_2808);
nor U2891 (N_2891,N_2835,N_2840);
nor U2892 (N_2892,N_2820,N_2834);
nor U2893 (N_2893,N_2805,N_2806);
nor U2894 (N_2894,N_2823,N_2812);
and U2895 (N_2895,N_2801,N_2828);
nor U2896 (N_2896,N_2828,N_2830);
xnor U2897 (N_2897,N_2830,N_2845);
and U2898 (N_2898,N_2838,N_2809);
nor U2899 (N_2899,N_2825,N_2828);
nor U2900 (N_2900,N_2858,N_2899);
nor U2901 (N_2901,N_2890,N_2883);
or U2902 (N_2902,N_2867,N_2882);
xnor U2903 (N_2903,N_2857,N_2880);
and U2904 (N_2904,N_2898,N_2864);
nand U2905 (N_2905,N_2896,N_2876);
xor U2906 (N_2906,N_2859,N_2866);
and U2907 (N_2907,N_2897,N_2868);
or U2908 (N_2908,N_2885,N_2872);
nor U2909 (N_2909,N_2887,N_2871);
nand U2910 (N_2910,N_2895,N_2894);
nand U2911 (N_2911,N_2874,N_2879);
nor U2912 (N_2912,N_2878,N_2853);
and U2913 (N_2913,N_2892,N_2850);
nor U2914 (N_2914,N_2854,N_2863);
nand U2915 (N_2915,N_2870,N_2893);
or U2916 (N_2916,N_2875,N_2856);
and U2917 (N_2917,N_2865,N_2851);
nor U2918 (N_2918,N_2873,N_2881);
or U2919 (N_2919,N_2855,N_2852);
xor U2920 (N_2920,N_2869,N_2888);
xnor U2921 (N_2921,N_2860,N_2886);
xnor U2922 (N_2922,N_2861,N_2884);
and U2923 (N_2923,N_2891,N_2889);
xor U2924 (N_2924,N_2862,N_2877);
and U2925 (N_2925,N_2859,N_2895);
nand U2926 (N_2926,N_2892,N_2871);
and U2927 (N_2927,N_2884,N_2883);
xnor U2928 (N_2928,N_2852,N_2854);
and U2929 (N_2929,N_2888,N_2894);
and U2930 (N_2930,N_2875,N_2895);
nand U2931 (N_2931,N_2899,N_2853);
nand U2932 (N_2932,N_2858,N_2855);
or U2933 (N_2933,N_2895,N_2866);
nand U2934 (N_2934,N_2874,N_2894);
nand U2935 (N_2935,N_2892,N_2882);
or U2936 (N_2936,N_2886,N_2851);
nor U2937 (N_2937,N_2885,N_2873);
xor U2938 (N_2938,N_2861,N_2890);
nand U2939 (N_2939,N_2851,N_2893);
and U2940 (N_2940,N_2868,N_2893);
nand U2941 (N_2941,N_2856,N_2871);
and U2942 (N_2942,N_2892,N_2874);
xnor U2943 (N_2943,N_2857,N_2873);
nand U2944 (N_2944,N_2892,N_2880);
nand U2945 (N_2945,N_2858,N_2866);
and U2946 (N_2946,N_2862,N_2884);
nand U2947 (N_2947,N_2852,N_2877);
or U2948 (N_2948,N_2887,N_2852);
nand U2949 (N_2949,N_2861,N_2886);
xnor U2950 (N_2950,N_2924,N_2917);
and U2951 (N_2951,N_2911,N_2947);
nor U2952 (N_2952,N_2934,N_2916);
nor U2953 (N_2953,N_2939,N_2919);
and U2954 (N_2954,N_2935,N_2933);
and U2955 (N_2955,N_2936,N_2925);
xnor U2956 (N_2956,N_2913,N_2941);
and U2957 (N_2957,N_2909,N_2942);
and U2958 (N_2958,N_2902,N_2927);
and U2959 (N_2959,N_2948,N_2932);
or U2960 (N_2960,N_2944,N_2904);
and U2961 (N_2961,N_2921,N_2906);
nand U2962 (N_2962,N_2945,N_2930);
xnor U2963 (N_2963,N_2910,N_2923);
nand U2964 (N_2964,N_2914,N_2949);
and U2965 (N_2965,N_2943,N_2907);
nand U2966 (N_2966,N_2915,N_2918);
nand U2967 (N_2967,N_2940,N_2901);
and U2968 (N_2968,N_2929,N_2905);
xnor U2969 (N_2969,N_2937,N_2928);
xor U2970 (N_2970,N_2926,N_2900);
xnor U2971 (N_2971,N_2903,N_2920);
nor U2972 (N_2972,N_2922,N_2938);
or U2973 (N_2973,N_2912,N_2931);
or U2974 (N_2974,N_2946,N_2908);
nand U2975 (N_2975,N_2908,N_2929);
and U2976 (N_2976,N_2915,N_2900);
xnor U2977 (N_2977,N_2924,N_2939);
nor U2978 (N_2978,N_2907,N_2942);
xnor U2979 (N_2979,N_2916,N_2902);
nand U2980 (N_2980,N_2932,N_2947);
nand U2981 (N_2981,N_2935,N_2941);
nor U2982 (N_2982,N_2912,N_2947);
nand U2983 (N_2983,N_2903,N_2917);
and U2984 (N_2984,N_2936,N_2922);
xor U2985 (N_2985,N_2911,N_2933);
or U2986 (N_2986,N_2909,N_2949);
or U2987 (N_2987,N_2933,N_2904);
nor U2988 (N_2988,N_2914,N_2941);
nor U2989 (N_2989,N_2912,N_2915);
or U2990 (N_2990,N_2908,N_2931);
nor U2991 (N_2991,N_2911,N_2917);
xor U2992 (N_2992,N_2939,N_2910);
and U2993 (N_2993,N_2934,N_2948);
xnor U2994 (N_2994,N_2916,N_2928);
nor U2995 (N_2995,N_2911,N_2908);
and U2996 (N_2996,N_2911,N_2926);
nor U2997 (N_2997,N_2906,N_2940);
or U2998 (N_2998,N_2948,N_2917);
and U2999 (N_2999,N_2912,N_2906);
nand UO_0 (O_0,N_2970,N_2983);
nand UO_1 (O_1,N_2968,N_2974);
nor UO_2 (O_2,N_2952,N_2991);
xnor UO_3 (O_3,N_2999,N_2967);
nor UO_4 (O_4,N_2997,N_2988);
or UO_5 (O_5,N_2956,N_2984);
or UO_6 (O_6,N_2963,N_2978);
or UO_7 (O_7,N_2966,N_2990);
and UO_8 (O_8,N_2964,N_2965);
nor UO_9 (O_9,N_2996,N_2969);
nor UO_10 (O_10,N_2961,N_2962);
nor UO_11 (O_11,N_2987,N_2973);
xnor UO_12 (O_12,N_2959,N_2951);
nor UO_13 (O_13,N_2995,N_2981);
nand UO_14 (O_14,N_2994,N_2986);
nand UO_15 (O_15,N_2979,N_2958);
xnor UO_16 (O_16,N_2975,N_2960);
and UO_17 (O_17,N_2998,N_2950);
xor UO_18 (O_18,N_2982,N_2976);
nor UO_19 (O_19,N_2953,N_2957);
and UO_20 (O_20,N_2993,N_2992);
nand UO_21 (O_21,N_2971,N_2954);
nand UO_22 (O_22,N_2985,N_2989);
and UO_23 (O_23,N_2972,N_2980);
nor UO_24 (O_24,N_2977,N_2955);
and UO_25 (O_25,N_2984,N_2959);
xnor UO_26 (O_26,N_2957,N_2952);
and UO_27 (O_27,N_2984,N_2960);
and UO_28 (O_28,N_2981,N_2996);
and UO_29 (O_29,N_2988,N_2966);
and UO_30 (O_30,N_2995,N_2970);
or UO_31 (O_31,N_2998,N_2968);
and UO_32 (O_32,N_2984,N_2979);
and UO_33 (O_33,N_2988,N_2950);
nand UO_34 (O_34,N_2979,N_2968);
and UO_35 (O_35,N_2969,N_2991);
or UO_36 (O_36,N_2973,N_2960);
and UO_37 (O_37,N_2981,N_2997);
and UO_38 (O_38,N_2985,N_2956);
xor UO_39 (O_39,N_2997,N_2959);
xnor UO_40 (O_40,N_2950,N_2979);
or UO_41 (O_41,N_2962,N_2988);
nand UO_42 (O_42,N_2993,N_2964);
nor UO_43 (O_43,N_2958,N_2960);
nand UO_44 (O_44,N_2959,N_2967);
nor UO_45 (O_45,N_2997,N_2957);
xnor UO_46 (O_46,N_2983,N_2978);
xor UO_47 (O_47,N_2950,N_2977);
nor UO_48 (O_48,N_2967,N_2971);
nand UO_49 (O_49,N_2970,N_2980);
or UO_50 (O_50,N_2984,N_2974);
nand UO_51 (O_51,N_2995,N_2967);
or UO_52 (O_52,N_2958,N_2970);
xnor UO_53 (O_53,N_2983,N_2985);
or UO_54 (O_54,N_2983,N_2982);
nand UO_55 (O_55,N_2978,N_2966);
nor UO_56 (O_56,N_2973,N_2996);
nand UO_57 (O_57,N_2971,N_2988);
nor UO_58 (O_58,N_2988,N_2982);
xor UO_59 (O_59,N_2965,N_2995);
nand UO_60 (O_60,N_2990,N_2961);
or UO_61 (O_61,N_2985,N_2980);
nand UO_62 (O_62,N_2980,N_2969);
nor UO_63 (O_63,N_2984,N_2972);
xor UO_64 (O_64,N_2998,N_2953);
nor UO_65 (O_65,N_2997,N_2994);
or UO_66 (O_66,N_2957,N_2990);
nand UO_67 (O_67,N_2972,N_2977);
nor UO_68 (O_68,N_2992,N_2995);
or UO_69 (O_69,N_2993,N_2979);
or UO_70 (O_70,N_2969,N_2962);
nand UO_71 (O_71,N_2981,N_2956);
xor UO_72 (O_72,N_2988,N_2976);
and UO_73 (O_73,N_2954,N_2986);
nand UO_74 (O_74,N_2968,N_2971);
xor UO_75 (O_75,N_2965,N_2957);
nand UO_76 (O_76,N_2972,N_2982);
and UO_77 (O_77,N_2951,N_2967);
nor UO_78 (O_78,N_2954,N_2974);
and UO_79 (O_79,N_2964,N_2994);
xor UO_80 (O_80,N_2980,N_2977);
nor UO_81 (O_81,N_2965,N_2991);
xnor UO_82 (O_82,N_2962,N_2973);
and UO_83 (O_83,N_2950,N_2974);
or UO_84 (O_84,N_2986,N_2999);
nor UO_85 (O_85,N_2980,N_2987);
nor UO_86 (O_86,N_2987,N_2983);
and UO_87 (O_87,N_2966,N_2994);
or UO_88 (O_88,N_2995,N_2958);
and UO_89 (O_89,N_2963,N_2972);
nor UO_90 (O_90,N_2993,N_2965);
nor UO_91 (O_91,N_2962,N_2997);
or UO_92 (O_92,N_2973,N_2974);
nor UO_93 (O_93,N_2984,N_2991);
nand UO_94 (O_94,N_2971,N_2974);
nand UO_95 (O_95,N_2965,N_2955);
nand UO_96 (O_96,N_2985,N_2954);
nor UO_97 (O_97,N_2997,N_2973);
nor UO_98 (O_98,N_2997,N_2977);
nor UO_99 (O_99,N_2957,N_2964);
nand UO_100 (O_100,N_2974,N_2999);
or UO_101 (O_101,N_2980,N_2954);
nor UO_102 (O_102,N_2968,N_2981);
nand UO_103 (O_103,N_2966,N_2975);
nand UO_104 (O_104,N_2959,N_2998);
nand UO_105 (O_105,N_2977,N_2991);
or UO_106 (O_106,N_2994,N_2990);
nand UO_107 (O_107,N_2976,N_2968);
or UO_108 (O_108,N_2973,N_2959);
and UO_109 (O_109,N_2979,N_2955);
nand UO_110 (O_110,N_2990,N_2952);
nor UO_111 (O_111,N_2993,N_2954);
nor UO_112 (O_112,N_2967,N_2953);
and UO_113 (O_113,N_2959,N_2964);
or UO_114 (O_114,N_2955,N_2964);
or UO_115 (O_115,N_2981,N_2952);
and UO_116 (O_116,N_2979,N_2980);
nand UO_117 (O_117,N_2957,N_2958);
or UO_118 (O_118,N_2989,N_2964);
and UO_119 (O_119,N_2961,N_2978);
and UO_120 (O_120,N_2976,N_2984);
xnor UO_121 (O_121,N_2963,N_2971);
nor UO_122 (O_122,N_2959,N_2955);
and UO_123 (O_123,N_2970,N_2982);
and UO_124 (O_124,N_2997,N_2976);
and UO_125 (O_125,N_2951,N_2992);
xor UO_126 (O_126,N_2998,N_2958);
nor UO_127 (O_127,N_2992,N_2965);
xor UO_128 (O_128,N_2960,N_2986);
nor UO_129 (O_129,N_2994,N_2982);
xor UO_130 (O_130,N_2966,N_2956);
and UO_131 (O_131,N_2974,N_2962);
nand UO_132 (O_132,N_2956,N_2990);
nand UO_133 (O_133,N_2978,N_2979);
and UO_134 (O_134,N_2987,N_2975);
nand UO_135 (O_135,N_2996,N_2988);
nor UO_136 (O_136,N_2967,N_2997);
and UO_137 (O_137,N_2991,N_2957);
nor UO_138 (O_138,N_2958,N_2950);
nor UO_139 (O_139,N_2953,N_2966);
nand UO_140 (O_140,N_2957,N_2968);
xnor UO_141 (O_141,N_2997,N_2960);
and UO_142 (O_142,N_2977,N_2966);
nor UO_143 (O_143,N_2992,N_2988);
and UO_144 (O_144,N_2978,N_2951);
nor UO_145 (O_145,N_2960,N_2993);
nor UO_146 (O_146,N_2979,N_2953);
xnor UO_147 (O_147,N_2981,N_2963);
nor UO_148 (O_148,N_2969,N_2985);
xor UO_149 (O_149,N_2970,N_2975);
xor UO_150 (O_150,N_2961,N_2968);
and UO_151 (O_151,N_2978,N_2999);
xor UO_152 (O_152,N_2951,N_2976);
nor UO_153 (O_153,N_2951,N_2955);
and UO_154 (O_154,N_2987,N_2968);
or UO_155 (O_155,N_2950,N_2996);
and UO_156 (O_156,N_2995,N_2960);
nor UO_157 (O_157,N_2985,N_2966);
and UO_158 (O_158,N_2990,N_2999);
xor UO_159 (O_159,N_2981,N_2951);
or UO_160 (O_160,N_2971,N_2959);
xor UO_161 (O_161,N_2975,N_2964);
nand UO_162 (O_162,N_2966,N_2969);
or UO_163 (O_163,N_2982,N_2981);
nand UO_164 (O_164,N_2953,N_2964);
nand UO_165 (O_165,N_2993,N_2970);
or UO_166 (O_166,N_2995,N_2987);
or UO_167 (O_167,N_2950,N_2970);
nor UO_168 (O_168,N_2993,N_2968);
nor UO_169 (O_169,N_2955,N_2971);
or UO_170 (O_170,N_2978,N_2990);
or UO_171 (O_171,N_2975,N_2980);
xor UO_172 (O_172,N_2985,N_2960);
and UO_173 (O_173,N_2992,N_2963);
and UO_174 (O_174,N_2970,N_2961);
or UO_175 (O_175,N_2967,N_2988);
nor UO_176 (O_176,N_2965,N_2985);
or UO_177 (O_177,N_2982,N_2966);
nor UO_178 (O_178,N_2953,N_2984);
nor UO_179 (O_179,N_2960,N_2964);
xnor UO_180 (O_180,N_2976,N_2952);
xor UO_181 (O_181,N_2978,N_2971);
nor UO_182 (O_182,N_2958,N_2954);
xor UO_183 (O_183,N_2967,N_2954);
nand UO_184 (O_184,N_2957,N_2971);
nor UO_185 (O_185,N_2962,N_2986);
xnor UO_186 (O_186,N_2986,N_2961);
nor UO_187 (O_187,N_2966,N_2973);
and UO_188 (O_188,N_2972,N_2988);
and UO_189 (O_189,N_2989,N_2950);
nand UO_190 (O_190,N_2992,N_2991);
nand UO_191 (O_191,N_2994,N_2961);
nand UO_192 (O_192,N_2989,N_2983);
or UO_193 (O_193,N_2958,N_2978);
and UO_194 (O_194,N_2973,N_2983);
nor UO_195 (O_195,N_2982,N_2959);
or UO_196 (O_196,N_2973,N_2963);
xnor UO_197 (O_197,N_2999,N_2987);
and UO_198 (O_198,N_2991,N_2998);
and UO_199 (O_199,N_2991,N_2955);
or UO_200 (O_200,N_2950,N_2986);
xnor UO_201 (O_201,N_2965,N_2967);
nand UO_202 (O_202,N_2960,N_2976);
or UO_203 (O_203,N_2989,N_2966);
nor UO_204 (O_204,N_2994,N_2985);
xor UO_205 (O_205,N_2960,N_2981);
nand UO_206 (O_206,N_2990,N_2987);
nor UO_207 (O_207,N_2976,N_2967);
or UO_208 (O_208,N_2984,N_2981);
or UO_209 (O_209,N_2988,N_2964);
xnor UO_210 (O_210,N_2968,N_2991);
xor UO_211 (O_211,N_2974,N_2998);
xor UO_212 (O_212,N_2978,N_2965);
nand UO_213 (O_213,N_2955,N_2952);
or UO_214 (O_214,N_2998,N_2973);
nand UO_215 (O_215,N_2993,N_2990);
xnor UO_216 (O_216,N_2968,N_2986);
nand UO_217 (O_217,N_2994,N_2983);
and UO_218 (O_218,N_2979,N_2957);
nor UO_219 (O_219,N_2970,N_2992);
xor UO_220 (O_220,N_2962,N_2955);
or UO_221 (O_221,N_2971,N_2953);
nand UO_222 (O_222,N_2971,N_2950);
nor UO_223 (O_223,N_2975,N_2968);
and UO_224 (O_224,N_2968,N_2952);
or UO_225 (O_225,N_2963,N_2969);
nor UO_226 (O_226,N_2978,N_2977);
nand UO_227 (O_227,N_2958,N_2985);
nor UO_228 (O_228,N_2961,N_2975);
xor UO_229 (O_229,N_2956,N_2968);
and UO_230 (O_230,N_2989,N_2995);
nand UO_231 (O_231,N_2958,N_2980);
and UO_232 (O_232,N_2973,N_2957);
nand UO_233 (O_233,N_2963,N_2995);
or UO_234 (O_234,N_2954,N_2961);
xnor UO_235 (O_235,N_2972,N_2951);
or UO_236 (O_236,N_2961,N_2964);
or UO_237 (O_237,N_2987,N_2985);
or UO_238 (O_238,N_2962,N_2953);
nand UO_239 (O_239,N_2992,N_2955);
nor UO_240 (O_240,N_2999,N_2964);
nand UO_241 (O_241,N_2990,N_2960);
and UO_242 (O_242,N_2989,N_2978);
and UO_243 (O_243,N_2987,N_2976);
or UO_244 (O_244,N_2980,N_2993);
nor UO_245 (O_245,N_2973,N_2969);
nor UO_246 (O_246,N_2956,N_2950);
or UO_247 (O_247,N_2995,N_2983);
and UO_248 (O_248,N_2955,N_2982);
and UO_249 (O_249,N_2951,N_2965);
xor UO_250 (O_250,N_2981,N_2965);
xnor UO_251 (O_251,N_2970,N_2979);
nor UO_252 (O_252,N_2956,N_2965);
or UO_253 (O_253,N_2990,N_2996);
nand UO_254 (O_254,N_2981,N_2999);
and UO_255 (O_255,N_2974,N_2981);
xor UO_256 (O_256,N_2973,N_2988);
xor UO_257 (O_257,N_2950,N_2954);
nor UO_258 (O_258,N_2977,N_2951);
and UO_259 (O_259,N_2991,N_2966);
nand UO_260 (O_260,N_2997,N_2996);
or UO_261 (O_261,N_2978,N_2953);
and UO_262 (O_262,N_2970,N_2972);
or UO_263 (O_263,N_2995,N_2979);
nor UO_264 (O_264,N_2958,N_2984);
nand UO_265 (O_265,N_2955,N_2968);
nor UO_266 (O_266,N_2985,N_2991);
xnor UO_267 (O_267,N_2966,N_2976);
or UO_268 (O_268,N_2967,N_2958);
xnor UO_269 (O_269,N_2957,N_2995);
nand UO_270 (O_270,N_2977,N_2994);
nand UO_271 (O_271,N_2993,N_2988);
nor UO_272 (O_272,N_2985,N_2950);
nor UO_273 (O_273,N_2991,N_2963);
nor UO_274 (O_274,N_2974,N_2956);
nor UO_275 (O_275,N_2996,N_2974);
nand UO_276 (O_276,N_2985,N_2998);
xnor UO_277 (O_277,N_2957,N_2950);
nor UO_278 (O_278,N_2969,N_2968);
nor UO_279 (O_279,N_2992,N_2968);
or UO_280 (O_280,N_2970,N_2977);
nor UO_281 (O_281,N_2997,N_2969);
or UO_282 (O_282,N_2965,N_2996);
nor UO_283 (O_283,N_2994,N_2993);
and UO_284 (O_284,N_2951,N_2962);
nor UO_285 (O_285,N_2963,N_2953);
nor UO_286 (O_286,N_2969,N_2954);
nand UO_287 (O_287,N_2999,N_2969);
nor UO_288 (O_288,N_2952,N_2975);
and UO_289 (O_289,N_2968,N_2999);
and UO_290 (O_290,N_2974,N_2979);
and UO_291 (O_291,N_2953,N_2958);
and UO_292 (O_292,N_2958,N_2951);
or UO_293 (O_293,N_2990,N_2995);
or UO_294 (O_294,N_2954,N_2979);
and UO_295 (O_295,N_2999,N_2950);
nor UO_296 (O_296,N_2968,N_2972);
and UO_297 (O_297,N_2968,N_2966);
nand UO_298 (O_298,N_2964,N_2990);
nor UO_299 (O_299,N_2989,N_2961);
xor UO_300 (O_300,N_2963,N_2989);
nand UO_301 (O_301,N_2963,N_2954);
and UO_302 (O_302,N_2956,N_2953);
and UO_303 (O_303,N_2995,N_2997);
or UO_304 (O_304,N_2963,N_2993);
nand UO_305 (O_305,N_2999,N_2977);
nand UO_306 (O_306,N_2984,N_2967);
or UO_307 (O_307,N_2979,N_2959);
nor UO_308 (O_308,N_2961,N_2952);
or UO_309 (O_309,N_2985,N_2961);
and UO_310 (O_310,N_2965,N_2977);
or UO_311 (O_311,N_2976,N_2958);
xnor UO_312 (O_312,N_2971,N_2964);
xor UO_313 (O_313,N_2992,N_2983);
and UO_314 (O_314,N_2990,N_2972);
nand UO_315 (O_315,N_2987,N_2981);
nand UO_316 (O_316,N_2998,N_2952);
nor UO_317 (O_317,N_2969,N_2978);
and UO_318 (O_318,N_2998,N_2969);
and UO_319 (O_319,N_2979,N_2998);
xnor UO_320 (O_320,N_2958,N_2987);
nor UO_321 (O_321,N_2996,N_2972);
xnor UO_322 (O_322,N_2994,N_2992);
and UO_323 (O_323,N_2970,N_2959);
and UO_324 (O_324,N_2969,N_2951);
nor UO_325 (O_325,N_2954,N_2984);
nor UO_326 (O_326,N_2951,N_2970);
or UO_327 (O_327,N_2974,N_2990);
nand UO_328 (O_328,N_2969,N_2971);
xnor UO_329 (O_329,N_2964,N_2982);
and UO_330 (O_330,N_2992,N_2978);
or UO_331 (O_331,N_2953,N_2960);
and UO_332 (O_332,N_2991,N_2951);
nand UO_333 (O_333,N_2961,N_2979);
nor UO_334 (O_334,N_2994,N_2952);
xnor UO_335 (O_335,N_2956,N_2955);
and UO_336 (O_336,N_2960,N_2954);
or UO_337 (O_337,N_2994,N_2955);
nor UO_338 (O_338,N_2966,N_2984);
and UO_339 (O_339,N_2976,N_2994);
and UO_340 (O_340,N_2972,N_2978);
or UO_341 (O_341,N_2999,N_2972);
nor UO_342 (O_342,N_2983,N_2953);
or UO_343 (O_343,N_2961,N_2980);
and UO_344 (O_344,N_2989,N_2986);
and UO_345 (O_345,N_2963,N_2964);
nor UO_346 (O_346,N_2952,N_2969);
and UO_347 (O_347,N_2977,N_2960);
and UO_348 (O_348,N_2962,N_2954);
nand UO_349 (O_349,N_2987,N_2972);
nand UO_350 (O_350,N_2981,N_2993);
nand UO_351 (O_351,N_2999,N_2957);
or UO_352 (O_352,N_2951,N_2952);
and UO_353 (O_353,N_2968,N_2962);
nand UO_354 (O_354,N_2966,N_2964);
nand UO_355 (O_355,N_2961,N_2956);
nor UO_356 (O_356,N_2974,N_2953);
and UO_357 (O_357,N_2981,N_2967);
or UO_358 (O_358,N_2975,N_2979);
nor UO_359 (O_359,N_2994,N_2953);
or UO_360 (O_360,N_2955,N_2974);
or UO_361 (O_361,N_2979,N_2963);
or UO_362 (O_362,N_2959,N_2953);
or UO_363 (O_363,N_2992,N_2958);
xor UO_364 (O_364,N_2960,N_2980);
nand UO_365 (O_365,N_2953,N_2976);
and UO_366 (O_366,N_2999,N_2975);
xor UO_367 (O_367,N_2975,N_2983);
or UO_368 (O_368,N_2987,N_2974);
or UO_369 (O_369,N_2963,N_2974);
and UO_370 (O_370,N_2963,N_2965);
and UO_371 (O_371,N_2967,N_2970);
or UO_372 (O_372,N_2966,N_2980);
nor UO_373 (O_373,N_2962,N_2971);
nand UO_374 (O_374,N_2992,N_2967);
nand UO_375 (O_375,N_2962,N_2964);
xnor UO_376 (O_376,N_2954,N_2996);
nor UO_377 (O_377,N_2993,N_2969);
or UO_378 (O_378,N_2995,N_2993);
or UO_379 (O_379,N_2961,N_2993);
and UO_380 (O_380,N_2969,N_2958);
nand UO_381 (O_381,N_2970,N_2996);
xnor UO_382 (O_382,N_2982,N_2987);
nor UO_383 (O_383,N_2997,N_2954);
nand UO_384 (O_384,N_2966,N_2951);
xnor UO_385 (O_385,N_2993,N_2953);
xnor UO_386 (O_386,N_2969,N_2977);
xnor UO_387 (O_387,N_2980,N_2995);
and UO_388 (O_388,N_2972,N_2997);
nor UO_389 (O_389,N_2973,N_2965);
xor UO_390 (O_390,N_2995,N_2999);
or UO_391 (O_391,N_2954,N_2998);
and UO_392 (O_392,N_2961,N_2955);
or UO_393 (O_393,N_2994,N_2962);
nor UO_394 (O_394,N_2997,N_2965);
xor UO_395 (O_395,N_2972,N_2985);
nand UO_396 (O_396,N_2994,N_2971);
xnor UO_397 (O_397,N_2969,N_2970);
xnor UO_398 (O_398,N_2983,N_2993);
nand UO_399 (O_399,N_2952,N_2970);
nor UO_400 (O_400,N_2952,N_2977);
xnor UO_401 (O_401,N_2994,N_2959);
or UO_402 (O_402,N_2988,N_2983);
nor UO_403 (O_403,N_2972,N_2973);
xor UO_404 (O_404,N_2998,N_2984);
or UO_405 (O_405,N_2963,N_2986);
nor UO_406 (O_406,N_2955,N_2978);
nand UO_407 (O_407,N_2984,N_2950);
and UO_408 (O_408,N_2955,N_2996);
xnor UO_409 (O_409,N_2956,N_2994);
xnor UO_410 (O_410,N_2958,N_2973);
nand UO_411 (O_411,N_2989,N_2953);
xor UO_412 (O_412,N_2990,N_2970);
nand UO_413 (O_413,N_2985,N_2952);
xor UO_414 (O_414,N_2973,N_2954);
nand UO_415 (O_415,N_2985,N_2967);
nor UO_416 (O_416,N_2980,N_2982);
xnor UO_417 (O_417,N_2953,N_2955);
and UO_418 (O_418,N_2960,N_2959);
or UO_419 (O_419,N_2980,N_2963);
nand UO_420 (O_420,N_2950,N_2981);
xnor UO_421 (O_421,N_2986,N_2965);
nor UO_422 (O_422,N_2999,N_2979);
and UO_423 (O_423,N_2969,N_2994);
nor UO_424 (O_424,N_2988,N_2991);
and UO_425 (O_425,N_2964,N_2956);
nand UO_426 (O_426,N_2994,N_2965);
or UO_427 (O_427,N_2956,N_2952);
and UO_428 (O_428,N_2965,N_2983);
and UO_429 (O_429,N_2990,N_2959);
nor UO_430 (O_430,N_2994,N_2996);
nor UO_431 (O_431,N_2954,N_2989);
or UO_432 (O_432,N_2973,N_2980);
nor UO_433 (O_433,N_2985,N_2964);
or UO_434 (O_434,N_2963,N_2983);
and UO_435 (O_435,N_2999,N_2994);
nand UO_436 (O_436,N_2972,N_2969);
nand UO_437 (O_437,N_2956,N_2983);
nor UO_438 (O_438,N_2976,N_2985);
nor UO_439 (O_439,N_2981,N_2955);
nand UO_440 (O_440,N_2956,N_2959);
nor UO_441 (O_441,N_2985,N_2997);
and UO_442 (O_442,N_2980,N_2974);
xor UO_443 (O_443,N_2960,N_2999);
or UO_444 (O_444,N_2959,N_2996);
nor UO_445 (O_445,N_2957,N_2954);
and UO_446 (O_446,N_2962,N_2952);
nand UO_447 (O_447,N_2997,N_2958);
or UO_448 (O_448,N_2996,N_2960);
or UO_449 (O_449,N_2952,N_2986);
xor UO_450 (O_450,N_2980,N_2997);
and UO_451 (O_451,N_2952,N_2984);
xnor UO_452 (O_452,N_2982,N_2956);
xnor UO_453 (O_453,N_2959,N_2975);
nor UO_454 (O_454,N_2988,N_2975);
and UO_455 (O_455,N_2988,N_2984);
xor UO_456 (O_456,N_2974,N_2957);
xnor UO_457 (O_457,N_2955,N_2987);
nand UO_458 (O_458,N_2990,N_2986);
or UO_459 (O_459,N_2996,N_2971);
or UO_460 (O_460,N_2957,N_2967);
or UO_461 (O_461,N_2956,N_2986);
nand UO_462 (O_462,N_2980,N_2951);
or UO_463 (O_463,N_2955,N_2957);
nand UO_464 (O_464,N_2958,N_2975);
xor UO_465 (O_465,N_2970,N_2999);
nor UO_466 (O_466,N_2974,N_2982);
nand UO_467 (O_467,N_2970,N_2981);
xor UO_468 (O_468,N_2987,N_2959);
nor UO_469 (O_469,N_2977,N_2998);
and UO_470 (O_470,N_2967,N_2996);
and UO_471 (O_471,N_2957,N_2981);
nor UO_472 (O_472,N_2975,N_2989);
or UO_473 (O_473,N_2990,N_2981);
xor UO_474 (O_474,N_2979,N_2983);
nand UO_475 (O_475,N_2954,N_2982);
and UO_476 (O_476,N_2965,N_2988);
nand UO_477 (O_477,N_2963,N_2999);
and UO_478 (O_478,N_2969,N_2987);
nand UO_479 (O_479,N_2984,N_2983);
xnor UO_480 (O_480,N_2984,N_2989);
nand UO_481 (O_481,N_2960,N_2971);
xor UO_482 (O_482,N_2970,N_2964);
nor UO_483 (O_483,N_2988,N_2957);
or UO_484 (O_484,N_2980,N_2991);
xor UO_485 (O_485,N_2982,N_2984);
nor UO_486 (O_486,N_2959,N_2962);
nand UO_487 (O_487,N_2974,N_2960);
or UO_488 (O_488,N_2989,N_2977);
or UO_489 (O_489,N_2972,N_2993);
and UO_490 (O_490,N_2952,N_2967);
and UO_491 (O_491,N_2952,N_2966);
or UO_492 (O_492,N_2970,N_2963);
and UO_493 (O_493,N_2958,N_2996);
and UO_494 (O_494,N_2971,N_2951);
nor UO_495 (O_495,N_2959,N_2961);
and UO_496 (O_496,N_2987,N_2961);
and UO_497 (O_497,N_2993,N_2985);
xor UO_498 (O_498,N_2966,N_2955);
or UO_499 (O_499,N_2991,N_2967);
endmodule