module basic_1500_15000_2000_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_164,In_1155);
nor U1 (N_1,In_969,In_653);
or U2 (N_2,In_89,In_370);
nor U3 (N_3,In_910,In_966);
nor U4 (N_4,In_1188,In_1207);
or U5 (N_5,In_1237,In_744);
and U6 (N_6,In_987,In_142);
nor U7 (N_7,In_1395,In_1439);
nand U8 (N_8,In_162,In_1114);
or U9 (N_9,In_1320,In_464);
nor U10 (N_10,In_230,In_1105);
and U11 (N_11,In_156,In_1380);
nor U12 (N_12,In_440,In_1092);
or U13 (N_13,In_1441,In_338);
or U14 (N_14,In_480,In_1473);
xor U15 (N_15,In_256,In_1219);
and U16 (N_16,In_898,In_258);
nor U17 (N_17,In_14,In_229);
or U18 (N_18,In_246,In_677);
nand U19 (N_19,In_38,In_260);
nand U20 (N_20,In_1257,In_130);
nor U21 (N_21,In_885,In_163);
nand U22 (N_22,In_176,In_105);
nor U23 (N_23,In_947,In_1338);
nand U24 (N_24,In_1429,In_1341);
or U25 (N_25,In_921,In_414);
or U26 (N_26,In_812,In_1321);
or U27 (N_27,In_1098,In_709);
nor U28 (N_28,In_347,In_915);
and U29 (N_29,In_1012,In_1040);
or U30 (N_30,In_594,In_834);
or U31 (N_31,In_1252,In_962);
and U32 (N_32,In_1293,In_682);
xor U33 (N_33,In_447,In_1397);
nor U34 (N_34,In_1280,In_542);
xor U35 (N_35,In_134,In_1262);
and U36 (N_36,In_330,In_832);
and U37 (N_37,In_761,In_1294);
xor U38 (N_38,In_58,In_1110);
or U39 (N_39,In_614,In_143);
nor U40 (N_40,In_1408,In_92);
nand U41 (N_41,In_1327,In_1425);
nor U42 (N_42,In_1011,In_1119);
nand U43 (N_43,In_666,In_505);
and U44 (N_44,In_1416,In_301);
xnor U45 (N_45,In_263,In_1363);
nand U46 (N_46,In_663,In_1185);
and U47 (N_47,In_506,In_765);
nand U48 (N_48,In_76,In_1041);
nor U49 (N_49,In_40,In_1485);
nand U50 (N_50,In_46,In_729);
nand U51 (N_51,In_39,In_387);
nand U52 (N_52,In_1230,In_552);
xor U53 (N_53,In_79,In_169);
nor U54 (N_54,In_826,In_860);
nand U55 (N_55,In_689,In_897);
xor U56 (N_56,In_1169,In_868);
xnor U57 (N_57,In_920,In_1287);
and U58 (N_58,In_109,In_596);
or U59 (N_59,In_1042,In_1392);
or U60 (N_60,In_1153,In_1051);
and U61 (N_61,In_408,In_439);
or U62 (N_62,In_1196,In_120);
xor U63 (N_63,In_65,In_803);
nand U64 (N_64,In_31,In_168);
and U65 (N_65,In_787,In_157);
nand U66 (N_66,In_1118,In_1282);
and U67 (N_67,In_784,In_170);
xnor U68 (N_68,In_1140,In_716);
nand U69 (N_69,In_607,In_1102);
nand U70 (N_70,In_1091,In_304);
nor U71 (N_71,In_753,In_904);
xnor U72 (N_72,In_1306,In_715);
nor U73 (N_73,In_61,In_652);
xnor U74 (N_74,In_1399,In_686);
and U75 (N_75,In_205,In_1220);
nand U76 (N_76,In_838,In_366);
nand U77 (N_77,In_118,In_990);
or U78 (N_78,In_140,In_422);
nand U79 (N_79,In_911,In_1029);
or U80 (N_80,In_1034,In_1036);
nor U81 (N_81,In_353,In_1284);
xor U82 (N_82,In_1240,In_566);
nor U83 (N_83,In_1386,In_488);
or U84 (N_84,In_1424,In_858);
and U85 (N_85,In_1404,In_1212);
nor U86 (N_86,In_467,In_285);
or U87 (N_87,In_679,In_411);
xor U88 (N_88,In_953,In_828);
nand U89 (N_89,In_786,In_329);
nor U90 (N_90,In_1097,In_691);
xor U91 (N_91,In_327,In_863);
and U92 (N_92,In_1088,In_1239);
and U93 (N_93,In_444,In_1455);
xor U94 (N_94,In_208,In_597);
nor U95 (N_95,In_27,In_1382);
nand U96 (N_96,In_1411,In_23);
and U97 (N_97,In_1182,In_474);
and U98 (N_98,In_537,In_373);
or U99 (N_99,In_982,In_1044);
xor U100 (N_100,In_397,In_1347);
and U101 (N_101,In_276,In_351);
or U102 (N_102,In_1497,In_903);
nand U103 (N_103,In_1020,In_577);
xnor U104 (N_104,In_1204,In_1215);
nand U105 (N_105,In_18,In_487);
nand U106 (N_106,In_405,In_644);
and U107 (N_107,In_1146,In_348);
or U108 (N_108,In_1434,In_1470);
or U109 (N_109,In_575,In_764);
and U110 (N_110,In_1054,In_1197);
nor U111 (N_111,In_981,In_572);
and U112 (N_112,In_1383,In_323);
nor U113 (N_113,In_1006,In_974);
or U114 (N_114,In_889,In_269);
nor U115 (N_115,In_426,In_1475);
xor U116 (N_116,In_382,In_934);
nor U117 (N_117,In_1431,In_1192);
and U118 (N_118,In_410,In_1353);
or U119 (N_119,In_96,In_855);
or U120 (N_120,In_1414,In_99);
or U121 (N_121,In_12,In_559);
or U122 (N_122,In_565,In_512);
or U123 (N_123,In_1229,In_17);
and U124 (N_124,In_1141,In_1448);
nand U125 (N_125,In_539,In_1325);
xor U126 (N_126,In_215,In_888);
and U127 (N_127,In_665,In_775);
nand U128 (N_128,In_621,In_504);
or U129 (N_129,In_106,In_1365);
or U130 (N_130,In_554,In_191);
or U131 (N_131,In_7,In_83);
or U132 (N_132,In_1168,In_958);
xnor U133 (N_133,In_478,In_1162);
nor U134 (N_134,In_1303,In_155);
nand U135 (N_135,In_290,In_154);
nand U136 (N_136,In_995,In_736);
nand U137 (N_137,In_690,In_1461);
or U138 (N_138,In_259,In_1205);
nor U139 (N_139,In_707,In_453);
nand U140 (N_140,In_1276,In_948);
xor U141 (N_141,In_454,In_1202);
or U142 (N_142,In_362,In_67);
or U143 (N_143,In_695,In_943);
and U144 (N_144,In_1055,In_1076);
and U145 (N_145,In_561,In_1050);
xnor U146 (N_146,In_312,In_827);
or U147 (N_147,In_908,In_1243);
nor U148 (N_148,In_590,In_203);
and U149 (N_149,In_1158,In_1357);
nor U150 (N_150,In_267,In_902);
and U151 (N_151,In_49,In_610);
or U152 (N_152,In_459,In_726);
nor U153 (N_153,In_1173,In_808);
xnor U154 (N_154,In_125,In_739);
xnor U155 (N_155,In_905,In_1016);
xnor U156 (N_156,In_694,In_961);
xor U157 (N_157,In_421,In_692);
nor U158 (N_158,In_510,In_669);
nand U159 (N_159,In_1305,In_1270);
xnor U160 (N_160,In_873,In_317);
nor U161 (N_161,In_1242,In_104);
and U162 (N_162,In_28,In_69);
nand U163 (N_163,In_917,In_791);
xnor U164 (N_164,In_697,In_207);
and U165 (N_165,In_306,In_980);
nor U166 (N_166,In_967,In_1444);
and U167 (N_167,In_245,In_1260);
nor U168 (N_168,In_159,In_428);
nor U169 (N_169,In_706,In_318);
or U170 (N_170,In_1032,In_448);
or U171 (N_171,In_196,In_634);
xor U172 (N_172,In_1261,In_1269);
or U173 (N_173,In_138,In_399);
nand U174 (N_174,In_1334,In_1060);
nor U175 (N_175,In_303,In_1391);
or U176 (N_176,In_293,In_342);
nor U177 (N_177,In_1130,In_821);
and U178 (N_178,In_26,In_678);
xnor U179 (N_179,In_1389,In_1449);
xor U180 (N_180,In_675,In_641);
xor U181 (N_181,In_1175,In_1376);
and U182 (N_182,In_713,In_37);
nand U183 (N_183,In_625,In_1275);
or U184 (N_184,In_704,In_647);
nor U185 (N_185,In_853,In_1329);
xor U186 (N_186,In_305,In_1154);
nand U187 (N_187,In_384,In_320);
nor U188 (N_188,In_1206,In_355);
and U189 (N_189,In_1106,In_358);
nor U190 (N_190,In_1156,In_438);
nand U191 (N_191,In_396,In_1493);
and U192 (N_192,In_298,In_1422);
nand U193 (N_193,In_97,In_785);
or U194 (N_194,In_291,In_667);
xor U195 (N_195,In_1074,In_486);
nand U196 (N_196,In_1007,In_328);
and U197 (N_197,In_296,In_1132);
nand U198 (N_198,In_72,In_1001);
nor U199 (N_199,In_899,In_13);
or U200 (N_200,In_606,In_1332);
and U201 (N_201,In_287,In_107);
xor U202 (N_202,In_1405,In_361);
and U203 (N_203,In_238,In_643);
xnor U204 (N_204,In_740,In_1316);
xor U205 (N_205,In_225,In_1472);
nand U206 (N_206,In_1069,In_1238);
nor U207 (N_207,In_1131,In_1281);
and U208 (N_208,In_1124,In_839);
or U209 (N_209,In_6,In_758);
nand U210 (N_210,In_1174,In_972);
xnor U211 (N_211,In_752,In_993);
or U212 (N_212,In_137,In_1423);
xor U213 (N_213,In_1375,In_1171);
nor U214 (N_214,In_1300,In_135);
nand U215 (N_215,In_485,In_1120);
and U216 (N_216,In_699,In_870);
and U217 (N_217,In_1498,In_940);
xor U218 (N_218,In_971,In_1013);
and U219 (N_219,In_95,In_901);
or U220 (N_220,In_1138,In_1268);
and U221 (N_221,In_153,In_1234);
or U222 (N_222,In_681,In_618);
xnor U223 (N_223,In_582,In_284);
nor U224 (N_224,In_774,In_569);
nor U225 (N_225,In_592,In_1043);
nand U226 (N_226,In_720,In_1285);
and U227 (N_227,In_42,In_1186);
nand U228 (N_228,In_1116,In_1496);
nand U229 (N_229,In_178,In_450);
or U230 (N_230,In_1189,In_683);
or U231 (N_231,In_1494,In_1048);
nand U232 (N_232,In_1247,In_1021);
nand U233 (N_233,In_710,In_345);
nor U234 (N_234,In_241,In_534);
nor U235 (N_235,In_145,In_657);
and U236 (N_236,In_509,In_550);
xor U237 (N_237,In_892,In_400);
xnor U238 (N_238,In_451,In_1368);
nand U239 (N_239,In_1364,In_1167);
or U240 (N_240,In_136,In_1079);
or U241 (N_241,In_956,In_1481);
nand U242 (N_242,In_456,In_711);
or U243 (N_243,In_1031,In_1142);
and U244 (N_244,In_684,In_623);
xor U245 (N_245,In_211,In_166);
xor U246 (N_246,In_100,In_1297);
and U247 (N_247,In_47,In_435);
nand U248 (N_248,In_824,In_1312);
nand U249 (N_249,In_1396,In_864);
nand U250 (N_250,In_1343,In_1370);
xnor U251 (N_251,In_167,In_831);
and U252 (N_252,In_535,In_991);
or U253 (N_253,In_635,In_514);
nor U254 (N_254,In_760,In_639);
xnor U255 (N_255,In_270,In_1463);
or U256 (N_256,In_1198,In_835);
or U257 (N_257,In_1165,In_1217);
or U258 (N_258,In_231,In_22);
or U259 (N_259,In_1467,In_1214);
nand U260 (N_260,In_1253,In_584);
nor U261 (N_261,In_1177,In_423);
nand U262 (N_262,In_173,In_471);
and U263 (N_263,In_593,In_141);
xnor U264 (N_264,In_806,In_468);
xor U265 (N_265,In_763,In_979);
nand U266 (N_266,In_965,In_1135);
nand U267 (N_267,In_3,In_1213);
and U268 (N_268,In_656,In_1352);
xor U269 (N_269,In_782,In_392);
or U270 (N_270,In_165,In_1336);
nor U271 (N_271,In_19,In_1199);
and U272 (N_272,In_796,In_262);
nand U273 (N_273,In_210,In_1466);
and U274 (N_274,In_1344,In_180);
and U275 (N_275,In_4,In_771);
or U276 (N_276,In_724,In_1170);
nor U277 (N_277,In_802,In_326);
xor U278 (N_278,In_294,In_402);
nand U279 (N_279,In_805,In_676);
xor U280 (N_280,In_574,In_475);
and U281 (N_281,In_543,In_696);
or U282 (N_282,In_360,In_29);
xnor U283 (N_283,In_1264,In_363);
xor U284 (N_284,In_769,In_344);
xor U285 (N_285,In_1258,In_346);
and U286 (N_286,In_236,In_1228);
xnor U287 (N_287,In_1190,In_1317);
or U288 (N_288,In_1419,In_533);
or U289 (N_289,In_1180,In_395);
nand U290 (N_290,In_1053,In_132);
and U291 (N_291,In_209,In_491);
xnor U292 (N_292,In_9,In_466);
nor U293 (N_293,In_64,In_718);
nor U294 (N_294,In_548,In_1447);
nand U295 (N_295,In_1236,In_242);
or U296 (N_296,In_1296,In_1277);
and U297 (N_297,In_161,In_1350);
or U298 (N_298,In_202,In_1273);
nand U299 (N_299,In_30,In_1085);
nand U300 (N_300,In_742,In_755);
or U301 (N_301,In_1271,In_1349);
xnor U302 (N_302,In_1499,In_1417);
and U303 (N_303,In_1224,In_190);
nor U304 (N_304,In_497,In_374);
or U305 (N_305,In_252,In_1468);
xor U306 (N_306,In_449,In_1379);
or U307 (N_307,In_1412,In_1326);
and U308 (N_308,In_1436,In_1272);
nand U309 (N_309,In_484,In_63);
xnor U310 (N_310,In_1469,In_1099);
xnor U311 (N_311,In_531,In_388);
nand U312 (N_312,In_1288,In_1028);
and U313 (N_313,In_1356,In_197);
nand U314 (N_314,In_126,In_1301);
nand U315 (N_315,In_662,In_1433);
and U316 (N_316,In_212,In_1047);
and U317 (N_317,In_978,In_629);
or U318 (N_318,In_1359,In_1160);
or U319 (N_319,In_266,In_1266);
nand U320 (N_320,In_600,In_0);
nor U321 (N_321,In_275,In_232);
or U322 (N_322,In_1018,In_364);
xor U323 (N_323,In_1390,In_833);
and U324 (N_324,In_822,In_174);
nand U325 (N_325,In_340,In_1378);
nand U326 (N_326,In_890,In_856);
or U327 (N_327,In_730,In_1250);
or U328 (N_328,In_315,In_770);
nand U329 (N_329,In_617,In_406);
nand U330 (N_330,In_56,In_1456);
nand U331 (N_331,In_490,In_220);
xnor U332 (N_332,In_1005,In_53);
or U333 (N_333,In_412,In_265);
and U334 (N_334,In_78,In_1195);
xnor U335 (N_335,In_309,In_283);
nor U336 (N_336,In_1394,In_177);
xnor U337 (N_337,In_900,In_98);
xor U338 (N_338,In_576,In_473);
nor U339 (N_339,In_1420,In_268);
or U340 (N_340,In_1454,In_352);
nand U341 (N_341,In_1176,In_564);
nand U342 (N_342,In_48,In_847);
xnor U343 (N_343,In_1314,In_1490);
xor U344 (N_344,In_1015,In_933);
and U345 (N_345,In_1115,In_88);
or U346 (N_346,In_529,In_723);
xor U347 (N_347,In_878,In_460);
or U348 (N_348,In_55,In_333);
nor U349 (N_349,In_337,In_425);
or U350 (N_350,In_70,In_465);
or U351 (N_351,In_804,In_811);
nor U352 (N_352,In_1452,In_372);
xor U353 (N_353,In_1178,In_1355);
nor U354 (N_354,In_1415,In_273);
nand U355 (N_355,In_1299,In_124);
and U356 (N_356,In_1017,In_1111);
and U357 (N_357,In_369,In_1410);
or U358 (N_358,In_640,In_526);
nor U359 (N_359,In_1159,In_861);
or U360 (N_360,In_799,In_217);
xnor U361 (N_361,In_1346,In_813);
and U362 (N_362,In_588,In_1232);
nand U363 (N_363,In_341,In_619);
nand U364 (N_364,In_558,In_302);
or U365 (N_365,In_45,In_1492);
nand U366 (N_366,In_280,In_521);
nand U367 (N_367,In_365,In_5);
nor U368 (N_368,In_527,In_825);
xor U369 (N_369,In_1077,In_759);
or U370 (N_370,In_809,In_181);
and U371 (N_371,In_1061,In_185);
or U372 (N_372,In_913,In_240);
nor U373 (N_373,In_646,In_85);
nand U374 (N_374,In_222,In_658);
nand U375 (N_375,In_1126,In_1478);
nand U376 (N_376,In_1335,In_792);
nand U377 (N_377,In_798,In_1438);
nor U378 (N_378,In_1129,In_1487);
and U379 (N_379,In_386,In_532);
and U380 (N_380,In_213,In_1388);
xor U381 (N_381,In_642,In_1231);
nand U382 (N_382,In_429,In_829);
and U383 (N_383,In_158,In_1121);
nor U384 (N_384,In_865,In_728);
nor U385 (N_385,In_224,In_939);
nor U386 (N_386,In_988,In_339);
and U387 (N_387,In_931,In_489);
nor U388 (N_388,In_923,In_1324);
or U389 (N_389,In_1484,In_616);
or U390 (N_390,In_493,In_630);
and U391 (N_391,In_1402,In_1458);
xnor U392 (N_392,In_627,In_472);
or U393 (N_393,In_1049,In_498);
or U394 (N_394,In_876,In_1128);
and U395 (N_395,In_1244,In_1109);
and U396 (N_396,In_1112,In_117);
or U397 (N_397,In_964,In_1451);
nor U398 (N_398,In_1440,In_1265);
nand U399 (N_399,In_750,In_1211);
xor U400 (N_400,In_551,In_1090);
xnor U401 (N_401,In_122,In_516);
nor U402 (N_402,In_248,In_445);
or U403 (N_403,In_175,In_147);
nor U404 (N_404,In_1249,In_380);
and U405 (N_405,In_906,In_1400);
and U406 (N_406,In_651,In_1457);
xor U407 (N_407,In_247,In_768);
nand U408 (N_408,In_1369,In_80);
nor U409 (N_409,In_114,In_1080);
xnor U410 (N_410,In_243,In_1446);
nor U411 (N_411,In_960,In_549);
nor U412 (N_412,In_547,In_1075);
nor U413 (N_413,In_778,In_857);
xor U414 (N_414,In_82,In_1427);
nand U415 (N_415,In_452,In_872);
nand U416 (N_416,In_1056,In_693);
nor U417 (N_417,In_818,In_705);
or U418 (N_418,In_25,In_1371);
or U419 (N_419,In_846,In_968);
and U420 (N_420,In_119,In_34);
and U421 (N_421,In_1331,In_1078);
nor U422 (N_422,In_1103,In_198);
xor U423 (N_423,In_457,In_688);
nand U424 (N_424,In_354,In_571);
or U425 (N_425,In_1179,In_999);
nand U426 (N_426,In_1495,In_830);
nand U427 (N_427,In_866,In_583);
xnor U428 (N_428,In_1100,In_815);
and U429 (N_429,In_1113,In_307);
xor U430 (N_430,In_455,In_469);
nand U431 (N_431,In_883,In_845);
nand U432 (N_432,In_233,In_1318);
or U433 (N_433,In_1354,In_843);
nand U434 (N_434,In_536,In_101);
or U435 (N_435,In_1127,In_633);
nor U436 (N_436,In_404,In_1218);
xor U437 (N_437,In_1151,In_1315);
or U438 (N_438,In_1381,In_1038);
nor U439 (N_439,In_985,In_741);
nand U440 (N_440,In_1366,In_371);
nor U441 (N_441,In_187,In_416);
and U442 (N_442,In_68,In_602);
and U443 (N_443,In_21,In_393);
or U444 (N_444,In_334,In_128);
nor U445 (N_445,In_150,In_195);
nor U446 (N_446,In_375,In_522);
and U447 (N_447,In_570,In_499);
and U448 (N_448,In_1225,In_1330);
xor U449 (N_449,In_1309,In_797);
nor U450 (N_450,In_997,In_378);
nand U451 (N_451,In_751,In_501);
and U452 (N_452,In_895,In_544);
or U453 (N_453,In_1307,In_540);
nand U454 (N_454,In_102,In_601);
xor U455 (N_455,In_1471,In_567);
nand U456 (N_456,In_1345,In_615);
nand U457 (N_457,In_1030,In_146);
nand U458 (N_458,In_733,In_343);
or U459 (N_459,In_1241,In_1248);
nor U460 (N_460,In_367,In_470);
xor U461 (N_461,In_20,In_311);
and U462 (N_462,In_1187,In_171);
xnor U463 (N_463,In_541,In_314);
nand U464 (N_464,In_800,In_325);
xnor U465 (N_465,In_1342,In_508);
and U466 (N_466,In_996,In_772);
and U467 (N_467,In_1278,In_881);
nor U468 (N_468,In_261,In_789);
or U469 (N_469,In_568,In_1062);
and U470 (N_470,In_193,In_708);
and U471 (N_471,In_952,In_1442);
xor U472 (N_472,In_219,In_87);
nor U473 (N_473,In_44,In_757);
nor U474 (N_474,In_1094,In_1009);
nand U475 (N_475,In_1026,In_1019);
nand U476 (N_476,In_74,In_520);
and U477 (N_477,In_886,In_441);
or U478 (N_478,In_893,In_1201);
xor U479 (N_479,In_737,In_1256);
nor U480 (N_480,In_816,In_916);
and U481 (N_481,In_585,In_1037);
nor U482 (N_482,In_1067,In_1147);
xor U483 (N_483,In_670,In_869);
or U484 (N_484,In_1377,In_52);
or U485 (N_485,In_433,In_1286);
xor U486 (N_486,In_182,In_235);
nor U487 (N_487,In_1184,In_1000);
nor U488 (N_488,In_732,In_680);
and U489 (N_489,In_249,In_1246);
and U490 (N_490,In_477,In_1039);
xnor U491 (N_491,In_668,In_935);
nand U492 (N_492,In_1073,In_936);
and U493 (N_493,In_738,In_1323);
xor U494 (N_494,In_108,In_867);
and U495 (N_495,In_581,In_73);
nor U496 (N_496,In_776,In_722);
xor U497 (N_497,In_415,In_1052);
nor U498 (N_498,In_401,In_1254);
xor U499 (N_499,In_32,In_1025);
or U500 (N_500,In_578,In_664);
or U501 (N_501,In_60,In_989);
xnor U502 (N_502,In_189,In_1125);
and U503 (N_503,In_674,In_1333);
xor U504 (N_504,In_1304,In_1477);
or U505 (N_505,In_560,In_90);
and U506 (N_506,In_525,In_461);
nor U507 (N_507,In_1137,In_862);
nand U508 (N_508,In_949,In_942);
or U509 (N_509,In_1134,In_712);
and U510 (N_510,In_1292,In_1157);
or U511 (N_511,In_432,In_385);
and U512 (N_512,In_24,In_1372);
or U513 (N_513,In_1166,In_919);
or U514 (N_514,In_794,In_957);
xor U515 (N_515,In_1374,In_1133);
xnor U516 (N_516,In_745,In_648);
nand U517 (N_517,In_887,In_281);
nor U518 (N_518,In_1123,In_10);
nand U519 (N_519,In_655,In_661);
xor U520 (N_520,In_702,In_43);
xnor U521 (N_521,In_1406,In_1459);
or U522 (N_522,In_295,In_672);
nor U523 (N_523,In_875,In_963);
nor U524 (N_524,In_734,In_660);
nor U525 (N_525,In_1474,In_563);
or U526 (N_526,In_1003,In_1491);
nand U527 (N_527,In_852,In_1183);
xnor U528 (N_528,In_994,In_925);
xnor U529 (N_529,In_780,In_1095);
nand U530 (N_530,In_192,In_1066);
or U531 (N_531,In_1328,In_1403);
and U532 (N_532,In_523,In_59);
nand U533 (N_533,In_255,In_1081);
nor U534 (N_534,In_1172,In_1082);
or U535 (N_535,In_700,In_112);
nand U536 (N_536,In_1384,In_75);
or U537 (N_537,In_649,In_1339);
xor U538 (N_538,In_1267,In_1453);
xnor U539 (N_539,In_139,In_1022);
xnor U540 (N_540,In_253,In_703);
xnor U541 (N_541,In_1222,In_1437);
and U542 (N_542,In_319,In_727);
nand U543 (N_543,In_36,In_859);
nand U544 (N_544,In_1083,In_496);
nor U545 (N_545,In_1409,In_795);
xnor U546 (N_546,In_1401,In_1148);
and U547 (N_547,In_1430,In_1362);
nand U548 (N_548,In_316,In_945);
or U549 (N_549,In_216,In_1483);
nor U550 (N_550,In_580,In_206);
and U551 (N_551,In_1164,In_277);
nor U552 (N_552,In_1035,In_41);
and U553 (N_553,In_1057,In_1263);
or U554 (N_554,In_914,In_437);
xnor U555 (N_555,In_781,In_292);
or U556 (N_556,In_659,In_927);
nand U557 (N_557,In_970,In_907);
xnor U558 (N_558,In_1322,In_186);
nor U559 (N_559,In_272,In_1460);
xor U560 (N_560,In_390,In_598);
nand U561 (N_561,In_793,In_836);
nor U562 (N_562,In_1251,In_144);
xnor U563 (N_563,In_1360,In_519);
nand U564 (N_564,In_714,In_1398);
or U565 (N_565,In_1058,In_1071);
nand U566 (N_566,In_624,In_84);
xnor U567 (N_567,In_116,In_86);
and U568 (N_568,In_1107,In_1351);
or U569 (N_569,In_562,In_62);
nor U570 (N_570,In_1208,In_420);
or U571 (N_571,In_511,In_503);
or U572 (N_572,In_1428,In_929);
nand U573 (N_573,In_476,In_376);
nand U574 (N_574,In_762,In_719);
xor U575 (N_575,In_16,In_1108);
nand U576 (N_576,In_973,In_819);
nor U577 (N_577,In_591,In_810);
xnor U578 (N_578,In_842,In_984);
nand U579 (N_579,In_479,In_1033);
nand U580 (N_580,In_731,In_1348);
or U581 (N_581,In_626,In_1139);
nor U582 (N_582,In_871,In_928);
xnor U583 (N_583,In_517,In_528);
nor U584 (N_584,In_848,In_81);
or U585 (N_585,In_172,In_1);
or U586 (N_586,In_115,In_959);
xor U587 (N_587,In_513,In_1337);
nand U588 (N_588,In_308,In_538);
nor U589 (N_589,In_424,In_1221);
xnor U590 (N_590,In_431,In_1150);
and U591 (N_591,In_234,In_383);
xor U592 (N_592,In_66,In_1302);
nand U593 (N_593,In_1298,In_524);
nor U594 (N_594,In_121,In_1274);
nand U595 (N_595,In_419,In_698);
or U596 (N_596,In_160,In_1283);
xor U597 (N_597,In_77,In_944);
nor U598 (N_598,In_637,In_111);
and U599 (N_599,In_123,In_557);
nor U600 (N_600,In_1340,In_608);
nor U601 (N_601,In_199,In_636);
or U602 (N_602,In_777,In_183);
and U603 (N_603,In_1464,In_434);
xnor U604 (N_604,In_1435,In_926);
nor U605 (N_605,In_611,In_188);
xnor U606 (N_606,In_1136,In_1358);
xnor U607 (N_607,In_1482,In_620);
xor U608 (N_608,In_271,In_1216);
nor U609 (N_609,In_300,In_127);
nor U610 (N_610,In_879,In_50);
and U611 (N_611,In_1145,In_223);
nor U612 (N_612,In_894,In_1223);
or U613 (N_613,In_1235,In_279);
nand U614 (N_614,In_756,In_264);
nand U615 (N_615,In_204,In_113);
xor U616 (N_616,In_1361,In_612);
xor U617 (N_617,In_1144,In_443);
nand U618 (N_618,In_1065,In_278);
or U619 (N_619,In_1191,In_874);
nand U620 (N_620,In_442,In_1295);
nand U621 (N_621,In_33,In_103);
nor U622 (N_622,In_587,In_976);
nand U623 (N_623,In_51,In_609);
xnor U624 (N_624,In_1004,In_324);
and U625 (N_625,In_518,In_599);
nor U626 (N_626,In_403,In_1089);
or U627 (N_627,In_1407,In_1385);
nor U628 (N_628,In_622,In_1194);
nor U629 (N_629,In_244,In_1093);
nor U630 (N_630,In_349,In_1122);
nand U631 (N_631,In_983,In_1226);
nand U632 (N_632,In_766,In_71);
xnor U633 (N_633,In_462,In_951);
and U634 (N_634,In_357,In_1101);
or U635 (N_635,In_1421,In_1152);
nand U636 (N_636,In_310,In_1443);
xnor U637 (N_637,In_2,In_823);
xor U638 (N_638,In_1068,In_377);
nor U639 (N_639,In_638,In_877);
and U640 (N_640,In_941,In_586);
or U641 (N_641,In_148,In_436);
and U642 (N_642,In_1480,In_1087);
xnor U643 (N_643,In_1024,In_977);
xor U644 (N_644,In_409,In_1002);
nor U645 (N_645,In_110,In_801);
xnor U646 (N_646,In_251,In_1426);
nand U647 (N_647,In_299,In_1289);
xnor U648 (N_648,In_226,In_790);
xnor U649 (N_649,In_1193,In_413);
nor U650 (N_650,In_1393,In_555);
and U651 (N_651,In_918,In_1200);
or U652 (N_652,In_937,In_912);
nand U653 (N_653,In_313,In_507);
and U654 (N_654,In_1117,In_35);
xor U655 (N_655,In_350,In_93);
nor U656 (N_656,In_1104,In_1311);
nor U657 (N_657,In_840,In_381);
or U658 (N_658,In_500,In_54);
xor U659 (N_659,In_228,In_149);
nor U660 (N_660,In_546,In_1418);
and U661 (N_661,In_613,In_882);
or U662 (N_662,In_717,In_654);
or U663 (N_663,In_950,In_992);
nor U664 (N_664,In_773,In_909);
nor U665 (N_665,In_553,In_214);
or U666 (N_666,In_398,In_297);
nor U667 (N_667,In_430,In_955);
or U668 (N_668,In_1387,In_282);
and U669 (N_669,In_850,In_891);
or U670 (N_670,In_417,In_407);
xnor U671 (N_671,In_8,In_1096);
nand U672 (N_672,In_1059,In_1064);
nor U673 (N_673,In_129,In_335);
or U674 (N_674,In_767,In_57);
nor U675 (N_675,In_1290,In_880);
nor U676 (N_676,In_844,In_239);
nor U677 (N_677,In_1367,In_841);
xnor U678 (N_678,In_687,In_1486);
nand U679 (N_679,In_184,In_817);
and U680 (N_680,In_1233,In_356);
or U681 (N_681,In_783,In_368);
or U682 (N_682,In_394,In_896);
and U683 (N_683,In_227,In_237);
nand U684 (N_684,In_1259,In_91);
and U685 (N_685,In_579,In_747);
and U686 (N_686,In_218,In_735);
nand U687 (N_687,In_946,In_701);
and U688 (N_688,In_1255,In_746);
nand U689 (N_689,In_589,In_391);
or U690 (N_690,In_837,In_200);
nand U691 (N_691,In_1070,In_379);
nor U692 (N_692,In_1310,In_650);
and U693 (N_693,In_998,In_286);
nor U694 (N_694,In_494,In_975);
nand U695 (N_695,In_632,In_1373);
nor U696 (N_696,In_807,In_849);
and U697 (N_697,In_1210,In_1149);
nand U698 (N_698,In_788,In_94);
or U699 (N_699,In_463,In_545);
or U700 (N_700,In_603,In_605);
or U701 (N_701,In_502,In_152);
or U702 (N_702,In_483,In_1313);
and U703 (N_703,In_322,In_15);
xnor U704 (N_704,In_1308,In_1027);
nand U705 (N_705,In_721,In_250);
nand U706 (N_706,In_336,In_954);
xor U707 (N_707,In_932,In_820);
nand U708 (N_708,In_1319,In_631);
and U709 (N_709,In_754,In_1045);
or U710 (N_710,In_11,In_1209);
or U711 (N_711,In_725,In_1143);
and U712 (N_712,In_1413,In_495);
nor U713 (N_713,In_930,In_685);
nor U714 (N_714,In_1245,In_1488);
nand U715 (N_715,In_254,In_133);
and U716 (N_716,In_748,In_1181);
and U717 (N_717,In_427,In_1163);
or U718 (N_718,In_515,In_151);
xor U719 (N_719,In_595,In_1072);
and U720 (N_720,In_628,In_673);
and U721 (N_721,In_1479,In_814);
nand U722 (N_722,In_671,In_851);
and U723 (N_723,In_922,In_924);
or U724 (N_724,In_779,In_257);
xnor U725 (N_725,In_221,In_1046);
nand U726 (N_726,In_446,In_131);
and U727 (N_727,In_986,In_1465);
xor U728 (N_728,In_331,In_274);
nand U729 (N_729,In_573,In_194);
nand U730 (N_730,In_938,In_1432);
and U731 (N_731,In_1008,In_556);
xnor U732 (N_732,In_458,In_1445);
nor U733 (N_733,In_1476,In_288);
nor U734 (N_734,In_1086,In_645);
and U735 (N_735,In_359,In_482);
or U736 (N_736,In_1010,In_289);
or U737 (N_737,In_201,In_1063);
or U738 (N_738,In_332,In_1023);
nand U739 (N_739,In_481,In_1161);
nor U740 (N_740,In_321,In_1203);
xnor U741 (N_741,In_1450,In_492);
and U742 (N_742,In_743,In_1227);
nand U743 (N_743,In_1462,In_884);
or U744 (N_744,In_854,In_1279);
and U745 (N_745,In_418,In_179);
nand U746 (N_746,In_604,In_1291);
nor U747 (N_747,In_1014,In_1084);
nand U748 (N_748,In_1489,In_530);
nand U749 (N_749,In_389,In_749);
nand U750 (N_750,In_295,In_956);
nand U751 (N_751,In_790,In_1484);
and U752 (N_752,In_656,In_753);
or U753 (N_753,In_271,In_1443);
nor U754 (N_754,In_759,In_1405);
xor U755 (N_755,In_854,In_219);
xnor U756 (N_756,In_659,In_792);
or U757 (N_757,In_482,In_521);
nor U758 (N_758,In_278,In_1448);
xnor U759 (N_759,In_796,In_388);
xor U760 (N_760,In_113,In_571);
xnor U761 (N_761,In_523,In_1282);
nor U762 (N_762,In_1468,In_284);
or U763 (N_763,In_639,In_1469);
and U764 (N_764,In_770,In_650);
and U765 (N_765,In_522,In_1268);
nor U766 (N_766,In_1023,In_1164);
and U767 (N_767,In_1110,In_1396);
or U768 (N_768,In_980,In_1423);
nand U769 (N_769,In_759,In_49);
xor U770 (N_770,In_607,In_994);
xor U771 (N_771,In_36,In_779);
and U772 (N_772,In_560,In_892);
and U773 (N_773,In_286,In_5);
and U774 (N_774,In_281,In_546);
xnor U775 (N_775,In_535,In_88);
and U776 (N_776,In_1204,In_750);
or U777 (N_777,In_330,In_1372);
nand U778 (N_778,In_74,In_1318);
xnor U779 (N_779,In_1080,In_67);
nor U780 (N_780,In_529,In_36);
xnor U781 (N_781,In_1113,In_1268);
nand U782 (N_782,In_1332,In_1228);
nand U783 (N_783,In_816,In_1469);
or U784 (N_784,In_823,In_1355);
or U785 (N_785,In_493,In_901);
and U786 (N_786,In_616,In_198);
and U787 (N_787,In_284,In_779);
xor U788 (N_788,In_1341,In_171);
xnor U789 (N_789,In_1232,In_1238);
nand U790 (N_790,In_1239,In_469);
nor U791 (N_791,In_316,In_994);
nor U792 (N_792,In_1337,In_834);
nor U793 (N_793,In_908,In_981);
and U794 (N_794,In_384,In_406);
or U795 (N_795,In_1387,In_842);
xnor U796 (N_796,In_575,In_292);
xor U797 (N_797,In_1074,In_516);
nor U798 (N_798,In_1378,In_272);
nor U799 (N_799,In_774,In_1440);
nand U800 (N_800,In_344,In_901);
xnor U801 (N_801,In_940,In_1284);
or U802 (N_802,In_241,In_225);
nand U803 (N_803,In_858,In_1230);
nand U804 (N_804,In_929,In_574);
nor U805 (N_805,In_1213,In_885);
xor U806 (N_806,In_936,In_452);
nand U807 (N_807,In_703,In_1013);
xnor U808 (N_808,In_480,In_668);
nor U809 (N_809,In_850,In_277);
nand U810 (N_810,In_914,In_18);
nor U811 (N_811,In_623,In_1392);
nand U812 (N_812,In_1231,In_236);
nor U813 (N_813,In_1130,In_39);
or U814 (N_814,In_404,In_591);
nor U815 (N_815,In_1377,In_454);
nor U816 (N_816,In_850,In_474);
xnor U817 (N_817,In_823,In_552);
nand U818 (N_818,In_1162,In_1393);
xor U819 (N_819,In_590,In_127);
xor U820 (N_820,In_1459,In_1190);
or U821 (N_821,In_983,In_349);
and U822 (N_822,In_1115,In_581);
or U823 (N_823,In_1432,In_1266);
nand U824 (N_824,In_577,In_1);
nor U825 (N_825,In_183,In_1380);
nand U826 (N_826,In_1154,In_1120);
or U827 (N_827,In_1334,In_316);
xor U828 (N_828,In_277,In_308);
xor U829 (N_829,In_415,In_65);
or U830 (N_830,In_59,In_381);
or U831 (N_831,In_440,In_767);
nor U832 (N_832,In_1243,In_633);
or U833 (N_833,In_363,In_901);
nand U834 (N_834,In_822,In_100);
or U835 (N_835,In_115,In_557);
xor U836 (N_836,In_890,In_1315);
xor U837 (N_837,In_38,In_1449);
or U838 (N_838,In_215,In_251);
xnor U839 (N_839,In_752,In_1277);
and U840 (N_840,In_1491,In_995);
and U841 (N_841,In_858,In_815);
xor U842 (N_842,In_1040,In_1378);
or U843 (N_843,In_666,In_266);
and U844 (N_844,In_467,In_911);
and U845 (N_845,In_1389,In_1068);
nor U846 (N_846,In_1463,In_328);
or U847 (N_847,In_938,In_859);
and U848 (N_848,In_627,In_1360);
and U849 (N_849,In_1433,In_637);
and U850 (N_850,In_317,In_379);
nand U851 (N_851,In_217,In_573);
or U852 (N_852,In_866,In_1335);
nor U853 (N_853,In_269,In_504);
and U854 (N_854,In_439,In_1187);
xnor U855 (N_855,In_1428,In_425);
nor U856 (N_856,In_878,In_1036);
nand U857 (N_857,In_528,In_1225);
nand U858 (N_858,In_1061,In_572);
xnor U859 (N_859,In_650,In_555);
xor U860 (N_860,In_249,In_254);
or U861 (N_861,In_871,In_452);
or U862 (N_862,In_1075,In_310);
nand U863 (N_863,In_808,In_992);
xnor U864 (N_864,In_944,In_606);
xor U865 (N_865,In_76,In_766);
and U866 (N_866,In_353,In_859);
and U867 (N_867,In_1291,In_318);
and U868 (N_868,In_439,In_320);
xor U869 (N_869,In_184,In_1001);
xor U870 (N_870,In_839,In_1391);
nor U871 (N_871,In_1077,In_408);
or U872 (N_872,In_372,In_1139);
nor U873 (N_873,In_873,In_598);
or U874 (N_874,In_1048,In_1132);
nand U875 (N_875,In_996,In_1330);
xor U876 (N_876,In_919,In_990);
nor U877 (N_877,In_1171,In_482);
xor U878 (N_878,In_1119,In_658);
or U879 (N_879,In_943,In_466);
nor U880 (N_880,In_1469,In_1089);
or U881 (N_881,In_777,In_536);
nand U882 (N_882,In_1046,In_457);
and U883 (N_883,In_1211,In_997);
or U884 (N_884,In_1063,In_794);
nand U885 (N_885,In_1222,In_305);
nor U886 (N_886,In_242,In_386);
or U887 (N_887,In_1067,In_79);
and U888 (N_888,In_1144,In_190);
nand U889 (N_889,In_1250,In_737);
or U890 (N_890,In_1447,In_162);
nand U891 (N_891,In_848,In_726);
xor U892 (N_892,In_186,In_1116);
nand U893 (N_893,In_1011,In_1156);
xor U894 (N_894,In_551,In_594);
xnor U895 (N_895,In_762,In_211);
nor U896 (N_896,In_467,In_1043);
or U897 (N_897,In_103,In_53);
nand U898 (N_898,In_1268,In_491);
nand U899 (N_899,In_919,In_79);
nor U900 (N_900,In_1026,In_878);
or U901 (N_901,In_1069,In_1257);
xor U902 (N_902,In_1182,In_712);
nand U903 (N_903,In_992,In_86);
xor U904 (N_904,In_762,In_549);
xnor U905 (N_905,In_1405,In_347);
nor U906 (N_906,In_1008,In_746);
and U907 (N_907,In_1408,In_928);
nor U908 (N_908,In_175,In_722);
and U909 (N_909,In_1098,In_757);
and U910 (N_910,In_793,In_1170);
xnor U911 (N_911,In_827,In_1489);
nand U912 (N_912,In_375,In_1312);
xnor U913 (N_913,In_1,In_699);
xnor U914 (N_914,In_359,In_1328);
xor U915 (N_915,In_629,In_504);
xnor U916 (N_916,In_1373,In_2);
and U917 (N_917,In_792,In_1309);
and U918 (N_918,In_760,In_771);
and U919 (N_919,In_451,In_1422);
nand U920 (N_920,In_1250,In_193);
and U921 (N_921,In_1243,In_587);
or U922 (N_922,In_196,In_144);
nand U923 (N_923,In_1002,In_996);
and U924 (N_924,In_657,In_1220);
or U925 (N_925,In_1338,In_1187);
xor U926 (N_926,In_548,In_96);
and U927 (N_927,In_955,In_1318);
nand U928 (N_928,In_110,In_1347);
nand U929 (N_929,In_1456,In_1346);
nor U930 (N_930,In_592,In_164);
xnor U931 (N_931,In_158,In_299);
xnor U932 (N_932,In_1168,In_131);
nor U933 (N_933,In_323,In_955);
nor U934 (N_934,In_187,In_159);
xor U935 (N_935,In_342,In_981);
or U936 (N_936,In_437,In_115);
and U937 (N_937,In_861,In_972);
nor U938 (N_938,In_148,In_191);
nand U939 (N_939,In_1333,In_300);
and U940 (N_940,In_1368,In_1422);
and U941 (N_941,In_437,In_743);
nor U942 (N_942,In_813,In_22);
and U943 (N_943,In_216,In_1272);
nand U944 (N_944,In_501,In_1370);
nand U945 (N_945,In_1205,In_113);
nand U946 (N_946,In_1422,In_500);
xnor U947 (N_947,In_1165,In_581);
nand U948 (N_948,In_884,In_213);
or U949 (N_949,In_582,In_987);
xnor U950 (N_950,In_762,In_242);
and U951 (N_951,In_1122,In_1098);
and U952 (N_952,In_1117,In_561);
nor U953 (N_953,In_52,In_1168);
and U954 (N_954,In_1219,In_391);
nand U955 (N_955,In_1299,In_929);
nor U956 (N_956,In_288,In_699);
nor U957 (N_957,In_92,In_894);
xor U958 (N_958,In_881,In_810);
xor U959 (N_959,In_334,In_1182);
and U960 (N_960,In_404,In_575);
or U961 (N_961,In_171,In_1064);
nor U962 (N_962,In_1166,In_791);
and U963 (N_963,In_1319,In_982);
or U964 (N_964,In_1334,In_91);
xor U965 (N_965,In_917,In_1062);
or U966 (N_966,In_208,In_1127);
and U967 (N_967,In_607,In_924);
xor U968 (N_968,In_786,In_1339);
or U969 (N_969,In_626,In_1049);
and U970 (N_970,In_822,In_906);
nand U971 (N_971,In_433,In_467);
nand U972 (N_972,In_1098,In_1458);
or U973 (N_973,In_1278,In_109);
nand U974 (N_974,In_422,In_1424);
or U975 (N_975,In_1495,In_197);
or U976 (N_976,In_448,In_427);
nand U977 (N_977,In_413,In_1459);
nor U978 (N_978,In_796,In_1115);
nand U979 (N_979,In_1260,In_1030);
or U980 (N_980,In_630,In_527);
and U981 (N_981,In_205,In_1030);
nand U982 (N_982,In_1026,In_303);
nor U983 (N_983,In_1402,In_1467);
nand U984 (N_984,In_702,In_1350);
or U985 (N_985,In_52,In_826);
or U986 (N_986,In_1148,In_670);
nor U987 (N_987,In_357,In_1361);
nand U988 (N_988,In_1048,In_1310);
or U989 (N_989,In_1411,In_932);
or U990 (N_990,In_578,In_939);
or U991 (N_991,In_299,In_1365);
nand U992 (N_992,In_39,In_632);
or U993 (N_993,In_186,In_1024);
xor U994 (N_994,In_377,In_1307);
xor U995 (N_995,In_153,In_57);
nand U996 (N_996,In_1124,In_564);
xor U997 (N_997,In_349,In_832);
or U998 (N_998,In_467,In_365);
nand U999 (N_999,In_444,In_1454);
xor U1000 (N_1000,In_271,In_1109);
or U1001 (N_1001,In_1087,In_1202);
xor U1002 (N_1002,In_1014,In_267);
nand U1003 (N_1003,In_1392,In_1337);
xor U1004 (N_1004,In_1016,In_1034);
nor U1005 (N_1005,In_1439,In_899);
nor U1006 (N_1006,In_369,In_1064);
nand U1007 (N_1007,In_834,In_567);
or U1008 (N_1008,In_1253,In_823);
nor U1009 (N_1009,In_695,In_1089);
or U1010 (N_1010,In_314,In_1129);
xnor U1011 (N_1011,In_761,In_671);
and U1012 (N_1012,In_860,In_1436);
and U1013 (N_1013,In_1068,In_1250);
and U1014 (N_1014,In_1085,In_449);
or U1015 (N_1015,In_746,In_1486);
and U1016 (N_1016,In_210,In_304);
or U1017 (N_1017,In_1238,In_1247);
nand U1018 (N_1018,In_235,In_580);
and U1019 (N_1019,In_1138,In_177);
nand U1020 (N_1020,In_549,In_1164);
nand U1021 (N_1021,In_1448,In_1366);
or U1022 (N_1022,In_1313,In_596);
xor U1023 (N_1023,In_905,In_1187);
and U1024 (N_1024,In_810,In_312);
or U1025 (N_1025,In_790,In_433);
or U1026 (N_1026,In_1039,In_266);
and U1027 (N_1027,In_1333,In_737);
or U1028 (N_1028,In_1186,In_1298);
xnor U1029 (N_1029,In_771,In_1338);
nand U1030 (N_1030,In_244,In_1339);
xor U1031 (N_1031,In_1112,In_1190);
nand U1032 (N_1032,In_656,In_168);
or U1033 (N_1033,In_893,In_273);
and U1034 (N_1034,In_1073,In_583);
nand U1035 (N_1035,In_1256,In_267);
nor U1036 (N_1036,In_1374,In_901);
and U1037 (N_1037,In_1341,In_445);
nor U1038 (N_1038,In_275,In_776);
nor U1039 (N_1039,In_228,In_848);
xor U1040 (N_1040,In_746,In_967);
nand U1041 (N_1041,In_1082,In_1033);
or U1042 (N_1042,In_75,In_209);
and U1043 (N_1043,In_775,In_340);
or U1044 (N_1044,In_963,In_1240);
and U1045 (N_1045,In_678,In_226);
nand U1046 (N_1046,In_144,In_486);
or U1047 (N_1047,In_1295,In_851);
and U1048 (N_1048,In_139,In_115);
nor U1049 (N_1049,In_980,In_1031);
nand U1050 (N_1050,In_860,In_1247);
nand U1051 (N_1051,In_739,In_1488);
nand U1052 (N_1052,In_1186,In_234);
and U1053 (N_1053,In_1296,In_1245);
and U1054 (N_1054,In_1033,In_1437);
nor U1055 (N_1055,In_1362,In_1372);
nor U1056 (N_1056,In_1035,In_93);
or U1057 (N_1057,In_1429,In_255);
nor U1058 (N_1058,In_437,In_515);
nand U1059 (N_1059,In_1167,In_10);
and U1060 (N_1060,In_323,In_303);
and U1061 (N_1061,In_479,In_1292);
or U1062 (N_1062,In_1252,In_20);
or U1063 (N_1063,In_1445,In_869);
xor U1064 (N_1064,In_594,In_314);
nor U1065 (N_1065,In_1325,In_1304);
and U1066 (N_1066,In_1384,In_436);
nor U1067 (N_1067,In_861,In_998);
and U1068 (N_1068,In_1243,In_1428);
and U1069 (N_1069,In_1309,In_253);
nor U1070 (N_1070,In_229,In_149);
nand U1071 (N_1071,In_567,In_628);
nor U1072 (N_1072,In_287,In_180);
xor U1073 (N_1073,In_700,In_1445);
nor U1074 (N_1074,In_1319,In_1288);
nor U1075 (N_1075,In_231,In_1117);
and U1076 (N_1076,In_924,In_740);
and U1077 (N_1077,In_826,In_343);
and U1078 (N_1078,In_1002,In_1018);
nand U1079 (N_1079,In_586,In_695);
nand U1080 (N_1080,In_92,In_1106);
and U1081 (N_1081,In_1205,In_126);
xnor U1082 (N_1082,In_682,In_208);
xnor U1083 (N_1083,In_407,In_1098);
or U1084 (N_1084,In_124,In_601);
xnor U1085 (N_1085,In_519,In_227);
or U1086 (N_1086,In_1168,In_355);
nand U1087 (N_1087,In_35,In_1328);
nand U1088 (N_1088,In_271,In_717);
nand U1089 (N_1089,In_624,In_283);
xnor U1090 (N_1090,In_1452,In_352);
or U1091 (N_1091,In_1420,In_371);
nand U1092 (N_1092,In_273,In_662);
nor U1093 (N_1093,In_1329,In_944);
nor U1094 (N_1094,In_1442,In_660);
and U1095 (N_1095,In_1163,In_1310);
or U1096 (N_1096,In_390,In_1303);
and U1097 (N_1097,In_1408,In_126);
xnor U1098 (N_1098,In_355,In_1102);
nor U1099 (N_1099,In_1390,In_1064);
nand U1100 (N_1100,In_51,In_958);
and U1101 (N_1101,In_1461,In_1095);
nand U1102 (N_1102,In_372,In_1172);
or U1103 (N_1103,In_866,In_773);
and U1104 (N_1104,In_1195,In_440);
and U1105 (N_1105,In_995,In_765);
and U1106 (N_1106,In_124,In_1151);
or U1107 (N_1107,In_139,In_414);
nor U1108 (N_1108,In_307,In_898);
nand U1109 (N_1109,In_835,In_643);
nor U1110 (N_1110,In_777,In_724);
xnor U1111 (N_1111,In_837,In_814);
nand U1112 (N_1112,In_1232,In_340);
nand U1113 (N_1113,In_1368,In_901);
or U1114 (N_1114,In_139,In_768);
xor U1115 (N_1115,In_536,In_697);
xnor U1116 (N_1116,In_1186,In_95);
nand U1117 (N_1117,In_164,In_170);
or U1118 (N_1118,In_639,In_1030);
or U1119 (N_1119,In_173,In_1404);
and U1120 (N_1120,In_1054,In_917);
and U1121 (N_1121,In_836,In_11);
or U1122 (N_1122,In_617,In_1052);
and U1123 (N_1123,In_481,In_474);
xor U1124 (N_1124,In_966,In_1067);
or U1125 (N_1125,In_22,In_852);
nor U1126 (N_1126,In_940,In_368);
and U1127 (N_1127,In_928,In_854);
nor U1128 (N_1128,In_1257,In_237);
or U1129 (N_1129,In_503,In_1134);
nor U1130 (N_1130,In_1427,In_791);
or U1131 (N_1131,In_565,In_428);
xor U1132 (N_1132,In_377,In_1442);
xnor U1133 (N_1133,In_598,In_1385);
nor U1134 (N_1134,In_50,In_195);
xor U1135 (N_1135,In_212,In_752);
nor U1136 (N_1136,In_705,In_1470);
xor U1137 (N_1137,In_991,In_1352);
and U1138 (N_1138,In_515,In_290);
and U1139 (N_1139,In_100,In_409);
nand U1140 (N_1140,In_226,In_929);
and U1141 (N_1141,In_726,In_352);
and U1142 (N_1142,In_736,In_810);
or U1143 (N_1143,In_1287,In_1384);
xnor U1144 (N_1144,In_641,In_1475);
xnor U1145 (N_1145,In_589,In_536);
nor U1146 (N_1146,In_1456,In_599);
or U1147 (N_1147,In_1387,In_461);
or U1148 (N_1148,In_1010,In_663);
xor U1149 (N_1149,In_738,In_1040);
nand U1150 (N_1150,In_201,In_1420);
and U1151 (N_1151,In_979,In_976);
or U1152 (N_1152,In_967,In_81);
nand U1153 (N_1153,In_1433,In_515);
or U1154 (N_1154,In_768,In_355);
and U1155 (N_1155,In_1259,In_757);
nand U1156 (N_1156,In_567,In_369);
and U1157 (N_1157,In_692,In_633);
and U1158 (N_1158,In_1221,In_1460);
or U1159 (N_1159,In_1029,In_691);
nand U1160 (N_1160,In_149,In_1450);
and U1161 (N_1161,In_1475,In_505);
xnor U1162 (N_1162,In_382,In_92);
and U1163 (N_1163,In_420,In_190);
nor U1164 (N_1164,In_1235,In_575);
nand U1165 (N_1165,In_1451,In_759);
nor U1166 (N_1166,In_445,In_970);
nor U1167 (N_1167,In_231,In_248);
and U1168 (N_1168,In_632,In_276);
nor U1169 (N_1169,In_1133,In_1149);
nor U1170 (N_1170,In_1405,In_939);
nor U1171 (N_1171,In_944,In_1403);
nand U1172 (N_1172,In_756,In_1439);
xor U1173 (N_1173,In_76,In_1222);
nand U1174 (N_1174,In_715,In_1081);
nor U1175 (N_1175,In_578,In_388);
xor U1176 (N_1176,In_867,In_597);
nand U1177 (N_1177,In_482,In_766);
nand U1178 (N_1178,In_376,In_1156);
nor U1179 (N_1179,In_1433,In_309);
nand U1180 (N_1180,In_1192,In_1241);
nor U1181 (N_1181,In_1106,In_1258);
or U1182 (N_1182,In_817,In_909);
nor U1183 (N_1183,In_238,In_740);
or U1184 (N_1184,In_1039,In_308);
nand U1185 (N_1185,In_1427,In_1290);
and U1186 (N_1186,In_624,In_1138);
or U1187 (N_1187,In_1309,In_848);
xor U1188 (N_1188,In_548,In_909);
nor U1189 (N_1189,In_468,In_1463);
or U1190 (N_1190,In_1364,In_139);
nor U1191 (N_1191,In_73,In_193);
nor U1192 (N_1192,In_1081,In_654);
nor U1193 (N_1193,In_1127,In_1242);
nor U1194 (N_1194,In_932,In_100);
nor U1195 (N_1195,In_62,In_639);
and U1196 (N_1196,In_327,In_1400);
and U1197 (N_1197,In_969,In_1392);
xnor U1198 (N_1198,In_1288,In_1378);
nor U1199 (N_1199,In_1198,In_553);
and U1200 (N_1200,In_1029,In_242);
nor U1201 (N_1201,In_431,In_1139);
or U1202 (N_1202,In_743,In_1378);
or U1203 (N_1203,In_1418,In_113);
xor U1204 (N_1204,In_461,In_193);
or U1205 (N_1205,In_633,In_195);
nor U1206 (N_1206,In_1387,In_444);
xor U1207 (N_1207,In_621,In_525);
nand U1208 (N_1208,In_559,In_79);
or U1209 (N_1209,In_679,In_1374);
and U1210 (N_1210,In_912,In_1220);
xnor U1211 (N_1211,In_612,In_313);
and U1212 (N_1212,In_1410,In_1471);
nor U1213 (N_1213,In_718,In_615);
nor U1214 (N_1214,In_1319,In_361);
nor U1215 (N_1215,In_228,In_111);
or U1216 (N_1216,In_66,In_143);
nand U1217 (N_1217,In_690,In_931);
and U1218 (N_1218,In_439,In_52);
nand U1219 (N_1219,In_1197,In_1274);
or U1220 (N_1220,In_438,In_587);
and U1221 (N_1221,In_460,In_791);
or U1222 (N_1222,In_491,In_664);
nand U1223 (N_1223,In_259,In_788);
or U1224 (N_1224,In_787,In_220);
nand U1225 (N_1225,In_907,In_692);
or U1226 (N_1226,In_1336,In_322);
nor U1227 (N_1227,In_1239,In_47);
or U1228 (N_1228,In_470,In_1279);
xor U1229 (N_1229,In_459,In_1342);
nand U1230 (N_1230,In_1458,In_1141);
nand U1231 (N_1231,In_751,In_898);
nand U1232 (N_1232,In_928,In_271);
nor U1233 (N_1233,In_188,In_1313);
or U1234 (N_1234,In_726,In_690);
nand U1235 (N_1235,In_567,In_1193);
nand U1236 (N_1236,In_536,In_505);
nand U1237 (N_1237,In_937,In_1477);
nor U1238 (N_1238,In_576,In_593);
and U1239 (N_1239,In_1201,In_956);
nor U1240 (N_1240,In_1350,In_1256);
nor U1241 (N_1241,In_1301,In_1153);
or U1242 (N_1242,In_1406,In_1183);
xnor U1243 (N_1243,In_1052,In_636);
xnor U1244 (N_1244,In_367,In_1133);
nand U1245 (N_1245,In_354,In_66);
and U1246 (N_1246,In_1488,In_962);
xnor U1247 (N_1247,In_913,In_1138);
or U1248 (N_1248,In_844,In_287);
nor U1249 (N_1249,In_552,In_17);
and U1250 (N_1250,In_615,In_1040);
nand U1251 (N_1251,In_1342,In_1092);
nand U1252 (N_1252,In_1248,In_424);
or U1253 (N_1253,In_441,In_578);
xnor U1254 (N_1254,In_1419,In_830);
nor U1255 (N_1255,In_890,In_1129);
xnor U1256 (N_1256,In_1219,In_678);
nand U1257 (N_1257,In_525,In_1367);
and U1258 (N_1258,In_925,In_155);
xnor U1259 (N_1259,In_1203,In_302);
or U1260 (N_1260,In_18,In_458);
xor U1261 (N_1261,In_403,In_460);
xor U1262 (N_1262,In_261,In_94);
or U1263 (N_1263,In_914,In_173);
or U1264 (N_1264,In_172,In_1077);
xor U1265 (N_1265,In_845,In_1075);
nor U1266 (N_1266,In_361,In_1409);
xnor U1267 (N_1267,In_906,In_162);
nor U1268 (N_1268,In_1466,In_1309);
xnor U1269 (N_1269,In_779,In_227);
and U1270 (N_1270,In_532,In_185);
nand U1271 (N_1271,In_1347,In_11);
or U1272 (N_1272,In_169,In_381);
and U1273 (N_1273,In_789,In_1433);
and U1274 (N_1274,In_846,In_1145);
and U1275 (N_1275,In_1135,In_83);
xor U1276 (N_1276,In_1054,In_62);
xor U1277 (N_1277,In_195,In_137);
and U1278 (N_1278,In_278,In_510);
nand U1279 (N_1279,In_24,In_1294);
xnor U1280 (N_1280,In_995,In_1354);
xnor U1281 (N_1281,In_250,In_42);
xor U1282 (N_1282,In_54,In_1471);
nand U1283 (N_1283,In_553,In_869);
and U1284 (N_1284,In_1063,In_646);
nor U1285 (N_1285,In_1165,In_1472);
and U1286 (N_1286,In_1042,In_478);
or U1287 (N_1287,In_41,In_834);
or U1288 (N_1288,In_380,In_256);
xor U1289 (N_1289,In_103,In_353);
or U1290 (N_1290,In_42,In_1022);
and U1291 (N_1291,In_78,In_777);
xnor U1292 (N_1292,In_870,In_646);
or U1293 (N_1293,In_212,In_483);
or U1294 (N_1294,In_203,In_207);
nand U1295 (N_1295,In_613,In_261);
or U1296 (N_1296,In_1277,In_249);
nand U1297 (N_1297,In_298,In_432);
nand U1298 (N_1298,In_1266,In_1475);
xor U1299 (N_1299,In_1246,In_1263);
nor U1300 (N_1300,In_408,In_47);
xor U1301 (N_1301,In_1162,In_1050);
nor U1302 (N_1302,In_1312,In_296);
nand U1303 (N_1303,In_785,In_880);
nand U1304 (N_1304,In_580,In_682);
or U1305 (N_1305,In_870,In_963);
nor U1306 (N_1306,In_802,In_1462);
or U1307 (N_1307,In_1344,In_1395);
or U1308 (N_1308,In_1273,In_596);
nand U1309 (N_1309,In_1341,In_139);
xnor U1310 (N_1310,In_1224,In_153);
xor U1311 (N_1311,In_1296,In_861);
nor U1312 (N_1312,In_1135,In_881);
nor U1313 (N_1313,In_210,In_1185);
xor U1314 (N_1314,In_366,In_1368);
nor U1315 (N_1315,In_911,In_886);
nor U1316 (N_1316,In_1452,In_1382);
nor U1317 (N_1317,In_515,In_251);
nor U1318 (N_1318,In_728,In_1186);
nor U1319 (N_1319,In_1023,In_1038);
nand U1320 (N_1320,In_932,In_1389);
or U1321 (N_1321,In_855,In_617);
and U1322 (N_1322,In_268,In_1301);
nor U1323 (N_1323,In_190,In_72);
and U1324 (N_1324,In_714,In_954);
nand U1325 (N_1325,In_1397,In_11);
xnor U1326 (N_1326,In_1359,In_1196);
xor U1327 (N_1327,In_571,In_426);
nand U1328 (N_1328,In_574,In_954);
nor U1329 (N_1329,In_367,In_1159);
or U1330 (N_1330,In_1360,In_1297);
nand U1331 (N_1331,In_1041,In_1315);
or U1332 (N_1332,In_1018,In_944);
nor U1333 (N_1333,In_140,In_639);
xnor U1334 (N_1334,In_817,In_727);
nand U1335 (N_1335,In_1095,In_154);
or U1336 (N_1336,In_1352,In_1069);
xnor U1337 (N_1337,In_227,In_762);
and U1338 (N_1338,In_1474,In_1398);
or U1339 (N_1339,In_211,In_531);
or U1340 (N_1340,In_848,In_929);
or U1341 (N_1341,In_332,In_343);
or U1342 (N_1342,In_1267,In_920);
nand U1343 (N_1343,In_742,In_1052);
or U1344 (N_1344,In_1050,In_901);
nand U1345 (N_1345,In_405,In_951);
xnor U1346 (N_1346,In_1131,In_1417);
and U1347 (N_1347,In_1230,In_1031);
nand U1348 (N_1348,In_794,In_384);
or U1349 (N_1349,In_848,In_843);
nor U1350 (N_1350,In_793,In_632);
nand U1351 (N_1351,In_223,In_238);
xor U1352 (N_1352,In_473,In_578);
nand U1353 (N_1353,In_678,In_28);
nor U1354 (N_1354,In_1040,In_82);
nand U1355 (N_1355,In_1131,In_1183);
nor U1356 (N_1356,In_907,In_1180);
xnor U1357 (N_1357,In_950,In_988);
nand U1358 (N_1358,In_1240,In_676);
nor U1359 (N_1359,In_1174,In_950);
xor U1360 (N_1360,In_157,In_832);
xnor U1361 (N_1361,In_1076,In_36);
nor U1362 (N_1362,In_1006,In_474);
nor U1363 (N_1363,In_780,In_828);
xor U1364 (N_1364,In_1499,In_890);
xor U1365 (N_1365,In_1247,In_1026);
and U1366 (N_1366,In_1037,In_19);
xnor U1367 (N_1367,In_149,In_42);
nand U1368 (N_1368,In_390,In_1121);
nand U1369 (N_1369,In_225,In_1143);
nor U1370 (N_1370,In_0,In_474);
or U1371 (N_1371,In_257,In_1047);
and U1372 (N_1372,In_324,In_851);
or U1373 (N_1373,In_123,In_874);
and U1374 (N_1374,In_1219,In_53);
or U1375 (N_1375,In_406,In_32);
or U1376 (N_1376,In_1170,In_1487);
or U1377 (N_1377,In_19,In_1105);
nor U1378 (N_1378,In_656,In_1033);
and U1379 (N_1379,In_383,In_1076);
xor U1380 (N_1380,In_648,In_6);
nor U1381 (N_1381,In_195,In_1177);
nand U1382 (N_1382,In_173,In_593);
nand U1383 (N_1383,In_941,In_334);
xnor U1384 (N_1384,In_1015,In_411);
nand U1385 (N_1385,In_1051,In_1346);
xor U1386 (N_1386,In_364,In_1476);
xor U1387 (N_1387,In_1462,In_1002);
nor U1388 (N_1388,In_1421,In_1088);
nor U1389 (N_1389,In_18,In_1214);
nor U1390 (N_1390,In_935,In_1120);
and U1391 (N_1391,In_1312,In_4);
and U1392 (N_1392,In_618,In_1262);
nand U1393 (N_1393,In_67,In_1488);
and U1394 (N_1394,In_949,In_937);
and U1395 (N_1395,In_308,In_1326);
and U1396 (N_1396,In_324,In_1055);
or U1397 (N_1397,In_1008,In_196);
or U1398 (N_1398,In_1269,In_1075);
nor U1399 (N_1399,In_1388,In_1448);
xnor U1400 (N_1400,In_1236,In_1064);
and U1401 (N_1401,In_1207,In_589);
nand U1402 (N_1402,In_691,In_273);
xor U1403 (N_1403,In_443,In_456);
and U1404 (N_1404,In_199,In_961);
xor U1405 (N_1405,In_307,In_454);
or U1406 (N_1406,In_762,In_962);
nor U1407 (N_1407,In_450,In_773);
xor U1408 (N_1408,In_62,In_1366);
or U1409 (N_1409,In_227,In_452);
nor U1410 (N_1410,In_1282,In_673);
and U1411 (N_1411,In_1032,In_387);
nand U1412 (N_1412,In_137,In_94);
and U1413 (N_1413,In_1249,In_756);
nand U1414 (N_1414,In_717,In_1366);
xnor U1415 (N_1415,In_412,In_607);
and U1416 (N_1416,In_399,In_1113);
xnor U1417 (N_1417,In_934,In_1452);
nand U1418 (N_1418,In_1064,In_504);
nand U1419 (N_1419,In_346,In_145);
or U1420 (N_1420,In_1311,In_1478);
nor U1421 (N_1421,In_1105,In_861);
and U1422 (N_1422,In_398,In_323);
nand U1423 (N_1423,In_265,In_335);
nand U1424 (N_1424,In_1174,In_778);
xnor U1425 (N_1425,In_1154,In_520);
nor U1426 (N_1426,In_693,In_523);
or U1427 (N_1427,In_660,In_3);
nand U1428 (N_1428,In_1439,In_1075);
nand U1429 (N_1429,In_398,In_504);
or U1430 (N_1430,In_329,In_1131);
xor U1431 (N_1431,In_459,In_1208);
xnor U1432 (N_1432,In_949,In_18);
xnor U1433 (N_1433,In_1007,In_95);
nor U1434 (N_1434,In_339,In_1076);
nor U1435 (N_1435,In_610,In_1153);
xnor U1436 (N_1436,In_758,In_412);
xor U1437 (N_1437,In_248,In_323);
xnor U1438 (N_1438,In_1087,In_29);
and U1439 (N_1439,In_120,In_1141);
or U1440 (N_1440,In_1337,In_93);
and U1441 (N_1441,In_470,In_1165);
and U1442 (N_1442,In_130,In_1272);
xnor U1443 (N_1443,In_1317,In_397);
and U1444 (N_1444,In_47,In_1191);
and U1445 (N_1445,In_52,In_548);
xor U1446 (N_1446,In_1171,In_311);
or U1447 (N_1447,In_737,In_945);
and U1448 (N_1448,In_758,In_260);
xnor U1449 (N_1449,In_671,In_467);
nor U1450 (N_1450,In_991,In_1200);
and U1451 (N_1451,In_594,In_1467);
nand U1452 (N_1452,In_847,In_1311);
or U1453 (N_1453,In_1267,In_1409);
nand U1454 (N_1454,In_1237,In_1085);
xor U1455 (N_1455,In_1083,In_1325);
nand U1456 (N_1456,In_1486,In_639);
and U1457 (N_1457,In_773,In_422);
nand U1458 (N_1458,In_503,In_1475);
nand U1459 (N_1459,In_654,In_1185);
and U1460 (N_1460,In_958,In_971);
xnor U1461 (N_1461,In_594,In_700);
and U1462 (N_1462,In_944,In_1202);
nor U1463 (N_1463,In_1335,In_164);
nand U1464 (N_1464,In_82,In_650);
or U1465 (N_1465,In_1011,In_679);
or U1466 (N_1466,In_150,In_1345);
or U1467 (N_1467,In_1405,In_966);
nand U1468 (N_1468,In_540,In_49);
or U1469 (N_1469,In_109,In_708);
nor U1470 (N_1470,In_871,In_334);
nor U1471 (N_1471,In_1044,In_382);
nand U1472 (N_1472,In_433,In_225);
nor U1473 (N_1473,In_1107,In_321);
nand U1474 (N_1474,In_630,In_1404);
nor U1475 (N_1475,In_585,In_302);
xor U1476 (N_1476,In_513,In_225);
nor U1477 (N_1477,In_1330,In_1479);
nor U1478 (N_1478,In_1279,In_792);
or U1479 (N_1479,In_1382,In_512);
nand U1480 (N_1480,In_633,In_378);
nor U1481 (N_1481,In_1037,In_158);
nand U1482 (N_1482,In_964,In_335);
and U1483 (N_1483,In_61,In_504);
nor U1484 (N_1484,In_471,In_612);
nor U1485 (N_1485,In_1401,In_1115);
and U1486 (N_1486,In_1429,In_189);
and U1487 (N_1487,In_414,In_532);
nor U1488 (N_1488,In_877,In_193);
nand U1489 (N_1489,In_1124,In_1373);
nor U1490 (N_1490,In_614,In_392);
or U1491 (N_1491,In_861,In_0);
and U1492 (N_1492,In_543,In_113);
nand U1493 (N_1493,In_62,In_1039);
nand U1494 (N_1494,In_821,In_35);
nand U1495 (N_1495,In_432,In_1441);
or U1496 (N_1496,In_925,In_773);
nand U1497 (N_1497,In_67,In_318);
nand U1498 (N_1498,In_455,In_451);
nand U1499 (N_1499,In_153,In_454);
xor U1500 (N_1500,In_1055,In_191);
or U1501 (N_1501,In_977,In_305);
xnor U1502 (N_1502,In_500,In_638);
nand U1503 (N_1503,In_936,In_1251);
xnor U1504 (N_1504,In_299,In_635);
nor U1505 (N_1505,In_47,In_53);
and U1506 (N_1506,In_114,In_645);
nor U1507 (N_1507,In_1202,In_1333);
and U1508 (N_1508,In_1093,In_390);
and U1509 (N_1509,In_215,In_568);
nand U1510 (N_1510,In_62,In_208);
or U1511 (N_1511,In_909,In_1257);
or U1512 (N_1512,In_1207,In_1230);
or U1513 (N_1513,In_757,In_985);
nor U1514 (N_1514,In_744,In_456);
nor U1515 (N_1515,In_191,In_199);
nor U1516 (N_1516,In_522,In_1203);
nand U1517 (N_1517,In_1077,In_769);
or U1518 (N_1518,In_524,In_813);
nand U1519 (N_1519,In_533,In_1189);
xor U1520 (N_1520,In_1238,In_415);
nand U1521 (N_1521,In_486,In_569);
nor U1522 (N_1522,In_1336,In_499);
xnor U1523 (N_1523,In_1263,In_743);
nand U1524 (N_1524,In_1012,In_287);
nor U1525 (N_1525,In_725,In_952);
xnor U1526 (N_1526,In_206,In_1111);
nor U1527 (N_1527,In_400,In_923);
or U1528 (N_1528,In_1235,In_452);
and U1529 (N_1529,In_491,In_373);
or U1530 (N_1530,In_1022,In_1263);
nand U1531 (N_1531,In_358,In_566);
and U1532 (N_1532,In_246,In_103);
and U1533 (N_1533,In_933,In_864);
nor U1534 (N_1534,In_1048,In_113);
or U1535 (N_1535,In_1130,In_95);
and U1536 (N_1536,In_1060,In_1050);
nor U1537 (N_1537,In_1035,In_664);
and U1538 (N_1538,In_1005,In_1358);
nand U1539 (N_1539,In_210,In_1146);
nand U1540 (N_1540,In_829,In_309);
nand U1541 (N_1541,In_816,In_325);
nand U1542 (N_1542,In_937,In_356);
or U1543 (N_1543,In_156,In_539);
xor U1544 (N_1544,In_69,In_1071);
xor U1545 (N_1545,In_1434,In_215);
nand U1546 (N_1546,In_3,In_851);
nand U1547 (N_1547,In_262,In_1212);
xor U1548 (N_1548,In_1200,In_1388);
or U1549 (N_1549,In_602,In_476);
xnor U1550 (N_1550,In_655,In_1214);
xor U1551 (N_1551,In_165,In_398);
nand U1552 (N_1552,In_344,In_1491);
nand U1553 (N_1553,In_236,In_1368);
nand U1554 (N_1554,In_106,In_1469);
or U1555 (N_1555,In_1292,In_702);
nand U1556 (N_1556,In_1343,In_1285);
nand U1557 (N_1557,In_122,In_1234);
xnor U1558 (N_1558,In_1218,In_1337);
xnor U1559 (N_1559,In_160,In_637);
nand U1560 (N_1560,In_391,In_586);
nor U1561 (N_1561,In_1367,In_1200);
and U1562 (N_1562,In_485,In_967);
nor U1563 (N_1563,In_5,In_101);
and U1564 (N_1564,In_735,In_1494);
or U1565 (N_1565,In_55,In_633);
xor U1566 (N_1566,In_1484,In_1385);
nor U1567 (N_1567,In_592,In_1419);
nor U1568 (N_1568,In_789,In_764);
nor U1569 (N_1569,In_260,In_644);
and U1570 (N_1570,In_1264,In_1202);
nor U1571 (N_1571,In_215,In_1043);
nand U1572 (N_1572,In_514,In_1323);
nor U1573 (N_1573,In_564,In_537);
nand U1574 (N_1574,In_292,In_93);
or U1575 (N_1575,In_1160,In_1173);
xnor U1576 (N_1576,In_1131,In_817);
or U1577 (N_1577,In_1132,In_1495);
nand U1578 (N_1578,In_630,In_832);
nor U1579 (N_1579,In_657,In_120);
or U1580 (N_1580,In_616,In_246);
nand U1581 (N_1581,In_1003,In_757);
and U1582 (N_1582,In_707,In_587);
nor U1583 (N_1583,In_49,In_498);
or U1584 (N_1584,In_148,In_164);
or U1585 (N_1585,In_585,In_417);
or U1586 (N_1586,In_12,In_566);
nor U1587 (N_1587,In_1497,In_635);
nand U1588 (N_1588,In_1482,In_46);
and U1589 (N_1589,In_1032,In_263);
or U1590 (N_1590,In_1129,In_520);
nor U1591 (N_1591,In_1437,In_94);
xnor U1592 (N_1592,In_452,In_1384);
nor U1593 (N_1593,In_152,In_1256);
and U1594 (N_1594,In_1229,In_659);
or U1595 (N_1595,In_681,In_905);
nand U1596 (N_1596,In_417,In_653);
xor U1597 (N_1597,In_1108,In_566);
xnor U1598 (N_1598,In_477,In_181);
or U1599 (N_1599,In_856,In_1349);
or U1600 (N_1600,In_82,In_498);
xnor U1601 (N_1601,In_892,In_602);
nor U1602 (N_1602,In_371,In_795);
and U1603 (N_1603,In_511,In_495);
nor U1604 (N_1604,In_1202,In_272);
and U1605 (N_1605,In_81,In_330);
and U1606 (N_1606,In_740,In_762);
nand U1607 (N_1607,In_991,In_824);
or U1608 (N_1608,In_362,In_356);
or U1609 (N_1609,In_956,In_475);
or U1610 (N_1610,In_100,In_425);
nor U1611 (N_1611,In_281,In_1445);
nand U1612 (N_1612,In_1064,In_85);
or U1613 (N_1613,In_140,In_1323);
or U1614 (N_1614,In_1057,In_485);
nand U1615 (N_1615,In_1085,In_702);
nand U1616 (N_1616,In_644,In_1022);
or U1617 (N_1617,In_212,In_148);
nor U1618 (N_1618,In_465,In_343);
xnor U1619 (N_1619,In_1132,In_928);
nor U1620 (N_1620,In_161,In_837);
xor U1621 (N_1621,In_801,In_960);
xor U1622 (N_1622,In_914,In_1076);
nand U1623 (N_1623,In_1147,In_868);
and U1624 (N_1624,In_1191,In_1280);
or U1625 (N_1625,In_756,In_219);
and U1626 (N_1626,In_1312,In_418);
and U1627 (N_1627,In_670,In_755);
xor U1628 (N_1628,In_1396,In_322);
nand U1629 (N_1629,In_1280,In_858);
nor U1630 (N_1630,In_788,In_650);
xnor U1631 (N_1631,In_1133,In_641);
or U1632 (N_1632,In_271,In_543);
nand U1633 (N_1633,In_408,In_115);
nand U1634 (N_1634,In_1059,In_907);
nand U1635 (N_1635,In_285,In_616);
and U1636 (N_1636,In_391,In_1008);
xor U1637 (N_1637,In_323,In_1076);
and U1638 (N_1638,In_983,In_301);
or U1639 (N_1639,In_309,In_871);
nand U1640 (N_1640,In_377,In_897);
xnor U1641 (N_1641,In_1361,In_676);
xnor U1642 (N_1642,In_1272,In_482);
xnor U1643 (N_1643,In_321,In_1286);
nand U1644 (N_1644,In_129,In_681);
xor U1645 (N_1645,In_699,In_201);
and U1646 (N_1646,In_418,In_569);
xor U1647 (N_1647,In_394,In_1185);
nand U1648 (N_1648,In_943,In_517);
xor U1649 (N_1649,In_643,In_184);
nor U1650 (N_1650,In_14,In_447);
and U1651 (N_1651,In_457,In_194);
and U1652 (N_1652,In_1213,In_307);
nand U1653 (N_1653,In_239,In_870);
or U1654 (N_1654,In_79,In_1149);
or U1655 (N_1655,In_876,In_598);
and U1656 (N_1656,In_136,In_954);
nor U1657 (N_1657,In_41,In_1087);
or U1658 (N_1658,In_1264,In_877);
nor U1659 (N_1659,In_624,In_447);
or U1660 (N_1660,In_1117,In_1468);
and U1661 (N_1661,In_819,In_938);
nand U1662 (N_1662,In_1056,In_906);
nor U1663 (N_1663,In_684,In_267);
nand U1664 (N_1664,In_118,In_92);
or U1665 (N_1665,In_1494,In_762);
nor U1666 (N_1666,In_0,In_1474);
nand U1667 (N_1667,In_1306,In_1007);
or U1668 (N_1668,In_1245,In_1341);
or U1669 (N_1669,In_228,In_255);
nand U1670 (N_1670,In_247,In_1391);
nor U1671 (N_1671,In_948,In_992);
nor U1672 (N_1672,In_318,In_437);
nor U1673 (N_1673,In_1183,In_317);
and U1674 (N_1674,In_563,In_793);
nand U1675 (N_1675,In_1066,In_482);
nand U1676 (N_1676,In_342,In_1494);
or U1677 (N_1677,In_192,In_1019);
nor U1678 (N_1678,In_1306,In_617);
or U1679 (N_1679,In_366,In_87);
nor U1680 (N_1680,In_2,In_1440);
xnor U1681 (N_1681,In_1128,In_874);
and U1682 (N_1682,In_346,In_417);
nor U1683 (N_1683,In_1043,In_33);
nor U1684 (N_1684,In_863,In_1002);
nand U1685 (N_1685,In_1112,In_263);
nor U1686 (N_1686,In_1400,In_463);
nand U1687 (N_1687,In_1467,In_653);
xnor U1688 (N_1688,In_56,In_1188);
xor U1689 (N_1689,In_1169,In_920);
nand U1690 (N_1690,In_571,In_346);
nor U1691 (N_1691,In_140,In_982);
nand U1692 (N_1692,In_915,In_758);
nand U1693 (N_1693,In_31,In_1298);
nand U1694 (N_1694,In_689,In_771);
and U1695 (N_1695,In_314,In_1458);
or U1696 (N_1696,In_655,In_842);
nor U1697 (N_1697,In_1321,In_966);
nand U1698 (N_1698,In_912,In_1119);
and U1699 (N_1699,In_926,In_1117);
nor U1700 (N_1700,In_1455,In_115);
nor U1701 (N_1701,In_327,In_497);
or U1702 (N_1702,In_1306,In_901);
nor U1703 (N_1703,In_919,In_764);
nor U1704 (N_1704,In_1464,In_575);
and U1705 (N_1705,In_47,In_1241);
or U1706 (N_1706,In_1406,In_485);
and U1707 (N_1707,In_1470,In_1121);
nor U1708 (N_1708,In_621,In_1275);
or U1709 (N_1709,In_1466,In_776);
xnor U1710 (N_1710,In_650,In_1123);
nor U1711 (N_1711,In_141,In_410);
nand U1712 (N_1712,In_1097,In_1149);
nor U1713 (N_1713,In_659,In_748);
nor U1714 (N_1714,In_1303,In_538);
nand U1715 (N_1715,In_151,In_274);
or U1716 (N_1716,In_17,In_1124);
nand U1717 (N_1717,In_75,In_635);
nand U1718 (N_1718,In_73,In_163);
xnor U1719 (N_1719,In_203,In_84);
and U1720 (N_1720,In_647,In_354);
xnor U1721 (N_1721,In_907,In_110);
or U1722 (N_1722,In_383,In_246);
nor U1723 (N_1723,In_519,In_1445);
or U1724 (N_1724,In_868,In_1322);
and U1725 (N_1725,In_1492,In_1065);
and U1726 (N_1726,In_544,In_286);
and U1727 (N_1727,In_937,In_1281);
and U1728 (N_1728,In_563,In_155);
nand U1729 (N_1729,In_97,In_620);
xnor U1730 (N_1730,In_889,In_1370);
nor U1731 (N_1731,In_141,In_563);
xnor U1732 (N_1732,In_999,In_875);
nand U1733 (N_1733,In_772,In_218);
nand U1734 (N_1734,In_210,In_1370);
and U1735 (N_1735,In_281,In_421);
or U1736 (N_1736,In_839,In_671);
nor U1737 (N_1737,In_993,In_417);
xor U1738 (N_1738,In_1482,In_69);
or U1739 (N_1739,In_1120,In_864);
nor U1740 (N_1740,In_337,In_1279);
xnor U1741 (N_1741,In_831,In_1040);
or U1742 (N_1742,In_520,In_223);
nand U1743 (N_1743,In_1234,In_667);
nor U1744 (N_1744,In_1418,In_984);
or U1745 (N_1745,In_861,In_244);
and U1746 (N_1746,In_38,In_621);
nand U1747 (N_1747,In_731,In_1056);
nand U1748 (N_1748,In_471,In_860);
xnor U1749 (N_1749,In_815,In_340);
nand U1750 (N_1750,In_251,In_274);
and U1751 (N_1751,In_114,In_445);
nand U1752 (N_1752,In_222,In_855);
or U1753 (N_1753,In_1010,In_1180);
and U1754 (N_1754,In_342,In_801);
nor U1755 (N_1755,In_533,In_354);
nor U1756 (N_1756,In_1214,In_225);
xor U1757 (N_1757,In_501,In_873);
nand U1758 (N_1758,In_538,In_979);
nand U1759 (N_1759,In_516,In_709);
nand U1760 (N_1760,In_1079,In_574);
nor U1761 (N_1761,In_652,In_683);
and U1762 (N_1762,In_807,In_344);
xor U1763 (N_1763,In_897,In_1298);
nand U1764 (N_1764,In_1268,In_918);
xnor U1765 (N_1765,In_1204,In_1483);
and U1766 (N_1766,In_555,In_62);
nor U1767 (N_1767,In_154,In_936);
nand U1768 (N_1768,In_1050,In_1315);
nor U1769 (N_1769,In_437,In_138);
xor U1770 (N_1770,In_1229,In_649);
nand U1771 (N_1771,In_721,In_252);
nor U1772 (N_1772,In_547,In_617);
nor U1773 (N_1773,In_909,In_626);
and U1774 (N_1774,In_526,In_333);
or U1775 (N_1775,In_199,In_690);
and U1776 (N_1776,In_1215,In_345);
nand U1777 (N_1777,In_1464,In_359);
and U1778 (N_1778,In_170,In_567);
and U1779 (N_1779,In_1382,In_241);
or U1780 (N_1780,In_1405,In_1326);
and U1781 (N_1781,In_1177,In_623);
xor U1782 (N_1782,In_51,In_36);
nor U1783 (N_1783,In_1493,In_1319);
and U1784 (N_1784,In_665,In_577);
and U1785 (N_1785,In_531,In_1255);
or U1786 (N_1786,In_924,In_915);
nor U1787 (N_1787,In_966,In_716);
nor U1788 (N_1788,In_340,In_1268);
nand U1789 (N_1789,In_416,In_277);
and U1790 (N_1790,In_836,In_857);
nor U1791 (N_1791,In_204,In_195);
xnor U1792 (N_1792,In_621,In_788);
nand U1793 (N_1793,In_669,In_1479);
xor U1794 (N_1794,In_694,In_842);
nor U1795 (N_1795,In_738,In_1048);
and U1796 (N_1796,In_739,In_84);
and U1797 (N_1797,In_821,In_1073);
or U1798 (N_1798,In_1365,In_719);
xor U1799 (N_1799,In_1411,In_1405);
nor U1800 (N_1800,In_114,In_1050);
nand U1801 (N_1801,In_114,In_907);
xor U1802 (N_1802,In_1495,In_1454);
nand U1803 (N_1803,In_462,In_1327);
xnor U1804 (N_1804,In_641,In_1276);
and U1805 (N_1805,In_895,In_288);
and U1806 (N_1806,In_1056,In_264);
nand U1807 (N_1807,In_1130,In_819);
and U1808 (N_1808,In_497,In_683);
or U1809 (N_1809,In_491,In_251);
or U1810 (N_1810,In_64,In_917);
or U1811 (N_1811,In_1324,In_730);
and U1812 (N_1812,In_663,In_601);
or U1813 (N_1813,In_563,In_154);
nand U1814 (N_1814,In_1141,In_484);
or U1815 (N_1815,In_184,In_1419);
or U1816 (N_1816,In_565,In_1114);
nor U1817 (N_1817,In_1135,In_925);
nor U1818 (N_1818,In_1461,In_80);
nor U1819 (N_1819,In_379,In_1079);
xor U1820 (N_1820,In_819,In_711);
nand U1821 (N_1821,In_752,In_747);
xor U1822 (N_1822,In_731,In_426);
xor U1823 (N_1823,In_1024,In_273);
nor U1824 (N_1824,In_1110,In_1018);
xnor U1825 (N_1825,In_712,In_727);
or U1826 (N_1826,In_1315,In_84);
or U1827 (N_1827,In_763,In_743);
nor U1828 (N_1828,In_31,In_789);
and U1829 (N_1829,In_1438,In_1036);
nor U1830 (N_1830,In_426,In_264);
xnor U1831 (N_1831,In_29,In_696);
nor U1832 (N_1832,In_805,In_972);
xnor U1833 (N_1833,In_882,In_143);
and U1834 (N_1834,In_803,In_55);
xor U1835 (N_1835,In_763,In_1084);
or U1836 (N_1836,In_297,In_1104);
xnor U1837 (N_1837,In_1361,In_619);
nor U1838 (N_1838,In_1196,In_25);
nor U1839 (N_1839,In_500,In_934);
xnor U1840 (N_1840,In_1434,In_1046);
nor U1841 (N_1841,In_838,In_1051);
nand U1842 (N_1842,In_385,In_777);
nand U1843 (N_1843,In_30,In_184);
nor U1844 (N_1844,In_1018,In_889);
nand U1845 (N_1845,In_1036,In_903);
and U1846 (N_1846,In_169,In_383);
nor U1847 (N_1847,In_1170,In_1216);
or U1848 (N_1848,In_577,In_1070);
or U1849 (N_1849,In_1297,In_375);
nor U1850 (N_1850,In_1479,In_561);
nand U1851 (N_1851,In_907,In_967);
xor U1852 (N_1852,In_276,In_459);
nor U1853 (N_1853,In_722,In_486);
nand U1854 (N_1854,In_1009,In_1202);
or U1855 (N_1855,In_1468,In_1452);
or U1856 (N_1856,In_472,In_1109);
or U1857 (N_1857,In_882,In_137);
and U1858 (N_1858,In_1388,In_292);
nor U1859 (N_1859,In_997,In_1345);
or U1860 (N_1860,In_76,In_234);
and U1861 (N_1861,In_694,In_174);
and U1862 (N_1862,In_651,In_1306);
or U1863 (N_1863,In_270,In_488);
or U1864 (N_1864,In_71,In_864);
xor U1865 (N_1865,In_662,In_895);
and U1866 (N_1866,In_32,In_1131);
xnor U1867 (N_1867,In_954,In_369);
xor U1868 (N_1868,In_1008,In_1327);
and U1869 (N_1869,In_735,In_302);
and U1870 (N_1870,In_1179,In_1130);
xnor U1871 (N_1871,In_491,In_524);
or U1872 (N_1872,In_1277,In_505);
nand U1873 (N_1873,In_689,In_549);
and U1874 (N_1874,In_1406,In_2);
xnor U1875 (N_1875,In_550,In_348);
and U1876 (N_1876,In_1298,In_517);
xnor U1877 (N_1877,In_1486,In_1323);
and U1878 (N_1878,In_604,In_1187);
nor U1879 (N_1879,In_820,In_636);
nand U1880 (N_1880,In_1215,In_1156);
xnor U1881 (N_1881,In_421,In_603);
and U1882 (N_1882,In_629,In_1313);
nand U1883 (N_1883,In_610,In_777);
or U1884 (N_1884,In_555,In_627);
xnor U1885 (N_1885,In_495,In_356);
nand U1886 (N_1886,In_943,In_662);
and U1887 (N_1887,In_904,In_497);
and U1888 (N_1888,In_726,In_98);
nand U1889 (N_1889,In_687,In_1048);
nand U1890 (N_1890,In_1295,In_1296);
nor U1891 (N_1891,In_430,In_468);
nand U1892 (N_1892,In_95,In_1267);
and U1893 (N_1893,In_676,In_206);
xnor U1894 (N_1894,In_813,In_915);
nand U1895 (N_1895,In_183,In_617);
and U1896 (N_1896,In_529,In_1210);
xor U1897 (N_1897,In_417,In_643);
nand U1898 (N_1898,In_580,In_111);
xnor U1899 (N_1899,In_491,In_121);
and U1900 (N_1900,In_1276,In_587);
nor U1901 (N_1901,In_208,In_914);
and U1902 (N_1902,In_850,In_732);
or U1903 (N_1903,In_488,In_636);
and U1904 (N_1904,In_808,In_866);
and U1905 (N_1905,In_860,In_330);
and U1906 (N_1906,In_554,In_718);
nand U1907 (N_1907,In_1222,In_970);
xor U1908 (N_1908,In_300,In_413);
and U1909 (N_1909,In_1371,In_515);
nor U1910 (N_1910,In_564,In_81);
nand U1911 (N_1911,In_850,In_1048);
nor U1912 (N_1912,In_1421,In_797);
xnor U1913 (N_1913,In_868,In_997);
nor U1914 (N_1914,In_764,In_883);
nand U1915 (N_1915,In_173,In_605);
nand U1916 (N_1916,In_1140,In_371);
xor U1917 (N_1917,In_901,In_802);
and U1918 (N_1918,In_1317,In_1283);
and U1919 (N_1919,In_739,In_1338);
nor U1920 (N_1920,In_368,In_1263);
and U1921 (N_1921,In_724,In_190);
xor U1922 (N_1922,In_1204,In_1115);
nor U1923 (N_1923,In_615,In_916);
and U1924 (N_1924,In_1231,In_721);
nor U1925 (N_1925,In_824,In_1095);
nor U1926 (N_1926,In_371,In_891);
xnor U1927 (N_1927,In_780,In_48);
nor U1928 (N_1928,In_549,In_477);
or U1929 (N_1929,In_863,In_140);
xnor U1930 (N_1930,In_1332,In_34);
nor U1931 (N_1931,In_825,In_845);
and U1932 (N_1932,In_868,In_559);
or U1933 (N_1933,In_869,In_143);
nand U1934 (N_1934,In_482,In_1281);
and U1935 (N_1935,In_41,In_1016);
nor U1936 (N_1936,In_980,In_401);
nand U1937 (N_1937,In_1245,In_9);
and U1938 (N_1938,In_5,In_482);
nand U1939 (N_1939,In_930,In_928);
nor U1940 (N_1940,In_889,In_1034);
or U1941 (N_1941,In_659,In_1002);
or U1942 (N_1942,In_155,In_1192);
and U1943 (N_1943,In_1056,In_1237);
nand U1944 (N_1944,In_674,In_946);
or U1945 (N_1945,In_1389,In_814);
and U1946 (N_1946,In_509,In_465);
and U1947 (N_1947,In_1115,In_62);
nand U1948 (N_1948,In_831,In_978);
and U1949 (N_1949,In_1237,In_751);
xnor U1950 (N_1950,In_185,In_945);
and U1951 (N_1951,In_1257,In_1189);
nand U1952 (N_1952,In_52,In_802);
and U1953 (N_1953,In_839,In_934);
nor U1954 (N_1954,In_440,In_353);
or U1955 (N_1955,In_842,In_70);
or U1956 (N_1956,In_534,In_1082);
and U1957 (N_1957,In_153,In_434);
xnor U1958 (N_1958,In_82,In_1046);
nor U1959 (N_1959,In_1355,In_1318);
nand U1960 (N_1960,In_279,In_535);
nand U1961 (N_1961,In_1238,In_1056);
nor U1962 (N_1962,In_458,In_148);
xor U1963 (N_1963,In_1114,In_193);
nand U1964 (N_1964,In_1445,In_1025);
or U1965 (N_1965,In_190,In_129);
nand U1966 (N_1966,In_1112,In_390);
or U1967 (N_1967,In_629,In_1371);
and U1968 (N_1968,In_490,In_272);
xor U1969 (N_1969,In_1176,In_342);
nand U1970 (N_1970,In_129,In_899);
or U1971 (N_1971,In_664,In_1429);
xor U1972 (N_1972,In_315,In_1268);
and U1973 (N_1973,In_723,In_1453);
nand U1974 (N_1974,In_828,In_717);
nor U1975 (N_1975,In_1296,In_1395);
nand U1976 (N_1976,In_612,In_1108);
nand U1977 (N_1977,In_784,In_952);
nor U1978 (N_1978,In_895,In_647);
and U1979 (N_1979,In_983,In_1439);
or U1980 (N_1980,In_359,In_177);
or U1981 (N_1981,In_323,In_371);
nand U1982 (N_1982,In_1281,In_330);
and U1983 (N_1983,In_452,In_1033);
and U1984 (N_1984,In_13,In_1203);
nand U1985 (N_1985,In_425,In_293);
nor U1986 (N_1986,In_1171,In_349);
and U1987 (N_1987,In_656,In_497);
nand U1988 (N_1988,In_1408,In_845);
or U1989 (N_1989,In_918,In_269);
or U1990 (N_1990,In_724,In_1386);
nor U1991 (N_1991,In_1095,In_1431);
xor U1992 (N_1992,In_1284,In_453);
xnor U1993 (N_1993,In_781,In_1119);
nand U1994 (N_1994,In_889,In_1178);
and U1995 (N_1995,In_1426,In_88);
nor U1996 (N_1996,In_932,In_102);
xor U1997 (N_1997,In_459,In_993);
nand U1998 (N_1998,In_1426,In_355);
nand U1999 (N_1999,In_670,In_762);
and U2000 (N_2000,In_511,In_997);
and U2001 (N_2001,In_212,In_56);
or U2002 (N_2002,In_773,In_243);
and U2003 (N_2003,In_671,In_715);
and U2004 (N_2004,In_1088,In_973);
xnor U2005 (N_2005,In_1164,In_156);
nand U2006 (N_2006,In_1174,In_22);
and U2007 (N_2007,In_1203,In_760);
nor U2008 (N_2008,In_279,In_1166);
nand U2009 (N_2009,In_1410,In_475);
or U2010 (N_2010,In_1061,In_1089);
or U2011 (N_2011,In_312,In_670);
nor U2012 (N_2012,In_660,In_1032);
nand U2013 (N_2013,In_137,In_79);
xor U2014 (N_2014,In_1232,In_270);
or U2015 (N_2015,In_1074,In_311);
nor U2016 (N_2016,In_126,In_617);
nand U2017 (N_2017,In_1152,In_300);
and U2018 (N_2018,In_73,In_421);
xor U2019 (N_2019,In_1401,In_64);
nor U2020 (N_2020,In_808,In_586);
nor U2021 (N_2021,In_304,In_1453);
nand U2022 (N_2022,In_755,In_824);
nor U2023 (N_2023,In_1470,In_1138);
or U2024 (N_2024,In_69,In_1311);
and U2025 (N_2025,In_113,In_1017);
nor U2026 (N_2026,In_109,In_517);
and U2027 (N_2027,In_969,In_46);
xor U2028 (N_2028,In_131,In_477);
or U2029 (N_2029,In_1142,In_558);
or U2030 (N_2030,In_1061,In_1049);
nor U2031 (N_2031,In_165,In_855);
and U2032 (N_2032,In_1416,In_1280);
nand U2033 (N_2033,In_1431,In_508);
nand U2034 (N_2034,In_25,In_332);
nor U2035 (N_2035,In_99,In_579);
and U2036 (N_2036,In_416,In_1139);
or U2037 (N_2037,In_419,In_1226);
xor U2038 (N_2038,In_31,In_596);
or U2039 (N_2039,In_528,In_578);
nand U2040 (N_2040,In_1249,In_72);
nand U2041 (N_2041,In_829,In_410);
nand U2042 (N_2042,In_1069,In_657);
xor U2043 (N_2043,In_1496,In_1060);
or U2044 (N_2044,In_597,In_317);
or U2045 (N_2045,In_492,In_556);
nand U2046 (N_2046,In_1185,In_511);
nand U2047 (N_2047,In_1083,In_1192);
nand U2048 (N_2048,In_1448,In_329);
xnor U2049 (N_2049,In_747,In_299);
nor U2050 (N_2050,In_265,In_743);
nor U2051 (N_2051,In_930,In_273);
nor U2052 (N_2052,In_16,In_1419);
and U2053 (N_2053,In_1109,In_1202);
nor U2054 (N_2054,In_912,In_1202);
nand U2055 (N_2055,In_318,In_945);
nor U2056 (N_2056,In_1255,In_1185);
xnor U2057 (N_2057,In_1068,In_622);
nand U2058 (N_2058,In_952,In_1193);
and U2059 (N_2059,In_1148,In_171);
xor U2060 (N_2060,In_308,In_844);
and U2061 (N_2061,In_1468,In_1342);
and U2062 (N_2062,In_1371,In_300);
nor U2063 (N_2063,In_584,In_698);
or U2064 (N_2064,In_436,In_1312);
nor U2065 (N_2065,In_1325,In_445);
or U2066 (N_2066,In_923,In_179);
nand U2067 (N_2067,In_39,In_877);
xor U2068 (N_2068,In_1258,In_655);
or U2069 (N_2069,In_249,In_854);
or U2070 (N_2070,In_1179,In_260);
nor U2071 (N_2071,In_1480,In_363);
nor U2072 (N_2072,In_1207,In_1238);
and U2073 (N_2073,In_924,In_243);
xnor U2074 (N_2074,In_854,In_1122);
or U2075 (N_2075,In_909,In_1126);
nand U2076 (N_2076,In_775,In_182);
nand U2077 (N_2077,In_40,In_1117);
or U2078 (N_2078,In_678,In_133);
xnor U2079 (N_2079,In_1252,In_243);
nor U2080 (N_2080,In_783,In_1229);
nand U2081 (N_2081,In_1029,In_345);
nand U2082 (N_2082,In_1400,In_885);
xor U2083 (N_2083,In_232,In_376);
and U2084 (N_2084,In_778,In_1178);
xnor U2085 (N_2085,In_1431,In_647);
nand U2086 (N_2086,In_610,In_873);
nor U2087 (N_2087,In_1299,In_1283);
nand U2088 (N_2088,In_1393,In_305);
nor U2089 (N_2089,In_163,In_1454);
and U2090 (N_2090,In_94,In_545);
and U2091 (N_2091,In_1498,In_1146);
nand U2092 (N_2092,In_1121,In_644);
or U2093 (N_2093,In_214,In_413);
nand U2094 (N_2094,In_172,In_92);
and U2095 (N_2095,In_1212,In_874);
and U2096 (N_2096,In_544,In_800);
nor U2097 (N_2097,In_141,In_1193);
and U2098 (N_2098,In_110,In_1340);
nor U2099 (N_2099,In_245,In_753);
nand U2100 (N_2100,In_388,In_70);
nor U2101 (N_2101,In_766,In_388);
xnor U2102 (N_2102,In_737,In_1066);
nor U2103 (N_2103,In_62,In_436);
nand U2104 (N_2104,In_23,In_891);
xnor U2105 (N_2105,In_308,In_413);
or U2106 (N_2106,In_848,In_1142);
and U2107 (N_2107,In_256,In_503);
or U2108 (N_2108,In_342,In_288);
or U2109 (N_2109,In_763,In_1421);
or U2110 (N_2110,In_594,In_402);
xnor U2111 (N_2111,In_13,In_1070);
nand U2112 (N_2112,In_960,In_506);
xor U2113 (N_2113,In_99,In_721);
or U2114 (N_2114,In_541,In_269);
and U2115 (N_2115,In_1431,In_436);
and U2116 (N_2116,In_813,In_1426);
and U2117 (N_2117,In_159,In_1322);
xor U2118 (N_2118,In_907,In_16);
xnor U2119 (N_2119,In_72,In_1369);
nand U2120 (N_2120,In_696,In_275);
or U2121 (N_2121,In_837,In_1393);
nand U2122 (N_2122,In_1277,In_659);
nor U2123 (N_2123,In_1083,In_583);
and U2124 (N_2124,In_831,In_386);
nand U2125 (N_2125,In_1299,In_532);
nand U2126 (N_2126,In_495,In_1412);
xor U2127 (N_2127,In_242,In_59);
and U2128 (N_2128,In_1483,In_1223);
xnor U2129 (N_2129,In_1192,In_1392);
nand U2130 (N_2130,In_1134,In_129);
nand U2131 (N_2131,In_1083,In_403);
and U2132 (N_2132,In_565,In_230);
xor U2133 (N_2133,In_490,In_751);
nor U2134 (N_2134,In_51,In_654);
xor U2135 (N_2135,In_56,In_1077);
and U2136 (N_2136,In_766,In_1074);
or U2137 (N_2137,In_358,In_58);
or U2138 (N_2138,In_386,In_1008);
xor U2139 (N_2139,In_172,In_860);
nand U2140 (N_2140,In_1090,In_258);
or U2141 (N_2141,In_518,In_101);
nor U2142 (N_2142,In_1392,In_966);
and U2143 (N_2143,In_281,In_914);
nor U2144 (N_2144,In_821,In_804);
or U2145 (N_2145,In_1087,In_670);
xor U2146 (N_2146,In_146,In_959);
nand U2147 (N_2147,In_859,In_700);
xnor U2148 (N_2148,In_977,In_82);
or U2149 (N_2149,In_456,In_392);
and U2150 (N_2150,In_498,In_688);
and U2151 (N_2151,In_1318,In_574);
or U2152 (N_2152,In_259,In_357);
or U2153 (N_2153,In_1154,In_803);
and U2154 (N_2154,In_861,In_336);
xor U2155 (N_2155,In_529,In_1055);
and U2156 (N_2156,In_56,In_404);
or U2157 (N_2157,In_448,In_880);
nand U2158 (N_2158,In_324,In_810);
nand U2159 (N_2159,In_1373,In_752);
and U2160 (N_2160,In_1373,In_908);
and U2161 (N_2161,In_178,In_517);
xnor U2162 (N_2162,In_503,In_1267);
nor U2163 (N_2163,In_321,In_338);
and U2164 (N_2164,In_132,In_1342);
or U2165 (N_2165,In_724,In_1030);
xor U2166 (N_2166,In_336,In_315);
and U2167 (N_2167,In_1018,In_289);
and U2168 (N_2168,In_1218,In_603);
nand U2169 (N_2169,In_1228,In_1317);
or U2170 (N_2170,In_374,In_778);
nand U2171 (N_2171,In_1080,In_945);
xnor U2172 (N_2172,In_197,In_433);
nand U2173 (N_2173,In_1059,In_832);
or U2174 (N_2174,In_438,In_1063);
and U2175 (N_2175,In_271,In_1036);
nand U2176 (N_2176,In_106,In_1203);
and U2177 (N_2177,In_1198,In_1246);
or U2178 (N_2178,In_983,In_1058);
and U2179 (N_2179,In_648,In_618);
nor U2180 (N_2180,In_778,In_730);
and U2181 (N_2181,In_1437,In_809);
nand U2182 (N_2182,In_969,In_1263);
xnor U2183 (N_2183,In_1229,In_1284);
xor U2184 (N_2184,In_249,In_1014);
nand U2185 (N_2185,In_171,In_582);
xor U2186 (N_2186,In_437,In_1408);
nor U2187 (N_2187,In_1195,In_451);
and U2188 (N_2188,In_1189,In_1152);
xnor U2189 (N_2189,In_187,In_287);
nand U2190 (N_2190,In_997,In_1038);
nand U2191 (N_2191,In_216,In_321);
nand U2192 (N_2192,In_1158,In_935);
xor U2193 (N_2193,In_629,In_561);
nand U2194 (N_2194,In_485,In_1329);
or U2195 (N_2195,In_726,In_283);
nand U2196 (N_2196,In_1395,In_1108);
and U2197 (N_2197,In_1015,In_255);
xor U2198 (N_2198,In_730,In_414);
xnor U2199 (N_2199,In_241,In_1053);
xnor U2200 (N_2200,In_1167,In_1324);
nor U2201 (N_2201,In_798,In_671);
and U2202 (N_2202,In_414,In_28);
nor U2203 (N_2203,In_717,In_1174);
nor U2204 (N_2204,In_126,In_1167);
xor U2205 (N_2205,In_349,In_454);
and U2206 (N_2206,In_973,In_150);
nor U2207 (N_2207,In_616,In_120);
and U2208 (N_2208,In_1201,In_706);
nor U2209 (N_2209,In_1018,In_959);
nor U2210 (N_2210,In_339,In_1242);
or U2211 (N_2211,In_1244,In_674);
nor U2212 (N_2212,In_1206,In_1027);
xor U2213 (N_2213,In_896,In_988);
nor U2214 (N_2214,In_417,In_1108);
nor U2215 (N_2215,In_319,In_741);
nor U2216 (N_2216,In_900,In_823);
nor U2217 (N_2217,In_1046,In_1386);
nor U2218 (N_2218,In_623,In_1172);
or U2219 (N_2219,In_746,In_980);
nand U2220 (N_2220,In_485,In_540);
or U2221 (N_2221,In_812,In_791);
nand U2222 (N_2222,In_1117,In_533);
nand U2223 (N_2223,In_1389,In_1471);
and U2224 (N_2224,In_673,In_1167);
nor U2225 (N_2225,In_715,In_171);
nand U2226 (N_2226,In_650,In_1284);
xnor U2227 (N_2227,In_1437,In_1483);
or U2228 (N_2228,In_119,In_133);
nor U2229 (N_2229,In_943,In_801);
and U2230 (N_2230,In_794,In_59);
nor U2231 (N_2231,In_367,In_574);
xor U2232 (N_2232,In_892,In_940);
nor U2233 (N_2233,In_574,In_237);
and U2234 (N_2234,In_1287,In_577);
or U2235 (N_2235,In_764,In_1069);
xor U2236 (N_2236,In_765,In_574);
or U2237 (N_2237,In_727,In_1159);
or U2238 (N_2238,In_100,In_222);
nor U2239 (N_2239,In_1210,In_889);
xnor U2240 (N_2240,In_1309,In_786);
xor U2241 (N_2241,In_1454,In_307);
nor U2242 (N_2242,In_271,In_1462);
and U2243 (N_2243,In_200,In_1337);
and U2244 (N_2244,In_126,In_1053);
and U2245 (N_2245,In_576,In_1125);
xnor U2246 (N_2246,In_506,In_119);
nor U2247 (N_2247,In_1339,In_776);
and U2248 (N_2248,In_1010,In_1317);
nand U2249 (N_2249,In_935,In_704);
or U2250 (N_2250,In_837,In_1167);
nand U2251 (N_2251,In_999,In_572);
and U2252 (N_2252,In_51,In_791);
and U2253 (N_2253,In_1299,In_1497);
and U2254 (N_2254,In_172,In_656);
nor U2255 (N_2255,In_37,In_827);
nor U2256 (N_2256,In_592,In_890);
nand U2257 (N_2257,In_548,In_433);
or U2258 (N_2258,In_548,In_1204);
xnor U2259 (N_2259,In_98,In_904);
and U2260 (N_2260,In_1351,In_1281);
and U2261 (N_2261,In_1034,In_489);
nand U2262 (N_2262,In_723,In_784);
and U2263 (N_2263,In_1286,In_796);
xnor U2264 (N_2264,In_679,In_297);
nor U2265 (N_2265,In_927,In_1328);
xor U2266 (N_2266,In_188,In_934);
and U2267 (N_2267,In_1113,In_679);
nor U2268 (N_2268,In_763,In_1048);
xnor U2269 (N_2269,In_1441,In_743);
nor U2270 (N_2270,In_602,In_1286);
and U2271 (N_2271,In_440,In_1024);
xor U2272 (N_2272,In_1392,In_578);
and U2273 (N_2273,In_1360,In_681);
xnor U2274 (N_2274,In_1191,In_1225);
nand U2275 (N_2275,In_831,In_1248);
and U2276 (N_2276,In_1045,In_96);
nor U2277 (N_2277,In_1161,In_110);
nor U2278 (N_2278,In_1392,In_219);
and U2279 (N_2279,In_529,In_751);
xor U2280 (N_2280,In_1385,In_252);
xor U2281 (N_2281,In_422,In_687);
or U2282 (N_2282,In_659,In_802);
and U2283 (N_2283,In_517,In_500);
or U2284 (N_2284,In_400,In_807);
nor U2285 (N_2285,In_115,In_1175);
nor U2286 (N_2286,In_397,In_1280);
and U2287 (N_2287,In_382,In_722);
and U2288 (N_2288,In_771,In_487);
xor U2289 (N_2289,In_1443,In_54);
xor U2290 (N_2290,In_242,In_1276);
nand U2291 (N_2291,In_779,In_344);
xor U2292 (N_2292,In_968,In_1380);
xor U2293 (N_2293,In_925,In_859);
nor U2294 (N_2294,In_1457,In_139);
and U2295 (N_2295,In_910,In_807);
nor U2296 (N_2296,In_811,In_261);
and U2297 (N_2297,In_404,In_59);
nor U2298 (N_2298,In_720,In_216);
and U2299 (N_2299,In_886,In_1002);
or U2300 (N_2300,In_1176,In_1478);
and U2301 (N_2301,In_1320,In_52);
and U2302 (N_2302,In_165,In_15);
or U2303 (N_2303,In_1399,In_1227);
nand U2304 (N_2304,In_305,In_1096);
nor U2305 (N_2305,In_764,In_529);
and U2306 (N_2306,In_361,In_701);
nand U2307 (N_2307,In_721,In_699);
and U2308 (N_2308,In_348,In_1206);
nor U2309 (N_2309,In_805,In_645);
and U2310 (N_2310,In_827,In_176);
nand U2311 (N_2311,In_319,In_1139);
nand U2312 (N_2312,In_1330,In_1220);
nor U2313 (N_2313,In_1249,In_1384);
nand U2314 (N_2314,In_270,In_1257);
xor U2315 (N_2315,In_1262,In_481);
or U2316 (N_2316,In_1069,In_1437);
xnor U2317 (N_2317,In_53,In_339);
xnor U2318 (N_2318,In_148,In_1245);
and U2319 (N_2319,In_9,In_1158);
nor U2320 (N_2320,In_278,In_1208);
and U2321 (N_2321,In_268,In_1397);
and U2322 (N_2322,In_121,In_316);
xnor U2323 (N_2323,In_628,In_1003);
nor U2324 (N_2324,In_1357,In_824);
or U2325 (N_2325,In_1117,In_607);
xor U2326 (N_2326,In_26,In_645);
nand U2327 (N_2327,In_855,In_723);
and U2328 (N_2328,In_10,In_381);
and U2329 (N_2329,In_537,In_1341);
nor U2330 (N_2330,In_805,In_498);
xor U2331 (N_2331,In_486,In_775);
and U2332 (N_2332,In_1318,In_1071);
xor U2333 (N_2333,In_626,In_921);
or U2334 (N_2334,In_1036,In_708);
or U2335 (N_2335,In_1473,In_390);
xnor U2336 (N_2336,In_603,In_1449);
or U2337 (N_2337,In_1289,In_353);
nand U2338 (N_2338,In_707,In_28);
xor U2339 (N_2339,In_1011,In_24);
or U2340 (N_2340,In_738,In_882);
nand U2341 (N_2341,In_130,In_427);
xor U2342 (N_2342,In_67,In_1125);
nor U2343 (N_2343,In_993,In_533);
xnor U2344 (N_2344,In_500,In_1157);
xnor U2345 (N_2345,In_1286,In_1018);
or U2346 (N_2346,In_803,In_667);
or U2347 (N_2347,In_1318,In_370);
xor U2348 (N_2348,In_460,In_1447);
xnor U2349 (N_2349,In_537,In_447);
nor U2350 (N_2350,In_778,In_1164);
xor U2351 (N_2351,In_698,In_1452);
and U2352 (N_2352,In_909,In_644);
and U2353 (N_2353,In_1466,In_1341);
nand U2354 (N_2354,In_593,In_1341);
nor U2355 (N_2355,In_956,In_291);
or U2356 (N_2356,In_301,In_135);
nor U2357 (N_2357,In_979,In_353);
and U2358 (N_2358,In_212,In_591);
xnor U2359 (N_2359,In_1196,In_282);
nor U2360 (N_2360,In_1108,In_830);
nand U2361 (N_2361,In_742,In_1471);
xor U2362 (N_2362,In_554,In_1216);
or U2363 (N_2363,In_264,In_313);
nand U2364 (N_2364,In_1069,In_28);
or U2365 (N_2365,In_1397,In_669);
xnor U2366 (N_2366,In_1132,In_1323);
nor U2367 (N_2367,In_427,In_354);
xnor U2368 (N_2368,In_156,In_1464);
and U2369 (N_2369,In_274,In_1456);
xnor U2370 (N_2370,In_842,In_382);
xnor U2371 (N_2371,In_869,In_1017);
nand U2372 (N_2372,In_773,In_29);
nor U2373 (N_2373,In_1159,In_301);
nor U2374 (N_2374,In_846,In_949);
nand U2375 (N_2375,In_1107,In_160);
nand U2376 (N_2376,In_616,In_1487);
xnor U2377 (N_2377,In_7,In_1002);
nor U2378 (N_2378,In_190,In_1342);
or U2379 (N_2379,In_1259,In_307);
xnor U2380 (N_2380,In_1302,In_1111);
nor U2381 (N_2381,In_1499,In_390);
and U2382 (N_2382,In_452,In_1422);
and U2383 (N_2383,In_1230,In_321);
or U2384 (N_2384,In_952,In_370);
and U2385 (N_2385,In_368,In_1257);
or U2386 (N_2386,In_983,In_958);
or U2387 (N_2387,In_583,In_1322);
and U2388 (N_2388,In_22,In_625);
nor U2389 (N_2389,In_138,In_1230);
nand U2390 (N_2390,In_296,In_603);
and U2391 (N_2391,In_798,In_1357);
nor U2392 (N_2392,In_208,In_1266);
xor U2393 (N_2393,In_1246,In_266);
nand U2394 (N_2394,In_1164,In_1297);
nand U2395 (N_2395,In_831,In_383);
or U2396 (N_2396,In_611,In_705);
and U2397 (N_2397,In_1243,In_1301);
nand U2398 (N_2398,In_644,In_318);
nand U2399 (N_2399,In_1025,In_145);
or U2400 (N_2400,In_157,In_548);
nand U2401 (N_2401,In_998,In_245);
xnor U2402 (N_2402,In_225,In_1191);
nand U2403 (N_2403,In_71,In_947);
xnor U2404 (N_2404,In_223,In_10);
and U2405 (N_2405,In_285,In_472);
nand U2406 (N_2406,In_1387,In_64);
xnor U2407 (N_2407,In_1463,In_24);
or U2408 (N_2408,In_1153,In_608);
and U2409 (N_2409,In_72,In_536);
or U2410 (N_2410,In_841,In_347);
and U2411 (N_2411,In_843,In_139);
nand U2412 (N_2412,In_1282,In_44);
and U2413 (N_2413,In_985,In_1164);
and U2414 (N_2414,In_135,In_323);
or U2415 (N_2415,In_230,In_395);
nor U2416 (N_2416,In_633,In_525);
or U2417 (N_2417,In_327,In_270);
nand U2418 (N_2418,In_1125,In_714);
xor U2419 (N_2419,In_861,In_109);
or U2420 (N_2420,In_1225,In_1278);
or U2421 (N_2421,In_1010,In_313);
xor U2422 (N_2422,In_299,In_420);
and U2423 (N_2423,In_647,In_748);
nand U2424 (N_2424,In_944,In_1270);
and U2425 (N_2425,In_738,In_339);
xnor U2426 (N_2426,In_275,In_865);
nor U2427 (N_2427,In_694,In_349);
nand U2428 (N_2428,In_675,In_700);
and U2429 (N_2429,In_1358,In_465);
xnor U2430 (N_2430,In_901,In_1242);
nor U2431 (N_2431,In_1297,In_660);
nand U2432 (N_2432,In_1322,In_150);
xor U2433 (N_2433,In_1366,In_1098);
nand U2434 (N_2434,In_1112,In_573);
nor U2435 (N_2435,In_705,In_1131);
or U2436 (N_2436,In_978,In_1427);
nand U2437 (N_2437,In_737,In_968);
and U2438 (N_2438,In_1428,In_280);
nand U2439 (N_2439,In_824,In_500);
nor U2440 (N_2440,In_435,In_1009);
nand U2441 (N_2441,In_791,In_41);
or U2442 (N_2442,In_903,In_1403);
or U2443 (N_2443,In_1104,In_461);
nand U2444 (N_2444,In_351,In_62);
and U2445 (N_2445,In_945,In_491);
or U2446 (N_2446,In_962,In_1384);
nor U2447 (N_2447,In_932,In_289);
nor U2448 (N_2448,In_82,In_692);
and U2449 (N_2449,In_1103,In_210);
and U2450 (N_2450,In_423,In_1239);
nor U2451 (N_2451,In_265,In_880);
xnor U2452 (N_2452,In_190,In_4);
nor U2453 (N_2453,In_1155,In_835);
xnor U2454 (N_2454,In_17,In_1451);
nor U2455 (N_2455,In_1287,In_1305);
xnor U2456 (N_2456,In_1443,In_1277);
or U2457 (N_2457,In_502,In_279);
nand U2458 (N_2458,In_279,In_498);
and U2459 (N_2459,In_1026,In_1440);
nor U2460 (N_2460,In_638,In_888);
xor U2461 (N_2461,In_1247,In_1390);
xor U2462 (N_2462,In_225,In_228);
and U2463 (N_2463,In_325,In_861);
xnor U2464 (N_2464,In_72,In_1036);
and U2465 (N_2465,In_907,In_386);
or U2466 (N_2466,In_890,In_3);
nand U2467 (N_2467,In_865,In_1340);
xor U2468 (N_2468,In_1239,In_8);
nor U2469 (N_2469,In_524,In_357);
nand U2470 (N_2470,In_1408,In_386);
or U2471 (N_2471,In_894,In_1498);
xnor U2472 (N_2472,In_1340,In_1215);
nand U2473 (N_2473,In_502,In_1334);
and U2474 (N_2474,In_977,In_980);
and U2475 (N_2475,In_118,In_451);
nand U2476 (N_2476,In_1294,In_192);
and U2477 (N_2477,In_1468,In_163);
xor U2478 (N_2478,In_53,In_1413);
and U2479 (N_2479,In_813,In_1207);
nand U2480 (N_2480,In_105,In_68);
nand U2481 (N_2481,In_410,In_1022);
xor U2482 (N_2482,In_429,In_629);
or U2483 (N_2483,In_621,In_382);
nor U2484 (N_2484,In_174,In_914);
or U2485 (N_2485,In_1196,In_1005);
nand U2486 (N_2486,In_817,In_1378);
and U2487 (N_2487,In_670,In_697);
or U2488 (N_2488,In_1486,In_1417);
or U2489 (N_2489,In_691,In_703);
or U2490 (N_2490,In_72,In_288);
nor U2491 (N_2491,In_160,In_758);
or U2492 (N_2492,In_1070,In_1114);
and U2493 (N_2493,In_48,In_1171);
and U2494 (N_2494,In_1453,In_355);
and U2495 (N_2495,In_1446,In_1105);
xor U2496 (N_2496,In_1374,In_1197);
nor U2497 (N_2497,In_221,In_1442);
nor U2498 (N_2498,In_940,In_1420);
nor U2499 (N_2499,In_861,In_1204);
nor U2500 (N_2500,In_984,In_375);
xnor U2501 (N_2501,In_1329,In_1334);
nor U2502 (N_2502,In_1019,In_18);
nand U2503 (N_2503,In_1214,In_1454);
nand U2504 (N_2504,In_151,In_802);
nor U2505 (N_2505,In_531,In_447);
xnor U2506 (N_2506,In_103,In_833);
nand U2507 (N_2507,In_310,In_69);
nand U2508 (N_2508,In_21,In_1000);
nand U2509 (N_2509,In_1414,In_471);
or U2510 (N_2510,In_50,In_1325);
and U2511 (N_2511,In_915,In_1041);
xor U2512 (N_2512,In_628,In_1444);
nand U2513 (N_2513,In_109,In_203);
nor U2514 (N_2514,In_1015,In_1162);
nand U2515 (N_2515,In_859,In_1465);
nand U2516 (N_2516,In_67,In_431);
nand U2517 (N_2517,In_262,In_693);
xor U2518 (N_2518,In_1179,In_1292);
and U2519 (N_2519,In_994,In_897);
xnor U2520 (N_2520,In_1223,In_1163);
nor U2521 (N_2521,In_473,In_18);
and U2522 (N_2522,In_902,In_1157);
xnor U2523 (N_2523,In_1252,In_1098);
or U2524 (N_2524,In_763,In_452);
or U2525 (N_2525,In_620,In_804);
or U2526 (N_2526,In_556,In_1420);
nor U2527 (N_2527,In_340,In_1017);
or U2528 (N_2528,In_581,In_396);
xnor U2529 (N_2529,In_578,In_265);
xor U2530 (N_2530,In_542,In_187);
nand U2531 (N_2531,In_176,In_1392);
or U2532 (N_2532,In_295,In_93);
or U2533 (N_2533,In_279,In_398);
nand U2534 (N_2534,In_1201,In_29);
xor U2535 (N_2535,In_191,In_749);
and U2536 (N_2536,In_670,In_337);
nor U2537 (N_2537,In_1329,In_756);
nor U2538 (N_2538,In_292,In_904);
nor U2539 (N_2539,In_552,In_60);
nor U2540 (N_2540,In_1317,In_841);
or U2541 (N_2541,In_1488,In_161);
and U2542 (N_2542,In_858,In_610);
nor U2543 (N_2543,In_424,In_448);
nand U2544 (N_2544,In_724,In_1131);
xor U2545 (N_2545,In_527,In_410);
nor U2546 (N_2546,In_832,In_593);
and U2547 (N_2547,In_214,In_76);
or U2548 (N_2548,In_72,In_871);
nor U2549 (N_2549,In_418,In_1245);
xnor U2550 (N_2550,In_1175,In_1295);
xor U2551 (N_2551,In_873,In_636);
and U2552 (N_2552,In_1047,In_561);
xor U2553 (N_2553,In_47,In_95);
nand U2554 (N_2554,In_549,In_312);
and U2555 (N_2555,In_1206,In_637);
xnor U2556 (N_2556,In_622,In_210);
xnor U2557 (N_2557,In_1202,In_1496);
and U2558 (N_2558,In_14,In_772);
or U2559 (N_2559,In_210,In_608);
or U2560 (N_2560,In_470,In_898);
nand U2561 (N_2561,In_522,In_694);
and U2562 (N_2562,In_1330,In_90);
or U2563 (N_2563,In_236,In_395);
nand U2564 (N_2564,In_300,In_291);
xnor U2565 (N_2565,In_559,In_1270);
and U2566 (N_2566,In_224,In_765);
xor U2567 (N_2567,In_1188,In_33);
nor U2568 (N_2568,In_191,In_470);
xnor U2569 (N_2569,In_971,In_1302);
or U2570 (N_2570,In_500,In_1247);
or U2571 (N_2571,In_31,In_60);
nor U2572 (N_2572,In_847,In_1387);
and U2573 (N_2573,In_333,In_1036);
or U2574 (N_2574,In_1397,In_510);
and U2575 (N_2575,In_1087,In_494);
xor U2576 (N_2576,In_1371,In_883);
nand U2577 (N_2577,In_1356,In_1250);
or U2578 (N_2578,In_1068,In_876);
nor U2579 (N_2579,In_358,In_486);
nand U2580 (N_2580,In_657,In_152);
nor U2581 (N_2581,In_1299,In_980);
nand U2582 (N_2582,In_283,In_1188);
xnor U2583 (N_2583,In_1370,In_1089);
xnor U2584 (N_2584,In_171,In_222);
nor U2585 (N_2585,In_1149,In_1475);
or U2586 (N_2586,In_1099,In_1037);
or U2587 (N_2587,In_172,In_1214);
nor U2588 (N_2588,In_1384,In_1361);
and U2589 (N_2589,In_1112,In_36);
and U2590 (N_2590,In_311,In_636);
and U2591 (N_2591,In_1310,In_83);
nand U2592 (N_2592,In_555,In_702);
xor U2593 (N_2593,In_1173,In_1218);
xor U2594 (N_2594,In_460,In_1140);
nor U2595 (N_2595,In_69,In_1057);
nand U2596 (N_2596,In_342,In_763);
or U2597 (N_2597,In_1311,In_982);
and U2598 (N_2598,In_1194,In_514);
nor U2599 (N_2599,In_878,In_945);
xor U2600 (N_2600,In_0,In_354);
or U2601 (N_2601,In_761,In_711);
nor U2602 (N_2602,In_402,In_382);
and U2603 (N_2603,In_1466,In_1102);
nand U2604 (N_2604,In_777,In_702);
and U2605 (N_2605,In_1210,In_441);
and U2606 (N_2606,In_1038,In_11);
nand U2607 (N_2607,In_497,In_144);
and U2608 (N_2608,In_300,In_122);
nand U2609 (N_2609,In_1382,In_295);
xor U2610 (N_2610,In_1083,In_123);
xor U2611 (N_2611,In_1392,In_823);
nand U2612 (N_2612,In_1475,In_938);
or U2613 (N_2613,In_1249,In_157);
and U2614 (N_2614,In_1429,In_1490);
nor U2615 (N_2615,In_1018,In_592);
or U2616 (N_2616,In_338,In_1429);
and U2617 (N_2617,In_741,In_153);
and U2618 (N_2618,In_254,In_1161);
nor U2619 (N_2619,In_240,In_179);
and U2620 (N_2620,In_514,In_1404);
or U2621 (N_2621,In_694,In_83);
and U2622 (N_2622,In_144,In_913);
or U2623 (N_2623,In_770,In_36);
nor U2624 (N_2624,In_113,In_325);
xor U2625 (N_2625,In_596,In_582);
nand U2626 (N_2626,In_715,In_631);
or U2627 (N_2627,In_437,In_550);
xnor U2628 (N_2628,In_505,In_393);
nor U2629 (N_2629,In_935,In_639);
nor U2630 (N_2630,In_106,In_1454);
xnor U2631 (N_2631,In_89,In_1050);
nor U2632 (N_2632,In_1106,In_417);
nor U2633 (N_2633,In_1151,In_177);
or U2634 (N_2634,In_515,In_1205);
and U2635 (N_2635,In_687,In_992);
nand U2636 (N_2636,In_1070,In_1474);
nor U2637 (N_2637,In_971,In_869);
or U2638 (N_2638,In_1334,In_350);
nand U2639 (N_2639,In_927,In_466);
xor U2640 (N_2640,In_898,In_1398);
and U2641 (N_2641,In_1345,In_1171);
and U2642 (N_2642,In_1047,In_260);
xnor U2643 (N_2643,In_1405,In_29);
or U2644 (N_2644,In_1289,In_1076);
and U2645 (N_2645,In_138,In_1082);
and U2646 (N_2646,In_361,In_1130);
xor U2647 (N_2647,In_759,In_1423);
nor U2648 (N_2648,In_200,In_1);
nand U2649 (N_2649,In_72,In_534);
or U2650 (N_2650,In_620,In_1399);
nor U2651 (N_2651,In_591,In_1169);
nor U2652 (N_2652,In_1012,In_1225);
nand U2653 (N_2653,In_167,In_1462);
or U2654 (N_2654,In_1253,In_1150);
nor U2655 (N_2655,In_1255,In_816);
and U2656 (N_2656,In_959,In_1166);
nand U2657 (N_2657,In_660,In_732);
nor U2658 (N_2658,In_107,In_1132);
nand U2659 (N_2659,In_1236,In_594);
or U2660 (N_2660,In_522,In_539);
or U2661 (N_2661,In_398,In_69);
nand U2662 (N_2662,In_220,In_229);
and U2663 (N_2663,In_282,In_1355);
and U2664 (N_2664,In_379,In_76);
nor U2665 (N_2665,In_507,In_324);
nand U2666 (N_2666,In_1409,In_86);
nand U2667 (N_2667,In_193,In_803);
or U2668 (N_2668,In_731,In_1399);
or U2669 (N_2669,In_345,In_575);
and U2670 (N_2670,In_209,In_586);
xnor U2671 (N_2671,In_694,In_1257);
nor U2672 (N_2672,In_207,In_106);
or U2673 (N_2673,In_1292,In_1036);
nand U2674 (N_2674,In_136,In_438);
and U2675 (N_2675,In_965,In_1379);
and U2676 (N_2676,In_1381,In_1410);
or U2677 (N_2677,In_655,In_766);
nor U2678 (N_2678,In_1393,In_109);
nand U2679 (N_2679,In_1281,In_1189);
or U2680 (N_2680,In_1008,In_1265);
or U2681 (N_2681,In_689,In_870);
nand U2682 (N_2682,In_230,In_710);
xnor U2683 (N_2683,In_569,In_1425);
nand U2684 (N_2684,In_389,In_617);
nand U2685 (N_2685,In_859,In_1205);
nor U2686 (N_2686,In_130,In_879);
nor U2687 (N_2687,In_842,In_1228);
nor U2688 (N_2688,In_464,In_1445);
and U2689 (N_2689,In_618,In_1009);
and U2690 (N_2690,In_1420,In_1109);
nor U2691 (N_2691,In_1427,In_1108);
xnor U2692 (N_2692,In_919,In_123);
or U2693 (N_2693,In_1419,In_442);
nor U2694 (N_2694,In_547,In_960);
and U2695 (N_2695,In_365,In_830);
and U2696 (N_2696,In_676,In_1133);
nand U2697 (N_2697,In_1096,In_1467);
xor U2698 (N_2698,In_865,In_1199);
or U2699 (N_2699,In_621,In_445);
xnor U2700 (N_2700,In_1055,In_1366);
or U2701 (N_2701,In_717,In_1293);
nor U2702 (N_2702,In_217,In_666);
and U2703 (N_2703,In_151,In_121);
nor U2704 (N_2704,In_726,In_1061);
xnor U2705 (N_2705,In_1158,In_932);
nor U2706 (N_2706,In_626,In_936);
nand U2707 (N_2707,In_909,In_1139);
nand U2708 (N_2708,In_126,In_212);
nand U2709 (N_2709,In_202,In_514);
nor U2710 (N_2710,In_520,In_201);
nand U2711 (N_2711,In_189,In_362);
nand U2712 (N_2712,In_1454,In_1156);
xor U2713 (N_2713,In_46,In_706);
nor U2714 (N_2714,In_1460,In_1461);
or U2715 (N_2715,In_356,In_86);
nand U2716 (N_2716,In_145,In_926);
and U2717 (N_2717,In_286,In_969);
and U2718 (N_2718,In_304,In_1117);
and U2719 (N_2719,In_656,In_648);
xor U2720 (N_2720,In_811,In_1407);
and U2721 (N_2721,In_165,In_1274);
xor U2722 (N_2722,In_1156,In_1276);
nor U2723 (N_2723,In_141,In_887);
xnor U2724 (N_2724,In_575,In_144);
xnor U2725 (N_2725,In_422,In_1378);
and U2726 (N_2726,In_219,In_1332);
xnor U2727 (N_2727,In_1339,In_1459);
and U2728 (N_2728,In_1424,In_827);
nor U2729 (N_2729,In_1489,In_502);
nor U2730 (N_2730,In_147,In_820);
and U2731 (N_2731,In_74,In_1082);
nor U2732 (N_2732,In_1039,In_1387);
and U2733 (N_2733,In_1317,In_1034);
and U2734 (N_2734,In_118,In_535);
xor U2735 (N_2735,In_940,In_362);
nand U2736 (N_2736,In_1374,In_1068);
nor U2737 (N_2737,In_681,In_657);
xnor U2738 (N_2738,In_4,In_1249);
nand U2739 (N_2739,In_360,In_650);
xnor U2740 (N_2740,In_1369,In_977);
or U2741 (N_2741,In_622,In_916);
and U2742 (N_2742,In_294,In_530);
nand U2743 (N_2743,In_687,In_496);
xnor U2744 (N_2744,In_1025,In_394);
or U2745 (N_2745,In_593,In_564);
nor U2746 (N_2746,In_1153,In_732);
xnor U2747 (N_2747,In_1285,In_1090);
or U2748 (N_2748,In_777,In_804);
or U2749 (N_2749,In_1158,In_1495);
or U2750 (N_2750,In_1432,In_849);
nand U2751 (N_2751,In_1267,In_212);
nor U2752 (N_2752,In_778,In_1390);
and U2753 (N_2753,In_1451,In_9);
and U2754 (N_2754,In_1191,In_1339);
nor U2755 (N_2755,In_1380,In_1422);
and U2756 (N_2756,In_1313,In_852);
and U2757 (N_2757,In_1035,In_457);
nand U2758 (N_2758,In_591,In_1308);
and U2759 (N_2759,In_1294,In_1024);
nand U2760 (N_2760,In_870,In_1254);
or U2761 (N_2761,In_1317,In_723);
xor U2762 (N_2762,In_1461,In_995);
or U2763 (N_2763,In_764,In_600);
or U2764 (N_2764,In_63,In_42);
nor U2765 (N_2765,In_73,In_666);
nor U2766 (N_2766,In_689,In_398);
or U2767 (N_2767,In_1255,In_841);
nor U2768 (N_2768,In_1373,In_821);
nor U2769 (N_2769,In_221,In_292);
xor U2770 (N_2770,In_700,In_67);
and U2771 (N_2771,In_656,In_1126);
nor U2772 (N_2772,In_250,In_472);
xor U2773 (N_2773,In_157,In_674);
xnor U2774 (N_2774,In_362,In_466);
nor U2775 (N_2775,In_1403,In_1269);
xnor U2776 (N_2776,In_584,In_782);
or U2777 (N_2777,In_638,In_886);
nand U2778 (N_2778,In_1397,In_1377);
and U2779 (N_2779,In_889,In_308);
and U2780 (N_2780,In_714,In_890);
xnor U2781 (N_2781,In_40,In_1188);
nand U2782 (N_2782,In_570,In_872);
nor U2783 (N_2783,In_951,In_1293);
or U2784 (N_2784,In_159,In_536);
or U2785 (N_2785,In_588,In_905);
and U2786 (N_2786,In_1396,In_1156);
nor U2787 (N_2787,In_1328,In_1237);
nand U2788 (N_2788,In_844,In_664);
xnor U2789 (N_2789,In_17,In_722);
nand U2790 (N_2790,In_771,In_812);
or U2791 (N_2791,In_1350,In_122);
nand U2792 (N_2792,In_380,In_470);
or U2793 (N_2793,In_1307,In_281);
or U2794 (N_2794,In_282,In_1344);
nor U2795 (N_2795,In_352,In_732);
and U2796 (N_2796,In_975,In_283);
or U2797 (N_2797,In_660,In_1138);
or U2798 (N_2798,In_841,In_892);
nor U2799 (N_2799,In_29,In_979);
xor U2800 (N_2800,In_1227,In_980);
xnor U2801 (N_2801,In_371,In_1152);
xor U2802 (N_2802,In_1009,In_1327);
or U2803 (N_2803,In_508,In_1466);
xor U2804 (N_2804,In_604,In_865);
and U2805 (N_2805,In_320,In_175);
nand U2806 (N_2806,In_1108,In_1342);
nor U2807 (N_2807,In_790,In_1229);
nor U2808 (N_2808,In_1272,In_856);
nand U2809 (N_2809,In_1172,In_191);
or U2810 (N_2810,In_1475,In_1108);
and U2811 (N_2811,In_986,In_1145);
and U2812 (N_2812,In_1128,In_1405);
and U2813 (N_2813,In_1006,In_39);
and U2814 (N_2814,In_351,In_1277);
and U2815 (N_2815,In_133,In_567);
nand U2816 (N_2816,In_1377,In_1362);
xnor U2817 (N_2817,In_27,In_970);
nor U2818 (N_2818,In_1444,In_123);
nor U2819 (N_2819,In_180,In_576);
nand U2820 (N_2820,In_1449,In_233);
and U2821 (N_2821,In_198,In_219);
xnor U2822 (N_2822,In_1119,In_665);
and U2823 (N_2823,In_1388,In_1258);
nand U2824 (N_2824,In_144,In_479);
or U2825 (N_2825,In_1238,In_1291);
xor U2826 (N_2826,In_1135,In_373);
or U2827 (N_2827,In_401,In_360);
nor U2828 (N_2828,In_924,In_545);
xor U2829 (N_2829,In_1280,In_335);
nand U2830 (N_2830,In_1193,In_336);
nor U2831 (N_2831,In_156,In_328);
nand U2832 (N_2832,In_1381,In_961);
and U2833 (N_2833,In_542,In_646);
or U2834 (N_2834,In_896,In_866);
nor U2835 (N_2835,In_874,In_55);
and U2836 (N_2836,In_1212,In_449);
or U2837 (N_2837,In_207,In_285);
and U2838 (N_2838,In_890,In_1389);
xnor U2839 (N_2839,In_973,In_1467);
nand U2840 (N_2840,In_1173,In_822);
nor U2841 (N_2841,In_822,In_101);
and U2842 (N_2842,In_355,In_653);
and U2843 (N_2843,In_666,In_421);
nor U2844 (N_2844,In_1160,In_820);
nor U2845 (N_2845,In_1252,In_224);
and U2846 (N_2846,In_120,In_153);
and U2847 (N_2847,In_419,In_1321);
nand U2848 (N_2848,In_148,In_71);
nor U2849 (N_2849,In_373,In_400);
nand U2850 (N_2850,In_608,In_436);
and U2851 (N_2851,In_46,In_1304);
nor U2852 (N_2852,In_620,In_780);
xor U2853 (N_2853,In_139,In_634);
nor U2854 (N_2854,In_1002,In_859);
and U2855 (N_2855,In_204,In_10);
xnor U2856 (N_2856,In_900,In_852);
nor U2857 (N_2857,In_1118,In_529);
xnor U2858 (N_2858,In_1177,In_304);
nor U2859 (N_2859,In_127,In_966);
and U2860 (N_2860,In_605,In_393);
or U2861 (N_2861,In_529,In_539);
nor U2862 (N_2862,In_625,In_1086);
and U2863 (N_2863,In_1302,In_61);
xnor U2864 (N_2864,In_1104,In_1057);
xor U2865 (N_2865,In_1025,In_450);
and U2866 (N_2866,In_332,In_1048);
or U2867 (N_2867,In_761,In_486);
or U2868 (N_2868,In_1066,In_1367);
xor U2869 (N_2869,In_105,In_583);
or U2870 (N_2870,In_901,In_1103);
xnor U2871 (N_2871,In_213,In_336);
xnor U2872 (N_2872,In_990,In_572);
xnor U2873 (N_2873,In_1359,In_914);
and U2874 (N_2874,In_665,In_435);
nor U2875 (N_2875,In_276,In_1240);
nor U2876 (N_2876,In_740,In_187);
xnor U2877 (N_2877,In_313,In_637);
and U2878 (N_2878,In_1448,In_1377);
xor U2879 (N_2879,In_1026,In_876);
nor U2880 (N_2880,In_645,In_1149);
nand U2881 (N_2881,In_25,In_151);
and U2882 (N_2882,In_10,In_345);
nor U2883 (N_2883,In_880,In_1381);
and U2884 (N_2884,In_48,In_250);
or U2885 (N_2885,In_1440,In_419);
nor U2886 (N_2886,In_1454,In_896);
and U2887 (N_2887,In_201,In_1100);
xor U2888 (N_2888,In_177,In_1058);
and U2889 (N_2889,In_304,In_362);
or U2890 (N_2890,In_1056,In_1335);
nor U2891 (N_2891,In_238,In_1460);
or U2892 (N_2892,In_13,In_872);
and U2893 (N_2893,In_1092,In_198);
xnor U2894 (N_2894,In_1309,In_1344);
and U2895 (N_2895,In_1163,In_1057);
xor U2896 (N_2896,In_1496,In_1224);
nand U2897 (N_2897,In_878,In_1309);
and U2898 (N_2898,In_546,In_522);
nor U2899 (N_2899,In_1056,In_1201);
nor U2900 (N_2900,In_703,In_840);
xor U2901 (N_2901,In_1124,In_1445);
and U2902 (N_2902,In_1178,In_841);
and U2903 (N_2903,In_774,In_77);
nand U2904 (N_2904,In_698,In_86);
nor U2905 (N_2905,In_376,In_389);
nor U2906 (N_2906,In_737,In_718);
xnor U2907 (N_2907,In_639,In_380);
nand U2908 (N_2908,In_722,In_629);
nand U2909 (N_2909,In_637,In_1438);
and U2910 (N_2910,In_1485,In_9);
nand U2911 (N_2911,In_466,In_360);
or U2912 (N_2912,In_23,In_1227);
nor U2913 (N_2913,In_662,In_689);
and U2914 (N_2914,In_165,In_1255);
and U2915 (N_2915,In_1305,In_124);
nor U2916 (N_2916,In_935,In_498);
xor U2917 (N_2917,In_1343,In_713);
xor U2918 (N_2918,In_865,In_188);
and U2919 (N_2919,In_1272,In_808);
and U2920 (N_2920,In_1041,In_1392);
nand U2921 (N_2921,In_1254,In_1133);
nor U2922 (N_2922,In_876,In_839);
nor U2923 (N_2923,In_859,In_233);
or U2924 (N_2924,In_424,In_473);
nand U2925 (N_2925,In_811,In_199);
and U2926 (N_2926,In_210,In_1154);
and U2927 (N_2927,In_1355,In_28);
and U2928 (N_2928,In_368,In_141);
nand U2929 (N_2929,In_1301,In_634);
xor U2930 (N_2930,In_257,In_688);
nand U2931 (N_2931,In_42,In_198);
xor U2932 (N_2932,In_680,In_234);
nand U2933 (N_2933,In_1275,In_1307);
xnor U2934 (N_2934,In_998,In_228);
nand U2935 (N_2935,In_524,In_574);
nand U2936 (N_2936,In_1257,In_1414);
nor U2937 (N_2937,In_1469,In_900);
xor U2938 (N_2938,In_846,In_370);
nor U2939 (N_2939,In_1326,In_1299);
or U2940 (N_2940,In_518,In_1296);
nand U2941 (N_2941,In_38,In_1400);
nor U2942 (N_2942,In_4,In_1287);
and U2943 (N_2943,In_629,In_1208);
or U2944 (N_2944,In_331,In_813);
or U2945 (N_2945,In_1343,In_31);
nand U2946 (N_2946,In_643,In_1445);
nor U2947 (N_2947,In_1436,In_575);
nand U2948 (N_2948,In_822,In_275);
nor U2949 (N_2949,In_1045,In_1);
nor U2950 (N_2950,In_225,In_1042);
nor U2951 (N_2951,In_1160,In_1145);
nor U2952 (N_2952,In_339,In_1073);
and U2953 (N_2953,In_734,In_694);
nand U2954 (N_2954,In_1388,In_1348);
or U2955 (N_2955,In_1329,In_50);
nor U2956 (N_2956,In_1431,In_1334);
or U2957 (N_2957,In_1302,In_524);
or U2958 (N_2958,In_554,In_1426);
xor U2959 (N_2959,In_1007,In_423);
or U2960 (N_2960,In_178,In_1105);
xor U2961 (N_2961,In_393,In_806);
or U2962 (N_2962,In_109,In_631);
or U2963 (N_2963,In_523,In_1281);
xor U2964 (N_2964,In_648,In_1007);
nor U2965 (N_2965,In_611,In_929);
and U2966 (N_2966,In_670,In_185);
and U2967 (N_2967,In_360,In_85);
or U2968 (N_2968,In_160,In_1429);
nor U2969 (N_2969,In_639,In_690);
xor U2970 (N_2970,In_785,In_627);
nor U2971 (N_2971,In_1037,In_489);
and U2972 (N_2972,In_246,In_351);
nor U2973 (N_2973,In_237,In_110);
and U2974 (N_2974,In_459,In_508);
xor U2975 (N_2975,In_124,In_155);
xor U2976 (N_2976,In_122,In_695);
and U2977 (N_2977,In_944,In_1126);
xor U2978 (N_2978,In_1061,In_1170);
nor U2979 (N_2979,In_147,In_20);
and U2980 (N_2980,In_846,In_1362);
xor U2981 (N_2981,In_51,In_952);
nor U2982 (N_2982,In_709,In_1199);
and U2983 (N_2983,In_1297,In_140);
xor U2984 (N_2984,In_1394,In_620);
nand U2985 (N_2985,In_248,In_444);
nor U2986 (N_2986,In_697,In_460);
xnor U2987 (N_2987,In_885,In_130);
or U2988 (N_2988,In_829,In_565);
nor U2989 (N_2989,In_677,In_1234);
nand U2990 (N_2990,In_952,In_760);
nor U2991 (N_2991,In_633,In_1076);
nand U2992 (N_2992,In_547,In_205);
xnor U2993 (N_2993,In_897,In_1033);
or U2994 (N_2994,In_1477,In_1285);
xnor U2995 (N_2995,In_1304,In_825);
or U2996 (N_2996,In_529,In_1003);
nor U2997 (N_2997,In_747,In_275);
nand U2998 (N_2998,In_1139,In_196);
and U2999 (N_2999,In_1056,In_23);
nand U3000 (N_3000,N_766,N_2874);
or U3001 (N_3001,N_1021,N_1432);
nor U3002 (N_3002,N_2598,N_2901);
nand U3003 (N_3003,N_2805,N_2581);
or U3004 (N_3004,N_112,N_30);
xnor U3005 (N_3005,N_489,N_2129);
or U3006 (N_3006,N_2984,N_1273);
xor U3007 (N_3007,N_2462,N_6);
xor U3008 (N_3008,N_744,N_2387);
and U3009 (N_3009,N_1075,N_2491);
and U3010 (N_3010,N_1934,N_222);
nor U3011 (N_3011,N_2839,N_331);
nor U3012 (N_3012,N_596,N_384);
and U3013 (N_3013,N_834,N_1914);
xnor U3014 (N_3014,N_2599,N_2687);
nor U3015 (N_3015,N_93,N_2006);
or U3016 (N_3016,N_767,N_519);
and U3017 (N_3017,N_2047,N_994);
and U3018 (N_3018,N_1718,N_1197);
xor U3019 (N_3019,N_1611,N_820);
and U3020 (N_3020,N_1307,N_2394);
xnor U3021 (N_3021,N_975,N_2423);
and U3022 (N_3022,N_2681,N_2001);
or U3023 (N_3023,N_1685,N_1347);
nand U3024 (N_3024,N_1101,N_409);
nor U3025 (N_3025,N_2999,N_2054);
nor U3026 (N_3026,N_2079,N_238);
or U3027 (N_3027,N_2171,N_2186);
nor U3028 (N_3028,N_522,N_1560);
nor U3029 (N_3029,N_143,N_429);
or U3030 (N_3030,N_1779,N_2773);
nand U3031 (N_3031,N_45,N_2700);
xor U3032 (N_3032,N_1696,N_2362);
or U3033 (N_3033,N_598,N_1688);
and U3034 (N_3034,N_534,N_1339);
and U3035 (N_3035,N_1567,N_2502);
and U3036 (N_3036,N_1707,N_1742);
or U3037 (N_3037,N_2865,N_2673);
xor U3038 (N_3038,N_1580,N_1951);
or U3039 (N_3039,N_2489,N_2657);
xnor U3040 (N_3040,N_1698,N_504);
nand U3041 (N_3041,N_769,N_746);
and U3042 (N_3042,N_1584,N_869);
nand U3043 (N_3043,N_2081,N_2671);
and U3044 (N_3044,N_1073,N_548);
xor U3045 (N_3045,N_661,N_2490);
nor U3046 (N_3046,N_179,N_2090);
and U3047 (N_3047,N_1806,N_458);
and U3048 (N_3048,N_776,N_1332);
xnor U3049 (N_3049,N_1755,N_590);
xnor U3050 (N_3050,N_898,N_2842);
or U3051 (N_3051,N_1917,N_672);
and U3052 (N_3052,N_2796,N_56);
nand U3053 (N_3053,N_2416,N_1081);
nor U3054 (N_3054,N_1777,N_2468);
or U3055 (N_3055,N_2167,N_1165);
or U3056 (N_3056,N_2688,N_1336);
nor U3057 (N_3057,N_609,N_2937);
nor U3058 (N_3058,N_209,N_2528);
and U3059 (N_3059,N_2152,N_271);
xor U3060 (N_3060,N_2968,N_1299);
and U3061 (N_3061,N_211,N_68);
or U3062 (N_3062,N_91,N_1470);
and U3063 (N_3063,N_2093,N_1618);
or U3064 (N_3064,N_1943,N_2544);
xor U3065 (N_3065,N_1158,N_1818);
or U3066 (N_3066,N_1897,N_1515);
and U3067 (N_3067,N_33,N_58);
nor U3068 (N_3068,N_582,N_2885);
nand U3069 (N_3069,N_150,N_2941);
or U3070 (N_3070,N_1061,N_2385);
nand U3071 (N_3071,N_2082,N_796);
nor U3072 (N_3072,N_76,N_2086);
and U3073 (N_3073,N_1553,N_1517);
nor U3074 (N_3074,N_2738,N_963);
and U3075 (N_3075,N_968,N_1913);
nand U3076 (N_3076,N_2748,N_1366);
or U3077 (N_3077,N_587,N_2721);
nor U3078 (N_3078,N_2443,N_1911);
xor U3079 (N_3079,N_871,N_248);
xnor U3080 (N_3080,N_185,N_2140);
nor U3081 (N_3081,N_5,N_1781);
nand U3082 (N_3082,N_1100,N_1672);
or U3083 (N_3083,N_390,N_2520);
or U3084 (N_3084,N_203,N_1801);
and U3085 (N_3085,N_1422,N_1286);
nor U3086 (N_3086,N_1119,N_1014);
and U3087 (N_3087,N_1555,N_2065);
nand U3088 (N_3088,N_1334,N_1945);
or U3089 (N_3089,N_2908,N_1773);
nor U3090 (N_3090,N_147,N_407);
nor U3091 (N_3091,N_2378,N_1350);
xnor U3092 (N_3092,N_98,N_278);
nor U3093 (N_3093,N_1739,N_2612);
or U3094 (N_3094,N_570,N_2098);
nand U3095 (N_3095,N_1167,N_1844);
xor U3096 (N_3096,N_2891,N_110);
nand U3097 (N_3097,N_1084,N_547);
xnor U3098 (N_3098,N_755,N_1868);
nor U3099 (N_3099,N_2932,N_155);
and U3100 (N_3100,N_2393,N_1658);
nor U3101 (N_3101,N_1207,N_2441);
or U3102 (N_3102,N_311,N_877);
nor U3103 (N_3103,N_473,N_657);
xor U3104 (N_3104,N_236,N_794);
nor U3105 (N_3105,N_856,N_892);
xnor U3106 (N_3106,N_723,N_1820);
and U3107 (N_3107,N_509,N_2388);
and U3108 (N_3108,N_2445,N_2312);
nand U3109 (N_3109,N_328,N_1068);
nand U3110 (N_3110,N_1033,N_2234);
and U3111 (N_3111,N_2960,N_40);
nand U3112 (N_3112,N_1343,N_2741);
or U3113 (N_3113,N_2419,N_2094);
nor U3114 (N_3114,N_1709,N_1208);
and U3115 (N_3115,N_1931,N_1702);
nand U3116 (N_3116,N_213,N_272);
or U3117 (N_3117,N_2498,N_2303);
nor U3118 (N_3118,N_1259,N_693);
nor U3119 (N_3119,N_2812,N_102);
nor U3120 (N_3120,N_2449,N_1850);
or U3121 (N_3121,N_475,N_2780);
xor U3122 (N_3122,N_2621,N_2845);
or U3123 (N_3123,N_2567,N_1621);
nor U3124 (N_3124,N_101,N_1487);
nor U3125 (N_3125,N_1012,N_2340);
nand U3126 (N_3126,N_1046,N_1364);
or U3127 (N_3127,N_826,N_2558);
and U3128 (N_3128,N_2304,N_690);
or U3129 (N_3129,N_1842,N_403);
nand U3130 (N_3130,N_550,N_330);
xnor U3131 (N_3131,N_1851,N_1804);
and U3132 (N_3132,N_173,N_2803);
nand U3133 (N_3133,N_1904,N_471);
and U3134 (N_3134,N_574,N_1916);
nand U3135 (N_3135,N_2726,N_1024);
nor U3136 (N_3136,N_2043,N_955);
nor U3137 (N_3137,N_1652,N_1276);
nand U3138 (N_3138,N_741,N_1952);
nor U3139 (N_3139,N_2760,N_43);
xnor U3140 (N_3140,N_1978,N_2483);
nand U3141 (N_3141,N_2176,N_2231);
nand U3142 (N_3142,N_1977,N_2871);
nor U3143 (N_3143,N_2837,N_891);
xor U3144 (N_3144,N_2359,N_1695);
nand U3145 (N_3145,N_180,N_916);
and U3146 (N_3146,N_385,N_564);
or U3147 (N_3147,N_764,N_2946);
nor U3148 (N_3148,N_2218,N_402);
or U3149 (N_3149,N_1973,N_487);
xor U3150 (N_3150,N_947,N_760);
nand U3151 (N_3151,N_616,N_608);
nor U3152 (N_3152,N_34,N_2683);
and U3153 (N_3153,N_2616,N_1132);
nand U3154 (N_3154,N_1057,N_309);
xnor U3155 (N_3155,N_1991,N_233);
or U3156 (N_3156,N_1306,N_1845);
xor U3157 (N_3157,N_901,N_2827);
nor U3158 (N_3158,N_1264,N_466);
nand U3159 (N_3159,N_1648,N_1503);
xor U3160 (N_3160,N_2767,N_2434);
or U3161 (N_3161,N_449,N_601);
or U3162 (N_3162,N_1636,N_1232);
nand U3163 (N_3163,N_1243,N_1554);
and U3164 (N_3164,N_2466,N_115);
nand U3165 (N_3165,N_1280,N_1310);
xor U3166 (N_3166,N_1242,N_2314);
xor U3167 (N_3167,N_1939,N_1179);
or U3168 (N_3168,N_531,N_630);
and U3169 (N_3169,N_1035,N_1400);
nand U3170 (N_3170,N_2686,N_1661);
and U3171 (N_3171,N_2912,N_2788);
xnor U3172 (N_3172,N_658,N_715);
xor U3173 (N_3173,N_2059,N_1980);
nand U3174 (N_3174,N_365,N_2809);
and U3175 (N_3175,N_1687,N_1572);
and U3176 (N_3176,N_2644,N_636);
nor U3177 (N_3177,N_1782,N_2372);
nor U3178 (N_3178,N_1417,N_1274);
xnor U3179 (N_3179,N_2847,N_1608);
nor U3180 (N_3180,N_2238,N_1159);
nand U3181 (N_3181,N_2624,N_2428);
and U3182 (N_3182,N_227,N_2617);
nand U3183 (N_3183,N_540,N_950);
xnor U3184 (N_3184,N_1896,N_2768);
and U3185 (N_3185,N_1963,N_2219);
or U3186 (N_3186,N_2403,N_740);
nand U3187 (N_3187,N_1301,N_1494);
nor U3188 (N_3188,N_1093,N_2830);
or U3189 (N_3189,N_1293,N_1041);
nand U3190 (N_3190,N_1747,N_2030);
nand U3191 (N_3191,N_1326,N_2050);
nor U3192 (N_3192,N_2506,N_2893);
nand U3193 (N_3193,N_2501,N_844);
xnor U3194 (N_3194,N_1095,N_2783);
xnor U3195 (N_3195,N_1632,N_2778);
nand U3196 (N_3196,N_825,N_2537);
nand U3197 (N_3197,N_1361,N_1113);
or U3198 (N_3198,N_762,N_1337);
xor U3199 (N_3199,N_1331,N_2370);
nand U3200 (N_3200,N_1313,N_2316);
or U3201 (N_3201,N_1481,N_1717);
xnor U3202 (N_3202,N_1708,N_1901);
xor U3203 (N_3203,N_1415,N_461);
xnor U3204 (N_3204,N_2199,N_474);
xnor U3205 (N_3205,N_1955,N_139);
xor U3206 (N_3206,N_1817,N_1226);
and U3207 (N_3207,N_2744,N_2677);
xor U3208 (N_3208,N_771,N_836);
nor U3209 (N_3209,N_1691,N_1087);
nor U3210 (N_3210,N_952,N_1822);
or U3211 (N_3211,N_1394,N_1783);
nor U3212 (N_3212,N_843,N_939);
nand U3213 (N_3213,N_187,N_557);
or U3214 (N_3214,N_703,N_100);
or U3215 (N_3215,N_541,N_419);
nor U3216 (N_3216,N_346,N_2763);
or U3217 (N_3217,N_1947,N_82);
or U3218 (N_3218,N_2333,N_35);
or U3219 (N_3219,N_2251,N_431);
xnor U3220 (N_3220,N_2009,N_2775);
and U3221 (N_3221,N_1209,N_2797);
nor U3222 (N_3222,N_2573,N_2203);
xor U3223 (N_3223,N_502,N_219);
and U3224 (N_3224,N_2239,N_2368);
and U3225 (N_3225,N_1144,N_1813);
nand U3226 (N_3226,N_62,N_230);
nand U3227 (N_3227,N_1460,N_2255);
xor U3228 (N_3228,N_2046,N_2751);
or U3229 (N_3229,N_1794,N_1941);
nand U3230 (N_3230,N_2354,N_1557);
nor U3231 (N_3231,N_2880,N_1492);
and U3232 (N_3232,N_435,N_2833);
xnor U3233 (N_3233,N_2456,N_2246);
or U3234 (N_3234,N_846,N_2150);
nand U3235 (N_3235,N_621,N_1859);
nand U3236 (N_3236,N_861,N_1040);
nor U3237 (N_3237,N_49,N_2352);
and U3238 (N_3238,N_2452,N_2109);
xor U3239 (N_3239,N_2976,N_711);
nand U3240 (N_3240,N_2335,N_283);
and U3241 (N_3241,N_1060,N_61);
or U3242 (N_3242,N_2052,N_1328);
and U3243 (N_3243,N_1885,N_641);
and U3244 (N_3244,N_677,N_2714);
nand U3245 (N_3245,N_1335,N_1118);
or U3246 (N_3246,N_2019,N_1835);
nor U3247 (N_3247,N_1296,N_581);
nor U3248 (N_3248,N_1305,N_592);
nand U3249 (N_3249,N_446,N_2791);
xnor U3250 (N_3250,N_1959,N_1292);
or U3251 (N_3251,N_2217,N_1569);
or U3252 (N_3252,N_2522,N_1713);
and U3253 (N_3253,N_2867,N_1103);
nor U3254 (N_3254,N_1204,N_1072);
xor U3255 (N_3255,N_104,N_2824);
or U3256 (N_3256,N_316,N_2647);
xor U3257 (N_3257,N_2407,N_759);
or U3258 (N_3258,N_255,N_1744);
nor U3259 (N_3259,N_270,N_2012);
and U3260 (N_3260,N_1112,N_1614);
or U3261 (N_3261,N_2172,N_2922);
nor U3262 (N_3262,N_152,N_618);
and U3263 (N_3263,N_2464,N_1121);
and U3264 (N_3264,N_2776,N_2425);
and U3265 (N_3265,N_1252,N_2702);
nor U3266 (N_3266,N_1593,N_650);
nor U3267 (N_3267,N_731,N_498);
and U3268 (N_3268,N_1847,N_1201);
or U3269 (N_3269,N_467,N_2602);
xor U3270 (N_3270,N_1124,N_1260);
or U3271 (N_3271,N_1427,N_2669);
and U3272 (N_3272,N_935,N_2132);
nand U3273 (N_3273,N_1027,N_2730);
nor U3274 (N_3274,N_2758,N_2073);
nor U3275 (N_3275,N_998,N_2816);
nor U3276 (N_3276,N_1171,N_2703);
xor U3277 (N_3277,N_78,N_638);
or U3278 (N_3278,N_951,N_1969);
nand U3279 (N_3279,N_917,N_896);
or U3280 (N_3280,N_606,N_1472);
and U3281 (N_3281,N_38,N_28);
xor U3282 (N_3282,N_1382,N_1541);
and U3283 (N_3283,N_1266,N_2561);
and U3284 (N_3284,N_1441,N_2247);
and U3285 (N_3285,N_1219,N_2613);
and U3286 (N_3286,N_2543,N_2244);
xnor U3287 (N_3287,N_2972,N_2765);
nor U3288 (N_3288,N_2695,N_221);
nand U3289 (N_3289,N_779,N_1458);
nor U3290 (N_3290,N_1,N_1324);
xnor U3291 (N_3291,N_2424,N_399);
xor U3292 (N_3292,N_1856,N_1876);
nor U3293 (N_3293,N_2056,N_310);
or U3294 (N_3294,N_351,N_1798);
and U3295 (N_3295,N_822,N_1297);
or U3296 (N_3296,N_734,N_728);
nand U3297 (N_3297,N_1589,N_1511);
nor U3298 (N_3298,N_2795,N_1053);
xnor U3299 (N_3299,N_456,N_727);
or U3300 (N_3300,N_1774,N_2655);
nor U3301 (N_3301,N_1290,N_459);
and U3302 (N_3302,N_1873,N_239);
and U3303 (N_3303,N_1490,N_1352);
nand U3304 (N_3304,N_1176,N_664);
and U3305 (N_3305,N_2485,N_2574);
and U3306 (N_3306,N_685,N_516);
nor U3307 (N_3307,N_51,N_1368);
and U3308 (N_3308,N_1650,N_2945);
xnor U3309 (N_3309,N_726,N_527);
xor U3310 (N_3310,N_284,N_863);
or U3311 (N_3311,N_2422,N_265);
nor U3312 (N_3312,N_1406,N_1237);
nor U3313 (N_3313,N_44,N_496);
or U3314 (N_3314,N_2162,N_517);
or U3315 (N_3315,N_2580,N_195);
nor U3316 (N_3316,N_1551,N_26);
nor U3317 (N_3317,N_2292,N_980);
and U3318 (N_3318,N_1890,N_324);
and U3319 (N_3319,N_2072,N_312);
nand U3320 (N_3320,N_1321,N_974);
and U3321 (N_3321,N_1816,N_1376);
or U3322 (N_3322,N_2310,N_973);
xnor U3323 (N_3323,N_438,N_2928);
or U3324 (N_3324,N_494,N_2823);
nand U3325 (N_3325,N_1711,N_602);
or U3326 (N_3326,N_1545,N_162);
nor U3327 (N_3327,N_2894,N_756);
nor U3328 (N_3328,N_160,N_931);
or U3329 (N_3329,N_249,N_580);
nand U3330 (N_3330,N_996,N_2849);
and U3331 (N_3331,N_2481,N_387);
xnor U3332 (N_3332,N_2963,N_671);
or U3333 (N_3333,N_1277,N_1058);
xnor U3334 (N_3334,N_1797,N_2062);
xnor U3335 (N_3335,N_1814,N_2565);
nor U3336 (N_3336,N_2646,N_937);
nand U3337 (N_3337,N_2343,N_1220);
and U3338 (N_3338,N_1079,N_1875);
or U3339 (N_3339,N_2998,N_1123);
nor U3340 (N_3340,N_1715,N_1236);
and U3341 (N_3341,N_455,N_669);
nand U3342 (N_3342,N_828,N_1495);
xnor U3343 (N_3343,N_2144,N_2044);
nor U3344 (N_3344,N_2575,N_235);
and U3345 (N_3345,N_1907,N_2037);
nor U3346 (N_3346,N_1283,N_563);
nor U3347 (N_3347,N_382,N_2027);
and U3348 (N_3348,N_194,N_1910);
xor U3349 (N_3349,N_1750,N_865);
and U3350 (N_3350,N_90,N_717);
nor U3351 (N_3351,N_1455,N_1086);
nand U3352 (N_3352,N_136,N_1054);
and U3353 (N_3353,N_1600,N_1327);
nor U3354 (N_3354,N_2774,N_2678);
and U3355 (N_3355,N_640,N_2228);
or U3356 (N_3356,N_2493,N_1651);
nor U3357 (N_3357,N_114,N_2545);
xnor U3358 (N_3358,N_588,N_543);
or U3359 (N_3359,N_1358,N_2592);
and U3360 (N_3360,N_2259,N_149);
or U3361 (N_3361,N_2318,N_1378);
and U3362 (N_3362,N_2420,N_2770);
xnor U3363 (N_3363,N_1793,N_2392);
xor U3364 (N_3364,N_1294,N_1461);
and U3365 (N_3365,N_2915,N_2366);
or U3366 (N_3366,N_1138,N_806);
nor U3367 (N_3367,N_1537,N_2273);
nand U3368 (N_3368,N_1741,N_2252);
nand U3369 (N_3369,N_2802,N_1796);
or U3370 (N_3370,N_542,N_2662);
nand U3371 (N_3371,N_785,N_1878);
nand U3372 (N_3372,N_1125,N_1463);
and U3373 (N_3373,N_1091,N_2642);
nor U3374 (N_3374,N_148,N_2974);
xor U3375 (N_3375,N_1539,N_2206);
and U3376 (N_3376,N_361,N_545);
nand U3377 (N_3377,N_2717,N_436);
or U3378 (N_3378,N_48,N_1833);
nand U3379 (N_3379,N_1933,N_2177);
nand U3380 (N_3380,N_2858,N_2028);
xor U3381 (N_3381,N_2131,N_1405);
nand U3382 (N_3382,N_634,N_457);
or U3383 (N_3383,N_1172,N_610);
or U3384 (N_3384,N_2679,N_287);
or U3385 (N_3385,N_1972,N_1202);
and U3386 (N_3386,N_1961,N_1666);
nor U3387 (N_3387,N_1949,N_873);
nor U3388 (N_3388,N_1190,N_183);
xor U3389 (N_3389,N_1623,N_2288);
nor U3390 (N_3390,N_1036,N_925);
xnor U3391 (N_3391,N_2418,N_945);
xnor U3392 (N_3392,N_840,N_477);
nand U3393 (N_3393,N_626,N_1697);
nor U3394 (N_3394,N_2672,N_1767);
and U3395 (N_3395,N_2959,N_922);
or U3396 (N_3396,N_1213,N_2952);
or U3397 (N_3397,N_2204,N_1383);
or U3398 (N_3398,N_481,N_1631);
nor U3399 (N_3399,N_2691,N_279);
nor U3400 (N_3400,N_301,N_2848);
xnor U3401 (N_3401,N_408,N_1089);
xnor U3402 (N_3402,N_2336,N_2554);
or U3403 (N_3403,N_1133,N_2486);
and U3404 (N_3404,N_560,N_275);
or U3405 (N_3405,N_2437,N_2718);
nor U3406 (N_3406,N_2693,N_1871);
nor U3407 (N_3407,N_1185,N_2249);
nor U3408 (N_3408,N_1126,N_37);
and U3409 (N_3409,N_2188,N_478);
xor U3410 (N_3410,N_16,N_644);
and U3411 (N_3411,N_454,N_2223);
nor U3412 (N_3412,N_2562,N_874);
nor U3413 (N_3413,N_24,N_2101);
and U3414 (N_3414,N_42,N_320);
nand U3415 (N_3415,N_1419,N_862);
and U3416 (N_3416,N_1177,N_2270);
or U3417 (N_3417,N_1265,N_607);
nand U3418 (N_3418,N_1606,N_134);
xor U3419 (N_3419,N_2376,N_2771);
and U3420 (N_3420,N_1444,N_2862);
or U3421 (N_3421,N_364,N_1412);
nand U3422 (N_3422,N_2185,N_629);
or U3423 (N_3423,N_2163,N_2311);
xor U3424 (N_3424,N_2148,N_1690);
nor U3425 (N_3425,N_888,N_750);
nor U3426 (N_3426,N_1740,N_2519);
nand U3427 (N_3427,N_262,N_997);
and U3428 (N_3428,N_1693,N_2619);
nor U3429 (N_3429,N_864,N_1080);
nor U3430 (N_3430,N_1604,N_959);
or U3431 (N_3431,N_2825,N_2384);
xor U3432 (N_3432,N_1319,N_289);
and U3433 (N_3433,N_347,N_1409);
nand U3434 (N_3434,N_1748,N_1625);
or U3435 (N_3435,N_2080,N_1404);
and U3436 (N_3436,N_2852,N_2237);
or U3437 (N_3437,N_2828,N_247);
or U3438 (N_3438,N_1078,N_157);
nand U3439 (N_3439,N_525,N_2367);
or U3440 (N_3440,N_1393,N_52);
nand U3441 (N_3441,N_903,N_2048);
and U3442 (N_3442,N_1971,N_2954);
nand U3443 (N_3443,N_999,N_2358);
or U3444 (N_3444,N_1626,N_366);
nand U3445 (N_3445,N_411,N_1262);
and U3446 (N_3446,N_423,N_85);
or U3447 (N_3447,N_1578,N_2942);
and U3448 (N_3448,N_899,N_2977);
and U3449 (N_3449,N_1946,N_1373);
xnor U3450 (N_3450,N_2705,N_2479);
and U3451 (N_3451,N_2016,N_710);
and U3452 (N_3452,N_1194,N_2451);
or U3453 (N_3453,N_2742,N_2787);
nor U3454 (N_3454,N_1643,N_1645);
nor U3455 (N_3455,N_821,N_538);
nor U3456 (N_3456,N_2197,N_1445);
and U3457 (N_3457,N_2690,N_1639);
nor U3458 (N_3458,N_1413,N_1789);
or U3459 (N_3459,N_374,N_2426);
nor U3460 (N_3460,N_850,N_957);
nor U3461 (N_3461,N_2421,N_954);
nand U3462 (N_3462,N_2969,N_128);
nand U3463 (N_3463,N_428,N_2542);
nor U3464 (N_3464,N_117,N_1281);
or U3465 (N_3465,N_642,N_2914);
or U3466 (N_3466,N_897,N_1716);
and U3467 (N_3467,N_909,N_1867);
xnor U3468 (N_3468,N_1304,N_1870);
and U3469 (N_3469,N_2173,N_295);
and U3470 (N_3470,N_1549,N_1023);
nand U3471 (N_3471,N_837,N_1615);
and U3472 (N_3472,N_2241,N_2463);
nand U3473 (N_3473,N_2179,N_47);
and U3474 (N_3474,N_562,N_1104);
xor U3475 (N_3475,N_323,N_445);
or U3476 (N_3476,N_604,N_1340);
xor U3477 (N_3477,N_559,N_1375);
or U3478 (N_3478,N_599,N_232);
or U3479 (N_3479,N_2448,N_924);
or U3480 (N_3480,N_1065,N_2038);
or U3481 (N_3481,N_1882,N_2040);
or U3482 (N_3482,N_824,N_371);
nand U3483 (N_3483,N_2118,N_1186);
or U3484 (N_3484,N_2844,N_2649);
nor U3485 (N_3485,N_1725,N_377);
xnor U3486 (N_3486,N_1325,N_1451);
xor U3487 (N_3487,N_2684,N_218);
and U3488 (N_3488,N_1586,N_1162);
or U3489 (N_3489,N_1956,N_2290);
xor U3490 (N_3490,N_804,N_1314);
nand U3491 (N_3491,N_2540,N_192);
xor U3492 (N_3492,N_1214,N_2017);
nand U3493 (N_3493,N_1096,N_2709);
nor U3494 (N_3494,N_2815,N_628);
nor U3495 (N_3495,N_956,N_2757);
and U3496 (N_3496,N_2650,N_165);
nor U3497 (N_3497,N_1088,N_1392);
and U3498 (N_3498,N_2088,N_1732);
nor U3499 (N_3499,N_1538,N_967);
or U3500 (N_3500,N_497,N_1734);
xnor U3501 (N_3501,N_2135,N_1523);
nor U3502 (N_3502,N_2471,N_1601);
nor U3503 (N_3503,N_362,N_2453);
xor U3504 (N_3504,N_2351,N_1221);
and U3505 (N_3505,N_2878,N_1520);
and U3506 (N_3506,N_881,N_2532);
and U3507 (N_3507,N_1902,N_1988);
xnor U3508 (N_3508,N_652,N_1482);
or U3509 (N_3509,N_1998,N_73);
nor U3510 (N_3510,N_2470,N_2725);
nand U3511 (N_3511,N_175,N_653);
xnor U3512 (N_3512,N_2117,N_551);
or U3513 (N_3513,N_732,N_2139);
or U3514 (N_3514,N_1527,N_513);
nor U3515 (N_3515,N_912,N_830);
nand U3516 (N_3516,N_2391,N_388);
xnor U3517 (N_3517,N_2454,N_2232);
nor U3518 (N_3518,N_2563,N_635);
xor U3519 (N_3519,N_1628,N_1735);
nor U3520 (N_3520,N_966,N_1838);
xnor U3521 (N_3521,N_1116,N_2353);
xnor U3522 (N_3522,N_2436,N_813);
xnor U3523 (N_3523,N_345,N_2057);
nand U3524 (N_3524,N_1056,N_1019);
xnor U3525 (N_3525,N_1927,N_783);
nand U3526 (N_3526,N_752,N_1244);
xor U3527 (N_3527,N_1028,N_810);
or U3528 (N_3528,N_1408,N_1227);
nand U3529 (N_3529,N_1083,N_2921);
and U3530 (N_3530,N_2697,N_2723);
nor U3531 (N_3531,N_2634,N_1948);
xor U3532 (N_3532,N_894,N_882);
nand U3533 (N_3533,N_1136,N_2810);
or U3534 (N_3534,N_74,N_962);
and U3535 (N_3535,N_1094,N_2003);
xnor U3536 (N_3536,N_1151,N_1908);
nor U3537 (N_3537,N_395,N_1448);
nor U3538 (N_3538,N_2786,N_14);
and U3539 (N_3539,N_1823,N_2762);
nor U3540 (N_3540,N_748,N_13);
or U3541 (N_3541,N_257,N_2444);
xor U3542 (N_3542,N_2752,N_172);
xor U3543 (N_3543,N_2410,N_1987);
or U3544 (N_3544,N_342,N_1456);
nor U3545 (N_3545,N_2517,N_355);
or U3546 (N_3546,N_2317,N_425);
xnor U3547 (N_3547,N_1267,N_141);
or U3548 (N_3548,N_2790,N_860);
nor U3549 (N_3549,N_571,N_736);
xor U3550 (N_3550,N_611,N_2704);
nand U3551 (N_3551,N_65,N_1924);
xnor U3552 (N_3552,N_226,N_1316);
and U3553 (N_3553,N_2973,N_55);
nand U3554 (N_3554,N_2594,N_2382);
nand U3555 (N_3555,N_2990,N_2821);
nand U3556 (N_3556,N_2497,N_406);
and U3557 (N_3557,N_987,N_2374);
or U3558 (N_3558,N_692,N_1760);
nor U3559 (N_3559,N_2077,N_2332);
nand U3560 (N_3560,N_1174,N_613);
and U3561 (N_3561,N_2549,N_1107);
and U3562 (N_3562,N_1686,N_178);
nand U3563 (N_3563,N_790,N_1535);
xor U3564 (N_3564,N_2983,N_2682);
and U3565 (N_3565,N_2411,N_1889);
and U3566 (N_3566,N_41,N_204);
and U3567 (N_3567,N_370,N_932);
and U3568 (N_3568,N_2198,N_2801);
or U3569 (N_3569,N_432,N_2670);
or U3570 (N_3570,N_462,N_2084);
xor U3571 (N_3571,N_349,N_1649);
nor U3572 (N_3572,N_1909,N_679);
nor U3573 (N_3573,N_2935,N_2071);
xor U3574 (N_3574,N_2018,N_1714);
xnor U3575 (N_3575,N_441,N_1329);
nand U3576 (N_3576,N_1429,N_933);
or U3577 (N_3577,N_1563,N_1756);
nand U3578 (N_3578,N_1930,N_972);
or U3579 (N_3579,N_2630,N_709);
nand U3580 (N_3580,N_1982,N_1966);
nor U3581 (N_3581,N_198,N_2338);
nand U3582 (N_3582,N_1164,N_1102);
nand U3583 (N_3583,N_849,N_400);
xor U3584 (N_3584,N_1152,N_2781);
xor U3585 (N_3585,N_886,N_1646);
and U3586 (N_3586,N_1884,N_2526);
or U3587 (N_3587,N_2339,N_2857);
xor U3588 (N_3588,N_437,N_1810);
xnor U3589 (N_3589,N_521,N_67);
or U3590 (N_3590,N_1425,N_880);
and U3591 (N_3591,N_649,N_1513);
and U3592 (N_3592,N_1200,N_2987);
xnor U3593 (N_3593,N_243,N_1938);
xor U3594 (N_3594,N_1670,N_1001);
nand U3595 (N_3595,N_2579,N_1986);
nand U3596 (N_3596,N_1067,N_2296);
nor U3597 (N_3597,N_763,N_1762);
or U3598 (N_3598,N_2205,N_1459);
or U3599 (N_3599,N_904,N_1807);
or U3600 (N_3600,N_720,N_121);
nor U3601 (N_3601,N_2123,N_2355);
and U3602 (N_3602,N_367,N_1270);
and U3603 (N_3603,N_2895,N_2663);
nor U3604 (N_3604,N_2794,N_743);
nand U3605 (N_3605,N_1426,N_1731);
nand U3606 (N_3606,N_673,N_1852);
nor U3607 (N_3607,N_2527,N_159);
nand U3608 (N_3608,N_1043,N_27);
or U3609 (N_3609,N_1768,N_2034);
or U3610 (N_3610,N_920,N_2638);
or U3611 (N_3611,N_174,N_2923);
nand U3612 (N_3612,N_1524,N_857);
nand U3613 (N_3613,N_1547,N_1320);
nand U3614 (N_3614,N_1753,N_2138);
nor U3615 (N_3615,N_2322,N_1598);
or U3616 (N_3616,N_512,N_1016);
nand U3617 (N_3617,N_631,N_1500);
nand U3618 (N_3618,N_2089,N_1674);
or U3619 (N_3619,N_2873,N_1240);
and U3620 (N_3620,N_958,N_2277);
or U3621 (N_3621,N_176,N_702);
nand U3622 (N_3622,N_847,N_137);
xnor U3623 (N_3623,N_2566,N_1721);
or U3624 (N_3624,N_2550,N_855);
nor U3625 (N_3625,N_2329,N_2728);
and U3626 (N_3626,N_1263,N_1788);
nand U3627 (N_3627,N_1241,N_1255);
nor U3628 (N_3628,N_1430,N_697);
xnor U3629 (N_3629,N_123,N_1020);
and U3630 (N_3630,N_2525,N_142);
xor U3631 (N_3631,N_439,N_2078);
nor U3632 (N_3632,N_2518,N_1477);
and U3633 (N_3633,N_444,N_1407);
nand U3634 (N_3634,N_1984,N_1724);
and U3635 (N_3635,N_495,N_383);
or U3636 (N_3636,N_81,N_867);
nor U3637 (N_3637,N_1011,N_103);
and U3638 (N_3638,N_2882,N_18);
and U3639 (N_3639,N_708,N_651);
or U3640 (N_3640,N_2263,N_1855);
nor U3641 (N_3641,N_1926,N_2800);
and U3642 (N_3642,N_1387,N_1225);
nand U3643 (N_3643,N_2007,N_1609);
or U3644 (N_3644,N_1157,N_2021);
nand U3645 (N_3645,N_1542,N_948);
and U3646 (N_3646,N_2720,N_424);
nand U3647 (N_3647,N_1275,N_2902);
nor U3648 (N_3648,N_2590,N_2291);
nor U3649 (N_3649,N_984,N_1218);
or U3650 (N_3650,N_2779,N_694);
nand U3651 (N_3651,N_196,N_2108);
xor U3652 (N_3652,N_2210,N_21);
or U3653 (N_3653,N_2804,N_1681);
nor U3654 (N_3654,N_25,N_1860);
nand U3655 (N_3655,N_885,N_707);
xnor U3656 (N_3656,N_39,N_724);
and U3657 (N_3657,N_1992,N_2813);
xor U3658 (N_3658,N_225,N_2930);
xnor U3659 (N_3659,N_273,N_2597);
nand U3660 (N_3660,N_22,N_2835);
nand U3661 (N_3661,N_906,N_2276);
xor U3662 (N_3662,N_164,N_373);
xnor U3663 (N_3663,N_1866,N_1210);
or U3664 (N_3664,N_1345,N_1092);
xnor U3665 (N_3665,N_1997,N_1215);
nor U3666 (N_3666,N_1704,N_1278);
and U3667 (N_3667,N_815,N_2271);
nor U3668 (N_3668,N_140,N_572);
or U3669 (N_3669,N_4,N_1574);
nor U3670 (N_3670,N_1433,N_2851);
nand U3671 (N_3671,N_624,N_1269);
xor U3672 (N_3672,N_2499,N_126);
and U3673 (N_3673,N_1981,N_961);
nor U3674 (N_3674,N_259,N_2735);
nand U3675 (N_3675,N_443,N_2166);
and U3676 (N_3676,N_1367,N_2534);
nor U3677 (N_3677,N_511,N_772);
nor U3678 (N_3678,N_721,N_2785);
and U3679 (N_3679,N_1754,N_2295);
and U3680 (N_3680,N_2261,N_1638);
xnor U3681 (N_3681,N_391,N_214);
xnor U3682 (N_3682,N_1333,N_1468);
or U3683 (N_3683,N_1447,N_2666);
xor U3684 (N_3684,N_280,N_2130);
nand U3685 (N_3685,N_1780,N_1139);
and U3686 (N_3686,N_1131,N_2157);
or U3687 (N_3687,N_2267,N_182);
nor U3688 (N_3688,N_167,N_1443);
xor U3689 (N_3689,N_2412,N_1017);
or U3690 (N_3690,N_854,N_818);
nor U3691 (N_3691,N_1710,N_337);
nand U3692 (N_3692,N_1667,N_802);
nand U3693 (N_3693,N_1010,N_2096);
xnor U3694 (N_3694,N_1752,N_77);
or U3695 (N_3695,N_1983,N_1839);
and U3696 (N_3696,N_1117,N_2287);
and U3697 (N_3697,N_2899,N_2482);
or U3698 (N_3698,N_851,N_2610);
nor U3699 (N_3699,N_1359,N_2603);
nand U3700 (N_3700,N_2137,N_217);
and U3701 (N_3701,N_946,N_2538);
or U3702 (N_3702,N_832,N_1288);
nor U3703 (N_3703,N_1428,N_2840);
or U3704 (N_3704,N_1418,N_2216);
xor U3705 (N_3705,N_682,N_2593);
and U3706 (N_3706,N_1925,N_812);
or U3707 (N_3707,N_2807,N_2400);
xnor U3708 (N_3708,N_161,N_990);
xor U3709 (N_3709,N_87,N_2749);
nand U3710 (N_3710,N_1390,N_1489);
and U3711 (N_3711,N_2248,N_1525);
and U3712 (N_3712,N_2377,N_299);
nand U3713 (N_3713,N_2654,N_2903);
xnor U3714 (N_3714,N_2253,N_668);
and U3715 (N_3715,N_805,N_2986);
nand U3716 (N_3716,N_50,N_2472);
or U3717 (N_3717,N_133,N_2626);
nor U3718 (N_3718,N_695,N_2181);
nand U3719 (N_3719,N_1474,N_2282);
and U3720 (N_3720,N_2458,N_2661);
xnor U3721 (N_3721,N_2793,N_0);
and U3722 (N_3722,N_2643,N_2478);
nor U3723 (N_3723,N_656,N_1629);
nand U3724 (N_3724,N_2531,N_2427);
nand U3725 (N_3725,N_2365,N_2064);
nand U3726 (N_3726,N_2306,N_2831);
nand U3727 (N_3727,N_2888,N_1905);
nor U3728 (N_3728,N_1414,N_2026);
nand U3729 (N_3729,N_911,N_2521);
or U3730 (N_3730,N_2125,N_2147);
nor U3731 (N_3731,N_936,N_442);
or U3732 (N_3732,N_754,N_2045);
nand U3733 (N_3733,N_2722,N_1450);
and U3734 (N_3734,N_1191,N_1800);
nand U3735 (N_3735,N_1254,N_1038);
nor U3736 (N_3736,N_1562,N_2307);
and U3737 (N_3737,N_1828,N_2967);
xor U3738 (N_3738,N_2348,N_451);
and U3739 (N_3739,N_2529,N_2736);
and U3740 (N_3740,N_1802,N_1829);
nand U3741 (N_3741,N_417,N_1641);
xor U3742 (N_3742,N_537,N_2629);
nor U3743 (N_3743,N_941,N_113);
and U3744 (N_3744,N_637,N_360);
nand U3745 (N_3745,N_1808,N_730);
nor U3746 (N_3746,N_281,N_1424);
nand U3747 (N_3747,N_2864,N_1869);
and U3748 (N_3748,N_705,N_2379);
nor U3749 (N_3749,N_1247,N_1771);
and U3750 (N_3750,N_2076,N_2841);
or U3751 (N_3751,N_1233,N_2719);
xor U3752 (N_3752,N_2872,N_2927);
or U3753 (N_3753,N_1935,N_823);
and U3754 (N_3754,N_119,N_2740);
nand U3755 (N_3755,N_2694,N_1071);
nor U3756 (N_3756,N_940,N_1311);
xnor U3757 (N_3757,N_890,N_2953);
xor U3758 (N_3758,N_2881,N_2051);
xor U3759 (N_3759,N_1923,N_2910);
nand U3760 (N_3760,N_2233,N_792);
xor U3761 (N_3761,N_1395,N_2401);
xor U3762 (N_3762,N_2260,N_296);
or U3763 (N_3763,N_577,N_1624);
xor U3764 (N_3764,N_1587,N_553);
xnor U3765 (N_3765,N_1703,N_2155);
nand U3766 (N_3766,N_2201,N_2406);
and U3767 (N_3767,N_492,N_1737);
nor U3768 (N_3768,N_1386,N_71);
and U3769 (N_3769,N_207,N_2105);
nor U3770 (N_3770,N_1389,N_930);
nor U3771 (N_3771,N_875,N_2879);
or U3772 (N_3772,N_1211,N_500);
xnor U3773 (N_3773,N_1349,N_953);
and U3774 (N_3774,N_2883,N_1381);
nor U3775 (N_3775,N_453,N_322);
nand U3776 (N_3776,N_242,N_2822);
nand U3777 (N_3777,N_1843,N_277);
and U3778 (N_3778,N_1356,N_1289);
nor U3779 (N_3779,N_1423,N_1728);
xnor U3780 (N_3780,N_1238,N_2936);
xnor U3781 (N_3781,N_1958,N_2658);
and U3782 (N_3782,N_202,N_2389);
xor U3783 (N_3783,N_612,N_2754);
nor U3784 (N_3784,N_926,N_53);
nor U3785 (N_3785,N_1677,N_1954);
or U3786 (N_3786,N_2706,N_2192);
nor U3787 (N_3787,N_2608,N_1886);
and U3788 (N_3788,N_472,N_1003);
nor U3789 (N_3789,N_2811,N_2305);
and U3790 (N_3790,N_923,N_2254);
nor U3791 (N_3791,N_546,N_625);
and U3792 (N_3792,N_1683,N_1565);
xor U3793 (N_3793,N_2455,N_171);
nor U3794 (N_3794,N_491,N_23);
nor U3795 (N_3795,N_2174,N_2279);
nand U3796 (N_3796,N_507,N_2692);
xnor U3797 (N_3797,N_1025,N_895);
nor U3798 (N_3798,N_2067,N_398);
nor U3799 (N_3799,N_2402,N_1351);
nand U3800 (N_3800,N_1528,N_1746);
nor U3801 (N_3801,N_706,N_835);
nand U3802 (N_3802,N_554,N_2334);
nor U3803 (N_3803,N_158,N_2484);
nor U3804 (N_3804,N_2262,N_2087);
or U3805 (N_3805,N_2235,N_910);
nor U3806 (N_3806,N_2777,N_291);
or U3807 (N_3807,N_2906,N_808);
xor U3808 (N_3808,N_2014,N_1540);
xnor U3809 (N_3809,N_1006,N_2460);
or U3810 (N_3810,N_2230,N_757);
and U3811 (N_3811,N_1064,N_978);
nor U3812 (N_3812,N_2390,N_659);
nand U3813 (N_3813,N_2539,N_991);
xor U3814 (N_3814,N_1974,N_2178);
or U3815 (N_3815,N_1355,N_1561);
nand U3816 (N_3816,N_2503,N_2035);
or U3817 (N_3817,N_1588,N_2190);
or U3818 (N_3818,N_32,N_793);
nor U3819 (N_3819,N_2215,N_1396);
xor U3820 (N_3820,N_1501,N_1130);
xnor U3821 (N_3821,N_1594,N_340);
nor U3822 (N_3822,N_2947,N_1205);
and U3823 (N_3823,N_1438,N_94);
nor U3824 (N_3824,N_782,N_1599);
nand U3825 (N_3825,N_59,N_1543);
or U3826 (N_3826,N_983,N_2141);
and U3827 (N_3827,N_2962,N_2467);
or U3828 (N_3828,N_908,N_10);
or U3829 (N_3829,N_1573,N_2746);
or U3830 (N_3830,N_2220,N_415);
and U3831 (N_3831,N_1217,N_1007);
nand U3832 (N_3832,N_992,N_1848);
nand U3833 (N_3833,N_2508,N_2274);
nand U3834 (N_3834,N_1516,N_1673);
or U3835 (N_3835,N_156,N_1642);
nand U3836 (N_3836,N_883,N_1239);
nor U3837 (N_3837,N_92,N_1295);
nand U3838 (N_3838,N_1187,N_2008);
nand U3839 (N_3839,N_336,N_893);
nor U3840 (N_3840,N_1505,N_918);
nor U3841 (N_3841,N_240,N_1583);
or U3842 (N_3842,N_566,N_1464);
and U3843 (N_3843,N_200,N_1198);
xor U3844 (N_3844,N_1603,N_1454);
nor U3845 (N_3845,N_2733,N_584);
and U3846 (N_3846,N_2020,N_1786);
xor U3847 (N_3847,N_859,N_258);
xnor U3848 (N_3848,N_2931,N_2438);
nand U3849 (N_3849,N_681,N_985);
nand U3850 (N_3850,N_2716,N_2469);
or U3851 (N_3851,N_452,N_915);
xor U3852 (N_3852,N_2734,N_1815);
nor U3853 (N_3853,N_1607,N_2587);
xnor U3854 (N_3854,N_463,N_2031);
nor U3855 (N_3855,N_565,N_814);
nor U3856 (N_3856,N_2281,N_359);
nor U3857 (N_3857,N_1042,N_256);
xnor U3858 (N_3858,N_2321,N_1853);
nand U3859 (N_3859,N_788,N_2195);
nor U3860 (N_3860,N_2011,N_2510);
nor U3861 (N_3861,N_2727,N_2648);
or U3862 (N_3862,N_2476,N_2896);
and U3863 (N_3863,N_1519,N_1865);
nor U3864 (N_3864,N_1964,N_1059);
nor U3865 (N_3865,N_879,N_2505);
nand U3866 (N_3866,N_2364,N_64);
or U3867 (N_3867,N_1679,N_1861);
or U3868 (N_3868,N_1622,N_389);
nor U3869 (N_3869,N_1579,N_1656);
and U3870 (N_3870,N_2100,N_2949);
nand U3871 (N_3871,N_2154,N_206);
nor U3872 (N_3872,N_66,N_1531);
and U3873 (N_3873,N_1928,N_1298);
xnor U3874 (N_3874,N_845,N_2504);
or U3875 (N_3875,N_2509,N_263);
xor U3876 (N_3876,N_1880,N_1895);
or U3877 (N_3877,N_594,N_3);
xor U3878 (N_3878,N_1249,N_689);
and U3879 (N_3879,N_1013,N_1660);
nand U3880 (N_3880,N_2136,N_1077);
xnor U3881 (N_3881,N_2225,N_858);
xnor U3882 (N_3882,N_1995,N_1493);
nand U3883 (N_3883,N_2656,N_1471);
nand U3884 (N_3884,N_1827,N_276);
and U3885 (N_3885,N_597,N_1348);
xnor U3886 (N_3886,N_1354,N_878);
nor U3887 (N_3887,N_2829,N_1680);
and U3888 (N_3888,N_514,N_344);
xnor U3889 (N_3889,N_2582,N_789);
or U3890 (N_3890,N_1145,N_786);
and U3891 (N_3891,N_341,N_1581);
nor U3892 (N_3892,N_237,N_1821);
nand U3893 (N_3893,N_2951,N_2124);
or U3894 (N_3894,N_2536,N_2982);
nand U3895 (N_3895,N_2068,N_751);
xor U3896 (N_3896,N_2861,N_2060);
or U3897 (N_3897,N_737,N_303);
or U3898 (N_3898,N_2004,N_1772);
or U3899 (N_3899,N_191,N_1486);
nand U3900 (N_3900,N_615,N_2632);
xnor U3901 (N_3901,N_166,N_2515);
xnor U3902 (N_3902,N_2121,N_1129);
or U3903 (N_3903,N_1993,N_1887);
nor U3904 (N_3904,N_96,N_1114);
and U3905 (N_3905,N_704,N_1391);
or U3906 (N_3906,N_780,N_2289);
nand U3907 (N_3907,N_662,N_1824);
and U3908 (N_3908,N_1950,N_1944);
and U3909 (N_3909,N_1612,N_2395);
xnor U3910 (N_3910,N_568,N_515);
nor U3911 (N_3911,N_1671,N_2600);
nor U3912 (N_3912,N_2552,N_483);
nand U3913 (N_3913,N_1953,N_297);
and U3914 (N_3914,N_536,N_1437);
or U3915 (N_3915,N_11,N_1439);
or U3916 (N_3916,N_1775,N_2069);
and U3917 (N_3917,N_338,N_2535);
nor U3918 (N_3918,N_1689,N_1647);
or U3919 (N_3919,N_797,N_1811);
xor U3920 (N_3920,N_2667,N_1312);
nand U3921 (N_3921,N_111,N_868);
or U3922 (N_3922,N_308,N_70);
nor U3923 (N_3923,N_2911,N_1776);
nor U3924 (N_3924,N_2369,N_2889);
xor U3925 (N_3925,N_1282,N_2494);
or U3926 (N_3926,N_350,N_1467);
and U3927 (N_3927,N_1510,N_2058);
nor U3928 (N_3928,N_2513,N_354);
and U3929 (N_3929,N_2955,N_2578);
nand U3930 (N_3930,N_348,N_210);
or U3931 (N_3931,N_2156,N_1893);
and U3932 (N_3932,N_2909,N_1182);
nor U3933 (N_3933,N_2652,N_305);
and U3934 (N_3934,N_2856,N_1435);
and U3935 (N_3935,N_2584,N_2112);
xnor U3936 (N_3936,N_1898,N_2696);
nor U3937 (N_3937,N_2116,N_253);
and U3938 (N_3938,N_1769,N_2091);
xnor U3939 (N_3939,N_220,N_683);
xor U3940 (N_3940,N_1142,N_758);
xnor U3941 (N_3941,N_977,N_2200);
nor U3942 (N_3942,N_1318,N_2553);
nand U3943 (N_3943,N_2325,N_2995);
nor U3944 (N_3944,N_2211,N_648);
xnor U3945 (N_3945,N_1416,N_523);
and U3946 (N_3946,N_2053,N_2442);
and U3947 (N_3947,N_1342,N_464);
nand U3948 (N_3948,N_1730,N_949);
xnor U3949 (N_3949,N_1706,N_2913);
xor U3950 (N_3950,N_2743,N_7);
xnor U3951 (N_3951,N_2819,N_725);
nand U3952 (N_3952,N_1962,N_2350);
and U3953 (N_3953,N_2769,N_1985);
or U3954 (N_3954,N_460,N_1719);
or U3955 (N_3955,N_282,N_2375);
and U3956 (N_3956,N_1018,N_1809);
nor U3957 (N_3957,N_2347,N_942);
or U3958 (N_3958,N_2843,N_2227);
xnor U3959 (N_3959,N_396,N_2589);
nor U3960 (N_3960,N_675,N_450);
nand U3961 (N_3961,N_2897,N_1488);
nor U3962 (N_3962,N_95,N_1877);
xnor U3963 (N_3963,N_394,N_1592);
and U3964 (N_3964,N_1705,N_319);
nor U3965 (N_3965,N_1514,N_2242);
or U3966 (N_3966,N_1206,N_300);
and U3967 (N_3967,N_386,N_2061);
and U3968 (N_3968,N_405,N_1970);
nand U3969 (N_3969,N_839,N_1140);
xnor U3970 (N_3970,N_228,N_2659);
nor U3971 (N_3971,N_1184,N_1008);
or U3972 (N_3972,N_567,N_979);
and U3973 (N_3973,N_1682,N_1250);
or U3974 (N_3974,N_1291,N_2622);
xor U3975 (N_3975,N_201,N_2866);
or U3976 (N_3976,N_2461,N_2104);
nor U3977 (N_3977,N_2640,N_1109);
xor U3978 (N_3978,N_2099,N_1149);
or U3979 (N_3979,N_1385,N_1929);
xor U3980 (N_3980,N_2488,N_964);
nor U3981 (N_3981,N_2143,N_2916);
and U3982 (N_3982,N_872,N_1751);
xnor U3983 (N_3983,N_2168,N_1533);
nor U3984 (N_3984,N_1440,N_469);
nand U3985 (N_3985,N_1122,N_188);
nor U3986 (N_3986,N_2187,N_2925);
or U3987 (N_3987,N_189,N_643);
nor U3988 (N_3988,N_2789,N_2319);
nand U3989 (N_3989,N_1663,N_1229);
xor U3990 (N_3990,N_1577,N_2404);
nor U3991 (N_3991,N_2413,N_1476);
xor U3992 (N_3992,N_99,N_2323);
nand U3993 (N_3993,N_1315,N_2756);
or U3994 (N_3994,N_1353,N_2397);
and U3995 (N_3995,N_678,N_2607);
nor U3996 (N_3996,N_1410,N_2023);
nor U3997 (N_3997,N_1996,N_2556);
nor U3998 (N_3998,N_129,N_1883);
nand U3999 (N_3999,N_122,N_2417);
and U4000 (N_4000,N_1568,N_1398);
nand U4001 (N_4001,N_2063,N_2715);
xor U4002 (N_4002,N_2134,N_943);
xnor U4003 (N_4003,N_1787,N_800);
nor U4004 (N_4004,N_852,N_1617);
nor U4005 (N_4005,N_1825,N_1374);
or U4006 (N_4006,N_1317,N_2929);
or U4007 (N_4007,N_1181,N_326);
or U4008 (N_4008,N_1284,N_619);
or U4009 (N_4009,N_2836,N_1662);
and U4010 (N_4010,N_2158,N_397);
xor U4011 (N_4011,N_1189,N_2487);
or U4012 (N_4012,N_1957,N_2175);
nand U4013 (N_4013,N_46,N_2939);
nand U4014 (N_4014,N_913,N_1633);
or U4015 (N_4015,N_476,N_212);
xor U4016 (N_4016,N_1479,N_2886);
nand U4017 (N_4017,N_696,N_315);
and U4018 (N_4018,N_120,N_1738);
xnor U4019 (N_4019,N_292,N_2533);
nor U4020 (N_4020,N_866,N_241);
and U4021 (N_4021,N_1235,N_2991);
and U4022 (N_4022,N_208,N_1039);
nor U4023 (N_4023,N_2475,N_1223);
or U4024 (N_4024,N_2905,N_372);
nand U4025 (N_4025,N_1212,N_586);
nor U4026 (N_4026,N_1532,N_1676);
or U4027 (N_4027,N_2808,N_1610);
nor U4028 (N_4028,N_639,N_181);
and U4029 (N_4029,N_907,N_1341);
nand U4030 (N_4030,N_2568,N_2875);
nor U4031 (N_4031,N_1720,N_368);
or U4032 (N_4032,N_1469,N_2940);
nor U4033 (N_4033,N_2293,N_1522);
nor U4034 (N_4034,N_430,N_1231);
and U4035 (N_4035,N_2924,N_2614);
or U4036 (N_4036,N_2265,N_1402);
and U4037 (N_4037,N_2585,N_1110);
nor U4038 (N_4038,N_2943,N_1120);
nand U4039 (N_4039,N_2110,N_1224);
nor U4040 (N_4040,N_1654,N_986);
xor U4041 (N_4041,N_80,N_733);
nand U4042 (N_4042,N_2586,N_343);
or U4043 (N_4043,N_1322,N_1790);
nor U4044 (N_4044,N_1188,N_2184);
nand U4045 (N_4045,N_1785,N_1699);
or U4046 (N_4046,N_2473,N_593);
nor U4047 (N_4047,N_2283,N_97);
or U4048 (N_4048,N_2764,N_713);
xor U4049 (N_4049,N_2814,N_378);
nand U4050 (N_4050,N_2029,N_413);
nor U4051 (N_4051,N_108,N_317);
nor U4052 (N_4052,N_2191,N_1074);
nor U4053 (N_4053,N_2122,N_701);
xnor U4054 (N_4054,N_1544,N_1506);
or U4055 (N_4055,N_1245,N_1300);
and U4056 (N_4056,N_2798,N_2636);
nor U4057 (N_4057,N_186,N_381);
and U4058 (N_4058,N_2588,N_304);
and U4059 (N_4059,N_184,N_2919);
and U4060 (N_4060,N_1193,N_17);
and U4061 (N_4061,N_1279,N_2300);
and U4062 (N_4062,N_645,N_1937);
and U4063 (N_4063,N_1127,N_1484);
nand U4064 (N_4064,N_1763,N_2164);
xor U4065 (N_4065,N_2548,N_2961);
and U4066 (N_4066,N_2337,N_1653);
and U4067 (N_4067,N_817,N_72);
nor U4068 (N_4068,N_1591,N_306);
or U4069 (N_4069,N_2772,N_532);
nand U4070 (N_4070,N_753,N_1692);
and U4071 (N_4071,N_393,N_2685);
nor U4072 (N_4072,N_666,N_1090);
nand U4073 (N_4073,N_976,N_1498);
and U4074 (N_4074,N_2194,N_595);
xnor U4075 (N_4075,N_1360,N_600);
nor U4076 (N_4076,N_2817,N_2222);
and U4077 (N_4077,N_1420,N_314);
nor U4078 (N_4078,N_2732,N_2381);
and U4079 (N_4079,N_1044,N_485);
and U4080 (N_4080,N_982,N_2541);
nor U4081 (N_4081,N_1150,N_151);
and U4082 (N_4082,N_2609,N_118);
nand U4083 (N_4083,N_1529,N_1989);
nor U4084 (N_4084,N_1936,N_488);
xnor U4085 (N_4085,N_1063,N_2625);
and U4086 (N_4086,N_2214,N_2111);
xnor U4087 (N_4087,N_2944,N_1434);
nand U4088 (N_4088,N_286,N_1228);
or U4089 (N_4089,N_307,N_2102);
nand U4090 (N_4090,N_1168,N_2530);
or U4091 (N_4091,N_2430,N_960);
and U4092 (N_4092,N_1919,N_1154);
nand U4093 (N_4093,N_2707,N_927);
nand U4094 (N_4094,N_2386,N_2326);
nor U4095 (N_4095,N_1891,N_965);
nand U4096 (N_4096,N_2103,N_105);
nor U4097 (N_4097,N_2623,N_589);
nor U4098 (N_4098,N_266,N_1370);
xnor U4099 (N_4099,N_778,N_484);
or U4100 (N_4100,N_2092,N_2346);
or U4101 (N_4101,N_1082,N_884);
xnor U4102 (N_4102,N_1764,N_841);
and U4103 (N_4103,N_2414,N_2933);
nor U4104 (N_4104,N_9,N_774);
and U4105 (N_4105,N_1990,N_2591);
nand U4106 (N_4106,N_2611,N_440);
or U4107 (N_4107,N_505,N_1874);
nand U4108 (N_4108,N_2396,N_603);
or U4109 (N_4109,N_614,N_2739);
or U4110 (N_4110,N_493,N_1854);
nand U4111 (N_4111,N_1222,N_1590);
and U4112 (N_4112,N_84,N_2363);
nand U4113 (N_4113,N_2855,N_2015);
or U4114 (N_4114,N_1372,N_2275);
and U4115 (N_4115,N_1761,N_1812);
xnor U4116 (N_4116,N_2605,N_2036);
xor U4117 (N_4117,N_1736,N_2850);
or U4118 (N_4118,N_1637,N_2868);
and U4119 (N_4119,N_1285,N_1362);
nand U4120 (N_4120,N_2806,N_2258);
xor U4121 (N_4121,N_1832,N_2920);
nor U4122 (N_4122,N_2429,N_2918);
nor U4123 (N_4123,N_1881,N_2066);
and U4124 (N_4124,N_2022,N_583);
or U4125 (N_4125,N_1766,N_2309);
xnor U4126 (N_4126,N_510,N_2860);
or U4127 (N_4127,N_739,N_2245);
and U4128 (N_4128,N_1457,N_1141);
and U4129 (N_4129,N_1045,N_1616);
nand U4130 (N_4130,N_2606,N_2890);
nand U4131 (N_4131,N_914,N_2900);
or U4132 (N_4132,N_2380,N_2165);
or U4133 (N_4133,N_2480,N_2269);
or U4134 (N_4134,N_2075,N_2405);
nor U4135 (N_4135,N_900,N_2766);
xor U4136 (N_4136,N_2547,N_2877);
xor U4137 (N_4137,N_1888,N_1258);
nor U4138 (N_4138,N_131,N_2457);
xor U4139 (N_4139,N_2971,N_807);
nor U4140 (N_4140,N_1055,N_775);
nand U4141 (N_4141,N_334,N_1668);
or U4142 (N_4142,N_2755,N_2492);
or U4143 (N_4143,N_838,N_520);
nand U4144 (N_4144,N_829,N_480);
nor U4145 (N_4145,N_1192,N_718);
and U4146 (N_4146,N_1004,N_2361);
and U4147 (N_4147,N_1403,N_902);
nand U4148 (N_4148,N_1831,N_1330);
xor U4149 (N_4149,N_1115,N_1846);
nor U4150 (N_4150,N_1180,N_2938);
nand U4151 (N_4151,N_993,N_2979);
nor U4152 (N_4152,N_2383,N_1585);
nor U4153 (N_4153,N_2324,N_1526);
nor U4154 (N_4154,N_135,N_1365);
or U4155 (N_4155,N_2615,N_2285);
xor U4156 (N_4156,N_2268,N_375);
and U4157 (N_4157,N_1976,N_163);
and U4158 (N_4158,N_2115,N_654);
xnor U4159 (N_4159,N_1712,N_2884);
and U4160 (N_4160,N_2170,N_19);
xnor U4161 (N_4161,N_2032,N_1069);
and U4162 (N_4162,N_197,N_2278);
nor U4163 (N_4163,N_2224,N_1199);
nand U4164 (N_4164,N_2761,N_1146);
nor U4165 (N_4165,N_549,N_1462);
or U4166 (N_4166,N_2495,N_1302);
nand U4167 (N_4167,N_1965,N_1380);
or U4168 (N_4168,N_1849,N_2142);
and U4169 (N_4169,N_2956,N_2651);
nor U4170 (N_4170,N_622,N_2221);
and U4171 (N_4171,N_2555,N_2645);
or U4172 (N_4172,N_2859,N_1559);
and U4173 (N_4173,N_154,N_434);
nand U4174 (N_4174,N_1261,N_1701);
and U4175 (N_4175,N_2863,N_1743);
nand U4176 (N_4176,N_357,N_569);
or U4177 (N_4177,N_1512,N_700);
nor U4178 (N_4178,N_2792,N_919);
xnor U4179 (N_4179,N_2331,N_1166);
xnor U4180 (N_4180,N_8,N_981);
and U4181 (N_4181,N_1452,N_1253);
or U4182 (N_4182,N_1942,N_244);
xor U4183 (N_4183,N_663,N_1499);
or U4184 (N_4184,N_1723,N_420);
nand U4185 (N_4185,N_1234,N_2196);
nor U4186 (N_4186,N_124,N_2013);
and U4187 (N_4187,N_1729,N_418);
nand U4188 (N_4188,N_486,N_1918);
xnor U4189 (N_4189,N_2753,N_1872);
and U4190 (N_4190,N_1548,N_2981);
nor U4191 (N_4191,N_1106,N_870);
nor U4192 (N_4192,N_1085,N_1509);
nand U4193 (N_4193,N_254,N_1203);
or U4194 (N_4194,N_325,N_716);
nand U4195 (N_4195,N_1630,N_989);
or U4196 (N_4196,N_1640,N_971);
xor U4197 (N_4197,N_1694,N_1496);
nand U4198 (N_4198,N_2571,N_2846);
nor U4199 (N_4199,N_1246,N_1346);
nand U4200 (N_4200,N_798,N_138);
or U4201 (N_4201,N_1994,N_422);
nand U4202 (N_4202,N_2576,N_2557);
or U4203 (N_4203,N_579,N_1449);
nand U4204 (N_4204,N_2133,N_1862);
nand U4205 (N_4205,N_2917,N_620);
xor U4206 (N_4206,N_2948,N_801);
or U4207 (N_4207,N_1384,N_799);
nor U4208 (N_4208,N_578,N_1830);
nand U4209 (N_4209,N_2970,N_1644);
nor U4210 (N_4210,N_770,N_2898);
nand U4211 (N_4211,N_591,N_251);
nor U4212 (N_4212,N_714,N_392);
nor U4213 (N_4213,N_1502,N_2569);
or U4214 (N_4214,N_1900,N_833);
and U4215 (N_4215,N_2373,N_379);
and U4216 (N_4216,N_2272,N_2474);
xor U4217 (N_4217,N_1508,N_1147);
nand U4218 (N_4218,N_777,N_1903);
nand U4219 (N_4219,N_765,N_687);
or U4220 (N_4220,N_1634,N_827);
and U4221 (N_4221,N_660,N_2120);
nor U4222 (N_4222,N_109,N_2820);
nand U4223 (N_4223,N_2106,N_928);
or U4224 (N_4224,N_526,N_1196);
or U4225 (N_4225,N_2631,N_1047);
and U4226 (N_4226,N_2854,N_2356);
or U4227 (N_4227,N_2618,N_2371);
nand U4228 (N_4228,N_2985,N_1805);
xnor U4229 (N_4229,N_1536,N_2256);
nand U4230 (N_4230,N_1128,N_1834);
or U4231 (N_4231,N_54,N_223);
xor U4232 (N_4232,N_376,N_1722);
nand U4233 (N_4233,N_1143,N_2266);
nand U4234 (N_4234,N_132,N_2207);
nor U4235 (N_4235,N_1148,N_2523);
nor U4236 (N_4236,N_250,N_468);
nor U4237 (N_4237,N_2711,N_524);
xor U4238 (N_4238,N_2989,N_1726);
and U4239 (N_4239,N_2298,N_216);
nand U4240 (N_4240,N_1344,N_699);
nand U4241 (N_4241,N_2447,N_2978);
nor U4242 (N_4242,N_2025,N_269);
and U4243 (N_4243,N_127,N_130);
or U4244 (N_4244,N_988,N_2049);
and U4245 (N_4245,N_1411,N_1778);
nand U4246 (N_4246,N_447,N_2477);
and U4247 (N_4247,N_2055,N_2818);
xor U4248 (N_4248,N_2330,N_2993);
nor U4249 (N_4249,N_2926,N_2126);
and U4250 (N_4250,N_1156,N_2349);
nor U4251 (N_4251,N_1371,N_1575);
xnor U4252 (N_4252,N_773,N_632);
and U4253 (N_4253,N_1858,N_2183);
or U4254 (N_4254,N_199,N_1507);
nor U4255 (N_4255,N_2119,N_2907);
nand U4256 (N_4256,N_1338,N_2342);
and U4257 (N_4257,N_2731,N_1066);
and U4258 (N_4258,N_416,N_1216);
xnor U4259 (N_4259,N_2564,N_1675);
and U4260 (N_4260,N_905,N_1303);
and U4261 (N_4261,N_1550,N_921);
nand U4262 (N_4262,N_2996,N_2344);
or U4263 (N_4263,N_2750,N_1534);
nand U4264 (N_4264,N_934,N_781);
xor U4265 (N_4265,N_329,N_944);
and U4266 (N_4266,N_89,N_2674);
xnor U4267 (N_4267,N_2496,N_1022);
or U4268 (N_4268,N_246,N_2729);
or U4269 (N_4269,N_2958,N_2675);
and U4270 (N_4270,N_1169,N_2799);
or U4271 (N_4271,N_1108,N_2360);
nor U4272 (N_4272,N_2934,N_1363);
xnor U4273 (N_4273,N_2980,N_2724);
and U4274 (N_4274,N_1749,N_2151);
or U4275 (N_4275,N_1921,N_1070);
and U4276 (N_4276,N_146,N_170);
or U4277 (N_4277,N_585,N_1518);
nand U4278 (N_4278,N_2236,N_2465);
or U4279 (N_4279,N_2745,N_2992);
nor U4280 (N_4280,N_2965,N_1799);
and U4281 (N_4281,N_1175,N_302);
and U4282 (N_4282,N_1759,N_617);
or U4283 (N_4283,N_1473,N_533);
and U4284 (N_4284,N_889,N_722);
nand U4285 (N_4285,N_2964,N_426);
or U4286 (N_4286,N_2202,N_2097);
xor U4287 (N_4287,N_1613,N_60);
xnor U4288 (N_4288,N_2627,N_267);
or U4289 (N_4289,N_1491,N_2264);
xor U4290 (N_4290,N_2637,N_2433);
xor U4291 (N_4291,N_2439,N_665);
nor U4292 (N_4292,N_2668,N_106);
nor U4293 (N_4293,N_2070,N_1015);
and U4294 (N_4294,N_791,N_15);
and U4295 (N_4295,N_938,N_747);
nand U4296 (N_4296,N_887,N_2737);
nand U4297 (N_4297,N_1257,N_1478);
and U4298 (N_4298,N_2153,N_352);
nand U4299 (N_4299,N_2975,N_2);
xor U4300 (N_4300,N_647,N_1836);
or U4301 (N_4301,N_290,N_627);
nor U4302 (N_4302,N_1421,N_2341);
xnor U4303 (N_4303,N_1879,N_1657);
xor U4304 (N_4304,N_2182,N_1857);
and U4305 (N_4305,N_2193,N_1619);
nand U4306 (N_4306,N_1049,N_1727);
nor U4307 (N_4307,N_809,N_2161);
xnor U4308 (N_4308,N_555,N_2286);
xor U4309 (N_4309,N_205,N_12);
nor U4310 (N_4310,N_1230,N_2280);
or U4311 (N_4311,N_36,N_313);
nand U4312 (N_4312,N_2327,N_1308);
and U4313 (N_4313,N_1399,N_1002);
nand U4314 (N_4314,N_2966,N_544);
or U4315 (N_4315,N_623,N_680);
xor U4316 (N_4316,N_2127,N_421);
nor U4317 (N_4317,N_2665,N_260);
or U4318 (N_4318,N_2551,N_633);
xnor U4319 (N_4319,N_433,N_1357);
nand U4320 (N_4320,N_1431,N_768);
and U4321 (N_4321,N_1627,N_1521);
nand U4322 (N_4322,N_2209,N_2297);
xnor U4323 (N_4323,N_1446,N_1979);
nand U4324 (N_4324,N_876,N_499);
nand U4325 (N_4325,N_1864,N_2415);
xor U4326 (N_4326,N_1388,N_1048);
or U4327 (N_4327,N_2113,N_1178);
and U4328 (N_4328,N_1967,N_1251);
nor U4329 (N_4329,N_268,N_969);
and U4330 (N_4330,N_1899,N_2039);
nand U4331 (N_4331,N_2834,N_738);
nand U4332 (N_4332,N_2010,N_2641);
nand U4333 (N_4333,N_1602,N_2435);
nand U4334 (N_4334,N_2887,N_1436);
or U4335 (N_4335,N_63,N_929);
xor U4336 (N_4336,N_2320,N_298);
or U4337 (N_4337,N_2653,N_2159);
and U4338 (N_4338,N_1841,N_1571);
nand U4339 (N_4339,N_848,N_1795);
nand U4340 (N_4340,N_2516,N_75);
nor U4341 (N_4341,N_1453,N_2595);
nand U4342 (N_4342,N_153,N_116);
nand U4343 (N_4343,N_465,N_288);
or U4344 (N_4344,N_1552,N_745);
and U4345 (N_4345,N_2085,N_1757);
and U4346 (N_4346,N_831,N_2892);
nor U4347 (N_4347,N_2713,N_2149);
nor U4348 (N_4348,N_2146,N_1595);
or U4349 (N_4349,N_1268,N_1745);
xor U4350 (N_4350,N_1397,N_1256);
or U4351 (N_4351,N_1975,N_1111);
xor U4352 (N_4352,N_2500,N_285);
nor U4353 (N_4353,N_1826,N_2583);
or U4354 (N_4354,N_1134,N_1483);
xnor U4355 (N_4355,N_1480,N_1052);
or U4356 (N_4356,N_1605,N_1922);
and U4357 (N_4357,N_529,N_2328);
xnor U4358 (N_4358,N_2041,N_1442);
nand U4359 (N_4359,N_2432,N_1894);
nor U4360 (N_4360,N_2994,N_215);
and U4361 (N_4361,N_412,N_2832);
xor U4362 (N_4362,N_2699,N_995);
nand U4363 (N_4363,N_1009,N_1597);
xor U4364 (N_4364,N_490,N_332);
or U4365 (N_4365,N_719,N_482);
nor U4366 (N_4366,N_1465,N_803);
nand U4367 (N_4367,N_363,N_1863);
nand U4368 (N_4368,N_1765,N_528);
or U4369 (N_4369,N_2698,N_2095);
nand U4370 (N_4370,N_2226,N_1369);
or U4371 (N_4371,N_561,N_573);
nor U4372 (N_4372,N_261,N_1678);
or U4373 (N_4373,N_1029,N_427);
xnor U4374 (N_4374,N_508,N_2189);
nand U4375 (N_4375,N_2689,N_2570);
nor U4376 (N_4376,N_339,N_1635);
and U4377 (N_4377,N_735,N_686);
xnor U4378 (N_4378,N_1504,N_1475);
or U4379 (N_4379,N_2459,N_2083);
or U4380 (N_4380,N_1906,N_970);
xnor U4381 (N_4381,N_2408,N_1183);
nand U4382 (N_4382,N_2559,N_1665);
and U4383 (N_4383,N_2301,N_1596);
nor U4384 (N_4384,N_274,N_575);
and U4385 (N_4385,N_2514,N_729);
or U4386 (N_4386,N_506,N_2572);
nand U4387 (N_4387,N_1700,N_245);
and U4388 (N_4388,N_1005,N_1098);
xor U4389 (N_4389,N_79,N_556);
and U4390 (N_4390,N_1000,N_294);
nor U4391 (N_4391,N_1915,N_558);
xnor U4392 (N_4392,N_1659,N_369);
or U4393 (N_4393,N_1999,N_670);
and U4394 (N_4394,N_2398,N_691);
xnor U4395 (N_4395,N_2212,N_190);
nand U4396 (N_4396,N_1032,N_2042);
xor U4397 (N_4397,N_193,N_688);
nand U4398 (N_4398,N_1034,N_1576);
nor U4399 (N_4399,N_2169,N_742);
nand U4400 (N_4400,N_2628,N_1137);
nor U4401 (N_4401,N_2710,N_1272);
xnor U4402 (N_4402,N_2284,N_31);
xnor U4403 (N_4403,N_674,N_83);
nor U4404 (N_4404,N_321,N_2904);
nor U4405 (N_4405,N_1530,N_2431);
nand U4406 (N_4406,N_1912,N_1026);
nor U4407 (N_4407,N_2601,N_698);
xor U4408 (N_4408,N_448,N_1287);
nand U4409 (N_4409,N_1758,N_1932);
or U4410 (N_4410,N_264,N_539);
or U4411 (N_4411,N_358,N_69);
and U4412 (N_4412,N_252,N_676);
and U4413 (N_4413,N_811,N_2450);
and U4414 (N_4414,N_2950,N_168);
xnor U4415 (N_4415,N_2712,N_353);
and U4416 (N_4416,N_1155,N_646);
nand U4417 (N_4417,N_1803,N_20);
xnor U4418 (N_4418,N_2620,N_1153);
xnor U4419 (N_4419,N_1940,N_2524);
nand U4420 (N_4420,N_2033,N_2240);
xor U4421 (N_4421,N_1379,N_1669);
xnor U4422 (N_4422,N_2299,N_1497);
or U4423 (N_4423,N_380,N_2005);
nand U4424 (N_4424,N_2853,N_1620);
and U4425 (N_4425,N_1791,N_1792);
or U4426 (N_4426,N_57,N_1920);
nor U4427 (N_4427,N_853,N_2664);
nor U4428 (N_4428,N_1037,N_819);
and U4429 (N_4429,N_1076,N_335);
nand U4430 (N_4430,N_2596,N_2409);
nand U4431 (N_4431,N_2229,N_1105);
nand U4432 (N_4432,N_1566,N_1770);
and U4433 (N_4433,N_605,N_518);
or U4434 (N_4434,N_2357,N_327);
nor U4435 (N_4435,N_144,N_293);
nor U4436 (N_4436,N_749,N_2997);
or U4437 (N_4437,N_2294,N_1485);
or U4438 (N_4438,N_1960,N_1170);
nand U4439 (N_4439,N_88,N_2313);
nor U4440 (N_4440,N_1664,N_234);
nand U4441 (N_4441,N_125,N_2747);
xnor U4442 (N_4442,N_1784,N_787);
xor U4443 (N_4443,N_2446,N_2000);
nor U4444 (N_4444,N_318,N_2114);
nand U4445 (N_4445,N_503,N_2560);
or U4446 (N_4446,N_1031,N_1050);
or U4447 (N_4447,N_1570,N_177);
and U4448 (N_4448,N_2660,N_1401);
nor U4449 (N_4449,N_2145,N_795);
nand U4450 (N_4450,N_29,N_2680);
or U4451 (N_4451,N_2160,N_1173);
xor U4452 (N_4452,N_655,N_145);
xnor U4453 (N_4453,N_552,N_2826);
xor U4454 (N_4454,N_2577,N_2512);
or U4455 (N_4455,N_86,N_231);
nand U4456 (N_4456,N_1097,N_1163);
and U4457 (N_4457,N_2876,N_2869);
xor U4458 (N_4458,N_2957,N_169);
nand U4459 (N_4459,N_2243,N_2838);
nor U4460 (N_4460,N_1558,N_479);
or U4461 (N_4461,N_1030,N_2345);
nand U4462 (N_4462,N_401,N_501);
or U4463 (N_4463,N_1195,N_1556);
and U4464 (N_4464,N_1248,N_1968);
nand U4465 (N_4465,N_224,N_2440);
and U4466 (N_4466,N_404,N_1135);
nand U4467 (N_4467,N_2639,N_2180);
nor U4468 (N_4468,N_2604,N_684);
or U4469 (N_4469,N_2708,N_1323);
xnor U4470 (N_4470,N_2507,N_2208);
or U4471 (N_4471,N_410,N_2399);
and U4472 (N_4472,N_2546,N_107);
xor U4473 (N_4473,N_2074,N_2870);
or U4474 (N_4474,N_2511,N_2002);
or U4475 (N_4475,N_2759,N_842);
or U4476 (N_4476,N_2250,N_530);
xor U4477 (N_4477,N_576,N_1160);
xor U4478 (N_4478,N_1733,N_1271);
and U4479 (N_4479,N_2633,N_1546);
xnor U4480 (N_4480,N_470,N_333);
nor U4481 (N_4481,N_1684,N_1062);
xnor U4482 (N_4482,N_1564,N_1466);
nand U4483 (N_4483,N_2988,N_1840);
xor U4484 (N_4484,N_816,N_761);
xnor U4485 (N_4485,N_2635,N_2107);
nor U4486 (N_4486,N_229,N_1892);
or U4487 (N_4487,N_2784,N_1051);
nor U4488 (N_4488,N_1161,N_1377);
nand U4489 (N_4489,N_2128,N_784);
or U4490 (N_4490,N_667,N_712);
nor U4491 (N_4491,N_2676,N_414);
and U4492 (N_4492,N_2308,N_1655);
xor U4493 (N_4493,N_356,N_535);
or U4494 (N_4494,N_1819,N_2024);
and U4495 (N_4495,N_2782,N_1582);
xnor U4496 (N_4496,N_2701,N_2302);
nor U4497 (N_4497,N_2315,N_1099);
nand U4498 (N_4498,N_2257,N_1309);
and U4499 (N_4499,N_2213,N_1837);
nand U4500 (N_4500,N_1118,N_2335);
nor U4501 (N_4501,N_679,N_6);
nor U4502 (N_4502,N_977,N_2909);
xor U4503 (N_4503,N_155,N_71);
nand U4504 (N_4504,N_1360,N_2863);
nand U4505 (N_4505,N_878,N_2173);
and U4506 (N_4506,N_891,N_644);
nor U4507 (N_4507,N_1730,N_2172);
nor U4508 (N_4508,N_1107,N_772);
and U4509 (N_4509,N_1359,N_1932);
nor U4510 (N_4510,N_2481,N_1106);
nand U4511 (N_4511,N_2075,N_2644);
and U4512 (N_4512,N_2846,N_1809);
and U4513 (N_4513,N_543,N_1731);
nand U4514 (N_4514,N_1075,N_2158);
xnor U4515 (N_4515,N_1479,N_220);
or U4516 (N_4516,N_1089,N_721);
nor U4517 (N_4517,N_2926,N_1501);
xor U4518 (N_4518,N_2385,N_195);
or U4519 (N_4519,N_2523,N_2092);
nand U4520 (N_4520,N_2161,N_2950);
or U4521 (N_4521,N_174,N_232);
xor U4522 (N_4522,N_349,N_1133);
and U4523 (N_4523,N_103,N_60);
or U4524 (N_4524,N_940,N_1580);
and U4525 (N_4525,N_1783,N_2897);
nand U4526 (N_4526,N_927,N_1645);
nor U4527 (N_4527,N_250,N_2343);
or U4528 (N_4528,N_1480,N_1840);
xnor U4529 (N_4529,N_2583,N_1023);
nor U4530 (N_4530,N_423,N_1536);
nor U4531 (N_4531,N_2700,N_494);
and U4532 (N_4532,N_1923,N_107);
xnor U4533 (N_4533,N_1205,N_769);
xnor U4534 (N_4534,N_1825,N_1443);
nand U4535 (N_4535,N_1674,N_2683);
or U4536 (N_4536,N_2539,N_382);
or U4537 (N_4537,N_2843,N_2437);
nand U4538 (N_4538,N_1801,N_2204);
and U4539 (N_4539,N_2553,N_580);
xnor U4540 (N_4540,N_2495,N_2126);
and U4541 (N_4541,N_1538,N_2358);
xor U4542 (N_4542,N_947,N_156);
nand U4543 (N_4543,N_718,N_2615);
nand U4544 (N_4544,N_2651,N_424);
or U4545 (N_4545,N_841,N_538);
and U4546 (N_4546,N_1839,N_124);
xor U4547 (N_4547,N_151,N_2391);
xnor U4548 (N_4548,N_2226,N_1832);
nand U4549 (N_4549,N_982,N_2261);
or U4550 (N_4550,N_1165,N_447);
xnor U4551 (N_4551,N_492,N_2314);
or U4552 (N_4552,N_126,N_530);
nor U4553 (N_4553,N_978,N_2125);
nor U4554 (N_4554,N_2236,N_2658);
and U4555 (N_4555,N_117,N_2280);
nand U4556 (N_4556,N_2013,N_1175);
xor U4557 (N_4557,N_475,N_2920);
or U4558 (N_4558,N_718,N_2055);
or U4559 (N_4559,N_2467,N_426);
nor U4560 (N_4560,N_2462,N_1232);
and U4561 (N_4561,N_915,N_1878);
or U4562 (N_4562,N_1637,N_985);
or U4563 (N_4563,N_1051,N_2723);
xor U4564 (N_4564,N_588,N_620);
nand U4565 (N_4565,N_883,N_1841);
xnor U4566 (N_4566,N_442,N_2103);
or U4567 (N_4567,N_2445,N_1648);
nor U4568 (N_4568,N_1725,N_512);
xor U4569 (N_4569,N_1639,N_2827);
xnor U4570 (N_4570,N_1977,N_2720);
or U4571 (N_4571,N_1652,N_1162);
and U4572 (N_4572,N_1432,N_2379);
or U4573 (N_4573,N_2590,N_614);
nor U4574 (N_4574,N_2206,N_1024);
and U4575 (N_4575,N_2010,N_799);
nand U4576 (N_4576,N_2932,N_2975);
nand U4577 (N_4577,N_837,N_914);
xor U4578 (N_4578,N_1528,N_2954);
nor U4579 (N_4579,N_273,N_1169);
nor U4580 (N_4580,N_1606,N_409);
nand U4581 (N_4581,N_2545,N_2825);
or U4582 (N_4582,N_223,N_2365);
nand U4583 (N_4583,N_1333,N_1300);
or U4584 (N_4584,N_1299,N_1120);
nand U4585 (N_4585,N_578,N_75);
nor U4586 (N_4586,N_761,N_297);
and U4587 (N_4587,N_51,N_238);
nand U4588 (N_4588,N_845,N_680);
nor U4589 (N_4589,N_834,N_278);
nor U4590 (N_4590,N_609,N_1767);
nor U4591 (N_4591,N_1694,N_2992);
or U4592 (N_4592,N_1896,N_2608);
nand U4593 (N_4593,N_1700,N_1528);
and U4594 (N_4594,N_275,N_251);
xor U4595 (N_4595,N_1716,N_2044);
nand U4596 (N_4596,N_1773,N_2729);
xnor U4597 (N_4597,N_1344,N_1098);
or U4598 (N_4598,N_1541,N_180);
and U4599 (N_4599,N_2186,N_1952);
nand U4600 (N_4600,N_1052,N_2385);
nor U4601 (N_4601,N_776,N_2585);
or U4602 (N_4602,N_2150,N_1673);
or U4603 (N_4603,N_1083,N_2602);
xor U4604 (N_4604,N_2642,N_1614);
nand U4605 (N_4605,N_2324,N_2230);
or U4606 (N_4606,N_2684,N_739);
and U4607 (N_4607,N_304,N_976);
nor U4608 (N_4608,N_2536,N_2651);
or U4609 (N_4609,N_563,N_38);
nand U4610 (N_4610,N_1071,N_1638);
or U4611 (N_4611,N_2928,N_91);
nor U4612 (N_4612,N_2870,N_1130);
xnor U4613 (N_4613,N_1745,N_2909);
nor U4614 (N_4614,N_2968,N_1268);
nor U4615 (N_4615,N_2794,N_2957);
and U4616 (N_4616,N_49,N_2985);
or U4617 (N_4617,N_729,N_1252);
nor U4618 (N_4618,N_2368,N_1732);
and U4619 (N_4619,N_595,N_880);
xnor U4620 (N_4620,N_1367,N_88);
nand U4621 (N_4621,N_2117,N_766);
or U4622 (N_4622,N_1006,N_2254);
nor U4623 (N_4623,N_1063,N_2776);
nand U4624 (N_4624,N_1464,N_2971);
nand U4625 (N_4625,N_656,N_2436);
nor U4626 (N_4626,N_681,N_23);
xor U4627 (N_4627,N_19,N_103);
and U4628 (N_4628,N_2016,N_38);
nor U4629 (N_4629,N_719,N_1720);
and U4630 (N_4630,N_1661,N_2755);
nand U4631 (N_4631,N_1990,N_308);
nor U4632 (N_4632,N_425,N_2201);
nand U4633 (N_4633,N_2712,N_389);
xnor U4634 (N_4634,N_2071,N_2481);
or U4635 (N_4635,N_2602,N_2229);
and U4636 (N_4636,N_2201,N_1287);
xor U4637 (N_4637,N_2836,N_67);
or U4638 (N_4638,N_2906,N_2441);
and U4639 (N_4639,N_648,N_951);
nand U4640 (N_4640,N_2285,N_917);
nor U4641 (N_4641,N_1080,N_1382);
nand U4642 (N_4642,N_1758,N_131);
nor U4643 (N_4643,N_2784,N_1714);
and U4644 (N_4644,N_1938,N_839);
xnor U4645 (N_4645,N_1043,N_667);
and U4646 (N_4646,N_2825,N_1286);
or U4647 (N_4647,N_1800,N_279);
nand U4648 (N_4648,N_2216,N_2084);
xnor U4649 (N_4649,N_968,N_2430);
nor U4650 (N_4650,N_395,N_1203);
or U4651 (N_4651,N_932,N_2843);
nand U4652 (N_4652,N_360,N_1987);
nand U4653 (N_4653,N_676,N_2478);
and U4654 (N_4654,N_1698,N_2764);
or U4655 (N_4655,N_2537,N_110);
nand U4656 (N_4656,N_1091,N_2376);
nor U4657 (N_4657,N_947,N_66);
or U4658 (N_4658,N_1186,N_1519);
and U4659 (N_4659,N_2602,N_1107);
xnor U4660 (N_4660,N_772,N_1943);
xnor U4661 (N_4661,N_175,N_2458);
xnor U4662 (N_4662,N_2503,N_723);
nand U4663 (N_4663,N_2691,N_1787);
or U4664 (N_4664,N_1052,N_2363);
nor U4665 (N_4665,N_2554,N_114);
nor U4666 (N_4666,N_1225,N_2991);
or U4667 (N_4667,N_2190,N_1907);
and U4668 (N_4668,N_351,N_2878);
nor U4669 (N_4669,N_1177,N_1917);
nand U4670 (N_4670,N_1625,N_321);
and U4671 (N_4671,N_2875,N_1186);
nor U4672 (N_4672,N_1284,N_1153);
xor U4673 (N_4673,N_1031,N_1409);
nor U4674 (N_4674,N_1306,N_2749);
and U4675 (N_4675,N_2891,N_1207);
or U4676 (N_4676,N_2709,N_1482);
or U4677 (N_4677,N_1304,N_1461);
and U4678 (N_4678,N_1478,N_1045);
xnor U4679 (N_4679,N_2255,N_1107);
nor U4680 (N_4680,N_473,N_2832);
nor U4681 (N_4681,N_2976,N_1876);
or U4682 (N_4682,N_1843,N_2047);
nand U4683 (N_4683,N_288,N_518);
or U4684 (N_4684,N_1889,N_1785);
nand U4685 (N_4685,N_1605,N_1537);
or U4686 (N_4686,N_529,N_1428);
and U4687 (N_4687,N_829,N_537);
and U4688 (N_4688,N_496,N_1918);
or U4689 (N_4689,N_2766,N_2670);
and U4690 (N_4690,N_2035,N_881);
or U4691 (N_4691,N_1787,N_2698);
or U4692 (N_4692,N_825,N_37);
nor U4693 (N_4693,N_83,N_69);
nand U4694 (N_4694,N_503,N_981);
xor U4695 (N_4695,N_1602,N_2392);
nor U4696 (N_4696,N_729,N_971);
nand U4697 (N_4697,N_1505,N_1459);
and U4698 (N_4698,N_2464,N_2757);
nand U4699 (N_4699,N_1039,N_2719);
nor U4700 (N_4700,N_2280,N_783);
nor U4701 (N_4701,N_236,N_674);
and U4702 (N_4702,N_1060,N_14);
or U4703 (N_4703,N_1515,N_105);
or U4704 (N_4704,N_346,N_1600);
nor U4705 (N_4705,N_418,N_134);
xor U4706 (N_4706,N_392,N_1120);
nand U4707 (N_4707,N_2687,N_384);
nor U4708 (N_4708,N_2925,N_673);
nand U4709 (N_4709,N_2203,N_462);
xor U4710 (N_4710,N_1275,N_314);
nand U4711 (N_4711,N_781,N_1026);
xor U4712 (N_4712,N_1491,N_2992);
and U4713 (N_4713,N_2097,N_1461);
nor U4714 (N_4714,N_629,N_70);
xnor U4715 (N_4715,N_2760,N_2224);
nand U4716 (N_4716,N_1387,N_993);
xnor U4717 (N_4717,N_220,N_696);
nor U4718 (N_4718,N_728,N_1803);
nand U4719 (N_4719,N_71,N_546);
xnor U4720 (N_4720,N_2853,N_811);
or U4721 (N_4721,N_2985,N_1875);
or U4722 (N_4722,N_1890,N_2396);
nand U4723 (N_4723,N_455,N_794);
or U4724 (N_4724,N_2874,N_661);
nand U4725 (N_4725,N_1161,N_870);
and U4726 (N_4726,N_1318,N_2938);
xnor U4727 (N_4727,N_2163,N_771);
and U4728 (N_4728,N_1126,N_1218);
nand U4729 (N_4729,N_679,N_1514);
xnor U4730 (N_4730,N_1016,N_140);
and U4731 (N_4731,N_936,N_126);
and U4732 (N_4732,N_1140,N_2898);
and U4733 (N_4733,N_2197,N_2471);
nor U4734 (N_4734,N_2255,N_1634);
and U4735 (N_4735,N_2077,N_59);
nor U4736 (N_4736,N_349,N_1190);
nor U4737 (N_4737,N_1571,N_1473);
nand U4738 (N_4738,N_2320,N_1693);
or U4739 (N_4739,N_1217,N_2927);
and U4740 (N_4740,N_1182,N_2296);
nor U4741 (N_4741,N_2999,N_553);
xor U4742 (N_4742,N_2762,N_2569);
nand U4743 (N_4743,N_1593,N_344);
and U4744 (N_4744,N_2400,N_785);
or U4745 (N_4745,N_1530,N_548);
and U4746 (N_4746,N_2479,N_1119);
or U4747 (N_4747,N_1221,N_210);
xnor U4748 (N_4748,N_2858,N_2797);
nor U4749 (N_4749,N_14,N_1496);
and U4750 (N_4750,N_862,N_1494);
xnor U4751 (N_4751,N_546,N_2539);
and U4752 (N_4752,N_2936,N_446);
and U4753 (N_4753,N_1951,N_2843);
nor U4754 (N_4754,N_1832,N_2235);
nor U4755 (N_4755,N_1657,N_764);
nor U4756 (N_4756,N_2086,N_2178);
nor U4757 (N_4757,N_2482,N_2988);
or U4758 (N_4758,N_388,N_361);
nor U4759 (N_4759,N_355,N_1970);
or U4760 (N_4760,N_2412,N_1077);
nand U4761 (N_4761,N_1711,N_1677);
xor U4762 (N_4762,N_2835,N_996);
and U4763 (N_4763,N_66,N_2703);
xor U4764 (N_4764,N_2394,N_2116);
or U4765 (N_4765,N_1731,N_848);
nand U4766 (N_4766,N_626,N_284);
nor U4767 (N_4767,N_68,N_2315);
or U4768 (N_4768,N_2080,N_2694);
and U4769 (N_4769,N_1125,N_988);
or U4770 (N_4770,N_2432,N_205);
nor U4771 (N_4771,N_1517,N_113);
and U4772 (N_4772,N_1086,N_50);
nor U4773 (N_4773,N_511,N_437);
nand U4774 (N_4774,N_487,N_1150);
and U4775 (N_4775,N_1693,N_264);
or U4776 (N_4776,N_803,N_603);
and U4777 (N_4777,N_1662,N_1568);
and U4778 (N_4778,N_306,N_445);
nor U4779 (N_4779,N_1310,N_1613);
and U4780 (N_4780,N_895,N_2340);
or U4781 (N_4781,N_1561,N_2192);
and U4782 (N_4782,N_90,N_2081);
nor U4783 (N_4783,N_2395,N_535);
and U4784 (N_4784,N_57,N_1771);
nor U4785 (N_4785,N_455,N_552);
nand U4786 (N_4786,N_2917,N_1550);
and U4787 (N_4787,N_1254,N_1403);
nand U4788 (N_4788,N_1620,N_150);
nand U4789 (N_4789,N_732,N_1132);
or U4790 (N_4790,N_2188,N_2215);
and U4791 (N_4791,N_1169,N_671);
nor U4792 (N_4792,N_1916,N_306);
xnor U4793 (N_4793,N_1861,N_56);
nor U4794 (N_4794,N_2924,N_1445);
nor U4795 (N_4795,N_716,N_1800);
and U4796 (N_4796,N_738,N_1320);
and U4797 (N_4797,N_1855,N_1411);
and U4798 (N_4798,N_2308,N_273);
and U4799 (N_4799,N_2024,N_23);
or U4800 (N_4800,N_501,N_552);
nor U4801 (N_4801,N_126,N_2651);
nand U4802 (N_4802,N_1741,N_2666);
nand U4803 (N_4803,N_1477,N_726);
and U4804 (N_4804,N_1037,N_1766);
or U4805 (N_4805,N_2445,N_470);
nor U4806 (N_4806,N_2507,N_2321);
and U4807 (N_4807,N_1202,N_2461);
nand U4808 (N_4808,N_259,N_1300);
nand U4809 (N_4809,N_2290,N_772);
nor U4810 (N_4810,N_2567,N_1037);
nand U4811 (N_4811,N_2670,N_2568);
nor U4812 (N_4812,N_2727,N_417);
and U4813 (N_4813,N_322,N_2758);
or U4814 (N_4814,N_1859,N_2644);
xor U4815 (N_4815,N_1015,N_1598);
nor U4816 (N_4816,N_701,N_1533);
xor U4817 (N_4817,N_520,N_2336);
and U4818 (N_4818,N_2015,N_570);
or U4819 (N_4819,N_500,N_1919);
and U4820 (N_4820,N_1899,N_1134);
or U4821 (N_4821,N_564,N_2125);
nor U4822 (N_4822,N_1984,N_500);
nor U4823 (N_4823,N_2290,N_547);
and U4824 (N_4824,N_642,N_1933);
nor U4825 (N_4825,N_2242,N_2888);
nand U4826 (N_4826,N_2440,N_2408);
or U4827 (N_4827,N_1926,N_2418);
xor U4828 (N_4828,N_2722,N_1519);
nor U4829 (N_4829,N_717,N_1002);
nor U4830 (N_4830,N_1139,N_2112);
nand U4831 (N_4831,N_2878,N_846);
and U4832 (N_4832,N_228,N_1521);
and U4833 (N_4833,N_1592,N_451);
or U4834 (N_4834,N_1724,N_1753);
nor U4835 (N_4835,N_2887,N_2582);
and U4836 (N_4836,N_981,N_901);
xor U4837 (N_4837,N_1504,N_2732);
nor U4838 (N_4838,N_541,N_2815);
xnor U4839 (N_4839,N_1749,N_595);
or U4840 (N_4840,N_1491,N_1486);
and U4841 (N_4841,N_2451,N_673);
nand U4842 (N_4842,N_1873,N_1204);
nor U4843 (N_4843,N_1577,N_1310);
nor U4844 (N_4844,N_1620,N_2228);
nand U4845 (N_4845,N_585,N_2472);
nor U4846 (N_4846,N_2737,N_2726);
xor U4847 (N_4847,N_1462,N_2145);
xnor U4848 (N_4848,N_2286,N_1610);
nand U4849 (N_4849,N_1528,N_1032);
or U4850 (N_4850,N_2328,N_2373);
nor U4851 (N_4851,N_2286,N_1444);
nor U4852 (N_4852,N_2291,N_578);
xor U4853 (N_4853,N_1452,N_2730);
and U4854 (N_4854,N_2377,N_60);
or U4855 (N_4855,N_1298,N_371);
or U4856 (N_4856,N_256,N_2351);
nand U4857 (N_4857,N_805,N_177);
and U4858 (N_4858,N_1272,N_307);
nor U4859 (N_4859,N_2452,N_702);
nor U4860 (N_4860,N_240,N_1996);
or U4861 (N_4861,N_2797,N_449);
or U4862 (N_4862,N_1134,N_2483);
or U4863 (N_4863,N_1437,N_2669);
or U4864 (N_4864,N_809,N_2125);
xor U4865 (N_4865,N_871,N_2086);
xor U4866 (N_4866,N_810,N_277);
xnor U4867 (N_4867,N_2619,N_937);
xnor U4868 (N_4868,N_1856,N_1123);
xor U4869 (N_4869,N_2372,N_2261);
and U4870 (N_4870,N_1045,N_414);
nand U4871 (N_4871,N_476,N_1471);
nor U4872 (N_4872,N_265,N_275);
nor U4873 (N_4873,N_52,N_897);
nor U4874 (N_4874,N_2558,N_1317);
nor U4875 (N_4875,N_1038,N_2002);
xnor U4876 (N_4876,N_2638,N_2348);
or U4877 (N_4877,N_1973,N_2788);
nand U4878 (N_4878,N_839,N_1305);
and U4879 (N_4879,N_1942,N_670);
or U4880 (N_4880,N_2122,N_1573);
and U4881 (N_4881,N_637,N_1549);
or U4882 (N_4882,N_2335,N_1855);
xor U4883 (N_4883,N_2615,N_1702);
xor U4884 (N_4884,N_1721,N_1805);
nor U4885 (N_4885,N_280,N_1477);
nor U4886 (N_4886,N_544,N_701);
nor U4887 (N_4887,N_2504,N_681);
xor U4888 (N_4888,N_1670,N_1144);
nand U4889 (N_4889,N_509,N_1522);
nor U4890 (N_4890,N_1655,N_2536);
and U4891 (N_4891,N_1828,N_307);
nor U4892 (N_4892,N_412,N_1058);
xor U4893 (N_4893,N_1080,N_2750);
nand U4894 (N_4894,N_658,N_232);
and U4895 (N_4895,N_2348,N_1575);
and U4896 (N_4896,N_1593,N_1501);
xor U4897 (N_4897,N_1185,N_2378);
xor U4898 (N_4898,N_837,N_1203);
xor U4899 (N_4899,N_69,N_1368);
or U4900 (N_4900,N_368,N_2971);
xnor U4901 (N_4901,N_378,N_2493);
nor U4902 (N_4902,N_2745,N_2218);
or U4903 (N_4903,N_330,N_614);
or U4904 (N_4904,N_1888,N_2763);
or U4905 (N_4905,N_2218,N_1897);
nand U4906 (N_4906,N_629,N_2088);
nor U4907 (N_4907,N_438,N_2733);
or U4908 (N_4908,N_1895,N_297);
nand U4909 (N_4909,N_1976,N_2362);
nor U4910 (N_4910,N_1364,N_1293);
nor U4911 (N_4911,N_2183,N_643);
xnor U4912 (N_4912,N_359,N_531);
xor U4913 (N_4913,N_1395,N_2817);
nor U4914 (N_4914,N_1443,N_2348);
nand U4915 (N_4915,N_1067,N_1328);
and U4916 (N_4916,N_1465,N_1470);
or U4917 (N_4917,N_1535,N_822);
or U4918 (N_4918,N_2352,N_2711);
or U4919 (N_4919,N_1460,N_340);
and U4920 (N_4920,N_2143,N_1405);
nor U4921 (N_4921,N_2292,N_1174);
and U4922 (N_4922,N_1695,N_2826);
nor U4923 (N_4923,N_463,N_1023);
and U4924 (N_4924,N_2970,N_153);
nor U4925 (N_4925,N_1413,N_961);
xor U4926 (N_4926,N_1598,N_825);
and U4927 (N_4927,N_1483,N_1538);
xor U4928 (N_4928,N_2844,N_2008);
nor U4929 (N_4929,N_1762,N_453);
and U4930 (N_4930,N_2928,N_2365);
nor U4931 (N_4931,N_256,N_2974);
and U4932 (N_4932,N_1269,N_2038);
nand U4933 (N_4933,N_2136,N_1575);
xor U4934 (N_4934,N_763,N_1555);
and U4935 (N_4935,N_2714,N_2913);
nor U4936 (N_4936,N_1905,N_1231);
or U4937 (N_4937,N_2206,N_152);
xor U4938 (N_4938,N_2851,N_502);
nand U4939 (N_4939,N_2292,N_162);
or U4940 (N_4940,N_1222,N_128);
and U4941 (N_4941,N_2806,N_2350);
nor U4942 (N_4942,N_2065,N_84);
nor U4943 (N_4943,N_735,N_2295);
or U4944 (N_4944,N_2259,N_2520);
nand U4945 (N_4945,N_73,N_2782);
xnor U4946 (N_4946,N_788,N_1231);
nand U4947 (N_4947,N_247,N_573);
xnor U4948 (N_4948,N_1282,N_2161);
or U4949 (N_4949,N_1580,N_2275);
nand U4950 (N_4950,N_2582,N_2525);
or U4951 (N_4951,N_587,N_2079);
xor U4952 (N_4952,N_1431,N_833);
nand U4953 (N_4953,N_2494,N_2110);
or U4954 (N_4954,N_573,N_963);
xnor U4955 (N_4955,N_2790,N_949);
nor U4956 (N_4956,N_2172,N_84);
nand U4957 (N_4957,N_1301,N_313);
nand U4958 (N_4958,N_942,N_2501);
nor U4959 (N_4959,N_2852,N_730);
or U4960 (N_4960,N_692,N_2112);
nand U4961 (N_4961,N_1254,N_59);
and U4962 (N_4962,N_1871,N_1181);
nand U4963 (N_4963,N_2515,N_2779);
or U4964 (N_4964,N_1720,N_2712);
nand U4965 (N_4965,N_2120,N_250);
nand U4966 (N_4966,N_474,N_2728);
xnor U4967 (N_4967,N_2245,N_115);
xor U4968 (N_4968,N_2075,N_1758);
and U4969 (N_4969,N_2648,N_2889);
nor U4970 (N_4970,N_690,N_2329);
and U4971 (N_4971,N_124,N_61);
or U4972 (N_4972,N_2397,N_702);
nand U4973 (N_4973,N_1818,N_2180);
nor U4974 (N_4974,N_2917,N_2795);
or U4975 (N_4975,N_2793,N_1187);
nand U4976 (N_4976,N_735,N_399);
and U4977 (N_4977,N_2379,N_880);
nor U4978 (N_4978,N_783,N_1324);
nor U4979 (N_4979,N_848,N_928);
xor U4980 (N_4980,N_1169,N_1834);
nor U4981 (N_4981,N_1059,N_1441);
nor U4982 (N_4982,N_2228,N_1814);
nor U4983 (N_4983,N_2576,N_606);
and U4984 (N_4984,N_326,N_1885);
nor U4985 (N_4985,N_2187,N_1351);
and U4986 (N_4986,N_2717,N_1051);
and U4987 (N_4987,N_216,N_2674);
nand U4988 (N_4988,N_1660,N_954);
xnor U4989 (N_4989,N_1130,N_2460);
xnor U4990 (N_4990,N_1726,N_1999);
xor U4991 (N_4991,N_1570,N_390);
nor U4992 (N_4992,N_2519,N_962);
or U4993 (N_4993,N_2413,N_992);
nand U4994 (N_4994,N_504,N_774);
xor U4995 (N_4995,N_2119,N_2656);
and U4996 (N_4996,N_2522,N_480);
nand U4997 (N_4997,N_1281,N_217);
nor U4998 (N_4998,N_218,N_2723);
and U4999 (N_4999,N_2112,N_1766);
xor U5000 (N_5000,N_2950,N_1999);
xor U5001 (N_5001,N_1185,N_2362);
xnor U5002 (N_5002,N_1414,N_2857);
and U5003 (N_5003,N_2792,N_313);
or U5004 (N_5004,N_2629,N_2049);
and U5005 (N_5005,N_1362,N_1991);
and U5006 (N_5006,N_79,N_953);
nor U5007 (N_5007,N_1671,N_1280);
xnor U5008 (N_5008,N_878,N_558);
nor U5009 (N_5009,N_2883,N_2153);
or U5010 (N_5010,N_1521,N_2236);
xnor U5011 (N_5011,N_434,N_1715);
or U5012 (N_5012,N_896,N_2683);
or U5013 (N_5013,N_826,N_337);
or U5014 (N_5014,N_1731,N_2355);
xor U5015 (N_5015,N_1641,N_1080);
or U5016 (N_5016,N_1427,N_2861);
or U5017 (N_5017,N_1556,N_347);
xnor U5018 (N_5018,N_2614,N_704);
nand U5019 (N_5019,N_2,N_2705);
nor U5020 (N_5020,N_1337,N_779);
nand U5021 (N_5021,N_201,N_1740);
and U5022 (N_5022,N_856,N_2982);
nand U5023 (N_5023,N_2153,N_2925);
nand U5024 (N_5024,N_1320,N_2129);
xnor U5025 (N_5025,N_982,N_1366);
nand U5026 (N_5026,N_2655,N_2099);
nor U5027 (N_5027,N_2686,N_639);
nor U5028 (N_5028,N_194,N_2920);
or U5029 (N_5029,N_723,N_1775);
xnor U5030 (N_5030,N_1192,N_1617);
nor U5031 (N_5031,N_195,N_1567);
xnor U5032 (N_5032,N_2059,N_1119);
and U5033 (N_5033,N_87,N_2800);
or U5034 (N_5034,N_1307,N_2881);
or U5035 (N_5035,N_303,N_289);
xnor U5036 (N_5036,N_2795,N_2906);
xnor U5037 (N_5037,N_2639,N_1729);
and U5038 (N_5038,N_2513,N_1416);
and U5039 (N_5039,N_368,N_1454);
nor U5040 (N_5040,N_483,N_186);
nor U5041 (N_5041,N_1498,N_807);
or U5042 (N_5042,N_1373,N_826);
or U5043 (N_5043,N_1821,N_79);
xnor U5044 (N_5044,N_2531,N_2450);
xor U5045 (N_5045,N_1082,N_1875);
nand U5046 (N_5046,N_834,N_2964);
or U5047 (N_5047,N_1783,N_10);
nor U5048 (N_5048,N_1,N_887);
nand U5049 (N_5049,N_127,N_418);
or U5050 (N_5050,N_1417,N_470);
nand U5051 (N_5051,N_221,N_1127);
nor U5052 (N_5052,N_127,N_1060);
nor U5053 (N_5053,N_1939,N_1728);
or U5054 (N_5054,N_300,N_2844);
nand U5055 (N_5055,N_2441,N_1834);
or U5056 (N_5056,N_1229,N_1333);
nor U5057 (N_5057,N_837,N_808);
xor U5058 (N_5058,N_2353,N_2461);
xor U5059 (N_5059,N_218,N_2846);
and U5060 (N_5060,N_2683,N_452);
and U5061 (N_5061,N_320,N_1291);
or U5062 (N_5062,N_1560,N_551);
nor U5063 (N_5063,N_1639,N_395);
or U5064 (N_5064,N_2944,N_2281);
nand U5065 (N_5065,N_468,N_513);
nor U5066 (N_5066,N_1634,N_2595);
nand U5067 (N_5067,N_983,N_391);
and U5068 (N_5068,N_424,N_1878);
xor U5069 (N_5069,N_1451,N_175);
xor U5070 (N_5070,N_2513,N_1977);
xor U5071 (N_5071,N_316,N_2190);
xnor U5072 (N_5072,N_2956,N_945);
and U5073 (N_5073,N_2338,N_1005);
or U5074 (N_5074,N_2705,N_2837);
nor U5075 (N_5075,N_2427,N_2022);
nor U5076 (N_5076,N_1008,N_803);
xnor U5077 (N_5077,N_597,N_954);
nand U5078 (N_5078,N_1582,N_1366);
nand U5079 (N_5079,N_197,N_879);
nand U5080 (N_5080,N_1233,N_1438);
and U5081 (N_5081,N_2449,N_2155);
and U5082 (N_5082,N_2246,N_1764);
nor U5083 (N_5083,N_2457,N_1362);
nor U5084 (N_5084,N_1764,N_664);
nand U5085 (N_5085,N_2367,N_1837);
and U5086 (N_5086,N_2700,N_1164);
nor U5087 (N_5087,N_1611,N_1277);
nor U5088 (N_5088,N_157,N_2550);
nor U5089 (N_5089,N_1059,N_121);
xnor U5090 (N_5090,N_2100,N_1621);
nor U5091 (N_5091,N_1972,N_2450);
and U5092 (N_5092,N_262,N_1733);
xor U5093 (N_5093,N_1120,N_1696);
nor U5094 (N_5094,N_1583,N_242);
or U5095 (N_5095,N_2551,N_678);
and U5096 (N_5096,N_86,N_282);
and U5097 (N_5097,N_2555,N_1277);
xor U5098 (N_5098,N_18,N_182);
nor U5099 (N_5099,N_2679,N_2597);
nand U5100 (N_5100,N_1123,N_2235);
or U5101 (N_5101,N_2350,N_990);
or U5102 (N_5102,N_2057,N_2917);
nand U5103 (N_5103,N_1456,N_2978);
xor U5104 (N_5104,N_418,N_1275);
or U5105 (N_5105,N_1697,N_1056);
nor U5106 (N_5106,N_966,N_35);
xnor U5107 (N_5107,N_1136,N_2012);
xnor U5108 (N_5108,N_2934,N_1795);
nand U5109 (N_5109,N_1591,N_1975);
nor U5110 (N_5110,N_368,N_52);
and U5111 (N_5111,N_427,N_1166);
nand U5112 (N_5112,N_51,N_2119);
and U5113 (N_5113,N_930,N_250);
nand U5114 (N_5114,N_2388,N_2507);
and U5115 (N_5115,N_1261,N_810);
and U5116 (N_5116,N_1710,N_2332);
nor U5117 (N_5117,N_2911,N_699);
xor U5118 (N_5118,N_580,N_2703);
and U5119 (N_5119,N_1107,N_1582);
nor U5120 (N_5120,N_2561,N_854);
and U5121 (N_5121,N_532,N_2030);
xor U5122 (N_5122,N_2153,N_2970);
or U5123 (N_5123,N_2537,N_265);
nor U5124 (N_5124,N_1119,N_2687);
and U5125 (N_5125,N_235,N_1936);
or U5126 (N_5126,N_67,N_2906);
nor U5127 (N_5127,N_2327,N_2449);
or U5128 (N_5128,N_1480,N_1237);
and U5129 (N_5129,N_1306,N_1620);
and U5130 (N_5130,N_2249,N_2476);
nor U5131 (N_5131,N_452,N_2797);
or U5132 (N_5132,N_2015,N_1433);
nand U5133 (N_5133,N_2932,N_1511);
nor U5134 (N_5134,N_1351,N_581);
and U5135 (N_5135,N_914,N_2966);
and U5136 (N_5136,N_1777,N_1297);
and U5137 (N_5137,N_2446,N_421);
xor U5138 (N_5138,N_254,N_2431);
nor U5139 (N_5139,N_2410,N_533);
nand U5140 (N_5140,N_466,N_2022);
xor U5141 (N_5141,N_488,N_1282);
and U5142 (N_5142,N_2968,N_1627);
and U5143 (N_5143,N_933,N_2889);
nor U5144 (N_5144,N_1448,N_2697);
and U5145 (N_5145,N_325,N_1018);
or U5146 (N_5146,N_1442,N_2187);
nand U5147 (N_5147,N_2787,N_1607);
nor U5148 (N_5148,N_2218,N_1300);
and U5149 (N_5149,N_998,N_1082);
nor U5150 (N_5150,N_610,N_1977);
nor U5151 (N_5151,N_585,N_962);
xor U5152 (N_5152,N_164,N_2890);
nand U5153 (N_5153,N_2438,N_1409);
and U5154 (N_5154,N_2366,N_1051);
or U5155 (N_5155,N_2983,N_2922);
or U5156 (N_5156,N_2024,N_786);
nand U5157 (N_5157,N_67,N_931);
nor U5158 (N_5158,N_570,N_2505);
and U5159 (N_5159,N_2373,N_1193);
nand U5160 (N_5160,N_1264,N_369);
and U5161 (N_5161,N_1599,N_870);
nand U5162 (N_5162,N_1939,N_1271);
nor U5163 (N_5163,N_2450,N_2729);
nand U5164 (N_5164,N_2750,N_2293);
nor U5165 (N_5165,N_494,N_933);
nor U5166 (N_5166,N_107,N_2672);
and U5167 (N_5167,N_1074,N_705);
nand U5168 (N_5168,N_1531,N_1027);
nand U5169 (N_5169,N_397,N_1720);
and U5170 (N_5170,N_1169,N_1421);
and U5171 (N_5171,N_488,N_2090);
xor U5172 (N_5172,N_585,N_1525);
nor U5173 (N_5173,N_1002,N_248);
nand U5174 (N_5174,N_123,N_2261);
nand U5175 (N_5175,N_180,N_521);
and U5176 (N_5176,N_668,N_1342);
nand U5177 (N_5177,N_2994,N_660);
nand U5178 (N_5178,N_988,N_2905);
nand U5179 (N_5179,N_1457,N_1022);
or U5180 (N_5180,N_44,N_1442);
and U5181 (N_5181,N_2459,N_95);
or U5182 (N_5182,N_2279,N_2295);
and U5183 (N_5183,N_2303,N_570);
or U5184 (N_5184,N_1891,N_475);
xor U5185 (N_5185,N_852,N_254);
and U5186 (N_5186,N_571,N_1559);
and U5187 (N_5187,N_633,N_1823);
and U5188 (N_5188,N_1944,N_2868);
xor U5189 (N_5189,N_2523,N_1939);
xnor U5190 (N_5190,N_1085,N_2607);
nor U5191 (N_5191,N_2287,N_164);
and U5192 (N_5192,N_989,N_1175);
nand U5193 (N_5193,N_724,N_1740);
or U5194 (N_5194,N_1370,N_2949);
nand U5195 (N_5195,N_658,N_1607);
nand U5196 (N_5196,N_1483,N_1110);
xor U5197 (N_5197,N_2367,N_2024);
nand U5198 (N_5198,N_1911,N_1076);
nor U5199 (N_5199,N_199,N_967);
or U5200 (N_5200,N_585,N_2954);
nor U5201 (N_5201,N_1723,N_2252);
nor U5202 (N_5202,N_648,N_115);
xor U5203 (N_5203,N_2199,N_654);
or U5204 (N_5204,N_984,N_1404);
or U5205 (N_5205,N_1963,N_2906);
xor U5206 (N_5206,N_368,N_74);
and U5207 (N_5207,N_444,N_2832);
and U5208 (N_5208,N_415,N_2524);
nor U5209 (N_5209,N_1739,N_807);
nor U5210 (N_5210,N_1760,N_1841);
or U5211 (N_5211,N_845,N_889);
nand U5212 (N_5212,N_961,N_919);
and U5213 (N_5213,N_1677,N_1379);
and U5214 (N_5214,N_687,N_50);
or U5215 (N_5215,N_2629,N_763);
nand U5216 (N_5216,N_1004,N_1843);
xor U5217 (N_5217,N_1020,N_2822);
nand U5218 (N_5218,N_161,N_1634);
nand U5219 (N_5219,N_1231,N_652);
xor U5220 (N_5220,N_2322,N_1372);
and U5221 (N_5221,N_2912,N_975);
nor U5222 (N_5222,N_2911,N_999);
nand U5223 (N_5223,N_1492,N_2149);
nand U5224 (N_5224,N_129,N_1100);
and U5225 (N_5225,N_823,N_1704);
or U5226 (N_5226,N_2867,N_1627);
or U5227 (N_5227,N_1496,N_343);
nor U5228 (N_5228,N_922,N_1555);
xor U5229 (N_5229,N_817,N_1766);
or U5230 (N_5230,N_621,N_2902);
xnor U5231 (N_5231,N_2768,N_689);
xor U5232 (N_5232,N_1842,N_798);
and U5233 (N_5233,N_461,N_278);
or U5234 (N_5234,N_2413,N_396);
nand U5235 (N_5235,N_940,N_2935);
nand U5236 (N_5236,N_978,N_2665);
and U5237 (N_5237,N_1838,N_2983);
or U5238 (N_5238,N_758,N_1063);
or U5239 (N_5239,N_958,N_728);
nand U5240 (N_5240,N_526,N_2705);
xor U5241 (N_5241,N_1609,N_1760);
nor U5242 (N_5242,N_1708,N_1297);
and U5243 (N_5243,N_1284,N_232);
or U5244 (N_5244,N_1955,N_2442);
and U5245 (N_5245,N_904,N_279);
or U5246 (N_5246,N_1711,N_407);
and U5247 (N_5247,N_1413,N_1534);
nand U5248 (N_5248,N_2906,N_1199);
or U5249 (N_5249,N_2738,N_2572);
and U5250 (N_5250,N_207,N_2436);
xnor U5251 (N_5251,N_1079,N_2273);
nand U5252 (N_5252,N_162,N_2276);
and U5253 (N_5253,N_2091,N_391);
xor U5254 (N_5254,N_554,N_1080);
or U5255 (N_5255,N_2842,N_636);
nor U5256 (N_5256,N_139,N_1);
nor U5257 (N_5257,N_483,N_2054);
nand U5258 (N_5258,N_917,N_1718);
nor U5259 (N_5259,N_1087,N_1004);
and U5260 (N_5260,N_1208,N_688);
or U5261 (N_5261,N_831,N_1170);
nor U5262 (N_5262,N_2006,N_2129);
or U5263 (N_5263,N_1370,N_1467);
or U5264 (N_5264,N_855,N_2330);
nand U5265 (N_5265,N_1833,N_2975);
nor U5266 (N_5266,N_1416,N_1000);
nand U5267 (N_5267,N_990,N_2501);
nor U5268 (N_5268,N_53,N_2764);
nand U5269 (N_5269,N_1289,N_819);
nor U5270 (N_5270,N_498,N_506);
nor U5271 (N_5271,N_953,N_739);
and U5272 (N_5272,N_2423,N_165);
or U5273 (N_5273,N_1309,N_1400);
nand U5274 (N_5274,N_3,N_1142);
xor U5275 (N_5275,N_2156,N_893);
nor U5276 (N_5276,N_1931,N_2016);
and U5277 (N_5277,N_612,N_1708);
or U5278 (N_5278,N_2942,N_449);
nand U5279 (N_5279,N_918,N_291);
nor U5280 (N_5280,N_2630,N_24);
or U5281 (N_5281,N_491,N_2699);
xnor U5282 (N_5282,N_2043,N_467);
xnor U5283 (N_5283,N_190,N_1653);
xnor U5284 (N_5284,N_1386,N_2507);
nor U5285 (N_5285,N_2019,N_2666);
or U5286 (N_5286,N_589,N_2231);
xor U5287 (N_5287,N_2817,N_2139);
nor U5288 (N_5288,N_2869,N_302);
or U5289 (N_5289,N_554,N_2113);
and U5290 (N_5290,N_508,N_810);
nand U5291 (N_5291,N_1469,N_1103);
and U5292 (N_5292,N_1984,N_2133);
and U5293 (N_5293,N_2345,N_69);
and U5294 (N_5294,N_1823,N_594);
xnor U5295 (N_5295,N_986,N_2572);
xor U5296 (N_5296,N_1455,N_2868);
and U5297 (N_5297,N_853,N_1197);
xor U5298 (N_5298,N_2818,N_2817);
or U5299 (N_5299,N_1693,N_2440);
and U5300 (N_5300,N_1399,N_2491);
nor U5301 (N_5301,N_715,N_1250);
nor U5302 (N_5302,N_1596,N_1269);
xnor U5303 (N_5303,N_464,N_668);
and U5304 (N_5304,N_946,N_1268);
xnor U5305 (N_5305,N_1626,N_2092);
nand U5306 (N_5306,N_2839,N_2538);
xnor U5307 (N_5307,N_962,N_2540);
xnor U5308 (N_5308,N_1780,N_2960);
nor U5309 (N_5309,N_730,N_573);
nand U5310 (N_5310,N_1338,N_2809);
nor U5311 (N_5311,N_333,N_1610);
or U5312 (N_5312,N_2950,N_1110);
nand U5313 (N_5313,N_707,N_2272);
xor U5314 (N_5314,N_2592,N_1023);
xor U5315 (N_5315,N_2263,N_418);
nor U5316 (N_5316,N_370,N_1462);
xnor U5317 (N_5317,N_1484,N_2303);
nor U5318 (N_5318,N_1585,N_2331);
nor U5319 (N_5319,N_2995,N_1605);
nand U5320 (N_5320,N_2246,N_648);
nand U5321 (N_5321,N_1445,N_2719);
nand U5322 (N_5322,N_1250,N_671);
nand U5323 (N_5323,N_1209,N_2211);
and U5324 (N_5324,N_2026,N_1323);
xor U5325 (N_5325,N_882,N_2257);
nor U5326 (N_5326,N_540,N_2948);
and U5327 (N_5327,N_370,N_2675);
nand U5328 (N_5328,N_1217,N_1403);
xor U5329 (N_5329,N_230,N_2346);
or U5330 (N_5330,N_462,N_1169);
and U5331 (N_5331,N_2893,N_69);
nor U5332 (N_5332,N_1060,N_847);
nor U5333 (N_5333,N_2422,N_1766);
nand U5334 (N_5334,N_213,N_230);
nor U5335 (N_5335,N_1141,N_1655);
and U5336 (N_5336,N_2918,N_2048);
and U5337 (N_5337,N_296,N_1259);
nor U5338 (N_5338,N_1087,N_2420);
or U5339 (N_5339,N_585,N_1966);
xnor U5340 (N_5340,N_2776,N_1852);
and U5341 (N_5341,N_1084,N_1600);
nand U5342 (N_5342,N_707,N_362);
xnor U5343 (N_5343,N_1676,N_1492);
nand U5344 (N_5344,N_1921,N_922);
nor U5345 (N_5345,N_352,N_1360);
or U5346 (N_5346,N_2506,N_557);
xnor U5347 (N_5347,N_752,N_1090);
nand U5348 (N_5348,N_298,N_1943);
nor U5349 (N_5349,N_1444,N_1818);
nor U5350 (N_5350,N_2602,N_2580);
nand U5351 (N_5351,N_1078,N_1992);
and U5352 (N_5352,N_1512,N_37);
or U5353 (N_5353,N_1296,N_1281);
nand U5354 (N_5354,N_1917,N_259);
nand U5355 (N_5355,N_2341,N_2363);
xor U5356 (N_5356,N_1159,N_399);
xor U5357 (N_5357,N_2662,N_273);
nor U5358 (N_5358,N_1505,N_1282);
xnor U5359 (N_5359,N_2679,N_1824);
nand U5360 (N_5360,N_2340,N_1005);
or U5361 (N_5361,N_1218,N_1195);
nor U5362 (N_5362,N_2585,N_1048);
nand U5363 (N_5363,N_1996,N_1774);
or U5364 (N_5364,N_2558,N_233);
nor U5365 (N_5365,N_2558,N_307);
nand U5366 (N_5366,N_2163,N_1829);
or U5367 (N_5367,N_630,N_42);
nand U5368 (N_5368,N_435,N_987);
and U5369 (N_5369,N_2186,N_1313);
nor U5370 (N_5370,N_633,N_2585);
and U5371 (N_5371,N_2245,N_901);
or U5372 (N_5372,N_1789,N_826);
nor U5373 (N_5373,N_1282,N_1483);
nor U5374 (N_5374,N_1534,N_2922);
and U5375 (N_5375,N_1900,N_2961);
nor U5376 (N_5376,N_1872,N_2330);
or U5377 (N_5377,N_2223,N_117);
nand U5378 (N_5378,N_1961,N_1130);
or U5379 (N_5379,N_64,N_566);
xor U5380 (N_5380,N_594,N_2748);
nor U5381 (N_5381,N_558,N_2924);
or U5382 (N_5382,N_1388,N_957);
xor U5383 (N_5383,N_2175,N_2519);
nand U5384 (N_5384,N_2165,N_1222);
or U5385 (N_5385,N_143,N_2382);
nor U5386 (N_5386,N_744,N_252);
nor U5387 (N_5387,N_788,N_2957);
nand U5388 (N_5388,N_1994,N_2018);
or U5389 (N_5389,N_1535,N_40);
and U5390 (N_5390,N_425,N_812);
xnor U5391 (N_5391,N_482,N_566);
or U5392 (N_5392,N_2474,N_679);
nand U5393 (N_5393,N_2057,N_1868);
nand U5394 (N_5394,N_2761,N_2835);
or U5395 (N_5395,N_388,N_946);
or U5396 (N_5396,N_2204,N_2529);
and U5397 (N_5397,N_2255,N_2477);
or U5398 (N_5398,N_1356,N_2527);
nor U5399 (N_5399,N_1,N_235);
nand U5400 (N_5400,N_2489,N_1212);
or U5401 (N_5401,N_1639,N_1745);
or U5402 (N_5402,N_2074,N_1516);
nor U5403 (N_5403,N_8,N_1250);
nor U5404 (N_5404,N_1811,N_2118);
xor U5405 (N_5405,N_901,N_2709);
xnor U5406 (N_5406,N_1216,N_1739);
and U5407 (N_5407,N_1618,N_1925);
nand U5408 (N_5408,N_813,N_1527);
or U5409 (N_5409,N_2654,N_1418);
and U5410 (N_5410,N_279,N_1817);
nor U5411 (N_5411,N_2310,N_2734);
nor U5412 (N_5412,N_2535,N_2668);
and U5413 (N_5413,N_1666,N_482);
or U5414 (N_5414,N_686,N_1746);
or U5415 (N_5415,N_2963,N_2266);
and U5416 (N_5416,N_104,N_1113);
nand U5417 (N_5417,N_1096,N_1362);
or U5418 (N_5418,N_335,N_2519);
nand U5419 (N_5419,N_362,N_412);
xor U5420 (N_5420,N_935,N_272);
nor U5421 (N_5421,N_2184,N_29);
nor U5422 (N_5422,N_1325,N_2998);
nand U5423 (N_5423,N_770,N_539);
xnor U5424 (N_5424,N_1768,N_1719);
xnor U5425 (N_5425,N_1806,N_2346);
xnor U5426 (N_5426,N_1729,N_1091);
and U5427 (N_5427,N_292,N_476);
xnor U5428 (N_5428,N_1186,N_1744);
nand U5429 (N_5429,N_2641,N_1670);
or U5430 (N_5430,N_703,N_888);
nand U5431 (N_5431,N_1228,N_2426);
nand U5432 (N_5432,N_557,N_2933);
and U5433 (N_5433,N_2786,N_244);
xnor U5434 (N_5434,N_1054,N_2625);
and U5435 (N_5435,N_2804,N_664);
xor U5436 (N_5436,N_1274,N_1629);
nand U5437 (N_5437,N_404,N_1670);
xor U5438 (N_5438,N_2589,N_676);
and U5439 (N_5439,N_1394,N_1057);
nand U5440 (N_5440,N_1917,N_615);
or U5441 (N_5441,N_1367,N_1071);
xor U5442 (N_5442,N_1236,N_2507);
xor U5443 (N_5443,N_1923,N_2753);
nand U5444 (N_5444,N_2474,N_548);
nand U5445 (N_5445,N_1819,N_2786);
xor U5446 (N_5446,N_1721,N_640);
or U5447 (N_5447,N_965,N_2408);
nor U5448 (N_5448,N_1171,N_1525);
and U5449 (N_5449,N_623,N_1283);
and U5450 (N_5450,N_2569,N_2731);
nand U5451 (N_5451,N_829,N_1031);
nor U5452 (N_5452,N_2906,N_1562);
nand U5453 (N_5453,N_2596,N_582);
nor U5454 (N_5454,N_332,N_89);
nand U5455 (N_5455,N_2345,N_24);
nand U5456 (N_5456,N_898,N_1458);
xnor U5457 (N_5457,N_186,N_404);
xor U5458 (N_5458,N_1455,N_1296);
or U5459 (N_5459,N_1331,N_1646);
nand U5460 (N_5460,N_2819,N_2279);
or U5461 (N_5461,N_1318,N_1408);
or U5462 (N_5462,N_936,N_949);
nor U5463 (N_5463,N_2139,N_928);
nor U5464 (N_5464,N_148,N_158);
nand U5465 (N_5465,N_429,N_1958);
nor U5466 (N_5466,N_1207,N_2092);
or U5467 (N_5467,N_2416,N_1976);
xnor U5468 (N_5468,N_415,N_622);
nand U5469 (N_5469,N_2407,N_2133);
xnor U5470 (N_5470,N_391,N_340);
nor U5471 (N_5471,N_2699,N_2338);
and U5472 (N_5472,N_1562,N_2451);
nand U5473 (N_5473,N_743,N_268);
and U5474 (N_5474,N_1382,N_645);
xor U5475 (N_5475,N_383,N_117);
or U5476 (N_5476,N_1174,N_678);
nand U5477 (N_5477,N_1289,N_1824);
nand U5478 (N_5478,N_2828,N_1373);
xor U5479 (N_5479,N_2217,N_1471);
nor U5480 (N_5480,N_1731,N_531);
or U5481 (N_5481,N_2182,N_1387);
nand U5482 (N_5482,N_1972,N_2766);
and U5483 (N_5483,N_868,N_2518);
or U5484 (N_5484,N_1139,N_543);
or U5485 (N_5485,N_1355,N_492);
or U5486 (N_5486,N_2365,N_2755);
and U5487 (N_5487,N_2531,N_1942);
and U5488 (N_5488,N_2453,N_966);
nand U5489 (N_5489,N_42,N_76);
nand U5490 (N_5490,N_137,N_1997);
or U5491 (N_5491,N_1443,N_732);
or U5492 (N_5492,N_217,N_290);
or U5493 (N_5493,N_2607,N_1375);
and U5494 (N_5494,N_2433,N_1375);
or U5495 (N_5495,N_1211,N_476);
nand U5496 (N_5496,N_2713,N_702);
xor U5497 (N_5497,N_2964,N_654);
xor U5498 (N_5498,N_2799,N_2727);
or U5499 (N_5499,N_2590,N_2455);
xor U5500 (N_5500,N_1908,N_1882);
nor U5501 (N_5501,N_962,N_1342);
xnor U5502 (N_5502,N_1395,N_1426);
nand U5503 (N_5503,N_1495,N_841);
or U5504 (N_5504,N_1150,N_1222);
or U5505 (N_5505,N_2981,N_1409);
xnor U5506 (N_5506,N_2651,N_1957);
and U5507 (N_5507,N_77,N_1330);
nand U5508 (N_5508,N_391,N_1522);
nand U5509 (N_5509,N_2891,N_1593);
xnor U5510 (N_5510,N_1821,N_2925);
nand U5511 (N_5511,N_1312,N_775);
or U5512 (N_5512,N_2642,N_1905);
and U5513 (N_5513,N_139,N_1140);
nand U5514 (N_5514,N_2378,N_890);
nor U5515 (N_5515,N_2846,N_1112);
or U5516 (N_5516,N_1652,N_1455);
nor U5517 (N_5517,N_1565,N_1971);
nand U5518 (N_5518,N_1809,N_2875);
or U5519 (N_5519,N_2197,N_635);
nand U5520 (N_5520,N_1412,N_2719);
xnor U5521 (N_5521,N_764,N_733);
nand U5522 (N_5522,N_2357,N_66);
and U5523 (N_5523,N_2366,N_425);
or U5524 (N_5524,N_2163,N_2052);
or U5525 (N_5525,N_1518,N_1830);
nor U5526 (N_5526,N_476,N_2190);
and U5527 (N_5527,N_707,N_2989);
or U5528 (N_5528,N_1142,N_2353);
nor U5529 (N_5529,N_2504,N_2329);
nor U5530 (N_5530,N_1295,N_157);
nand U5531 (N_5531,N_1279,N_101);
nor U5532 (N_5532,N_2597,N_1591);
nor U5533 (N_5533,N_2905,N_814);
or U5534 (N_5534,N_1823,N_796);
nand U5535 (N_5535,N_8,N_2054);
or U5536 (N_5536,N_612,N_1149);
or U5537 (N_5537,N_457,N_1773);
and U5538 (N_5538,N_1228,N_808);
or U5539 (N_5539,N_1496,N_2319);
xor U5540 (N_5540,N_2526,N_1058);
nand U5541 (N_5541,N_1361,N_494);
and U5542 (N_5542,N_1866,N_2226);
or U5543 (N_5543,N_992,N_1947);
xnor U5544 (N_5544,N_2886,N_1106);
xnor U5545 (N_5545,N_791,N_2268);
xor U5546 (N_5546,N_745,N_669);
or U5547 (N_5547,N_2783,N_855);
nor U5548 (N_5548,N_2950,N_2486);
xor U5549 (N_5549,N_1475,N_669);
nand U5550 (N_5550,N_2661,N_2259);
or U5551 (N_5551,N_2032,N_315);
xor U5552 (N_5552,N_1376,N_1505);
nor U5553 (N_5553,N_1446,N_1793);
nand U5554 (N_5554,N_410,N_352);
xor U5555 (N_5555,N_967,N_991);
xnor U5556 (N_5556,N_1218,N_388);
nand U5557 (N_5557,N_1030,N_2440);
and U5558 (N_5558,N_1862,N_2968);
nor U5559 (N_5559,N_2230,N_2615);
nor U5560 (N_5560,N_2546,N_852);
and U5561 (N_5561,N_2306,N_2508);
and U5562 (N_5562,N_199,N_59);
nand U5563 (N_5563,N_1476,N_1472);
or U5564 (N_5564,N_1960,N_2501);
xor U5565 (N_5565,N_2416,N_644);
or U5566 (N_5566,N_2278,N_2381);
or U5567 (N_5567,N_1795,N_2961);
xnor U5568 (N_5568,N_2820,N_1312);
nor U5569 (N_5569,N_583,N_1764);
nor U5570 (N_5570,N_1768,N_2117);
or U5571 (N_5571,N_2905,N_2976);
and U5572 (N_5572,N_2063,N_868);
or U5573 (N_5573,N_2648,N_1618);
nand U5574 (N_5574,N_430,N_2543);
xnor U5575 (N_5575,N_1663,N_2314);
nor U5576 (N_5576,N_677,N_2496);
xor U5577 (N_5577,N_557,N_2921);
and U5578 (N_5578,N_2274,N_1009);
and U5579 (N_5579,N_660,N_2365);
or U5580 (N_5580,N_1215,N_2766);
and U5581 (N_5581,N_2703,N_654);
nor U5582 (N_5582,N_2566,N_1774);
nand U5583 (N_5583,N_1649,N_542);
and U5584 (N_5584,N_141,N_799);
nand U5585 (N_5585,N_2459,N_2835);
nor U5586 (N_5586,N_2556,N_363);
nand U5587 (N_5587,N_375,N_2209);
and U5588 (N_5588,N_1380,N_2918);
xnor U5589 (N_5589,N_1104,N_21);
nand U5590 (N_5590,N_405,N_2299);
xor U5591 (N_5591,N_2774,N_602);
nand U5592 (N_5592,N_2707,N_1742);
nand U5593 (N_5593,N_1805,N_312);
xor U5594 (N_5594,N_2079,N_1482);
nor U5595 (N_5595,N_1871,N_1662);
or U5596 (N_5596,N_1231,N_364);
and U5597 (N_5597,N_2661,N_1028);
nor U5598 (N_5598,N_1484,N_4);
and U5599 (N_5599,N_414,N_1353);
and U5600 (N_5600,N_1064,N_1205);
nand U5601 (N_5601,N_2404,N_1428);
or U5602 (N_5602,N_137,N_766);
and U5603 (N_5603,N_86,N_1705);
nor U5604 (N_5604,N_195,N_1131);
nor U5605 (N_5605,N_1126,N_2602);
nor U5606 (N_5606,N_426,N_600);
nor U5607 (N_5607,N_157,N_352);
nor U5608 (N_5608,N_1969,N_1994);
nand U5609 (N_5609,N_1843,N_619);
and U5610 (N_5610,N_2707,N_2574);
nand U5611 (N_5611,N_2445,N_2124);
and U5612 (N_5612,N_1649,N_140);
xor U5613 (N_5613,N_2016,N_174);
nor U5614 (N_5614,N_1111,N_1533);
xnor U5615 (N_5615,N_1084,N_1668);
nor U5616 (N_5616,N_2185,N_2303);
or U5617 (N_5617,N_2150,N_1250);
xnor U5618 (N_5618,N_1487,N_1780);
or U5619 (N_5619,N_1319,N_1104);
nand U5620 (N_5620,N_697,N_2956);
or U5621 (N_5621,N_582,N_393);
xor U5622 (N_5622,N_113,N_157);
nor U5623 (N_5623,N_2450,N_504);
nand U5624 (N_5624,N_359,N_1729);
nand U5625 (N_5625,N_2564,N_593);
or U5626 (N_5626,N_765,N_2628);
xor U5627 (N_5627,N_1181,N_2523);
and U5628 (N_5628,N_2095,N_821);
or U5629 (N_5629,N_2581,N_2270);
xor U5630 (N_5630,N_2249,N_2411);
and U5631 (N_5631,N_1172,N_1547);
xor U5632 (N_5632,N_2448,N_133);
xnor U5633 (N_5633,N_2710,N_1618);
xnor U5634 (N_5634,N_2057,N_773);
nor U5635 (N_5635,N_1459,N_42);
nor U5636 (N_5636,N_2367,N_73);
or U5637 (N_5637,N_2188,N_1139);
or U5638 (N_5638,N_63,N_1459);
nor U5639 (N_5639,N_1389,N_265);
xnor U5640 (N_5640,N_818,N_1825);
xnor U5641 (N_5641,N_1332,N_264);
nand U5642 (N_5642,N_729,N_2150);
and U5643 (N_5643,N_395,N_2361);
and U5644 (N_5644,N_1942,N_1466);
nor U5645 (N_5645,N_347,N_492);
and U5646 (N_5646,N_1068,N_963);
nand U5647 (N_5647,N_1297,N_1282);
nand U5648 (N_5648,N_963,N_482);
nor U5649 (N_5649,N_2776,N_766);
nor U5650 (N_5650,N_990,N_2251);
xor U5651 (N_5651,N_1510,N_2594);
xnor U5652 (N_5652,N_2765,N_1361);
nor U5653 (N_5653,N_1530,N_1510);
nand U5654 (N_5654,N_481,N_1332);
xnor U5655 (N_5655,N_129,N_656);
or U5656 (N_5656,N_1949,N_863);
xor U5657 (N_5657,N_999,N_2809);
or U5658 (N_5658,N_2660,N_2423);
or U5659 (N_5659,N_2631,N_1204);
or U5660 (N_5660,N_2925,N_2634);
nand U5661 (N_5661,N_167,N_2801);
and U5662 (N_5662,N_498,N_2745);
nor U5663 (N_5663,N_225,N_121);
or U5664 (N_5664,N_1388,N_39);
nor U5665 (N_5665,N_1196,N_1121);
and U5666 (N_5666,N_1609,N_429);
nand U5667 (N_5667,N_947,N_1559);
or U5668 (N_5668,N_1677,N_610);
xor U5669 (N_5669,N_770,N_1450);
nor U5670 (N_5670,N_830,N_59);
nor U5671 (N_5671,N_1454,N_772);
nor U5672 (N_5672,N_977,N_2834);
and U5673 (N_5673,N_2390,N_2913);
and U5674 (N_5674,N_642,N_2394);
or U5675 (N_5675,N_2824,N_2390);
or U5676 (N_5676,N_677,N_880);
or U5677 (N_5677,N_81,N_1195);
and U5678 (N_5678,N_289,N_1732);
xor U5679 (N_5679,N_2304,N_2513);
or U5680 (N_5680,N_1755,N_2710);
or U5681 (N_5681,N_2218,N_2470);
and U5682 (N_5682,N_475,N_1046);
or U5683 (N_5683,N_1501,N_2218);
and U5684 (N_5684,N_354,N_1535);
and U5685 (N_5685,N_240,N_417);
and U5686 (N_5686,N_964,N_676);
nor U5687 (N_5687,N_2364,N_663);
nand U5688 (N_5688,N_1000,N_1168);
xnor U5689 (N_5689,N_274,N_2784);
nand U5690 (N_5690,N_1003,N_2444);
nor U5691 (N_5691,N_1456,N_2082);
and U5692 (N_5692,N_504,N_2346);
nand U5693 (N_5693,N_8,N_557);
xor U5694 (N_5694,N_1728,N_545);
nand U5695 (N_5695,N_1553,N_469);
or U5696 (N_5696,N_1372,N_338);
nand U5697 (N_5697,N_2123,N_982);
or U5698 (N_5698,N_1800,N_1645);
or U5699 (N_5699,N_1295,N_1945);
xor U5700 (N_5700,N_307,N_1855);
nand U5701 (N_5701,N_1911,N_794);
and U5702 (N_5702,N_1995,N_1094);
and U5703 (N_5703,N_2371,N_636);
and U5704 (N_5704,N_247,N_1315);
or U5705 (N_5705,N_1054,N_812);
or U5706 (N_5706,N_1734,N_1026);
and U5707 (N_5707,N_2330,N_1792);
xnor U5708 (N_5708,N_1511,N_2160);
nand U5709 (N_5709,N_1789,N_796);
xor U5710 (N_5710,N_2583,N_1373);
or U5711 (N_5711,N_1023,N_2044);
nand U5712 (N_5712,N_1599,N_2598);
xnor U5713 (N_5713,N_97,N_1029);
nand U5714 (N_5714,N_1606,N_789);
and U5715 (N_5715,N_2639,N_377);
xnor U5716 (N_5716,N_359,N_2394);
xor U5717 (N_5717,N_116,N_576);
and U5718 (N_5718,N_2566,N_1478);
or U5719 (N_5719,N_2441,N_2541);
nand U5720 (N_5720,N_1209,N_1274);
xnor U5721 (N_5721,N_2757,N_1980);
nor U5722 (N_5722,N_1913,N_292);
xor U5723 (N_5723,N_1579,N_1055);
or U5724 (N_5724,N_652,N_2206);
nand U5725 (N_5725,N_2018,N_1301);
or U5726 (N_5726,N_388,N_782);
or U5727 (N_5727,N_2764,N_2965);
nand U5728 (N_5728,N_2770,N_22);
nor U5729 (N_5729,N_604,N_232);
xnor U5730 (N_5730,N_960,N_893);
and U5731 (N_5731,N_1398,N_38);
xor U5732 (N_5732,N_685,N_69);
or U5733 (N_5733,N_1575,N_758);
xor U5734 (N_5734,N_1341,N_1348);
nor U5735 (N_5735,N_2016,N_1585);
nand U5736 (N_5736,N_2742,N_1486);
and U5737 (N_5737,N_890,N_1886);
nand U5738 (N_5738,N_1028,N_2180);
nand U5739 (N_5739,N_2992,N_1640);
xor U5740 (N_5740,N_2424,N_441);
and U5741 (N_5741,N_2743,N_2099);
nand U5742 (N_5742,N_2022,N_1060);
nor U5743 (N_5743,N_1392,N_1615);
nor U5744 (N_5744,N_528,N_2216);
and U5745 (N_5745,N_2647,N_1577);
and U5746 (N_5746,N_432,N_414);
xnor U5747 (N_5747,N_2909,N_1561);
or U5748 (N_5748,N_1079,N_989);
or U5749 (N_5749,N_2686,N_2337);
xor U5750 (N_5750,N_2821,N_2734);
nand U5751 (N_5751,N_1632,N_1463);
and U5752 (N_5752,N_2262,N_2415);
and U5753 (N_5753,N_2920,N_1319);
and U5754 (N_5754,N_1008,N_1006);
nor U5755 (N_5755,N_2583,N_1351);
xor U5756 (N_5756,N_1012,N_1597);
nand U5757 (N_5757,N_291,N_1863);
nor U5758 (N_5758,N_2511,N_2928);
and U5759 (N_5759,N_1640,N_91);
nand U5760 (N_5760,N_2458,N_2841);
nand U5761 (N_5761,N_1384,N_209);
nand U5762 (N_5762,N_1049,N_2695);
or U5763 (N_5763,N_57,N_1799);
nor U5764 (N_5764,N_97,N_1058);
and U5765 (N_5765,N_824,N_2427);
nor U5766 (N_5766,N_2125,N_1270);
xor U5767 (N_5767,N_2969,N_2645);
or U5768 (N_5768,N_487,N_677);
or U5769 (N_5769,N_855,N_388);
xor U5770 (N_5770,N_299,N_2478);
or U5771 (N_5771,N_209,N_520);
and U5772 (N_5772,N_2429,N_1209);
nand U5773 (N_5773,N_2782,N_1338);
and U5774 (N_5774,N_366,N_1918);
and U5775 (N_5775,N_1307,N_801);
and U5776 (N_5776,N_1735,N_2603);
or U5777 (N_5777,N_686,N_2765);
or U5778 (N_5778,N_1885,N_979);
nor U5779 (N_5779,N_2172,N_2016);
or U5780 (N_5780,N_2640,N_460);
and U5781 (N_5781,N_2661,N_2484);
or U5782 (N_5782,N_2801,N_1343);
xor U5783 (N_5783,N_2650,N_2024);
and U5784 (N_5784,N_2499,N_2721);
or U5785 (N_5785,N_568,N_1313);
nor U5786 (N_5786,N_1875,N_2210);
xnor U5787 (N_5787,N_2940,N_1942);
or U5788 (N_5788,N_1562,N_1389);
nand U5789 (N_5789,N_2308,N_48);
and U5790 (N_5790,N_2047,N_2655);
or U5791 (N_5791,N_2601,N_999);
xnor U5792 (N_5792,N_260,N_1841);
xnor U5793 (N_5793,N_1938,N_2754);
and U5794 (N_5794,N_987,N_2652);
xnor U5795 (N_5795,N_1965,N_2799);
xor U5796 (N_5796,N_1925,N_2436);
nand U5797 (N_5797,N_854,N_399);
and U5798 (N_5798,N_1736,N_1241);
and U5799 (N_5799,N_2887,N_2770);
and U5800 (N_5800,N_2225,N_2229);
nor U5801 (N_5801,N_1427,N_149);
nand U5802 (N_5802,N_1229,N_956);
and U5803 (N_5803,N_2327,N_218);
nor U5804 (N_5804,N_2469,N_1608);
nor U5805 (N_5805,N_1726,N_1691);
nor U5806 (N_5806,N_2615,N_2192);
or U5807 (N_5807,N_1127,N_599);
nor U5808 (N_5808,N_706,N_1486);
and U5809 (N_5809,N_512,N_1021);
nor U5810 (N_5810,N_2116,N_1890);
nor U5811 (N_5811,N_2466,N_732);
xnor U5812 (N_5812,N_663,N_1992);
or U5813 (N_5813,N_1285,N_139);
nor U5814 (N_5814,N_557,N_527);
or U5815 (N_5815,N_2662,N_2070);
nor U5816 (N_5816,N_1865,N_576);
or U5817 (N_5817,N_1763,N_2924);
and U5818 (N_5818,N_1833,N_709);
nand U5819 (N_5819,N_944,N_1454);
and U5820 (N_5820,N_2770,N_2793);
and U5821 (N_5821,N_220,N_420);
xnor U5822 (N_5822,N_863,N_574);
xnor U5823 (N_5823,N_982,N_78);
or U5824 (N_5824,N_2664,N_1606);
xnor U5825 (N_5825,N_2021,N_1270);
nand U5826 (N_5826,N_2271,N_2595);
and U5827 (N_5827,N_167,N_1679);
xor U5828 (N_5828,N_826,N_754);
nand U5829 (N_5829,N_2491,N_322);
or U5830 (N_5830,N_1057,N_821);
or U5831 (N_5831,N_282,N_272);
xnor U5832 (N_5832,N_1854,N_2401);
xor U5833 (N_5833,N_1631,N_1459);
nor U5834 (N_5834,N_1377,N_841);
or U5835 (N_5835,N_1411,N_24);
xor U5836 (N_5836,N_535,N_2100);
nor U5837 (N_5837,N_314,N_1614);
or U5838 (N_5838,N_725,N_2753);
nor U5839 (N_5839,N_1914,N_2994);
xnor U5840 (N_5840,N_2976,N_1971);
or U5841 (N_5841,N_1112,N_736);
nand U5842 (N_5842,N_606,N_890);
xnor U5843 (N_5843,N_2147,N_2801);
nand U5844 (N_5844,N_1540,N_410);
and U5845 (N_5845,N_1391,N_736);
xor U5846 (N_5846,N_525,N_1941);
nand U5847 (N_5847,N_1978,N_701);
nand U5848 (N_5848,N_342,N_594);
xnor U5849 (N_5849,N_854,N_246);
nor U5850 (N_5850,N_231,N_1631);
xnor U5851 (N_5851,N_1120,N_325);
or U5852 (N_5852,N_1871,N_2811);
xor U5853 (N_5853,N_670,N_1406);
or U5854 (N_5854,N_2159,N_901);
xnor U5855 (N_5855,N_774,N_616);
nand U5856 (N_5856,N_2853,N_303);
nand U5857 (N_5857,N_1614,N_2362);
xnor U5858 (N_5858,N_1216,N_1136);
and U5859 (N_5859,N_2644,N_1016);
or U5860 (N_5860,N_2016,N_1932);
or U5861 (N_5861,N_2758,N_2349);
and U5862 (N_5862,N_361,N_491);
or U5863 (N_5863,N_2823,N_573);
or U5864 (N_5864,N_366,N_1083);
or U5865 (N_5865,N_2315,N_1591);
nor U5866 (N_5866,N_2346,N_229);
or U5867 (N_5867,N_2376,N_1255);
nor U5868 (N_5868,N_221,N_2045);
nor U5869 (N_5869,N_709,N_2239);
nand U5870 (N_5870,N_1434,N_1138);
nand U5871 (N_5871,N_2552,N_19);
and U5872 (N_5872,N_2672,N_940);
and U5873 (N_5873,N_924,N_2175);
or U5874 (N_5874,N_2660,N_1237);
nand U5875 (N_5875,N_1012,N_2295);
xnor U5876 (N_5876,N_2204,N_2629);
nor U5877 (N_5877,N_349,N_2079);
nand U5878 (N_5878,N_1881,N_2397);
xor U5879 (N_5879,N_829,N_1819);
xor U5880 (N_5880,N_931,N_1497);
nor U5881 (N_5881,N_2301,N_2541);
and U5882 (N_5882,N_1622,N_1241);
xor U5883 (N_5883,N_2934,N_1197);
nor U5884 (N_5884,N_1579,N_2883);
and U5885 (N_5885,N_615,N_2422);
nand U5886 (N_5886,N_976,N_2517);
xnor U5887 (N_5887,N_354,N_2811);
nand U5888 (N_5888,N_112,N_2762);
or U5889 (N_5889,N_1131,N_1796);
nor U5890 (N_5890,N_942,N_2047);
or U5891 (N_5891,N_691,N_1421);
and U5892 (N_5892,N_824,N_225);
or U5893 (N_5893,N_1941,N_2523);
xnor U5894 (N_5894,N_1993,N_1481);
xnor U5895 (N_5895,N_2354,N_1762);
or U5896 (N_5896,N_2246,N_2006);
nand U5897 (N_5897,N_785,N_1539);
and U5898 (N_5898,N_459,N_1839);
xor U5899 (N_5899,N_1106,N_157);
and U5900 (N_5900,N_1004,N_833);
xor U5901 (N_5901,N_1108,N_1041);
nor U5902 (N_5902,N_453,N_559);
nor U5903 (N_5903,N_2925,N_2949);
and U5904 (N_5904,N_941,N_2055);
xor U5905 (N_5905,N_1807,N_2925);
and U5906 (N_5906,N_1237,N_2701);
or U5907 (N_5907,N_713,N_2061);
and U5908 (N_5908,N_567,N_1665);
and U5909 (N_5909,N_2509,N_2249);
nor U5910 (N_5910,N_1313,N_2732);
and U5911 (N_5911,N_731,N_1353);
xor U5912 (N_5912,N_485,N_1739);
or U5913 (N_5913,N_1483,N_1984);
nand U5914 (N_5914,N_711,N_1627);
or U5915 (N_5915,N_2587,N_817);
or U5916 (N_5916,N_2943,N_889);
and U5917 (N_5917,N_2118,N_2675);
or U5918 (N_5918,N_1230,N_851);
nand U5919 (N_5919,N_2733,N_1438);
or U5920 (N_5920,N_8,N_135);
or U5921 (N_5921,N_1521,N_2943);
nand U5922 (N_5922,N_2434,N_1585);
nor U5923 (N_5923,N_2835,N_2600);
or U5924 (N_5924,N_1756,N_2335);
and U5925 (N_5925,N_2815,N_2608);
and U5926 (N_5926,N_1104,N_2491);
nand U5927 (N_5927,N_1244,N_2398);
nand U5928 (N_5928,N_2251,N_1752);
nor U5929 (N_5929,N_1527,N_1589);
nand U5930 (N_5930,N_523,N_2491);
nor U5931 (N_5931,N_2485,N_558);
and U5932 (N_5932,N_1058,N_209);
or U5933 (N_5933,N_601,N_2469);
nand U5934 (N_5934,N_710,N_371);
nand U5935 (N_5935,N_1956,N_2426);
xor U5936 (N_5936,N_2181,N_2509);
and U5937 (N_5937,N_780,N_1326);
xnor U5938 (N_5938,N_494,N_1163);
nor U5939 (N_5939,N_2823,N_2465);
xor U5940 (N_5940,N_2320,N_2020);
nand U5941 (N_5941,N_336,N_968);
nand U5942 (N_5942,N_374,N_2927);
nor U5943 (N_5943,N_1863,N_1474);
or U5944 (N_5944,N_504,N_2920);
xnor U5945 (N_5945,N_2239,N_1071);
nand U5946 (N_5946,N_1463,N_2889);
or U5947 (N_5947,N_2662,N_526);
nor U5948 (N_5948,N_860,N_1983);
or U5949 (N_5949,N_0,N_108);
nand U5950 (N_5950,N_1119,N_699);
or U5951 (N_5951,N_778,N_2384);
and U5952 (N_5952,N_2376,N_1424);
xnor U5953 (N_5953,N_1826,N_2240);
xor U5954 (N_5954,N_64,N_50);
or U5955 (N_5955,N_562,N_2961);
nor U5956 (N_5956,N_737,N_2398);
or U5957 (N_5957,N_1256,N_439);
and U5958 (N_5958,N_1604,N_1763);
nand U5959 (N_5959,N_432,N_1691);
xor U5960 (N_5960,N_675,N_1949);
or U5961 (N_5961,N_2103,N_113);
xor U5962 (N_5962,N_2460,N_2562);
and U5963 (N_5963,N_1077,N_670);
nor U5964 (N_5964,N_635,N_273);
nand U5965 (N_5965,N_811,N_1179);
nor U5966 (N_5966,N_64,N_2137);
xnor U5967 (N_5967,N_2611,N_1654);
or U5968 (N_5968,N_613,N_2254);
xnor U5969 (N_5969,N_1110,N_1220);
nor U5970 (N_5970,N_1880,N_50);
xor U5971 (N_5971,N_2145,N_634);
xnor U5972 (N_5972,N_2527,N_2427);
and U5973 (N_5973,N_1212,N_343);
nor U5974 (N_5974,N_858,N_2739);
nand U5975 (N_5975,N_2846,N_1831);
or U5976 (N_5976,N_946,N_577);
xor U5977 (N_5977,N_2629,N_2038);
or U5978 (N_5978,N_1307,N_107);
and U5979 (N_5979,N_2835,N_1137);
or U5980 (N_5980,N_2420,N_2869);
and U5981 (N_5981,N_322,N_1665);
nand U5982 (N_5982,N_1343,N_1228);
xor U5983 (N_5983,N_603,N_186);
or U5984 (N_5984,N_2626,N_347);
nor U5985 (N_5985,N_1310,N_2549);
nor U5986 (N_5986,N_1884,N_1424);
and U5987 (N_5987,N_2335,N_2043);
nand U5988 (N_5988,N_1730,N_688);
nor U5989 (N_5989,N_1560,N_2256);
nand U5990 (N_5990,N_1669,N_358);
and U5991 (N_5991,N_2763,N_1795);
nand U5992 (N_5992,N_2416,N_655);
nand U5993 (N_5993,N_2126,N_2107);
xnor U5994 (N_5994,N_231,N_1126);
and U5995 (N_5995,N_2855,N_1216);
and U5996 (N_5996,N_1607,N_1731);
nor U5997 (N_5997,N_2340,N_1023);
nand U5998 (N_5998,N_889,N_207);
nor U5999 (N_5999,N_2941,N_778);
or U6000 (N_6000,N_3292,N_3507);
xnor U6001 (N_6001,N_5771,N_5138);
nor U6002 (N_6002,N_3181,N_4949);
nor U6003 (N_6003,N_3733,N_4494);
xor U6004 (N_6004,N_3314,N_3684);
and U6005 (N_6005,N_3248,N_4327);
and U6006 (N_6006,N_3360,N_4778);
nand U6007 (N_6007,N_3755,N_4332);
or U6008 (N_6008,N_4013,N_5052);
nor U6009 (N_6009,N_4873,N_4884);
xor U6010 (N_6010,N_4426,N_5691);
nand U6011 (N_6011,N_5146,N_5063);
nor U6012 (N_6012,N_3571,N_3361);
xor U6013 (N_6013,N_5089,N_5974);
nand U6014 (N_6014,N_4608,N_5364);
xnor U6015 (N_6015,N_4093,N_5024);
nor U6016 (N_6016,N_4680,N_3878);
nor U6017 (N_6017,N_4509,N_4697);
or U6018 (N_6018,N_3928,N_4307);
nor U6019 (N_6019,N_5312,N_4811);
nand U6020 (N_6020,N_4367,N_3669);
nand U6021 (N_6021,N_3392,N_5406);
nor U6022 (N_6022,N_3862,N_5445);
xor U6023 (N_6023,N_4766,N_5207);
or U6024 (N_6024,N_4254,N_4591);
nand U6025 (N_6025,N_4381,N_3494);
and U6026 (N_6026,N_3947,N_4663);
xnor U6027 (N_6027,N_4049,N_4097);
and U6028 (N_6028,N_3979,N_3382);
or U6029 (N_6029,N_4495,N_3816);
nand U6030 (N_6030,N_3994,N_3830);
nor U6031 (N_6031,N_4530,N_5893);
nor U6032 (N_6032,N_5096,N_5431);
xor U6033 (N_6033,N_4890,N_5056);
xor U6034 (N_6034,N_5291,N_5922);
or U6035 (N_6035,N_4443,N_5323);
or U6036 (N_6036,N_4649,N_3868);
and U6037 (N_6037,N_3982,N_5214);
and U6038 (N_6038,N_4127,N_3347);
nand U6039 (N_6039,N_4893,N_5812);
nand U6040 (N_6040,N_5444,N_5514);
nor U6041 (N_6041,N_3333,N_3045);
nor U6042 (N_6042,N_5506,N_4411);
xor U6043 (N_6043,N_5318,N_5645);
and U6044 (N_6044,N_5826,N_4704);
or U6045 (N_6045,N_3387,N_5757);
xnor U6046 (N_6046,N_3728,N_5171);
nand U6047 (N_6047,N_5767,N_5695);
nor U6048 (N_6048,N_5789,N_3604);
nor U6049 (N_6049,N_3964,N_4405);
or U6050 (N_6050,N_5702,N_5047);
nor U6051 (N_6051,N_3231,N_4971);
xor U6052 (N_6052,N_4669,N_5053);
and U6053 (N_6053,N_5865,N_5864);
or U6054 (N_6054,N_3534,N_5519);
nand U6055 (N_6055,N_5746,N_3552);
nand U6056 (N_6056,N_3154,N_5688);
and U6057 (N_6057,N_5629,N_3495);
and U6058 (N_6058,N_4109,N_4805);
or U6059 (N_6059,N_5128,N_5566);
nand U6060 (N_6060,N_5238,N_3601);
nand U6061 (N_6061,N_4939,N_5015);
nand U6062 (N_6062,N_5689,N_3431);
nand U6063 (N_6063,N_5124,N_3636);
or U6064 (N_6064,N_3024,N_5496);
nor U6065 (N_6065,N_4456,N_5577);
nand U6066 (N_6066,N_4902,N_3734);
or U6067 (N_6067,N_3567,N_3528);
xnor U6068 (N_6068,N_5429,N_3648);
or U6069 (N_6069,N_3704,N_3961);
nand U6070 (N_6070,N_5031,N_5191);
xnor U6071 (N_6071,N_4035,N_3933);
nor U6072 (N_6072,N_5930,N_4803);
nand U6073 (N_6073,N_3397,N_5665);
and U6074 (N_6074,N_5532,N_3771);
or U6075 (N_6075,N_4396,N_5565);
nand U6076 (N_6076,N_4115,N_3653);
and U6077 (N_6077,N_5973,N_4611);
nand U6078 (N_6078,N_3168,N_5121);
and U6079 (N_6079,N_3038,N_3877);
nand U6080 (N_6080,N_4534,N_5280);
nand U6081 (N_6081,N_5180,N_3004);
or U6082 (N_6082,N_4918,N_4785);
or U6083 (N_6083,N_3092,N_5265);
or U6084 (N_6084,N_5725,N_5741);
nand U6085 (N_6085,N_5260,N_3677);
nor U6086 (N_6086,N_4906,N_5393);
and U6087 (N_6087,N_3536,N_3195);
and U6088 (N_6088,N_4600,N_5273);
and U6089 (N_6089,N_4603,N_4636);
nand U6090 (N_6090,N_5547,N_5244);
and U6091 (N_6091,N_3673,N_3237);
nand U6092 (N_6092,N_5655,N_4172);
and U6093 (N_6093,N_3535,N_3419);
or U6094 (N_6094,N_3707,N_4877);
and U6095 (N_6095,N_5742,N_5115);
xnor U6096 (N_6096,N_5871,N_3574);
nand U6097 (N_6097,N_4905,N_4291);
and U6098 (N_6098,N_3941,N_3517);
nand U6099 (N_6099,N_3548,N_5882);
nor U6100 (N_6100,N_4804,N_3859);
or U6101 (N_6101,N_5360,N_4794);
xor U6102 (N_6102,N_3581,N_5768);
or U6103 (N_6103,N_4769,N_5349);
or U6104 (N_6104,N_5550,N_3124);
xor U6105 (N_6105,N_5411,N_4650);
nand U6106 (N_6106,N_5996,N_4656);
or U6107 (N_6107,N_3950,N_4023);
nor U6108 (N_6108,N_4233,N_3336);
xnor U6109 (N_6109,N_3825,N_5723);
nor U6110 (N_6110,N_4505,N_4612);
and U6111 (N_6111,N_3269,N_4862);
and U6112 (N_6112,N_4853,N_3044);
or U6113 (N_6113,N_3254,N_4843);
nor U6114 (N_6114,N_4057,N_4928);
and U6115 (N_6115,N_5600,N_3630);
or U6116 (N_6116,N_4595,N_3803);
xor U6117 (N_6117,N_3132,N_3914);
nand U6118 (N_6118,N_4437,N_3641);
nor U6119 (N_6119,N_4101,N_3564);
xnor U6120 (N_6120,N_4496,N_3695);
or U6121 (N_6121,N_5734,N_5989);
nand U6122 (N_6122,N_3433,N_4406);
and U6123 (N_6123,N_4980,N_5716);
nor U6124 (N_6124,N_3430,N_4734);
xor U6125 (N_6125,N_4909,N_5717);
or U6126 (N_6126,N_5251,N_5888);
or U6127 (N_6127,N_4026,N_4130);
nand U6128 (N_6128,N_4310,N_5891);
or U6129 (N_6129,N_5542,N_5956);
xor U6130 (N_6130,N_4768,N_4226);
xnor U6131 (N_6131,N_5325,N_5857);
xor U6132 (N_6132,N_4576,N_3180);
and U6133 (N_6133,N_3876,N_4249);
nand U6134 (N_6134,N_4468,N_5963);
xnor U6135 (N_6135,N_3052,N_5525);
and U6136 (N_6136,N_5708,N_4925);
or U6137 (N_6137,N_4104,N_5567);
xnor U6138 (N_6138,N_4467,N_3139);
nand U6139 (N_6139,N_4086,N_4385);
nor U6140 (N_6140,N_5611,N_4347);
nor U6141 (N_6141,N_3227,N_4126);
xor U6142 (N_6142,N_3224,N_3870);
or U6143 (N_6143,N_3946,N_4683);
xnor U6144 (N_6144,N_3490,N_5476);
xor U6145 (N_6145,N_4724,N_4072);
or U6146 (N_6146,N_5537,N_3986);
xor U6147 (N_6147,N_4537,N_5553);
xor U6148 (N_6148,N_4485,N_4976);
xor U6149 (N_6149,N_5879,N_5668);
nor U6150 (N_6150,N_5198,N_5184);
and U6151 (N_6151,N_3306,N_3245);
nor U6152 (N_6152,N_3512,N_3988);
nor U6153 (N_6153,N_5042,N_5926);
nand U6154 (N_6154,N_5559,N_4229);
or U6155 (N_6155,N_5187,N_4914);
or U6156 (N_6156,N_4222,N_4465);
nor U6157 (N_6157,N_3896,N_4297);
and U6158 (N_6158,N_4434,N_3579);
and U6159 (N_6159,N_4190,N_5143);
or U6160 (N_6160,N_4507,N_4904);
xor U6161 (N_6161,N_5841,N_5833);
or U6162 (N_6162,N_5797,N_3573);
nand U6163 (N_6163,N_3133,N_3094);
nand U6164 (N_6164,N_3644,N_3294);
nor U6165 (N_6165,N_3839,N_4211);
nor U6166 (N_6166,N_3752,N_5202);
or U6167 (N_6167,N_5793,N_3748);
and U6168 (N_6168,N_4103,N_5100);
nand U6169 (N_6169,N_4299,N_4899);
nand U6170 (N_6170,N_4816,N_5382);
xor U6171 (N_6171,N_5275,N_3422);
xnor U6172 (N_6172,N_5549,N_5412);
xnor U6173 (N_6173,N_5731,N_3799);
nand U6174 (N_6174,N_5007,N_3034);
or U6175 (N_6175,N_3193,N_5610);
or U6176 (N_6176,N_3220,N_4008);
and U6177 (N_6177,N_4205,N_5212);
xnor U6178 (N_6178,N_5447,N_3781);
and U6179 (N_6179,N_4732,N_3190);
or U6180 (N_6180,N_5813,N_5872);
and U6181 (N_6181,N_5536,N_5483);
or U6182 (N_6182,N_3712,N_3940);
nand U6183 (N_6183,N_4316,N_5803);
nand U6184 (N_6184,N_3861,N_4635);
xnor U6185 (N_6185,N_3289,N_5590);
or U6186 (N_6186,N_5441,N_4851);
xnor U6187 (N_6187,N_4662,N_4060);
xor U6188 (N_6188,N_4464,N_5269);
nand U6189 (N_6189,N_5983,N_5898);
xnor U6190 (N_6190,N_3802,N_4184);
or U6191 (N_6191,N_3112,N_4753);
nor U6192 (N_6192,N_3867,N_3118);
nor U6193 (N_6193,N_4919,N_5173);
nor U6194 (N_6194,N_3499,N_3539);
xnor U6195 (N_6195,N_4675,N_5246);
nor U6196 (N_6196,N_3588,N_3957);
nor U6197 (N_6197,N_3339,N_3883);
nand U6198 (N_6198,N_5423,N_3332);
and U6199 (N_6199,N_5909,N_5924);
and U6200 (N_6200,N_5576,N_3123);
and U6201 (N_6201,N_5800,N_3087);
and U6202 (N_6202,N_4000,N_4374);
or U6203 (N_6203,N_4501,N_5675);
or U6204 (N_6204,N_4741,N_3892);
or U6205 (N_6205,N_3386,N_5092);
xor U6206 (N_6206,N_3683,N_4720);
and U6207 (N_6207,N_5563,N_4099);
and U6208 (N_6208,N_4538,N_4022);
and U6209 (N_6209,N_4053,N_4598);
nor U6210 (N_6210,N_5978,N_4395);
or U6211 (N_6211,N_5463,N_3807);
nor U6212 (N_6212,N_5527,N_5961);
xor U6213 (N_6213,N_5736,N_5966);
nand U6214 (N_6214,N_3889,N_4373);
or U6215 (N_6215,N_4874,N_4480);
nor U6216 (N_6216,N_3836,N_4784);
and U6217 (N_6217,N_4339,N_3182);
and U6218 (N_6218,N_3253,N_4214);
nor U6219 (N_6219,N_4071,N_4318);
xor U6220 (N_6220,N_3189,N_3186);
or U6221 (N_6221,N_4627,N_5418);
nand U6222 (N_6222,N_5132,N_4065);
or U6223 (N_6223,N_3760,N_4440);
xor U6224 (N_6224,N_5086,N_3596);
nand U6225 (N_6225,N_3155,N_3432);
or U6226 (N_6226,N_5125,N_4850);
and U6227 (N_6227,N_5233,N_5058);
nand U6228 (N_6228,N_3616,N_5883);
nor U6229 (N_6229,N_3925,N_4558);
xnor U6230 (N_6230,N_5938,N_4881);
xnor U6231 (N_6231,N_5127,N_3672);
nor U6232 (N_6232,N_4003,N_5947);
and U6233 (N_6233,N_5658,N_3675);
or U6234 (N_6234,N_3015,N_4116);
nand U6235 (N_6235,N_4353,N_3320);
xnor U6236 (N_6236,N_5054,N_3054);
and U6237 (N_6237,N_5510,N_5111);
and U6238 (N_6238,N_5846,N_4564);
nand U6239 (N_6239,N_5057,N_5150);
nand U6240 (N_6240,N_5439,N_4247);
nand U6241 (N_6241,N_5928,N_4380);
or U6242 (N_6242,N_3510,N_3486);
or U6243 (N_6243,N_3820,N_5578);
xnor U6244 (N_6244,N_3468,N_4751);
xor U6245 (N_6245,N_3362,N_4015);
nand U6246 (N_6246,N_4963,N_5616);
nand U6247 (N_6247,N_3886,N_4965);
nand U6248 (N_6248,N_3553,N_4552);
nor U6249 (N_6249,N_4189,N_5270);
xnor U6250 (N_6250,N_4819,N_4163);
or U6251 (N_6251,N_3225,N_4799);
or U6252 (N_6252,N_5038,N_3146);
or U6253 (N_6253,N_5209,N_3238);
nand U6254 (N_6254,N_5597,N_5461);
nor U6255 (N_6255,N_3282,N_3016);
nor U6256 (N_6256,N_4298,N_4364);
nor U6257 (N_6257,N_4333,N_5422);
or U6258 (N_6258,N_3716,N_5558);
nand U6259 (N_6259,N_4975,N_4516);
nand U6260 (N_6260,N_3984,N_5501);
xor U6261 (N_6261,N_3954,N_3444);
xnor U6262 (N_6262,N_5706,N_5845);
nor U6263 (N_6263,N_5779,N_3843);
and U6264 (N_6264,N_4712,N_5080);
nor U6265 (N_6265,N_5556,N_5607);
nor U6266 (N_6266,N_5452,N_3547);
and U6267 (N_6267,N_5427,N_5359);
nand U6268 (N_6268,N_5377,N_3801);
and U6269 (N_6269,N_5962,N_3256);
nor U6270 (N_6270,N_4498,N_5249);
nor U6271 (N_6271,N_5149,N_4394);
xnor U6272 (N_6272,N_3879,N_3584);
nand U6273 (N_6273,N_3334,N_3491);
xor U6274 (N_6274,N_3503,N_3809);
and U6275 (N_6275,N_3021,N_3855);
nor U6276 (N_6276,N_3600,N_4639);
xnor U6277 (N_6277,N_4442,N_5298);
and U6278 (N_6278,N_4688,N_5808);
and U6279 (N_6279,N_4482,N_3068);
and U6280 (N_6280,N_5314,N_4594);
xnor U6281 (N_6281,N_5315,N_4221);
nand U6282 (N_6282,N_4575,N_3773);
or U6283 (N_6283,N_4533,N_3980);
and U6284 (N_6284,N_5794,N_5224);
or U6285 (N_6285,N_3911,N_3219);
nand U6286 (N_6286,N_5859,N_4856);
nor U6287 (N_6287,N_5262,N_3624);
nor U6288 (N_6288,N_3597,N_5199);
and U6289 (N_6289,N_3291,N_4164);
nand U6290 (N_6290,N_4240,N_5862);
xnor U6291 (N_6291,N_4838,N_4593);
nor U6292 (N_6292,N_3632,N_5585);
xor U6293 (N_6293,N_3647,N_4759);
or U6294 (N_6294,N_4828,N_4752);
xor U6295 (N_6295,N_3960,N_3147);
nand U6296 (N_6296,N_3117,N_5321);
or U6297 (N_6297,N_5016,N_5489);
and U6298 (N_6298,N_3770,N_4666);
and U6299 (N_6299,N_4050,N_4266);
and U6300 (N_6300,N_5420,N_3390);
nand U6301 (N_6301,N_4416,N_4152);
nor U6302 (N_6302,N_4984,N_4346);
or U6303 (N_6303,N_3795,N_3818);
nand U6304 (N_6304,N_5440,N_5048);
and U6305 (N_6305,N_5105,N_3720);
xnor U6306 (N_6306,N_3711,N_4998);
xnor U6307 (N_6307,N_3049,N_5247);
or U6308 (N_6308,N_3909,N_3524);
and U6309 (N_6309,N_4895,N_5643);
or U6310 (N_6310,N_4772,N_5028);
or U6311 (N_6311,N_4055,N_3126);
nor U6312 (N_6312,N_4324,N_5261);
nand U6313 (N_6313,N_3834,N_5686);
nor U6314 (N_6314,N_3039,N_5030);
and U6315 (N_6315,N_5976,N_4774);
xor U6316 (N_6316,N_3963,N_5331);
nand U6317 (N_6317,N_5334,N_4541);
nor U6318 (N_6318,N_5448,N_4973);
xor U6319 (N_6319,N_5732,N_4710);
xnor U6320 (N_6320,N_3208,N_3369);
nor U6321 (N_6321,N_5304,N_3663);
nor U6322 (N_6322,N_3585,N_3939);
and U6323 (N_6323,N_3657,N_5534);
nand U6324 (N_6324,N_3128,N_4520);
or U6325 (N_6325,N_3797,N_5917);
nor U6326 (N_6326,N_3586,N_3860);
and U6327 (N_6327,N_5097,N_3767);
or U6328 (N_6328,N_3262,N_3266);
or U6329 (N_6329,N_3913,N_4356);
xor U6330 (N_6330,N_4641,N_4922);
or U6331 (N_6331,N_3625,N_5497);
xor U6332 (N_6332,N_4376,N_4755);
xor U6333 (N_6333,N_3810,N_5669);
or U6334 (N_6334,N_3204,N_4673);
nand U6335 (N_6335,N_4160,N_5851);
xor U6336 (N_6336,N_3152,N_5217);
xnor U6337 (N_6337,N_4502,N_4959);
xor U6338 (N_6338,N_3005,N_4589);
xor U6339 (N_6339,N_5329,N_4786);
and U6340 (N_6340,N_3456,N_5977);
or U6341 (N_6341,N_4714,N_4542);
nor U6342 (N_6342,N_3523,N_4891);
nand U6343 (N_6343,N_5613,N_3001);
xnor U6344 (N_6344,N_3281,N_3040);
or U6345 (N_6345,N_5894,N_4111);
nand U6346 (N_6346,N_3840,N_3633);
nand U6347 (N_6347,N_4342,N_5151);
xnor U6348 (N_6348,N_3140,N_5581);
xor U6349 (N_6349,N_3285,N_4349);
nand U6350 (N_6350,N_5798,N_3077);
nand U6351 (N_6351,N_4585,N_5009);
nor U6352 (N_6352,N_3451,N_5988);
nor U6353 (N_6353,N_5035,N_3022);
xnor U6354 (N_6354,N_5751,N_4609);
or U6355 (N_6355,N_4684,N_5625);
nand U6356 (N_6356,N_3295,N_4757);
or U6357 (N_6357,N_5230,N_3981);
xor U6358 (N_6358,N_5433,N_4698);
nor U6359 (N_6359,N_4117,N_4835);
nand U6360 (N_6360,N_5059,N_4739);
xnor U6361 (N_6361,N_5599,N_4045);
or U6362 (N_6362,N_3541,N_4671);
nor U6363 (N_6363,N_3283,N_3882);
xnor U6364 (N_6364,N_4849,N_5965);
xnor U6365 (N_6365,N_5698,N_5477);
nor U6366 (N_6366,N_5823,N_5679);
xor U6367 (N_6367,N_4889,N_4510);
nor U6368 (N_6368,N_5253,N_4308);
nor U6369 (N_6369,N_4281,N_5034);
nand U6370 (N_6370,N_4460,N_3342);
or U6371 (N_6371,N_4863,N_3097);
nand U6372 (N_6372,N_4942,N_4438);
or U6373 (N_6373,N_4279,N_5182);
xnor U6374 (N_6374,N_4679,N_5432);
nand U6375 (N_6375,N_3265,N_3837);
nor U6376 (N_6376,N_4210,N_3470);
or U6377 (N_6377,N_3041,N_3096);
and U6378 (N_6378,N_4454,N_5997);
and U6379 (N_6379,N_5093,N_4119);
and U6380 (N_6380,N_4936,N_5934);
nand U6381 (N_6381,N_3741,N_5667);
or U6382 (N_6382,N_4717,N_3165);
and U6383 (N_6383,N_5484,N_4536);
nand U6384 (N_6384,N_4602,N_3335);
or U6385 (N_6385,N_4133,N_3099);
xor U6386 (N_6386,N_5367,N_4244);
nand U6387 (N_6387,N_3628,N_4039);
or U6388 (N_6388,N_4178,N_5328);
nor U6389 (N_6389,N_4253,N_3305);
xnor U6390 (N_6390,N_3263,N_5868);
or U6391 (N_6391,N_5912,N_3206);
xor U6392 (N_6392,N_5861,N_5958);
nand U6393 (N_6393,N_3903,N_4319);
nand U6394 (N_6394,N_3131,N_3620);
or U6395 (N_6395,N_3977,N_4791);
and U6396 (N_6396,N_4660,N_3023);
or U6397 (N_6397,N_3176,N_4470);
nor U6398 (N_6398,N_3838,N_4392);
nand U6399 (N_6399,N_4232,N_5979);
or U6400 (N_6400,N_5266,N_3813);
or U6401 (N_6401,N_3638,N_5672);
nand U6402 (N_6402,N_4486,N_4449);
xnor U6403 (N_6403,N_3458,N_3153);
nand U6404 (N_6404,N_5417,N_3768);
or U6405 (N_6405,N_5903,N_4156);
and U6406 (N_6406,N_4958,N_3401);
or U6407 (N_6407,N_5579,N_5885);
and U6408 (N_6408,N_4883,N_4417);
nand U6409 (N_6409,N_5752,N_5758);
nor U6410 (N_6410,N_5221,N_3464);
and U6411 (N_6411,N_5719,N_3693);
nand U6412 (N_6412,N_4387,N_4623);
nand U6413 (N_6413,N_3806,N_4361);
nor U6414 (N_6414,N_4457,N_4568);
and U6415 (N_6415,N_5811,N_4458);
or U6416 (N_6416,N_4944,N_3095);
nor U6417 (N_6417,N_3384,N_4581);
xor U6418 (N_6418,N_3776,N_4667);
xnor U6419 (N_6419,N_4615,N_5967);
or U6420 (N_6420,N_4379,N_5913);
and U6421 (N_6421,N_3739,N_5620);
and U6422 (N_6422,N_5013,N_4605);
xnor U6423 (N_6423,N_4999,N_4617);
and U6424 (N_6424,N_5512,N_5470);
nor U6425 (N_6425,N_5941,N_5641);
nand U6426 (N_6426,N_4900,N_4582);
xnor U6427 (N_6427,N_3047,N_5019);
nor U6428 (N_6428,N_5819,N_3849);
xor U6429 (N_6429,N_5469,N_5396);
or U6430 (N_6430,N_5674,N_3798);
xor U6431 (N_6431,N_4224,N_4185);
xor U6432 (N_6432,N_5374,N_5206);
nor U6433 (N_6433,N_4265,N_5921);
nor U6434 (N_6434,N_4511,N_4020);
nor U6435 (N_6435,N_3053,N_4798);
and U6436 (N_6436,N_3061,N_5853);
nor U6437 (N_6437,N_5055,N_4446);
xnor U6438 (N_6438,N_5436,N_4122);
and U6439 (N_6439,N_3377,N_3679);
nor U6440 (N_6440,N_5095,N_3415);
and U6441 (N_6441,N_3970,N_3233);
or U6442 (N_6442,N_3250,N_4170);
nand U6443 (N_6443,N_3062,N_3697);
nor U6444 (N_6444,N_5710,N_3085);
nand U6445 (N_6445,N_3453,N_3396);
xor U6446 (N_6446,N_4390,N_5822);
nor U6447 (N_6447,N_3105,N_5073);
xor U6448 (N_6448,N_3481,N_3296);
nor U6449 (N_6449,N_4025,N_5159);
and U6450 (N_6450,N_5375,N_4961);
and U6451 (N_6451,N_5032,N_5687);
nor U6452 (N_6452,N_4158,N_4861);
nor U6453 (N_6453,N_5681,N_3763);
and U6454 (N_6454,N_5505,N_4746);
nor U6455 (N_6455,N_5937,N_5390);
and U6456 (N_6456,N_5877,N_4954);
nand U6457 (N_6457,N_4238,N_4886);
xor U6458 (N_6458,N_4738,N_4867);
and U6459 (N_6459,N_3850,N_4624);
nor U6460 (N_6460,N_3743,N_4304);
nor U6461 (N_6461,N_5932,N_4938);
nand U6462 (N_6462,N_3615,N_4400);
nand U6463 (N_6463,N_5907,N_4584);
nor U6464 (N_6464,N_3513,N_5156);
nor U6465 (N_6465,N_5152,N_5737);
and U6466 (N_6466,N_3119,N_5906);
nand U6467 (N_6467,N_5615,N_5088);
nand U6468 (N_6468,N_3448,N_3302);
or U6469 (N_6469,N_5139,N_3527);
and U6470 (N_6470,N_4682,N_3301);
nand U6471 (N_6471,N_4758,N_5993);
or U6472 (N_6472,N_5378,N_4577);
nor U6473 (N_6473,N_3187,N_3719);
xor U6474 (N_6474,N_5749,N_5474);
or U6475 (N_6475,N_3999,N_3530);
or U6476 (N_6476,N_4112,N_4393);
nor U6477 (N_6477,N_5591,N_4329);
nor U6478 (N_6478,N_4652,N_3671);
nor U6479 (N_6479,N_3661,N_3804);
nor U6480 (N_6480,N_3215,N_5188);
nand U6481 (N_6481,N_5113,N_4848);
or U6482 (N_6482,N_3948,N_5004);
and U6483 (N_6483,N_5666,N_3135);
xnor U6484 (N_6484,N_4787,N_3006);
and U6485 (N_6485,N_5168,N_4880);
and U6486 (N_6486,N_3368,N_5081);
nand U6487 (N_6487,N_4323,N_5735);
xor U6488 (N_6488,N_4780,N_3209);
nor U6489 (N_6489,N_4033,N_3323);
xor U6490 (N_6490,N_3778,N_3148);
xnor U6491 (N_6491,N_3354,N_5942);
xnor U6492 (N_6492,N_3691,N_5493);
nor U6493 (N_6493,N_4145,N_4330);
xnor U6494 (N_6494,N_3279,N_3300);
or U6495 (N_6495,N_4929,N_4996);
xor U6496 (N_6496,N_4822,N_4220);
and U6497 (N_6497,N_5226,N_4365);
nand U6498 (N_6498,N_3353,N_3731);
or U6499 (N_6499,N_4063,N_4744);
nand U6500 (N_6500,N_5825,N_5012);
nand U6501 (N_6501,N_4988,N_4872);
or U6502 (N_6502,N_3990,N_5720);
nor U6503 (N_6503,N_3446,N_3326);
or U6504 (N_6504,N_3461,N_3032);
xnor U6505 (N_6505,N_4814,N_5231);
xor U6506 (N_6506,N_4545,N_5606);
nor U6507 (N_6507,N_3502,N_3303);
nor U6508 (N_6508,N_5229,N_5248);
nand U6509 (N_6509,N_4225,N_4337);
xor U6510 (N_6510,N_5023,N_4830);
and U6511 (N_6511,N_3580,N_3084);
and U6512 (N_6512,N_3428,N_3462);
and U6513 (N_6513,N_5381,N_4102);
nand U6514 (N_6514,N_3409,N_5968);
and U6515 (N_6515,N_3542,N_5394);
or U6516 (N_6516,N_5889,N_5764);
xor U6517 (N_6517,N_5502,N_4713);
nor U6518 (N_6518,N_3786,N_4017);
nor U6519 (N_6519,N_4066,N_3765);
xor U6520 (N_6520,N_5582,N_5564);
xnor U6521 (N_6521,N_5425,N_5046);
or U6522 (N_6522,N_3975,N_4421);
or U6523 (N_6523,N_4910,N_3389);
nor U6524 (N_6524,N_5745,N_3592);
xnor U6525 (N_6525,N_4219,N_3560);
nor U6526 (N_6526,N_4960,N_3101);
nor U6527 (N_6527,N_5385,N_4203);
xor U6528 (N_6528,N_4548,N_4021);
nor U6529 (N_6529,N_4808,N_5972);
xor U6530 (N_6530,N_4549,N_5428);
xor U6531 (N_6531,N_3210,N_4275);
and U6532 (N_6532,N_4789,N_5663);
nand U6533 (N_6533,N_5008,N_3315);
or U6534 (N_6534,N_5650,N_4571);
nand U6535 (N_6535,N_4523,N_3487);
xnor U6536 (N_6536,N_5852,N_5204);
and U6537 (N_6537,N_5694,N_5239);
nand U6538 (N_6538,N_3758,N_3247);
nand U6539 (N_6539,N_5507,N_3316);
xor U6540 (N_6540,N_5175,N_4286);
and U6541 (N_6541,N_5001,N_4653);
nand U6542 (N_6542,N_4543,N_5189);
and U6543 (N_6543,N_4864,N_5902);
nor U6544 (N_6544,N_4098,N_4661);
and U6545 (N_6545,N_5761,N_5292);
nand U6546 (N_6546,N_3750,N_4648);
nor U6547 (N_6547,N_4557,N_5660);
xnor U6548 (N_6548,N_5504,N_5025);
nor U6549 (N_6549,N_4424,N_5772);
and U6550 (N_6550,N_5085,N_5987);
and U6551 (N_6551,N_4198,N_5548);
or U6552 (N_6552,N_5068,N_5712);
nor U6553 (N_6553,N_5061,N_4041);
and U6554 (N_6554,N_3983,N_5991);
nand U6555 (N_6555,N_3589,N_4363);
and U6556 (N_6556,N_5442,N_4729);
and U6557 (N_6557,N_4273,N_5358);
nor U6558 (N_6558,N_3011,N_3835);
nand U6559 (N_6559,N_4974,N_5104);
or U6560 (N_6560,N_5368,N_4425);
nand U6561 (N_6561,N_4478,N_4670);
and U6562 (N_6562,N_5994,N_4208);
xnor U6563 (N_6563,N_3922,N_3532);
or U6564 (N_6564,N_5855,N_4242);
nand U6565 (N_6565,N_4472,N_5365);
and U6566 (N_6566,N_4427,N_5410);
xnor U6567 (N_6567,N_5520,N_5210);
nand U6568 (N_6568,N_4271,N_5067);
xnor U6569 (N_6569,N_4091,N_5466);
xnor U6570 (N_6570,N_4444,N_3078);
nand U6571 (N_6571,N_3884,N_4689);
nor U6572 (N_6572,N_3607,N_3971);
nand U6573 (N_6573,N_5322,N_3505);
and U6574 (N_6574,N_3293,N_3070);
or U6575 (N_6575,N_5490,N_5680);
nand U6576 (N_6576,N_4166,N_4833);
nor U6577 (N_6577,N_5572,N_3642);
or U6578 (N_6578,N_4572,N_3191);
xor U6579 (N_6579,N_5157,N_5729);
nand U6580 (N_6580,N_5870,N_3506);
or U6581 (N_6581,N_3364,N_3649);
nand U6582 (N_6582,N_4168,N_3640);
and U6583 (N_6583,N_4311,N_4412);
xnor U6584 (N_6584,N_3325,N_3145);
nand U6585 (N_6585,N_4121,N_4727);
xnor U6586 (N_6586,N_4701,N_4707);
xnor U6587 (N_6587,N_4012,N_5457);
or U6588 (N_6588,N_4408,N_3402);
nor U6589 (N_6589,N_5194,N_5069);
or U6590 (N_6590,N_3002,N_4181);
and U6591 (N_6591,N_3637,N_3658);
nor U6592 (N_6592,N_4451,N_5041);
nand U6593 (N_6593,N_4825,N_3793);
and U6594 (N_6594,N_4842,N_3365);
nor U6595 (N_6595,N_4907,N_4815);
xnor U6596 (N_6596,N_3471,N_4760);
nand U6597 (N_6597,N_3929,N_4728);
nor U6598 (N_6598,N_3582,N_5743);
nor U6599 (N_6599,N_4990,N_3897);
xnor U6600 (N_6600,N_5446,N_3033);
xnor U6601 (N_6601,N_3891,N_3489);
nand U6602 (N_6602,N_3894,N_4212);
and U6603 (N_6603,N_5817,N_4439);
or U6604 (N_6604,N_4546,N_3475);
nand U6605 (N_6605,N_4631,N_5843);
nand U6606 (N_6606,N_4837,N_5363);
or U6607 (N_6607,N_3966,N_5642);
xor U6608 (N_6608,N_5551,N_5594);
and U6609 (N_6609,N_3356,N_5166);
or U6610 (N_6610,N_4413,N_3160);
nand U6611 (N_6611,N_5170,N_5144);
nand U6612 (N_6612,N_4606,N_3504);
nand U6613 (N_6613,N_3890,N_5398);
or U6614 (N_6614,N_4551,N_3944);
or U6615 (N_6615,N_5543,N_3609);
nor U6616 (N_6616,N_5593,N_4176);
or U6617 (N_6617,N_4586,N_5356);
or U6618 (N_6618,N_5632,N_3412);
and U6619 (N_6619,N_3357,N_5475);
nand U6620 (N_6620,N_5522,N_5287);
and U6621 (N_6621,N_4908,N_5503);
and U6622 (N_6622,N_3598,N_4040);
and U6623 (N_6623,N_5316,N_3348);
nand U6624 (N_6624,N_5371,N_4228);
xnor U6625 (N_6625,N_5709,N_3162);
or U6626 (N_6626,N_4664,N_5765);
or U6627 (N_6627,N_4357,N_5043);
nand U6628 (N_6628,N_5380,N_3469);
xor U6629 (N_6629,N_3550,N_3346);
and U6630 (N_6630,N_3667,N_3901);
and U6631 (N_6631,N_4522,N_4865);
and U6632 (N_6632,N_4430,N_3692);
nor U6633 (N_6633,N_4118,N_4621);
xor U6634 (N_6634,N_3157,N_3910);
nand U6635 (N_6635,N_5277,N_3822);
and U6636 (N_6636,N_3953,N_3817);
nor U6637 (N_6637,N_3149,N_4935);
or U6638 (N_6638,N_4255,N_5300);
nand U6639 (N_6639,N_4933,N_5366);
xor U6640 (N_6640,N_4284,N_5060);
xnor U6641 (N_6641,N_4618,N_5999);
xnor U6642 (N_6642,N_4058,N_5847);
and U6643 (N_6643,N_3071,N_5234);
nor U6644 (N_6644,N_5814,N_3590);
and U6645 (N_6645,N_5109,N_5286);
nand U6646 (N_6646,N_4730,N_3985);
nand U6647 (N_6647,N_4646,N_5916);
and U6648 (N_6648,N_5279,N_4450);
or U6649 (N_6649,N_5886,N_4917);
xnor U6650 (N_6650,N_3962,N_5165);
xor U6651 (N_6651,N_4686,N_4554);
nand U6652 (N_6652,N_3488,N_3327);
and U6653 (N_6653,N_4695,N_3965);
and U6654 (N_6654,N_3103,N_3218);
xor U6655 (N_6655,N_5228,N_5627);
xnor U6656 (N_6656,N_3277,N_4923);
and U6657 (N_6657,N_5701,N_5858);
nor U6658 (N_6658,N_3583,N_5509);
nor U6659 (N_6659,N_4700,N_5555);
and U6660 (N_6660,N_3746,N_4005);
xnor U6661 (N_6661,N_4312,N_4204);
nor U6662 (N_6662,N_4479,N_5571);
nor U6663 (N_6663,N_4341,N_3497);
xor U6664 (N_6664,N_4930,N_5324);
xor U6665 (N_6665,N_5915,N_4616);
xor U6666 (N_6666,N_3723,N_4706);
nor U6667 (N_6667,N_3100,N_5535);
nand U6668 (N_6668,N_5670,N_5951);
or U6669 (N_6669,N_5964,N_4067);
nor U6670 (N_6670,N_5320,N_5449);
and U6671 (N_6671,N_5773,N_3407);
or U6672 (N_6672,N_4038,N_4481);
nor U6673 (N_6673,N_3367,N_4423);
nor U6674 (N_6674,N_5079,N_5690);
nor U6675 (N_6675,N_5637,N_3819);
nand U6676 (N_6676,N_4604,N_3427);
nand U6677 (N_6677,N_3611,N_3603);
or U6678 (N_6678,N_3166,N_3429);
nor U6679 (N_6679,N_5078,N_4257);
nand U6680 (N_6680,N_5982,N_5980);
nand U6681 (N_6681,N_5101,N_5795);
nor U6682 (N_6682,N_3436,N_3902);
xor U6683 (N_6683,N_3866,N_4500);
or U6684 (N_6684,N_5087,N_3915);
nor U6685 (N_6685,N_5064,N_4513);
and U6686 (N_6686,N_3058,N_3411);
nand U6687 (N_6687,N_4945,N_5383);
or U6688 (N_6688,N_5309,N_5386);
xor U6689 (N_6689,N_3474,N_3519);
or U6690 (N_6690,N_5361,N_5414);
or U6691 (N_6691,N_5010,N_3930);
nand U6692 (N_6692,N_3477,N_3359);
or U6693 (N_6693,N_3251,N_3618);
or U6694 (N_6694,N_3352,N_3904);
nor U6695 (N_6695,N_3438,N_5659);
or U6696 (N_6696,N_3845,N_3319);
and U6697 (N_6697,N_4587,N_4042);
and U6698 (N_6698,N_4716,N_3945);
or U6699 (N_6699,N_3252,N_3899);
xnor U6700 (N_6700,N_3163,N_4715);
nand U6701 (N_6701,N_3156,N_5589);
and U6702 (N_6702,N_3388,N_5218);
or U6703 (N_6703,N_5437,N_4338);
nand U6704 (N_6704,N_5598,N_3304);
xnor U6705 (N_6705,N_4027,N_4547);
and U6706 (N_6706,N_3403,N_3179);
nor U6707 (N_6707,N_4167,N_5975);
nand U6708 (N_6708,N_5575,N_4981);
or U6709 (N_6709,N_3702,N_5478);
nand U6710 (N_6710,N_3110,N_4262);
nand U6711 (N_6711,N_3559,N_4818);
xnor U6712 (N_6712,N_4644,N_3395);
xor U6713 (N_6713,N_3205,N_4628);
and U6714 (N_6714,N_3847,N_5240);
or U6715 (N_6715,N_3623,N_4681);
xor U6716 (N_6716,N_3479,N_4209);
nand U6717 (N_6717,N_3383,N_5177);
or U6718 (N_6718,N_4570,N_3833);
or U6719 (N_6719,N_4241,N_4519);
or U6720 (N_6720,N_5245,N_4657);
nor U6721 (N_6721,N_4740,N_3223);
and U6722 (N_6722,N_3645,N_3668);
or U6723 (N_6723,N_5219,N_5945);
xor U6724 (N_6724,N_3805,N_5608);
nand U6725 (N_6725,N_5959,N_4737);
and U6726 (N_6726,N_3619,N_3167);
or U6727 (N_6727,N_5281,N_4821);
nand U6728 (N_6728,N_5801,N_5554);
or U6729 (N_6729,N_5804,N_3013);
nor U6730 (N_6730,N_5753,N_4092);
and U6731 (N_6731,N_3699,N_3212);
nand U6732 (N_6732,N_4199,N_3230);
or U6733 (N_6733,N_3116,N_3268);
xor U6734 (N_6734,N_3241,N_4702);
nor U6735 (N_6735,N_3090,N_5142);
or U6736 (N_6736,N_5341,N_4969);
xnor U6737 (N_6737,N_4399,N_4947);
xnor U6738 (N_6738,N_5222,N_4800);
nor U6739 (N_6739,N_4326,N_5002);
and U6740 (N_6740,N_4061,N_5102);
or U6741 (N_6741,N_5404,N_3236);
or U6742 (N_6742,N_3400,N_5402);
nand U6743 (N_6743,N_4882,N_3827);
nand U6744 (N_6744,N_4555,N_3107);
and U6745 (N_6745,N_4985,N_4149);
and U6746 (N_6746,N_4953,N_3873);
nand U6747 (N_6747,N_4633,N_4951);
or U6748 (N_6748,N_4544,N_5353);
and U6749 (N_6749,N_5918,N_4231);
nand U6750 (N_6750,N_4410,N_5203);
nor U6751 (N_6751,N_5950,N_5274);
nor U6752 (N_6752,N_3151,N_4832);
and U6753 (N_6753,N_4401,N_4995);
xor U6754 (N_6754,N_4144,N_3662);
or U6755 (N_6755,N_3955,N_5271);
xnor U6756 (N_6756,N_4004,N_3072);
nand U6757 (N_6757,N_5464,N_5639);
and U6758 (N_6758,N_5283,N_4692);
and U6759 (N_6759,N_5568,N_5225);
nand U6760 (N_6760,N_4177,N_3972);
nand U6761 (N_6761,N_5617,N_4369);
and U6762 (N_6762,N_3780,N_5408);
nor U6763 (N_6763,N_5117,N_5647);
and U6764 (N_6764,N_4920,N_4200);
or U6765 (N_6765,N_4082,N_3518);
xor U6766 (N_6766,N_5153,N_3614);
xor U6767 (N_6767,N_4081,N_3688);
or U6768 (N_6768,N_5721,N_3627);
and U6769 (N_6769,N_4565,N_3551);
and U6770 (N_6770,N_4246,N_4321);
nor U6771 (N_6771,N_4354,N_5662);
xor U6772 (N_6772,N_5570,N_5454);
or U6773 (N_6773,N_4088,N_5112);
nor U6774 (N_6774,N_3246,N_5940);
or U6775 (N_6775,N_3183,N_5296);
and U6776 (N_6776,N_5401,N_4620);
nor U6777 (N_6777,N_3555,N_4110);
or U6778 (N_6778,N_5327,N_4124);
or U6779 (N_6779,N_3457,N_4524);
or U6780 (N_6780,N_3274,N_3740);
nand U6781 (N_6781,N_4322,N_4845);
or U6782 (N_6782,N_3605,N_4064);
nor U6783 (N_6783,N_4274,N_4371);
and U6784 (N_6784,N_4763,N_4937);
or U6785 (N_6785,N_3102,N_5866);
or U6786 (N_6786,N_4912,N_4043);
or U6787 (N_6787,N_3060,N_3450);
or U6788 (N_6788,N_4876,N_5785);
and U6789 (N_6789,N_3035,N_4313);
xor U6790 (N_6790,N_5626,N_5372);
nand U6791 (N_6791,N_3076,N_4512);
nand U6792 (N_6792,N_5491,N_4296);
xnor U6793 (N_6793,N_3138,N_4694);
nor U6794 (N_6794,N_4788,N_5145);
and U6795 (N_6795,N_5174,N_5123);
nor U6796 (N_6796,N_3404,N_3549);
and U6797 (N_6797,N_3122,N_5416);
xor U6798 (N_6798,N_5684,N_4532);
nand U6799 (N_6799,N_4658,N_3730);
and U6800 (N_6800,N_4632,N_3312);
or U6801 (N_6801,N_4154,N_3445);
and U6802 (N_6802,N_3372,N_5106);
xnor U6803 (N_6803,N_3785,N_5933);
or U6804 (N_6804,N_3114,N_3442);
nor U6805 (N_6805,N_3083,N_5434);
and U6806 (N_6806,N_5809,N_3680);
and U6807 (N_6807,N_3426,N_5584);
nor U6808 (N_6808,N_3144,N_3987);
or U6809 (N_6809,N_5971,N_5821);
nor U6810 (N_6810,N_3027,N_4404);
or U6811 (N_6811,N_3055,N_5727);
xnor U6812 (N_6812,N_4001,N_5498);
xnor U6813 (N_6813,N_4802,N_4743);
nand U6814 (N_6814,N_5596,N_5103);
nand U6815 (N_6815,N_4762,N_3184);
and U6816 (N_6816,N_5920,N_5276);
xor U6817 (N_6817,N_5678,N_5133);
and U6818 (N_6818,N_3969,N_5901);
or U6819 (N_6819,N_4795,N_5492);
or U6820 (N_6820,N_3814,N_4964);
or U6821 (N_6821,N_5237,N_5759);
nor U6822 (N_6822,N_4134,N_4141);
or U6823 (N_6823,N_4659,N_5389);
nor U6824 (N_6824,N_4783,N_4645);
and U6825 (N_6825,N_4801,N_3343);
or U6826 (N_6826,N_4377,N_4894);
or U6827 (N_6827,N_5172,N_3467);
or U6828 (N_6828,N_4372,N_4175);
nand U6829 (N_6829,N_5740,N_5897);
and U6830 (N_6830,N_4469,N_4483);
xor U6831 (N_6831,N_5969,N_5459);
and U6832 (N_6832,N_5039,N_4809);
or U6833 (N_6833,N_4153,N_3178);
xnor U6834 (N_6834,N_4407,N_3460);
nand U6835 (N_6835,N_5692,N_5835);
nand U6836 (N_6836,N_4136,N_3602);
or U6837 (N_6837,N_3322,N_4642);
xnor U6838 (N_6838,N_3566,N_5703);
nor U6839 (N_6839,N_4272,N_4982);
and U6840 (N_6840,N_5777,N_3106);
or U6841 (N_6841,N_3243,N_5313);
and U6842 (N_6842,N_3271,N_3213);
nor U6843 (N_6843,N_5333,N_3036);
and U6844 (N_6844,N_5622,N_3565);
and U6845 (N_6845,N_4194,N_3345);
xnor U6846 (N_6846,N_3028,N_5472);
nand U6847 (N_6847,N_3313,N_5045);
nand U6848 (N_6848,N_5302,N_3441);
or U6849 (N_6849,N_4761,N_5635);
nand U6850 (N_6850,N_3515,N_3920);
nor U6851 (N_6851,N_3449,N_4559);
and U6852 (N_6852,N_5839,N_5301);
nor U6853 (N_6853,N_4215,N_5307);
nand U6854 (N_6854,N_4352,N_3498);
xor U6855 (N_6855,N_4950,N_5354);
xnor U6856 (N_6856,N_3088,N_4846);
xor U6857 (N_6857,N_5456,N_4047);
or U6858 (N_6858,N_3713,N_4108);
or U6859 (N_6859,N_4129,N_3065);
xnor U6860 (N_6860,N_5049,N_3575);
and U6861 (N_6861,N_5108,N_3508);
nand U6862 (N_6862,N_4687,N_4159);
nand U6863 (N_6863,N_3783,N_5419);
nand U6864 (N_6864,N_5370,N_4462);
nor U6865 (N_6865,N_3385,N_3393);
nand U6866 (N_6866,N_5040,N_4062);
nand U6867 (N_6867,N_4492,N_5881);
and U6868 (N_6868,N_5130,N_3993);
xor U6869 (N_6869,N_3973,N_5196);
xor U6870 (N_6870,N_5526,N_5282);
nor U6871 (N_6871,N_4288,N_5557);
and U6872 (N_6872,N_3829,N_4368);
and U6873 (N_6873,N_5754,N_5952);
xnor U6874 (N_6874,N_3792,N_3545);
or U6875 (N_6875,N_3736,N_3482);
xnor U6876 (N_6876,N_5943,N_5388);
and U6877 (N_6877,N_4328,N_3452);
nor U6878 (N_6878,N_3073,N_4016);
and U6879 (N_6879,N_3175,N_5513);
nand U6880 (N_6880,N_4599,N_4087);
nor U6881 (N_6881,N_3751,N_5580);
or U6882 (N_6882,N_3874,N_3374);
xnor U6883 (N_6883,N_4989,N_3111);
nor U6884 (N_6884,N_3007,N_3344);
xnor U6885 (N_6885,N_5426,N_3745);
or U6886 (N_6886,N_5707,N_5424);
xnor U6887 (N_6887,N_3042,N_3544);
nand U6888 (N_6888,N_4403,N_3610);
and U6889 (N_6889,N_5673,N_3423);
and U6890 (N_6890,N_3408,N_4432);
or U6891 (N_6891,N_4143,N_3943);
xor U6892 (N_6892,N_5601,N_3905);
nor U6893 (N_6893,N_4535,N_4336);
or U6894 (N_6894,N_3594,N_4827);
nor U6895 (N_6895,N_3612,N_3161);
nand U6896 (N_6896,N_3134,N_5774);
or U6897 (N_6897,N_3823,N_5815);
nand U6898 (N_6898,N_5290,N_3067);
nor U6899 (N_6899,N_5756,N_3196);
nand U6900 (N_6900,N_4054,N_4011);
nor U6901 (N_6901,N_4428,N_5284);
xnor U6902 (N_6902,N_4236,N_4260);
and U6903 (N_6903,N_4216,N_3756);
xnor U6904 (N_6904,N_4810,N_4431);
or U6905 (N_6905,N_5487,N_3927);
and U6906 (N_6906,N_5392,N_5697);
xor U6907 (N_6907,N_4578,N_3264);
nand U6908 (N_6908,N_3249,N_5243);
or U6909 (N_6909,N_5141,N_3934);
and U6910 (N_6910,N_5197,N_4250);
xnor U6911 (N_6911,N_4409,N_4866);
nand U6912 (N_6912,N_3473,N_4915);
nand U6913 (N_6913,N_5726,N_4084);
nor U6914 (N_6914,N_5998,N_4796);
nand U6915 (N_6915,N_5376,N_3188);
nor U6916 (N_6916,N_3164,N_5421);
or U6917 (N_6917,N_4002,N_4733);
or U6918 (N_6918,N_5644,N_5255);
and U6919 (N_6919,N_3558,N_3715);
or U6920 (N_6920,N_4709,N_4588);
nor U6921 (N_6921,N_3660,N_5914);
and U6922 (N_6922,N_3222,N_3735);
or U6923 (N_6923,N_3398,N_3221);
or U6924 (N_6924,N_5011,N_3405);
or U6925 (N_6925,N_4493,N_4916);
nand U6926 (N_6926,N_3777,N_3371);
nor U6927 (N_6927,N_4292,N_4083);
or U6928 (N_6928,N_5241,N_5714);
and U6929 (N_6929,N_5592,N_4448);
nand U6930 (N_6930,N_5711,N_3130);
xor U6931 (N_6931,N_5890,N_3127);
xnor U6932 (N_6932,N_3821,N_5515);
xor U6933 (N_6933,N_5223,N_5155);
xnor U6934 (N_6934,N_3666,N_3349);
xnor U6935 (N_6935,N_5345,N_3056);
and U6936 (N_6936,N_3789,N_4270);
and U6937 (N_6937,N_3137,N_3521);
xnor U6938 (N_6938,N_5854,N_5467);
and U6939 (N_6939,N_3561,N_4488);
or U6940 (N_6940,N_5587,N_4282);
nand U6941 (N_6941,N_4173,N_5799);
nand U6942 (N_6942,N_4295,N_4300);
nor U6943 (N_6943,N_4765,N_4781);
xnor U6944 (N_6944,N_5288,N_5844);
and U6945 (N_6945,N_3514,N_4875);
nand U6946 (N_6946,N_5486,N_4484);
nor U6947 (N_6947,N_3533,N_3496);
or U6948 (N_6948,N_4779,N_4305);
xor U6949 (N_6949,N_3172,N_3439);
nor U6950 (N_6950,N_4267,N_5521);
or U6951 (N_6951,N_3309,N_4151);
and U6952 (N_6952,N_4473,N_5154);
nand U6953 (N_6953,N_4790,N_4601);
or U6954 (N_6954,N_3848,N_5880);
or U6955 (N_6955,N_5788,N_4840);
nand U6956 (N_6956,N_3917,N_3587);
or U6957 (N_6957,N_4114,N_3727);
and U6958 (N_6958,N_4165,N_4508);
nor U6959 (N_6959,N_4665,N_3141);
nand U6960 (N_6960,N_4719,N_5699);
or U6961 (N_6961,N_4573,N_4384);
nand U6962 (N_6962,N_3143,N_4841);
nor U6963 (N_6963,N_5485,N_4069);
and U6964 (N_6964,N_3297,N_3936);
nor U6965 (N_6965,N_5098,N_5310);
and U6966 (N_6966,N_3764,N_3080);
and U6967 (N_6967,N_3951,N_4870);
and U6968 (N_6968,N_3000,N_5923);
nand U6969 (N_6969,N_4094,N_5523);
nor U6970 (N_6970,N_4854,N_5399);
xnor U6971 (N_6971,N_5739,N_3516);
nor U6972 (N_6972,N_4489,N_4596);
nor U6973 (N_6973,N_4217,N_5693);
nor U6974 (N_6974,N_3841,N_4775);
nand U6975 (N_6975,N_5254,N_3808);
nand U6976 (N_6976,N_5992,N_5905);
nor U6977 (N_6977,N_5831,N_4622);
xor U6978 (N_6978,N_5860,N_3284);
nor U6979 (N_6979,N_3199,N_3959);
nand U6980 (N_6980,N_4192,N_4174);
and U6981 (N_6981,N_3043,N_3826);
xor U6982 (N_6982,N_4824,N_5652);
or U6983 (N_6983,N_5395,N_5494);
nand U6984 (N_6984,N_5373,N_5946);
nand U6985 (N_6985,N_3562,N_4477);
nor U6986 (N_6986,N_3893,N_5696);
xnor U6987 (N_6987,N_3846,N_4638);
nor U6988 (N_6988,N_5347,N_3455);
and U6989 (N_6989,N_3863,N_4491);
nand U6990 (N_6990,N_5114,N_5352);
or U6991 (N_6991,N_4358,N_4590);
or U6992 (N_6992,N_5235,N_5544);
nand U6993 (N_6993,N_5193,N_3420);
nand U6994 (N_6994,N_3978,N_5211);
and U6995 (N_6995,N_4239,N_3617);
nand U6996 (N_6996,N_5541,N_5935);
nor U6997 (N_6997,N_3725,N_3378);
and U6998 (N_6998,N_3492,N_4183);
nor U6999 (N_6999,N_3577,N_4052);
xor U7000 (N_7000,N_5350,N_5829);
xor U7001 (N_7001,N_5413,N_5263);
nand U7002 (N_7002,N_4452,N_5529);
nor U7003 (N_7003,N_4504,N_5289);
xor U7004 (N_7004,N_5850,N_4014);
and U7005 (N_7005,N_3394,N_3125);
and U7006 (N_7006,N_4792,N_3775);
nand U7007 (N_7007,N_4767,N_5634);
or U7008 (N_7008,N_4475,N_4823);
and U7009 (N_7009,N_4580,N_5863);
and U7010 (N_7010,N_3216,N_5403);
xor U7011 (N_7011,N_4726,N_4514);
or U7012 (N_7012,N_3081,N_3280);
nor U7013 (N_7013,N_5021,N_5718);
xor U7014 (N_7014,N_5094,N_4223);
nand U7015 (N_7015,N_3864,N_3075);
nor U7016 (N_7016,N_4315,N_3570);
and U7017 (N_7017,N_4839,N_4090);
nand U7018 (N_7018,N_3478,N_3578);
nor U7019 (N_7019,N_4521,N_4674);
nor U7020 (N_7020,N_5026,N_4793);
xor U7021 (N_7021,N_4952,N_3443);
xor U7022 (N_7022,N_3790,N_3772);
nor U7023 (N_7023,N_3086,N_3009);
nor U7024 (N_7024,N_5636,N_4335);
xnor U7025 (N_7025,N_4946,N_4647);
xnor U7026 (N_7026,N_4029,N_5887);
or U7027 (N_7027,N_4139,N_5397);
xor U7028 (N_7028,N_3413,N_4317);
or U7029 (N_7029,N_4820,N_4024);
nor U7030 (N_7030,N_5602,N_4986);
nor U7031 (N_7031,N_4155,N_5460);
or U7032 (N_7032,N_3665,N_3643);
nand U7033 (N_7033,N_4858,N_5830);
nand U7034 (N_7034,N_5136,N_3108);
nor U7035 (N_7035,N_4979,N_4871);
xor U7036 (N_7036,N_4776,N_5438);
nand U7037 (N_7037,N_4076,N_4362);
and U7038 (N_7038,N_3089,N_5939);
nor U7039 (N_7039,N_5824,N_4721);
and U7040 (N_7040,N_5264,N_3912);
xor U7041 (N_7041,N_4678,N_5840);
and U7042 (N_7042,N_5480,N_3710);
and U7043 (N_7043,N_3997,N_5682);
and U7044 (N_7044,N_3721,N_3942);
nor U7045 (N_7045,N_5676,N_4718);
xor U7046 (N_7046,N_5455,N_3093);
nor U7047 (N_7047,N_3779,N_4051);
xnor U7048 (N_7048,N_4966,N_5208);
nor U7049 (N_7049,N_4386,N_5070);
nand U7050 (N_7050,N_3656,N_5178);
xor U7051 (N_7051,N_3854,N_5781);
nand U7052 (N_7052,N_3995,N_5044);
or U7053 (N_7053,N_3169,N_3747);
and U7054 (N_7054,N_4878,N_3885);
nor U7055 (N_7055,N_4132,N_5766);
xnor U7056 (N_7056,N_3379,N_5985);
and U7057 (N_7057,N_3685,N_5256);
nor U7058 (N_7058,N_4180,N_4471);
or U7059 (N_7059,N_3290,N_4940);
xor U7060 (N_7060,N_4283,N_3968);
and U7061 (N_7061,N_5299,N_3046);
xor U7062 (N_7062,N_4569,N_5931);
xnor U7063 (N_7063,N_5656,N_5473);
and U7064 (N_7064,N_3120,N_4955);
and U7065 (N_7065,N_5232,N_4397);
nand U7066 (N_7066,N_5430,N_3239);
and U7067 (N_7067,N_4748,N_3674);
nor U7068 (N_7068,N_3476,N_3008);
xor U7069 (N_7069,N_3259,N_5633);
and U7070 (N_7070,N_5140,N_4855);
and U7071 (N_7071,N_3299,N_3406);
nor U7072 (N_7072,N_5780,N_4526);
nor U7073 (N_7073,N_5762,N_4293);
nor U7074 (N_7074,N_3853,N_3635);
nand U7075 (N_7075,N_5818,N_4359);
and U7076 (N_7076,N_4186,N_4325);
xnor U7077 (N_7077,N_5595,N_3724);
nor U7078 (N_7078,N_4531,N_5838);
xnor U7079 (N_7079,N_5990,N_4527);
xnor U7080 (N_7080,N_5415,N_5948);
nor U7081 (N_7081,N_5778,N_5257);
and U7082 (N_7082,N_4625,N_3421);
xnor U7083 (N_7083,N_3717,N_3538);
and U7084 (N_7084,N_4125,N_4073);
and U7085 (N_7085,N_5252,N_3520);
and U7086 (N_7086,N_5770,N_5763);
xnor U7087 (N_7087,N_5272,N_3906);
nand U7088 (N_7088,N_5192,N_4085);
or U7089 (N_7089,N_5683,N_5134);
xnor U7090 (N_7090,N_3842,N_5471);
nand U7091 (N_7091,N_3480,N_3918);
and U7092 (N_7092,N_3782,N_3706);
and U7093 (N_7093,N_4703,N_5126);
or U7094 (N_7094,N_3192,N_5297);
or U7095 (N_7095,N_5832,N_4696);
or U7096 (N_7096,N_5654,N_5267);
xnor U7097 (N_7097,N_4162,N_3976);
nor U7098 (N_7098,N_5065,N_5185);
xor U7099 (N_7099,N_3682,N_3463);
nor U7100 (N_7100,N_5653,N_4723);
nand U7101 (N_7101,N_4123,N_4529);
nor U7102 (N_7102,N_3276,N_4868);
nand U7103 (N_7103,N_4948,N_3255);
nor U7104 (N_7104,N_5176,N_5072);
and U7105 (N_7105,N_4230,N_4847);
xor U7106 (N_7106,N_3207,N_5236);
nor U7107 (N_7107,N_5200,N_5516);
xor U7108 (N_7108,N_3916,N_3150);
xnor U7109 (N_7109,N_4736,N_3307);
nor U7110 (N_7110,N_5755,N_5084);
and U7111 (N_7111,N_4191,N_5792);
xnor U7112 (N_7112,N_5524,N_4113);
nor U7113 (N_7113,N_4277,N_5326);
nand U7114 (N_7114,N_4836,N_4171);
and U7115 (N_7115,N_3852,N_3800);
nor U7116 (N_7116,N_3709,N_5605);
nor U7117 (N_7117,N_5167,N_5148);
nor U7118 (N_7118,N_3613,N_5628);
xor U7119 (N_7119,N_5790,N_4320);
and U7120 (N_7120,N_5339,N_3714);
and U7121 (N_7121,N_4056,N_3272);
xor U7122 (N_7122,N_4654,N_5258);
or U7123 (N_7123,N_3317,N_3742);
xnor U7124 (N_7124,N_3526,N_4921);
and U7125 (N_7125,N_3235,N_5848);
nor U7126 (N_7126,N_3330,N_3654);
or U7127 (N_7127,N_5107,N_3201);
or U7128 (N_7128,N_4926,N_4263);
or U7129 (N_7129,N_5715,N_4934);
xnor U7130 (N_7130,N_3857,N_4503);
xnor U7131 (N_7131,N_5730,N_3856);
or U7132 (N_7132,N_5482,N_3048);
and U7133 (N_7133,N_5869,N_3974);
xnor U7134 (N_7134,N_3872,N_4131);
and U7135 (N_7135,N_3288,N_3136);
nor U7136 (N_7136,N_4105,N_3257);
nor U7137 (N_7137,N_5250,N_4031);
or U7138 (N_7138,N_5294,N_4314);
nor U7139 (N_7139,N_4497,N_5624);
nand U7140 (N_7140,N_4006,N_4046);
and U7141 (N_7141,N_5357,N_5586);
xor U7142 (N_7142,N_5953,N_3556);
xnor U7143 (N_7143,N_5623,N_3051);
and U7144 (N_7144,N_4034,N_4829);
or U7145 (N_7145,N_3380,N_4968);
nor U7146 (N_7146,N_4375,N_3459);
and U7147 (N_7147,N_5828,N_3240);
xnor U7148 (N_7148,N_4566,N_3858);
xnor U7149 (N_7149,N_4146,N_3173);
nor U7150 (N_7150,N_3676,N_4285);
nor U7151 (N_7151,N_4261,N_5936);
nand U7152 (N_7152,N_3324,N_3286);
xnor U7153 (N_7153,N_5201,N_5649);
or U7154 (N_7154,N_4924,N_5343);
nand U7155 (N_7155,N_5295,N_3599);
nand U7156 (N_7156,N_4859,N_4927);
and U7157 (N_7157,N_3171,N_4309);
or U7158 (N_7158,N_4243,N_4070);
nor U7159 (N_7159,N_5552,N_4888);
nand U7160 (N_7160,N_4420,N_3417);
xor U7161 (N_7161,N_3091,N_4157);
and U7162 (N_7162,N_4896,N_3355);
and U7163 (N_7163,N_4515,N_5066);
nand U7164 (N_7164,N_4943,N_4474);
xor U7165 (N_7165,N_5820,N_3784);
nand U7166 (N_7166,N_3900,N_3919);
xnor U7167 (N_7167,N_3234,N_5604);
xor U7168 (N_7168,N_4079,N_5533);
and U7169 (N_7169,N_4574,N_4348);
or U7170 (N_7170,N_5603,N_3812);
nand U7171 (N_7171,N_3875,N_3531);
and U7172 (N_7172,N_5120,N_3761);
or U7173 (N_7173,N_5116,N_5205);
xnor U7174 (N_7174,N_4655,N_4048);
nand U7175 (N_7175,N_4834,N_3629);
nor U7176 (N_7176,N_5784,N_3026);
nor U7177 (N_7177,N_5574,N_4607);
nand U7178 (N_7178,N_4994,N_4391);
nand U7179 (N_7179,N_5435,N_4258);
or U7180 (N_7180,N_4812,N_4817);
nand U7181 (N_7181,N_4018,N_4294);
and U7182 (N_7182,N_4107,N_3197);
xor U7183 (N_7183,N_4028,N_4429);
nand U7184 (N_7184,N_4931,N_5531);
or U7185 (N_7185,N_5216,N_5986);
nand U7186 (N_7186,N_5163,N_4499);
xor U7187 (N_7187,N_4879,N_4562);
nor U7188 (N_7188,N_5311,N_5895);
and U7189 (N_7189,N_5348,N_3698);
or U7190 (N_7190,N_4782,N_5453);
and U7191 (N_7191,N_3522,N_4234);
xor U7192 (N_7192,N_5137,N_3703);
xor U7193 (N_7193,N_4813,N_3375);
nand U7194 (N_7194,N_3037,N_3991);
or U7195 (N_7195,N_3363,N_4764);
xnor U7196 (N_7196,N_5954,N_5949);
xnor U7197 (N_7197,N_3898,N_4676);
or U7198 (N_7198,N_5900,N_4213);
nor U7199 (N_7199,N_5082,N_3621);
or U7200 (N_7200,N_4887,N_3576);
and U7201 (N_7201,N_5450,N_3232);
nand U7202 (N_7202,N_5213,N_3104);
and U7203 (N_7203,N_5562,N_4560);
or U7204 (N_7204,N_3650,N_4036);
nor U7205 (N_7205,N_4278,N_5970);
nand U7206 (N_7206,N_4074,N_3029);
nand U7207 (N_7207,N_4161,N_5391);
or U7208 (N_7208,N_3718,N_5029);
or U7209 (N_7209,N_3753,N_3200);
nor U7210 (N_7210,N_4344,N_4366);
nand U7211 (N_7211,N_5638,N_3887);
nor U7212 (N_7212,N_3509,N_5330);
and U7213 (N_7213,N_5005,N_4128);
xnor U7214 (N_7214,N_4256,N_3967);
or U7215 (N_7215,N_3737,N_3529);
nand U7216 (N_7216,N_3174,N_5077);
xor U7217 (N_7217,N_5569,N_3952);
xor U7218 (N_7218,N_4901,N_3170);
or U7219 (N_7219,N_3937,N_3687);
and U7220 (N_7220,N_5337,N_5242);
xnor U7221 (N_7221,N_4264,N_4142);
nand U7222 (N_7222,N_4685,N_5135);
or U7223 (N_7223,N_3655,N_4668);
nor U7224 (N_7224,N_4735,N_5910);
or U7225 (N_7225,N_4553,N_3572);
nor U7226 (N_7226,N_4418,N_3895);
and U7227 (N_7227,N_4619,N_3749);
nor U7228 (N_7228,N_4280,N_5981);
nand U7229 (N_7229,N_4597,N_5769);
nor U7230 (N_7230,N_4967,N_3788);
xor U7231 (N_7231,N_5003,N_3729);
xnor U7232 (N_7232,N_3057,N_5856);
and U7233 (N_7233,N_3888,N_5849);
and U7234 (N_7234,N_5443,N_4414);
nor U7235 (N_7235,N_4248,N_3298);
xor U7236 (N_7236,N_4978,N_4218);
or U7237 (N_7237,N_5661,N_5308);
nand U7238 (N_7238,N_3311,N_3020);
and U7239 (N_7239,N_3063,N_5896);
nand U7240 (N_7240,N_4911,N_4251);
xnor U7241 (N_7241,N_3924,N_4201);
xor U7242 (N_7242,N_5842,N_3690);
nor U7243 (N_7243,N_3258,N_4019);
xnor U7244 (N_7244,N_3926,N_5083);
or U7245 (N_7245,N_3696,N_5657);
xor U7246 (N_7246,N_3003,N_5259);
nand U7247 (N_7247,N_5705,N_4777);
nor U7248 (N_7248,N_3129,N_4389);
and U7249 (N_7249,N_4435,N_5090);
xor U7250 (N_7250,N_4613,N_3794);
nand U7251 (N_7251,N_3066,N_3338);
xnor U7252 (N_7252,N_3109,N_3557);
and U7253 (N_7253,N_5786,N_5118);
xnor U7254 (N_7254,N_4991,N_4518);
nor U7255 (N_7255,N_5836,N_3472);
nor U7256 (N_7256,N_4148,N_4195);
or U7257 (N_7257,N_5546,N_4268);
nand U7258 (N_7258,N_5874,N_4691);
nand U7259 (N_7259,N_5614,N_3754);
or U7260 (N_7260,N_3689,N_5713);
nand U7261 (N_7261,N_3465,N_4957);
and U7262 (N_7262,N_3376,N_3082);
nor U7263 (N_7263,N_5319,N_4992);
and U7264 (N_7264,N_3935,N_5810);
nand U7265 (N_7265,N_5499,N_3851);
nand U7266 (N_7266,N_4749,N_3014);
nand U7267 (N_7267,N_5884,N_3708);
nand U7268 (N_7268,N_4044,N_5215);
xnor U7269 (N_7269,N_3275,N_3722);
and U7270 (N_7270,N_4629,N_5075);
or U7271 (N_7271,N_4898,N_5908);
xnor U7272 (N_7272,N_3328,N_3537);
xnor U7273 (N_7273,N_4885,N_3244);
nand U7274 (N_7274,N_4334,N_4826);
nand U7275 (N_7275,N_3525,N_3414);
nor U7276 (N_7276,N_5648,N_3554);
nor U7277 (N_7277,N_5588,N_4383);
xor U7278 (N_7278,N_4773,N_4289);
or U7279 (N_7279,N_4080,N_5834);
xnor U7280 (N_7280,N_5036,N_4436);
xor U7281 (N_7281,N_5609,N_5560);
or U7282 (N_7282,N_4182,N_3932);
and U7283 (N_7283,N_3340,N_5700);
or U7284 (N_7284,N_4528,N_3881);
or U7285 (N_7285,N_4077,N_4956);
nand U7286 (N_7286,N_3907,N_5827);
nor U7287 (N_7287,N_3766,N_4306);
nor U7288 (N_7288,N_5984,N_5807);
nand U7289 (N_7289,N_5899,N_5017);
nor U7290 (N_7290,N_4770,N_5540);
and U7291 (N_7291,N_3726,N_4711);
xor U7292 (N_7292,N_5183,N_4897);
nand U7293 (N_7293,N_3391,N_5677);
nor U7294 (N_7294,N_5775,N_3310);
and U7295 (N_7295,N_4030,N_4206);
nor U7296 (N_7296,N_4343,N_5362);
nor U7297 (N_7297,N_3159,N_4269);
nand U7298 (N_7298,N_5873,N_5179);
nand U7299 (N_7299,N_5186,N_3646);
or U7300 (N_7300,N_5518,N_5876);
xor U7301 (N_7301,N_4259,N_5583);
or U7302 (N_7302,N_4592,N_3217);
xnor U7303 (N_7303,N_4032,N_3273);
or U7304 (N_7304,N_4466,N_4993);
or U7305 (N_7305,N_4302,N_5878);
nor U7306 (N_7306,N_3018,N_3762);
nand U7307 (N_7307,N_5733,N_3996);
and U7308 (N_7308,N_3242,N_4626);
or U7309 (N_7309,N_4563,N_5782);
xnor U7310 (N_7310,N_4747,N_3701);
nand U7311 (N_7311,N_4290,N_4725);
and U7312 (N_7312,N_5511,N_5037);
or U7313 (N_7313,N_3652,N_3540);
and U7314 (N_7314,N_3501,N_3569);
nor U7315 (N_7315,N_3418,N_3198);
nand U7316 (N_7316,N_4476,N_5960);
nand U7317 (N_7317,N_3064,N_4677);
or U7318 (N_7318,N_3744,N_3203);
nand U7319 (N_7319,N_4120,N_4301);
nor U7320 (N_7320,N_5796,N_3543);
nor U7321 (N_7321,N_5014,N_4459);
nor U7322 (N_7322,N_5369,N_3681);
or U7323 (N_7323,N_5867,N_5530);
nand U7324 (N_7324,N_5169,N_5050);
and U7325 (N_7325,N_3267,N_4567);
nand U7326 (N_7326,N_3485,N_4179);
nand U7327 (N_7327,N_5664,N_4370);
and U7328 (N_7328,N_3113,N_5802);
nor U7329 (N_7329,N_4331,N_4490);
and U7330 (N_7330,N_4970,N_3484);
and U7331 (N_7331,N_3416,N_4517);
nand U7332 (N_7332,N_4075,N_3546);
and U7333 (N_7333,N_5387,N_5227);
nand U7334 (N_7334,N_5076,N_3634);
or U7335 (N_7335,N_5110,N_5062);
xor U7336 (N_7336,N_3511,N_4983);
nand U7337 (N_7337,N_3261,N_5190);
nor U7338 (N_7338,N_4742,N_4433);
xor U7339 (N_7339,N_3399,N_3958);
xor U7340 (N_7340,N_3074,N_5671);
xnor U7341 (N_7341,N_3500,N_5955);
xor U7342 (N_7342,N_3831,N_5573);
and U7343 (N_7343,N_3908,N_5162);
nand U7344 (N_7344,N_4360,N_3998);
nand U7345 (N_7345,N_3260,N_5495);
nand U7346 (N_7346,N_5305,N_4525);
nor U7347 (N_7347,N_3774,N_4731);
xnor U7348 (N_7348,N_3700,N_4402);
xor U7349 (N_7349,N_4441,N_5317);
nand U7350 (N_7350,N_5018,N_5342);
xor U7351 (N_7351,N_4188,N_4009);
and U7352 (N_7352,N_4640,N_4351);
xor U7353 (N_7353,N_3017,N_3329);
and U7354 (N_7354,N_5099,N_3595);
nor U7355 (N_7355,N_4708,N_4207);
nand U7356 (N_7356,N_4340,N_5160);
nor U7357 (N_7357,N_5640,N_4455);
and U7358 (N_7358,N_5646,N_5006);
or U7359 (N_7359,N_5783,N_4350);
xnor U7360 (N_7360,N_3639,N_4705);
and U7361 (N_7361,N_3992,N_4010);
nand U7362 (N_7362,N_4447,N_5033);
nand U7363 (N_7363,N_3791,N_5293);
nor U7364 (N_7364,N_3670,N_3185);
or U7365 (N_7365,N_5837,N_3651);
nand U7366 (N_7366,N_3435,N_3370);
and U7367 (N_7367,N_4059,N_5995);
or U7368 (N_7368,N_3956,N_3769);
nor U7369 (N_7369,N_3341,N_4169);
xor U7370 (N_7370,N_5071,N_3938);
and U7371 (N_7371,N_4237,N_5074);
xor U7372 (N_7372,N_3659,N_4630);
nand U7373 (N_7373,N_5220,N_3568);
and U7374 (N_7374,N_3031,N_4561);
xor U7375 (N_7375,N_5468,N_4579);
and U7376 (N_7376,N_3787,N_5619);
and U7377 (N_7377,N_5278,N_4461);
and U7378 (N_7378,N_5119,N_3321);
and U7379 (N_7379,N_5195,N_5508);
nand U7380 (N_7380,N_3989,N_5805);
nor U7381 (N_7381,N_5346,N_4398);
xnor U7382 (N_7382,N_5724,N_5351);
xor U7383 (N_7383,N_4643,N_4245);
nand U7384 (N_7384,N_4583,N_3738);
and U7385 (N_7385,N_4771,N_4202);
xor U7386 (N_7386,N_3177,N_4614);
or U7387 (N_7387,N_3351,N_3270);
and U7388 (N_7388,N_5488,N_4487);
nor U7389 (N_7389,N_5561,N_4932);
nor U7390 (N_7390,N_3228,N_5409);
nor U7391 (N_7391,N_4287,N_5500);
nor U7392 (N_7392,N_5027,N_3098);
nor U7393 (N_7393,N_4844,N_3434);
nand U7394 (N_7394,N_3373,N_5181);
xor U7395 (N_7395,N_4068,N_3194);
xor U7396 (N_7396,N_5957,N_5164);
and U7397 (N_7397,N_5336,N_4422);
and U7398 (N_7398,N_4137,N_5744);
or U7399 (N_7399,N_5285,N_3308);
and U7400 (N_7400,N_5538,N_5631);
and U7401 (N_7401,N_5816,N_5618);
and U7402 (N_7402,N_4690,N_4672);
nand U7403 (N_7403,N_5750,N_4913);
nand U7404 (N_7404,N_3410,N_4903);
xnor U7405 (N_7405,N_4637,N_4754);
nand U7406 (N_7406,N_5904,N_4150);
nor U7407 (N_7407,N_3447,N_4892);
xnor U7408 (N_7408,N_5332,N_5338);
xnor U7409 (N_7409,N_4997,N_3229);
xor U7410 (N_7410,N_4382,N_3626);
nand U7411 (N_7411,N_4235,N_3591);
xnor U7412 (N_7412,N_5161,N_4345);
or U7413 (N_7413,N_5911,N_4756);
and U7414 (N_7414,N_3025,N_3815);
nand U7415 (N_7415,N_4276,N_4857);
xnor U7416 (N_7416,N_5122,N_5528);
and U7417 (N_7417,N_5407,N_3880);
nor U7418 (N_7418,N_4651,N_5651);
xnor U7419 (N_7419,N_3563,N_5728);
and U7420 (N_7420,N_5462,N_3757);
and U7421 (N_7421,N_3202,N_4187);
and U7422 (N_7422,N_5747,N_3454);
xor U7423 (N_7423,N_3158,N_5944);
and U7424 (N_7424,N_3921,N_5020);
nand U7425 (N_7425,N_4860,N_4100);
xor U7426 (N_7426,N_4962,N_5791);
nand U7427 (N_7427,N_4745,N_4693);
or U7428 (N_7428,N_5539,N_3142);
and U7429 (N_7429,N_3832,N_5306);
and U7430 (N_7430,N_3121,N_3012);
nor U7431 (N_7431,N_5131,N_5340);
and U7432 (N_7432,N_4797,N_5927);
nand U7433 (N_7433,N_3811,N_5379);
xor U7434 (N_7434,N_3824,N_4445);
nand U7435 (N_7435,N_3796,N_5158);
nor U7436 (N_7436,N_4078,N_3483);
nand U7437 (N_7437,N_5704,N_5268);
and U7438 (N_7438,N_4722,N_3019);
nor U7439 (N_7439,N_3115,N_5630);
or U7440 (N_7440,N_3079,N_4539);
nor U7441 (N_7441,N_3865,N_3425);
nand U7442 (N_7442,N_5355,N_3437);
and U7443 (N_7443,N_3705,N_4252);
xnor U7444 (N_7444,N_3424,N_5612);
or U7445 (N_7445,N_4540,N_3828);
xnor U7446 (N_7446,N_3631,N_3759);
xor U7447 (N_7447,N_4453,N_4140);
nor U7448 (N_7448,N_5738,N_3350);
nand U7449 (N_7449,N_5919,N_4634);
or U7450 (N_7450,N_5545,N_4750);
nor U7451 (N_7451,N_5787,N_3366);
nand U7452 (N_7452,N_3440,N_4941);
nor U7453 (N_7453,N_4196,N_4037);
nor U7454 (N_7454,N_3931,N_4138);
xor U7455 (N_7455,N_5685,N_4610);
or U7456 (N_7456,N_4095,N_3493);
and U7457 (N_7457,N_5129,N_5748);
or U7458 (N_7458,N_4869,N_5621);
nand U7459 (N_7459,N_5022,N_4303);
xnor U7460 (N_7460,N_3211,N_4831);
or U7461 (N_7461,N_5517,N_4415);
and U7462 (N_7462,N_3664,N_4506);
xor U7463 (N_7463,N_5458,N_4355);
or U7464 (N_7464,N_4106,N_4089);
and U7465 (N_7465,N_5925,N_5335);
nand U7466 (N_7466,N_4419,N_5451);
nor U7467 (N_7467,N_3381,N_3608);
nand U7468 (N_7468,N_5929,N_4007);
nand U7469 (N_7469,N_5722,N_4987);
xnor U7470 (N_7470,N_3869,N_4556);
and U7471 (N_7471,N_5344,N_3606);
and U7472 (N_7472,N_4193,N_5481);
nand U7473 (N_7473,N_3686,N_3593);
or U7474 (N_7474,N_3358,N_5405);
or U7475 (N_7475,N_3226,N_4806);
nor U7476 (N_7476,N_3732,N_5892);
nand U7477 (N_7477,N_5465,N_3214);
xnor U7478 (N_7478,N_5760,N_3278);
or U7479 (N_7479,N_5000,N_5776);
or U7480 (N_7480,N_4852,N_3694);
xor U7481 (N_7481,N_4197,N_3923);
nand U7482 (N_7482,N_3030,N_4977);
or U7483 (N_7483,N_5051,N_4388);
nand U7484 (N_7484,N_5875,N_3466);
or U7485 (N_7485,N_3871,N_5400);
xor U7486 (N_7486,N_5303,N_3622);
or U7487 (N_7487,N_4463,N_3331);
nor U7488 (N_7488,N_4147,N_4378);
xor U7489 (N_7489,N_3337,N_3844);
nand U7490 (N_7490,N_4096,N_3010);
or U7491 (N_7491,N_4135,N_3050);
and U7492 (N_7492,N_4227,N_3287);
and U7493 (N_7493,N_3678,N_3069);
nor U7494 (N_7494,N_5806,N_3949);
nand U7495 (N_7495,N_4699,N_4550);
xnor U7496 (N_7496,N_5479,N_3318);
and U7497 (N_7497,N_4972,N_5091);
xor U7498 (N_7498,N_5147,N_3059);
or U7499 (N_7499,N_5384,N_4807);
xnor U7500 (N_7500,N_5221,N_5793);
nand U7501 (N_7501,N_5672,N_3232);
nand U7502 (N_7502,N_3207,N_3297);
xor U7503 (N_7503,N_3019,N_5990);
xnor U7504 (N_7504,N_4731,N_5045);
xnor U7505 (N_7505,N_3373,N_4005);
and U7506 (N_7506,N_4703,N_4134);
or U7507 (N_7507,N_4177,N_5219);
nand U7508 (N_7508,N_4195,N_5535);
and U7509 (N_7509,N_5329,N_5068);
nor U7510 (N_7510,N_5683,N_3202);
and U7511 (N_7511,N_3429,N_3866);
and U7512 (N_7512,N_3285,N_5879);
or U7513 (N_7513,N_4761,N_4095);
or U7514 (N_7514,N_5459,N_5375);
nand U7515 (N_7515,N_4421,N_5806);
xnor U7516 (N_7516,N_3597,N_4106);
and U7517 (N_7517,N_5383,N_3322);
xor U7518 (N_7518,N_4869,N_5160);
and U7519 (N_7519,N_3998,N_3386);
and U7520 (N_7520,N_4316,N_5145);
nand U7521 (N_7521,N_4108,N_4110);
nor U7522 (N_7522,N_4249,N_5281);
xnor U7523 (N_7523,N_5503,N_4751);
or U7524 (N_7524,N_5116,N_3559);
and U7525 (N_7525,N_4200,N_4649);
and U7526 (N_7526,N_4254,N_3210);
and U7527 (N_7527,N_3711,N_4157);
xnor U7528 (N_7528,N_5220,N_3359);
nor U7529 (N_7529,N_5379,N_5885);
nand U7530 (N_7530,N_5122,N_3290);
and U7531 (N_7531,N_5668,N_3576);
and U7532 (N_7532,N_5762,N_5727);
nand U7533 (N_7533,N_4104,N_5096);
or U7534 (N_7534,N_5219,N_5200);
and U7535 (N_7535,N_4516,N_4205);
and U7536 (N_7536,N_5333,N_4905);
nor U7537 (N_7537,N_5592,N_5318);
nor U7538 (N_7538,N_4182,N_5162);
nand U7539 (N_7539,N_5725,N_3804);
or U7540 (N_7540,N_4456,N_3737);
or U7541 (N_7541,N_3275,N_5404);
nand U7542 (N_7542,N_3041,N_5178);
nand U7543 (N_7543,N_3122,N_4358);
xor U7544 (N_7544,N_4731,N_4152);
and U7545 (N_7545,N_3658,N_4020);
nor U7546 (N_7546,N_5339,N_5083);
and U7547 (N_7547,N_5247,N_3327);
or U7548 (N_7548,N_4176,N_3170);
nand U7549 (N_7549,N_3411,N_4630);
and U7550 (N_7550,N_5612,N_3477);
nor U7551 (N_7551,N_4261,N_3640);
xor U7552 (N_7552,N_3159,N_5606);
or U7553 (N_7553,N_4625,N_3880);
nand U7554 (N_7554,N_4940,N_4166);
nand U7555 (N_7555,N_5639,N_3157);
and U7556 (N_7556,N_4858,N_5273);
nor U7557 (N_7557,N_4327,N_4903);
nand U7558 (N_7558,N_5997,N_3009);
and U7559 (N_7559,N_3005,N_4152);
nand U7560 (N_7560,N_4516,N_4064);
and U7561 (N_7561,N_4527,N_4925);
xnor U7562 (N_7562,N_4558,N_3629);
nand U7563 (N_7563,N_5665,N_4371);
nor U7564 (N_7564,N_3729,N_5100);
and U7565 (N_7565,N_3931,N_4566);
and U7566 (N_7566,N_3614,N_5818);
or U7567 (N_7567,N_3149,N_4195);
or U7568 (N_7568,N_5100,N_3637);
nor U7569 (N_7569,N_4214,N_5903);
or U7570 (N_7570,N_3754,N_4831);
nor U7571 (N_7571,N_3910,N_4280);
nand U7572 (N_7572,N_3417,N_5544);
nor U7573 (N_7573,N_4865,N_3488);
or U7574 (N_7574,N_3939,N_4158);
and U7575 (N_7575,N_5736,N_5054);
nor U7576 (N_7576,N_3605,N_3415);
or U7577 (N_7577,N_3768,N_4253);
or U7578 (N_7578,N_3525,N_4918);
and U7579 (N_7579,N_5630,N_5502);
xnor U7580 (N_7580,N_3512,N_4097);
and U7581 (N_7581,N_5777,N_3019);
or U7582 (N_7582,N_3115,N_5689);
nand U7583 (N_7583,N_5894,N_3497);
and U7584 (N_7584,N_4407,N_4949);
xnor U7585 (N_7585,N_3553,N_4722);
nand U7586 (N_7586,N_3317,N_4647);
and U7587 (N_7587,N_4365,N_3170);
and U7588 (N_7588,N_3898,N_3194);
nor U7589 (N_7589,N_3249,N_4909);
nor U7590 (N_7590,N_4954,N_3170);
xor U7591 (N_7591,N_5821,N_3427);
or U7592 (N_7592,N_4205,N_4706);
nand U7593 (N_7593,N_5497,N_3917);
and U7594 (N_7594,N_3510,N_4865);
or U7595 (N_7595,N_4848,N_3027);
and U7596 (N_7596,N_4051,N_5229);
nor U7597 (N_7597,N_4477,N_4833);
nor U7598 (N_7598,N_3369,N_5564);
nand U7599 (N_7599,N_4451,N_3461);
or U7600 (N_7600,N_5174,N_5881);
nand U7601 (N_7601,N_4291,N_3395);
and U7602 (N_7602,N_3496,N_5995);
or U7603 (N_7603,N_4075,N_3294);
and U7604 (N_7604,N_4493,N_5782);
nand U7605 (N_7605,N_5727,N_4056);
nand U7606 (N_7606,N_4213,N_4136);
and U7607 (N_7607,N_4748,N_5544);
nor U7608 (N_7608,N_3095,N_5632);
nor U7609 (N_7609,N_5159,N_4841);
xnor U7610 (N_7610,N_3136,N_5474);
nand U7611 (N_7611,N_3883,N_5710);
and U7612 (N_7612,N_5020,N_5162);
and U7613 (N_7613,N_3639,N_5505);
and U7614 (N_7614,N_3343,N_4100);
nand U7615 (N_7615,N_4870,N_3939);
nand U7616 (N_7616,N_4849,N_3038);
and U7617 (N_7617,N_4138,N_3844);
or U7618 (N_7618,N_4553,N_3053);
or U7619 (N_7619,N_3013,N_4343);
and U7620 (N_7620,N_3777,N_3361);
and U7621 (N_7621,N_3293,N_5468);
and U7622 (N_7622,N_5804,N_4320);
and U7623 (N_7623,N_5789,N_4410);
nand U7624 (N_7624,N_3502,N_4616);
nor U7625 (N_7625,N_3957,N_3302);
or U7626 (N_7626,N_4044,N_5869);
nor U7627 (N_7627,N_5811,N_5161);
nand U7628 (N_7628,N_3401,N_5893);
xor U7629 (N_7629,N_5271,N_3950);
and U7630 (N_7630,N_4591,N_3027);
or U7631 (N_7631,N_5378,N_4299);
nor U7632 (N_7632,N_4412,N_4519);
nand U7633 (N_7633,N_4623,N_4859);
nand U7634 (N_7634,N_4154,N_3817);
or U7635 (N_7635,N_3098,N_5004);
nor U7636 (N_7636,N_5838,N_5355);
or U7637 (N_7637,N_3901,N_3540);
xor U7638 (N_7638,N_4188,N_5252);
nor U7639 (N_7639,N_5143,N_4105);
or U7640 (N_7640,N_4405,N_3408);
or U7641 (N_7641,N_4742,N_5824);
and U7642 (N_7642,N_4100,N_3097);
or U7643 (N_7643,N_3574,N_5277);
nand U7644 (N_7644,N_5165,N_5558);
and U7645 (N_7645,N_5516,N_3104);
xor U7646 (N_7646,N_4570,N_3012);
and U7647 (N_7647,N_3082,N_4647);
xnor U7648 (N_7648,N_3106,N_3334);
xor U7649 (N_7649,N_3813,N_3574);
or U7650 (N_7650,N_4182,N_4530);
nand U7651 (N_7651,N_3009,N_4206);
nor U7652 (N_7652,N_4941,N_4815);
or U7653 (N_7653,N_3052,N_3884);
nor U7654 (N_7654,N_4644,N_3653);
nand U7655 (N_7655,N_5500,N_4500);
or U7656 (N_7656,N_4205,N_4978);
nand U7657 (N_7657,N_3407,N_3969);
xnor U7658 (N_7658,N_4752,N_3906);
nand U7659 (N_7659,N_5513,N_5517);
nor U7660 (N_7660,N_4093,N_4609);
nand U7661 (N_7661,N_5093,N_5160);
or U7662 (N_7662,N_5329,N_4628);
nor U7663 (N_7663,N_3617,N_3346);
xnor U7664 (N_7664,N_4260,N_3604);
nand U7665 (N_7665,N_3382,N_4147);
nor U7666 (N_7666,N_5586,N_3792);
nor U7667 (N_7667,N_4709,N_4242);
or U7668 (N_7668,N_3362,N_3184);
or U7669 (N_7669,N_4567,N_4622);
nand U7670 (N_7670,N_5163,N_4551);
and U7671 (N_7671,N_3548,N_3978);
xor U7672 (N_7672,N_4887,N_5949);
nor U7673 (N_7673,N_3823,N_5738);
or U7674 (N_7674,N_3931,N_4841);
nand U7675 (N_7675,N_5206,N_5384);
nor U7676 (N_7676,N_4071,N_4801);
xnor U7677 (N_7677,N_4372,N_5355);
nand U7678 (N_7678,N_4813,N_3939);
xnor U7679 (N_7679,N_5513,N_5391);
and U7680 (N_7680,N_5199,N_4170);
and U7681 (N_7681,N_3193,N_4725);
nand U7682 (N_7682,N_5590,N_3030);
xnor U7683 (N_7683,N_3680,N_4751);
and U7684 (N_7684,N_4312,N_3785);
xor U7685 (N_7685,N_4756,N_5164);
or U7686 (N_7686,N_4728,N_3017);
nor U7687 (N_7687,N_4519,N_3434);
nor U7688 (N_7688,N_5485,N_5005);
or U7689 (N_7689,N_5235,N_4781);
or U7690 (N_7690,N_3843,N_4821);
and U7691 (N_7691,N_5404,N_3156);
nand U7692 (N_7692,N_4240,N_3288);
or U7693 (N_7693,N_3681,N_3669);
nor U7694 (N_7694,N_4593,N_3617);
nor U7695 (N_7695,N_4648,N_4013);
nand U7696 (N_7696,N_3938,N_5443);
nand U7697 (N_7697,N_4952,N_3422);
or U7698 (N_7698,N_3416,N_3494);
and U7699 (N_7699,N_3770,N_4569);
nand U7700 (N_7700,N_3236,N_4056);
nand U7701 (N_7701,N_5221,N_3356);
xnor U7702 (N_7702,N_3673,N_3174);
or U7703 (N_7703,N_3624,N_4893);
nor U7704 (N_7704,N_3415,N_3867);
nor U7705 (N_7705,N_3151,N_3256);
xor U7706 (N_7706,N_4617,N_3503);
nor U7707 (N_7707,N_3344,N_4039);
nand U7708 (N_7708,N_3718,N_5416);
and U7709 (N_7709,N_4437,N_4887);
and U7710 (N_7710,N_5659,N_5437);
xor U7711 (N_7711,N_4677,N_3351);
or U7712 (N_7712,N_4570,N_4673);
nand U7713 (N_7713,N_4062,N_5583);
or U7714 (N_7714,N_5350,N_3867);
or U7715 (N_7715,N_3561,N_3170);
nand U7716 (N_7716,N_5422,N_4963);
nand U7717 (N_7717,N_4326,N_5972);
nand U7718 (N_7718,N_3013,N_5589);
xor U7719 (N_7719,N_5439,N_3170);
or U7720 (N_7720,N_5095,N_3984);
or U7721 (N_7721,N_5524,N_3953);
xor U7722 (N_7722,N_5123,N_4172);
nand U7723 (N_7723,N_5185,N_3059);
or U7724 (N_7724,N_5013,N_5090);
nand U7725 (N_7725,N_4119,N_5903);
and U7726 (N_7726,N_5943,N_3920);
and U7727 (N_7727,N_3951,N_5891);
or U7728 (N_7728,N_3490,N_4017);
or U7729 (N_7729,N_3019,N_4943);
and U7730 (N_7730,N_5468,N_5246);
and U7731 (N_7731,N_4754,N_5802);
xor U7732 (N_7732,N_5829,N_4490);
nor U7733 (N_7733,N_5580,N_3648);
nor U7734 (N_7734,N_5503,N_4235);
xor U7735 (N_7735,N_3529,N_4270);
and U7736 (N_7736,N_4196,N_3516);
xor U7737 (N_7737,N_4838,N_5414);
nand U7738 (N_7738,N_3222,N_5537);
nand U7739 (N_7739,N_3737,N_3659);
nand U7740 (N_7740,N_4823,N_4970);
or U7741 (N_7741,N_4041,N_3101);
nor U7742 (N_7742,N_4815,N_3795);
and U7743 (N_7743,N_5173,N_4836);
and U7744 (N_7744,N_5859,N_5989);
xnor U7745 (N_7745,N_5555,N_3488);
or U7746 (N_7746,N_3417,N_5779);
and U7747 (N_7747,N_4378,N_4511);
nand U7748 (N_7748,N_4811,N_5918);
nand U7749 (N_7749,N_4375,N_3619);
or U7750 (N_7750,N_3752,N_5011);
or U7751 (N_7751,N_3714,N_4169);
and U7752 (N_7752,N_4302,N_5971);
nor U7753 (N_7753,N_4341,N_5529);
xnor U7754 (N_7754,N_5215,N_3306);
nor U7755 (N_7755,N_4431,N_3339);
xor U7756 (N_7756,N_3702,N_3282);
nor U7757 (N_7757,N_3784,N_5835);
or U7758 (N_7758,N_4657,N_3118);
or U7759 (N_7759,N_5185,N_4338);
xor U7760 (N_7760,N_3288,N_5010);
nand U7761 (N_7761,N_3491,N_5567);
nand U7762 (N_7762,N_4570,N_5016);
nand U7763 (N_7763,N_5634,N_3575);
nand U7764 (N_7764,N_4565,N_4182);
xnor U7765 (N_7765,N_5931,N_5518);
xor U7766 (N_7766,N_3565,N_4075);
and U7767 (N_7767,N_4444,N_4386);
xnor U7768 (N_7768,N_4385,N_3770);
and U7769 (N_7769,N_4493,N_5013);
and U7770 (N_7770,N_5596,N_3672);
nor U7771 (N_7771,N_4859,N_5835);
or U7772 (N_7772,N_3274,N_3585);
xor U7773 (N_7773,N_4782,N_3794);
xor U7774 (N_7774,N_5102,N_5605);
and U7775 (N_7775,N_3487,N_3291);
xnor U7776 (N_7776,N_5035,N_5447);
nand U7777 (N_7777,N_4202,N_3971);
xor U7778 (N_7778,N_4516,N_4641);
nand U7779 (N_7779,N_4802,N_3309);
nand U7780 (N_7780,N_5012,N_4633);
and U7781 (N_7781,N_3367,N_4373);
and U7782 (N_7782,N_4835,N_4418);
xor U7783 (N_7783,N_4249,N_4748);
or U7784 (N_7784,N_3704,N_4152);
nand U7785 (N_7785,N_5037,N_3913);
nand U7786 (N_7786,N_5587,N_4791);
xor U7787 (N_7787,N_3314,N_5752);
and U7788 (N_7788,N_5296,N_4601);
nand U7789 (N_7789,N_3881,N_5329);
or U7790 (N_7790,N_4392,N_4945);
nand U7791 (N_7791,N_4350,N_4499);
nand U7792 (N_7792,N_3269,N_3164);
or U7793 (N_7793,N_5030,N_4828);
nand U7794 (N_7794,N_4220,N_4511);
and U7795 (N_7795,N_4445,N_3245);
nand U7796 (N_7796,N_4829,N_3237);
nor U7797 (N_7797,N_5705,N_5450);
or U7798 (N_7798,N_5968,N_3298);
or U7799 (N_7799,N_4525,N_4281);
nand U7800 (N_7800,N_4620,N_4726);
xnor U7801 (N_7801,N_5895,N_3341);
or U7802 (N_7802,N_4118,N_5169);
or U7803 (N_7803,N_5094,N_3230);
nand U7804 (N_7804,N_4639,N_3695);
xnor U7805 (N_7805,N_3526,N_4020);
nand U7806 (N_7806,N_5232,N_4203);
and U7807 (N_7807,N_5551,N_3713);
xor U7808 (N_7808,N_3159,N_5473);
or U7809 (N_7809,N_4023,N_5294);
and U7810 (N_7810,N_3390,N_5653);
nor U7811 (N_7811,N_3932,N_4867);
nor U7812 (N_7812,N_3184,N_4176);
and U7813 (N_7813,N_3345,N_3954);
nor U7814 (N_7814,N_4420,N_4707);
or U7815 (N_7815,N_3824,N_4464);
and U7816 (N_7816,N_5803,N_4522);
or U7817 (N_7817,N_4269,N_5203);
or U7818 (N_7818,N_5735,N_5684);
and U7819 (N_7819,N_3522,N_5148);
xnor U7820 (N_7820,N_3710,N_5532);
and U7821 (N_7821,N_3548,N_5799);
nand U7822 (N_7822,N_3939,N_5886);
or U7823 (N_7823,N_4353,N_5711);
xor U7824 (N_7824,N_3183,N_5503);
and U7825 (N_7825,N_3840,N_5960);
nor U7826 (N_7826,N_5823,N_5405);
xor U7827 (N_7827,N_5217,N_3867);
or U7828 (N_7828,N_4954,N_5927);
nor U7829 (N_7829,N_4066,N_3659);
xnor U7830 (N_7830,N_4353,N_5573);
xor U7831 (N_7831,N_5740,N_5265);
nand U7832 (N_7832,N_4523,N_5173);
xor U7833 (N_7833,N_5261,N_3108);
nor U7834 (N_7834,N_5443,N_3018);
nand U7835 (N_7835,N_5089,N_4572);
xor U7836 (N_7836,N_5041,N_3562);
and U7837 (N_7837,N_5776,N_4230);
xor U7838 (N_7838,N_3389,N_3809);
nor U7839 (N_7839,N_5987,N_4067);
xor U7840 (N_7840,N_5202,N_3021);
nor U7841 (N_7841,N_3518,N_3312);
xnor U7842 (N_7842,N_4986,N_3833);
or U7843 (N_7843,N_4640,N_5680);
or U7844 (N_7844,N_4647,N_4039);
nand U7845 (N_7845,N_3549,N_4886);
nor U7846 (N_7846,N_5014,N_5513);
nor U7847 (N_7847,N_5568,N_5700);
and U7848 (N_7848,N_4044,N_5745);
and U7849 (N_7849,N_3844,N_5612);
and U7850 (N_7850,N_5661,N_5077);
xnor U7851 (N_7851,N_4597,N_4311);
and U7852 (N_7852,N_4673,N_3532);
nand U7853 (N_7853,N_3788,N_4117);
xnor U7854 (N_7854,N_4492,N_3221);
nand U7855 (N_7855,N_3133,N_4965);
nor U7856 (N_7856,N_4568,N_3651);
nand U7857 (N_7857,N_4274,N_4525);
nand U7858 (N_7858,N_5270,N_3094);
xnor U7859 (N_7859,N_5148,N_3036);
xor U7860 (N_7860,N_4445,N_5419);
or U7861 (N_7861,N_3031,N_4627);
or U7862 (N_7862,N_4318,N_5129);
nor U7863 (N_7863,N_3922,N_4636);
nand U7864 (N_7864,N_4489,N_4586);
or U7865 (N_7865,N_3446,N_5244);
xor U7866 (N_7866,N_4377,N_5691);
nor U7867 (N_7867,N_3789,N_4437);
xor U7868 (N_7868,N_5939,N_4554);
and U7869 (N_7869,N_5479,N_4021);
xnor U7870 (N_7870,N_4789,N_3091);
xnor U7871 (N_7871,N_3408,N_3846);
nand U7872 (N_7872,N_5644,N_5802);
or U7873 (N_7873,N_4309,N_5991);
nor U7874 (N_7874,N_5459,N_3702);
nor U7875 (N_7875,N_3136,N_4802);
nand U7876 (N_7876,N_3109,N_4977);
or U7877 (N_7877,N_5313,N_5925);
nand U7878 (N_7878,N_4797,N_3574);
and U7879 (N_7879,N_5543,N_3904);
and U7880 (N_7880,N_3789,N_5203);
xnor U7881 (N_7881,N_5946,N_3950);
nand U7882 (N_7882,N_5895,N_3463);
xor U7883 (N_7883,N_5580,N_3505);
or U7884 (N_7884,N_5102,N_3686);
and U7885 (N_7885,N_3780,N_4560);
xnor U7886 (N_7886,N_5274,N_3411);
xnor U7887 (N_7887,N_3716,N_4668);
nor U7888 (N_7888,N_4780,N_3615);
nand U7889 (N_7889,N_5832,N_5134);
and U7890 (N_7890,N_3923,N_5738);
nand U7891 (N_7891,N_5251,N_4884);
xnor U7892 (N_7892,N_4312,N_3276);
or U7893 (N_7893,N_3494,N_4822);
or U7894 (N_7894,N_4097,N_5412);
or U7895 (N_7895,N_4392,N_3721);
or U7896 (N_7896,N_5625,N_4155);
nor U7897 (N_7897,N_5991,N_5039);
nand U7898 (N_7898,N_4315,N_5633);
and U7899 (N_7899,N_3510,N_3669);
nor U7900 (N_7900,N_5793,N_5690);
or U7901 (N_7901,N_5604,N_5252);
xor U7902 (N_7902,N_5414,N_5652);
and U7903 (N_7903,N_5335,N_4010);
nor U7904 (N_7904,N_5155,N_3891);
nand U7905 (N_7905,N_4168,N_4370);
xnor U7906 (N_7906,N_5377,N_5946);
nand U7907 (N_7907,N_3252,N_4569);
nand U7908 (N_7908,N_3741,N_3546);
nand U7909 (N_7909,N_5290,N_5717);
nand U7910 (N_7910,N_3436,N_5229);
xnor U7911 (N_7911,N_5569,N_5185);
or U7912 (N_7912,N_4108,N_4226);
or U7913 (N_7913,N_4090,N_3226);
or U7914 (N_7914,N_5185,N_3795);
xnor U7915 (N_7915,N_5338,N_5831);
and U7916 (N_7916,N_5817,N_3533);
xnor U7917 (N_7917,N_3311,N_5946);
and U7918 (N_7918,N_4882,N_4903);
or U7919 (N_7919,N_3220,N_3319);
and U7920 (N_7920,N_4771,N_4706);
nand U7921 (N_7921,N_5464,N_3477);
or U7922 (N_7922,N_4817,N_3611);
and U7923 (N_7923,N_4153,N_3950);
nor U7924 (N_7924,N_5994,N_4074);
nand U7925 (N_7925,N_5113,N_5440);
or U7926 (N_7926,N_4851,N_5948);
and U7927 (N_7927,N_5712,N_3811);
xnor U7928 (N_7928,N_5905,N_4385);
nor U7929 (N_7929,N_4691,N_3309);
and U7930 (N_7930,N_3038,N_3781);
nor U7931 (N_7931,N_3952,N_3999);
nor U7932 (N_7932,N_4978,N_3629);
xor U7933 (N_7933,N_3641,N_4304);
xor U7934 (N_7934,N_3435,N_5666);
or U7935 (N_7935,N_3057,N_5253);
xnor U7936 (N_7936,N_3633,N_4789);
nand U7937 (N_7937,N_4640,N_3782);
nor U7938 (N_7938,N_3666,N_3115);
or U7939 (N_7939,N_3003,N_4741);
and U7940 (N_7940,N_3432,N_5451);
and U7941 (N_7941,N_4131,N_4972);
xor U7942 (N_7942,N_4243,N_5739);
nand U7943 (N_7943,N_3434,N_5910);
nand U7944 (N_7944,N_3246,N_5622);
xor U7945 (N_7945,N_4015,N_5161);
nand U7946 (N_7946,N_3151,N_4161);
xnor U7947 (N_7947,N_5907,N_5530);
or U7948 (N_7948,N_4544,N_3423);
or U7949 (N_7949,N_3118,N_5197);
nor U7950 (N_7950,N_5933,N_5514);
and U7951 (N_7951,N_3091,N_5327);
and U7952 (N_7952,N_4995,N_5403);
xnor U7953 (N_7953,N_3449,N_4748);
xor U7954 (N_7954,N_5339,N_5871);
nor U7955 (N_7955,N_4605,N_5572);
or U7956 (N_7956,N_5991,N_5904);
xnor U7957 (N_7957,N_4829,N_5908);
or U7958 (N_7958,N_5236,N_4019);
or U7959 (N_7959,N_5042,N_3030);
or U7960 (N_7960,N_4754,N_5773);
nand U7961 (N_7961,N_4135,N_5842);
or U7962 (N_7962,N_3166,N_5403);
or U7963 (N_7963,N_5241,N_5472);
nand U7964 (N_7964,N_4790,N_5994);
nand U7965 (N_7965,N_4957,N_3955);
nor U7966 (N_7966,N_3333,N_5277);
xor U7967 (N_7967,N_5926,N_5752);
nand U7968 (N_7968,N_5814,N_4834);
or U7969 (N_7969,N_3538,N_5832);
or U7970 (N_7970,N_5317,N_3627);
and U7971 (N_7971,N_5491,N_4216);
nand U7972 (N_7972,N_5435,N_4283);
or U7973 (N_7973,N_4265,N_5385);
and U7974 (N_7974,N_3429,N_4256);
nand U7975 (N_7975,N_5088,N_3892);
and U7976 (N_7976,N_4166,N_5119);
nor U7977 (N_7977,N_5018,N_5225);
nand U7978 (N_7978,N_3156,N_3651);
and U7979 (N_7979,N_3550,N_5283);
or U7980 (N_7980,N_5125,N_4845);
nand U7981 (N_7981,N_3870,N_5674);
and U7982 (N_7982,N_5807,N_3169);
or U7983 (N_7983,N_3092,N_4301);
xnor U7984 (N_7984,N_4595,N_4853);
nor U7985 (N_7985,N_3589,N_3779);
nor U7986 (N_7986,N_3024,N_5502);
nor U7987 (N_7987,N_3430,N_5410);
nor U7988 (N_7988,N_5764,N_4624);
nand U7989 (N_7989,N_5718,N_3607);
or U7990 (N_7990,N_3528,N_4769);
and U7991 (N_7991,N_3862,N_4405);
nand U7992 (N_7992,N_4699,N_5266);
and U7993 (N_7993,N_3194,N_5522);
and U7994 (N_7994,N_5769,N_3720);
nand U7995 (N_7995,N_4691,N_3903);
or U7996 (N_7996,N_3624,N_4305);
or U7997 (N_7997,N_4810,N_5099);
or U7998 (N_7998,N_5366,N_5884);
xnor U7999 (N_7999,N_3010,N_5675);
nand U8000 (N_8000,N_4258,N_3934);
nand U8001 (N_8001,N_5162,N_4554);
and U8002 (N_8002,N_4676,N_5827);
and U8003 (N_8003,N_4341,N_5914);
nor U8004 (N_8004,N_4763,N_5680);
nor U8005 (N_8005,N_4766,N_5253);
xor U8006 (N_8006,N_5783,N_5830);
xor U8007 (N_8007,N_3188,N_4976);
or U8008 (N_8008,N_5188,N_5001);
and U8009 (N_8009,N_3449,N_4756);
or U8010 (N_8010,N_3739,N_3951);
and U8011 (N_8011,N_4482,N_5098);
nand U8012 (N_8012,N_3099,N_5438);
xor U8013 (N_8013,N_4721,N_4431);
xnor U8014 (N_8014,N_5010,N_5130);
and U8015 (N_8015,N_5959,N_4878);
nor U8016 (N_8016,N_5026,N_5061);
and U8017 (N_8017,N_3425,N_4475);
and U8018 (N_8018,N_4232,N_3894);
or U8019 (N_8019,N_5953,N_3668);
and U8020 (N_8020,N_5791,N_5903);
nor U8021 (N_8021,N_3182,N_5595);
xor U8022 (N_8022,N_4831,N_3599);
nor U8023 (N_8023,N_3311,N_4674);
nor U8024 (N_8024,N_5865,N_5147);
nand U8025 (N_8025,N_4173,N_4339);
nor U8026 (N_8026,N_4966,N_5054);
nor U8027 (N_8027,N_5459,N_3062);
and U8028 (N_8028,N_3251,N_4228);
nand U8029 (N_8029,N_5805,N_4917);
or U8030 (N_8030,N_5152,N_3575);
nand U8031 (N_8031,N_3071,N_5995);
xor U8032 (N_8032,N_3903,N_5649);
nand U8033 (N_8033,N_5839,N_3539);
xnor U8034 (N_8034,N_5902,N_3299);
and U8035 (N_8035,N_5932,N_5069);
and U8036 (N_8036,N_5718,N_5217);
nor U8037 (N_8037,N_3994,N_3316);
xor U8038 (N_8038,N_3307,N_4673);
nand U8039 (N_8039,N_5042,N_3545);
nor U8040 (N_8040,N_5211,N_5050);
nor U8041 (N_8041,N_5460,N_3216);
xor U8042 (N_8042,N_5568,N_4281);
xor U8043 (N_8043,N_3374,N_5788);
or U8044 (N_8044,N_5504,N_5656);
and U8045 (N_8045,N_5767,N_5635);
and U8046 (N_8046,N_4982,N_3306);
or U8047 (N_8047,N_4410,N_3045);
xor U8048 (N_8048,N_4823,N_3136);
nand U8049 (N_8049,N_3272,N_3792);
and U8050 (N_8050,N_3562,N_3079);
and U8051 (N_8051,N_3614,N_3599);
and U8052 (N_8052,N_4774,N_3686);
xor U8053 (N_8053,N_4667,N_3324);
or U8054 (N_8054,N_5075,N_3251);
xnor U8055 (N_8055,N_4417,N_3752);
and U8056 (N_8056,N_3887,N_3303);
xor U8057 (N_8057,N_3399,N_5773);
and U8058 (N_8058,N_5637,N_5877);
or U8059 (N_8059,N_5958,N_3495);
nor U8060 (N_8060,N_4416,N_4071);
nor U8061 (N_8061,N_5139,N_5290);
xor U8062 (N_8062,N_5472,N_4177);
nand U8063 (N_8063,N_4826,N_5184);
nor U8064 (N_8064,N_5900,N_5108);
or U8065 (N_8065,N_3175,N_5416);
or U8066 (N_8066,N_3953,N_4151);
xor U8067 (N_8067,N_5704,N_5593);
nand U8068 (N_8068,N_3908,N_4176);
nor U8069 (N_8069,N_5283,N_5253);
xnor U8070 (N_8070,N_5884,N_5248);
xnor U8071 (N_8071,N_4016,N_5537);
or U8072 (N_8072,N_3640,N_5533);
xor U8073 (N_8073,N_4914,N_4973);
or U8074 (N_8074,N_5452,N_4886);
and U8075 (N_8075,N_3295,N_3121);
nand U8076 (N_8076,N_5622,N_3295);
xor U8077 (N_8077,N_5424,N_4793);
or U8078 (N_8078,N_4833,N_5462);
or U8079 (N_8079,N_4209,N_5687);
xor U8080 (N_8080,N_3867,N_4532);
nand U8081 (N_8081,N_5408,N_4758);
or U8082 (N_8082,N_4206,N_3689);
or U8083 (N_8083,N_3109,N_3669);
xor U8084 (N_8084,N_3482,N_5481);
or U8085 (N_8085,N_3741,N_5084);
nand U8086 (N_8086,N_3509,N_4470);
or U8087 (N_8087,N_3331,N_3269);
nor U8088 (N_8088,N_3507,N_4420);
nor U8089 (N_8089,N_3610,N_5367);
and U8090 (N_8090,N_5652,N_3841);
xnor U8091 (N_8091,N_4895,N_3188);
and U8092 (N_8092,N_3393,N_3673);
or U8093 (N_8093,N_5300,N_3384);
or U8094 (N_8094,N_3854,N_5078);
or U8095 (N_8095,N_4217,N_5406);
or U8096 (N_8096,N_4734,N_3438);
nor U8097 (N_8097,N_3344,N_3617);
and U8098 (N_8098,N_5939,N_5033);
and U8099 (N_8099,N_3109,N_5525);
and U8100 (N_8100,N_5618,N_3518);
and U8101 (N_8101,N_5972,N_4535);
xor U8102 (N_8102,N_3790,N_3649);
nand U8103 (N_8103,N_5084,N_4521);
nor U8104 (N_8104,N_4494,N_3256);
and U8105 (N_8105,N_3339,N_4436);
nor U8106 (N_8106,N_5991,N_4830);
nor U8107 (N_8107,N_5675,N_3861);
or U8108 (N_8108,N_5347,N_5154);
nor U8109 (N_8109,N_3588,N_4506);
nand U8110 (N_8110,N_3561,N_5596);
and U8111 (N_8111,N_5785,N_5764);
xnor U8112 (N_8112,N_5225,N_4002);
nor U8113 (N_8113,N_5330,N_3005);
nor U8114 (N_8114,N_3797,N_3739);
xor U8115 (N_8115,N_4761,N_5191);
or U8116 (N_8116,N_4894,N_4142);
nand U8117 (N_8117,N_3907,N_3198);
xor U8118 (N_8118,N_4460,N_5669);
nor U8119 (N_8119,N_4398,N_3085);
or U8120 (N_8120,N_4496,N_5271);
nor U8121 (N_8121,N_3113,N_4508);
and U8122 (N_8122,N_4523,N_4892);
xor U8123 (N_8123,N_4506,N_3376);
xor U8124 (N_8124,N_5071,N_3354);
nor U8125 (N_8125,N_4646,N_3148);
nor U8126 (N_8126,N_5508,N_4327);
or U8127 (N_8127,N_5077,N_4282);
and U8128 (N_8128,N_3139,N_3023);
nor U8129 (N_8129,N_3430,N_4098);
and U8130 (N_8130,N_3576,N_3647);
nand U8131 (N_8131,N_4856,N_4151);
xnor U8132 (N_8132,N_3235,N_3142);
or U8133 (N_8133,N_5551,N_4627);
nand U8134 (N_8134,N_3458,N_3384);
or U8135 (N_8135,N_4040,N_3592);
nor U8136 (N_8136,N_3828,N_3213);
xnor U8137 (N_8137,N_4773,N_5091);
or U8138 (N_8138,N_5531,N_3357);
or U8139 (N_8139,N_3770,N_5850);
nand U8140 (N_8140,N_3234,N_5690);
or U8141 (N_8141,N_4135,N_4783);
nand U8142 (N_8142,N_3788,N_4588);
or U8143 (N_8143,N_3747,N_4149);
xor U8144 (N_8144,N_5674,N_4124);
or U8145 (N_8145,N_4212,N_5169);
and U8146 (N_8146,N_4241,N_3021);
nand U8147 (N_8147,N_5236,N_4345);
or U8148 (N_8148,N_4930,N_5246);
and U8149 (N_8149,N_3876,N_3445);
or U8150 (N_8150,N_5050,N_5613);
or U8151 (N_8151,N_4519,N_5351);
xor U8152 (N_8152,N_4894,N_3186);
or U8153 (N_8153,N_4240,N_4404);
or U8154 (N_8154,N_4277,N_4089);
and U8155 (N_8155,N_3247,N_3743);
nand U8156 (N_8156,N_4949,N_4611);
nor U8157 (N_8157,N_4791,N_3320);
nand U8158 (N_8158,N_3592,N_5450);
nand U8159 (N_8159,N_5483,N_5268);
or U8160 (N_8160,N_5781,N_4574);
or U8161 (N_8161,N_4083,N_3695);
or U8162 (N_8162,N_4151,N_4041);
nand U8163 (N_8163,N_5250,N_3716);
nand U8164 (N_8164,N_5365,N_4601);
nand U8165 (N_8165,N_5519,N_5560);
nand U8166 (N_8166,N_5211,N_3503);
nor U8167 (N_8167,N_5576,N_3478);
nor U8168 (N_8168,N_4639,N_3659);
and U8169 (N_8169,N_4953,N_5789);
nor U8170 (N_8170,N_5456,N_4375);
and U8171 (N_8171,N_4910,N_5588);
and U8172 (N_8172,N_5554,N_3459);
and U8173 (N_8173,N_3013,N_3162);
and U8174 (N_8174,N_4572,N_5652);
and U8175 (N_8175,N_4449,N_4045);
nor U8176 (N_8176,N_3943,N_5866);
and U8177 (N_8177,N_3996,N_3418);
nor U8178 (N_8178,N_4622,N_3052);
nor U8179 (N_8179,N_3032,N_3952);
nor U8180 (N_8180,N_5900,N_3499);
and U8181 (N_8181,N_4633,N_4974);
or U8182 (N_8182,N_5330,N_3443);
and U8183 (N_8183,N_5436,N_5848);
or U8184 (N_8184,N_5605,N_4056);
or U8185 (N_8185,N_3019,N_5488);
nor U8186 (N_8186,N_4375,N_4456);
or U8187 (N_8187,N_3280,N_5475);
nand U8188 (N_8188,N_3673,N_3196);
and U8189 (N_8189,N_5422,N_3246);
nand U8190 (N_8190,N_3303,N_5481);
or U8191 (N_8191,N_3908,N_3220);
nand U8192 (N_8192,N_4555,N_4055);
nand U8193 (N_8193,N_5901,N_5609);
nand U8194 (N_8194,N_4297,N_5903);
or U8195 (N_8195,N_4043,N_5779);
or U8196 (N_8196,N_4819,N_4872);
or U8197 (N_8197,N_5801,N_3425);
nand U8198 (N_8198,N_4664,N_3198);
xnor U8199 (N_8199,N_3956,N_4138);
nand U8200 (N_8200,N_5899,N_3193);
nor U8201 (N_8201,N_5521,N_4025);
nand U8202 (N_8202,N_4514,N_5041);
or U8203 (N_8203,N_4388,N_4657);
nor U8204 (N_8204,N_4157,N_5149);
or U8205 (N_8205,N_4029,N_3190);
xnor U8206 (N_8206,N_3069,N_5527);
and U8207 (N_8207,N_5914,N_5890);
nand U8208 (N_8208,N_5946,N_5607);
nor U8209 (N_8209,N_3842,N_4305);
or U8210 (N_8210,N_3094,N_5859);
or U8211 (N_8211,N_5055,N_4138);
xnor U8212 (N_8212,N_4983,N_3555);
or U8213 (N_8213,N_3100,N_4059);
or U8214 (N_8214,N_5756,N_3518);
xor U8215 (N_8215,N_3074,N_4127);
xor U8216 (N_8216,N_4246,N_3501);
and U8217 (N_8217,N_5634,N_3049);
and U8218 (N_8218,N_4020,N_5235);
and U8219 (N_8219,N_4810,N_5587);
and U8220 (N_8220,N_5438,N_5685);
nand U8221 (N_8221,N_3531,N_3878);
nand U8222 (N_8222,N_5786,N_3939);
nand U8223 (N_8223,N_5570,N_4539);
nor U8224 (N_8224,N_4660,N_5385);
and U8225 (N_8225,N_3883,N_3764);
xnor U8226 (N_8226,N_4696,N_4831);
or U8227 (N_8227,N_5631,N_5768);
and U8228 (N_8228,N_5151,N_4747);
nand U8229 (N_8229,N_4612,N_3363);
or U8230 (N_8230,N_4573,N_5319);
xor U8231 (N_8231,N_3768,N_4554);
xnor U8232 (N_8232,N_5810,N_4371);
nor U8233 (N_8233,N_3585,N_5401);
nand U8234 (N_8234,N_3418,N_3819);
nand U8235 (N_8235,N_5478,N_5291);
or U8236 (N_8236,N_4528,N_4675);
xor U8237 (N_8237,N_4936,N_5756);
nor U8238 (N_8238,N_4358,N_3916);
and U8239 (N_8239,N_5292,N_3729);
xnor U8240 (N_8240,N_4215,N_3044);
nor U8241 (N_8241,N_4940,N_3176);
xnor U8242 (N_8242,N_4205,N_3385);
xnor U8243 (N_8243,N_5523,N_5396);
nor U8244 (N_8244,N_4348,N_3402);
and U8245 (N_8245,N_4691,N_4269);
or U8246 (N_8246,N_4471,N_3876);
or U8247 (N_8247,N_4463,N_3511);
nor U8248 (N_8248,N_5746,N_3629);
and U8249 (N_8249,N_4076,N_3313);
nand U8250 (N_8250,N_4787,N_3069);
nor U8251 (N_8251,N_3244,N_3817);
and U8252 (N_8252,N_5477,N_4303);
nand U8253 (N_8253,N_4388,N_3564);
nor U8254 (N_8254,N_3878,N_4846);
xor U8255 (N_8255,N_5283,N_3646);
xnor U8256 (N_8256,N_4743,N_4361);
and U8257 (N_8257,N_3085,N_4565);
or U8258 (N_8258,N_4984,N_3201);
or U8259 (N_8259,N_5577,N_3951);
and U8260 (N_8260,N_3260,N_4956);
xnor U8261 (N_8261,N_4198,N_3808);
and U8262 (N_8262,N_4917,N_3269);
nor U8263 (N_8263,N_3192,N_4229);
and U8264 (N_8264,N_4085,N_3441);
nand U8265 (N_8265,N_3889,N_3146);
nand U8266 (N_8266,N_3777,N_5635);
and U8267 (N_8267,N_4274,N_4979);
or U8268 (N_8268,N_5921,N_4878);
nor U8269 (N_8269,N_4183,N_3593);
nand U8270 (N_8270,N_4466,N_5298);
and U8271 (N_8271,N_4106,N_5903);
and U8272 (N_8272,N_5394,N_5508);
and U8273 (N_8273,N_3114,N_3012);
xnor U8274 (N_8274,N_4888,N_3086);
nand U8275 (N_8275,N_3490,N_4266);
nand U8276 (N_8276,N_4340,N_4590);
and U8277 (N_8277,N_3335,N_4873);
xor U8278 (N_8278,N_5344,N_3596);
or U8279 (N_8279,N_4276,N_5299);
xnor U8280 (N_8280,N_5640,N_5833);
or U8281 (N_8281,N_5142,N_4066);
and U8282 (N_8282,N_4507,N_3959);
and U8283 (N_8283,N_4963,N_4205);
nand U8284 (N_8284,N_4625,N_4603);
or U8285 (N_8285,N_4116,N_4351);
xor U8286 (N_8286,N_5075,N_4595);
nand U8287 (N_8287,N_4374,N_4247);
xnor U8288 (N_8288,N_5119,N_4690);
xor U8289 (N_8289,N_3097,N_4997);
xor U8290 (N_8290,N_3515,N_4903);
nor U8291 (N_8291,N_5818,N_5160);
nor U8292 (N_8292,N_5549,N_4310);
or U8293 (N_8293,N_5592,N_4863);
nand U8294 (N_8294,N_4849,N_3471);
or U8295 (N_8295,N_5977,N_5026);
or U8296 (N_8296,N_3582,N_4765);
nand U8297 (N_8297,N_5197,N_3171);
nor U8298 (N_8298,N_4441,N_4541);
or U8299 (N_8299,N_5838,N_5569);
xnor U8300 (N_8300,N_4932,N_5810);
nor U8301 (N_8301,N_5070,N_4910);
or U8302 (N_8302,N_3922,N_3986);
or U8303 (N_8303,N_5789,N_3178);
or U8304 (N_8304,N_3125,N_5703);
or U8305 (N_8305,N_5438,N_4255);
and U8306 (N_8306,N_3854,N_3699);
nand U8307 (N_8307,N_4297,N_5551);
xnor U8308 (N_8308,N_3558,N_4291);
or U8309 (N_8309,N_4236,N_4769);
and U8310 (N_8310,N_5930,N_5812);
or U8311 (N_8311,N_3453,N_4877);
and U8312 (N_8312,N_3581,N_5060);
and U8313 (N_8313,N_3616,N_5524);
and U8314 (N_8314,N_5505,N_3183);
or U8315 (N_8315,N_3903,N_4915);
and U8316 (N_8316,N_5142,N_3867);
and U8317 (N_8317,N_5201,N_4308);
nor U8318 (N_8318,N_5456,N_4967);
and U8319 (N_8319,N_5035,N_3186);
xnor U8320 (N_8320,N_5089,N_3618);
and U8321 (N_8321,N_3929,N_3045);
and U8322 (N_8322,N_5543,N_4554);
xnor U8323 (N_8323,N_5825,N_5125);
nor U8324 (N_8324,N_4835,N_3553);
or U8325 (N_8325,N_5401,N_5370);
nor U8326 (N_8326,N_3559,N_5607);
or U8327 (N_8327,N_5749,N_3260);
nor U8328 (N_8328,N_3721,N_3540);
xnor U8329 (N_8329,N_5923,N_4832);
xnor U8330 (N_8330,N_5056,N_4251);
nand U8331 (N_8331,N_3530,N_3241);
xnor U8332 (N_8332,N_3127,N_5797);
xnor U8333 (N_8333,N_5389,N_3135);
or U8334 (N_8334,N_4877,N_3715);
nand U8335 (N_8335,N_5633,N_3752);
xnor U8336 (N_8336,N_3708,N_3615);
nor U8337 (N_8337,N_3680,N_4832);
nor U8338 (N_8338,N_4333,N_4427);
xor U8339 (N_8339,N_4872,N_3465);
nand U8340 (N_8340,N_3799,N_4141);
xnor U8341 (N_8341,N_5594,N_4706);
xnor U8342 (N_8342,N_3944,N_3613);
or U8343 (N_8343,N_4146,N_5272);
nor U8344 (N_8344,N_5922,N_4046);
xnor U8345 (N_8345,N_4157,N_3448);
nor U8346 (N_8346,N_5343,N_5186);
or U8347 (N_8347,N_4838,N_4088);
and U8348 (N_8348,N_5944,N_5438);
xor U8349 (N_8349,N_5969,N_3666);
or U8350 (N_8350,N_5187,N_4942);
and U8351 (N_8351,N_3249,N_3343);
nor U8352 (N_8352,N_5520,N_5926);
or U8353 (N_8353,N_4398,N_5526);
xor U8354 (N_8354,N_4780,N_3373);
xnor U8355 (N_8355,N_4983,N_5712);
nor U8356 (N_8356,N_5319,N_5486);
xnor U8357 (N_8357,N_3494,N_4715);
xnor U8358 (N_8358,N_5693,N_3594);
xnor U8359 (N_8359,N_4976,N_5633);
nor U8360 (N_8360,N_5762,N_4771);
xnor U8361 (N_8361,N_3214,N_3520);
and U8362 (N_8362,N_5906,N_3407);
nand U8363 (N_8363,N_3776,N_3601);
nand U8364 (N_8364,N_3782,N_5731);
or U8365 (N_8365,N_4454,N_3414);
or U8366 (N_8366,N_3167,N_5319);
xor U8367 (N_8367,N_5765,N_3696);
xnor U8368 (N_8368,N_4713,N_5038);
xnor U8369 (N_8369,N_4221,N_3225);
nor U8370 (N_8370,N_4704,N_5010);
and U8371 (N_8371,N_5043,N_5871);
xnor U8372 (N_8372,N_3059,N_4463);
xnor U8373 (N_8373,N_4945,N_5190);
nand U8374 (N_8374,N_4339,N_5652);
nor U8375 (N_8375,N_5991,N_5220);
xnor U8376 (N_8376,N_5963,N_3481);
xor U8377 (N_8377,N_5893,N_3041);
nand U8378 (N_8378,N_5382,N_4011);
or U8379 (N_8379,N_3917,N_3650);
and U8380 (N_8380,N_5856,N_4177);
and U8381 (N_8381,N_5979,N_5421);
nor U8382 (N_8382,N_4417,N_4889);
xor U8383 (N_8383,N_4865,N_5388);
and U8384 (N_8384,N_3322,N_5615);
xor U8385 (N_8385,N_5761,N_4064);
and U8386 (N_8386,N_5989,N_3159);
xor U8387 (N_8387,N_4795,N_5171);
nand U8388 (N_8388,N_3890,N_4729);
and U8389 (N_8389,N_3717,N_3981);
nand U8390 (N_8390,N_4452,N_5945);
nor U8391 (N_8391,N_4653,N_3047);
nor U8392 (N_8392,N_5213,N_4731);
nand U8393 (N_8393,N_5177,N_5592);
nand U8394 (N_8394,N_3213,N_5350);
xor U8395 (N_8395,N_3114,N_3584);
and U8396 (N_8396,N_5590,N_5411);
nor U8397 (N_8397,N_3849,N_4342);
and U8398 (N_8398,N_5206,N_4826);
nand U8399 (N_8399,N_4429,N_5297);
nor U8400 (N_8400,N_3771,N_4043);
nor U8401 (N_8401,N_3268,N_4674);
and U8402 (N_8402,N_5668,N_4328);
and U8403 (N_8403,N_5157,N_5390);
xor U8404 (N_8404,N_3892,N_4414);
nor U8405 (N_8405,N_3838,N_4861);
xor U8406 (N_8406,N_5342,N_5325);
or U8407 (N_8407,N_4944,N_3913);
nand U8408 (N_8408,N_3332,N_3261);
and U8409 (N_8409,N_5289,N_4630);
nand U8410 (N_8410,N_5401,N_5321);
nand U8411 (N_8411,N_4976,N_4978);
nor U8412 (N_8412,N_4548,N_5888);
nand U8413 (N_8413,N_5157,N_4130);
nor U8414 (N_8414,N_5681,N_4114);
or U8415 (N_8415,N_4213,N_3567);
xor U8416 (N_8416,N_4834,N_4646);
nor U8417 (N_8417,N_4674,N_5830);
nor U8418 (N_8418,N_5980,N_4278);
nand U8419 (N_8419,N_4821,N_3807);
nand U8420 (N_8420,N_3011,N_3093);
xnor U8421 (N_8421,N_4860,N_3015);
nor U8422 (N_8422,N_3211,N_4553);
xnor U8423 (N_8423,N_3139,N_3661);
or U8424 (N_8424,N_5439,N_3435);
nor U8425 (N_8425,N_4774,N_3629);
nor U8426 (N_8426,N_3914,N_5019);
xor U8427 (N_8427,N_4912,N_5219);
nor U8428 (N_8428,N_3513,N_5566);
or U8429 (N_8429,N_5217,N_4749);
nand U8430 (N_8430,N_3984,N_5906);
and U8431 (N_8431,N_3686,N_4749);
or U8432 (N_8432,N_5153,N_4707);
xor U8433 (N_8433,N_4726,N_5519);
and U8434 (N_8434,N_3982,N_4050);
and U8435 (N_8435,N_3765,N_3347);
and U8436 (N_8436,N_5022,N_3479);
nand U8437 (N_8437,N_4710,N_4199);
nor U8438 (N_8438,N_3096,N_3114);
or U8439 (N_8439,N_4830,N_3907);
nor U8440 (N_8440,N_4968,N_3954);
nor U8441 (N_8441,N_4201,N_4334);
and U8442 (N_8442,N_3621,N_3737);
and U8443 (N_8443,N_4742,N_4300);
xor U8444 (N_8444,N_5166,N_5963);
xnor U8445 (N_8445,N_5862,N_5219);
or U8446 (N_8446,N_3750,N_5078);
or U8447 (N_8447,N_5152,N_5055);
nand U8448 (N_8448,N_4709,N_4361);
nand U8449 (N_8449,N_5873,N_4597);
and U8450 (N_8450,N_4331,N_5802);
xor U8451 (N_8451,N_4151,N_4075);
or U8452 (N_8452,N_3635,N_4084);
xor U8453 (N_8453,N_4358,N_3364);
xnor U8454 (N_8454,N_5972,N_3171);
nand U8455 (N_8455,N_4741,N_5316);
nor U8456 (N_8456,N_5592,N_5064);
xnor U8457 (N_8457,N_4718,N_3140);
and U8458 (N_8458,N_4842,N_3981);
and U8459 (N_8459,N_5198,N_5573);
or U8460 (N_8460,N_3860,N_3760);
nand U8461 (N_8461,N_4046,N_4324);
and U8462 (N_8462,N_4904,N_3797);
nand U8463 (N_8463,N_4850,N_4787);
nand U8464 (N_8464,N_3899,N_5823);
or U8465 (N_8465,N_5513,N_3192);
nand U8466 (N_8466,N_3423,N_3879);
xnor U8467 (N_8467,N_5236,N_4321);
or U8468 (N_8468,N_3083,N_5117);
or U8469 (N_8469,N_3164,N_4661);
xor U8470 (N_8470,N_5272,N_4900);
nand U8471 (N_8471,N_3585,N_5725);
nor U8472 (N_8472,N_3699,N_4727);
nor U8473 (N_8473,N_5936,N_5749);
or U8474 (N_8474,N_4421,N_5014);
or U8475 (N_8475,N_5354,N_4379);
nor U8476 (N_8476,N_5935,N_4009);
or U8477 (N_8477,N_5705,N_5618);
nor U8478 (N_8478,N_5488,N_4643);
and U8479 (N_8479,N_5419,N_3108);
or U8480 (N_8480,N_3880,N_5427);
nor U8481 (N_8481,N_4651,N_4863);
or U8482 (N_8482,N_5552,N_5220);
or U8483 (N_8483,N_4248,N_5252);
and U8484 (N_8484,N_4365,N_3851);
nor U8485 (N_8485,N_5895,N_4165);
and U8486 (N_8486,N_4202,N_3684);
and U8487 (N_8487,N_5995,N_5661);
nand U8488 (N_8488,N_3253,N_4115);
and U8489 (N_8489,N_4075,N_5115);
and U8490 (N_8490,N_4614,N_5778);
or U8491 (N_8491,N_5012,N_3530);
and U8492 (N_8492,N_3959,N_3900);
or U8493 (N_8493,N_3466,N_4979);
or U8494 (N_8494,N_5603,N_4110);
nor U8495 (N_8495,N_4826,N_5108);
nand U8496 (N_8496,N_3710,N_3931);
xor U8497 (N_8497,N_4886,N_5883);
nand U8498 (N_8498,N_5788,N_4989);
xnor U8499 (N_8499,N_3879,N_3478);
or U8500 (N_8500,N_3065,N_4609);
or U8501 (N_8501,N_5655,N_4992);
xnor U8502 (N_8502,N_4368,N_5751);
and U8503 (N_8503,N_5030,N_3832);
xor U8504 (N_8504,N_5227,N_5399);
xnor U8505 (N_8505,N_3722,N_4609);
xnor U8506 (N_8506,N_5612,N_3932);
nor U8507 (N_8507,N_5508,N_4984);
xor U8508 (N_8508,N_5920,N_3318);
or U8509 (N_8509,N_4010,N_5058);
or U8510 (N_8510,N_4816,N_3491);
nand U8511 (N_8511,N_4686,N_3771);
xor U8512 (N_8512,N_3116,N_3567);
xor U8513 (N_8513,N_5128,N_5427);
nand U8514 (N_8514,N_4035,N_5048);
and U8515 (N_8515,N_4460,N_4117);
nor U8516 (N_8516,N_4764,N_3076);
xnor U8517 (N_8517,N_4529,N_5301);
and U8518 (N_8518,N_3783,N_5798);
nor U8519 (N_8519,N_4276,N_3867);
or U8520 (N_8520,N_4110,N_3082);
nand U8521 (N_8521,N_4075,N_4780);
and U8522 (N_8522,N_4888,N_3468);
nor U8523 (N_8523,N_3335,N_5886);
and U8524 (N_8524,N_4881,N_5225);
xor U8525 (N_8525,N_3162,N_5665);
xnor U8526 (N_8526,N_5071,N_5443);
or U8527 (N_8527,N_3871,N_3717);
nor U8528 (N_8528,N_5966,N_5114);
nor U8529 (N_8529,N_3724,N_5529);
nor U8530 (N_8530,N_3791,N_3505);
nand U8531 (N_8531,N_5203,N_3377);
or U8532 (N_8532,N_3852,N_4933);
nor U8533 (N_8533,N_3278,N_3750);
or U8534 (N_8534,N_4497,N_4141);
nor U8535 (N_8535,N_3650,N_4186);
nand U8536 (N_8536,N_4530,N_3970);
nand U8537 (N_8537,N_5496,N_5737);
xor U8538 (N_8538,N_3250,N_5070);
nor U8539 (N_8539,N_5654,N_5150);
xnor U8540 (N_8540,N_4951,N_3194);
xnor U8541 (N_8541,N_3421,N_4291);
xnor U8542 (N_8542,N_5587,N_3101);
or U8543 (N_8543,N_3687,N_5152);
and U8544 (N_8544,N_5824,N_3573);
nand U8545 (N_8545,N_4810,N_5727);
xor U8546 (N_8546,N_4904,N_3610);
nand U8547 (N_8547,N_4096,N_5140);
and U8548 (N_8548,N_5582,N_3464);
nand U8549 (N_8549,N_3993,N_4974);
and U8550 (N_8550,N_5873,N_3223);
xor U8551 (N_8551,N_4351,N_3785);
and U8552 (N_8552,N_5412,N_4994);
xor U8553 (N_8553,N_4418,N_5169);
or U8554 (N_8554,N_4278,N_3044);
nand U8555 (N_8555,N_5359,N_5903);
nor U8556 (N_8556,N_4565,N_3372);
or U8557 (N_8557,N_3912,N_3298);
nand U8558 (N_8558,N_4611,N_4413);
or U8559 (N_8559,N_4476,N_5426);
nor U8560 (N_8560,N_5285,N_4878);
and U8561 (N_8561,N_3080,N_5256);
xnor U8562 (N_8562,N_5227,N_3430);
xor U8563 (N_8563,N_3772,N_5874);
xor U8564 (N_8564,N_4226,N_4615);
xnor U8565 (N_8565,N_4359,N_3078);
xor U8566 (N_8566,N_5578,N_3700);
or U8567 (N_8567,N_4685,N_4750);
xor U8568 (N_8568,N_3612,N_3801);
or U8569 (N_8569,N_3245,N_5537);
nand U8570 (N_8570,N_5363,N_4091);
nor U8571 (N_8571,N_5801,N_5329);
xnor U8572 (N_8572,N_4399,N_5130);
or U8573 (N_8573,N_4581,N_5312);
and U8574 (N_8574,N_4967,N_4712);
and U8575 (N_8575,N_3647,N_4793);
xor U8576 (N_8576,N_4672,N_3710);
and U8577 (N_8577,N_3276,N_4579);
xnor U8578 (N_8578,N_4833,N_4044);
nand U8579 (N_8579,N_4993,N_5177);
nand U8580 (N_8580,N_5691,N_4388);
nand U8581 (N_8581,N_5461,N_4514);
xnor U8582 (N_8582,N_5100,N_4721);
or U8583 (N_8583,N_3646,N_5152);
nand U8584 (N_8584,N_3069,N_4902);
or U8585 (N_8585,N_5886,N_3593);
nand U8586 (N_8586,N_4469,N_3037);
and U8587 (N_8587,N_3272,N_5976);
nand U8588 (N_8588,N_4721,N_5592);
and U8589 (N_8589,N_4787,N_5756);
nand U8590 (N_8590,N_3213,N_4147);
or U8591 (N_8591,N_3231,N_4680);
nor U8592 (N_8592,N_4813,N_3070);
nand U8593 (N_8593,N_3411,N_5379);
nand U8594 (N_8594,N_4471,N_3971);
nand U8595 (N_8595,N_3492,N_3565);
or U8596 (N_8596,N_4414,N_3569);
and U8597 (N_8597,N_4055,N_5069);
or U8598 (N_8598,N_4522,N_5049);
xor U8599 (N_8599,N_4308,N_3649);
and U8600 (N_8600,N_3234,N_5029);
xnor U8601 (N_8601,N_3989,N_5985);
and U8602 (N_8602,N_3324,N_5164);
nand U8603 (N_8603,N_4849,N_4393);
xnor U8604 (N_8604,N_3272,N_5143);
and U8605 (N_8605,N_4959,N_3174);
or U8606 (N_8606,N_5443,N_5196);
and U8607 (N_8607,N_4486,N_3962);
and U8608 (N_8608,N_4374,N_5266);
or U8609 (N_8609,N_5563,N_5275);
nand U8610 (N_8610,N_5844,N_3430);
nor U8611 (N_8611,N_5272,N_4620);
nor U8612 (N_8612,N_4821,N_4360);
or U8613 (N_8613,N_4589,N_5293);
and U8614 (N_8614,N_3382,N_3387);
xnor U8615 (N_8615,N_4333,N_4419);
nand U8616 (N_8616,N_5684,N_3785);
nand U8617 (N_8617,N_5122,N_4171);
or U8618 (N_8618,N_4578,N_3968);
xor U8619 (N_8619,N_5060,N_3696);
xor U8620 (N_8620,N_4635,N_3014);
nand U8621 (N_8621,N_4779,N_4931);
or U8622 (N_8622,N_3057,N_5953);
and U8623 (N_8623,N_5221,N_3151);
or U8624 (N_8624,N_3126,N_4638);
nor U8625 (N_8625,N_4978,N_3314);
nand U8626 (N_8626,N_4932,N_3950);
and U8627 (N_8627,N_4296,N_5581);
and U8628 (N_8628,N_3678,N_5722);
nor U8629 (N_8629,N_4886,N_4397);
nor U8630 (N_8630,N_3348,N_5494);
or U8631 (N_8631,N_3337,N_4942);
nand U8632 (N_8632,N_5653,N_3437);
or U8633 (N_8633,N_4269,N_3474);
nor U8634 (N_8634,N_3727,N_3135);
xor U8635 (N_8635,N_3179,N_4536);
nand U8636 (N_8636,N_4399,N_3821);
and U8637 (N_8637,N_5925,N_4190);
xor U8638 (N_8638,N_3216,N_3214);
xor U8639 (N_8639,N_4434,N_4510);
and U8640 (N_8640,N_3294,N_4641);
nand U8641 (N_8641,N_4699,N_4668);
xor U8642 (N_8642,N_3023,N_4938);
xnor U8643 (N_8643,N_3234,N_3728);
and U8644 (N_8644,N_3456,N_4715);
and U8645 (N_8645,N_5135,N_4320);
nor U8646 (N_8646,N_5589,N_4887);
or U8647 (N_8647,N_4652,N_3960);
nand U8648 (N_8648,N_5161,N_5299);
nor U8649 (N_8649,N_3449,N_5627);
or U8650 (N_8650,N_5833,N_3042);
nor U8651 (N_8651,N_4874,N_5571);
xor U8652 (N_8652,N_4339,N_5070);
nand U8653 (N_8653,N_3483,N_3440);
and U8654 (N_8654,N_5605,N_3519);
and U8655 (N_8655,N_4965,N_5953);
nor U8656 (N_8656,N_4298,N_3954);
xor U8657 (N_8657,N_3929,N_5820);
nor U8658 (N_8658,N_4310,N_5194);
xor U8659 (N_8659,N_4916,N_3062);
or U8660 (N_8660,N_5071,N_4061);
and U8661 (N_8661,N_5504,N_3701);
xnor U8662 (N_8662,N_4087,N_4343);
and U8663 (N_8663,N_5982,N_4639);
nand U8664 (N_8664,N_4303,N_3803);
or U8665 (N_8665,N_4948,N_3683);
and U8666 (N_8666,N_5101,N_4333);
and U8667 (N_8667,N_5300,N_3610);
and U8668 (N_8668,N_4203,N_3907);
nand U8669 (N_8669,N_4240,N_3709);
xnor U8670 (N_8670,N_5668,N_4781);
and U8671 (N_8671,N_3775,N_5987);
nand U8672 (N_8672,N_5909,N_5814);
nand U8673 (N_8673,N_5820,N_5148);
nand U8674 (N_8674,N_4047,N_3862);
or U8675 (N_8675,N_5694,N_3309);
and U8676 (N_8676,N_4189,N_5796);
or U8677 (N_8677,N_5119,N_3296);
xor U8678 (N_8678,N_5950,N_4030);
nand U8679 (N_8679,N_3493,N_4334);
and U8680 (N_8680,N_4530,N_4718);
and U8681 (N_8681,N_3458,N_5699);
or U8682 (N_8682,N_5590,N_4954);
nor U8683 (N_8683,N_4803,N_5395);
nand U8684 (N_8684,N_5817,N_3294);
nand U8685 (N_8685,N_3424,N_4476);
nor U8686 (N_8686,N_5237,N_5634);
xnor U8687 (N_8687,N_4151,N_3338);
nor U8688 (N_8688,N_4867,N_4999);
xor U8689 (N_8689,N_3293,N_4226);
and U8690 (N_8690,N_5360,N_5533);
xnor U8691 (N_8691,N_3295,N_3525);
xor U8692 (N_8692,N_3848,N_3098);
nor U8693 (N_8693,N_5698,N_5454);
or U8694 (N_8694,N_3237,N_5826);
nand U8695 (N_8695,N_5449,N_4259);
xor U8696 (N_8696,N_4937,N_4754);
nor U8697 (N_8697,N_5346,N_5432);
nand U8698 (N_8698,N_3484,N_5552);
xnor U8699 (N_8699,N_5283,N_5518);
nor U8700 (N_8700,N_4065,N_4205);
nand U8701 (N_8701,N_4570,N_3105);
nand U8702 (N_8702,N_5928,N_4798);
and U8703 (N_8703,N_5385,N_4388);
nor U8704 (N_8704,N_3163,N_5736);
xor U8705 (N_8705,N_3386,N_4336);
xor U8706 (N_8706,N_5912,N_5404);
nor U8707 (N_8707,N_3116,N_4977);
nor U8708 (N_8708,N_3575,N_3184);
and U8709 (N_8709,N_3520,N_4479);
xor U8710 (N_8710,N_4329,N_5947);
or U8711 (N_8711,N_3578,N_3060);
nor U8712 (N_8712,N_3559,N_3627);
nor U8713 (N_8713,N_3011,N_4369);
nand U8714 (N_8714,N_4060,N_5150);
xnor U8715 (N_8715,N_4503,N_3253);
nand U8716 (N_8716,N_5871,N_3311);
nand U8717 (N_8717,N_3204,N_4433);
nor U8718 (N_8718,N_5505,N_3421);
and U8719 (N_8719,N_4316,N_5744);
xor U8720 (N_8720,N_5858,N_5836);
and U8721 (N_8721,N_5032,N_5921);
nand U8722 (N_8722,N_4217,N_5611);
nand U8723 (N_8723,N_4502,N_4258);
xnor U8724 (N_8724,N_5583,N_5752);
xor U8725 (N_8725,N_4104,N_5749);
xor U8726 (N_8726,N_3590,N_5580);
or U8727 (N_8727,N_3829,N_3281);
or U8728 (N_8728,N_5870,N_5505);
and U8729 (N_8729,N_3808,N_3950);
or U8730 (N_8730,N_5965,N_3944);
xnor U8731 (N_8731,N_4777,N_3077);
xnor U8732 (N_8732,N_5968,N_5072);
xor U8733 (N_8733,N_5652,N_3704);
nor U8734 (N_8734,N_4559,N_4909);
and U8735 (N_8735,N_4105,N_3153);
xnor U8736 (N_8736,N_4519,N_3661);
nand U8737 (N_8737,N_3020,N_4324);
or U8738 (N_8738,N_5609,N_4988);
nor U8739 (N_8739,N_5241,N_4656);
and U8740 (N_8740,N_5618,N_4018);
and U8741 (N_8741,N_3749,N_5976);
nor U8742 (N_8742,N_3126,N_5259);
or U8743 (N_8743,N_4182,N_3979);
xor U8744 (N_8744,N_3011,N_5778);
and U8745 (N_8745,N_3989,N_5908);
or U8746 (N_8746,N_4926,N_4373);
xnor U8747 (N_8747,N_4282,N_3572);
xor U8748 (N_8748,N_4444,N_3833);
and U8749 (N_8749,N_5336,N_3406);
and U8750 (N_8750,N_3514,N_5331);
or U8751 (N_8751,N_5537,N_4184);
or U8752 (N_8752,N_5686,N_5470);
nor U8753 (N_8753,N_4499,N_5821);
nor U8754 (N_8754,N_4863,N_3108);
nor U8755 (N_8755,N_5151,N_3071);
nand U8756 (N_8756,N_5423,N_3053);
or U8757 (N_8757,N_5143,N_3747);
nor U8758 (N_8758,N_4412,N_3893);
nor U8759 (N_8759,N_3499,N_4965);
and U8760 (N_8760,N_5553,N_5260);
and U8761 (N_8761,N_3175,N_5592);
nor U8762 (N_8762,N_3270,N_4395);
xor U8763 (N_8763,N_4180,N_4672);
nand U8764 (N_8764,N_5328,N_5302);
or U8765 (N_8765,N_4674,N_4237);
or U8766 (N_8766,N_3026,N_4300);
xnor U8767 (N_8767,N_5824,N_3039);
and U8768 (N_8768,N_4611,N_5630);
or U8769 (N_8769,N_3437,N_5790);
nor U8770 (N_8770,N_5415,N_5501);
xor U8771 (N_8771,N_4589,N_5854);
or U8772 (N_8772,N_5698,N_5233);
xnor U8773 (N_8773,N_4005,N_4472);
nor U8774 (N_8774,N_3979,N_3632);
or U8775 (N_8775,N_3235,N_5678);
and U8776 (N_8776,N_3549,N_4020);
nor U8777 (N_8777,N_3025,N_5382);
and U8778 (N_8778,N_3147,N_5747);
or U8779 (N_8779,N_3318,N_3558);
xor U8780 (N_8780,N_4936,N_5157);
xnor U8781 (N_8781,N_5096,N_4808);
or U8782 (N_8782,N_3797,N_5142);
nor U8783 (N_8783,N_3800,N_5115);
or U8784 (N_8784,N_5174,N_3227);
or U8785 (N_8785,N_4707,N_3904);
nor U8786 (N_8786,N_3202,N_5722);
or U8787 (N_8787,N_3738,N_5121);
and U8788 (N_8788,N_3567,N_3429);
nand U8789 (N_8789,N_3437,N_5089);
nor U8790 (N_8790,N_4926,N_3885);
xor U8791 (N_8791,N_4857,N_4087);
and U8792 (N_8792,N_4373,N_5040);
nor U8793 (N_8793,N_5421,N_3320);
or U8794 (N_8794,N_3621,N_3412);
xor U8795 (N_8795,N_5497,N_5476);
or U8796 (N_8796,N_4023,N_3881);
or U8797 (N_8797,N_5105,N_5355);
nor U8798 (N_8798,N_4219,N_4116);
nor U8799 (N_8799,N_4506,N_3204);
nor U8800 (N_8800,N_4384,N_5442);
or U8801 (N_8801,N_3882,N_3562);
and U8802 (N_8802,N_5859,N_3656);
xor U8803 (N_8803,N_4686,N_3190);
xnor U8804 (N_8804,N_3891,N_5942);
and U8805 (N_8805,N_5715,N_3982);
or U8806 (N_8806,N_5374,N_3847);
xnor U8807 (N_8807,N_5176,N_4575);
or U8808 (N_8808,N_5471,N_5800);
nand U8809 (N_8809,N_3445,N_4316);
nand U8810 (N_8810,N_4557,N_4890);
xor U8811 (N_8811,N_5817,N_4013);
and U8812 (N_8812,N_3459,N_4792);
and U8813 (N_8813,N_5071,N_5445);
nand U8814 (N_8814,N_4131,N_4713);
xor U8815 (N_8815,N_5260,N_5979);
xnor U8816 (N_8816,N_4396,N_4704);
xor U8817 (N_8817,N_4551,N_3215);
nor U8818 (N_8818,N_4365,N_4547);
or U8819 (N_8819,N_3576,N_4086);
or U8820 (N_8820,N_5772,N_5298);
and U8821 (N_8821,N_4194,N_5358);
xnor U8822 (N_8822,N_5534,N_3334);
nand U8823 (N_8823,N_3574,N_4399);
xnor U8824 (N_8824,N_5619,N_5715);
xor U8825 (N_8825,N_3350,N_5696);
nor U8826 (N_8826,N_4048,N_4264);
nor U8827 (N_8827,N_5864,N_3809);
nor U8828 (N_8828,N_4619,N_5585);
and U8829 (N_8829,N_5518,N_5595);
or U8830 (N_8830,N_3111,N_4716);
and U8831 (N_8831,N_4256,N_3890);
or U8832 (N_8832,N_4249,N_4311);
or U8833 (N_8833,N_4955,N_4141);
xor U8834 (N_8834,N_3879,N_3441);
xor U8835 (N_8835,N_4125,N_5366);
nand U8836 (N_8836,N_5548,N_5339);
and U8837 (N_8837,N_3662,N_4548);
xnor U8838 (N_8838,N_5634,N_5567);
nand U8839 (N_8839,N_3890,N_5612);
nor U8840 (N_8840,N_4948,N_4534);
and U8841 (N_8841,N_4798,N_3650);
and U8842 (N_8842,N_3460,N_4957);
nand U8843 (N_8843,N_4467,N_4945);
xor U8844 (N_8844,N_3143,N_4325);
nor U8845 (N_8845,N_3400,N_4194);
xor U8846 (N_8846,N_3464,N_5540);
xor U8847 (N_8847,N_4037,N_4467);
xnor U8848 (N_8848,N_5850,N_5181);
xor U8849 (N_8849,N_5470,N_3804);
xnor U8850 (N_8850,N_4736,N_3232);
xnor U8851 (N_8851,N_4869,N_5859);
and U8852 (N_8852,N_4279,N_5579);
xor U8853 (N_8853,N_4963,N_5509);
or U8854 (N_8854,N_5992,N_3079);
and U8855 (N_8855,N_4454,N_4928);
nand U8856 (N_8856,N_3037,N_3918);
xor U8857 (N_8857,N_3129,N_5797);
nand U8858 (N_8858,N_5037,N_3805);
xor U8859 (N_8859,N_3092,N_4215);
nor U8860 (N_8860,N_5362,N_5707);
and U8861 (N_8861,N_3010,N_3577);
xnor U8862 (N_8862,N_4966,N_5628);
nor U8863 (N_8863,N_4423,N_3220);
and U8864 (N_8864,N_3700,N_3968);
nor U8865 (N_8865,N_4773,N_3151);
and U8866 (N_8866,N_4211,N_5933);
or U8867 (N_8867,N_4972,N_3174);
nand U8868 (N_8868,N_4886,N_4634);
xnor U8869 (N_8869,N_3418,N_4950);
and U8870 (N_8870,N_4214,N_5791);
xnor U8871 (N_8871,N_5405,N_4523);
nand U8872 (N_8872,N_5952,N_5151);
nand U8873 (N_8873,N_5676,N_3478);
and U8874 (N_8874,N_3831,N_3685);
and U8875 (N_8875,N_5161,N_3356);
and U8876 (N_8876,N_3858,N_4592);
nand U8877 (N_8877,N_3743,N_5928);
nand U8878 (N_8878,N_3494,N_3977);
or U8879 (N_8879,N_4170,N_5065);
or U8880 (N_8880,N_4547,N_5982);
nor U8881 (N_8881,N_4229,N_5626);
nor U8882 (N_8882,N_5019,N_4204);
nor U8883 (N_8883,N_4128,N_4624);
and U8884 (N_8884,N_4107,N_5587);
and U8885 (N_8885,N_5479,N_5730);
xor U8886 (N_8886,N_5580,N_3690);
xnor U8887 (N_8887,N_4234,N_3597);
nor U8888 (N_8888,N_5088,N_3405);
nand U8889 (N_8889,N_4994,N_5900);
xnor U8890 (N_8890,N_5026,N_4335);
or U8891 (N_8891,N_3516,N_5546);
xor U8892 (N_8892,N_4071,N_5588);
nand U8893 (N_8893,N_4764,N_3200);
nand U8894 (N_8894,N_4028,N_5862);
and U8895 (N_8895,N_4385,N_5310);
nor U8896 (N_8896,N_3172,N_5720);
nor U8897 (N_8897,N_4126,N_3098);
xor U8898 (N_8898,N_4233,N_4683);
nand U8899 (N_8899,N_5350,N_4446);
xor U8900 (N_8900,N_3654,N_3037);
xor U8901 (N_8901,N_4976,N_3597);
nor U8902 (N_8902,N_3676,N_5092);
xor U8903 (N_8903,N_5256,N_3093);
and U8904 (N_8904,N_3375,N_3351);
nor U8905 (N_8905,N_5035,N_4441);
or U8906 (N_8906,N_3059,N_4164);
nor U8907 (N_8907,N_5824,N_3865);
nor U8908 (N_8908,N_4021,N_4642);
and U8909 (N_8909,N_5693,N_5497);
xnor U8910 (N_8910,N_3884,N_3006);
nor U8911 (N_8911,N_4686,N_4639);
or U8912 (N_8912,N_5397,N_5387);
nor U8913 (N_8913,N_3500,N_4632);
and U8914 (N_8914,N_3961,N_4204);
or U8915 (N_8915,N_3633,N_4336);
nor U8916 (N_8916,N_4602,N_3104);
nand U8917 (N_8917,N_5620,N_4812);
xnor U8918 (N_8918,N_5427,N_5249);
or U8919 (N_8919,N_4298,N_5358);
and U8920 (N_8920,N_5052,N_3522);
xor U8921 (N_8921,N_3353,N_4763);
nand U8922 (N_8922,N_5319,N_5490);
or U8923 (N_8923,N_5377,N_3799);
nand U8924 (N_8924,N_4720,N_5220);
and U8925 (N_8925,N_4250,N_3106);
nor U8926 (N_8926,N_4840,N_3261);
and U8927 (N_8927,N_3691,N_5218);
and U8928 (N_8928,N_5197,N_5514);
and U8929 (N_8929,N_5562,N_5089);
xor U8930 (N_8930,N_3085,N_5392);
nor U8931 (N_8931,N_3679,N_5502);
nor U8932 (N_8932,N_5932,N_4952);
nand U8933 (N_8933,N_4687,N_3701);
xor U8934 (N_8934,N_3433,N_5891);
and U8935 (N_8935,N_3537,N_4492);
nand U8936 (N_8936,N_5598,N_3070);
nand U8937 (N_8937,N_3900,N_5138);
nand U8938 (N_8938,N_3023,N_4785);
nor U8939 (N_8939,N_4674,N_5701);
and U8940 (N_8940,N_4684,N_4891);
xor U8941 (N_8941,N_5371,N_4939);
nand U8942 (N_8942,N_4706,N_4993);
or U8943 (N_8943,N_3088,N_4828);
nand U8944 (N_8944,N_5565,N_4502);
and U8945 (N_8945,N_5440,N_5304);
nand U8946 (N_8946,N_4774,N_5501);
nor U8947 (N_8947,N_5592,N_5392);
or U8948 (N_8948,N_4527,N_5193);
xor U8949 (N_8949,N_5669,N_5608);
and U8950 (N_8950,N_3903,N_5044);
nor U8951 (N_8951,N_5969,N_3141);
nand U8952 (N_8952,N_5441,N_3294);
or U8953 (N_8953,N_5395,N_3907);
nand U8954 (N_8954,N_5355,N_5853);
nand U8955 (N_8955,N_5832,N_5373);
nor U8956 (N_8956,N_5098,N_3284);
nor U8957 (N_8957,N_4805,N_3052);
and U8958 (N_8958,N_4498,N_4133);
xnor U8959 (N_8959,N_4548,N_4526);
or U8960 (N_8960,N_4527,N_3322);
nor U8961 (N_8961,N_5860,N_4469);
xnor U8962 (N_8962,N_3059,N_3622);
xnor U8963 (N_8963,N_4235,N_5272);
nor U8964 (N_8964,N_3605,N_4220);
nor U8965 (N_8965,N_4715,N_5227);
and U8966 (N_8966,N_5764,N_5177);
or U8967 (N_8967,N_5668,N_3997);
nor U8968 (N_8968,N_5544,N_5215);
xor U8969 (N_8969,N_5357,N_5704);
xnor U8970 (N_8970,N_5211,N_3999);
or U8971 (N_8971,N_5671,N_4173);
nand U8972 (N_8972,N_3064,N_3117);
xor U8973 (N_8973,N_3135,N_5445);
xor U8974 (N_8974,N_5777,N_5853);
nand U8975 (N_8975,N_5635,N_3774);
nand U8976 (N_8976,N_5492,N_4344);
or U8977 (N_8977,N_4109,N_5221);
or U8978 (N_8978,N_3752,N_3598);
or U8979 (N_8979,N_4627,N_5864);
xnor U8980 (N_8980,N_4293,N_3133);
nand U8981 (N_8981,N_4058,N_4290);
or U8982 (N_8982,N_3724,N_4463);
and U8983 (N_8983,N_3953,N_4043);
nand U8984 (N_8984,N_5015,N_4427);
nand U8985 (N_8985,N_5921,N_4973);
or U8986 (N_8986,N_5205,N_5857);
nor U8987 (N_8987,N_4182,N_4929);
nor U8988 (N_8988,N_4009,N_3817);
or U8989 (N_8989,N_3027,N_3409);
and U8990 (N_8990,N_5959,N_3133);
or U8991 (N_8991,N_4749,N_4394);
or U8992 (N_8992,N_5864,N_5464);
xnor U8993 (N_8993,N_5404,N_3160);
nand U8994 (N_8994,N_5827,N_4691);
nand U8995 (N_8995,N_4565,N_4599);
nor U8996 (N_8996,N_3828,N_5676);
and U8997 (N_8997,N_5440,N_4529);
xnor U8998 (N_8998,N_3423,N_3007);
or U8999 (N_8999,N_4157,N_3323);
and U9000 (N_9000,N_8277,N_7819);
or U9001 (N_9001,N_8354,N_7751);
nor U9002 (N_9002,N_6042,N_7344);
xor U9003 (N_9003,N_8875,N_8851);
and U9004 (N_9004,N_8585,N_7120);
or U9005 (N_9005,N_6528,N_7719);
or U9006 (N_9006,N_8809,N_6854);
and U9007 (N_9007,N_7671,N_8428);
or U9008 (N_9008,N_7174,N_8124);
nand U9009 (N_9009,N_8486,N_7706);
nand U9010 (N_9010,N_8186,N_7616);
xnor U9011 (N_9011,N_6776,N_8461);
and U9012 (N_9012,N_8546,N_6541);
nand U9013 (N_9013,N_7721,N_6791);
nor U9014 (N_9014,N_8456,N_7804);
nand U9015 (N_9015,N_7194,N_6437);
nor U9016 (N_9016,N_8121,N_8453);
or U9017 (N_9017,N_7187,N_6342);
xor U9018 (N_9018,N_8781,N_7938);
nand U9019 (N_9019,N_8129,N_8935);
xnor U9020 (N_9020,N_7210,N_8865);
and U9021 (N_9021,N_8949,N_7385);
or U9022 (N_9022,N_7366,N_7716);
nand U9023 (N_9023,N_6045,N_8928);
nor U9024 (N_9024,N_8696,N_8849);
or U9025 (N_9025,N_7907,N_6894);
nand U9026 (N_9026,N_6262,N_6185);
and U9027 (N_9027,N_6521,N_7283);
xor U9028 (N_9028,N_7461,N_7585);
nand U9029 (N_9029,N_7248,N_7891);
nor U9030 (N_9030,N_7323,N_7754);
nor U9031 (N_9031,N_7753,N_6626);
xor U9032 (N_9032,N_8263,N_6194);
or U9033 (N_9033,N_6552,N_6510);
xnor U9034 (N_9034,N_6344,N_6631);
and U9035 (N_9035,N_8424,N_7710);
or U9036 (N_9036,N_7551,N_8688);
or U9037 (N_9037,N_6607,N_6126);
nor U9038 (N_9038,N_7195,N_8429);
and U9039 (N_9039,N_8514,N_8068);
and U9040 (N_9040,N_6880,N_7137);
nand U9041 (N_9041,N_7528,N_8359);
nor U9042 (N_9042,N_7343,N_7578);
or U9043 (N_9043,N_6068,N_8330);
nand U9044 (N_9044,N_8468,N_6432);
nand U9045 (N_9045,N_6079,N_7491);
or U9046 (N_9046,N_6094,N_6622);
nand U9047 (N_9047,N_8582,N_8577);
nand U9048 (N_9048,N_7535,N_8113);
nand U9049 (N_9049,N_6861,N_7342);
nand U9050 (N_9050,N_8058,N_8265);
nor U9051 (N_9051,N_8300,N_8235);
nand U9052 (N_9052,N_7074,N_7552);
xor U9053 (N_9053,N_6551,N_6717);
nor U9054 (N_9054,N_6283,N_8361);
nor U9055 (N_9055,N_8798,N_6041);
nor U9056 (N_9056,N_7138,N_7615);
xor U9057 (N_9057,N_6462,N_6538);
nand U9058 (N_9058,N_8645,N_7212);
and U9059 (N_9059,N_6014,N_6915);
or U9060 (N_9060,N_8387,N_6003);
nor U9061 (N_9061,N_8431,N_7034);
or U9062 (N_9062,N_8727,N_6049);
xnor U9063 (N_9063,N_7944,N_6128);
xnor U9064 (N_9064,N_8139,N_8224);
or U9065 (N_9065,N_6250,N_6269);
and U9066 (N_9066,N_8894,N_6775);
or U9067 (N_9067,N_6946,N_6828);
and U9068 (N_9068,N_8826,N_7401);
and U9069 (N_9069,N_6714,N_6056);
nand U9070 (N_9070,N_8262,N_8906);
and U9071 (N_9071,N_7778,N_8519);
nor U9072 (N_9072,N_7258,N_6173);
nor U9073 (N_9073,N_8377,N_6089);
and U9074 (N_9074,N_8903,N_6325);
nand U9075 (N_9075,N_6756,N_8454);
xnor U9076 (N_9076,N_7843,N_8610);
or U9077 (N_9077,N_6291,N_8286);
xor U9078 (N_9078,N_8169,N_6028);
or U9079 (N_9079,N_7219,N_7260);
or U9080 (N_9080,N_6081,N_6215);
and U9081 (N_9081,N_8627,N_6361);
xor U9082 (N_9082,N_8747,N_6111);
and U9083 (N_9083,N_7699,N_8861);
nor U9084 (N_9084,N_6846,N_6588);
or U9085 (N_9085,N_7169,N_6759);
or U9086 (N_9086,N_7798,N_8685);
xnor U9087 (N_9087,N_6096,N_8467);
xor U9088 (N_9088,N_7351,N_8436);
xor U9089 (N_9089,N_8026,N_7823);
or U9090 (N_9090,N_8481,N_6720);
nand U9091 (N_9091,N_6800,N_7924);
nand U9092 (N_9092,N_6220,N_6282);
and U9093 (N_9093,N_7160,N_7294);
and U9094 (N_9094,N_7732,N_6316);
nor U9095 (N_9095,N_8273,N_6678);
nor U9096 (N_9096,N_8012,N_7129);
and U9097 (N_9097,N_6984,N_7325);
xnor U9098 (N_9098,N_6322,N_8567);
nand U9099 (N_9099,N_8166,N_6178);
xnor U9100 (N_9100,N_6749,N_6696);
or U9101 (N_9101,N_8938,N_7741);
or U9102 (N_9102,N_6442,N_8441);
or U9103 (N_9103,N_8478,N_6172);
and U9104 (N_9104,N_7257,N_8821);
nor U9105 (N_9105,N_7885,N_7613);
xnor U9106 (N_9106,N_8219,N_7322);
and U9107 (N_9107,N_7390,N_7950);
nand U9108 (N_9108,N_7000,N_8516);
nand U9109 (N_9109,N_6304,N_8417);
nor U9110 (N_9110,N_7740,N_7096);
nor U9111 (N_9111,N_8097,N_6149);
and U9112 (N_9112,N_8498,N_6624);
or U9113 (N_9113,N_7456,N_6670);
or U9114 (N_9114,N_6105,N_6928);
nor U9115 (N_9115,N_6779,N_8701);
xor U9116 (N_9116,N_8161,N_6916);
nor U9117 (N_9117,N_8563,N_8140);
and U9118 (N_9118,N_6612,N_6685);
nand U9119 (N_9119,N_6184,N_8187);
or U9120 (N_9120,N_7059,N_6988);
xnor U9121 (N_9121,N_7504,N_6723);
and U9122 (N_9122,N_6176,N_7463);
nand U9123 (N_9123,N_7156,N_6133);
nor U9124 (N_9124,N_7779,N_7735);
and U9125 (N_9125,N_7250,N_7775);
xnor U9126 (N_9126,N_8541,N_6958);
nor U9127 (N_9127,N_8050,N_7596);
or U9128 (N_9128,N_6444,N_7119);
or U9129 (N_9129,N_8116,N_8572);
xor U9130 (N_9130,N_7863,N_8170);
or U9131 (N_9131,N_8176,N_8053);
and U9132 (N_9132,N_8434,N_6054);
or U9133 (N_9133,N_8211,N_7889);
and U9134 (N_9134,N_6117,N_6691);
xor U9135 (N_9135,N_7689,N_8403);
nor U9136 (N_9136,N_6980,N_7302);
and U9137 (N_9137,N_8751,N_6561);
nor U9138 (N_9138,N_7115,N_6877);
or U9139 (N_9139,N_6533,N_6257);
nand U9140 (N_9140,N_6647,N_7972);
xor U9141 (N_9141,N_8643,N_7881);
or U9142 (N_9142,N_7375,N_7291);
nor U9143 (N_9143,N_8279,N_6290);
and U9144 (N_9144,N_8168,N_6968);
or U9145 (N_9145,N_8775,N_6844);
or U9146 (N_9146,N_7886,N_6120);
and U9147 (N_9147,N_7019,N_7705);
nor U9148 (N_9148,N_8379,N_7641);
and U9149 (N_9149,N_6687,N_8332);
nand U9150 (N_9150,N_8126,N_6908);
nand U9151 (N_9151,N_6356,N_8704);
nor U9152 (N_9152,N_7471,N_6926);
nor U9153 (N_9153,N_8762,N_8180);
and U9154 (N_9154,N_8163,N_6137);
nor U9155 (N_9155,N_8684,N_7009);
xnor U9156 (N_9156,N_6256,N_6548);
or U9157 (N_9157,N_8746,N_7029);
xnor U9158 (N_9158,N_8433,N_6506);
nand U9159 (N_9159,N_8096,N_7542);
nor U9160 (N_9160,N_8462,N_7109);
nor U9161 (N_9161,N_8583,N_6884);
nand U9162 (N_9162,N_7842,N_8082);
or U9163 (N_9163,N_7049,N_6627);
and U9164 (N_9164,N_7757,N_6864);
or U9165 (N_9165,N_7444,N_7702);
nand U9166 (N_9166,N_6848,N_8008);
xnor U9167 (N_9167,N_7569,N_7422);
xnor U9168 (N_9168,N_8995,N_7185);
and U9169 (N_9169,N_6298,N_6796);
xor U9170 (N_9170,N_7017,N_7232);
xnor U9171 (N_9171,N_7567,N_7234);
and U9172 (N_9172,N_8934,N_7176);
xor U9173 (N_9173,N_6721,N_8081);
nand U9174 (N_9174,N_8703,N_7799);
and U9175 (N_9175,N_7255,N_8918);
and U9176 (N_9176,N_6944,N_7562);
or U9177 (N_9177,N_8626,N_7420);
xnor U9178 (N_9178,N_8607,N_8349);
nand U9179 (N_9179,N_6722,N_6307);
nand U9180 (N_9180,N_6404,N_7624);
and U9181 (N_9181,N_6431,N_6196);
and U9182 (N_9182,N_7879,N_8063);
nor U9183 (N_9183,N_6684,N_6286);
nor U9184 (N_9184,N_7857,N_6456);
nand U9185 (N_9185,N_8569,N_6330);
nor U9186 (N_9186,N_7155,N_8499);
nor U9187 (N_9187,N_8900,N_7544);
nand U9188 (N_9188,N_6881,N_7594);
and U9189 (N_9189,N_7038,N_7680);
nor U9190 (N_9190,N_8657,N_7559);
and U9191 (N_9191,N_6012,N_7339);
xnor U9192 (N_9192,N_7919,N_7012);
nor U9193 (N_9193,N_6682,N_6353);
or U9194 (N_9194,N_7630,N_6130);
nand U9195 (N_9195,N_7039,N_6156);
nand U9196 (N_9196,N_6376,N_6385);
nor U9197 (N_9197,N_8828,N_7442);
or U9198 (N_9198,N_8641,N_7678);
nand U9199 (N_9199,N_6931,N_6331);
or U9200 (N_9200,N_7600,N_6009);
and U9201 (N_9201,N_7334,N_7411);
or U9202 (N_9202,N_8805,N_8697);
nand U9203 (N_9203,N_6150,N_6859);
or U9204 (N_9204,N_7646,N_8654);
or U9205 (N_9205,N_6950,N_6808);
nor U9206 (N_9206,N_8293,N_8554);
or U9207 (N_9207,N_6228,N_8831);
nand U9208 (N_9208,N_8267,N_7910);
nor U9209 (N_9209,N_6410,N_8590);
nand U9210 (N_9210,N_7618,N_7229);
nor U9211 (N_9211,N_7825,N_6430);
nor U9212 (N_9212,N_6597,N_7217);
or U9213 (N_9213,N_7828,N_8074);
and U9214 (N_9214,N_7902,N_8223);
xor U9215 (N_9215,N_8829,N_6729);
and U9216 (N_9216,N_7536,N_8042);
nor U9217 (N_9217,N_8413,N_6397);
xor U9218 (N_9218,N_6073,N_7146);
nand U9219 (N_9219,N_6428,N_7270);
nor U9220 (N_9220,N_8376,N_7981);
nor U9221 (N_9221,N_6845,N_7966);
or U9222 (N_9222,N_6490,N_8606);
or U9223 (N_9223,N_8717,N_8409);
nand U9224 (N_9224,N_8132,N_6413);
xnor U9225 (N_9225,N_6898,N_6144);
or U9226 (N_9226,N_6033,N_6809);
xor U9227 (N_9227,N_8108,N_8337);
nand U9228 (N_9228,N_6989,N_6666);
and U9229 (N_9229,N_6787,N_8856);
xnor U9230 (N_9230,N_8144,N_8303);
xnor U9231 (N_9231,N_7446,N_7999);
xor U9232 (N_9232,N_7426,N_6708);
nand U9233 (N_9233,N_8877,N_6365);
nand U9234 (N_9234,N_8924,N_7923);
xnor U9235 (N_9235,N_8494,N_7611);
xnor U9236 (N_9236,N_6731,N_7941);
xor U9237 (N_9237,N_6482,N_8886);
and U9238 (N_9238,N_6692,N_6166);
or U9239 (N_9239,N_8155,N_6230);
or U9240 (N_9240,N_7018,N_6399);
and U9241 (N_9241,N_8878,N_7755);
nor U9242 (N_9242,N_7116,N_6467);
nand U9243 (N_9243,N_8043,N_6268);
and U9244 (N_9244,N_7164,N_8987);
and U9245 (N_9245,N_7988,N_6941);
and U9246 (N_9246,N_8317,N_7952);
or U9247 (N_9247,N_7273,N_8771);
and U9248 (N_9248,N_7298,N_7020);
nand U9249 (N_9249,N_6386,N_7769);
and U9250 (N_9250,N_6662,N_8694);
xnor U9251 (N_9251,N_8136,N_6853);
and U9252 (N_9252,N_8037,N_6318);
or U9253 (N_9253,N_7350,N_8782);
or U9254 (N_9254,N_6632,N_7084);
nand U9255 (N_9255,N_6760,N_8619);
or U9256 (N_9256,N_7186,N_7466);
and U9257 (N_9257,N_6486,N_8416);
xnor U9258 (N_9258,N_6942,N_7657);
nand U9259 (N_9259,N_6499,N_7853);
or U9260 (N_9260,N_8573,N_8507);
xor U9261 (N_9261,N_8979,N_7718);
nor U9262 (N_9262,N_7895,N_7868);
nor U9263 (N_9263,N_7897,N_7309);
or U9264 (N_9264,N_7993,N_8713);
nor U9265 (N_9265,N_7336,N_6657);
nor U9266 (N_9266,N_7311,N_7151);
or U9267 (N_9267,N_8017,N_6157);
nand U9268 (N_9268,N_7122,N_7629);
nand U9269 (N_9269,N_7654,N_6636);
and U9270 (N_9270,N_8973,N_6677);
nor U9271 (N_9271,N_6640,N_7113);
and U9272 (N_9272,N_6147,N_6366);
xnor U9273 (N_9273,N_6160,N_6280);
and U9274 (N_9274,N_7381,N_8937);
nand U9275 (N_9275,N_6686,N_7290);
and U9276 (N_9276,N_6887,N_7956);
or U9277 (N_9277,N_7926,N_7335);
or U9278 (N_9278,N_6614,N_8653);
and U9279 (N_9279,N_8274,N_6681);
nor U9280 (N_9280,N_7154,N_6819);
nor U9281 (N_9281,N_6226,N_8051);
and U9282 (N_9282,N_8060,N_6998);
and U9283 (N_9283,N_8913,N_7748);
nand U9284 (N_9284,N_6782,N_7656);
xnor U9285 (N_9285,N_7180,N_6066);
xnor U9286 (N_9286,N_7384,N_8001);
nor U9287 (N_9287,N_7467,N_8493);
nor U9288 (N_9288,N_7098,N_7802);
and U9289 (N_9289,N_6567,N_6971);
and U9290 (N_9290,N_7346,N_8358);
and U9291 (N_9291,N_8339,N_8500);
nor U9292 (N_9292,N_6396,N_8266);
nor U9293 (N_9293,N_6234,N_8272);
xor U9294 (N_9294,N_7231,N_7410);
xor U9295 (N_9295,N_8504,N_8027);
nor U9296 (N_9296,N_7771,N_8908);
xnor U9297 (N_9297,N_7355,N_6812);
xor U9298 (N_9298,N_6159,N_6592);
nor U9299 (N_9299,N_7795,N_7175);
nor U9300 (N_9300,N_6763,N_6106);
nor U9301 (N_9301,N_6907,N_6634);
nand U9302 (N_9302,N_6996,N_8759);
or U9303 (N_9303,N_6453,N_8490);
nand U9304 (N_9304,N_8996,N_7511);
or U9305 (N_9305,N_6357,N_8820);
xnor U9306 (N_9306,N_7584,N_6843);
and U9307 (N_9307,N_7445,N_7141);
xor U9308 (N_9308,N_8767,N_8055);
xor U9309 (N_9309,N_7846,N_7221);
nand U9310 (N_9310,N_8810,N_8919);
and U9311 (N_9311,N_7582,N_6522);
and U9312 (N_9312,N_8693,N_8492);
and U9313 (N_9313,N_7677,N_7788);
xor U9314 (N_9314,N_8135,N_6387);
and U9315 (N_9315,N_7087,N_8232);
nand U9316 (N_9316,N_7685,N_6182);
or U9317 (N_9317,N_6868,N_6177);
nor U9318 (N_9318,N_8764,N_8098);
and U9319 (N_9319,N_6069,N_8482);
xnor U9320 (N_9320,N_7664,N_7661);
xnor U9321 (N_9321,N_6703,N_8639);
or U9322 (N_9322,N_6977,N_7898);
nor U9323 (N_9323,N_6934,N_6186);
nand U9324 (N_9324,N_7055,N_8664);
or U9325 (N_9325,N_7449,N_8811);
xnor U9326 (N_9326,N_8699,N_8411);
or U9327 (N_9327,N_7844,N_8106);
nor U9328 (N_9328,N_7126,N_8120);
xor U9329 (N_9329,N_6192,N_8306);
nor U9330 (N_9330,N_6730,N_7697);
and U9331 (N_9331,N_6002,N_6424);
nor U9332 (N_9332,N_6630,N_8871);
nor U9333 (N_9333,N_7808,N_6976);
and U9334 (N_9334,N_7419,N_8673);
nor U9335 (N_9335,N_6679,N_8816);
nand U9336 (N_9336,N_6450,N_8172);
or U9337 (N_9337,N_6956,N_8010);
nand U9338 (N_9338,N_6616,N_8438);
nor U9339 (N_9339,N_6860,N_7864);
or U9340 (N_9340,N_6825,N_7920);
xnor U9341 (N_9341,N_6171,N_6526);
nor U9342 (N_9342,N_8385,N_8034);
nand U9343 (N_9343,N_6535,N_7439);
and U9344 (N_9344,N_8648,N_8633);
nand U9345 (N_9345,N_7515,N_8257);
or U9346 (N_9346,N_7786,N_7082);
nand U9347 (N_9347,N_8715,N_7431);
nand U9348 (N_9348,N_8133,N_8927);
or U9349 (N_9349,N_6850,N_6964);
nor U9350 (N_9350,N_8275,N_8199);
nand U9351 (N_9351,N_8046,N_6062);
nand U9352 (N_9352,N_7905,N_7837);
nor U9353 (N_9353,N_6494,N_8845);
or U9354 (N_9354,N_7824,N_8800);
xor U9355 (N_9355,N_6893,N_7436);
nand U9356 (N_9356,N_8917,N_6264);
nand U9357 (N_9357,N_7162,N_8887);
and U9358 (N_9358,N_8197,N_8660);
or U9359 (N_9359,N_7502,N_6240);
and U9360 (N_9360,N_7806,N_6239);
nand U9361 (N_9361,N_8381,N_6460);
or U9362 (N_9362,N_7363,N_6855);
or U9363 (N_9363,N_7736,N_7784);
or U9364 (N_9364,N_7974,N_8517);
xor U9365 (N_9365,N_7599,N_8156);
nor U9366 (N_9366,N_7675,N_7731);
or U9367 (N_9367,N_6492,N_8785);
nand U9368 (N_9368,N_6905,N_6064);
nor U9369 (N_9369,N_7152,N_8819);
nand U9370 (N_9370,N_8677,N_8527);
or U9371 (N_9371,N_8920,N_6311);
or U9372 (N_9372,N_6707,N_7479);
xnor U9373 (N_9373,N_7866,N_7915);
nand U9374 (N_9374,N_8846,N_7933);
xor U9375 (N_9375,N_8579,N_6248);
nand U9376 (N_9376,N_7373,N_6013);
or U9377 (N_9377,N_6668,N_6109);
and U9378 (N_9378,N_7826,N_7516);
and U9379 (N_9379,N_8041,N_8445);
and U9380 (N_9380,N_6458,N_7768);
or U9381 (N_9381,N_6532,N_7610);
xnor U9382 (N_9382,N_7025,N_7807);
xor U9383 (N_9383,N_6131,N_7563);
and U9384 (N_9384,N_7522,N_7358);
or U9385 (N_9385,N_6414,N_7455);
or U9386 (N_9386,N_6175,N_8722);
or U9387 (N_9387,N_6767,N_8702);
and U9388 (N_9388,N_8794,N_6737);
nand U9389 (N_9389,N_6605,N_6732);
nor U9390 (N_9390,N_6549,N_7263);
xor U9391 (N_9391,N_7614,N_7961);
or U9392 (N_9392,N_8479,N_7333);
xor U9393 (N_9393,N_6470,N_7233);
and U9394 (N_9394,N_8580,N_8035);
and U9395 (N_9395,N_7111,N_7145);
xnor U9396 (N_9396,N_6856,N_7701);
xor U9397 (N_9397,N_6108,N_8608);
xor U9398 (N_9398,N_8833,N_7581);
xnor U9399 (N_9399,N_7117,N_8876);
and U9400 (N_9400,N_7166,N_6373);
nand U9401 (N_9401,N_8993,N_6305);
or U9402 (N_9402,N_7415,N_8812);
nor U9403 (N_9403,N_8078,N_6271);
xnor U9404 (N_9404,N_7653,N_7916);
xnor U9405 (N_9405,N_8218,N_7749);
or U9406 (N_9406,N_7723,N_6713);
or U9407 (N_9407,N_7447,N_7216);
or U9408 (N_9408,N_7670,N_7429);
nor U9409 (N_9409,N_8319,N_6895);
nor U9410 (N_9410,N_6099,N_7338);
xnor U9411 (N_9411,N_8921,N_7839);
and U9412 (N_9412,N_7524,N_8065);
nor U9413 (N_9413,N_6690,N_8191);
and U9414 (N_9414,N_7583,N_7061);
and U9415 (N_9415,N_8451,N_8965);
nor U9416 (N_9416,N_6000,N_8680);
and U9417 (N_9417,N_7900,N_6724);
xor U9418 (N_9418,N_6121,N_8054);
nand U9419 (N_9419,N_7712,N_8047);
and U9420 (N_9420,N_8893,N_8862);
xnor U9421 (N_9421,N_6923,N_8718);
nand U9422 (N_9422,N_7792,N_8575);
and U9423 (N_9423,N_7540,N_7829);
xor U9424 (N_9424,N_6781,N_7728);
nand U9425 (N_9425,N_8302,N_8450);
nand U9426 (N_9426,N_6446,N_7781);
xor U9427 (N_9427,N_8141,N_8881);
nor U9428 (N_9428,N_8804,N_8233);
nor U9429 (N_9429,N_8004,N_6116);
nand U9430 (N_9430,N_6488,N_7772);
and U9431 (N_9431,N_7158,N_8345);
and U9432 (N_9432,N_7561,N_7321);
xor U9433 (N_9433,N_6706,N_6416);
nand U9434 (N_9434,N_6583,N_6308);
nand U9435 (N_9435,N_7215,N_7400);
xnor U9436 (N_9436,N_7711,N_6259);
xnor U9437 (N_9437,N_8378,N_7128);
nor U9438 (N_9438,N_7545,N_6663);
or U9439 (N_9439,N_7539,N_8309);
xor U9440 (N_9440,N_6987,N_6151);
and U9441 (N_9441,N_6343,N_7265);
or U9442 (N_9442,N_7395,N_7733);
or U9443 (N_9443,N_6193,N_8926);
nand U9444 (N_9444,N_6261,N_6965);
and U9445 (N_9445,N_6803,N_7188);
nand U9446 (N_9446,N_6071,N_7238);
nand U9447 (N_9447,N_8591,N_6997);
or U9448 (N_9448,N_8220,N_8308);
xnor U9449 (N_9449,N_8547,N_6935);
nor U9450 (N_9450,N_6736,N_8734);
nand U9451 (N_9451,N_7573,N_7965);
xnor U9452 (N_9452,N_7903,N_6865);
and U9453 (N_9453,N_6032,N_8914);
nor U9454 (N_9454,N_7954,N_7996);
and U9455 (N_9455,N_7517,N_8629);
nor U9456 (N_9456,N_8615,N_7822);
or U9457 (N_9457,N_8085,N_8859);
xnor U9458 (N_9458,N_6537,N_8796);
or U9459 (N_9459,N_7153,N_7101);
nor U9460 (N_9460,N_8393,N_6281);
nor U9461 (N_9461,N_8522,N_8707);
and U9462 (N_9462,N_8057,N_7303);
nor U9463 (N_9463,N_8435,N_6578);
and U9464 (N_9464,N_6727,N_6858);
nor U9465 (N_9465,N_8976,N_6493);
and U9466 (N_9466,N_6031,N_6285);
xor U9467 (N_9467,N_6153,N_8644);
nor U9468 (N_9468,N_6862,N_7328);
or U9469 (N_9469,N_8780,N_6917);
nor U9470 (N_9470,N_7332,N_6718);
xnor U9471 (N_9471,N_7173,N_6745);
xnor U9472 (N_9472,N_7144,N_8988);
nor U9473 (N_9473,N_8088,N_8793);
nand U9474 (N_9474,N_8523,N_7345);
nand U9475 (N_9475,N_7713,N_6179);
nand U9476 (N_9476,N_7848,N_7013);
or U9477 (N_9477,N_8414,N_7251);
and U9478 (N_9478,N_7088,N_6871);
or U9479 (N_9479,N_8766,N_6061);
nand U9480 (N_9480,N_6203,N_8814);
or U9481 (N_9481,N_8666,N_6347);
xor U9482 (N_9482,N_7045,N_6279);
and U9483 (N_9483,N_7803,N_7026);
xor U9484 (N_9484,N_7560,N_8956);
nand U9485 (N_9485,N_7501,N_7565);
nand U9486 (N_9486,N_8880,N_8084);
or U9487 (N_9487,N_8755,N_7960);
and U9488 (N_9488,N_6419,N_7064);
and U9489 (N_9489,N_7612,N_6789);
nor U9490 (N_9490,N_6835,N_8278);
or U9491 (N_9491,N_7404,N_7812);
xnor U9492 (N_9492,N_6889,N_8807);
and U9493 (N_9493,N_8890,N_7925);
xor U9494 (N_9494,N_7150,N_7371);
nand U9495 (N_9495,N_6058,N_6478);
nor U9496 (N_9496,N_6757,N_6628);
nand U9497 (N_9497,N_6870,N_7183);
nor U9498 (N_9498,N_8036,N_7849);
nor U9499 (N_9499,N_8848,N_6799);
nor U9500 (N_9500,N_6902,N_7951);
or U9501 (N_9501,N_7377,N_7028);
or U9502 (N_9502,N_8075,N_8024);
or U9503 (N_9503,N_8896,N_6919);
nand U9504 (N_9504,N_7405,N_7810);
or U9505 (N_9505,N_6037,N_7546);
and U9506 (N_9506,N_6839,N_6332);
nand U9507 (N_9507,N_8748,N_6388);
nor U9508 (N_9508,N_6496,N_8315);
nand U9509 (N_9509,N_6086,N_6837);
xor U9510 (N_9510,N_7840,N_6829);
and U9511 (N_9511,N_6512,N_6065);
and U9512 (N_9512,N_7031,N_6480);
or U9513 (N_9513,N_6038,N_8100);
nor U9514 (N_9514,N_6556,N_7256);
and U9515 (N_9515,N_7314,N_6146);
nand U9516 (N_9516,N_6070,N_8947);
nor U9517 (N_9517,N_7094,N_8539);
nor U9518 (N_9518,N_8281,N_8143);
or U9519 (N_9519,N_7399,N_8066);
xnor U9520 (N_9520,N_6909,N_8930);
nor U9521 (N_9521,N_7425,N_8923);
xnor U9522 (N_9522,N_8353,N_8455);
xor U9523 (N_9523,N_7997,N_7021);
and U9524 (N_9524,N_7024,N_7976);
or U9525 (N_9525,N_6697,N_7738);
xnor U9526 (N_9526,N_8025,N_7714);
and U9527 (N_9527,N_6097,N_7440);
xnor U9528 (N_9528,N_6606,N_8245);
xnor U9529 (N_9529,N_8737,N_8242);
nor U9530 (N_9530,N_7036,N_7369);
or U9531 (N_9531,N_8825,N_8652);
nand U9532 (N_9532,N_6314,N_8375);
xor U9533 (N_9533,N_8588,N_7370);
xnor U9534 (N_9534,N_8671,N_8432);
nand U9535 (N_9535,N_6345,N_7845);
nand U9536 (N_9536,N_8231,N_8784);
or U9537 (N_9537,N_8264,N_8553);
and U9538 (N_9538,N_6026,N_8596);
nand U9539 (N_9539,N_7698,N_7037);
nor U9540 (N_9540,N_7527,N_8968);
nand U9541 (N_9541,N_6024,N_7362);
xnor U9542 (N_9542,N_8261,N_7764);
and U9543 (N_9543,N_6497,N_8350);
xnor U9544 (N_9544,N_6047,N_8327);
xor U9545 (N_9545,N_7131,N_7044);
or U9546 (N_9546,N_8774,N_7027);
nor U9547 (N_9547,N_6440,N_8367);
nand U9548 (N_9548,N_8312,N_6351);
or U9549 (N_9549,N_7693,N_6511);
nand U9550 (N_9550,N_7142,N_7402);
nand U9551 (N_9551,N_8735,N_7453);
and U9552 (N_9552,N_7245,N_7790);
and U9553 (N_9553,N_6403,N_8839);
or U9554 (N_9554,N_6082,N_6786);
nand U9555 (N_9555,N_8369,N_8071);
nor U9556 (N_9556,N_6407,N_6427);
or U9557 (N_9557,N_7070,N_6572);
xnor U9558 (N_9558,N_8562,N_7520);
or U9559 (N_9559,N_8912,N_6888);
nand U9560 (N_9560,N_7887,N_6479);
xor U9561 (N_9561,N_6629,N_6645);
xnor U9562 (N_9562,N_8898,N_8225);
and U9563 (N_9563,N_8534,N_6242);
or U9564 (N_9564,N_8310,N_7604);
and U9565 (N_9565,N_8397,N_7177);
and U9566 (N_9566,N_7745,N_8285);
nand U9567 (N_9567,N_7060,N_8983);
or U9568 (N_9568,N_8616,N_8368);
nor U9569 (N_9569,N_7484,N_8502);
xor U9570 (N_9570,N_6059,N_7625);
xnor U9571 (N_9571,N_6790,N_7132);
xnor U9572 (N_9572,N_7658,N_7576);
or U9573 (N_9573,N_8407,N_6542);
nor U9574 (N_9574,N_8147,N_7602);
and U9575 (N_9575,N_6401,N_7204);
and U9576 (N_9576,N_6728,N_7674);
nor U9577 (N_9577,N_8586,N_6609);
nor U9578 (N_9578,N_8488,N_6661);
nor U9579 (N_9579,N_7796,N_7742);
nor U9580 (N_9580,N_7190,N_7196);
and U9581 (N_9581,N_8858,N_8649);
and U9582 (N_9582,N_7949,N_7050);
or U9583 (N_9583,N_6973,N_7368);
nand U9584 (N_9584,N_8726,N_6051);
or U9585 (N_9585,N_6187,N_8691);
nor U9586 (N_9586,N_6251,N_6918);
nand U9587 (N_9587,N_7279,N_8844);
or U9588 (N_9588,N_6863,N_8611);
and U9589 (N_9589,N_8929,N_6165);
or U9590 (N_9590,N_7633,N_6986);
xnor U9591 (N_9591,N_8131,N_8067);
nor U9592 (N_9592,N_6320,N_8270);
nand U9593 (N_9593,N_7414,N_6152);
xnor U9594 (N_9594,N_8874,N_6788);
or U9595 (N_9595,N_8564,N_7310);
nand U9596 (N_9596,N_8110,N_6232);
and U9597 (N_9597,N_7356,N_7010);
nand U9598 (N_9598,N_8384,N_7063);
or U9599 (N_9599,N_8234,N_7409);
or U9600 (N_9600,N_8102,N_6374);
nor U9601 (N_9601,N_6590,N_7601);
or U9602 (N_9602,N_8902,N_6227);
nand U9603 (N_9603,N_7239,N_6772);
and U9604 (N_9604,N_7899,N_6360);
and U9605 (N_9605,N_7487,N_6025);
and U9606 (N_9606,N_8295,N_8405);
xnor U9607 (N_9607,N_8083,N_8749);
nor U9608 (N_9608,N_8721,N_7297);
and U9609 (N_9609,N_7472,N_7667);
nor U9610 (N_9610,N_6570,N_8059);
or U9611 (N_9611,N_6619,N_7413);
nor U9612 (N_9612,N_6752,N_6953);
xor U9613 (N_9613,N_6838,N_6602);
nor U9614 (N_9614,N_6010,N_7538);
nor U9615 (N_9615,N_6233,N_7112);
or U9616 (N_9616,N_8173,N_8003);
xnor U9617 (N_9617,N_8545,N_6435);
and U9618 (N_9618,N_7387,N_8552);
nand U9619 (N_9619,N_8736,N_6615);
and U9620 (N_9620,N_6266,N_7747);
or U9621 (N_9621,N_6395,N_6539);
nor U9622 (N_9622,N_6957,N_7433);
nand U9623 (N_9623,N_7114,N_8955);
nand U9624 (N_9624,N_7473,N_6508);
xor U9625 (N_9625,N_7638,N_8822);
xnor U9626 (N_9626,N_7856,N_6523);
nand U9627 (N_9627,N_7226,N_8980);
xor U9628 (N_9628,N_6170,N_7968);
nand U9629 (N_9629,N_7053,N_8948);
nand U9630 (N_9630,N_7354,N_7507);
and U9631 (N_9631,N_7509,N_7592);
xnor U9632 (N_9632,N_6180,N_6992);
nor U9633 (N_9633,N_8484,N_7133);
nor U9634 (N_9634,N_8540,N_6415);
and U9635 (N_9635,N_8195,N_6091);
or U9636 (N_9636,N_6929,N_8398);
nor U9637 (N_9637,N_7969,N_7652);
xnor U9638 (N_9638,N_8728,N_7095);
xnor U9639 (N_9639,N_7683,N_8214);
nand U9640 (N_9640,N_7259,N_7986);
nand U9641 (N_9641,N_6204,N_6655);
nand U9642 (N_9642,N_7326,N_6355);
nor U9643 (N_9643,N_6135,N_6341);
xor U9644 (N_9644,N_6247,N_7729);
nor U9645 (N_9645,N_7486,N_7148);
nand U9646 (N_9646,N_6334,N_6092);
xor U9647 (N_9647,N_7450,N_7572);
nand U9648 (N_9648,N_6048,N_7480);
nor U9649 (N_9649,N_6765,N_8897);
nor U9650 (N_9650,N_7505,N_7870);
xnor U9651 (N_9651,N_6005,N_8402);
or U9652 (N_9652,N_8356,N_7746);
and U9653 (N_9653,N_7835,N_8005);
and U9654 (N_9654,N_6698,N_7774);
nor U9655 (N_9655,N_6270,N_8679);
nor U9656 (N_9656,N_6358,N_7927);
or U9657 (N_9657,N_7942,N_7103);
nand U9658 (N_9658,N_6758,N_7032);
or U9659 (N_9659,N_8061,N_7979);
and U9660 (N_9660,N_7347,N_6044);
nor U9661 (N_9661,N_6574,N_8584);
nor U9662 (N_9662,N_8406,N_7330);
xor U9663 (N_9663,N_8395,N_7353);
xnor U9664 (N_9664,N_8631,N_7514);
xor U9665 (N_9665,N_7673,N_7285);
nand U9666 (N_9666,N_8524,N_7929);
nor U9667 (N_9667,N_8311,N_6505);
and U9668 (N_9668,N_6085,N_6938);
or U9669 (N_9669,N_7780,N_7734);
or U9670 (N_9670,N_7568,N_6362);
nand U9671 (N_9671,N_6317,N_8207);
nand U9672 (N_9672,N_8355,N_6183);
or U9673 (N_9673,N_6529,N_8485);
or U9674 (N_9674,N_8373,N_8473);
nand U9675 (N_9675,N_8548,N_6447);
or U9676 (N_9676,N_8305,N_6983);
xnor U9677 (N_9677,N_6903,N_8997);
nor U9678 (N_9678,N_7770,N_6525);
nor U9679 (N_9679,N_7523,N_8883);
xor U9680 (N_9680,N_7262,N_8154);
or U9681 (N_9681,N_8343,N_8093);
xnor U9682 (N_9682,N_8138,N_7306);
nor U9683 (N_9683,N_7865,N_8408);
nor U9684 (N_9684,N_6067,N_8550);
xnor U9685 (N_9685,N_7308,N_8421);
nand U9686 (N_9686,N_6489,N_7838);
xnor U9687 (N_9687,N_6673,N_8668);
nor U9688 (N_9688,N_7955,N_6313);
nand U9689 (N_9689,N_8249,N_6514);
and U9690 (N_9690,N_8152,N_8977);
or U9691 (N_9691,N_7275,N_8215);
nor U9692 (N_9692,N_7532,N_8932);
nand U9693 (N_9693,N_6252,N_6798);
nor U9694 (N_9694,N_8044,N_7883);
xor U9695 (N_9695,N_7388,N_6205);
nand U9696 (N_9696,N_8150,N_8117);
nand U9697 (N_9697,N_7935,N_7001);
and U9698 (N_9698,N_6201,N_8895);
xor U9699 (N_9699,N_6669,N_6940);
xnor U9700 (N_9700,N_7708,N_6975);
or U9701 (N_9701,N_7871,N_6582);
xnor U9702 (N_9702,N_7946,N_8260);
or U9703 (N_9703,N_8818,N_6181);
nor U9704 (N_9704,N_7163,N_7247);
xnor U9705 (N_9705,N_8425,N_6932);
or U9706 (N_9706,N_7643,N_7575);
nor U9707 (N_9707,N_6502,N_8282);
nor U9708 (N_9708,N_8208,N_7867);
nor U9709 (N_9709,N_7761,N_6140);
or U9710 (N_9710,N_8018,N_6123);
and U9711 (N_9711,N_6434,N_8291);
and U9712 (N_9712,N_8420,N_6555);
or U9713 (N_9713,N_8360,N_6891);
or U9714 (N_9714,N_7104,N_7574);
xnor U9715 (N_9715,N_8247,N_7170);
or U9716 (N_9716,N_8571,N_8316);
xnor U9717 (N_9717,N_8423,N_7282);
nor U9718 (N_9718,N_8951,N_6952);
nand U9719 (N_9719,N_8401,N_7288);
or U9720 (N_9720,N_6223,N_7977);
nor U9721 (N_9721,N_8415,N_7073);
nand U9722 (N_9722,N_6164,N_7789);
xnor U9723 (N_9723,N_7904,N_6595);
nand U9724 (N_9724,N_7490,N_6560);
nand U9725 (N_9725,N_6463,N_6218);
and U9726 (N_9726,N_8763,N_8324);
and U9727 (N_9727,N_8738,N_7317);
or U9728 (N_9728,N_8860,N_7284);
nor U9729 (N_9729,N_8399,N_6519);
nor U9730 (N_9730,N_7737,N_7834);
or U9731 (N_9731,N_6674,N_6158);
nor U9732 (N_9732,N_8374,N_8840);
nand U9733 (N_9733,N_7859,N_7662);
xor U9734 (N_9734,N_6238,N_6491);
or U9735 (N_9735,N_8033,N_6221);
and U9736 (N_9736,N_6142,N_7106);
nor U9737 (N_9737,N_8808,N_8497);
and U9738 (N_9738,N_7526,N_7640);
and U9739 (N_9739,N_6004,N_6300);
or U9740 (N_9740,N_8729,N_6744);
xnor U9741 (N_9741,N_7130,N_7634);
nor U9742 (N_9742,N_7743,N_8122);
nor U9743 (N_9743,N_6036,N_8513);
or U9744 (N_9744,N_8465,N_6925);
nor U9745 (N_9745,N_7531,N_6327);
nor U9746 (N_9746,N_7593,N_6822);
nand U9747 (N_9747,N_6075,N_6716);
or U9748 (N_9748,N_7932,N_8683);
or U9749 (N_9749,N_7454,N_7553);
or U9750 (N_9750,N_7165,N_6814);
nand U9751 (N_9751,N_7644,N_8581);
xnor U9752 (N_9752,N_6603,N_7393);
nor U9753 (N_9753,N_8014,N_8175);
and U9754 (N_9754,N_7460,N_6621);
nand U9755 (N_9755,N_7506,N_7002);
or U9756 (N_9756,N_7570,N_8189);
nor U9757 (N_9757,N_6011,N_8364);
and U9758 (N_9758,N_6110,N_8984);
or U9759 (N_9759,N_8463,N_6132);
and U9760 (N_9760,N_7072,N_6995);
nor U9761 (N_9761,N_8019,N_8298);
nor U9762 (N_9762,N_6801,N_8959);
and U9763 (N_9763,N_8506,N_8427);
and U9764 (N_9764,N_7475,N_8183);
or U9765 (N_9765,N_6573,N_8276);
nand U9766 (N_9766,N_8164,N_6195);
nor U9767 (N_9767,N_6098,N_6558);
xnor U9768 (N_9768,N_6167,N_8258);
nand U9769 (N_9769,N_6680,N_7051);
xnor U9770 (N_9770,N_6750,N_6006);
xnor U9771 (N_9771,N_6637,N_7266);
nand U9772 (N_9772,N_6465,N_7530);
xnor U9773 (N_9773,N_8733,N_6875);
or U9774 (N_9774,N_8363,N_7277);
or U9775 (N_9775,N_6598,N_7086);
xnor U9776 (N_9776,N_8777,N_6979);
xor U9777 (N_9777,N_6235,N_7296);
or U9778 (N_9778,N_7428,N_7645);
or U9779 (N_9779,N_6947,N_7909);
xor U9780 (N_9780,N_6417,N_7497);
xnor U9781 (N_9781,N_6377,N_8030);
xnor U9782 (N_9782,N_6474,N_8789);
nor U9783 (N_9783,N_6461,N_7301);
xnor U9784 (N_9784,N_7124,N_8576);
xnor U9785 (N_9785,N_8127,N_7533);
or U9786 (N_9786,N_6885,N_7208);
xor U9787 (N_9787,N_7319,N_8304);
nand U9788 (N_9788,N_7182,N_6297);
and U9789 (N_9789,N_7985,N_8770);
nand U9790 (N_9790,N_7006,N_8076);
xor U9791 (N_9791,N_8873,N_7318);
or U9792 (N_9792,N_8213,N_8941);
nand U9793 (N_9793,N_7207,N_8203);
and U9794 (N_9794,N_7139,N_7287);
or U9795 (N_9795,N_6276,N_8978);
nand U9796 (N_9796,N_7571,N_8194);
nand U9797 (N_9797,N_8192,N_7123);
xor U9798 (N_9798,N_7852,N_6229);
xnor U9799 (N_9799,N_8483,N_8595);
xnor U9800 (N_9800,N_7665,N_6970);
and U9801 (N_9801,N_8157,N_7482);
and U9802 (N_9802,N_6301,N_6466);
nand U9803 (N_9803,N_6390,N_7894);
and U9804 (N_9804,N_8957,N_7882);
nor U9805 (N_9805,N_6699,N_6258);
and U9806 (N_9806,N_8678,N_6352);
and U9807 (N_9807,N_8841,N_8389);
nand U9808 (N_9808,N_6600,N_8669);
and U9809 (N_9809,N_6644,N_7901);
or U9810 (N_9810,N_8032,N_8942);
or U9811 (N_9811,N_7205,N_7348);
nand U9812 (N_9812,N_8006,N_6949);
or U9813 (N_9813,N_8501,N_8458);
nand U9814 (N_9814,N_8239,N_8602);
and U9815 (N_9815,N_6169,N_6920);
xor U9816 (N_9816,N_6774,N_7642);
or U9817 (N_9817,N_7209,N_8297);
nor U9818 (N_9818,N_8325,N_8982);
or U9819 (N_9819,N_6601,N_8322);
nor U9820 (N_9820,N_6087,N_6393);
and U9821 (N_9821,N_6339,N_6326);
nand U9822 (N_9822,N_8145,N_6021);
nand U9823 (N_9823,N_6441,N_8799);
or U9824 (N_9824,N_7669,N_6579);
xor U9825 (N_9825,N_8842,N_8111);
nor U9826 (N_9826,N_8592,N_8806);
and U9827 (N_9827,N_8675,N_6659);
or U9828 (N_9828,N_8365,N_7438);
nand U9829 (N_9829,N_7289,N_7519);
xor U9830 (N_9830,N_8531,N_6817);
or U9831 (N_9831,N_6930,N_7760);
nor U9832 (N_9832,N_6524,N_7237);
and U9833 (N_9833,N_8039,N_8410);
nand U9834 (N_9834,N_8109,N_6249);
or U9835 (N_9835,N_6007,N_7191);
nor U9836 (N_9836,N_6309,N_6338);
nand U9837 (N_9837,N_8761,N_8511);
xor U9838 (N_9838,N_7380,N_6473);
nor U9839 (N_9839,N_7416,N_8510);
nor U9840 (N_9840,N_6321,N_6323);
xnor U9841 (N_9841,N_7292,N_7992);
nor U9842 (N_9842,N_7841,N_8489);
xnor U9843 (N_9843,N_6999,N_6445);
and U9844 (N_9844,N_8299,N_7430);
and U9845 (N_9845,N_8508,N_7649);
and U9846 (N_9846,N_8447,N_8536);
nor U9847 (N_9847,N_6294,N_8753);
or U9848 (N_9848,N_6023,N_7758);
xor U9849 (N_9849,N_6275,N_6274);
and U9850 (N_9850,N_8773,N_7830);
or U9851 (N_9851,N_7280,N_6484);
xor U9852 (N_9852,N_7016,N_8158);
and U9853 (N_9853,N_6063,N_6734);
nor U9854 (N_9854,N_6554,N_6874);
or U9855 (N_9855,N_8013,N_6936);
or U9856 (N_9856,N_8460,N_7090);
or U9857 (N_9857,N_6378,N_6982);
nor U9858 (N_9858,N_7488,N_6141);
and U9859 (N_9859,N_6501,N_7293);
and U9860 (N_9860,N_8294,N_6700);
and U9861 (N_9861,N_6939,N_6733);
or U9862 (N_9862,N_8255,N_8986);
or U9863 (N_9863,N_6421,N_8357);
nand U9864 (N_9864,N_7071,N_7099);
nand U9865 (N_9865,N_7127,N_7329);
nor U9866 (N_9866,N_7476,N_6764);
xnor U9867 (N_9867,N_8070,N_7206);
nand U9868 (N_9868,N_8529,N_6124);
or U9869 (N_9869,N_6016,N_7783);
nand U9870 (N_9870,N_8663,N_7459);
nand U9871 (N_9871,N_7727,N_8137);
xnor U9872 (N_9872,N_7874,N_6810);
nor U9873 (N_9873,N_6773,N_6985);
nand U9874 (N_9874,N_6293,N_7046);
or U9875 (N_9875,N_7948,N_8095);
nor U9876 (N_9876,N_7550,N_8020);
xor U9877 (N_9877,N_8744,N_8651);
or U9878 (N_9878,N_7286,N_6516);
and U9879 (N_9879,N_8787,N_7418);
nand U9880 (N_9880,N_8028,N_6095);
nor U9881 (N_9881,N_8797,N_7352);
nor U9882 (N_9882,N_6245,N_8618);
and U9883 (N_9883,N_7655,N_8370);
nor U9884 (N_9884,N_6793,N_7557);
xor U9885 (N_9885,N_6625,N_8835);
and U9886 (N_9886,N_6638,N_7564);
nor U9887 (N_9887,N_8803,N_7767);
or U9888 (N_9888,N_8177,N_6216);
or U9889 (N_9889,N_8179,N_6969);
xnor U9890 (N_9890,N_6129,N_6959);
and U9891 (N_9891,N_7587,N_8178);
nor U9892 (N_9892,N_6741,N_6815);
nor U9893 (N_9893,N_6816,N_7108);
nor U9894 (N_9894,N_8783,N_8532);
xnor U9895 (N_9895,N_8439,N_8185);
nor U9896 (N_9896,N_8321,N_8256);
xnor U9897 (N_9897,N_8760,N_7408);
and U9898 (N_9898,N_6755,N_6569);
or U9899 (N_9899,N_7007,N_6217);
nor U9900 (N_9900,N_7022,N_6425);
or U9901 (N_9901,N_6797,N_8491);
xor U9902 (N_9902,N_7548,N_7220);
nand U9903 (N_9903,N_7469,N_7242);
nor U9904 (N_9904,N_7496,N_6557);
nand U9905 (N_9905,N_8528,N_6587);
and U9906 (N_9906,N_6022,N_7791);
and U9907 (N_9907,N_6544,N_7441);
nand U9908 (N_9908,N_8830,N_8665);
or U9909 (N_9909,N_8950,N_6495);
xnor U9910 (N_9910,N_8412,N_6335);
xor U9911 (N_9911,N_8624,N_6704);
or U9912 (N_9912,N_7271,N_8558);
nor U9913 (N_9913,N_6611,N_6849);
and U9914 (N_9914,N_6702,N_8521);
xor U9915 (N_9915,N_8765,N_8943);
and U9916 (N_9916,N_7023,N_7715);
or U9917 (N_9917,N_7912,N_8772);
or U9918 (N_9918,N_6927,N_8868);
or U9919 (N_9919,N_8991,N_7075);
xor U9920 (N_9920,N_8340,N_6102);
xor U9921 (N_9921,N_8444,N_8716);
and U9922 (N_9922,N_7147,N_7717);
nor U9923 (N_9923,N_8457,N_6077);
and U9924 (N_9924,N_7065,N_6943);
xnor U9925 (N_9925,N_6100,N_7800);
nor U9926 (N_9926,N_8972,N_8636);
and U9927 (N_9927,N_8940,N_7978);
nand U9928 (N_9928,N_6543,N_8720);
nor U9929 (N_9929,N_6960,N_6476);
and U9930 (N_9930,N_7386,N_7134);
xnor U9931 (N_9931,N_6576,N_7939);
nor U9932 (N_9932,N_7991,N_7435);
nor U9933 (N_9933,N_7884,N_8128);
nand U9934 (N_9934,N_7485,N_8834);
nand U9935 (N_9935,N_8640,N_8676);
nor U9936 (N_9936,N_7831,N_8062);
and U9937 (N_9937,N_6246,N_8614);
nand U9938 (N_9938,N_6802,N_7577);
nand U9939 (N_9939,N_7650,N_8366);
and U9940 (N_9940,N_8904,N_8252);
xnor U9941 (N_9941,N_8193,N_7421);
nor U9942 (N_9942,N_8538,N_6751);
nor U9943 (N_9943,N_6076,N_6785);
or U9944 (N_9944,N_7589,N_8092);
nor U9945 (N_9945,N_7281,N_6531);
xnor U9946 (N_9946,N_8525,N_6651);
xor U9947 (N_9947,N_7092,N_6211);
or U9948 (N_9948,N_6443,N_8867);
nand U9949 (N_9949,N_8599,N_7043);
nor U9950 (N_9950,N_6284,N_6540);
xnor U9951 (N_9951,N_7821,N_8090);
or U9952 (N_9952,N_7218,N_6517);
nor U9953 (N_9953,N_6833,N_7236);
or U9954 (N_9954,N_6711,N_7608);
nand U9955 (N_9955,N_6214,N_6719);
and U9956 (N_9956,N_8658,N_6794);
or U9957 (N_9957,N_6383,N_6113);
and U9958 (N_9958,N_7192,N_8112);
nor U9959 (N_9959,N_6869,N_7962);
xnor U9960 (N_9960,N_6340,N_7253);
xnor U9961 (N_9961,N_8740,N_6255);
and U9962 (N_9962,N_8530,N_7691);
xnor U9963 (N_9963,N_8852,N_7627);
nor U9964 (N_9964,N_6090,N_6212);
or U9965 (N_9965,N_8642,N_8474);
and U9966 (N_9966,N_7254,N_7272);
nor U9967 (N_9967,N_7668,N_8817);
xnor U9968 (N_9968,N_7928,N_7397);
xnor U9969 (N_9969,N_8888,N_7537);
nor U9970 (N_9970,N_7042,N_8542);
xnor U9971 (N_9971,N_6423,N_6804);
nor U9972 (N_9972,N_6043,N_8205);
nor U9973 (N_9973,N_6832,N_8732);
and U9974 (N_9974,N_8843,N_8079);
or U9975 (N_9975,N_6807,N_8509);
nor U9976 (N_9976,N_6429,N_7873);
nor U9977 (N_9977,N_7659,N_8568);
or U9978 (N_9978,N_6139,N_7637);
and U9979 (N_9979,N_6018,N_8011);
nand U9980 (N_9980,N_8709,N_8725);
nand U9981 (N_9981,N_6675,N_8967);
or U9982 (N_9982,N_8475,N_6504);
or U9983 (N_9983,N_8296,N_6876);
and U9984 (N_9984,N_6748,N_8971);
nand U9985 (N_9985,N_7223,N_7500);
or U9986 (N_9986,N_7860,N_6513);
and U9987 (N_9987,N_6391,N_6236);
or U9988 (N_9988,N_6477,N_8990);
nor U9989 (N_9989,N_8174,N_8243);
xor U9990 (N_9990,N_7980,N_8198);
and U9991 (N_9991,N_6289,N_7851);
xnor U9992 (N_9992,N_7312,N_6599);
nand U9993 (N_9993,N_7709,N_8301);
nand U9994 (N_9994,N_8561,N_6897);
xor U9995 (N_9995,N_7198,N_7383);
and U9996 (N_9996,N_7695,N_8227);
and U9997 (N_9997,N_8719,N_7744);
and U9998 (N_9998,N_7750,N_6620);
or U9999 (N_9999,N_8362,N_7773);
or U10000 (N_10000,N_8637,N_7621);
nand U10001 (N_10001,N_6610,N_6818);
xor U10002 (N_10002,N_7058,N_8118);
nand U10003 (N_10003,N_7110,N_7588);
or U10004 (N_10004,N_6641,N_7357);
and U10005 (N_10005,N_7003,N_7994);
nand U10006 (N_10006,N_6197,N_7663);
xnor U10007 (N_10007,N_7041,N_8788);
xnor U10008 (N_10008,N_7143,N_8114);
or U10009 (N_10009,N_7498,N_8565);
nand U10010 (N_10010,N_6046,N_6581);
xnor U10011 (N_10011,N_6712,N_8689);
nand U10012 (N_10012,N_6472,N_8072);
and U10013 (N_10013,N_7015,N_6402);
nor U10014 (N_10014,N_8341,N_8259);
xnor U10015 (N_10015,N_6972,N_6664);
xnor U10016 (N_10016,N_8724,N_6649);
or U10017 (N_10017,N_7225,N_6823);
xor U10018 (N_10018,N_7917,N_7739);
nand U10019 (N_10019,N_6743,N_7464);
and U10020 (N_10020,N_7930,N_6913);
or U10021 (N_10021,N_6545,N_8007);
nand U10022 (N_10022,N_8049,N_8000);
nor U10023 (N_10023,N_6225,N_8656);
nand U10024 (N_10024,N_6020,N_7547);
or U10025 (N_10025,N_8605,N_7434);
and U10026 (N_10026,N_8741,N_6379);
nor U10027 (N_10027,N_8603,N_6296);
xnor U10028 (N_10028,N_6584,N_6080);
or U10029 (N_10029,N_6125,N_7931);
nor U10030 (N_10030,N_6550,N_6019);
nand U10031 (N_10031,N_7077,N_8125);
or U10032 (N_10032,N_8884,N_8149);
and U10033 (N_10033,N_8549,N_8945);
and U10034 (N_10034,N_7756,N_8442);
nor U10035 (N_10035,N_8655,N_8016);
nand U10036 (N_10036,N_6324,N_6694);
nand U10037 (N_10037,N_8210,N_8739);
or U10038 (N_10038,N_6336,N_6892);
or U10039 (N_10039,N_7982,N_8612);
nor U10040 (N_10040,N_7937,N_7448);
nor U10041 (N_10041,N_6665,N_6392);
or U10042 (N_10042,N_8228,N_7213);
and U10043 (N_10043,N_6190,N_6667);
nand U10044 (N_10044,N_6993,N_7973);
xnor U10045 (N_10045,N_6371,N_6653);
and U10046 (N_10046,N_7462,N_6329);
and U10047 (N_10047,N_7085,N_7816);
xor U10048 (N_10048,N_7474,N_8250);
xor U10049 (N_10049,N_8023,N_7730);
nand U10050 (N_10050,N_8520,N_7011);
nand U10051 (N_10051,N_6852,N_8371);
nor U10052 (N_10052,N_6202,N_6872);
nand U10053 (N_10053,N_7417,N_6811);
xnor U10054 (N_10054,N_7181,N_6074);
xnor U10055 (N_10055,N_8165,N_7959);
nand U10056 (N_10056,N_8335,N_8086);
nor U10057 (N_10057,N_8838,N_6754);
and U10058 (N_10058,N_8091,N_7091);
nor U10059 (N_10059,N_7382,N_7069);
and U10060 (N_10060,N_6104,N_6689);
nor U10061 (N_10061,N_7047,N_7679);
nor U10062 (N_10062,N_6319,N_7035);
or U10063 (N_10063,N_7376,N_8776);
xor U10064 (N_10064,N_7171,N_6163);
xor U10065 (N_10065,N_7159,N_8472);
and U10066 (N_10066,N_6451,N_7622);
nand U10067 (N_10067,N_7696,N_8892);
xnor U10068 (N_10068,N_8404,N_6792);
and U10069 (N_10069,N_7222,N_7451);
or U10070 (N_10070,N_6994,N_8604);
nor U10071 (N_10071,N_8646,N_6981);
xor U10072 (N_10072,N_7579,N_6265);
or U10073 (N_10073,N_8939,N_8559);
nand U10074 (N_10074,N_8674,N_7499);
nor U10075 (N_10075,N_7676,N_8960);
and U10076 (N_10076,N_6035,N_6780);
nand U10077 (N_10077,N_8123,N_8756);
or U10078 (N_10078,N_7364,N_8745);
and U10079 (N_10079,N_8621,N_6906);
nor U10080 (N_10080,N_7682,N_6398);
nor U10081 (N_10081,N_8687,N_7057);
or U10082 (N_10082,N_8690,N_6683);
nor U10083 (N_10083,N_8824,N_6559);
nand U10084 (N_10084,N_8323,N_7631);
and U10085 (N_10085,N_8911,N_6596);
or U10086 (N_10086,N_8832,N_7617);
and U10087 (N_10087,N_8418,N_6406);
nand U10088 (N_10088,N_6840,N_8710);
xnor U10089 (N_10089,N_6405,N_7687);
nor U10090 (N_10090,N_6515,N_8879);
nand U10091 (N_10091,N_6509,N_6050);
nor U10092 (N_10092,N_8708,N_6118);
xnor U10093 (N_10093,N_7457,N_8578);
and U10094 (N_10094,N_8692,N_6122);
nor U10095 (N_10095,N_6198,N_8964);
xnor U10096 (N_10096,N_6346,N_6547);
nor U10097 (N_10097,N_6890,N_6878);
or U10098 (N_10098,N_7836,N_6433);
xor U10099 (N_10099,N_6771,N_6857);
and U10100 (N_10100,N_7083,N_8672);
nor U10101 (N_10101,N_6842,N_6455);
nand U10102 (N_10102,N_8352,N_6219);
xnor U10103 (N_10103,N_6224,N_8107);
and U10104 (N_10104,N_7752,N_8670);
xor U10105 (N_10105,N_6372,N_7878);
or U10106 (N_10106,N_8338,N_8382);
nor U10107 (N_10107,N_7510,N_8515);
xor U10108 (N_10108,N_6040,N_7940);
nand U10109 (N_10109,N_6337,N_6438);
xnor U10110 (N_10110,N_6563,N_6851);
and U10111 (N_10111,N_6093,N_7660);
or U10112 (N_10112,N_7359,N_7406);
xnor U10113 (N_10113,N_7858,N_6188);
nand U10114 (N_10114,N_7004,N_8634);
xnor U10115 (N_10115,N_6847,N_8847);
nand U10116 (N_10116,N_6083,N_7797);
and U10117 (N_10117,N_6746,N_6370);
and U10118 (N_10118,N_6027,N_8854);
nand U10119 (N_10119,N_6200,N_7341);
nand U10120 (N_10120,N_7549,N_7097);
nor U10121 (N_10121,N_6408,N_7040);
nand U10122 (N_10122,N_8351,N_7193);
xor U10123 (N_10123,N_8589,N_7876);
and U10124 (N_10124,N_7628,N_8130);
nand U10125 (N_10125,N_8778,N_8853);
or U10126 (N_10126,N_8907,N_8518);
or U10127 (N_10127,N_6974,N_8850);
or U10128 (N_10128,N_6633,N_8855);
and U10129 (N_10129,N_7503,N_7518);
xnor U10130 (N_10130,N_6639,N_7722);
or U10131 (N_10131,N_8533,N_8466);
and U10132 (N_10132,N_7763,N_6978);
nand U10133 (N_10133,N_8029,N_7990);
nand U10134 (N_10134,N_7033,N_8864);
nand U10135 (N_10135,N_8101,N_6546);
and U10136 (N_10136,N_8240,N_7793);
or U10137 (N_10137,N_7135,N_8916);
nand U10138 (N_10138,N_6208,N_7513);
nand U10139 (N_10139,N_6769,N_8103);
xor U10140 (N_10140,N_6693,N_7398);
nand U10141 (N_10141,N_8313,N_8962);
or U10142 (N_10142,N_8237,N_8989);
nor U10143 (N_10143,N_8714,N_7809);
and U10144 (N_10144,N_8909,N_8667);
xor U10145 (N_10145,N_7947,N_8966);
nand U10146 (N_10146,N_8437,N_8863);
and U10147 (N_10147,N_6873,N_8394);
nand U10148 (N_10148,N_8206,N_8200);
xor U10149 (N_10149,N_6701,N_7700);
or U10150 (N_10150,N_7782,N_7609);
nor U10151 (N_10151,N_7235,N_7785);
xnor U10152 (N_10152,N_7970,N_6695);
xor U10153 (N_10153,N_8757,N_6418);
or U10154 (N_10154,N_8038,N_7815);
nor U10155 (N_10155,N_8700,N_7315);
xnor U10156 (N_10156,N_7877,N_6088);
nor U10157 (N_10157,N_7465,N_6299);
xor U10158 (N_10158,N_7320,N_8148);
or U10159 (N_10159,N_8574,N_6753);
and U10160 (N_10160,N_6127,N_6824);
and U10161 (N_10161,N_8638,N_7211);
xor U10162 (N_10162,N_8146,N_7647);
and U10163 (N_10163,N_6739,N_6821);
or U10164 (N_10164,N_7855,N_7125);
xnor U10165 (N_10165,N_6436,N_6030);
and U10166 (N_10166,N_7918,N_8661);
xor U10167 (N_10167,N_7269,N_6805);
and U10168 (N_10168,N_7896,N_8537);
or U10169 (N_10169,N_8769,N_7636);
and U10170 (N_10170,N_7391,N_6658);
and U10171 (N_10171,N_7299,N_7875);
nor U10172 (N_10172,N_6367,N_8347);
nor U10173 (N_10173,N_7267,N_6306);
or U10174 (N_10174,N_8598,N_6107);
and U10175 (N_10175,N_6483,N_7331);
xnor U10176 (N_10176,N_6961,N_6740);
nor U10177 (N_10177,N_8961,N_7847);
xor U10178 (N_10178,N_7424,N_8196);
and U10179 (N_10179,N_7278,N_8476);
nor U10180 (N_10180,N_8396,N_7827);
nor U10181 (N_10181,N_8400,N_8212);
xnor U10182 (N_10182,N_8998,N_8449);
nand U10183 (N_10183,N_6145,N_6189);
xnor U10184 (N_10184,N_8944,N_6409);
and U10185 (N_10185,N_7246,N_7008);
or U10186 (N_10186,N_8925,N_8551);
nor U10187 (N_10187,N_6464,N_6726);
or U10188 (N_10188,N_8226,N_8380);
nand U10189 (N_10189,N_8099,N_6585);
and U10190 (N_10190,N_8184,N_7817);
and U10191 (N_10191,N_6882,N_7943);
and U10192 (N_10192,N_8115,N_8326);
nand U10193 (N_10193,N_8836,N_6866);
and U10194 (N_10194,N_6914,N_8009);
xnor U10195 (N_10195,N_7541,N_8280);
xnor U10196 (N_10196,N_6143,N_6162);
and U10197 (N_10197,N_7274,N_8597);
xnor U10198 (N_10198,N_8503,N_8080);
and U10199 (N_10199,N_8650,N_6292);
xnor U10200 (N_10200,N_6715,N_8975);
nand U10201 (N_10201,N_6826,N_7759);
and U10202 (N_10202,N_7521,N_6520);
or U10203 (N_10203,N_7987,N_7850);
nor U10204 (N_10204,N_6288,N_7598);
and U10205 (N_10205,N_6057,N_8815);
and U10206 (N_10206,N_6778,N_8872);
xor U10207 (N_10207,N_7556,N_6795);
or U10208 (N_10208,N_8630,N_7481);
nor U10209 (N_10209,N_7100,N_8314);
or U10210 (N_10210,N_8985,N_6830);
nand U10211 (N_10211,N_6034,N_6966);
nand U10212 (N_10212,N_7958,N_8217);
and U10213 (N_10213,N_8344,N_7054);
nand U10214 (N_10214,N_6738,N_6302);
or U10215 (N_10215,N_6148,N_8471);
or U10216 (N_10216,N_7200,N_6963);
nor U10217 (N_10217,N_7304,N_7443);
nor U10218 (N_10218,N_7525,N_8329);
nand U10219 (N_10219,N_8202,N_6955);
or U10220 (N_10220,N_7888,N_6886);
nand U10221 (N_10221,N_7403,N_7833);
or U10222 (N_10222,N_8963,N_8448);
or U10223 (N_10223,N_7984,N_7921);
and U10224 (N_10224,N_7508,N_6210);
xor U10225 (N_10225,N_7623,N_6207);
and U10226 (N_10226,N_8320,N_7365);
and U10227 (N_10227,N_7964,N_7995);
nor U10228 (N_10228,N_6017,N_8331);
nand U10229 (N_10229,N_7692,N_6154);
xor U10230 (N_10230,N_7316,N_8495);
xor U10231 (N_10231,N_6836,N_6475);
or U10232 (N_10232,N_8905,N_6577);
nor U10233 (N_10233,N_7492,N_6222);
nand U10234 (N_10234,N_6348,N_7427);
xor U10235 (N_10235,N_8283,N_8544);
nand U10236 (N_10236,N_6688,N_8570);
nor U10237 (N_10237,N_8134,N_7360);
xor U10238 (N_10238,N_8336,N_6333);
nand U10239 (N_10239,N_7228,N_7586);
xnor U10240 (N_10240,N_8505,N_7607);
and U10241 (N_10241,N_7264,N_7543);
nor U10242 (N_10242,N_8031,N_6015);
xnor U10243 (N_10243,N_6101,N_8742);
or U10244 (N_10244,N_6747,N_6469);
nor U10245 (N_10245,N_8682,N_6725);
or U10246 (N_10246,N_7189,N_7922);
nand U10247 (N_10247,N_6672,N_6368);
nor U10248 (N_10248,N_6277,N_6770);
nor U10249 (N_10249,N_8958,N_7605);
nand U10250 (N_10250,N_8974,N_8271);
and U10251 (N_10251,N_6593,N_7688);
nor U10252 (N_10252,N_6623,N_6119);
nand U10253 (N_10253,N_6967,N_7534);
nand U10254 (N_10254,N_8248,N_6161);
nand U10255 (N_10255,N_8910,N_8857);
or U10256 (N_10256,N_7597,N_7911);
nor U10257 (N_10257,N_7300,N_7906);
xnor U10258 (N_10258,N_8698,N_6652);
nor U10259 (N_10259,N_6813,N_8094);
nor U10260 (N_10260,N_8188,N_7394);
xor U10261 (N_10261,N_7566,N_7672);
xnor U10262 (N_10262,N_8229,N_7725);
xnor U10263 (N_10263,N_8802,N_8470);
or U10264 (N_10264,N_7892,N_8933);
nand U10265 (N_10265,N_6053,N_8623);
xnor U10266 (N_10266,N_8142,N_7080);
xnor U10267 (N_10267,N_6642,N_7197);
nand U10268 (N_10268,N_6899,N_6206);
nand U10269 (N_10269,N_6112,N_7243);
xnor U10270 (N_10270,N_6635,N_8477);
and U10271 (N_10271,N_7378,N_6267);
and U10272 (N_10272,N_7340,N_7724);
xnor U10273 (N_10273,N_8104,N_8601);
xnor U10274 (N_10274,N_8002,N_6951);
xor U10275 (N_10275,N_7494,N_8021);
xnor U10276 (N_10276,N_8292,N_8222);
nand U10277 (N_10277,N_7407,N_8587);
and U10278 (N_10278,N_8954,N_8159);
nor U10279 (N_10279,N_8885,N_6457);
and U10280 (N_10280,N_7396,N_8786);
xnor U10281 (N_10281,N_6777,N_6910);
nor U10282 (N_10282,N_6841,N_6705);
and U10283 (N_10283,N_8089,N_7862);
nor U10284 (N_10284,N_6589,N_8452);
xnor U10285 (N_10285,N_7452,N_8535);
and U10286 (N_10286,N_8870,N_8386);
xor U10287 (N_10287,N_8662,N_6575);
nor U10288 (N_10288,N_6411,N_8069);
xnor U10289 (N_10289,N_6507,N_8236);
nand U10290 (N_10290,N_6389,N_7305);
xnor U10291 (N_10291,N_7529,N_7081);
or U10292 (N_10292,N_7140,N_6381);
and U10293 (N_10293,N_8827,N_6155);
nor U10294 (N_10294,N_6359,N_8837);
nand U10295 (N_10295,N_7957,N_8015);
xor U10296 (N_10296,N_8073,N_7107);
or U10297 (N_10297,N_8560,N_7214);
nand U10298 (N_10298,N_6761,N_8869);
xor U10299 (N_10299,N_7118,N_8048);
xor U10300 (N_10300,N_7945,N_6191);
xnor U10301 (N_10301,N_7178,N_7787);
nand U10302 (N_10302,N_8526,N_6536);
or U10303 (N_10303,N_8201,N_6498);
nand U10304 (N_10304,N_6962,N_6650);
xnor U10305 (N_10305,N_7201,N_7062);
and U10306 (N_10306,N_8077,N_7975);
nor U10307 (N_10307,N_7989,N_6273);
or U10308 (N_10308,N_8730,N_7327);
xnor U10309 (N_10309,N_6586,N_6834);
and U10310 (N_10310,N_6924,N_8635);
nand U10311 (N_10311,N_8711,N_7078);
nand U10312 (N_10312,N_6363,N_7483);
and U10313 (N_10313,N_7066,N_8241);
nor U10314 (N_10314,N_7241,N_6883);
nand U10315 (N_10315,N_6806,N_8952);
nor U10316 (N_10316,N_6613,N_6879);
and U10317 (N_10317,N_7639,N_8706);
xor U10318 (N_10318,N_7324,N_8659);
or U10319 (N_10319,N_6487,N_8899);
xnor U10320 (N_10320,N_6762,N_7252);
xnor U10321 (N_10321,N_7495,N_6735);
xor U10322 (N_10322,N_7392,N_8328);
or U10323 (N_10323,N_8750,N_8392);
and U10324 (N_10324,N_6287,N_7694);
xor U10325 (N_10325,N_7093,N_6459);
xor U10326 (N_10326,N_8119,N_6412);
nand U10327 (N_10327,N_6503,N_6420);
and U10328 (N_10328,N_8969,N_6594);
and U10329 (N_10329,N_8512,N_6263);
and U10330 (N_10330,N_8209,N_7554);
nor U10331 (N_10331,N_6646,N_6768);
and U10332 (N_10332,N_8268,N_8953);
nor U10333 (N_10333,N_6710,N_7056);
xor U10334 (N_10334,N_7493,N_6912);
nand U10335 (N_10335,N_8625,N_6867);
nand U10336 (N_10336,N_7068,N_7869);
or U10337 (N_10337,N_7765,N_8758);
xnor U10338 (N_10338,N_7014,N_7666);
and U10339 (N_10339,N_8221,N_6375);
xnor U10340 (N_10340,N_6921,N_7890);
xor U10341 (N_10341,N_6052,N_7936);
nand U10342 (N_10342,N_7686,N_8390);
nor U10343 (N_10343,N_8723,N_7726);
nand U10344 (N_10344,N_6213,N_8153);
or U10345 (N_10345,N_6369,N_7313);
xnor U10346 (N_10346,N_8882,N_7379);
or U10347 (N_10347,N_6400,N_8813);
and U10348 (N_10348,N_7606,N_7861);
or U10349 (N_10349,N_8768,N_7030);
and U10350 (N_10350,N_6709,N_8391);
or U10351 (N_10351,N_8891,N_8936);
nand U10352 (N_10352,N_7105,N_6901);
and U10353 (N_10353,N_7908,N_7635);
nand U10354 (N_10354,N_7230,N_8342);
and U10355 (N_10355,N_6933,N_7458);
xnor U10356 (N_10356,N_7704,N_8284);
xor U10357 (N_10357,N_8752,N_6904);
nand U10358 (N_10358,N_8480,N_8622);
and U10359 (N_10359,N_8647,N_7203);
or U10360 (N_10360,N_8426,N_7720);
and U10361 (N_10361,N_6618,N_6922);
or U10362 (N_10362,N_8922,N_6527);
xnor U10363 (N_10363,N_7832,N_7648);
xor U10364 (N_10364,N_8543,N_6656);
or U10365 (N_10365,N_6565,N_7651);
xnor U10366 (N_10366,N_8171,N_7580);
or U10367 (N_10367,N_6029,N_7555);
and U10368 (N_10368,N_6500,N_8056);
nand U10369 (N_10369,N_8269,N_7076);
nor U10370 (N_10370,N_7067,N_7690);
or U10371 (N_10371,N_7814,N_7470);
and U10372 (N_10372,N_6439,N_7489);
nor U10373 (N_10373,N_7052,N_7307);
or U10374 (N_10374,N_8981,N_8705);
nor U10375 (N_10375,N_8040,N_8045);
or U10376 (N_10376,N_7626,N_6568);
and U10377 (N_10377,N_7872,N_8889);
xor U10378 (N_10378,N_7168,N_8712);
xor U10379 (N_10379,N_6315,N_7893);
and U10380 (N_10380,N_8105,N_6896);
xnor U10381 (N_10381,N_7276,N_8052);
nor U10382 (N_10382,N_8594,N_8216);
or U10383 (N_10383,N_7590,N_7136);
xnor U10384 (N_10384,N_6660,N_6237);
and U10385 (N_10385,N_7880,N_6564);
and U10386 (N_10386,N_8064,N_8801);
nand U10387 (N_10387,N_6948,N_6608);
xor U10388 (N_10388,N_6231,N_7240);
nor U10389 (N_10389,N_6422,N_7349);
xor U10390 (N_10390,N_6530,N_6134);
nor U10391 (N_10391,N_6937,N_6448);
nand U10392 (N_10392,N_8970,N_6254);
and U10393 (N_10393,N_8496,N_7967);
nand U10394 (N_10394,N_6783,N_7227);
nor U10395 (N_10395,N_7249,N_8681);
and U10396 (N_10396,N_8372,N_8754);
nand U10397 (N_10397,N_7971,N_7478);
xnor U10398 (N_10398,N_6676,N_6827);
or U10399 (N_10399,N_7374,N_6328);
and U10400 (N_10400,N_8290,N_6001);
and U10401 (N_10401,N_7591,N_7295);
nand U10402 (N_10402,N_6295,N_7477);
xnor U10403 (N_10403,N_7801,N_6990);
or U10404 (N_10404,N_6078,N_8600);
and U10405 (N_10405,N_6991,N_6136);
or U10406 (N_10406,N_6449,N_8469);
or U10407 (N_10407,N_8422,N_8238);
nand U10408 (N_10408,N_7048,N_8999);
nor U10409 (N_10409,N_7367,N_8915);
xnor U10410 (N_10410,N_8791,N_7707);
or U10411 (N_10411,N_7179,N_8254);
or U10412 (N_10412,N_6384,N_8230);
xnor U10413 (N_10413,N_8566,N_8246);
and U10414 (N_10414,N_6244,N_8695);
nand U10415 (N_10415,N_6518,N_6591);
or U10416 (N_10416,N_6039,N_8160);
or U10417 (N_10417,N_7811,N_7005);
nand U10418 (N_10418,N_7261,N_7703);
or U10419 (N_10419,N_8087,N_8307);
xnor U10420 (N_10420,N_6310,N_7412);
or U10421 (N_10421,N_6354,N_8823);
xnor U10422 (N_10422,N_6253,N_7684);
xnor U10423 (N_10423,N_7632,N_8348);
nand U10424 (N_10424,N_7794,N_7854);
nand U10425 (N_10425,N_6380,N_7766);
nor U10426 (N_10426,N_7934,N_8383);
or U10427 (N_10427,N_8334,N_8251);
xor U10428 (N_10428,N_8628,N_8632);
and U10429 (N_10429,N_7558,N_7372);
nor U10430 (N_10430,N_6468,N_8931);
nand U10431 (N_10431,N_6168,N_6243);
xnor U10432 (N_10432,N_7102,N_6654);
or U10433 (N_10433,N_7777,N_8779);
xor U10434 (N_10434,N_7998,N_7983);
xnor U10435 (N_10435,N_8743,N_8151);
and U10436 (N_10436,N_8459,N_6382);
and U10437 (N_10437,N_6272,N_8446);
nor U10438 (N_10438,N_6485,N_6303);
nor U10439 (N_10439,N_6571,N_7199);
or U10440 (N_10440,N_7603,N_6671);
xnor U10441 (N_10441,N_7468,N_8557);
or U10442 (N_10442,N_8430,N_8617);
or U10443 (N_10443,N_7172,N_8487);
and U10444 (N_10444,N_6566,N_8901);
xnor U10445 (N_10445,N_7423,N_6260);
or U10446 (N_10446,N_6945,N_8253);
xnor U10447 (N_10447,N_6481,N_6209);
and U10448 (N_10448,N_6831,N_7157);
or U10449 (N_10449,N_7167,N_6742);
and U10450 (N_10450,N_8443,N_7813);
nand U10451 (N_10451,N_6055,N_7389);
nand U10452 (N_10452,N_7202,N_7913);
and U10453 (N_10453,N_6114,N_7595);
xor U10454 (N_10454,N_8333,N_7820);
nand U10455 (N_10455,N_6766,N_8686);
nor U10456 (N_10456,N_6643,N_8318);
nor U10457 (N_10457,N_6954,N_6241);
or U10458 (N_10458,N_7620,N_6471);
and U10459 (N_10459,N_8792,N_8620);
xnor U10460 (N_10460,N_7089,N_8609);
xor U10461 (N_10461,N_7512,N_7776);
or U10462 (N_10462,N_7361,N_7619);
and U10463 (N_10463,N_7184,N_6278);
xor U10464 (N_10464,N_7963,N_8162);
or U10465 (N_10465,N_8946,N_6648);
nor U10466 (N_10466,N_8190,N_8464);
nand U10467 (N_10467,N_7121,N_8795);
nor U10468 (N_10468,N_6452,N_8287);
nor U10469 (N_10469,N_7818,N_7161);
nor U10470 (N_10470,N_6553,N_6103);
and U10471 (N_10471,N_8593,N_6900);
or U10472 (N_10472,N_7762,N_6534);
and U10473 (N_10473,N_8346,N_8204);
and U10474 (N_10474,N_6349,N_7268);
or U10475 (N_10475,N_6911,N_7337);
or U10476 (N_10476,N_6426,N_6072);
nor U10477 (N_10477,N_7079,N_6562);
and U10478 (N_10478,N_7437,N_6604);
nor U10479 (N_10479,N_8613,N_6394);
or U10480 (N_10480,N_6454,N_6820);
nor U10481 (N_10481,N_7244,N_6580);
nor U10482 (N_10482,N_6364,N_8288);
xor U10483 (N_10483,N_6060,N_8419);
nor U10484 (N_10484,N_8388,N_6174);
or U10485 (N_10485,N_6312,N_6115);
or U10486 (N_10486,N_8731,N_8181);
nand U10487 (N_10487,N_8022,N_6084);
nor U10488 (N_10488,N_8866,N_7681);
or U10489 (N_10489,N_7224,N_7953);
and U10490 (N_10490,N_6784,N_8182);
nor U10491 (N_10491,N_8790,N_7149);
xnor U10492 (N_10492,N_8244,N_6138);
or U10493 (N_10493,N_7805,N_8440);
and U10494 (N_10494,N_6008,N_8556);
nand U10495 (N_10495,N_8555,N_8992);
or U10496 (N_10496,N_7914,N_7432);
and U10497 (N_10497,N_8167,N_8994);
and U10498 (N_10498,N_6350,N_6617);
and U10499 (N_10499,N_8289,N_6199);
nor U10500 (N_10500,N_8281,N_8915);
and U10501 (N_10501,N_8785,N_8332);
and U10502 (N_10502,N_7788,N_6541);
nand U10503 (N_10503,N_7916,N_8102);
or U10504 (N_10504,N_6666,N_7225);
nor U10505 (N_10505,N_7819,N_7978);
xnor U10506 (N_10506,N_6849,N_8980);
nor U10507 (N_10507,N_7213,N_6798);
nand U10508 (N_10508,N_7922,N_7633);
xnor U10509 (N_10509,N_7298,N_7442);
and U10510 (N_10510,N_8255,N_8206);
and U10511 (N_10511,N_6977,N_7601);
and U10512 (N_10512,N_6660,N_8842);
nand U10513 (N_10513,N_6660,N_8777);
nand U10514 (N_10514,N_7353,N_8097);
or U10515 (N_10515,N_7362,N_8261);
and U10516 (N_10516,N_6137,N_8356);
nor U10517 (N_10517,N_8299,N_8553);
and U10518 (N_10518,N_7199,N_6325);
or U10519 (N_10519,N_7201,N_8401);
nor U10520 (N_10520,N_8215,N_8595);
and U10521 (N_10521,N_6106,N_6280);
or U10522 (N_10522,N_7266,N_8924);
nand U10523 (N_10523,N_6821,N_8578);
xor U10524 (N_10524,N_6297,N_6015);
xnor U10525 (N_10525,N_7275,N_8584);
xor U10526 (N_10526,N_6586,N_8967);
nand U10527 (N_10527,N_8097,N_6305);
or U10528 (N_10528,N_8785,N_8114);
and U10529 (N_10529,N_6695,N_6404);
or U10530 (N_10530,N_8877,N_6057);
nor U10531 (N_10531,N_8147,N_8778);
xnor U10532 (N_10532,N_8929,N_8998);
nor U10533 (N_10533,N_8361,N_8196);
nand U10534 (N_10534,N_8457,N_7075);
and U10535 (N_10535,N_6489,N_7501);
nand U10536 (N_10536,N_8837,N_7894);
xnor U10537 (N_10537,N_8621,N_6574);
xnor U10538 (N_10538,N_7839,N_6795);
or U10539 (N_10539,N_6634,N_6524);
nand U10540 (N_10540,N_8067,N_7936);
nor U10541 (N_10541,N_6453,N_6284);
xnor U10542 (N_10542,N_6255,N_6358);
or U10543 (N_10543,N_7879,N_6232);
or U10544 (N_10544,N_8061,N_8773);
nor U10545 (N_10545,N_8336,N_8098);
or U10546 (N_10546,N_7462,N_8676);
nand U10547 (N_10547,N_7482,N_8644);
nand U10548 (N_10548,N_7646,N_6495);
xnor U10549 (N_10549,N_8263,N_8798);
xnor U10550 (N_10550,N_6626,N_8310);
nand U10551 (N_10551,N_7811,N_8815);
nand U10552 (N_10552,N_8700,N_7066);
xnor U10553 (N_10553,N_8076,N_8067);
and U10554 (N_10554,N_7500,N_7420);
and U10555 (N_10555,N_7604,N_8450);
or U10556 (N_10556,N_6921,N_6726);
nor U10557 (N_10557,N_7006,N_8046);
and U10558 (N_10558,N_7123,N_6637);
or U10559 (N_10559,N_8488,N_8537);
xor U10560 (N_10560,N_6270,N_8520);
xnor U10561 (N_10561,N_7451,N_7855);
and U10562 (N_10562,N_8126,N_6371);
nand U10563 (N_10563,N_6415,N_6326);
or U10564 (N_10564,N_8582,N_7730);
nand U10565 (N_10565,N_6867,N_8016);
xnor U10566 (N_10566,N_6068,N_8096);
or U10567 (N_10567,N_6366,N_7430);
nand U10568 (N_10568,N_8403,N_6359);
nand U10569 (N_10569,N_8534,N_8761);
and U10570 (N_10570,N_7663,N_8314);
nand U10571 (N_10571,N_8233,N_8421);
or U10572 (N_10572,N_6835,N_6450);
and U10573 (N_10573,N_6891,N_7325);
nor U10574 (N_10574,N_8105,N_6710);
nand U10575 (N_10575,N_7961,N_6485);
nand U10576 (N_10576,N_7656,N_7568);
or U10577 (N_10577,N_7912,N_8324);
xnor U10578 (N_10578,N_7056,N_8189);
nor U10579 (N_10579,N_7002,N_6719);
nor U10580 (N_10580,N_8225,N_6864);
nand U10581 (N_10581,N_7906,N_6468);
nand U10582 (N_10582,N_6477,N_8021);
and U10583 (N_10583,N_7174,N_8343);
nor U10584 (N_10584,N_8836,N_7825);
and U10585 (N_10585,N_8981,N_7291);
xnor U10586 (N_10586,N_7280,N_7715);
or U10587 (N_10587,N_6456,N_8678);
nor U10588 (N_10588,N_7561,N_7668);
xor U10589 (N_10589,N_6434,N_7023);
nor U10590 (N_10590,N_7970,N_6469);
and U10591 (N_10591,N_6595,N_6830);
nand U10592 (N_10592,N_7138,N_7284);
xnor U10593 (N_10593,N_8196,N_8365);
or U10594 (N_10594,N_8154,N_7090);
nor U10595 (N_10595,N_7853,N_7740);
nor U10596 (N_10596,N_6535,N_6671);
nand U10597 (N_10597,N_8516,N_6414);
nand U10598 (N_10598,N_8346,N_7074);
nor U10599 (N_10599,N_7250,N_7899);
nand U10600 (N_10600,N_6600,N_6798);
nor U10601 (N_10601,N_8463,N_7806);
and U10602 (N_10602,N_8902,N_6913);
xor U10603 (N_10603,N_7960,N_6792);
and U10604 (N_10604,N_6540,N_6646);
nand U10605 (N_10605,N_7811,N_8089);
nand U10606 (N_10606,N_8097,N_8323);
nor U10607 (N_10607,N_7694,N_8689);
nand U10608 (N_10608,N_8623,N_6461);
xor U10609 (N_10609,N_6855,N_7409);
nor U10610 (N_10610,N_7645,N_7093);
or U10611 (N_10611,N_7983,N_6102);
and U10612 (N_10612,N_7381,N_8390);
nor U10613 (N_10613,N_6173,N_7947);
nand U10614 (N_10614,N_7881,N_7854);
nor U10615 (N_10615,N_8566,N_6931);
or U10616 (N_10616,N_6127,N_8717);
or U10617 (N_10617,N_7949,N_7253);
nor U10618 (N_10618,N_6718,N_6033);
and U10619 (N_10619,N_7253,N_7457);
nand U10620 (N_10620,N_6933,N_7253);
nand U10621 (N_10621,N_8412,N_7399);
xnor U10622 (N_10622,N_8211,N_6297);
nand U10623 (N_10623,N_8527,N_6700);
xor U10624 (N_10624,N_7365,N_8835);
or U10625 (N_10625,N_7224,N_7973);
and U10626 (N_10626,N_7012,N_6536);
xor U10627 (N_10627,N_6228,N_6969);
or U10628 (N_10628,N_8775,N_8321);
nand U10629 (N_10629,N_7008,N_8206);
and U10630 (N_10630,N_8964,N_8242);
and U10631 (N_10631,N_7504,N_8332);
and U10632 (N_10632,N_6681,N_6984);
xnor U10633 (N_10633,N_8566,N_6164);
or U10634 (N_10634,N_7951,N_7576);
or U10635 (N_10635,N_8798,N_8444);
nand U10636 (N_10636,N_7627,N_8980);
xor U10637 (N_10637,N_6642,N_6572);
or U10638 (N_10638,N_7730,N_7253);
nand U10639 (N_10639,N_6374,N_8821);
and U10640 (N_10640,N_6990,N_6367);
nor U10641 (N_10641,N_7332,N_6555);
or U10642 (N_10642,N_8298,N_8062);
xor U10643 (N_10643,N_6556,N_7480);
xnor U10644 (N_10644,N_8887,N_6806);
xor U10645 (N_10645,N_6692,N_7775);
or U10646 (N_10646,N_8925,N_8461);
xor U10647 (N_10647,N_7462,N_6149);
nor U10648 (N_10648,N_8373,N_7284);
and U10649 (N_10649,N_8922,N_7865);
nand U10650 (N_10650,N_6343,N_7006);
and U10651 (N_10651,N_8563,N_6155);
xnor U10652 (N_10652,N_7204,N_6337);
nand U10653 (N_10653,N_7982,N_6753);
nor U10654 (N_10654,N_8686,N_8961);
or U10655 (N_10655,N_6138,N_6599);
or U10656 (N_10656,N_6850,N_8277);
xor U10657 (N_10657,N_6409,N_7694);
and U10658 (N_10658,N_7582,N_7531);
or U10659 (N_10659,N_6260,N_6622);
nand U10660 (N_10660,N_6133,N_7071);
or U10661 (N_10661,N_6438,N_7479);
nor U10662 (N_10662,N_6718,N_6369);
nor U10663 (N_10663,N_6829,N_6548);
or U10664 (N_10664,N_8465,N_7938);
xnor U10665 (N_10665,N_8414,N_7719);
or U10666 (N_10666,N_8980,N_8858);
or U10667 (N_10667,N_6011,N_7547);
or U10668 (N_10668,N_6285,N_7542);
or U10669 (N_10669,N_6207,N_7032);
or U10670 (N_10670,N_8169,N_8081);
and U10671 (N_10671,N_6924,N_7496);
nand U10672 (N_10672,N_7126,N_6993);
nand U10673 (N_10673,N_6521,N_8773);
nand U10674 (N_10674,N_7247,N_7207);
xor U10675 (N_10675,N_7761,N_6293);
or U10676 (N_10676,N_7970,N_8511);
or U10677 (N_10677,N_6525,N_7737);
or U10678 (N_10678,N_6913,N_7470);
xor U10679 (N_10679,N_6554,N_8230);
xnor U10680 (N_10680,N_8853,N_6437);
nor U10681 (N_10681,N_8281,N_8380);
nor U10682 (N_10682,N_8277,N_8126);
nand U10683 (N_10683,N_8036,N_7099);
xnor U10684 (N_10684,N_7517,N_7890);
nor U10685 (N_10685,N_7639,N_6360);
xor U10686 (N_10686,N_6226,N_8202);
xnor U10687 (N_10687,N_6623,N_7223);
or U10688 (N_10688,N_6684,N_8017);
xor U10689 (N_10689,N_7553,N_6110);
nor U10690 (N_10690,N_7965,N_6693);
or U10691 (N_10691,N_6492,N_7231);
nor U10692 (N_10692,N_7665,N_8072);
nand U10693 (N_10693,N_7392,N_8330);
and U10694 (N_10694,N_7220,N_8586);
or U10695 (N_10695,N_6187,N_6786);
nand U10696 (N_10696,N_7785,N_7810);
and U10697 (N_10697,N_8878,N_8046);
or U10698 (N_10698,N_8387,N_6185);
or U10699 (N_10699,N_7097,N_6875);
nand U10700 (N_10700,N_6130,N_7718);
nand U10701 (N_10701,N_7507,N_7086);
xnor U10702 (N_10702,N_6333,N_7687);
nand U10703 (N_10703,N_7041,N_6296);
xnor U10704 (N_10704,N_7385,N_8722);
and U10705 (N_10705,N_6202,N_7251);
nor U10706 (N_10706,N_7614,N_8456);
and U10707 (N_10707,N_8377,N_7608);
xor U10708 (N_10708,N_6937,N_6358);
xnor U10709 (N_10709,N_7555,N_8947);
nor U10710 (N_10710,N_7258,N_6198);
nand U10711 (N_10711,N_6570,N_8277);
nand U10712 (N_10712,N_7224,N_7037);
or U10713 (N_10713,N_8624,N_6558);
nand U10714 (N_10714,N_7456,N_7199);
xnor U10715 (N_10715,N_8323,N_8301);
xnor U10716 (N_10716,N_7458,N_7659);
nor U10717 (N_10717,N_7639,N_8338);
nor U10718 (N_10718,N_8783,N_8804);
nand U10719 (N_10719,N_8812,N_7335);
or U10720 (N_10720,N_6409,N_6719);
nand U10721 (N_10721,N_7301,N_7570);
xor U10722 (N_10722,N_8000,N_7195);
nor U10723 (N_10723,N_8070,N_8853);
nand U10724 (N_10724,N_8099,N_7159);
and U10725 (N_10725,N_7656,N_7147);
nor U10726 (N_10726,N_7944,N_6864);
nand U10727 (N_10727,N_6728,N_6156);
nor U10728 (N_10728,N_6663,N_7485);
nand U10729 (N_10729,N_7225,N_7255);
xnor U10730 (N_10730,N_6407,N_6955);
nor U10731 (N_10731,N_8698,N_8997);
and U10732 (N_10732,N_8377,N_7706);
and U10733 (N_10733,N_6165,N_6157);
xor U10734 (N_10734,N_7427,N_8507);
nand U10735 (N_10735,N_6594,N_6115);
or U10736 (N_10736,N_7016,N_8261);
and U10737 (N_10737,N_8886,N_8336);
nor U10738 (N_10738,N_8853,N_8761);
nor U10739 (N_10739,N_6656,N_6235);
xor U10740 (N_10740,N_6283,N_8574);
or U10741 (N_10741,N_6189,N_8776);
and U10742 (N_10742,N_6844,N_8840);
xor U10743 (N_10743,N_7008,N_6783);
xor U10744 (N_10744,N_6940,N_7223);
or U10745 (N_10745,N_7537,N_8686);
xnor U10746 (N_10746,N_8979,N_8382);
xnor U10747 (N_10747,N_6640,N_7495);
or U10748 (N_10748,N_6808,N_7213);
and U10749 (N_10749,N_8511,N_8914);
or U10750 (N_10750,N_6382,N_8256);
xor U10751 (N_10751,N_6364,N_7037);
or U10752 (N_10752,N_8863,N_7364);
nand U10753 (N_10753,N_8140,N_7764);
nand U10754 (N_10754,N_6995,N_7040);
nor U10755 (N_10755,N_8734,N_8563);
or U10756 (N_10756,N_6629,N_7377);
or U10757 (N_10757,N_7264,N_8811);
or U10758 (N_10758,N_6466,N_6154);
and U10759 (N_10759,N_7998,N_8603);
or U10760 (N_10760,N_8423,N_6147);
nor U10761 (N_10761,N_7285,N_7439);
and U10762 (N_10762,N_7363,N_8668);
nor U10763 (N_10763,N_8117,N_6906);
xnor U10764 (N_10764,N_8384,N_6457);
nand U10765 (N_10765,N_7872,N_7319);
or U10766 (N_10766,N_7089,N_6791);
nand U10767 (N_10767,N_7368,N_7583);
nand U10768 (N_10768,N_6372,N_6053);
or U10769 (N_10769,N_6992,N_8337);
xnor U10770 (N_10770,N_8417,N_6485);
xnor U10771 (N_10771,N_6380,N_8244);
nor U10772 (N_10772,N_8679,N_8880);
and U10773 (N_10773,N_6499,N_8402);
nand U10774 (N_10774,N_6093,N_8140);
nand U10775 (N_10775,N_6834,N_6220);
nand U10776 (N_10776,N_8505,N_7455);
or U10777 (N_10777,N_8985,N_8687);
nand U10778 (N_10778,N_8118,N_6886);
or U10779 (N_10779,N_6975,N_6007);
or U10780 (N_10780,N_8823,N_7587);
and U10781 (N_10781,N_7705,N_7771);
nor U10782 (N_10782,N_8958,N_7470);
and U10783 (N_10783,N_6858,N_7426);
or U10784 (N_10784,N_8580,N_6031);
xor U10785 (N_10785,N_6010,N_8608);
nor U10786 (N_10786,N_8375,N_6270);
nor U10787 (N_10787,N_6923,N_7158);
nor U10788 (N_10788,N_8958,N_7502);
xnor U10789 (N_10789,N_6250,N_7419);
nor U10790 (N_10790,N_7807,N_6385);
nand U10791 (N_10791,N_7584,N_6890);
and U10792 (N_10792,N_7073,N_6353);
or U10793 (N_10793,N_8811,N_8506);
nand U10794 (N_10794,N_8377,N_8868);
and U10795 (N_10795,N_8072,N_7647);
and U10796 (N_10796,N_8768,N_7941);
or U10797 (N_10797,N_6471,N_6225);
or U10798 (N_10798,N_7186,N_8558);
and U10799 (N_10799,N_6420,N_8235);
nor U10800 (N_10800,N_6714,N_6547);
and U10801 (N_10801,N_8091,N_6663);
nor U10802 (N_10802,N_8483,N_8838);
and U10803 (N_10803,N_8653,N_7515);
or U10804 (N_10804,N_8960,N_7781);
nand U10805 (N_10805,N_8307,N_6346);
nor U10806 (N_10806,N_8253,N_7706);
nor U10807 (N_10807,N_8618,N_8437);
or U10808 (N_10808,N_6164,N_8874);
nand U10809 (N_10809,N_6414,N_6279);
nor U10810 (N_10810,N_7840,N_8217);
nor U10811 (N_10811,N_7923,N_6846);
xor U10812 (N_10812,N_8811,N_6993);
or U10813 (N_10813,N_8863,N_6689);
nor U10814 (N_10814,N_6494,N_8245);
and U10815 (N_10815,N_8208,N_6781);
nor U10816 (N_10816,N_7304,N_6092);
nor U10817 (N_10817,N_7032,N_6175);
and U10818 (N_10818,N_7020,N_6988);
nand U10819 (N_10819,N_7375,N_8810);
or U10820 (N_10820,N_8804,N_8901);
and U10821 (N_10821,N_6261,N_8868);
nand U10822 (N_10822,N_6639,N_7847);
nor U10823 (N_10823,N_7709,N_7600);
xnor U10824 (N_10824,N_7694,N_7008);
nand U10825 (N_10825,N_7498,N_8327);
or U10826 (N_10826,N_7892,N_6100);
nand U10827 (N_10827,N_6210,N_7130);
or U10828 (N_10828,N_8709,N_6078);
xor U10829 (N_10829,N_6993,N_8312);
nor U10830 (N_10830,N_8034,N_6965);
or U10831 (N_10831,N_6968,N_8378);
or U10832 (N_10832,N_6409,N_8504);
and U10833 (N_10833,N_8598,N_8094);
or U10834 (N_10834,N_7560,N_7819);
nand U10835 (N_10835,N_7795,N_8644);
xnor U10836 (N_10836,N_7385,N_8436);
nor U10837 (N_10837,N_7698,N_7868);
nor U10838 (N_10838,N_7329,N_8951);
and U10839 (N_10839,N_6772,N_6968);
and U10840 (N_10840,N_6343,N_8473);
and U10841 (N_10841,N_6884,N_8794);
nand U10842 (N_10842,N_8070,N_6983);
xor U10843 (N_10843,N_6255,N_8564);
xor U10844 (N_10844,N_7985,N_8351);
nand U10845 (N_10845,N_8986,N_7654);
nor U10846 (N_10846,N_6583,N_6125);
and U10847 (N_10847,N_6948,N_6902);
nand U10848 (N_10848,N_6082,N_7320);
nor U10849 (N_10849,N_8221,N_6135);
xnor U10850 (N_10850,N_8797,N_6309);
nor U10851 (N_10851,N_8064,N_8656);
or U10852 (N_10852,N_8274,N_6841);
and U10853 (N_10853,N_8587,N_8269);
xor U10854 (N_10854,N_6858,N_6168);
and U10855 (N_10855,N_6716,N_7091);
and U10856 (N_10856,N_7829,N_8572);
nor U10857 (N_10857,N_6088,N_6379);
nor U10858 (N_10858,N_6586,N_6975);
nor U10859 (N_10859,N_6233,N_6153);
nor U10860 (N_10860,N_7555,N_8884);
and U10861 (N_10861,N_7407,N_8461);
xnor U10862 (N_10862,N_6671,N_8311);
and U10863 (N_10863,N_7531,N_6848);
nor U10864 (N_10864,N_8164,N_7113);
xor U10865 (N_10865,N_6004,N_7901);
xor U10866 (N_10866,N_7743,N_6434);
and U10867 (N_10867,N_7525,N_8475);
and U10868 (N_10868,N_8356,N_8428);
and U10869 (N_10869,N_6454,N_8901);
and U10870 (N_10870,N_8811,N_7275);
or U10871 (N_10871,N_6755,N_7236);
nor U10872 (N_10872,N_8951,N_7543);
or U10873 (N_10873,N_8535,N_6459);
and U10874 (N_10874,N_8833,N_6126);
nor U10875 (N_10875,N_6404,N_6970);
xnor U10876 (N_10876,N_7338,N_6976);
and U10877 (N_10877,N_8923,N_7566);
xnor U10878 (N_10878,N_7074,N_7413);
nand U10879 (N_10879,N_7692,N_6112);
nor U10880 (N_10880,N_7908,N_7135);
nor U10881 (N_10881,N_8952,N_8446);
or U10882 (N_10882,N_7584,N_6106);
nor U10883 (N_10883,N_7105,N_7222);
nand U10884 (N_10884,N_8743,N_8978);
and U10885 (N_10885,N_6623,N_6851);
nor U10886 (N_10886,N_7638,N_6677);
nand U10887 (N_10887,N_8230,N_8111);
or U10888 (N_10888,N_8107,N_7812);
nand U10889 (N_10889,N_8054,N_6552);
nor U10890 (N_10890,N_6206,N_7693);
nand U10891 (N_10891,N_7339,N_7562);
nor U10892 (N_10892,N_8898,N_7653);
nor U10893 (N_10893,N_6436,N_6867);
xor U10894 (N_10894,N_8285,N_8516);
and U10895 (N_10895,N_6416,N_6802);
and U10896 (N_10896,N_6149,N_6870);
or U10897 (N_10897,N_8936,N_7093);
xnor U10898 (N_10898,N_8664,N_7132);
nor U10899 (N_10899,N_6829,N_7635);
nor U10900 (N_10900,N_6340,N_7337);
and U10901 (N_10901,N_8671,N_7570);
xor U10902 (N_10902,N_7507,N_6083);
or U10903 (N_10903,N_6201,N_7712);
nand U10904 (N_10904,N_7465,N_6174);
or U10905 (N_10905,N_7114,N_8536);
xnor U10906 (N_10906,N_8160,N_7004);
xnor U10907 (N_10907,N_7696,N_8408);
xor U10908 (N_10908,N_7456,N_6777);
or U10909 (N_10909,N_8361,N_6487);
and U10910 (N_10910,N_8110,N_8065);
nand U10911 (N_10911,N_8204,N_6801);
and U10912 (N_10912,N_6052,N_8850);
nor U10913 (N_10913,N_6289,N_6917);
nor U10914 (N_10914,N_6716,N_8248);
xnor U10915 (N_10915,N_8370,N_8975);
nor U10916 (N_10916,N_8623,N_6859);
nand U10917 (N_10917,N_8756,N_8982);
nand U10918 (N_10918,N_7020,N_8965);
or U10919 (N_10919,N_8726,N_7942);
nand U10920 (N_10920,N_7316,N_7705);
nor U10921 (N_10921,N_6303,N_6966);
and U10922 (N_10922,N_7563,N_6542);
nand U10923 (N_10923,N_7216,N_7906);
and U10924 (N_10924,N_6492,N_7924);
xor U10925 (N_10925,N_6625,N_6532);
nand U10926 (N_10926,N_7289,N_7420);
nor U10927 (N_10927,N_7654,N_7172);
and U10928 (N_10928,N_8691,N_8990);
xnor U10929 (N_10929,N_8289,N_7042);
xor U10930 (N_10930,N_7755,N_8302);
or U10931 (N_10931,N_6151,N_6552);
nand U10932 (N_10932,N_6442,N_6607);
or U10933 (N_10933,N_8509,N_6280);
or U10934 (N_10934,N_6986,N_8554);
nand U10935 (N_10935,N_8213,N_6642);
xnor U10936 (N_10936,N_6361,N_6723);
and U10937 (N_10937,N_7255,N_8622);
xnor U10938 (N_10938,N_6923,N_6986);
nand U10939 (N_10939,N_7478,N_6337);
nor U10940 (N_10940,N_7775,N_8664);
and U10941 (N_10941,N_8062,N_7429);
xor U10942 (N_10942,N_8754,N_7395);
nand U10943 (N_10943,N_6594,N_6890);
or U10944 (N_10944,N_6687,N_6300);
nor U10945 (N_10945,N_6034,N_8743);
nor U10946 (N_10946,N_7961,N_8551);
xor U10947 (N_10947,N_8563,N_7387);
xnor U10948 (N_10948,N_6690,N_8411);
nor U10949 (N_10949,N_8305,N_6541);
and U10950 (N_10950,N_8608,N_8152);
nor U10951 (N_10951,N_8981,N_6971);
nor U10952 (N_10952,N_7309,N_8665);
xor U10953 (N_10953,N_7335,N_7089);
nor U10954 (N_10954,N_8486,N_7526);
nand U10955 (N_10955,N_8033,N_7179);
and U10956 (N_10956,N_7521,N_8384);
or U10957 (N_10957,N_6854,N_8836);
nand U10958 (N_10958,N_6581,N_7290);
xnor U10959 (N_10959,N_8051,N_8431);
nor U10960 (N_10960,N_8696,N_6631);
xnor U10961 (N_10961,N_8984,N_7782);
nand U10962 (N_10962,N_8603,N_6350);
nor U10963 (N_10963,N_7258,N_6986);
xor U10964 (N_10964,N_6453,N_7559);
nand U10965 (N_10965,N_7602,N_6136);
xnor U10966 (N_10966,N_6296,N_8725);
or U10967 (N_10967,N_8520,N_6352);
or U10968 (N_10968,N_7462,N_6798);
nor U10969 (N_10969,N_6238,N_8428);
or U10970 (N_10970,N_7821,N_7357);
or U10971 (N_10971,N_8947,N_6156);
xor U10972 (N_10972,N_6150,N_6309);
or U10973 (N_10973,N_8607,N_8823);
or U10974 (N_10974,N_6529,N_7881);
xor U10975 (N_10975,N_6659,N_7546);
and U10976 (N_10976,N_8391,N_8923);
nor U10977 (N_10977,N_6802,N_8427);
nand U10978 (N_10978,N_6600,N_8535);
and U10979 (N_10979,N_7850,N_8572);
or U10980 (N_10980,N_8014,N_7210);
xor U10981 (N_10981,N_6263,N_6647);
xnor U10982 (N_10982,N_8290,N_6874);
nand U10983 (N_10983,N_8828,N_7315);
xor U10984 (N_10984,N_6952,N_8041);
nor U10985 (N_10985,N_7272,N_8916);
or U10986 (N_10986,N_8130,N_7527);
nand U10987 (N_10987,N_7892,N_6825);
nand U10988 (N_10988,N_7347,N_8248);
or U10989 (N_10989,N_6825,N_7528);
nand U10990 (N_10990,N_7643,N_7977);
nand U10991 (N_10991,N_6279,N_7836);
nand U10992 (N_10992,N_8918,N_6943);
nand U10993 (N_10993,N_6864,N_8171);
xor U10994 (N_10994,N_8128,N_8983);
nor U10995 (N_10995,N_6280,N_7336);
nand U10996 (N_10996,N_8781,N_7222);
and U10997 (N_10997,N_6485,N_6055);
and U10998 (N_10998,N_7237,N_7644);
nand U10999 (N_10999,N_7624,N_8227);
xor U11000 (N_11000,N_8822,N_6709);
xnor U11001 (N_11001,N_8931,N_8850);
xor U11002 (N_11002,N_7775,N_7829);
nor U11003 (N_11003,N_7025,N_6553);
nand U11004 (N_11004,N_8287,N_8572);
and U11005 (N_11005,N_7345,N_6178);
xnor U11006 (N_11006,N_8164,N_8144);
and U11007 (N_11007,N_8444,N_7152);
nor U11008 (N_11008,N_6930,N_8014);
or U11009 (N_11009,N_8927,N_7268);
nor U11010 (N_11010,N_7921,N_6418);
xor U11011 (N_11011,N_7804,N_6130);
xor U11012 (N_11012,N_8213,N_7772);
xor U11013 (N_11013,N_7128,N_6936);
nor U11014 (N_11014,N_6997,N_7004);
xnor U11015 (N_11015,N_6168,N_6504);
xor U11016 (N_11016,N_8866,N_8160);
and U11017 (N_11017,N_7875,N_8691);
or U11018 (N_11018,N_8489,N_7541);
and U11019 (N_11019,N_7723,N_6045);
and U11020 (N_11020,N_6019,N_7328);
xnor U11021 (N_11021,N_7992,N_7448);
nand U11022 (N_11022,N_7189,N_8388);
or U11023 (N_11023,N_7470,N_7219);
or U11024 (N_11024,N_7616,N_7827);
or U11025 (N_11025,N_6174,N_6277);
xor U11026 (N_11026,N_6385,N_7467);
nand U11027 (N_11027,N_6889,N_7886);
or U11028 (N_11028,N_8263,N_8254);
or U11029 (N_11029,N_6934,N_8127);
and U11030 (N_11030,N_6601,N_8591);
or U11031 (N_11031,N_8488,N_7244);
or U11032 (N_11032,N_8711,N_6466);
xnor U11033 (N_11033,N_6406,N_6695);
nand U11034 (N_11034,N_8373,N_7367);
and U11035 (N_11035,N_7039,N_6566);
and U11036 (N_11036,N_7037,N_8666);
and U11037 (N_11037,N_6723,N_6469);
xor U11038 (N_11038,N_8127,N_8467);
xnor U11039 (N_11039,N_8439,N_7557);
or U11040 (N_11040,N_8118,N_8810);
or U11041 (N_11041,N_8048,N_6190);
and U11042 (N_11042,N_7954,N_8694);
or U11043 (N_11043,N_6675,N_6770);
xnor U11044 (N_11044,N_7874,N_7658);
nand U11045 (N_11045,N_7600,N_6152);
or U11046 (N_11046,N_6462,N_7128);
nand U11047 (N_11047,N_7219,N_6343);
or U11048 (N_11048,N_7486,N_7839);
or U11049 (N_11049,N_6068,N_8092);
nand U11050 (N_11050,N_7740,N_7750);
nand U11051 (N_11051,N_8839,N_8347);
nand U11052 (N_11052,N_6262,N_6663);
or U11053 (N_11053,N_6779,N_8396);
and U11054 (N_11054,N_6378,N_7047);
xnor U11055 (N_11055,N_6022,N_8029);
nand U11056 (N_11056,N_7632,N_7438);
and U11057 (N_11057,N_7499,N_6273);
nor U11058 (N_11058,N_8706,N_6044);
xnor U11059 (N_11059,N_7967,N_6525);
or U11060 (N_11060,N_7457,N_8121);
or U11061 (N_11061,N_6585,N_6289);
and U11062 (N_11062,N_8738,N_8575);
nor U11063 (N_11063,N_7491,N_6717);
and U11064 (N_11064,N_8307,N_8876);
xnor U11065 (N_11065,N_7927,N_7279);
or U11066 (N_11066,N_7496,N_7899);
nand U11067 (N_11067,N_8952,N_7693);
nand U11068 (N_11068,N_8205,N_8921);
or U11069 (N_11069,N_7579,N_7361);
or U11070 (N_11070,N_6740,N_8776);
xor U11071 (N_11071,N_6888,N_7196);
and U11072 (N_11072,N_6352,N_6109);
xnor U11073 (N_11073,N_8248,N_6305);
xnor U11074 (N_11074,N_7480,N_8858);
nor U11075 (N_11075,N_7824,N_6908);
nand U11076 (N_11076,N_8300,N_6925);
or U11077 (N_11077,N_7684,N_8852);
xor U11078 (N_11078,N_6538,N_7832);
xor U11079 (N_11079,N_8955,N_6596);
nand U11080 (N_11080,N_7241,N_6775);
nand U11081 (N_11081,N_7569,N_6947);
xnor U11082 (N_11082,N_7731,N_8287);
nor U11083 (N_11083,N_8243,N_8130);
nand U11084 (N_11084,N_8881,N_8627);
xnor U11085 (N_11085,N_8240,N_7614);
nor U11086 (N_11086,N_6522,N_7810);
nor U11087 (N_11087,N_7125,N_6525);
and U11088 (N_11088,N_7090,N_6243);
or U11089 (N_11089,N_8920,N_8174);
and U11090 (N_11090,N_7286,N_6690);
nand U11091 (N_11091,N_7990,N_6713);
xnor U11092 (N_11092,N_7407,N_8912);
and U11093 (N_11093,N_7699,N_8535);
nor U11094 (N_11094,N_7985,N_6336);
or U11095 (N_11095,N_8840,N_7540);
or U11096 (N_11096,N_7044,N_7329);
and U11097 (N_11097,N_8929,N_6966);
nand U11098 (N_11098,N_6467,N_8297);
and U11099 (N_11099,N_8832,N_8451);
nor U11100 (N_11100,N_8817,N_8632);
and U11101 (N_11101,N_8713,N_8343);
and U11102 (N_11102,N_7471,N_7073);
nand U11103 (N_11103,N_7182,N_8871);
nor U11104 (N_11104,N_6072,N_8149);
xnor U11105 (N_11105,N_6208,N_8214);
or U11106 (N_11106,N_7215,N_7624);
xnor U11107 (N_11107,N_7942,N_6372);
xnor U11108 (N_11108,N_8296,N_8554);
nand U11109 (N_11109,N_6651,N_6855);
nand U11110 (N_11110,N_7844,N_8072);
nand U11111 (N_11111,N_6622,N_6561);
xor U11112 (N_11112,N_8009,N_8976);
xnor U11113 (N_11113,N_7236,N_6855);
and U11114 (N_11114,N_7387,N_7543);
nor U11115 (N_11115,N_7992,N_8552);
nor U11116 (N_11116,N_8676,N_8112);
xnor U11117 (N_11117,N_6277,N_7424);
xnor U11118 (N_11118,N_8919,N_7504);
nand U11119 (N_11119,N_6821,N_6153);
xor U11120 (N_11120,N_8183,N_6885);
nand U11121 (N_11121,N_7231,N_6186);
nand U11122 (N_11122,N_8192,N_7890);
nand U11123 (N_11123,N_7844,N_6035);
nand U11124 (N_11124,N_6055,N_6511);
or U11125 (N_11125,N_8114,N_8959);
and U11126 (N_11126,N_8785,N_7619);
xnor U11127 (N_11127,N_8064,N_6291);
nand U11128 (N_11128,N_7853,N_7215);
or U11129 (N_11129,N_6046,N_6157);
or U11130 (N_11130,N_8360,N_6431);
nor U11131 (N_11131,N_8309,N_8179);
or U11132 (N_11132,N_7328,N_7678);
nor U11133 (N_11133,N_6716,N_6134);
nor U11134 (N_11134,N_8719,N_6245);
and U11135 (N_11135,N_7530,N_8680);
nand U11136 (N_11136,N_6487,N_7011);
xnor U11137 (N_11137,N_7250,N_6653);
and U11138 (N_11138,N_8658,N_7043);
or U11139 (N_11139,N_6950,N_6722);
xor U11140 (N_11140,N_7983,N_7289);
and U11141 (N_11141,N_8105,N_7882);
or U11142 (N_11142,N_7607,N_6226);
or U11143 (N_11143,N_6823,N_7607);
xnor U11144 (N_11144,N_8241,N_6183);
and U11145 (N_11145,N_7840,N_7866);
nand U11146 (N_11146,N_7879,N_8260);
nor U11147 (N_11147,N_8517,N_7086);
and U11148 (N_11148,N_7028,N_8232);
xor U11149 (N_11149,N_7025,N_6062);
xnor U11150 (N_11150,N_7842,N_6399);
and U11151 (N_11151,N_8199,N_7795);
nor U11152 (N_11152,N_7579,N_8118);
and U11153 (N_11153,N_8905,N_7481);
nand U11154 (N_11154,N_8774,N_8284);
xnor U11155 (N_11155,N_6151,N_8982);
or U11156 (N_11156,N_8927,N_7456);
nand U11157 (N_11157,N_8945,N_6247);
xnor U11158 (N_11158,N_6517,N_7976);
or U11159 (N_11159,N_8957,N_7635);
nor U11160 (N_11160,N_6679,N_6201);
and U11161 (N_11161,N_8958,N_6417);
nand U11162 (N_11162,N_7440,N_8082);
or U11163 (N_11163,N_7225,N_7717);
nand U11164 (N_11164,N_6684,N_7793);
nor U11165 (N_11165,N_8001,N_7168);
nand U11166 (N_11166,N_6958,N_8129);
or U11167 (N_11167,N_6711,N_7805);
or U11168 (N_11168,N_7666,N_6820);
nand U11169 (N_11169,N_7808,N_7169);
nand U11170 (N_11170,N_8778,N_7632);
xor U11171 (N_11171,N_6213,N_8761);
xor U11172 (N_11172,N_7226,N_7471);
and U11173 (N_11173,N_7817,N_7456);
xnor U11174 (N_11174,N_6558,N_6630);
nand U11175 (N_11175,N_6662,N_7687);
nor U11176 (N_11176,N_6865,N_8926);
nor U11177 (N_11177,N_6076,N_8214);
or U11178 (N_11178,N_8843,N_7607);
nand U11179 (N_11179,N_7912,N_7863);
nor U11180 (N_11180,N_6641,N_6845);
nor U11181 (N_11181,N_7395,N_8455);
nand U11182 (N_11182,N_7564,N_6031);
and U11183 (N_11183,N_7296,N_7219);
xnor U11184 (N_11184,N_7856,N_8271);
nor U11185 (N_11185,N_7218,N_7526);
nor U11186 (N_11186,N_6311,N_7096);
xor U11187 (N_11187,N_7927,N_6058);
nand U11188 (N_11188,N_8275,N_6908);
nor U11189 (N_11189,N_8081,N_8082);
xor U11190 (N_11190,N_7741,N_6052);
and U11191 (N_11191,N_6030,N_6933);
nand U11192 (N_11192,N_7022,N_8735);
or U11193 (N_11193,N_8916,N_8045);
nand U11194 (N_11194,N_8709,N_7789);
xnor U11195 (N_11195,N_6412,N_7847);
nand U11196 (N_11196,N_6056,N_7108);
nor U11197 (N_11197,N_6423,N_6691);
and U11198 (N_11198,N_6649,N_7925);
or U11199 (N_11199,N_8253,N_8149);
or U11200 (N_11200,N_7380,N_8539);
or U11201 (N_11201,N_7679,N_8531);
and U11202 (N_11202,N_8937,N_6255);
or U11203 (N_11203,N_8235,N_8915);
nor U11204 (N_11204,N_6528,N_8022);
nand U11205 (N_11205,N_7410,N_6003);
nor U11206 (N_11206,N_8227,N_8901);
nor U11207 (N_11207,N_6045,N_8851);
nand U11208 (N_11208,N_7069,N_8590);
nor U11209 (N_11209,N_8216,N_6906);
and U11210 (N_11210,N_8091,N_8158);
or U11211 (N_11211,N_8458,N_6677);
and U11212 (N_11212,N_6231,N_7365);
xor U11213 (N_11213,N_7356,N_8608);
nor U11214 (N_11214,N_6713,N_7049);
xor U11215 (N_11215,N_6731,N_7585);
and U11216 (N_11216,N_8680,N_6488);
nand U11217 (N_11217,N_7228,N_8625);
nand U11218 (N_11218,N_6624,N_7207);
or U11219 (N_11219,N_6358,N_7635);
and U11220 (N_11220,N_7546,N_7439);
or U11221 (N_11221,N_7798,N_6186);
or U11222 (N_11222,N_8671,N_8427);
and U11223 (N_11223,N_8764,N_8719);
nand U11224 (N_11224,N_8048,N_7992);
xor U11225 (N_11225,N_7210,N_6075);
or U11226 (N_11226,N_8416,N_7360);
xnor U11227 (N_11227,N_6757,N_8636);
and U11228 (N_11228,N_8632,N_6086);
nor U11229 (N_11229,N_7321,N_6695);
nand U11230 (N_11230,N_8453,N_8165);
nand U11231 (N_11231,N_8666,N_7328);
or U11232 (N_11232,N_8003,N_6175);
nand U11233 (N_11233,N_6745,N_8273);
nor U11234 (N_11234,N_7614,N_8448);
xor U11235 (N_11235,N_8641,N_8276);
nand U11236 (N_11236,N_6205,N_8983);
nand U11237 (N_11237,N_7152,N_7442);
nor U11238 (N_11238,N_6351,N_6878);
nor U11239 (N_11239,N_8817,N_7406);
nand U11240 (N_11240,N_6476,N_6148);
xnor U11241 (N_11241,N_6813,N_7343);
nand U11242 (N_11242,N_7869,N_7233);
and U11243 (N_11243,N_7414,N_8716);
xor U11244 (N_11244,N_7310,N_8952);
nand U11245 (N_11245,N_8393,N_7242);
nand U11246 (N_11246,N_6962,N_7335);
or U11247 (N_11247,N_7615,N_8771);
and U11248 (N_11248,N_6902,N_8677);
xnor U11249 (N_11249,N_7822,N_6721);
or U11250 (N_11250,N_8475,N_6100);
nand U11251 (N_11251,N_8924,N_6107);
and U11252 (N_11252,N_8747,N_8071);
or U11253 (N_11253,N_7598,N_8561);
xnor U11254 (N_11254,N_6202,N_6367);
nor U11255 (N_11255,N_8935,N_7889);
and U11256 (N_11256,N_7351,N_8065);
and U11257 (N_11257,N_8489,N_6349);
nor U11258 (N_11258,N_7633,N_6024);
xor U11259 (N_11259,N_8069,N_8573);
or U11260 (N_11260,N_8612,N_6818);
nand U11261 (N_11261,N_8975,N_8757);
xor U11262 (N_11262,N_8102,N_8792);
xnor U11263 (N_11263,N_8763,N_7428);
or U11264 (N_11264,N_8073,N_7254);
xnor U11265 (N_11265,N_7209,N_8994);
and U11266 (N_11266,N_8211,N_7808);
nand U11267 (N_11267,N_7644,N_7975);
xor U11268 (N_11268,N_8447,N_8425);
and U11269 (N_11269,N_6192,N_7479);
and U11270 (N_11270,N_8901,N_7268);
nand U11271 (N_11271,N_8002,N_6109);
nor U11272 (N_11272,N_6008,N_6658);
nor U11273 (N_11273,N_7261,N_8485);
or U11274 (N_11274,N_7273,N_7168);
nor U11275 (N_11275,N_7505,N_6077);
and U11276 (N_11276,N_7760,N_8207);
xor U11277 (N_11277,N_8112,N_7464);
nand U11278 (N_11278,N_6034,N_7276);
nand U11279 (N_11279,N_8657,N_7330);
nand U11280 (N_11280,N_6947,N_8681);
xnor U11281 (N_11281,N_8221,N_7119);
or U11282 (N_11282,N_6055,N_6967);
and U11283 (N_11283,N_8113,N_6315);
nor U11284 (N_11284,N_8760,N_6315);
and U11285 (N_11285,N_6932,N_8899);
xnor U11286 (N_11286,N_7057,N_7843);
nand U11287 (N_11287,N_8604,N_6701);
nor U11288 (N_11288,N_8779,N_6218);
and U11289 (N_11289,N_8116,N_6528);
nor U11290 (N_11290,N_8331,N_7740);
and U11291 (N_11291,N_8102,N_8107);
xnor U11292 (N_11292,N_7501,N_6055);
nor U11293 (N_11293,N_6301,N_8050);
nor U11294 (N_11294,N_7180,N_8724);
nand U11295 (N_11295,N_8874,N_6772);
or U11296 (N_11296,N_7597,N_6999);
or U11297 (N_11297,N_6972,N_6110);
xor U11298 (N_11298,N_6945,N_6050);
xor U11299 (N_11299,N_8728,N_8440);
nand U11300 (N_11300,N_7701,N_7628);
and U11301 (N_11301,N_7295,N_6067);
and U11302 (N_11302,N_6461,N_7877);
nand U11303 (N_11303,N_6024,N_7113);
or U11304 (N_11304,N_8210,N_6410);
nand U11305 (N_11305,N_8285,N_6823);
xor U11306 (N_11306,N_8096,N_6999);
or U11307 (N_11307,N_6983,N_6166);
and U11308 (N_11308,N_8337,N_7740);
nand U11309 (N_11309,N_7836,N_7260);
xnor U11310 (N_11310,N_7875,N_6574);
nand U11311 (N_11311,N_8757,N_6373);
nand U11312 (N_11312,N_6389,N_8859);
xnor U11313 (N_11313,N_7396,N_8403);
nand U11314 (N_11314,N_8095,N_6443);
nand U11315 (N_11315,N_8297,N_7972);
nand U11316 (N_11316,N_8699,N_7758);
nor U11317 (N_11317,N_8916,N_7770);
and U11318 (N_11318,N_8943,N_7816);
and U11319 (N_11319,N_6506,N_7115);
xor U11320 (N_11320,N_8976,N_6801);
or U11321 (N_11321,N_6533,N_8824);
nor U11322 (N_11322,N_7583,N_7611);
nor U11323 (N_11323,N_6693,N_8092);
nor U11324 (N_11324,N_7420,N_6849);
xnor U11325 (N_11325,N_8859,N_8798);
nor U11326 (N_11326,N_7208,N_8520);
or U11327 (N_11327,N_6691,N_6104);
and U11328 (N_11328,N_7254,N_8053);
nor U11329 (N_11329,N_8786,N_8327);
or U11330 (N_11330,N_7165,N_7996);
or U11331 (N_11331,N_6140,N_7762);
and U11332 (N_11332,N_6737,N_6817);
or U11333 (N_11333,N_8765,N_8281);
nor U11334 (N_11334,N_8639,N_8693);
nand U11335 (N_11335,N_6378,N_6042);
or U11336 (N_11336,N_6822,N_8488);
nor U11337 (N_11337,N_8288,N_8507);
and U11338 (N_11338,N_7207,N_7407);
nand U11339 (N_11339,N_7361,N_7833);
and U11340 (N_11340,N_7123,N_7296);
nand U11341 (N_11341,N_7033,N_7169);
xnor U11342 (N_11342,N_6349,N_7012);
and U11343 (N_11343,N_8767,N_7339);
and U11344 (N_11344,N_7664,N_6959);
xnor U11345 (N_11345,N_6549,N_6630);
or U11346 (N_11346,N_7333,N_6634);
xnor U11347 (N_11347,N_8055,N_6083);
nand U11348 (N_11348,N_7662,N_8290);
nand U11349 (N_11349,N_7592,N_6795);
xnor U11350 (N_11350,N_7198,N_7155);
nand U11351 (N_11351,N_7067,N_6521);
or U11352 (N_11352,N_6635,N_8923);
nor U11353 (N_11353,N_7822,N_8152);
xnor U11354 (N_11354,N_6768,N_7698);
nor U11355 (N_11355,N_8918,N_8025);
nor U11356 (N_11356,N_6661,N_6021);
and U11357 (N_11357,N_8363,N_7327);
and U11358 (N_11358,N_8243,N_6312);
and U11359 (N_11359,N_8225,N_8370);
nand U11360 (N_11360,N_8874,N_7625);
nor U11361 (N_11361,N_6392,N_7126);
and U11362 (N_11362,N_6618,N_6663);
nor U11363 (N_11363,N_7292,N_6039);
nand U11364 (N_11364,N_6607,N_8391);
xnor U11365 (N_11365,N_7692,N_6147);
and U11366 (N_11366,N_6229,N_7188);
and U11367 (N_11367,N_6424,N_7500);
and U11368 (N_11368,N_7681,N_7941);
nand U11369 (N_11369,N_6425,N_6962);
nand U11370 (N_11370,N_7130,N_8504);
xnor U11371 (N_11371,N_6644,N_6614);
or U11372 (N_11372,N_7140,N_6400);
and U11373 (N_11373,N_7823,N_7204);
nor U11374 (N_11374,N_6270,N_8413);
xor U11375 (N_11375,N_6613,N_7718);
nor U11376 (N_11376,N_7860,N_8098);
nand U11377 (N_11377,N_8303,N_8552);
nor U11378 (N_11378,N_6002,N_8694);
and U11379 (N_11379,N_6162,N_7911);
nor U11380 (N_11380,N_6011,N_8341);
and U11381 (N_11381,N_8259,N_8304);
nand U11382 (N_11382,N_6632,N_6228);
xnor U11383 (N_11383,N_7364,N_8541);
and U11384 (N_11384,N_7105,N_8157);
xor U11385 (N_11385,N_7014,N_6182);
and U11386 (N_11386,N_8291,N_6366);
xnor U11387 (N_11387,N_6929,N_6924);
or U11388 (N_11388,N_6224,N_7279);
and U11389 (N_11389,N_7186,N_6798);
xor U11390 (N_11390,N_6463,N_7270);
and U11391 (N_11391,N_6777,N_8123);
xor U11392 (N_11392,N_8870,N_7640);
xor U11393 (N_11393,N_8272,N_8768);
xor U11394 (N_11394,N_6318,N_8651);
nor U11395 (N_11395,N_6413,N_6251);
nor U11396 (N_11396,N_7696,N_6634);
xnor U11397 (N_11397,N_6232,N_8952);
xor U11398 (N_11398,N_7123,N_7578);
nor U11399 (N_11399,N_8112,N_6887);
and U11400 (N_11400,N_7723,N_6257);
or U11401 (N_11401,N_7017,N_6434);
xor U11402 (N_11402,N_7206,N_6397);
or U11403 (N_11403,N_8110,N_8461);
nor U11404 (N_11404,N_8215,N_6976);
xor U11405 (N_11405,N_7648,N_8531);
or U11406 (N_11406,N_8406,N_6888);
nor U11407 (N_11407,N_6119,N_6438);
nand U11408 (N_11408,N_8746,N_8575);
nor U11409 (N_11409,N_6330,N_6712);
and U11410 (N_11410,N_7339,N_6067);
and U11411 (N_11411,N_6933,N_6395);
nand U11412 (N_11412,N_7309,N_8344);
or U11413 (N_11413,N_8559,N_7924);
nand U11414 (N_11414,N_8357,N_6952);
nor U11415 (N_11415,N_7853,N_8380);
xor U11416 (N_11416,N_7341,N_7631);
nand U11417 (N_11417,N_7954,N_7696);
or U11418 (N_11418,N_6599,N_6814);
xor U11419 (N_11419,N_6789,N_6645);
xnor U11420 (N_11420,N_8031,N_7068);
or U11421 (N_11421,N_6988,N_8281);
xnor U11422 (N_11422,N_6306,N_7943);
or U11423 (N_11423,N_8531,N_8470);
xor U11424 (N_11424,N_8550,N_6654);
and U11425 (N_11425,N_6793,N_6068);
nor U11426 (N_11426,N_8925,N_7730);
nor U11427 (N_11427,N_8591,N_7833);
or U11428 (N_11428,N_7338,N_8711);
xor U11429 (N_11429,N_7735,N_8397);
nor U11430 (N_11430,N_7479,N_6745);
or U11431 (N_11431,N_8978,N_7169);
nand U11432 (N_11432,N_6035,N_8831);
nor U11433 (N_11433,N_6254,N_7770);
or U11434 (N_11434,N_6864,N_6609);
nor U11435 (N_11435,N_8935,N_6820);
nor U11436 (N_11436,N_7700,N_6303);
xnor U11437 (N_11437,N_6751,N_8299);
nor U11438 (N_11438,N_6901,N_6718);
xor U11439 (N_11439,N_6082,N_6551);
and U11440 (N_11440,N_6609,N_8392);
or U11441 (N_11441,N_6331,N_7908);
nand U11442 (N_11442,N_7691,N_6253);
nor U11443 (N_11443,N_7836,N_8927);
nor U11444 (N_11444,N_8419,N_6090);
nand U11445 (N_11445,N_7814,N_8765);
nor U11446 (N_11446,N_7152,N_7308);
or U11447 (N_11447,N_8315,N_7536);
or U11448 (N_11448,N_7991,N_6740);
nand U11449 (N_11449,N_8348,N_7068);
nor U11450 (N_11450,N_6960,N_8172);
or U11451 (N_11451,N_8592,N_6366);
nand U11452 (N_11452,N_7722,N_8959);
nor U11453 (N_11453,N_7757,N_7858);
and U11454 (N_11454,N_8265,N_8388);
xnor U11455 (N_11455,N_8056,N_8959);
and U11456 (N_11456,N_6348,N_8761);
and U11457 (N_11457,N_7219,N_6552);
nand U11458 (N_11458,N_7933,N_8825);
and U11459 (N_11459,N_7899,N_8404);
nand U11460 (N_11460,N_7379,N_6427);
nor U11461 (N_11461,N_6499,N_7719);
xnor U11462 (N_11462,N_6258,N_6003);
xor U11463 (N_11463,N_7155,N_7328);
nand U11464 (N_11464,N_6278,N_6999);
nand U11465 (N_11465,N_7455,N_7097);
and U11466 (N_11466,N_6664,N_8017);
nor U11467 (N_11467,N_6421,N_8095);
or U11468 (N_11468,N_7973,N_7082);
xor U11469 (N_11469,N_6191,N_6572);
xnor U11470 (N_11470,N_7773,N_8387);
and U11471 (N_11471,N_6365,N_8960);
nor U11472 (N_11472,N_6809,N_8408);
nor U11473 (N_11473,N_7186,N_7295);
nand U11474 (N_11474,N_7430,N_8388);
and U11475 (N_11475,N_8554,N_7590);
xor U11476 (N_11476,N_6220,N_6567);
or U11477 (N_11477,N_7490,N_6785);
or U11478 (N_11478,N_6882,N_8144);
xnor U11479 (N_11479,N_8316,N_7269);
nand U11480 (N_11480,N_6332,N_8265);
and U11481 (N_11481,N_8903,N_7277);
and U11482 (N_11482,N_8136,N_6681);
or U11483 (N_11483,N_8974,N_7978);
xnor U11484 (N_11484,N_6997,N_6127);
or U11485 (N_11485,N_7374,N_7210);
or U11486 (N_11486,N_6522,N_8719);
nand U11487 (N_11487,N_7133,N_8969);
or U11488 (N_11488,N_8896,N_8376);
or U11489 (N_11489,N_6709,N_6939);
xnor U11490 (N_11490,N_7235,N_6430);
or U11491 (N_11491,N_6534,N_7592);
xor U11492 (N_11492,N_6368,N_6485);
xnor U11493 (N_11493,N_7868,N_6188);
or U11494 (N_11494,N_7797,N_7594);
nor U11495 (N_11495,N_7089,N_8864);
xnor U11496 (N_11496,N_6332,N_7395);
or U11497 (N_11497,N_6700,N_6928);
nand U11498 (N_11498,N_7031,N_8308);
nor U11499 (N_11499,N_8199,N_6944);
and U11500 (N_11500,N_8298,N_7184);
nand U11501 (N_11501,N_8751,N_7035);
and U11502 (N_11502,N_8517,N_8000);
and U11503 (N_11503,N_7486,N_8711);
or U11504 (N_11504,N_6740,N_6358);
nand U11505 (N_11505,N_6283,N_6109);
nor U11506 (N_11506,N_6302,N_7214);
or U11507 (N_11507,N_7482,N_8623);
and U11508 (N_11508,N_7512,N_7056);
xor U11509 (N_11509,N_8356,N_7022);
nand U11510 (N_11510,N_8730,N_6474);
nor U11511 (N_11511,N_8922,N_8041);
and U11512 (N_11512,N_8126,N_7747);
nor U11513 (N_11513,N_8594,N_6075);
or U11514 (N_11514,N_6596,N_6782);
or U11515 (N_11515,N_6687,N_7080);
xnor U11516 (N_11516,N_6932,N_7290);
or U11517 (N_11517,N_6651,N_6379);
nor U11518 (N_11518,N_6810,N_8962);
xnor U11519 (N_11519,N_6015,N_6626);
nor U11520 (N_11520,N_7302,N_8054);
nand U11521 (N_11521,N_8099,N_7432);
nor U11522 (N_11522,N_7107,N_6735);
nand U11523 (N_11523,N_8103,N_6292);
and U11524 (N_11524,N_8991,N_6750);
and U11525 (N_11525,N_6602,N_7598);
xnor U11526 (N_11526,N_8913,N_8592);
xor U11527 (N_11527,N_8280,N_6649);
nor U11528 (N_11528,N_8706,N_7390);
and U11529 (N_11529,N_6150,N_8006);
and U11530 (N_11530,N_7129,N_6931);
xnor U11531 (N_11531,N_6967,N_8757);
xor U11532 (N_11532,N_8155,N_8938);
nand U11533 (N_11533,N_6746,N_8056);
xor U11534 (N_11534,N_8144,N_6699);
xnor U11535 (N_11535,N_8942,N_8732);
or U11536 (N_11536,N_7656,N_7066);
xnor U11537 (N_11537,N_6561,N_6346);
or U11538 (N_11538,N_7443,N_7636);
nand U11539 (N_11539,N_6685,N_7772);
nor U11540 (N_11540,N_6816,N_7420);
xor U11541 (N_11541,N_8120,N_8676);
nand U11542 (N_11542,N_7689,N_6170);
nor U11543 (N_11543,N_8187,N_8510);
nand U11544 (N_11544,N_7420,N_8324);
nor U11545 (N_11545,N_6238,N_7847);
and U11546 (N_11546,N_6993,N_8036);
xor U11547 (N_11547,N_6636,N_8019);
and U11548 (N_11548,N_7210,N_7375);
nand U11549 (N_11549,N_8949,N_8464);
xor U11550 (N_11550,N_8557,N_7899);
or U11551 (N_11551,N_6763,N_6099);
nand U11552 (N_11552,N_6803,N_8839);
xor U11553 (N_11553,N_6647,N_8483);
nor U11554 (N_11554,N_7641,N_8662);
nor U11555 (N_11555,N_7997,N_7681);
and U11556 (N_11556,N_8923,N_6045);
nand U11557 (N_11557,N_8809,N_7058);
and U11558 (N_11558,N_6869,N_8728);
nor U11559 (N_11559,N_6410,N_6682);
nand U11560 (N_11560,N_6156,N_8334);
xor U11561 (N_11561,N_6479,N_7300);
and U11562 (N_11562,N_6370,N_8596);
xnor U11563 (N_11563,N_6818,N_8022);
or U11564 (N_11564,N_8516,N_8778);
xor U11565 (N_11565,N_6520,N_6241);
nand U11566 (N_11566,N_7781,N_6651);
nor U11567 (N_11567,N_7453,N_8171);
nand U11568 (N_11568,N_8830,N_8351);
and U11569 (N_11569,N_8152,N_6212);
nor U11570 (N_11570,N_7552,N_8722);
nor U11571 (N_11571,N_8126,N_7978);
and U11572 (N_11572,N_7497,N_6477);
nor U11573 (N_11573,N_7535,N_7037);
and U11574 (N_11574,N_8727,N_8349);
or U11575 (N_11575,N_7756,N_8949);
and U11576 (N_11576,N_7551,N_6649);
nor U11577 (N_11577,N_6845,N_8496);
xor U11578 (N_11578,N_8844,N_8160);
nand U11579 (N_11579,N_6406,N_7066);
nor U11580 (N_11580,N_8228,N_8575);
xnor U11581 (N_11581,N_7219,N_8090);
or U11582 (N_11582,N_7369,N_6946);
nor U11583 (N_11583,N_8436,N_7693);
or U11584 (N_11584,N_7921,N_6885);
xor U11585 (N_11585,N_8582,N_8817);
nor U11586 (N_11586,N_6455,N_7417);
nor U11587 (N_11587,N_8298,N_7679);
nand U11588 (N_11588,N_7113,N_8578);
nand U11589 (N_11589,N_8451,N_6669);
xnor U11590 (N_11590,N_6931,N_8634);
nor U11591 (N_11591,N_8669,N_7977);
xor U11592 (N_11592,N_6556,N_6454);
and U11593 (N_11593,N_8129,N_6731);
and U11594 (N_11594,N_7381,N_6043);
or U11595 (N_11595,N_6961,N_7859);
nand U11596 (N_11596,N_8795,N_6755);
nor U11597 (N_11597,N_6012,N_7487);
or U11598 (N_11598,N_6118,N_8702);
nand U11599 (N_11599,N_6434,N_6344);
xnor U11600 (N_11600,N_7212,N_6452);
nand U11601 (N_11601,N_6549,N_7786);
and U11602 (N_11602,N_8885,N_7914);
xor U11603 (N_11603,N_7888,N_8337);
nor U11604 (N_11604,N_8652,N_8378);
or U11605 (N_11605,N_6465,N_7563);
nor U11606 (N_11606,N_8464,N_8790);
nor U11607 (N_11607,N_6823,N_6980);
nor U11608 (N_11608,N_6202,N_6724);
nand U11609 (N_11609,N_7424,N_8714);
or U11610 (N_11610,N_7860,N_7498);
and U11611 (N_11611,N_8888,N_8952);
xnor U11612 (N_11612,N_8286,N_7202);
or U11613 (N_11613,N_8962,N_6410);
and U11614 (N_11614,N_8059,N_8462);
xnor U11615 (N_11615,N_8287,N_8317);
xor U11616 (N_11616,N_8372,N_6902);
nor U11617 (N_11617,N_8281,N_6525);
or U11618 (N_11618,N_8832,N_8529);
and U11619 (N_11619,N_7946,N_7842);
and U11620 (N_11620,N_7028,N_8610);
or U11621 (N_11621,N_6810,N_6985);
xnor U11622 (N_11622,N_7913,N_7115);
nor U11623 (N_11623,N_6800,N_8923);
nor U11624 (N_11624,N_7110,N_6929);
or U11625 (N_11625,N_7579,N_6417);
xor U11626 (N_11626,N_6547,N_7436);
nor U11627 (N_11627,N_8236,N_6149);
nor U11628 (N_11628,N_8384,N_8681);
or U11629 (N_11629,N_7961,N_7702);
and U11630 (N_11630,N_6734,N_8607);
or U11631 (N_11631,N_6076,N_7034);
and U11632 (N_11632,N_6183,N_7825);
and U11633 (N_11633,N_8252,N_8041);
and U11634 (N_11634,N_6706,N_6917);
nor U11635 (N_11635,N_6402,N_7281);
nor U11636 (N_11636,N_8089,N_7544);
xnor U11637 (N_11637,N_7590,N_7387);
nand U11638 (N_11638,N_8609,N_6238);
and U11639 (N_11639,N_7277,N_6008);
or U11640 (N_11640,N_6046,N_7729);
xnor U11641 (N_11641,N_8565,N_8008);
or U11642 (N_11642,N_6140,N_6409);
nand U11643 (N_11643,N_6668,N_6303);
and U11644 (N_11644,N_6074,N_8721);
nor U11645 (N_11645,N_7543,N_7691);
nand U11646 (N_11646,N_8851,N_6075);
and U11647 (N_11647,N_8989,N_8393);
xnor U11648 (N_11648,N_6832,N_7487);
xnor U11649 (N_11649,N_8532,N_6958);
nand U11650 (N_11650,N_8467,N_6023);
and U11651 (N_11651,N_7717,N_6067);
xnor U11652 (N_11652,N_7504,N_8053);
xor U11653 (N_11653,N_6699,N_7125);
nor U11654 (N_11654,N_7801,N_7006);
or U11655 (N_11655,N_8353,N_8736);
xnor U11656 (N_11656,N_7304,N_6559);
and U11657 (N_11657,N_7972,N_6817);
nor U11658 (N_11658,N_7357,N_8131);
nand U11659 (N_11659,N_8026,N_6192);
and U11660 (N_11660,N_7536,N_7758);
xnor U11661 (N_11661,N_6495,N_6102);
and U11662 (N_11662,N_8191,N_7416);
and U11663 (N_11663,N_8675,N_6941);
nor U11664 (N_11664,N_8428,N_7795);
nor U11665 (N_11665,N_8275,N_8935);
xnor U11666 (N_11666,N_8097,N_6084);
nand U11667 (N_11667,N_8795,N_7717);
and U11668 (N_11668,N_8723,N_7435);
or U11669 (N_11669,N_6400,N_8126);
nand U11670 (N_11670,N_7978,N_7372);
xor U11671 (N_11671,N_8703,N_7828);
xor U11672 (N_11672,N_7793,N_8002);
xnor U11673 (N_11673,N_6994,N_6842);
nor U11674 (N_11674,N_6559,N_7758);
xnor U11675 (N_11675,N_8418,N_7105);
nor U11676 (N_11676,N_8744,N_6890);
nand U11677 (N_11677,N_6689,N_6942);
xnor U11678 (N_11678,N_6086,N_7183);
or U11679 (N_11679,N_6016,N_6056);
or U11680 (N_11680,N_7992,N_6522);
and U11681 (N_11681,N_6258,N_7892);
xor U11682 (N_11682,N_7810,N_7534);
nand U11683 (N_11683,N_6299,N_8872);
nand U11684 (N_11684,N_8925,N_8970);
nor U11685 (N_11685,N_7950,N_7687);
and U11686 (N_11686,N_7238,N_6218);
xor U11687 (N_11687,N_6229,N_8295);
and U11688 (N_11688,N_7219,N_8444);
nand U11689 (N_11689,N_8557,N_6543);
nand U11690 (N_11690,N_6228,N_8614);
xor U11691 (N_11691,N_7667,N_8595);
or U11692 (N_11692,N_7583,N_8343);
nor U11693 (N_11693,N_6655,N_8100);
nand U11694 (N_11694,N_7201,N_8521);
nand U11695 (N_11695,N_6433,N_8875);
nand U11696 (N_11696,N_7656,N_6793);
and U11697 (N_11697,N_8766,N_6790);
nor U11698 (N_11698,N_8096,N_6338);
and U11699 (N_11699,N_6387,N_7798);
and U11700 (N_11700,N_6969,N_7700);
and U11701 (N_11701,N_7038,N_7128);
nor U11702 (N_11702,N_8397,N_6657);
xnor U11703 (N_11703,N_7136,N_6792);
nand U11704 (N_11704,N_8840,N_8642);
or U11705 (N_11705,N_6288,N_7010);
or U11706 (N_11706,N_6883,N_7658);
xnor U11707 (N_11707,N_7598,N_7882);
xnor U11708 (N_11708,N_7483,N_8939);
nor U11709 (N_11709,N_6415,N_8064);
nor U11710 (N_11710,N_7823,N_6999);
or U11711 (N_11711,N_6787,N_6928);
and U11712 (N_11712,N_7888,N_6796);
or U11713 (N_11713,N_8423,N_6647);
or U11714 (N_11714,N_6591,N_8929);
nand U11715 (N_11715,N_8895,N_8398);
and U11716 (N_11716,N_8965,N_6764);
or U11717 (N_11717,N_6091,N_8029);
and U11718 (N_11718,N_8553,N_6486);
xor U11719 (N_11719,N_6231,N_6826);
nor U11720 (N_11720,N_6645,N_8859);
nor U11721 (N_11721,N_7708,N_8399);
nand U11722 (N_11722,N_6682,N_6106);
xnor U11723 (N_11723,N_8400,N_6319);
nor U11724 (N_11724,N_7732,N_7436);
nand U11725 (N_11725,N_8533,N_7794);
or U11726 (N_11726,N_7424,N_8601);
nand U11727 (N_11727,N_6308,N_8610);
xor U11728 (N_11728,N_8490,N_6043);
and U11729 (N_11729,N_7334,N_7885);
and U11730 (N_11730,N_7646,N_6744);
xnor U11731 (N_11731,N_6252,N_6343);
xor U11732 (N_11732,N_6741,N_7096);
nand U11733 (N_11733,N_7738,N_7908);
and U11734 (N_11734,N_7094,N_6536);
nand U11735 (N_11735,N_6451,N_6406);
and U11736 (N_11736,N_6488,N_7695);
xor U11737 (N_11737,N_7335,N_8619);
and U11738 (N_11738,N_7895,N_8930);
nand U11739 (N_11739,N_8382,N_8864);
and U11740 (N_11740,N_6592,N_6381);
xor U11741 (N_11741,N_8854,N_6463);
xnor U11742 (N_11742,N_7833,N_7150);
and U11743 (N_11743,N_6401,N_7025);
xnor U11744 (N_11744,N_6836,N_8820);
nand U11745 (N_11745,N_7207,N_7012);
nor U11746 (N_11746,N_8511,N_7857);
nor U11747 (N_11747,N_6453,N_6468);
xor U11748 (N_11748,N_8569,N_7757);
or U11749 (N_11749,N_6658,N_7917);
nor U11750 (N_11750,N_6681,N_7684);
xor U11751 (N_11751,N_6829,N_7909);
nand U11752 (N_11752,N_7487,N_6178);
or U11753 (N_11753,N_7115,N_8918);
nand U11754 (N_11754,N_7566,N_7793);
xor U11755 (N_11755,N_7060,N_8363);
xor U11756 (N_11756,N_8629,N_8724);
or U11757 (N_11757,N_7657,N_8170);
nor U11758 (N_11758,N_8719,N_6720);
xnor U11759 (N_11759,N_7914,N_6533);
or U11760 (N_11760,N_7371,N_7083);
nor U11761 (N_11761,N_7805,N_8780);
nor U11762 (N_11762,N_7487,N_8624);
xor U11763 (N_11763,N_7755,N_8960);
and U11764 (N_11764,N_7576,N_6982);
or U11765 (N_11765,N_7226,N_8230);
nand U11766 (N_11766,N_8347,N_8944);
xor U11767 (N_11767,N_8068,N_7963);
and U11768 (N_11768,N_7592,N_6465);
and U11769 (N_11769,N_7546,N_6589);
and U11770 (N_11770,N_8472,N_8990);
nand U11771 (N_11771,N_8921,N_8455);
or U11772 (N_11772,N_7941,N_7960);
nand U11773 (N_11773,N_6293,N_6113);
xnor U11774 (N_11774,N_8832,N_7011);
and U11775 (N_11775,N_7605,N_7065);
and U11776 (N_11776,N_6449,N_8691);
and U11777 (N_11777,N_7224,N_8009);
nand U11778 (N_11778,N_8044,N_6693);
nand U11779 (N_11779,N_6365,N_7755);
and U11780 (N_11780,N_8064,N_8205);
xor U11781 (N_11781,N_6467,N_6048);
nor U11782 (N_11782,N_6303,N_8574);
and U11783 (N_11783,N_7252,N_7655);
and U11784 (N_11784,N_6154,N_8524);
nand U11785 (N_11785,N_7503,N_6122);
and U11786 (N_11786,N_8646,N_7834);
or U11787 (N_11787,N_8753,N_6068);
xor U11788 (N_11788,N_7304,N_8605);
nor U11789 (N_11789,N_6468,N_6625);
and U11790 (N_11790,N_8635,N_7149);
nand U11791 (N_11791,N_8563,N_7293);
xnor U11792 (N_11792,N_8421,N_6147);
or U11793 (N_11793,N_8252,N_7832);
nor U11794 (N_11794,N_6477,N_6705);
nand U11795 (N_11795,N_6346,N_7105);
nor U11796 (N_11796,N_6151,N_7069);
nand U11797 (N_11797,N_7852,N_6388);
or U11798 (N_11798,N_8109,N_8582);
xor U11799 (N_11799,N_6314,N_8280);
nand U11800 (N_11800,N_7568,N_8773);
xor U11801 (N_11801,N_7600,N_7867);
nand U11802 (N_11802,N_7154,N_8877);
or U11803 (N_11803,N_8322,N_7437);
or U11804 (N_11804,N_8546,N_8630);
nor U11805 (N_11805,N_8690,N_6492);
xor U11806 (N_11806,N_6705,N_7398);
xor U11807 (N_11807,N_6294,N_6020);
nor U11808 (N_11808,N_7054,N_6796);
nand U11809 (N_11809,N_8950,N_8633);
xnor U11810 (N_11810,N_7821,N_7394);
nor U11811 (N_11811,N_7545,N_7892);
xnor U11812 (N_11812,N_7945,N_7847);
nor U11813 (N_11813,N_8594,N_6870);
and U11814 (N_11814,N_7899,N_8632);
or U11815 (N_11815,N_7436,N_6942);
or U11816 (N_11816,N_8183,N_6400);
and U11817 (N_11817,N_7587,N_7941);
nor U11818 (N_11818,N_6279,N_6822);
nand U11819 (N_11819,N_7240,N_6189);
and U11820 (N_11820,N_6618,N_8321);
or U11821 (N_11821,N_6950,N_7468);
or U11822 (N_11822,N_7209,N_8734);
nand U11823 (N_11823,N_6733,N_7096);
and U11824 (N_11824,N_6177,N_8551);
xnor U11825 (N_11825,N_6016,N_7132);
nor U11826 (N_11826,N_7633,N_8341);
or U11827 (N_11827,N_8717,N_6970);
nand U11828 (N_11828,N_6600,N_6141);
and U11829 (N_11829,N_6870,N_8354);
nor U11830 (N_11830,N_7971,N_8627);
or U11831 (N_11831,N_6625,N_6451);
nor U11832 (N_11832,N_6487,N_8459);
or U11833 (N_11833,N_8103,N_8634);
nor U11834 (N_11834,N_7195,N_7734);
nor U11835 (N_11835,N_8372,N_8871);
xnor U11836 (N_11836,N_6327,N_8030);
nor U11837 (N_11837,N_8981,N_8130);
nand U11838 (N_11838,N_8517,N_8871);
or U11839 (N_11839,N_8574,N_8190);
nor U11840 (N_11840,N_6197,N_7123);
or U11841 (N_11841,N_7215,N_7415);
or U11842 (N_11842,N_7975,N_6162);
nand U11843 (N_11843,N_7853,N_7306);
xor U11844 (N_11844,N_6698,N_7322);
xor U11845 (N_11845,N_8564,N_6635);
nand U11846 (N_11846,N_7909,N_8920);
nand U11847 (N_11847,N_6624,N_8481);
nand U11848 (N_11848,N_6326,N_8244);
nand U11849 (N_11849,N_7204,N_6051);
and U11850 (N_11850,N_6086,N_6198);
nor U11851 (N_11851,N_8658,N_8097);
nand U11852 (N_11852,N_6070,N_7967);
nor U11853 (N_11853,N_7426,N_8161);
nor U11854 (N_11854,N_8075,N_8514);
or U11855 (N_11855,N_6171,N_7696);
nand U11856 (N_11856,N_7308,N_7335);
xor U11857 (N_11857,N_8517,N_7471);
xnor U11858 (N_11858,N_6865,N_6712);
xor U11859 (N_11859,N_8279,N_7866);
nor U11860 (N_11860,N_6544,N_6384);
and U11861 (N_11861,N_7432,N_7686);
and U11862 (N_11862,N_6686,N_6669);
and U11863 (N_11863,N_8110,N_8179);
xor U11864 (N_11864,N_8423,N_8619);
nor U11865 (N_11865,N_6564,N_8109);
xnor U11866 (N_11866,N_8024,N_6998);
nor U11867 (N_11867,N_8483,N_6732);
xor U11868 (N_11868,N_8799,N_8647);
and U11869 (N_11869,N_7683,N_7750);
and U11870 (N_11870,N_6711,N_7831);
or U11871 (N_11871,N_8593,N_7520);
and U11872 (N_11872,N_7521,N_8738);
nor U11873 (N_11873,N_7795,N_8091);
nand U11874 (N_11874,N_7224,N_7097);
nor U11875 (N_11875,N_7665,N_7314);
and U11876 (N_11876,N_8044,N_8015);
nand U11877 (N_11877,N_8191,N_6696);
nor U11878 (N_11878,N_7916,N_6895);
nand U11879 (N_11879,N_8509,N_6616);
and U11880 (N_11880,N_7477,N_8887);
nor U11881 (N_11881,N_6094,N_7256);
nand U11882 (N_11882,N_7652,N_7966);
and U11883 (N_11883,N_8106,N_6970);
xor U11884 (N_11884,N_7402,N_8582);
nand U11885 (N_11885,N_7712,N_8114);
or U11886 (N_11886,N_6742,N_8930);
xor U11887 (N_11887,N_6765,N_8321);
xor U11888 (N_11888,N_6235,N_6399);
and U11889 (N_11889,N_7464,N_7365);
nor U11890 (N_11890,N_7001,N_7448);
or U11891 (N_11891,N_8832,N_8967);
nand U11892 (N_11892,N_6982,N_8301);
and U11893 (N_11893,N_7383,N_6857);
xor U11894 (N_11894,N_6949,N_8159);
nor U11895 (N_11895,N_7066,N_7810);
and U11896 (N_11896,N_8870,N_6068);
or U11897 (N_11897,N_8985,N_7779);
or U11898 (N_11898,N_7928,N_6716);
nand U11899 (N_11899,N_7131,N_6532);
xnor U11900 (N_11900,N_7157,N_8046);
or U11901 (N_11901,N_6101,N_8598);
xnor U11902 (N_11902,N_6574,N_8204);
nor U11903 (N_11903,N_8986,N_8114);
and U11904 (N_11904,N_7693,N_7926);
and U11905 (N_11905,N_7295,N_6339);
nor U11906 (N_11906,N_6969,N_7376);
and U11907 (N_11907,N_8239,N_7698);
nor U11908 (N_11908,N_7231,N_8518);
nand U11909 (N_11909,N_8249,N_8367);
nor U11910 (N_11910,N_8909,N_6337);
and U11911 (N_11911,N_7245,N_8317);
and U11912 (N_11912,N_6341,N_7289);
and U11913 (N_11913,N_7340,N_6360);
xnor U11914 (N_11914,N_6792,N_6659);
and U11915 (N_11915,N_7781,N_6614);
nor U11916 (N_11916,N_7730,N_6640);
and U11917 (N_11917,N_7360,N_6481);
and U11918 (N_11918,N_6774,N_8457);
and U11919 (N_11919,N_7441,N_6840);
nor U11920 (N_11920,N_6861,N_8139);
nand U11921 (N_11921,N_6844,N_8552);
or U11922 (N_11922,N_8266,N_6390);
nor U11923 (N_11923,N_8425,N_6907);
and U11924 (N_11924,N_6800,N_7229);
and U11925 (N_11925,N_6529,N_8162);
xor U11926 (N_11926,N_8377,N_8206);
xor U11927 (N_11927,N_7402,N_7924);
or U11928 (N_11928,N_6374,N_7430);
and U11929 (N_11929,N_7364,N_8045);
xnor U11930 (N_11930,N_8197,N_8136);
xor U11931 (N_11931,N_8183,N_8980);
and U11932 (N_11932,N_7368,N_8282);
nand U11933 (N_11933,N_6038,N_6448);
or U11934 (N_11934,N_6787,N_7227);
nor U11935 (N_11935,N_7343,N_6789);
or U11936 (N_11936,N_8781,N_7561);
or U11937 (N_11937,N_6634,N_8489);
or U11938 (N_11938,N_7803,N_6068);
and U11939 (N_11939,N_6475,N_6576);
nor U11940 (N_11940,N_6862,N_8515);
xnor U11941 (N_11941,N_8862,N_6253);
nand U11942 (N_11942,N_7916,N_6893);
and U11943 (N_11943,N_6650,N_8775);
xor U11944 (N_11944,N_6809,N_7025);
nand U11945 (N_11945,N_8138,N_7494);
nand U11946 (N_11946,N_7824,N_7697);
nand U11947 (N_11947,N_7014,N_8823);
nor U11948 (N_11948,N_6823,N_6335);
nand U11949 (N_11949,N_7505,N_6445);
or U11950 (N_11950,N_6426,N_7013);
nor U11951 (N_11951,N_7560,N_8962);
and U11952 (N_11952,N_7554,N_7149);
and U11953 (N_11953,N_8365,N_7834);
nand U11954 (N_11954,N_8743,N_8599);
or U11955 (N_11955,N_8141,N_6000);
or U11956 (N_11956,N_6458,N_8588);
or U11957 (N_11957,N_6204,N_6758);
nor U11958 (N_11958,N_6169,N_6367);
nand U11959 (N_11959,N_6099,N_6869);
nor U11960 (N_11960,N_7635,N_6016);
and U11961 (N_11961,N_7691,N_7139);
and U11962 (N_11962,N_7420,N_7852);
and U11963 (N_11963,N_6748,N_7406);
and U11964 (N_11964,N_7986,N_8097);
or U11965 (N_11965,N_6673,N_6170);
xor U11966 (N_11966,N_8442,N_8464);
and U11967 (N_11967,N_7545,N_6119);
nand U11968 (N_11968,N_7731,N_7798);
nand U11969 (N_11969,N_6709,N_8305);
xor U11970 (N_11970,N_7306,N_6812);
nand U11971 (N_11971,N_6338,N_6737);
and U11972 (N_11972,N_7316,N_6178);
nand U11973 (N_11973,N_7456,N_6389);
nand U11974 (N_11974,N_6100,N_7656);
nor U11975 (N_11975,N_7889,N_6712);
nand U11976 (N_11976,N_8794,N_8277);
xnor U11977 (N_11977,N_6261,N_7911);
nor U11978 (N_11978,N_7868,N_7125);
or U11979 (N_11979,N_6909,N_7177);
xnor U11980 (N_11980,N_7691,N_7820);
nand U11981 (N_11981,N_7307,N_6931);
or U11982 (N_11982,N_7337,N_6222);
or U11983 (N_11983,N_8506,N_8670);
xnor U11984 (N_11984,N_7745,N_7793);
or U11985 (N_11985,N_7592,N_6912);
nor U11986 (N_11986,N_6897,N_7326);
and U11987 (N_11987,N_8153,N_8628);
xor U11988 (N_11988,N_6256,N_8219);
or U11989 (N_11989,N_6682,N_6003);
nor U11990 (N_11990,N_6389,N_6995);
and U11991 (N_11991,N_7305,N_8308);
xor U11992 (N_11992,N_8665,N_8347);
nand U11993 (N_11993,N_7556,N_8727);
xor U11994 (N_11994,N_7824,N_7918);
xor U11995 (N_11995,N_8123,N_6883);
or U11996 (N_11996,N_8650,N_6251);
xor U11997 (N_11997,N_7599,N_8497);
nor U11998 (N_11998,N_7330,N_8221);
or U11999 (N_11999,N_6024,N_7434);
and U12000 (N_12000,N_10070,N_11186);
and U12001 (N_12001,N_10714,N_11076);
nor U12002 (N_12002,N_10901,N_10110);
nand U12003 (N_12003,N_9100,N_9622);
and U12004 (N_12004,N_9244,N_10596);
nand U12005 (N_12005,N_9549,N_10026);
xor U12006 (N_12006,N_11302,N_9394);
or U12007 (N_12007,N_9322,N_10570);
nor U12008 (N_12008,N_11546,N_10174);
and U12009 (N_12009,N_11697,N_9783);
nand U12010 (N_12010,N_10024,N_10525);
nand U12011 (N_12011,N_9345,N_11424);
nand U12012 (N_12012,N_11814,N_9854);
and U12013 (N_12013,N_10131,N_9996);
and U12014 (N_12014,N_9206,N_9369);
xnor U12015 (N_12015,N_11143,N_11763);
xor U12016 (N_12016,N_10078,N_10912);
and U12017 (N_12017,N_10454,N_11403);
xnor U12018 (N_12018,N_11364,N_9684);
nor U12019 (N_12019,N_9978,N_11477);
or U12020 (N_12020,N_10624,N_10499);
nor U12021 (N_12021,N_9513,N_9564);
nor U12022 (N_12022,N_11241,N_10075);
and U12023 (N_12023,N_11167,N_11960);
and U12024 (N_12024,N_9742,N_11385);
xnor U12025 (N_12025,N_10950,N_9005);
and U12026 (N_12026,N_10697,N_11058);
and U12027 (N_12027,N_9055,N_9190);
xnor U12028 (N_12028,N_9747,N_9392);
and U12029 (N_12029,N_9951,N_9601);
nand U12030 (N_12030,N_11715,N_11958);
and U12031 (N_12031,N_10173,N_11844);
nand U12032 (N_12032,N_10356,N_9624);
and U12033 (N_12033,N_11103,N_10620);
nor U12034 (N_12034,N_9305,N_10528);
nor U12035 (N_12035,N_9258,N_9480);
nand U12036 (N_12036,N_9659,N_11609);
or U12037 (N_12037,N_9265,N_9059);
xnor U12038 (N_12038,N_9066,N_10358);
nor U12039 (N_12039,N_9098,N_10723);
and U12040 (N_12040,N_10130,N_11415);
and U12041 (N_12041,N_9867,N_10015);
nand U12042 (N_12042,N_9671,N_11141);
and U12043 (N_12043,N_10524,N_11412);
or U12044 (N_12044,N_11976,N_11535);
nor U12045 (N_12045,N_11436,N_11102);
and U12046 (N_12046,N_9507,N_10664);
nand U12047 (N_12047,N_10868,N_11825);
xor U12048 (N_12048,N_9896,N_11848);
and U12049 (N_12049,N_9567,N_11421);
xnor U12050 (N_12050,N_9444,N_9638);
nor U12051 (N_12051,N_11975,N_11252);
or U12052 (N_12052,N_11195,N_11517);
nand U12053 (N_12053,N_11114,N_11692);
nand U12054 (N_12054,N_10818,N_10933);
nand U12055 (N_12055,N_11258,N_11482);
xor U12056 (N_12056,N_9554,N_9824);
and U12057 (N_12057,N_9210,N_9414);
or U12058 (N_12058,N_11784,N_11070);
and U12059 (N_12059,N_10772,N_11527);
or U12060 (N_12060,N_11084,N_10698);
and U12061 (N_12061,N_11718,N_9705);
and U12062 (N_12062,N_11497,N_10306);
and U12063 (N_12063,N_10521,N_11378);
nor U12064 (N_12064,N_9974,N_11232);
nand U12065 (N_12065,N_10971,N_9503);
or U12066 (N_12066,N_9016,N_11269);
nand U12067 (N_12067,N_10298,N_11164);
and U12068 (N_12068,N_10021,N_10321);
xnor U12069 (N_12069,N_10422,N_11351);
nand U12070 (N_12070,N_9211,N_9436);
xnor U12071 (N_12071,N_10065,N_10179);
xnor U12072 (N_12072,N_9730,N_10833);
and U12073 (N_12073,N_11465,N_10048);
xor U12074 (N_12074,N_11935,N_10458);
nor U12075 (N_12075,N_9559,N_11719);
xor U12076 (N_12076,N_10142,N_9221);
and U12077 (N_12077,N_11920,N_11035);
nor U12078 (N_12078,N_11365,N_9683);
and U12079 (N_12079,N_9933,N_9483);
nand U12080 (N_12080,N_11346,N_10307);
xor U12081 (N_12081,N_9844,N_10042);
xnor U12082 (N_12082,N_10480,N_11766);
or U12083 (N_12083,N_10583,N_11100);
nor U12084 (N_12084,N_10311,N_10397);
or U12085 (N_12085,N_9645,N_11292);
nand U12086 (N_12086,N_11328,N_10449);
nor U12087 (N_12087,N_10137,N_9508);
and U12088 (N_12088,N_11854,N_9868);
or U12089 (N_12089,N_10953,N_11587);
and U12090 (N_12090,N_11612,N_11870);
nor U12091 (N_12091,N_10739,N_10826);
xor U12092 (N_12092,N_9878,N_10039);
or U12093 (N_12093,N_11708,N_10495);
nor U12094 (N_12094,N_11998,N_11681);
nand U12095 (N_12095,N_10462,N_9900);
nor U12096 (N_12096,N_10045,N_9644);
xnor U12097 (N_12097,N_10588,N_9290);
and U12098 (N_12098,N_9164,N_11341);
nor U12099 (N_12099,N_10262,N_11754);
nand U12100 (N_12100,N_9312,N_9876);
nand U12101 (N_12101,N_10803,N_11600);
xor U12102 (N_12102,N_9101,N_9024);
xor U12103 (N_12103,N_9422,N_10692);
nor U12104 (N_12104,N_10657,N_9534);
and U12105 (N_12105,N_11877,N_11116);
nand U12106 (N_12106,N_10861,N_9156);
nand U12107 (N_12107,N_10081,N_9278);
xnor U12108 (N_12108,N_9769,N_11373);
nor U12109 (N_12109,N_9993,N_11282);
or U12110 (N_12110,N_10423,N_9701);
nand U12111 (N_12111,N_11501,N_9517);
and U12112 (N_12112,N_9755,N_11537);
xnor U12113 (N_12113,N_9126,N_9643);
xor U12114 (N_12114,N_9434,N_11912);
and U12115 (N_12115,N_10545,N_10910);
xor U12116 (N_12116,N_11499,N_11264);
and U12117 (N_12117,N_11205,N_9053);
or U12118 (N_12118,N_10202,N_9048);
or U12119 (N_12119,N_11223,N_10341);
nand U12120 (N_12120,N_9072,N_10194);
xnor U12121 (N_12121,N_11545,N_11340);
xor U12122 (N_12122,N_11027,N_11469);
nor U12123 (N_12123,N_9427,N_10176);
nand U12124 (N_12124,N_11307,N_11334);
nor U12125 (N_12125,N_11916,N_9541);
nor U12126 (N_12126,N_10169,N_10560);
or U12127 (N_12127,N_11795,N_11984);
nand U12128 (N_12128,N_9540,N_9964);
nor U12129 (N_12129,N_11742,N_11688);
xnor U12130 (N_12130,N_9197,N_9649);
nand U12131 (N_12131,N_11067,N_9668);
nand U12132 (N_12132,N_10970,N_9631);
xor U12133 (N_12133,N_9799,N_9665);
nor U12134 (N_12134,N_9527,N_10085);
xor U12135 (N_12135,N_9907,N_9883);
xor U12136 (N_12136,N_11714,N_10217);
nand U12137 (N_12137,N_10364,N_9308);
xor U12138 (N_12138,N_10814,N_11862);
and U12139 (N_12139,N_10730,N_9111);
nor U12140 (N_12140,N_11438,N_10291);
nand U12141 (N_12141,N_9025,N_9501);
and U12142 (N_12142,N_10726,N_11224);
and U12143 (N_12143,N_10822,N_9360);
or U12144 (N_12144,N_11213,N_9310);
and U12145 (N_12145,N_9218,N_10218);
nand U12146 (N_12146,N_10631,N_9944);
or U12147 (N_12147,N_9573,N_10537);
or U12148 (N_12148,N_11696,N_10770);
nand U12149 (N_12149,N_11214,N_9034);
or U12150 (N_12150,N_10133,N_9814);
nand U12151 (N_12151,N_10103,N_10675);
xnor U12152 (N_12152,N_11310,N_10198);
xnor U12153 (N_12153,N_11138,N_11734);
nor U12154 (N_12154,N_9620,N_11466);
nand U12155 (N_12155,N_9617,N_9056);
nor U12156 (N_12156,N_9796,N_11071);
and U12157 (N_12157,N_10378,N_9355);
and U12158 (N_12158,N_11124,N_10945);
xnor U12159 (N_12159,N_9982,N_10703);
xnor U12160 (N_12160,N_10641,N_11749);
nor U12161 (N_12161,N_11175,N_9932);
nand U12162 (N_12162,N_9677,N_11721);
or U12163 (N_12163,N_10416,N_11893);
and U12164 (N_12164,N_11416,N_10759);
or U12165 (N_12165,N_9589,N_10434);
and U12166 (N_12166,N_11352,N_11126);
nor U12167 (N_12167,N_9338,N_10143);
or U12168 (N_12168,N_11133,N_10731);
and U12169 (N_12169,N_10183,N_9882);
and U12170 (N_12170,N_11772,N_10411);
xor U12171 (N_12171,N_11685,N_9811);
nor U12172 (N_12172,N_10410,N_10832);
nor U12173 (N_12173,N_10186,N_10589);
and U12174 (N_12174,N_11171,N_11871);
nor U12175 (N_12175,N_10063,N_10448);
nand U12176 (N_12176,N_11115,N_11608);
xnor U12177 (N_12177,N_9260,N_11149);
xnor U12178 (N_12178,N_10461,N_9162);
or U12179 (N_12179,N_10542,N_11561);
xor U12180 (N_12180,N_9803,N_9832);
and U12181 (N_12181,N_10993,N_9008);
or U12182 (N_12182,N_10083,N_9716);
nand U12183 (N_12183,N_10853,N_11360);
and U12184 (N_12184,N_10430,N_11025);
and U12185 (N_12185,N_10598,N_10577);
and U12186 (N_12186,N_11383,N_10195);
nor U12187 (N_12187,N_10090,N_11247);
nor U12188 (N_12188,N_9858,N_10764);
nor U12189 (N_12189,N_9981,N_11142);
and U12190 (N_12190,N_11644,N_11228);
xor U12191 (N_12191,N_10964,N_10827);
nor U12192 (N_12192,N_11250,N_10118);
or U12193 (N_12193,N_11859,N_11940);
or U12194 (N_12194,N_11240,N_9909);
xnor U12195 (N_12195,N_10909,N_9830);
or U12196 (N_12196,N_9767,N_10967);
nand U12197 (N_12197,N_9550,N_10302);
and U12198 (N_12198,N_10960,N_10767);
nor U12199 (N_12199,N_9324,N_11538);
nand U12200 (N_12200,N_10666,N_10595);
or U12201 (N_12201,N_11081,N_9724);
and U12202 (N_12202,N_9577,N_11691);
or U12203 (N_12203,N_11362,N_11625);
or U12204 (N_12204,N_11462,N_11583);
and U12205 (N_12205,N_9081,N_9575);
xor U12206 (N_12206,N_9425,N_11369);
nor U12207 (N_12207,N_9592,N_10211);
or U12208 (N_12208,N_9328,N_11621);
and U12209 (N_12209,N_10443,N_10421);
and U12210 (N_12210,N_10694,N_11646);
or U12211 (N_12211,N_9842,N_10288);
xnor U12212 (N_12212,N_10023,N_11379);
nand U12213 (N_12213,N_9354,N_10144);
xor U12214 (N_12214,N_11557,N_11181);
nor U12215 (N_12215,N_9363,N_10928);
and U12216 (N_12216,N_11518,N_11648);
nand U12217 (N_12217,N_10471,N_10673);
xor U12218 (N_12218,N_11390,N_9366);
or U12219 (N_12219,N_10308,N_9253);
nand U12220 (N_12220,N_11633,N_10988);
nor U12221 (N_12221,N_10609,N_9795);
nand U12222 (N_12222,N_11919,N_11093);
or U12223 (N_12223,N_10225,N_10985);
xnor U12224 (N_12224,N_10141,N_10957);
and U12225 (N_12225,N_10856,N_10293);
and U12226 (N_12226,N_9569,N_9772);
nor U12227 (N_12227,N_9424,N_9154);
and U12228 (N_12228,N_10648,N_9296);
nor U12229 (N_12229,N_10013,N_9042);
or U12230 (N_12230,N_9222,N_11426);
or U12231 (N_12231,N_11040,N_10236);
xnor U12232 (N_12232,N_11942,N_10066);
nand U12233 (N_12233,N_10256,N_10937);
nand U12234 (N_12234,N_10071,N_10088);
or U12235 (N_12235,N_11288,N_11530);
or U12236 (N_12236,N_11690,N_11377);
xor U12237 (N_12237,N_9556,N_10830);
xnor U12238 (N_12238,N_10955,N_10239);
nor U12239 (N_12239,N_10270,N_9160);
nor U12240 (N_12240,N_9561,N_11253);
and U12241 (N_12241,N_9188,N_9050);
and U12242 (N_12242,N_10167,N_10485);
nor U12243 (N_12243,N_11885,N_9365);
and U12244 (N_12244,N_10760,N_10328);
xor U12245 (N_12245,N_10136,N_10392);
nor U12246 (N_12246,N_10687,N_10628);
xnor U12247 (N_12247,N_9039,N_9405);
or U12248 (N_12248,N_9725,N_10644);
or U12249 (N_12249,N_11061,N_10880);
xnor U12250 (N_12250,N_9330,N_11617);
or U12251 (N_12251,N_9471,N_11078);
nor U12252 (N_12252,N_11913,N_11227);
or U12253 (N_12253,N_10189,N_11259);
or U12254 (N_12254,N_11925,N_9407);
and U12255 (N_12255,N_9793,N_11125);
nand U12256 (N_12256,N_11575,N_9606);
and U12257 (N_12257,N_11911,N_9686);
xnor U12258 (N_12258,N_10372,N_10774);
or U12259 (N_12259,N_9863,N_10089);
and U12260 (N_12260,N_11505,N_9737);
nor U12261 (N_12261,N_10080,N_9040);
nor U12262 (N_12262,N_11393,N_11872);
and U12263 (N_12263,N_9536,N_9410);
xor U12264 (N_12264,N_11931,N_11120);
nor U12265 (N_12265,N_11597,N_11155);
or U12266 (N_12266,N_11525,N_10248);
xnor U12267 (N_12267,N_9490,N_10701);
xor U12268 (N_12268,N_9605,N_11978);
and U12269 (N_12269,N_11679,N_10974);
nor U12270 (N_12270,N_9255,N_9022);
nor U12271 (N_12271,N_10860,N_10296);
and U12272 (N_12272,N_10247,N_10643);
and U12273 (N_12273,N_11325,N_11090);
and U12274 (N_12274,N_11347,N_9217);
nand U12275 (N_12275,N_11513,N_11866);
nand U12276 (N_12276,N_10191,N_10517);
nand U12277 (N_12277,N_11305,N_11219);
xnor U12278 (N_12278,N_11986,N_10403);
nor U12279 (N_12279,N_10655,N_10310);
xnor U12280 (N_12280,N_10158,N_10851);
and U12281 (N_12281,N_10446,N_11079);
xnor U12282 (N_12282,N_10459,N_9297);
nand U12283 (N_12283,N_9073,N_10990);
nor U12284 (N_12284,N_9179,N_10742);
or U12285 (N_12285,N_10309,N_10736);
nand U12286 (N_12286,N_11666,N_9857);
nand U12287 (N_12287,N_11011,N_9037);
nor U12288 (N_12288,N_9834,N_9949);
nand U12289 (N_12289,N_9697,N_9486);
and U12290 (N_12290,N_9903,N_10559);
or U12291 (N_12291,N_11407,N_10228);
nand U12292 (N_12292,N_9504,N_9367);
nor U12293 (N_12293,N_9240,N_11570);
nor U12294 (N_12294,N_10414,N_9060);
or U12295 (N_12295,N_10523,N_10235);
nor U12296 (N_12296,N_10798,N_10650);
or U12297 (N_12297,N_11522,N_11112);
or U12298 (N_12298,N_11961,N_9359);
nand U12299 (N_12299,N_11726,N_9770);
nand U12300 (N_12300,N_11442,N_9927);
and U12301 (N_12301,N_9177,N_10242);
and U12302 (N_12302,N_11689,N_10575);
and U12303 (N_12303,N_9199,N_9380);
nand U12304 (N_12304,N_11674,N_11451);
nand U12305 (N_12305,N_10243,N_10223);
nand U12306 (N_12306,N_11770,N_9242);
nand U12307 (N_12307,N_11943,N_10546);
and U12308 (N_12308,N_10640,N_10882);
or U12309 (N_12309,N_9890,N_11890);
and U12310 (N_12310,N_11713,N_10787);
nor U12311 (N_12311,N_10301,N_10263);
nor U12312 (N_12312,N_9674,N_11900);
xnor U12313 (N_12313,N_9560,N_10145);
or U12314 (N_12314,N_9509,N_9362);
or U12315 (N_12315,N_11370,N_10484);
and U12316 (N_12316,N_9170,N_10418);
and U12317 (N_12317,N_10255,N_9849);
xor U12318 (N_12318,N_10233,N_10785);
or U12319 (N_12319,N_10053,N_10608);
xor U12320 (N_12320,N_9489,N_11454);
nand U12321 (N_12321,N_10407,N_10058);
and U12322 (N_12322,N_10452,N_11565);
xnor U12323 (N_12323,N_11645,N_11993);
or U12324 (N_12324,N_11662,N_10313);
or U12325 (N_12325,N_9994,N_9453);
xnor U12326 (N_12326,N_9827,N_11658);
and U12327 (N_12327,N_10312,N_11192);
nor U12328 (N_12328,N_9914,N_10958);
xnor U12329 (N_12329,N_9514,N_11934);
xor U12330 (N_12330,N_9061,N_10722);
and U12331 (N_12331,N_9930,N_10371);
nor U12332 (N_12332,N_11521,N_11456);
xor U12333 (N_12333,N_9463,N_9722);
nand U12334 (N_12334,N_9381,N_9484);
nand U12335 (N_12335,N_10333,N_9011);
nand U12336 (N_12336,N_10894,N_11483);
nand U12337 (N_12337,N_10269,N_11170);
or U12338 (N_12338,N_10922,N_10016);
xor U12339 (N_12339,N_10476,N_9572);
xor U12340 (N_12340,N_10916,N_10483);
nor U12341 (N_12341,N_9368,N_11262);
or U12342 (N_12342,N_9754,N_10508);
nand U12343 (N_12343,N_9374,N_9460);
or U12344 (N_12344,N_10797,N_10445);
or U12345 (N_12345,N_11845,N_10734);
nor U12346 (N_12346,N_10899,N_10547);
or U12347 (N_12347,N_9891,N_10938);
nand U12348 (N_12348,N_9348,N_9880);
or U12349 (N_12349,N_9421,N_10699);
or U12350 (N_12350,N_10511,N_11254);
nor U12351 (N_12351,N_11296,N_11243);
nor U12352 (N_12352,N_11684,N_11459);
nand U12353 (N_12353,N_11199,N_9472);
and U12354 (N_12354,N_9917,N_11601);
or U12355 (N_12355,N_10890,N_10586);
nor U12356 (N_12356,N_10616,N_11190);
and U12357 (N_12357,N_11837,N_9710);
xor U12358 (N_12358,N_11122,N_11344);
or U12359 (N_12359,N_10331,N_11847);
and U12360 (N_12360,N_11965,N_9478);
and U12361 (N_12361,N_9702,N_11405);
xnor U12362 (N_12362,N_10467,N_11406);
nand U12363 (N_12363,N_10388,N_10297);
or U12364 (N_12364,N_10763,N_10206);
nor U12365 (N_12365,N_11515,N_11467);
xnor U12366 (N_12366,N_11826,N_9398);
xor U12367 (N_12367,N_10592,N_10164);
xnor U12368 (N_12368,N_10468,N_10134);
nor U12369 (N_12369,N_11794,N_10304);
or U12370 (N_12370,N_10553,N_9545);
nand U12371 (N_12371,N_11797,N_11812);
or U12372 (N_12372,N_9189,N_11717);
xnor U12373 (N_12373,N_9113,N_10062);
and U12374 (N_12374,N_10219,N_10896);
xor U12375 (N_12375,N_11703,N_11151);
nor U12376 (N_12376,N_9646,N_9828);
nand U12377 (N_12377,N_10744,N_10649);
nand U12378 (N_12378,N_10847,N_11273);
or U12379 (N_12379,N_10897,N_10925);
nor U12380 (N_12380,N_10056,N_11147);
or U12381 (N_12381,N_9157,N_10120);
xor U12382 (N_12382,N_11823,N_9377);
or U12383 (N_12383,N_9329,N_9279);
nand U12384 (N_12384,N_11777,N_9955);
or U12385 (N_12385,N_9127,N_9339);
xor U12386 (N_12386,N_11672,N_9528);
nor U12387 (N_12387,N_10823,N_9630);
nor U12388 (N_12388,N_10662,N_11676);
nor U12389 (N_12389,N_10983,N_11723);
xnor U12390 (N_12390,N_10824,N_10781);
nand U12391 (N_12391,N_11957,N_9216);
and U12392 (N_12392,N_10613,N_9069);
nand U12393 (N_12393,N_10166,N_10018);
nand U12394 (N_12394,N_10050,N_9798);
nor U12395 (N_12395,N_11979,N_9611);
and U12396 (N_12396,N_11833,N_11381);
nor U12397 (N_12397,N_10230,N_10610);
nor U12398 (N_12398,N_10582,N_10815);
or U12399 (N_12399,N_11470,N_9739);
xor U12400 (N_12400,N_10124,N_10921);
xnor U12401 (N_12401,N_9736,N_9812);
and U12402 (N_12402,N_9479,N_10852);
or U12403 (N_12403,N_11211,N_10557);
xor U12404 (N_12404,N_9007,N_10320);
and U12405 (N_12405,N_10754,N_11182);
nor U12406 (N_12406,N_10385,N_10659);
or U12407 (N_12407,N_9787,N_11108);
nand U12408 (N_12408,N_10779,N_10954);
xnor U12409 (N_12409,N_10246,N_11301);
xor U12410 (N_12410,N_9859,N_11386);
and U12411 (N_12411,N_9985,N_10874);
nand U12412 (N_12412,N_10634,N_11059);
or U12413 (N_12413,N_11235,N_10902);
xnor U12414 (N_12414,N_11775,N_10911);
nand U12415 (N_12415,N_9496,N_10425);
nand U12416 (N_12416,N_9726,N_11060);
nand U12417 (N_12417,N_9967,N_9017);
nand U12418 (N_12418,N_10600,N_9445);
or U12419 (N_12419,N_9920,N_10354);
xor U12420 (N_12420,N_11710,N_10929);
nor U12421 (N_12421,N_11539,N_10966);
and U12422 (N_12422,N_9992,N_10819);
or U12423 (N_12423,N_9838,N_9597);
or U12424 (N_12424,N_11808,N_9252);
or U12425 (N_12425,N_11568,N_9547);
or U12426 (N_12426,N_10335,N_11339);
or U12427 (N_12427,N_9987,N_10382);
nand U12428 (N_12428,N_10636,N_9235);
and U12429 (N_12429,N_10404,N_9581);
xnor U12430 (N_12430,N_9320,N_10749);
and U12431 (N_12431,N_11113,N_11229);
xnor U12432 (N_12432,N_9228,N_11431);
nand U12433 (N_12433,N_9303,N_11453);
and U12434 (N_12434,N_10168,N_11397);
nand U12435 (N_12435,N_9306,N_9696);
and U12436 (N_12436,N_11769,N_10432);
nor U12437 (N_12437,N_11811,N_10941);
nor U12438 (N_12438,N_10156,N_10813);
and U12439 (N_12439,N_10107,N_9729);
or U12440 (N_12440,N_9451,N_11032);
or U12441 (N_12441,N_9706,N_10069);
nand U12442 (N_12442,N_11484,N_10405);
xor U12443 (N_12443,N_10030,N_9533);
or U12444 (N_12444,N_9984,N_10479);
and U12445 (N_12445,N_11485,N_9058);
or U12446 (N_12446,N_10345,N_9695);
nor U12447 (N_12447,N_9144,N_9588);
nand U12448 (N_12448,N_10936,N_10806);
xor U12449 (N_12449,N_11145,N_10326);
or U12450 (N_12450,N_11333,N_9450);
or U12451 (N_12451,N_11008,N_9571);
nor U12452 (N_12452,N_11051,N_10951);
nand U12453 (N_12453,N_10778,N_10535);
nor U12454 (N_12454,N_10682,N_10807);
nand U12455 (N_12455,N_10002,N_9474);
nor U12456 (N_12456,N_10623,N_11510);
nand U12457 (N_12457,N_9307,N_11999);
nand U12458 (N_12458,N_10098,N_11498);
xnor U12459 (N_12459,N_11836,N_11524);
or U12460 (N_12460,N_11156,N_9960);
xnor U12461 (N_12461,N_9986,N_9112);
or U12462 (N_12462,N_10172,N_11665);
or U12463 (N_12463,N_9777,N_10652);
and U12464 (N_12464,N_9723,N_11265);
nand U12465 (N_12465,N_11185,N_10935);
or U12466 (N_12466,N_10100,N_9775);
nor U12467 (N_12467,N_9064,N_9411);
or U12468 (N_12468,N_10677,N_9012);
or U12469 (N_12469,N_11969,N_10337);
nand U12470 (N_12470,N_10292,N_9602);
nor U12471 (N_12471,N_11380,N_11129);
and U12472 (N_12472,N_10717,N_9647);
xor U12473 (N_12473,N_9028,N_10907);
or U12474 (N_12474,N_10727,N_11136);
xor U12475 (N_12475,N_9897,N_10791);
xor U12476 (N_12476,N_11630,N_11007);
and U12477 (N_12477,N_10121,N_10630);
and U12478 (N_12478,N_9515,N_11727);
nor U12479 (N_12479,N_11968,N_9402);
nand U12480 (N_12480,N_10845,N_10339);
and U12481 (N_12481,N_11152,N_11495);
nor U12482 (N_12482,N_9873,N_9922);
or U12483 (N_12483,N_11637,N_9790);
or U12484 (N_12484,N_10109,N_9125);
nand U12485 (N_12485,N_10695,N_9087);
nand U12486 (N_12486,N_10688,N_10681);
xnor U12487 (N_12487,N_9839,N_11936);
xnor U12488 (N_12488,N_11852,N_9316);
xor U12489 (N_12489,N_9275,N_9760);
nor U12490 (N_12490,N_11983,N_10040);
xnor U12491 (N_12491,N_9247,N_9397);
nand U12492 (N_12492,N_9613,N_9670);
and U12493 (N_12493,N_9151,N_11560);
nand U12494 (N_12494,N_11460,N_10715);
nor U12495 (N_12495,N_10054,N_9114);
nor U12496 (N_12496,N_9709,N_11874);
xnor U12497 (N_12497,N_11016,N_10883);
and U12498 (N_12498,N_9107,N_11955);
nor U12499 (N_12499,N_11661,N_11663);
nor U12500 (N_12500,N_11440,N_10221);
nor U12501 (N_12501,N_11441,N_11980);
or U12502 (N_12502,N_9353,N_9884);
xor U12503 (N_12503,N_11620,N_11356);
and U12504 (N_12504,N_11554,N_11730);
or U12505 (N_12505,N_11653,N_11589);
nand U12506 (N_12506,N_11791,N_10908);
and U12507 (N_12507,N_9442,N_11239);
or U12508 (N_12508,N_11111,N_11768);
nand U12509 (N_12509,N_10436,N_9744);
xnor U12510 (N_12510,N_11366,N_9989);
nand U12511 (N_12511,N_9429,N_11263);
or U12512 (N_12512,N_11799,N_11720);
and U12513 (N_12513,N_11953,N_9289);
and U12514 (N_12514,N_11846,N_9990);
xor U12515 (N_12515,N_11187,N_11753);
xnor U12516 (N_12516,N_9959,N_11843);
and U12517 (N_12517,N_9166,N_11057);
and U12518 (N_12518,N_10618,N_10603);
or U12519 (N_12519,N_10705,N_10325);
and U12520 (N_12520,N_9800,N_10357);
or U12521 (N_12521,N_10319,N_9473);
nand U12522 (N_12522,N_10314,N_9500);
nor U12523 (N_12523,N_10888,N_10658);
nand U12524 (N_12524,N_10707,N_10572);
nand U12525 (N_12525,N_9929,N_10258);
and U12526 (N_12526,N_10552,N_11776);
nor U12527 (N_12527,N_11033,N_10286);
or U12528 (N_12528,N_11917,N_11809);
nor U12529 (N_12529,N_10565,N_9001);
and U12530 (N_12530,N_11207,N_10998);
nand U12531 (N_12531,N_10049,N_11086);
and U12532 (N_12532,N_11831,N_11873);
xnor U12533 (N_12533,N_10984,N_11197);
xor U12534 (N_12534,N_11266,N_9753);
nor U12535 (N_12535,N_9682,N_10713);
xnor U12536 (N_12536,N_9825,N_10601);
or U12537 (N_12537,N_9277,N_11650);
nand U12538 (N_12538,N_9950,N_11821);
and U12539 (N_12539,N_10633,N_10917);
and U12540 (N_12540,N_11687,N_10579);
or U12541 (N_12541,N_11367,N_9132);
and U12542 (N_12542,N_9945,N_11316);
nand U12543 (N_12543,N_11411,N_11906);
or U12544 (N_12544,N_11030,N_10303);
xnor U12545 (N_12545,N_9761,N_9083);
nand U12546 (N_12546,N_10660,N_10464);
and U12547 (N_12547,N_9401,N_10540);
and U12548 (N_12548,N_11329,N_10663);
and U12549 (N_12549,N_11504,N_10741);
or U12550 (N_12550,N_11274,N_11915);
nand U12551 (N_12551,N_11716,N_11104);
xor U12552 (N_12552,N_11902,N_11800);
nor U12553 (N_12553,N_11599,N_11249);
or U12554 (N_12554,N_9843,N_11285);
nor U12555 (N_12555,N_11813,N_9889);
nand U12556 (N_12556,N_10377,N_10825);
nor U12557 (N_12557,N_11686,N_9570);
and U12558 (N_12558,N_9282,N_9361);
nor U12559 (N_12559,N_11074,N_10783);
nor U12560 (N_12560,N_10061,N_10344);
or U12561 (N_12561,N_11771,N_9691);
nor U12562 (N_12562,N_10032,N_10412);
nand U12563 (N_12563,N_9626,N_10881);
nor U12564 (N_12564,N_9640,N_11174);
nor U12565 (N_12565,N_11203,N_11807);
nand U12566 (N_12566,N_11883,N_11448);
nand U12567 (N_12567,N_9309,N_9840);
nand U12568 (N_12568,N_9924,N_9948);
or U12569 (N_12569,N_11359,N_10439);
nor U12570 (N_12570,N_10866,N_9979);
or U12571 (N_12571,N_11829,N_11956);
and U12572 (N_12572,N_10606,N_10709);
nor U12573 (N_12573,N_11361,N_11491);
xnor U12574 (N_12574,N_10022,N_10531);
nand U12575 (N_12575,N_9234,N_11231);
and U12576 (N_12576,N_9776,N_9600);
and U12577 (N_12577,N_11628,N_10520);
or U12578 (N_12578,N_11306,N_10369);
xnor U12579 (N_12579,N_11037,N_11312);
nand U12580 (N_12580,N_10119,N_10775);
xnor U12581 (N_12581,N_10820,N_11695);
nor U12582 (N_12582,N_10667,N_10429);
nor U12583 (N_12583,N_10087,N_10346);
xor U12584 (N_12584,N_10376,N_9741);
or U12585 (N_12585,N_9721,N_9935);
nor U12586 (N_12586,N_10014,N_9735);
nor U12587 (N_12587,N_10808,N_11256);
or U12588 (N_12588,N_9163,N_10114);
xor U12589 (N_12589,N_9492,N_9009);
and U12590 (N_12590,N_11475,N_9095);
nor U12591 (N_12591,N_11432,N_10748);
nand U12592 (N_12592,N_9685,N_10758);
and U12593 (N_12593,N_10862,N_9464);
nand U12594 (N_12594,N_11750,N_9494);
nand U12595 (N_12595,N_11179,N_9146);
and U12596 (N_12596,N_10564,N_11314);
or U12597 (N_12597,N_9106,N_11506);
nor U12598 (N_12598,N_10626,N_9928);
xor U12599 (N_12599,N_11140,N_11413);
nor U12600 (N_12600,N_11295,N_11127);
xnor U12601 (N_12601,N_10277,N_10943);
xor U12602 (N_12602,N_9219,N_9763);
or U12603 (N_12603,N_11338,N_11134);
or U12604 (N_12604,N_11700,N_11212);
or U12605 (N_12605,N_9634,N_9273);
and U12606 (N_12606,N_11342,N_10393);
nor U12607 (N_12607,N_9227,N_9782);
nand U12608 (N_12608,N_11711,N_10503);
nand U12609 (N_12609,N_11349,N_10095);
xor U12610 (N_12610,N_10536,N_11667);
and U12611 (N_12611,N_11520,N_9676);
and U12612 (N_12612,N_10244,N_10457);
nand U12613 (N_12613,N_11158,N_10192);
xnor U12614 (N_12614,N_9816,N_11624);
and U12615 (N_12615,N_9806,N_10132);
or U12616 (N_12616,N_9860,N_10096);
and U12617 (N_12617,N_10267,N_10629);
xor U12618 (N_12618,N_10036,N_11160);
nor U12619 (N_12619,N_10322,N_9214);
and U12620 (N_12620,N_11891,N_11635);
and U12621 (N_12621,N_10543,N_11828);
xor U12622 (N_12622,N_9245,N_9433);
nand U12623 (N_12623,N_11579,N_9731);
nor U12624 (N_12624,N_10686,N_9565);
or U12625 (N_12625,N_11097,N_9233);
or U12626 (N_12626,N_11260,N_10597);
and U12627 (N_12627,N_10099,N_11042);
and U12628 (N_12628,N_10740,N_10501);
nand U12629 (N_12629,N_11876,N_9065);
xnor U12630 (N_12630,N_9610,N_10926);
nor U12631 (N_12631,N_11632,N_10538);
and U12632 (N_12632,N_9650,N_11294);
xor U12633 (N_12633,N_9975,N_10161);
nor U12634 (N_12634,N_11619,N_9874);
nor U12635 (N_12635,N_10059,N_10387);
and U12636 (N_12636,N_9013,N_10196);
xnor U12637 (N_12637,N_9455,N_10067);
xnor U12638 (N_12638,N_11204,N_9212);
xnor U12639 (N_12639,N_9980,N_9759);
nand U12640 (N_12640,N_10092,N_9419);
or U12641 (N_12641,N_10992,N_10879);
and U12642 (N_12642,N_9232,N_11080);
nor U12643 (N_12643,N_11372,N_11449);
nor U12644 (N_12644,N_11184,N_9373);
or U12645 (N_12645,N_10716,N_9661);
and U12646 (N_12646,N_10753,N_10469);
nor U12647 (N_12647,N_10463,N_9379);
or U12648 (N_12648,N_10619,N_11085);
or U12649 (N_12649,N_11603,N_10581);
xnor U12650 (N_12650,N_9118,N_9954);
nor U12651 (N_12651,N_9885,N_10227);
xnor U12652 (N_12652,N_11492,N_11875);
and U12653 (N_12653,N_10789,N_9030);
xnor U12654 (N_12654,N_11176,N_10777);
and U12655 (N_12655,N_10590,N_9616);
nor U12656 (N_12656,N_10129,N_10932);
nand U12657 (N_12657,N_10365,N_10029);
nor U12658 (N_12658,N_9872,N_9568);
and U12659 (N_12659,N_11180,N_10512);
nor U12660 (N_12660,N_10973,N_11962);
xor U12661 (N_12661,N_11106,N_10127);
or U12662 (N_12662,N_9408,N_9270);
nor U12663 (N_12663,N_10509,N_10602);
and U12664 (N_12664,N_11588,N_9399);
or U12665 (N_12665,N_9664,N_10282);
or U12666 (N_12666,N_11796,N_9043);
and U12667 (N_12667,N_9119,N_11026);
xor U12668 (N_12668,N_9000,N_10035);
nor U12669 (N_12669,N_11581,N_11447);
nor U12670 (N_12670,N_10647,N_11702);
and U12671 (N_12671,N_10380,N_9552);
and U12672 (N_12672,N_9003,N_10184);
nor U12673 (N_12673,N_10838,N_10737);
xnor U12674 (N_12674,N_11118,N_10842);
and U12675 (N_12675,N_10460,N_10481);
nor U12676 (N_12676,N_9078,N_10946);
xor U12677 (N_12677,N_11098,N_11778);
xnor U12678 (N_12678,N_9203,N_11945);
nor U12679 (N_12679,N_11892,N_9774);
nor U12680 (N_12680,N_9894,N_11668);
xnor U12681 (N_12681,N_9495,N_9145);
or U12682 (N_12682,N_11073,N_9809);
xor U12683 (N_12683,N_11946,N_11222);
and U12684 (N_12684,N_11324,N_10534);
xnor U12685 (N_12685,N_9621,N_11056);
or U12686 (N_12686,N_9619,N_11088);
or U12687 (N_12687,N_10359,N_10816);
and U12688 (N_12688,N_11894,N_9991);
nand U12689 (N_12689,N_9941,N_10621);
xor U12690 (N_12690,N_11707,N_11698);
xnor U12691 (N_12691,N_11994,N_9105);
nor U12692 (N_12692,N_11291,N_11068);
and U12693 (N_12693,N_11616,N_10300);
or U12694 (N_12694,N_10762,N_9680);
nand U12695 (N_12695,N_9877,N_11815);
xor U12696 (N_12696,N_9902,N_11861);
xnor U12697 (N_12697,N_10573,N_11092);
xnor U12698 (N_12698,N_11350,N_9498);
nand U12699 (N_12699,N_9915,N_11571);
nand U12700 (N_12700,N_10274,N_9356);
or U12701 (N_12701,N_10329,N_11767);
nor U12702 (N_12702,N_11226,N_9656);
or U12703 (N_12703,N_9181,N_9256);
and U12704 (N_12704,N_9443,N_9134);
nor U12705 (N_12705,N_10898,N_9269);
xnor U12706 (N_12706,N_11276,N_10755);
nand U12707 (N_12707,N_11172,N_10353);
nor U12708 (N_12708,N_9908,N_10077);
xor U12709 (N_12709,N_11196,N_10566);
nor U12710 (N_12710,N_10170,N_11782);
xor U12711 (N_12711,N_9182,N_9939);
nor U12712 (N_12712,N_9099,N_10214);
nand U12713 (N_12713,N_9391,N_10498);
nor U12714 (N_12714,N_11790,N_9237);
and U12715 (N_12715,N_10956,N_10844);
or U12716 (N_12716,N_11830,N_10224);
xnor U12717 (N_12717,N_11096,N_11014);
xnor U12718 (N_12718,N_9158,N_11508);
nor U12719 (N_12719,N_10746,N_10685);
or U12720 (N_12720,N_11914,N_9291);
nor U12721 (N_12721,N_9923,N_11146);
and U12722 (N_12722,N_10712,N_11881);
or U12723 (N_12723,N_11903,N_11981);
and U12724 (N_12724,N_11574,N_11209);
nor U12725 (N_12725,N_11835,N_11677);
xnor U12726 (N_12726,N_9633,N_9487);
xnor U12727 (N_12727,N_11006,N_10079);
nor U12728 (N_12728,N_11939,N_10729);
or U12729 (N_12729,N_10968,N_9693);
and U12730 (N_12730,N_10415,N_10097);
nand U12731 (N_12731,N_10318,N_10979);
or U12732 (N_12732,N_9584,N_10444);
xor U12733 (N_12733,N_9153,N_11801);
xnor U12734 (N_12734,N_11355,N_11683);
and U12735 (N_12735,N_10522,N_9449);
nand U12736 (N_12736,N_11951,N_11591);
or U12737 (N_12737,N_10074,N_11500);
or U12738 (N_12738,N_11055,N_11327);
xnor U12739 (N_12739,N_10863,N_11839);
nor U12740 (N_12740,N_9771,N_11215);
nor U12741 (N_12741,N_9070,N_10893);
and U12742 (N_12742,N_11017,N_11735);
nor U12743 (N_12743,N_11543,N_9171);
nand U12744 (N_12744,N_11286,N_11728);
nand U12745 (N_12745,N_11959,N_11188);
or U12746 (N_12746,N_9343,N_10997);
nor U12747 (N_12747,N_9447,N_10474);
xnor U12748 (N_12748,N_11077,N_9717);
xnor U12749 (N_12749,N_11330,N_11409);
nand U12750 (N_12750,N_11694,N_11275);
or U12751 (N_12751,N_11210,N_10265);
xor U12752 (N_12752,N_10155,N_9281);
and U12753 (N_12753,N_10900,N_9651);
nor U12754 (N_12754,N_11446,N_11206);
xor U12755 (N_12755,N_10064,N_9121);
nand U12756 (N_12756,N_10111,N_10281);
nor U12757 (N_12757,N_11682,N_11562);
xnor U12758 (N_12758,N_10691,N_9097);
or U12759 (N_12759,N_10556,N_9300);
xnor U12760 (N_12760,N_9836,N_10115);
or U12761 (N_12761,N_11110,N_11166);
nor U12762 (N_12762,N_11244,N_9502);
or U12763 (N_12763,N_9350,N_9272);
xor U12764 (N_12764,N_9267,N_11990);
or U12765 (N_12765,N_11394,N_10494);
nand U12766 (N_12766,N_9018,N_9254);
xor U12767 (N_12767,N_9919,N_10578);
or U12768 (N_12768,N_10413,N_11321);
nand U12769 (N_12769,N_10920,N_11198);
nand U12770 (N_12770,N_10394,N_9093);
nand U12771 (N_12771,N_11238,N_9538);
xnor U12772 (N_12772,N_10516,N_10987);
and U12773 (N_12773,N_9223,N_11907);
nand U12774 (N_12774,N_10751,N_11121);
nand U12775 (N_12775,N_11363,N_11109);
xor U12776 (N_12776,N_11331,N_9711);
xnor U12777 (N_12777,N_9315,N_9371);
nand U12778 (N_12778,N_9071,N_10980);
nand U12779 (N_12779,N_11908,N_9441);
nand U12780 (N_12780,N_10402,N_10148);
nand U12781 (N_12781,N_9732,N_9150);
and U12782 (N_12782,N_10773,N_11751);
nor U12783 (N_12783,N_10733,N_11150);
or U12784 (N_12784,N_11858,N_9912);
or U12785 (N_12785,N_9456,N_10361);
nor U12786 (N_12786,N_11793,N_11159);
or U12787 (N_12787,N_10163,N_9758);
nand U12788 (N_12788,N_10419,N_11308);
xor U12789 (N_12789,N_9285,N_10840);
nor U12790 (N_12790,N_9518,N_9109);
nand U12791 (N_12791,N_11028,N_9023);
nor U12792 (N_12792,N_9321,N_10708);
xor U12793 (N_12793,N_11132,N_10238);
and U12794 (N_12794,N_10904,N_9358);
nand U12795 (N_12795,N_10027,N_11613);
nand U12796 (N_12796,N_11473,N_10117);
nor U12797 (N_12797,N_9147,N_9301);
and U12798 (N_12798,N_11153,N_9614);
xor U12799 (N_12799,N_11487,N_11234);
or U12800 (N_12800,N_9704,N_9587);
or U12801 (N_12801,N_10804,N_11388);
xnor U12802 (N_12802,N_11082,N_11246);
and U12803 (N_12803,N_10431,N_10005);
or U12804 (N_12804,N_11566,N_9938);
xnor U12805 (N_12805,N_11278,N_11922);
xnor U12806 (N_12806,N_10794,N_9246);
nand U12807 (N_12807,N_10094,N_10724);
nand U12808 (N_12808,N_10507,N_9956);
or U12809 (N_12809,N_9403,N_11044);
nor U12810 (N_12810,N_9820,N_10193);
xnor U12811 (N_12811,N_10008,N_9006);
and U12812 (N_12812,N_9526,N_11533);
nand U12813 (N_12813,N_11189,N_11009);
or U12814 (N_12814,N_11706,N_10375);
or U12815 (N_12815,N_10315,N_11422);
xnor U12816 (N_12816,N_9094,N_10792);
nor U12817 (N_12817,N_9208,N_11985);
xor U12818 (N_12818,N_9014,N_10178);
nor U12819 (N_12819,N_11594,N_10470);
nand U12820 (N_12820,N_9027,N_9178);
and U12821 (N_12821,N_9995,N_9165);
or U12822 (N_12822,N_10940,N_10210);
xor U12823 (N_12823,N_10324,N_10962);
xor U12824 (N_12824,N_9506,N_9475);
and U12825 (N_12825,N_11396,N_10835);
nor U12826 (N_12826,N_10638,N_9700);
nand U12827 (N_12827,N_10719,N_9002);
nor U12828 (N_12828,N_9335,N_10475);
nor U12829 (N_12829,N_10251,N_11884);
nand U12830 (N_12830,N_10046,N_11941);
and U12831 (N_12831,N_9336,N_10020);
nand U12832 (N_12832,N_11511,N_11015);
nand U12833 (N_12833,N_10678,N_11789);
and U12834 (N_12834,N_9204,N_10867);
and U12835 (N_12835,N_10924,N_11038);
and U12836 (N_12836,N_11722,N_10750);
and U12837 (N_12837,N_10710,N_9342);
or U12838 (N_12838,N_11332,N_9488);
xnor U12839 (N_12839,N_11739,N_11803);
or U12840 (N_12840,N_9957,N_9653);
nand U12841 (N_12841,N_11281,N_9750);
or U12842 (N_12842,N_10383,N_9906);
nand U12843 (N_12843,N_10001,N_11401);
xor U12844 (N_12844,N_11992,N_10550);
xor U12845 (N_12845,N_10829,N_9752);
or U12846 (N_12846,N_11805,N_10409);
and U12847 (N_12847,N_9983,N_11450);
or U12848 (N_12848,N_11838,N_9047);
and U12849 (N_12849,N_9918,N_11649);
nand U12850 (N_12850,N_10106,N_11651);
nand U12851 (N_12851,N_11743,N_10280);
or U12852 (N_12852,N_10544,N_10752);
nand U12853 (N_12853,N_10187,N_11987);
or U12854 (N_12854,N_10440,N_10562);
xnor U12855 (N_12855,N_10433,N_11218);
nand U12856 (N_12856,N_10220,N_10212);
nand U12857 (N_12857,N_11320,N_10101);
or U12858 (N_12858,N_10625,N_11573);
nand U12859 (N_12859,N_11724,N_10961);
or U12860 (N_12860,N_9467,N_11954);
xor U12861 (N_12861,N_9708,N_9781);
xor U12862 (N_12862,N_11069,N_10398);
or U12863 (N_12863,N_10986,N_9831);
or U12864 (N_12864,N_9249,N_11904);
and U12865 (N_12865,N_9334,N_9689);
and U12866 (N_12866,N_11611,N_11343);
xnor U12867 (N_12867,N_11221,N_9961);
or U12868 (N_12868,N_10102,N_10780);
or U12869 (N_12869,N_9762,N_9855);
xnor U12870 (N_12870,N_11755,N_11834);
nor U12871 (N_12871,N_11563,N_9198);
nand U12872 (N_12872,N_9375,N_10253);
nor U12873 (N_12873,N_11003,N_9901);
nand U12874 (N_12874,N_10505,N_11896);
nor U12875 (N_12875,N_10848,N_9553);
and U12876 (N_12876,N_11744,N_11154);
nor U12877 (N_12877,N_9015,N_9388);
and U12878 (N_12878,N_9727,N_9940);
nor U12879 (N_12879,N_9376,N_11019);
or U12880 (N_12880,N_9977,N_11284);
nor U12881 (N_12881,N_11309,N_9738);
and U12882 (N_12882,N_11493,N_9248);
and U12883 (N_12883,N_11736,N_10841);
nor U12884 (N_12884,N_10349,N_9311);
or U12885 (N_12885,N_9293,N_10799);
and U12886 (N_12886,N_9520,N_11168);
nand U12887 (N_12887,N_10004,N_10237);
nand U12888 (N_12888,N_9299,N_11387);
xnor U12889 (N_12889,N_11010,N_11529);
nand U12890 (N_12890,N_10490,N_9623);
nor U12891 (N_12891,N_9169,N_10976);
nand U12892 (N_12892,N_11117,N_11592);
and U12893 (N_12893,N_9937,N_9797);
nor U12894 (N_12894,N_10877,N_9337);
nor U12895 (N_12895,N_10782,N_11034);
or U12896 (N_12896,N_10994,N_10279);
xor U12897 (N_12897,N_11582,N_10510);
xor U12898 (N_12898,N_11781,N_10295);
nor U12899 (N_12899,N_9084,N_10140);
nor U12900 (N_12900,N_9871,N_9148);
or U12901 (N_12901,N_9926,N_10506);
and U12902 (N_12902,N_9143,N_11013);
nor U12903 (N_12903,N_11841,N_11760);
nor U12904 (N_12904,N_9086,N_11423);
nor U12905 (N_12905,N_9332,N_11163);
xor U12906 (N_12906,N_9869,N_10496);
and U12907 (N_12907,N_9740,N_9173);
nand U12908 (N_12908,N_11478,N_10275);
and U12909 (N_12909,N_11382,N_9733);
xnor U12910 (N_12910,N_9172,N_11869);
nor U12911 (N_12911,N_11062,N_11849);
and U12912 (N_12912,N_9482,N_9129);
xor U12913 (N_12913,N_11066,N_9122);
nor U12914 (N_12914,N_11398,N_10278);
nor U12915 (N_12915,N_10028,N_11046);
or U12916 (N_12916,N_9666,N_10000);
and U12917 (N_12917,N_10390,N_9481);
and U12918 (N_12918,N_9438,N_11607);
and U12919 (N_12919,N_9537,N_10568);
and U12920 (N_12920,N_10112,N_10478);
xor U12921 (N_12921,N_9786,N_10989);
nand U12922 (N_12922,N_11947,N_10793);
nor U12923 (N_12923,N_9916,N_11220);
and U12924 (N_12924,N_10033,N_9516);
nor U12925 (N_12925,N_11918,N_9582);
nor U12926 (N_12926,N_11480,N_10456);
or U12927 (N_12927,N_10453,N_11457);
nand U12928 (N_12928,N_10563,N_10580);
nor U12929 (N_12929,N_10273,N_11656);
and U12930 (N_12930,N_11640,N_10513);
or U12931 (N_12931,N_11233,N_9505);
xnor U12932 (N_12932,N_9225,N_10391);
or U12933 (N_12933,N_9461,N_10533);
nand U12934 (N_12934,N_10646,N_9035);
nand U12935 (N_12935,N_9077,N_9694);
xnor U12936 (N_12936,N_10796,N_10914);
nand U12937 (N_12937,N_9524,N_10952);
and U12938 (N_12938,N_11860,N_10213);
nor U12939 (N_12939,N_10334,N_11012);
or U12940 (N_12940,N_10654,N_9681);
or U12941 (N_12941,N_9865,N_10831);
and U12942 (N_12942,N_10160,N_10472);
and U12943 (N_12943,N_9743,N_11402);
nand U12944 (N_12944,N_10204,N_11052);
or U12945 (N_12945,N_9642,N_10493);
and U12946 (N_12946,N_11399,N_11144);
nand U12947 (N_12947,N_10052,N_9213);
and U12948 (N_12948,N_9323,N_11289);
and U12949 (N_12949,N_11867,N_10135);
xor U12950 (N_12950,N_11200,N_9628);
nor U12951 (N_12951,N_11880,N_11297);
and U12952 (N_12952,N_9746,N_10891);
and U12953 (N_12953,N_11137,N_10706);
or U12954 (N_12954,N_9529,N_10931);
nand U12955 (N_12955,N_11322,N_9446);
xnor U12956 (N_12956,N_11183,N_9026);
nor U12957 (N_12957,N_10607,N_9349);
nor U12958 (N_12958,N_9522,N_9250);
xnor U12959 (N_12959,N_9662,N_10362);
nor U12960 (N_12960,N_10627,N_11732);
or U12961 (N_12961,N_9067,N_11191);
nand U12962 (N_12962,N_10718,N_11225);
and U12963 (N_12963,N_11279,N_11729);
nor U12964 (N_12964,N_9778,N_10492);
or U12965 (N_12965,N_10466,N_10585);
nor U12966 (N_12966,N_9525,N_10199);
xnor U12967 (N_12967,N_11490,N_9423);
xor U12968 (N_12968,N_11572,N_10010);
or U12969 (N_12969,N_10872,N_11705);
or U12970 (N_12970,N_10125,N_11773);
nand U12971 (N_12971,N_11693,N_10051);
nand U12972 (N_12972,N_11948,N_9104);
nor U12973 (N_12973,N_10271,N_9080);
nand U12974 (N_12974,N_9936,N_9720);
nand U12975 (N_12975,N_9236,N_10942);
xor U12976 (N_12976,N_10116,N_10222);
and U12977 (N_12977,N_9230,N_9712);
and U12978 (N_12978,N_11065,N_10702);
xor U12979 (N_12979,N_10154,N_10665);
nor U12980 (N_12980,N_10261,N_11123);
xor U12981 (N_12981,N_9578,N_10870);
and U12982 (N_12982,N_9357,N_10250);
xnor U12983 (N_12983,N_9045,N_11569);
and U12984 (N_12984,N_10229,N_10948);
nand U12985 (N_12985,N_10656,N_10368);
xnor U12986 (N_12986,N_10180,N_9318);
xor U12987 (N_12987,N_11786,N_10704);
and U12988 (N_12988,N_11354,N_11392);
nand U12989 (N_12989,N_9319,N_11765);
nand U12990 (N_12990,N_10370,N_10150);
nor U12991 (N_12991,N_9851,N_9428);
or U12992 (N_12992,N_10558,N_9031);
xor U12993 (N_12993,N_10240,N_10188);
nand U12994 (N_12994,N_9298,N_9140);
or U12995 (N_12995,N_11300,N_9892);
nor U12996 (N_12996,N_10201,N_9194);
nor U12997 (N_12997,N_11556,N_10903);
or U12998 (N_12998,N_9765,N_10821);
nand U12999 (N_12999,N_11802,N_11335);
or U13000 (N_13000,N_10895,N_11971);
and U13001 (N_13001,N_9603,N_9396);
or U13002 (N_13002,N_10519,N_11193);
or U13003 (N_13003,N_9333,N_10532);
nand U13004 (N_13004,N_10865,N_11287);
nand U13005 (N_13005,N_9768,N_9325);
xor U13006 (N_13006,N_11966,N_11745);
nor U13007 (N_13007,N_11540,N_10379);
or U13008 (N_13008,N_9861,N_10732);
nand U13009 (N_13009,N_11481,N_10864);
xor U13010 (N_13010,N_9898,N_11036);
nor U13011 (N_13011,N_10373,N_10232);
nor U13012 (N_13012,N_9757,N_10438);
or U13013 (N_13013,N_10386,N_11391);
nand U13014 (N_13014,N_11598,N_10019);
and U13015 (N_13015,N_11479,N_9523);
nor U13016 (N_13016,N_11910,N_10317);
or U13017 (N_13017,N_11089,N_9969);
and U13018 (N_13018,N_11201,N_10690);
xnor U13019 (N_13019,N_11208,N_9052);
or U13020 (N_13020,N_9152,N_9406);
xnor U13021 (N_13021,N_9351,N_11075);
xnor U13022 (N_13022,N_9822,N_10771);
or U13023 (N_13023,N_9004,N_11629);
xor U13024 (N_13024,N_11299,N_11237);
or U13025 (N_13025,N_9669,N_9751);
xnor U13026 (N_13026,N_11439,N_9715);
and U13027 (N_13027,N_11614,N_10738);
nand U13028 (N_13028,N_10639,N_9159);
or U13029 (N_13029,N_11471,N_9635);
or U13030 (N_13030,N_9497,N_11909);
or U13031 (N_13031,N_10614,N_9688);
xnor U13032 (N_13032,N_10555,N_9057);
and U13033 (N_13033,N_9657,N_11458);
and U13034 (N_13034,N_11277,N_9205);
nand U13035 (N_13035,N_11049,N_9804);
xor U13036 (N_13036,N_9137,N_11590);
xnor U13037 (N_13037,N_10396,N_10802);
or U13038 (N_13038,N_9791,N_9044);
xnor U13039 (N_13039,N_11905,N_10450);
nand U13040 (N_13040,N_10177,N_10800);
nand U13041 (N_13041,N_11758,N_10294);
or U13042 (N_13042,N_9819,N_10632);
nor U13043 (N_13043,N_10959,N_11963);
nor U13044 (N_13044,N_9703,N_9866);
nor U13045 (N_13045,N_11323,N_9192);
and U13046 (N_13046,N_11072,N_11022);
and U13047 (N_13047,N_10068,N_9385);
and U13048 (N_13048,N_10913,N_10347);
and U13049 (N_13049,N_11991,N_9226);
xor U13050 (N_13050,N_9543,N_9393);
nand U13051 (N_13051,N_11970,N_9511);
xnor U13052 (N_13052,N_10323,N_10886);
and U13053 (N_13053,N_9943,N_10795);
nand U13054 (N_13054,N_9294,N_9259);
xnor U13055 (N_13055,N_9627,N_9485);
nand U13056 (N_13056,N_10873,N_11618);
nor U13057 (N_13057,N_11888,N_11242);
nor U13058 (N_13058,N_9370,N_9810);
xnor U13059 (N_13059,N_9295,N_11271);
nand U13060 (N_13060,N_10185,N_11878);
nand U13061 (N_13061,N_10384,N_11169);
xor U13062 (N_13062,N_11641,N_11000);
or U13063 (N_13063,N_9593,N_9566);
or U13064 (N_13064,N_9200,N_11427);
or U13065 (N_13065,N_9679,N_10139);
nor U13066 (N_13066,N_10743,N_11748);
xnor U13067 (N_13067,N_11095,N_11358);
nor U13068 (N_13068,N_10529,N_10205);
and U13069 (N_13069,N_11091,N_9317);
or U13070 (N_13070,N_9020,N_9789);
or U13071 (N_13071,N_10676,N_9997);
or U13072 (N_13072,N_11455,N_9852);
and U13073 (N_13073,N_10181,N_10515);
nand U13074 (N_13074,N_10287,N_11552);
xnor U13075 (N_13075,N_9457,N_10031);
nand U13076 (N_13076,N_10784,N_11319);
xnor U13077 (N_13077,N_9224,N_11669);
and U13078 (N_13078,N_11548,N_11819);
and U13079 (N_13079,N_10599,N_9773);
xor U13080 (N_13080,N_10611,N_9562);
nand U13081 (N_13081,N_11336,N_11488);
and U13082 (N_13082,N_11400,N_9952);
nor U13083 (N_13083,N_10037,N_9063);
and U13084 (N_13084,N_9117,N_11559);
xor U13085 (N_13085,N_10576,N_11610);
or U13086 (N_13086,N_9075,N_11950);
nand U13087 (N_13087,N_10047,N_11532);
nor U13088 (N_13088,N_10594,N_9542);
xor U13089 (N_13089,N_9971,N_9390);
nor U13090 (N_13090,N_9378,N_9029);
or U13091 (N_13091,N_11670,N_10400);
xor U13092 (N_13092,N_10892,N_10420);
nor U13093 (N_13093,N_10905,N_10108);
and U13094 (N_13094,N_10488,N_9096);
xnor U13095 (N_13095,N_11425,N_11099);
nor U13096 (N_13096,N_11083,N_9314);
nor U13097 (N_13097,N_9400,N_10497);
and U13098 (N_13098,N_10442,N_11895);
and U13099 (N_13099,N_10105,N_9327);
and U13100 (N_13100,N_10348,N_9082);
and U13101 (N_13101,N_11486,N_9141);
nor U13102 (N_13102,N_9856,N_10571);
nand U13103 (N_13103,N_9202,N_10290);
nand U13104 (N_13104,N_9784,N_11712);
nor U13105 (N_13105,N_11507,N_10157);
nand U13106 (N_13106,N_11293,N_11928);
nand U13107 (N_13107,N_9284,N_10809);
nor U13108 (N_13108,N_10991,N_11041);
or U13109 (N_13109,N_11433,N_10128);
nand U13110 (N_13110,N_11938,N_10612);
or U13111 (N_13111,N_9521,N_9326);
and U13112 (N_13112,N_11148,N_10745);
and U13113 (N_13113,N_11857,N_9135);
nand U13114 (N_13114,N_9431,N_10996);
xnor U13115 (N_13115,N_10939,N_10651);
nor U13116 (N_13116,N_9658,N_11005);
xnor U13117 (N_13117,N_9599,N_10399);
and U13118 (N_13118,N_9220,N_11245);
and U13119 (N_13119,N_9785,N_10927);
and U13120 (N_13120,N_10768,N_9792);
nand U13121 (N_13121,N_9848,N_9641);
and U13122 (N_13122,N_10811,N_11967);
and U13123 (N_13123,N_9466,N_11756);
nand U13124 (N_13124,N_9352,N_10190);
or U13125 (N_13125,N_11926,N_11395);
nor U13126 (N_13126,N_9576,N_9131);
nor U13127 (N_13127,N_11818,N_9142);
nand U13128 (N_13128,N_10122,N_10541);
nor U13129 (N_13129,N_9609,N_11311);
nor U13130 (N_13130,N_9499,N_11326);
and U13131 (N_13131,N_10367,N_10711);
nor U13132 (N_13132,N_9905,N_11551);
xnor U13133 (N_13133,N_10854,N_9968);
or U13134 (N_13134,N_10395,N_9953);
nand U13135 (N_13135,N_10165,N_10441);
or U13136 (N_13136,N_9372,N_9185);
nand U13137 (N_13137,N_11952,N_9690);
or U13138 (N_13138,N_9713,N_9346);
nor U13139 (N_13139,N_9288,N_9972);
and U13140 (N_13140,N_10843,N_9826);
and U13141 (N_13141,N_11982,N_11105);
nor U13142 (N_13142,N_11853,N_11820);
xnor U13143 (N_13143,N_10884,N_11107);
xnor U13144 (N_13144,N_9102,N_9331);
and U13145 (N_13145,N_10700,N_10500);
nand U13146 (N_13146,N_9512,N_9618);
nor U13147 (N_13147,N_10171,N_10351);
nand U13148 (N_13148,N_11020,N_11832);
and U13149 (N_13149,N_9201,N_10417);
and U13150 (N_13150,N_10591,N_11615);
xnor U13151 (N_13151,N_9660,N_10919);
nor U13152 (N_13152,N_9215,N_10549);
nand U13153 (N_13153,N_9432,N_11050);
nand U13154 (N_13154,N_11973,N_11659);
and U13155 (N_13155,N_11779,N_10455);
xor U13156 (N_13156,N_9678,N_10934);
xor U13157 (N_13157,N_11418,N_11384);
xnor U13158 (N_13158,N_10257,N_9041);
and U13159 (N_13159,N_9594,N_11932);
nor U13160 (N_13160,N_10828,N_11725);
nand U13161 (N_13161,N_11747,N_10769);
and U13162 (N_13162,N_10093,N_10539);
nor U13163 (N_13163,N_10151,N_9698);
and U13164 (N_13164,N_11780,N_11901);
and U13165 (N_13165,N_9302,N_9585);
or U13166 (N_13166,N_9887,N_9583);
xor U13167 (N_13167,N_10147,N_9607);
xor U13168 (N_13168,N_10696,N_10548);
nand U13169 (N_13169,N_11921,N_11647);
nand U13170 (N_13170,N_9128,N_11063);
nand U13171 (N_13171,N_10408,N_10424);
and U13172 (N_13172,N_11810,N_9062);
nand U13173 (N_13173,N_9207,N_10072);
or U13174 (N_13174,N_9779,N_9864);
nand U13175 (N_13175,N_10669,N_11410);
xor U13176 (N_13176,N_11737,N_11787);
xnor U13177 (N_13177,N_11251,N_10234);
and U13178 (N_13178,N_10207,N_11865);
nor U13179 (N_13179,N_9531,N_9313);
nor U13180 (N_13180,N_9963,N_10834);
nand U13181 (N_13181,N_10680,N_10679);
nand U13182 (N_13182,N_11792,N_10981);
or U13183 (N_13183,N_9837,N_10683);
xnor U13184 (N_13184,N_9801,N_9266);
nand U13185 (N_13185,N_9384,N_10426);
nand U13186 (N_13186,N_11988,N_11496);
nor U13187 (N_13187,N_11764,N_9845);
nand U13188 (N_13188,N_9089,N_10104);
nor U13189 (N_13189,N_11636,N_10642);
nor U13190 (N_13190,N_10034,N_10363);
and U13191 (N_13191,N_10906,N_10197);
and U13192 (N_13192,N_11023,N_9191);
xor U13193 (N_13193,N_10527,N_10975);
xnor U13194 (N_13194,N_11627,N_11623);
nor U13195 (N_13195,N_9136,N_9364);
nor U13196 (N_13196,N_9175,N_10159);
nor U13197 (N_13197,N_10805,N_9807);
nor U13198 (N_13198,N_11544,N_11923);
xnor U13199 (N_13199,N_9632,N_9493);
nor U13200 (N_13200,N_9636,N_9794);
nand U13201 (N_13201,N_10857,N_10113);
nor U13202 (N_13202,N_10465,N_9231);
nand U13203 (N_13203,N_9563,N_11408);
xnor U13204 (N_13204,N_9970,N_9439);
and U13205 (N_13205,N_9596,N_10332);
nand U13206 (N_13206,N_10073,N_9021);
and U13207 (N_13207,N_10672,N_10152);
nor U13208 (N_13208,N_9186,N_11494);
nand U13209 (N_13209,N_9415,N_10878);
nor U13210 (N_13210,N_9276,N_9886);
nand U13211 (N_13211,N_10569,N_9699);
xor U13212 (N_13212,N_11054,N_9435);
and U13213 (N_13213,N_10126,N_11419);
or U13214 (N_13214,N_9413,N_10635);
nor U13215 (N_13215,N_11444,N_10209);
nor U13216 (N_13216,N_10437,N_9120);
xnor U13217 (N_13217,N_9074,N_10006);
nand U13218 (N_13218,N_11270,N_11822);
nand U13219 (N_13219,N_11476,N_9654);
or U13220 (N_13220,N_10427,N_10885);
nor U13221 (N_13221,N_10674,N_11045);
or U13222 (N_13222,N_10208,N_10268);
nand U13223 (N_13223,N_9823,N_11974);
and U13224 (N_13224,N_10138,N_11757);
or U13225 (N_13225,N_10876,N_10342);
xnor U13226 (N_13226,N_9539,N_11031);
and U13227 (N_13227,N_11536,N_9815);
or U13228 (N_13228,N_10567,N_11816);
or U13229 (N_13229,N_10338,N_10473);
and U13230 (N_13230,N_10285,N_11165);
and U13231 (N_13231,N_9243,N_10684);
and U13232 (N_13232,N_10305,N_10340);
and U13233 (N_13233,N_11577,N_9934);
and U13234 (N_13234,N_9167,N_11178);
xnor U13235 (N_13235,N_11759,N_10776);
nor U13236 (N_13236,N_9195,N_9881);
nor U13237 (N_13237,N_11043,N_11783);
nor U13238 (N_13238,N_10216,N_9340);
nor U13239 (N_13239,N_9174,N_11371);
xnor U13240 (N_13240,N_11997,N_11531);
nor U13241 (N_13241,N_9580,N_10790);
nor U13242 (N_13242,N_10162,N_11898);
nand U13243 (N_13243,N_11177,N_10728);
and U13244 (N_13244,N_9546,N_9579);
and U13245 (N_13245,N_11977,N_11029);
nor U13246 (N_13246,N_9183,N_10215);
nor U13247 (N_13247,N_10389,N_9079);
nand U13248 (N_13248,N_11680,N_9477);
and U13249 (N_13249,N_9046,N_10837);
nor U13250 (N_13250,N_10869,N_11261);
xor U13251 (N_13251,N_10352,N_11048);
xor U13252 (N_13252,N_11578,N_11989);
nand U13253 (N_13253,N_11298,N_10761);
and U13254 (N_13254,N_10447,N_10003);
nor U13255 (N_13255,N_10336,N_11564);
nand U13256 (N_13256,N_10366,N_10451);
xor U13257 (N_13257,N_10978,N_9049);
or U13258 (N_13258,N_9155,N_10043);
nor U13259 (N_13259,N_9999,N_10316);
and U13260 (N_13260,N_10551,N_9558);
nand U13261 (N_13261,N_9292,N_10668);
xnor U13262 (N_13262,N_10012,N_11002);
xnor U13263 (N_13263,N_9707,N_11502);
nand U13264 (N_13264,N_9133,N_11840);
xor U13265 (N_13265,N_10947,N_9667);
nand U13266 (N_13266,N_11368,N_10289);
xnor U13267 (N_13267,N_11267,N_9180);
nor U13268 (N_13268,N_9149,N_10995);
nor U13269 (N_13269,N_9850,N_9692);
nand U13270 (N_13270,N_9749,N_11937);
nor U13271 (N_13271,N_10374,N_10561);
nor U13272 (N_13272,N_9728,N_9942);
nand U13273 (N_13273,N_11996,N_9103);
nor U13274 (N_13274,N_11375,N_11523);
and U13275 (N_13275,N_11740,N_10574);
nand U13276 (N_13276,N_11788,N_9530);
and U13277 (N_13277,N_11353,N_11709);
or U13278 (N_13278,N_9092,N_11021);
or U13279 (N_13279,N_10965,N_10836);
xor U13280 (N_13280,N_10245,N_11675);
nor U13281 (N_13281,N_9459,N_9469);
nand U13282 (N_13282,N_10146,N_9130);
and U13283 (N_13283,N_10231,N_10044);
or U13284 (N_13284,N_11927,N_10812);
xnor U13285 (N_13285,N_11445,N_9604);
nand U13286 (N_13286,N_10360,N_10735);
nor U13287 (N_13287,N_10038,N_9586);
nand U13288 (N_13288,N_9462,N_11374);
xor U13289 (N_13289,N_10428,N_9387);
xor U13290 (N_13290,N_11701,N_9841);
nand U13291 (N_13291,N_9535,N_10153);
nand U13292 (N_13292,N_9947,N_10670);
nand U13293 (N_13293,N_11660,N_11863);
xor U13294 (N_13294,N_9115,N_11257);
and U13295 (N_13295,N_11376,N_11824);
or U13296 (N_13296,N_9718,N_9412);
nand U13297 (N_13297,N_10060,N_11855);
and U13298 (N_13298,N_9612,N_9675);
nor U13299 (N_13299,N_9931,N_11162);
and U13300 (N_13300,N_10009,N_10086);
xnor U13301 (N_13301,N_10788,N_9595);
nor U13302 (N_13302,N_9608,N_11586);
nor U13303 (N_13303,N_10482,N_11606);
nor U13304 (N_13304,N_10514,N_9976);
xnor U13305 (N_13305,N_9257,N_10637);
xor U13306 (N_13306,N_11899,N_9458);
xnor U13307 (N_13307,N_9280,N_11337);
and U13308 (N_13308,N_10381,N_11741);
xnor U13309 (N_13309,N_10200,N_11567);
nor U13310 (N_13310,N_10264,N_11526);
and U13311 (N_13311,N_11452,N_9899);
xnor U13312 (N_13312,N_11313,N_10526);
xor U13313 (N_13313,N_11428,N_9591);
or U13314 (N_13314,N_11101,N_11514);
xnor U13315 (N_13315,N_9241,N_9847);
nor U13316 (N_13316,N_10401,N_11157);
xnor U13317 (N_13317,N_9389,N_9088);
or U13318 (N_13318,N_9193,N_9862);
nand U13319 (N_13319,N_10817,N_11558);
nand U13320 (N_13320,N_9988,N_9383);
xnor U13321 (N_13321,N_11139,N_10944);
xnor U13322 (N_13322,N_11887,N_11283);
nor U13323 (N_13323,N_10327,N_10765);
nand U13324 (N_13324,N_11255,N_9264);
nand U13325 (N_13325,N_9590,N_9714);
nor U13326 (N_13326,N_10766,N_11654);
nor U13327 (N_13327,N_9032,N_10491);
and U13328 (N_13328,N_11217,N_11018);
xnor U13329 (N_13329,N_11348,N_10972);
xor U13330 (N_13330,N_10175,N_9913);
xnor U13331 (N_13331,N_10839,N_9629);
or U13332 (N_13332,N_9510,N_9239);
xor U13333 (N_13333,N_9532,N_10615);
nand U13334 (N_13334,N_10182,N_9416);
xnor U13335 (N_13335,N_11463,N_9085);
or U13336 (N_13336,N_10283,N_10554);
and U13337 (N_13337,N_11435,N_11785);
or U13338 (N_13338,N_10982,N_10057);
and U13339 (N_13339,N_11053,N_11194);
or U13340 (N_13340,N_11897,N_9966);
xor U13341 (N_13341,N_9187,N_9519);
nor U13342 (N_13342,N_11173,N_11429);
nor U13343 (N_13343,N_9748,N_11357);
nor U13344 (N_13344,N_11417,N_10887);
nor U13345 (N_13345,N_10617,N_11547);
and U13346 (N_13346,N_11472,N_11509);
xor U13347 (N_13347,N_11280,N_11119);
and U13348 (N_13348,N_10977,N_9452);
or U13349 (N_13349,N_9420,N_10661);
or U13350 (N_13350,N_9846,N_10299);
xor U13351 (N_13351,N_11135,N_10963);
or U13352 (N_13352,N_10725,N_10757);
or U13353 (N_13353,N_11774,N_11389);
and U13354 (N_13354,N_11626,N_9625);
xnor U13355 (N_13355,N_9010,N_9430);
xnor U13356 (N_13356,N_11236,N_9116);
or U13357 (N_13357,N_10747,N_9756);
xor U13358 (N_13358,N_11434,N_10011);
and U13359 (N_13359,N_9209,N_9161);
nor U13360 (N_13360,N_9076,N_11804);
and U13361 (N_13361,N_10123,N_9274);
or U13362 (N_13362,N_10489,N_10330);
nand U13363 (N_13363,N_11605,N_10259);
and U13364 (N_13364,N_11944,N_11345);
xnor U13365 (N_13365,N_9409,N_11879);
or U13366 (N_13366,N_10918,N_9652);
nand U13367 (N_13367,N_9470,N_11752);
or U13368 (N_13368,N_11964,N_11886);
xor U13369 (N_13369,N_10849,N_11856);
nor U13370 (N_13370,N_9544,N_9813);
nor U13371 (N_13371,N_10810,N_11678);
nor U13372 (N_13372,N_10343,N_11130);
xor U13373 (N_13373,N_11216,N_9054);
nor U13374 (N_13374,N_11584,N_9557);
and U13375 (N_13375,N_10252,N_10858);
nor U13376 (N_13376,N_10041,N_10149);
nor U13377 (N_13377,N_11024,N_9051);
or U13378 (N_13378,N_11949,N_10076);
nand U13379 (N_13379,N_9788,N_10855);
or U13380 (N_13380,N_10645,N_9286);
and U13381 (N_13381,N_11555,N_11929);
nand U13382 (N_13382,N_9853,N_10260);
xnor U13383 (N_13383,N_11549,N_11806);
and U13384 (N_13384,N_9888,N_9805);
and U13385 (N_13385,N_9802,N_9261);
or U13386 (N_13386,N_11761,N_10055);
xnor U13387 (N_13387,N_11827,N_9196);
xnor U13388 (N_13388,N_9833,N_11094);
and U13389 (N_13389,N_10622,N_9476);
nand U13390 (N_13390,N_10889,N_10406);
xnor U13391 (N_13391,N_11664,N_9283);
and U13392 (N_13392,N_11864,N_9615);
nor U13393 (N_13393,N_10082,N_10504);
xnor U13394 (N_13394,N_10272,N_10435);
and U13395 (N_13395,N_9895,N_9091);
nand U13396 (N_13396,N_11731,N_11699);
nor U13397 (N_13397,N_9184,N_11595);
or U13398 (N_13398,N_11461,N_11550);
and U13399 (N_13399,N_9574,N_11290);
nand U13400 (N_13400,N_11972,N_9238);
xor U13401 (N_13401,N_11580,N_10266);
nand U13402 (N_13402,N_11850,N_10355);
or U13403 (N_13403,N_11602,N_9110);
and U13404 (N_13404,N_9426,N_11230);
nand U13405 (N_13405,N_10689,N_9229);
xnor U13406 (N_13406,N_9946,N_11596);
and U13407 (N_13407,N_10518,N_11474);
xor U13408 (N_13408,N_9648,N_9973);
xnor U13409 (N_13409,N_9958,N_10226);
xnor U13410 (N_13410,N_10915,N_10969);
xor U13411 (N_13411,N_9673,N_10720);
or U13412 (N_13412,N_11039,N_10999);
xnor U13413 (N_13413,N_11631,N_10653);
nand U13414 (N_13414,N_11798,N_9139);
xor U13415 (N_13415,N_10007,N_9036);
nor U13416 (N_13416,N_10203,N_9168);
nor U13417 (N_13417,N_9893,N_11671);
and U13418 (N_13418,N_10949,N_10276);
or U13419 (N_13419,N_11087,N_10721);
nor U13420 (N_13420,N_9780,N_11414);
nor U13421 (N_13421,N_9911,N_11622);
xor U13422 (N_13422,N_9734,N_9068);
nor U13423 (N_13423,N_11519,N_9639);
and U13424 (N_13424,N_9904,N_11512);
nand U13425 (N_13425,N_10786,N_11430);
nor U13426 (N_13426,N_11673,N_9341);
xor U13427 (N_13427,N_10502,N_11528);
nor U13428 (N_13428,N_9404,N_9719);
nor U13429 (N_13429,N_11001,N_11882);
or U13430 (N_13430,N_9417,N_9766);
xor U13431 (N_13431,N_11995,N_11604);
and U13432 (N_13432,N_10487,N_11542);
and U13433 (N_13433,N_10859,N_11652);
xnor U13434 (N_13434,N_11064,N_11248);
nand U13435 (N_13435,N_11924,N_9879);
or U13436 (N_13436,N_9454,N_11304);
and U13437 (N_13437,N_11443,N_9663);
xnor U13438 (N_13438,N_9998,N_10584);
or U13439 (N_13439,N_10486,N_10025);
and U13440 (N_13440,N_11643,N_10850);
nor U13441 (N_13441,N_10284,N_10671);
and U13442 (N_13442,N_10871,N_11738);
or U13443 (N_13443,N_11642,N_11889);
nand U13444 (N_13444,N_11733,N_9655);
nor U13445 (N_13445,N_9108,N_9268);
nor U13446 (N_13446,N_10530,N_11851);
xor U13447 (N_13447,N_9395,N_10604);
xor U13448 (N_13448,N_9304,N_11746);
nand U13449 (N_13449,N_9465,N_10249);
nor U13450 (N_13450,N_11842,N_11541);
and U13451 (N_13451,N_9870,N_11303);
xor U13452 (N_13452,N_11576,N_9038);
and U13453 (N_13453,N_9835,N_9637);
xor U13454 (N_13454,N_9548,N_9124);
and U13455 (N_13455,N_11704,N_9382);
xor U13456 (N_13456,N_11464,N_9921);
or U13457 (N_13457,N_11762,N_9123);
nor U13458 (N_13458,N_11534,N_11657);
and U13459 (N_13459,N_11638,N_9468);
xnor U13460 (N_13460,N_9263,N_11004);
nand U13461 (N_13461,N_9287,N_10923);
and U13462 (N_13462,N_11553,N_10350);
and U13463 (N_13463,N_11317,N_9555);
xnor U13464 (N_13464,N_11585,N_10084);
xor U13465 (N_13465,N_9271,N_9925);
xor U13466 (N_13466,N_9821,N_10756);
nand U13467 (N_13467,N_11420,N_9033);
nand U13468 (N_13468,N_9386,N_11318);
xor U13469 (N_13469,N_11272,N_10605);
or U13470 (N_13470,N_9551,N_9808);
and U13471 (N_13471,N_10477,N_11047);
or U13472 (N_13472,N_9491,N_11516);
or U13473 (N_13473,N_9687,N_11930);
and U13474 (N_13474,N_11202,N_10091);
xnor U13475 (N_13475,N_10801,N_11817);
xor U13476 (N_13476,N_9764,N_11868);
xnor U13477 (N_13477,N_10254,N_9440);
nand U13478 (N_13478,N_9672,N_11161);
and U13479 (N_13479,N_9090,N_11128);
and U13480 (N_13480,N_9817,N_10693);
and U13481 (N_13481,N_10930,N_11437);
nor U13482 (N_13482,N_11503,N_10017);
nand U13483 (N_13483,N_9598,N_10846);
nand U13484 (N_13484,N_10241,N_10587);
nor U13485 (N_13485,N_9262,N_9448);
or U13486 (N_13486,N_11634,N_11639);
xor U13487 (N_13487,N_11489,N_11933);
xor U13488 (N_13488,N_9437,N_9176);
xor U13489 (N_13489,N_9829,N_9347);
and U13490 (N_13490,N_9875,N_11468);
nor U13491 (N_13491,N_11655,N_9344);
xor U13492 (N_13492,N_9910,N_9251);
and U13493 (N_13493,N_9818,N_10875);
and U13494 (N_13494,N_9019,N_9138);
or U13495 (N_13495,N_11593,N_9965);
nor U13496 (N_13496,N_9962,N_11404);
or U13497 (N_13497,N_9418,N_11131);
nor U13498 (N_13498,N_11315,N_10593);
and U13499 (N_13499,N_11268,N_9745);
xor U13500 (N_13500,N_9411,N_10341);
nor U13501 (N_13501,N_10254,N_10941);
nand U13502 (N_13502,N_11100,N_10220);
nand U13503 (N_13503,N_9941,N_10393);
nand U13504 (N_13504,N_11396,N_9989);
xnor U13505 (N_13505,N_9129,N_11780);
xnor U13506 (N_13506,N_11064,N_9964);
nand U13507 (N_13507,N_11940,N_10320);
or U13508 (N_13508,N_9363,N_10396);
or U13509 (N_13509,N_10566,N_9679);
or U13510 (N_13510,N_10237,N_11950);
and U13511 (N_13511,N_11518,N_11614);
nand U13512 (N_13512,N_9546,N_9581);
nand U13513 (N_13513,N_10159,N_9837);
nor U13514 (N_13514,N_11996,N_10323);
or U13515 (N_13515,N_11593,N_10490);
xnor U13516 (N_13516,N_9426,N_10963);
nor U13517 (N_13517,N_9132,N_11534);
nor U13518 (N_13518,N_9892,N_11361);
xor U13519 (N_13519,N_10077,N_9425);
or U13520 (N_13520,N_9123,N_10961);
xor U13521 (N_13521,N_9379,N_9173);
or U13522 (N_13522,N_11850,N_11924);
nand U13523 (N_13523,N_11652,N_10515);
nand U13524 (N_13524,N_11188,N_11217);
nor U13525 (N_13525,N_11099,N_9368);
nand U13526 (N_13526,N_11573,N_9260);
nand U13527 (N_13527,N_9563,N_9458);
and U13528 (N_13528,N_9513,N_10643);
xnor U13529 (N_13529,N_11295,N_11443);
nor U13530 (N_13530,N_11979,N_11910);
nand U13531 (N_13531,N_9729,N_9561);
or U13532 (N_13532,N_10745,N_10630);
or U13533 (N_13533,N_9222,N_10526);
nand U13534 (N_13534,N_11418,N_10771);
xor U13535 (N_13535,N_11169,N_11998);
or U13536 (N_13536,N_11652,N_9630);
nand U13537 (N_13537,N_10457,N_11383);
nor U13538 (N_13538,N_11122,N_11932);
and U13539 (N_13539,N_10840,N_9909);
nand U13540 (N_13540,N_10580,N_10449);
or U13541 (N_13541,N_9012,N_11599);
nand U13542 (N_13542,N_10365,N_9101);
xnor U13543 (N_13543,N_9880,N_10779);
nor U13544 (N_13544,N_10583,N_9413);
nor U13545 (N_13545,N_11651,N_10342);
or U13546 (N_13546,N_9784,N_11905);
and U13547 (N_13547,N_9087,N_9376);
or U13548 (N_13548,N_10284,N_9811);
xor U13549 (N_13549,N_11676,N_10851);
nand U13550 (N_13550,N_11096,N_10601);
and U13551 (N_13551,N_11905,N_10163);
or U13552 (N_13552,N_10214,N_9426);
nand U13553 (N_13553,N_11855,N_9549);
and U13554 (N_13554,N_11934,N_9794);
and U13555 (N_13555,N_10583,N_9397);
nand U13556 (N_13556,N_11459,N_10871);
xor U13557 (N_13557,N_10835,N_11579);
or U13558 (N_13558,N_9338,N_10347);
xor U13559 (N_13559,N_9534,N_11976);
nor U13560 (N_13560,N_11584,N_10700);
xnor U13561 (N_13561,N_9545,N_9279);
and U13562 (N_13562,N_10790,N_11945);
xor U13563 (N_13563,N_11393,N_10358);
and U13564 (N_13564,N_9224,N_11442);
nand U13565 (N_13565,N_11894,N_11840);
nand U13566 (N_13566,N_10007,N_9607);
and U13567 (N_13567,N_9183,N_10237);
and U13568 (N_13568,N_11073,N_9355);
or U13569 (N_13569,N_10939,N_11851);
nand U13570 (N_13570,N_10674,N_9147);
or U13571 (N_13571,N_11328,N_11926);
nor U13572 (N_13572,N_10543,N_10689);
or U13573 (N_13573,N_10692,N_11267);
and U13574 (N_13574,N_10693,N_9302);
and U13575 (N_13575,N_10417,N_11807);
or U13576 (N_13576,N_9678,N_11276);
nand U13577 (N_13577,N_9347,N_11492);
or U13578 (N_13578,N_10091,N_9554);
nor U13579 (N_13579,N_11109,N_10892);
nand U13580 (N_13580,N_11991,N_11787);
and U13581 (N_13581,N_10717,N_10319);
xnor U13582 (N_13582,N_9485,N_10877);
nand U13583 (N_13583,N_10125,N_11592);
and U13584 (N_13584,N_11393,N_10937);
nand U13585 (N_13585,N_11514,N_11382);
nor U13586 (N_13586,N_9772,N_9113);
and U13587 (N_13587,N_10968,N_11204);
or U13588 (N_13588,N_11957,N_10056);
and U13589 (N_13589,N_11327,N_10520);
xnor U13590 (N_13590,N_11685,N_9761);
or U13591 (N_13591,N_9242,N_11512);
nor U13592 (N_13592,N_11828,N_9085);
and U13593 (N_13593,N_9171,N_10662);
nor U13594 (N_13594,N_11302,N_10234);
nand U13595 (N_13595,N_11673,N_9012);
xnor U13596 (N_13596,N_10526,N_10564);
or U13597 (N_13597,N_10109,N_9285);
xor U13598 (N_13598,N_10127,N_11977);
or U13599 (N_13599,N_11983,N_9219);
xor U13600 (N_13600,N_9965,N_9306);
or U13601 (N_13601,N_9631,N_9161);
or U13602 (N_13602,N_9780,N_10852);
and U13603 (N_13603,N_9789,N_10054);
or U13604 (N_13604,N_9890,N_11246);
xnor U13605 (N_13605,N_9394,N_11977);
xnor U13606 (N_13606,N_9237,N_11557);
nor U13607 (N_13607,N_11002,N_9117);
or U13608 (N_13608,N_11786,N_9201);
nand U13609 (N_13609,N_10140,N_10492);
and U13610 (N_13610,N_11145,N_10593);
nand U13611 (N_13611,N_10415,N_10324);
nor U13612 (N_13612,N_9285,N_9129);
nor U13613 (N_13613,N_11695,N_11846);
and U13614 (N_13614,N_9236,N_9957);
or U13615 (N_13615,N_10220,N_11945);
nor U13616 (N_13616,N_11684,N_9136);
and U13617 (N_13617,N_9366,N_9200);
and U13618 (N_13618,N_10401,N_9355);
nor U13619 (N_13619,N_10423,N_10783);
and U13620 (N_13620,N_10587,N_9088);
nor U13621 (N_13621,N_11167,N_11363);
and U13622 (N_13622,N_9532,N_9251);
nor U13623 (N_13623,N_10799,N_10377);
and U13624 (N_13624,N_9641,N_10364);
or U13625 (N_13625,N_11874,N_11674);
nand U13626 (N_13626,N_11437,N_10312);
or U13627 (N_13627,N_11293,N_9775);
and U13628 (N_13628,N_9752,N_9719);
or U13629 (N_13629,N_11809,N_9873);
nand U13630 (N_13630,N_11548,N_11897);
nand U13631 (N_13631,N_9861,N_9165);
xor U13632 (N_13632,N_10636,N_10378);
nor U13633 (N_13633,N_11933,N_9833);
nor U13634 (N_13634,N_11043,N_11357);
or U13635 (N_13635,N_10590,N_9471);
nand U13636 (N_13636,N_11104,N_11957);
xnor U13637 (N_13637,N_11835,N_9168);
and U13638 (N_13638,N_9978,N_10996);
nor U13639 (N_13639,N_10775,N_10822);
nor U13640 (N_13640,N_11545,N_9393);
nand U13641 (N_13641,N_10386,N_10011);
and U13642 (N_13642,N_9441,N_11892);
or U13643 (N_13643,N_10899,N_10096);
xor U13644 (N_13644,N_9494,N_10365);
nor U13645 (N_13645,N_10577,N_10192);
nand U13646 (N_13646,N_11497,N_11859);
nand U13647 (N_13647,N_9268,N_10339);
nand U13648 (N_13648,N_10913,N_10094);
xnor U13649 (N_13649,N_11252,N_10337);
and U13650 (N_13650,N_11568,N_9807);
xnor U13651 (N_13651,N_10491,N_11454);
nor U13652 (N_13652,N_9134,N_9774);
and U13653 (N_13653,N_9903,N_11341);
and U13654 (N_13654,N_9756,N_10044);
or U13655 (N_13655,N_9471,N_11587);
xor U13656 (N_13656,N_11684,N_9168);
and U13657 (N_13657,N_9366,N_9577);
and U13658 (N_13658,N_10237,N_11540);
nor U13659 (N_13659,N_9712,N_10666);
nand U13660 (N_13660,N_10090,N_10490);
nand U13661 (N_13661,N_9083,N_11468);
xor U13662 (N_13662,N_11384,N_9512);
nor U13663 (N_13663,N_11791,N_11368);
or U13664 (N_13664,N_10779,N_10920);
nor U13665 (N_13665,N_9027,N_10656);
nand U13666 (N_13666,N_10058,N_9227);
nor U13667 (N_13667,N_9026,N_11013);
xor U13668 (N_13668,N_10287,N_10448);
nor U13669 (N_13669,N_10526,N_9525);
xnor U13670 (N_13670,N_10813,N_10848);
and U13671 (N_13671,N_9565,N_9858);
xnor U13672 (N_13672,N_11500,N_9411);
or U13673 (N_13673,N_10661,N_11917);
nand U13674 (N_13674,N_9012,N_11403);
nand U13675 (N_13675,N_10305,N_9287);
nor U13676 (N_13676,N_10476,N_9551);
and U13677 (N_13677,N_9251,N_11664);
or U13678 (N_13678,N_11233,N_9906);
nand U13679 (N_13679,N_10609,N_11601);
nand U13680 (N_13680,N_11371,N_11828);
nand U13681 (N_13681,N_9584,N_9383);
or U13682 (N_13682,N_10634,N_10958);
and U13683 (N_13683,N_9277,N_11909);
or U13684 (N_13684,N_10338,N_11312);
and U13685 (N_13685,N_9156,N_11950);
and U13686 (N_13686,N_11289,N_9626);
xor U13687 (N_13687,N_9812,N_11496);
nand U13688 (N_13688,N_9023,N_11352);
or U13689 (N_13689,N_10608,N_9253);
nand U13690 (N_13690,N_10041,N_11968);
nand U13691 (N_13691,N_11927,N_10766);
and U13692 (N_13692,N_11957,N_10106);
nor U13693 (N_13693,N_9107,N_9913);
or U13694 (N_13694,N_10642,N_10761);
nor U13695 (N_13695,N_10329,N_11008);
or U13696 (N_13696,N_9186,N_10834);
nand U13697 (N_13697,N_11273,N_9125);
nand U13698 (N_13698,N_11685,N_9507);
nand U13699 (N_13699,N_10155,N_10772);
xor U13700 (N_13700,N_9788,N_11105);
or U13701 (N_13701,N_9992,N_10241);
xnor U13702 (N_13702,N_11893,N_9864);
and U13703 (N_13703,N_10467,N_9802);
and U13704 (N_13704,N_10282,N_11449);
nand U13705 (N_13705,N_11176,N_11640);
nand U13706 (N_13706,N_10209,N_9734);
or U13707 (N_13707,N_10885,N_9747);
xnor U13708 (N_13708,N_10757,N_10607);
and U13709 (N_13709,N_9966,N_9746);
nand U13710 (N_13710,N_11022,N_10301);
xor U13711 (N_13711,N_11300,N_11846);
or U13712 (N_13712,N_9262,N_9692);
xnor U13713 (N_13713,N_9548,N_10920);
and U13714 (N_13714,N_10608,N_11525);
or U13715 (N_13715,N_11154,N_9082);
and U13716 (N_13716,N_10853,N_11707);
nor U13717 (N_13717,N_9395,N_10199);
nand U13718 (N_13718,N_10857,N_11689);
nand U13719 (N_13719,N_10951,N_11431);
nor U13720 (N_13720,N_10854,N_10813);
or U13721 (N_13721,N_11236,N_9100);
xor U13722 (N_13722,N_9899,N_9493);
xor U13723 (N_13723,N_9682,N_9918);
xor U13724 (N_13724,N_11398,N_9591);
nand U13725 (N_13725,N_10401,N_9378);
nand U13726 (N_13726,N_10666,N_9855);
xor U13727 (N_13727,N_10164,N_10230);
and U13728 (N_13728,N_10214,N_10917);
or U13729 (N_13729,N_11293,N_10013);
and U13730 (N_13730,N_9214,N_9490);
and U13731 (N_13731,N_11969,N_10670);
or U13732 (N_13732,N_11088,N_9070);
xnor U13733 (N_13733,N_10472,N_11470);
xor U13734 (N_13734,N_9082,N_9998);
nand U13735 (N_13735,N_9968,N_11455);
and U13736 (N_13736,N_10797,N_10364);
and U13737 (N_13737,N_11735,N_10375);
and U13738 (N_13738,N_9562,N_9075);
nor U13739 (N_13739,N_11989,N_11747);
or U13740 (N_13740,N_9969,N_10247);
nand U13741 (N_13741,N_9706,N_9551);
and U13742 (N_13742,N_11806,N_9483);
and U13743 (N_13743,N_10936,N_10060);
or U13744 (N_13744,N_11500,N_9049);
nand U13745 (N_13745,N_11735,N_10906);
nand U13746 (N_13746,N_9429,N_9358);
nor U13747 (N_13747,N_11581,N_11033);
xnor U13748 (N_13748,N_9142,N_11987);
xor U13749 (N_13749,N_9256,N_10163);
xor U13750 (N_13750,N_11497,N_10118);
xor U13751 (N_13751,N_9027,N_11923);
xnor U13752 (N_13752,N_9699,N_10403);
xnor U13753 (N_13753,N_10002,N_9400);
nand U13754 (N_13754,N_9273,N_10545);
or U13755 (N_13755,N_11026,N_9342);
nand U13756 (N_13756,N_10587,N_9877);
and U13757 (N_13757,N_10219,N_10276);
nand U13758 (N_13758,N_9139,N_11161);
and U13759 (N_13759,N_10845,N_11989);
xnor U13760 (N_13760,N_11052,N_9385);
nor U13761 (N_13761,N_9125,N_10739);
xnor U13762 (N_13762,N_9295,N_10172);
xor U13763 (N_13763,N_11139,N_11135);
xnor U13764 (N_13764,N_10463,N_11922);
nand U13765 (N_13765,N_9499,N_10473);
nor U13766 (N_13766,N_9066,N_9637);
nand U13767 (N_13767,N_11263,N_11133);
nor U13768 (N_13768,N_9326,N_9455);
nor U13769 (N_13769,N_10861,N_9483);
xor U13770 (N_13770,N_9908,N_9226);
and U13771 (N_13771,N_10367,N_9569);
xnor U13772 (N_13772,N_9711,N_9754);
or U13773 (N_13773,N_11882,N_10666);
nand U13774 (N_13774,N_9731,N_9775);
nand U13775 (N_13775,N_9894,N_10727);
xor U13776 (N_13776,N_9847,N_9075);
and U13777 (N_13777,N_11848,N_9421);
nand U13778 (N_13778,N_11437,N_9223);
nor U13779 (N_13779,N_9444,N_10953);
nand U13780 (N_13780,N_10129,N_9752);
and U13781 (N_13781,N_10391,N_10464);
nand U13782 (N_13782,N_11901,N_10223);
or U13783 (N_13783,N_9021,N_9614);
xnor U13784 (N_13784,N_11346,N_11092);
nor U13785 (N_13785,N_9160,N_11236);
xnor U13786 (N_13786,N_11450,N_10557);
xor U13787 (N_13787,N_11163,N_10842);
and U13788 (N_13788,N_10620,N_9501);
nand U13789 (N_13789,N_11330,N_11301);
nand U13790 (N_13790,N_11178,N_9028);
nand U13791 (N_13791,N_11471,N_9849);
nor U13792 (N_13792,N_9874,N_9218);
nor U13793 (N_13793,N_10709,N_10501);
nand U13794 (N_13794,N_9621,N_11607);
and U13795 (N_13795,N_10679,N_10511);
nand U13796 (N_13796,N_9499,N_11377);
or U13797 (N_13797,N_9750,N_10051);
and U13798 (N_13798,N_9058,N_10435);
and U13799 (N_13799,N_9548,N_10032);
and U13800 (N_13800,N_11210,N_9189);
nand U13801 (N_13801,N_10624,N_9613);
nand U13802 (N_13802,N_10741,N_11628);
or U13803 (N_13803,N_9929,N_11532);
and U13804 (N_13804,N_10558,N_9431);
or U13805 (N_13805,N_9436,N_11150);
or U13806 (N_13806,N_11524,N_9992);
and U13807 (N_13807,N_10051,N_10373);
nor U13808 (N_13808,N_10957,N_9308);
xor U13809 (N_13809,N_9530,N_9302);
and U13810 (N_13810,N_9974,N_9059);
xnor U13811 (N_13811,N_9116,N_9082);
or U13812 (N_13812,N_9226,N_9044);
xor U13813 (N_13813,N_11299,N_11082);
nor U13814 (N_13814,N_9360,N_11606);
nor U13815 (N_13815,N_10259,N_10786);
xnor U13816 (N_13816,N_11473,N_10298);
nand U13817 (N_13817,N_10104,N_10544);
and U13818 (N_13818,N_10958,N_10883);
or U13819 (N_13819,N_11040,N_11574);
and U13820 (N_13820,N_11771,N_10095);
nand U13821 (N_13821,N_10308,N_10691);
nand U13822 (N_13822,N_9808,N_10367);
and U13823 (N_13823,N_10969,N_9427);
and U13824 (N_13824,N_10348,N_11114);
nand U13825 (N_13825,N_11881,N_10639);
and U13826 (N_13826,N_11698,N_10802);
xor U13827 (N_13827,N_11475,N_11928);
nor U13828 (N_13828,N_9654,N_9541);
nor U13829 (N_13829,N_11669,N_11121);
and U13830 (N_13830,N_10199,N_11467);
xnor U13831 (N_13831,N_10545,N_11922);
nor U13832 (N_13832,N_10166,N_11904);
or U13833 (N_13833,N_11870,N_10981);
nor U13834 (N_13834,N_9761,N_11755);
nand U13835 (N_13835,N_9410,N_11149);
nand U13836 (N_13836,N_10513,N_10218);
xnor U13837 (N_13837,N_9329,N_11144);
nor U13838 (N_13838,N_11305,N_10520);
xnor U13839 (N_13839,N_9863,N_10366);
xor U13840 (N_13840,N_9039,N_11134);
nor U13841 (N_13841,N_9829,N_9002);
nor U13842 (N_13842,N_10801,N_10437);
and U13843 (N_13843,N_10028,N_10201);
and U13844 (N_13844,N_11968,N_10018);
and U13845 (N_13845,N_10838,N_9421);
xnor U13846 (N_13846,N_11206,N_11394);
nor U13847 (N_13847,N_9615,N_9867);
and U13848 (N_13848,N_9884,N_10510);
nand U13849 (N_13849,N_11846,N_10300);
or U13850 (N_13850,N_9707,N_10611);
and U13851 (N_13851,N_11434,N_10846);
nor U13852 (N_13852,N_10274,N_9755);
and U13853 (N_13853,N_11207,N_10433);
nor U13854 (N_13854,N_10271,N_11648);
nor U13855 (N_13855,N_10671,N_9471);
nor U13856 (N_13856,N_10253,N_11198);
or U13857 (N_13857,N_9078,N_11966);
nor U13858 (N_13858,N_9612,N_10095);
and U13859 (N_13859,N_11617,N_11946);
and U13860 (N_13860,N_9430,N_10230);
or U13861 (N_13861,N_10790,N_11717);
xor U13862 (N_13862,N_11019,N_9492);
or U13863 (N_13863,N_10434,N_11334);
and U13864 (N_13864,N_9393,N_10096);
nor U13865 (N_13865,N_10829,N_9916);
xnor U13866 (N_13866,N_10731,N_9736);
and U13867 (N_13867,N_11181,N_9928);
xnor U13868 (N_13868,N_10788,N_9374);
xor U13869 (N_13869,N_11632,N_9728);
or U13870 (N_13870,N_10671,N_11115);
or U13871 (N_13871,N_11682,N_11186);
nor U13872 (N_13872,N_9394,N_10761);
and U13873 (N_13873,N_9364,N_9165);
or U13874 (N_13874,N_10508,N_10921);
nand U13875 (N_13875,N_11955,N_11637);
or U13876 (N_13876,N_10092,N_10121);
and U13877 (N_13877,N_11105,N_10234);
or U13878 (N_13878,N_9116,N_11055);
nor U13879 (N_13879,N_9198,N_11445);
and U13880 (N_13880,N_10547,N_9457);
xnor U13881 (N_13881,N_11658,N_10772);
or U13882 (N_13882,N_9427,N_11939);
xor U13883 (N_13883,N_9576,N_11264);
nor U13884 (N_13884,N_10061,N_9813);
xnor U13885 (N_13885,N_9821,N_10762);
and U13886 (N_13886,N_11040,N_9701);
xor U13887 (N_13887,N_10278,N_10845);
and U13888 (N_13888,N_10752,N_11100);
or U13889 (N_13889,N_10470,N_10852);
xnor U13890 (N_13890,N_10774,N_10077);
and U13891 (N_13891,N_11710,N_9719);
xnor U13892 (N_13892,N_11327,N_11357);
nand U13893 (N_13893,N_11938,N_9027);
nand U13894 (N_13894,N_10289,N_9725);
or U13895 (N_13895,N_10282,N_9061);
nand U13896 (N_13896,N_10604,N_11281);
or U13897 (N_13897,N_9488,N_11869);
nor U13898 (N_13898,N_11293,N_9861);
xnor U13899 (N_13899,N_10942,N_10648);
nor U13900 (N_13900,N_11645,N_9284);
or U13901 (N_13901,N_10276,N_9827);
nand U13902 (N_13902,N_10071,N_10079);
nor U13903 (N_13903,N_10038,N_11766);
nand U13904 (N_13904,N_10752,N_11680);
or U13905 (N_13905,N_9940,N_10194);
nor U13906 (N_13906,N_11470,N_11036);
nand U13907 (N_13907,N_10608,N_11104);
nor U13908 (N_13908,N_11659,N_10126);
or U13909 (N_13909,N_10908,N_9701);
xnor U13910 (N_13910,N_9740,N_10144);
nand U13911 (N_13911,N_9484,N_10099);
or U13912 (N_13912,N_9231,N_10478);
and U13913 (N_13913,N_11249,N_10827);
nor U13914 (N_13914,N_11860,N_11915);
nor U13915 (N_13915,N_10928,N_10743);
nor U13916 (N_13916,N_9768,N_9974);
and U13917 (N_13917,N_11137,N_10649);
or U13918 (N_13918,N_10363,N_9564);
nand U13919 (N_13919,N_11779,N_9036);
and U13920 (N_13920,N_9007,N_9889);
nand U13921 (N_13921,N_10492,N_11640);
xor U13922 (N_13922,N_11361,N_10253);
nand U13923 (N_13923,N_9762,N_10064);
xnor U13924 (N_13924,N_10105,N_9275);
xor U13925 (N_13925,N_11693,N_9767);
or U13926 (N_13926,N_11371,N_10039);
nand U13927 (N_13927,N_10350,N_10767);
nor U13928 (N_13928,N_10205,N_10213);
or U13929 (N_13929,N_10607,N_10018);
nand U13930 (N_13930,N_9428,N_11719);
xnor U13931 (N_13931,N_11624,N_10326);
or U13932 (N_13932,N_11376,N_9980);
or U13933 (N_13933,N_9878,N_9057);
and U13934 (N_13934,N_9236,N_11363);
nor U13935 (N_13935,N_9540,N_9652);
nor U13936 (N_13936,N_10744,N_10435);
nand U13937 (N_13937,N_11303,N_10506);
nand U13938 (N_13938,N_9638,N_10035);
nor U13939 (N_13939,N_9060,N_10169);
and U13940 (N_13940,N_9985,N_11485);
or U13941 (N_13941,N_9679,N_9419);
or U13942 (N_13942,N_11918,N_9035);
nand U13943 (N_13943,N_9603,N_11958);
nor U13944 (N_13944,N_10248,N_10373);
and U13945 (N_13945,N_9087,N_9941);
nor U13946 (N_13946,N_11810,N_10983);
nand U13947 (N_13947,N_9727,N_11669);
xnor U13948 (N_13948,N_11228,N_11955);
or U13949 (N_13949,N_10555,N_11957);
nand U13950 (N_13950,N_10160,N_10747);
and U13951 (N_13951,N_10373,N_11348);
or U13952 (N_13952,N_10778,N_11629);
xnor U13953 (N_13953,N_11891,N_9944);
xor U13954 (N_13954,N_9004,N_10235);
nand U13955 (N_13955,N_9709,N_11972);
or U13956 (N_13956,N_10348,N_11593);
or U13957 (N_13957,N_11845,N_11071);
and U13958 (N_13958,N_11051,N_11311);
xor U13959 (N_13959,N_10842,N_9734);
and U13960 (N_13960,N_11683,N_11158);
or U13961 (N_13961,N_10837,N_9538);
or U13962 (N_13962,N_9191,N_10965);
nor U13963 (N_13963,N_11788,N_10074);
xor U13964 (N_13964,N_10247,N_9278);
xnor U13965 (N_13965,N_11883,N_10741);
xor U13966 (N_13966,N_9996,N_9946);
nor U13967 (N_13967,N_10153,N_9475);
or U13968 (N_13968,N_11587,N_10701);
nand U13969 (N_13969,N_10017,N_9961);
xor U13970 (N_13970,N_9533,N_9522);
nand U13971 (N_13971,N_11860,N_11105);
and U13972 (N_13972,N_10191,N_11176);
nand U13973 (N_13973,N_10970,N_10828);
or U13974 (N_13974,N_9508,N_11253);
nand U13975 (N_13975,N_11350,N_9128);
nor U13976 (N_13976,N_11332,N_9858);
and U13977 (N_13977,N_11859,N_10343);
nor U13978 (N_13978,N_11127,N_10417);
and U13979 (N_13979,N_9307,N_9291);
nand U13980 (N_13980,N_9053,N_9906);
and U13981 (N_13981,N_11711,N_9548);
or U13982 (N_13982,N_10247,N_9072);
xnor U13983 (N_13983,N_9722,N_9068);
or U13984 (N_13984,N_10986,N_11970);
and U13985 (N_13985,N_10457,N_9621);
and U13986 (N_13986,N_9706,N_9269);
nand U13987 (N_13987,N_9791,N_9451);
nand U13988 (N_13988,N_10518,N_11808);
and U13989 (N_13989,N_10417,N_10199);
xnor U13990 (N_13990,N_11080,N_9042);
or U13991 (N_13991,N_9949,N_9857);
or U13992 (N_13992,N_9451,N_10231);
xor U13993 (N_13993,N_11232,N_10595);
or U13994 (N_13994,N_10374,N_9660);
xnor U13995 (N_13995,N_9948,N_10349);
nor U13996 (N_13996,N_11701,N_11229);
nor U13997 (N_13997,N_9957,N_10626);
nor U13998 (N_13998,N_11247,N_11242);
nand U13999 (N_13999,N_9702,N_9133);
and U14000 (N_14000,N_10675,N_10232);
nor U14001 (N_14001,N_9836,N_10436);
nand U14002 (N_14002,N_11893,N_10057);
nand U14003 (N_14003,N_9031,N_10993);
nor U14004 (N_14004,N_11488,N_9382);
xor U14005 (N_14005,N_9704,N_11757);
nor U14006 (N_14006,N_9891,N_9907);
nand U14007 (N_14007,N_10975,N_11682);
nand U14008 (N_14008,N_10536,N_9773);
or U14009 (N_14009,N_9884,N_10643);
or U14010 (N_14010,N_9075,N_11414);
xor U14011 (N_14011,N_10884,N_9598);
nor U14012 (N_14012,N_11412,N_11990);
nand U14013 (N_14013,N_10794,N_9578);
and U14014 (N_14014,N_11293,N_10104);
xor U14015 (N_14015,N_10553,N_9347);
nand U14016 (N_14016,N_10489,N_9626);
or U14017 (N_14017,N_9864,N_11988);
nand U14018 (N_14018,N_10607,N_11690);
xor U14019 (N_14019,N_10395,N_11790);
nand U14020 (N_14020,N_10235,N_11900);
and U14021 (N_14021,N_10254,N_9500);
nor U14022 (N_14022,N_9502,N_9476);
and U14023 (N_14023,N_9124,N_11893);
nand U14024 (N_14024,N_10068,N_10177);
nor U14025 (N_14025,N_11705,N_9681);
or U14026 (N_14026,N_11421,N_10343);
nand U14027 (N_14027,N_9895,N_10200);
nand U14028 (N_14028,N_11850,N_11500);
nand U14029 (N_14029,N_11341,N_9662);
nor U14030 (N_14030,N_9997,N_9625);
or U14031 (N_14031,N_9932,N_9656);
or U14032 (N_14032,N_10827,N_9792);
or U14033 (N_14033,N_9312,N_10047);
nor U14034 (N_14034,N_11412,N_10334);
nor U14035 (N_14035,N_10831,N_10465);
or U14036 (N_14036,N_11450,N_9687);
and U14037 (N_14037,N_9032,N_10254);
or U14038 (N_14038,N_10431,N_11771);
and U14039 (N_14039,N_10978,N_11216);
or U14040 (N_14040,N_9522,N_10348);
nand U14041 (N_14041,N_11245,N_11559);
xor U14042 (N_14042,N_11883,N_10158);
nor U14043 (N_14043,N_10553,N_11473);
and U14044 (N_14044,N_10106,N_10735);
and U14045 (N_14045,N_10995,N_9610);
or U14046 (N_14046,N_10271,N_10785);
or U14047 (N_14047,N_11382,N_10873);
nand U14048 (N_14048,N_9014,N_9392);
nand U14049 (N_14049,N_11140,N_11889);
xnor U14050 (N_14050,N_11244,N_10072);
and U14051 (N_14051,N_10560,N_11837);
nor U14052 (N_14052,N_10091,N_10219);
nand U14053 (N_14053,N_9765,N_9559);
or U14054 (N_14054,N_10691,N_9648);
and U14055 (N_14055,N_11574,N_11055);
xnor U14056 (N_14056,N_10871,N_10200);
or U14057 (N_14057,N_10728,N_11784);
nor U14058 (N_14058,N_10335,N_9258);
xor U14059 (N_14059,N_10682,N_9809);
or U14060 (N_14060,N_9538,N_10916);
nor U14061 (N_14061,N_10972,N_10519);
nand U14062 (N_14062,N_10791,N_11161);
nand U14063 (N_14063,N_10558,N_10051);
xor U14064 (N_14064,N_9657,N_11218);
or U14065 (N_14065,N_9256,N_11196);
nand U14066 (N_14066,N_9860,N_9129);
or U14067 (N_14067,N_9868,N_11837);
xor U14068 (N_14068,N_9029,N_10888);
xor U14069 (N_14069,N_11182,N_10671);
or U14070 (N_14070,N_11287,N_10562);
and U14071 (N_14071,N_9956,N_11374);
nand U14072 (N_14072,N_9962,N_11918);
or U14073 (N_14073,N_11213,N_10197);
nor U14074 (N_14074,N_10793,N_10437);
or U14075 (N_14075,N_11119,N_9587);
nor U14076 (N_14076,N_10231,N_11643);
nand U14077 (N_14077,N_9111,N_9091);
nor U14078 (N_14078,N_9421,N_11944);
nand U14079 (N_14079,N_9027,N_10234);
or U14080 (N_14080,N_11807,N_9514);
nand U14081 (N_14081,N_10429,N_9624);
nor U14082 (N_14082,N_9923,N_11810);
and U14083 (N_14083,N_10555,N_11671);
nor U14084 (N_14084,N_11083,N_11072);
nor U14085 (N_14085,N_11320,N_9374);
or U14086 (N_14086,N_11849,N_11201);
or U14087 (N_14087,N_11517,N_9002);
or U14088 (N_14088,N_11856,N_9991);
or U14089 (N_14089,N_10397,N_9632);
or U14090 (N_14090,N_11107,N_11974);
and U14091 (N_14091,N_11807,N_10255);
nor U14092 (N_14092,N_10958,N_10408);
and U14093 (N_14093,N_9295,N_10390);
xnor U14094 (N_14094,N_11493,N_10039);
or U14095 (N_14095,N_10954,N_9681);
nand U14096 (N_14096,N_9313,N_10235);
or U14097 (N_14097,N_9341,N_9045);
and U14098 (N_14098,N_11406,N_10953);
xnor U14099 (N_14099,N_10706,N_11074);
nand U14100 (N_14100,N_11932,N_9750);
nand U14101 (N_14101,N_10452,N_10480);
nor U14102 (N_14102,N_11396,N_10230);
or U14103 (N_14103,N_10142,N_9441);
nor U14104 (N_14104,N_10513,N_10794);
or U14105 (N_14105,N_10087,N_11058);
nand U14106 (N_14106,N_11176,N_9020);
and U14107 (N_14107,N_9081,N_10632);
nand U14108 (N_14108,N_9644,N_9488);
nand U14109 (N_14109,N_9926,N_9305);
or U14110 (N_14110,N_9358,N_9940);
xnor U14111 (N_14111,N_10845,N_11625);
nor U14112 (N_14112,N_9499,N_9765);
or U14113 (N_14113,N_9377,N_11079);
xor U14114 (N_14114,N_10671,N_10419);
nor U14115 (N_14115,N_9481,N_10318);
xnor U14116 (N_14116,N_10480,N_10968);
nand U14117 (N_14117,N_11219,N_9934);
nor U14118 (N_14118,N_9159,N_9674);
nor U14119 (N_14119,N_10510,N_10156);
xnor U14120 (N_14120,N_9191,N_10090);
xnor U14121 (N_14121,N_11611,N_9128);
or U14122 (N_14122,N_9534,N_11755);
and U14123 (N_14123,N_11516,N_11276);
xor U14124 (N_14124,N_10621,N_9578);
and U14125 (N_14125,N_10975,N_10616);
nor U14126 (N_14126,N_10101,N_9194);
or U14127 (N_14127,N_11743,N_10786);
or U14128 (N_14128,N_11826,N_10412);
nor U14129 (N_14129,N_11681,N_9264);
nand U14130 (N_14130,N_10272,N_10811);
and U14131 (N_14131,N_10440,N_10098);
nor U14132 (N_14132,N_9411,N_9030);
nand U14133 (N_14133,N_11262,N_11385);
nand U14134 (N_14134,N_9644,N_9478);
or U14135 (N_14135,N_10084,N_10455);
and U14136 (N_14136,N_9415,N_10835);
or U14137 (N_14137,N_10926,N_10400);
nand U14138 (N_14138,N_9629,N_10274);
nand U14139 (N_14139,N_11246,N_10576);
or U14140 (N_14140,N_10788,N_10073);
nand U14141 (N_14141,N_11094,N_11333);
nor U14142 (N_14142,N_10071,N_10592);
and U14143 (N_14143,N_10393,N_9667);
nor U14144 (N_14144,N_10995,N_9005);
nor U14145 (N_14145,N_10567,N_9475);
or U14146 (N_14146,N_11793,N_10248);
or U14147 (N_14147,N_9939,N_9024);
xnor U14148 (N_14148,N_9916,N_11829);
or U14149 (N_14149,N_10638,N_10849);
xnor U14150 (N_14150,N_10313,N_9939);
or U14151 (N_14151,N_10425,N_11584);
nor U14152 (N_14152,N_10110,N_11442);
or U14153 (N_14153,N_11314,N_10959);
nand U14154 (N_14154,N_11328,N_10706);
and U14155 (N_14155,N_11590,N_10371);
xnor U14156 (N_14156,N_11061,N_11752);
nor U14157 (N_14157,N_9299,N_9795);
or U14158 (N_14158,N_9276,N_10272);
and U14159 (N_14159,N_11497,N_10938);
or U14160 (N_14160,N_10538,N_11228);
and U14161 (N_14161,N_11971,N_10433);
nand U14162 (N_14162,N_10747,N_11737);
nand U14163 (N_14163,N_11034,N_10932);
nor U14164 (N_14164,N_9960,N_9951);
nor U14165 (N_14165,N_9963,N_9196);
xor U14166 (N_14166,N_9109,N_9900);
and U14167 (N_14167,N_10963,N_11439);
or U14168 (N_14168,N_11977,N_10636);
nand U14169 (N_14169,N_9596,N_11872);
and U14170 (N_14170,N_11665,N_9427);
and U14171 (N_14171,N_11340,N_9853);
or U14172 (N_14172,N_9770,N_10207);
nor U14173 (N_14173,N_11605,N_11074);
xnor U14174 (N_14174,N_9659,N_11407);
nand U14175 (N_14175,N_9599,N_10291);
xor U14176 (N_14176,N_11797,N_10785);
and U14177 (N_14177,N_11584,N_9909);
and U14178 (N_14178,N_11428,N_9530);
xnor U14179 (N_14179,N_11895,N_10713);
nand U14180 (N_14180,N_10020,N_10130);
nor U14181 (N_14181,N_11590,N_9977);
nand U14182 (N_14182,N_10731,N_11922);
or U14183 (N_14183,N_9826,N_10016);
or U14184 (N_14184,N_9023,N_10465);
nand U14185 (N_14185,N_9303,N_9215);
xnor U14186 (N_14186,N_11162,N_10464);
and U14187 (N_14187,N_11740,N_10751);
nor U14188 (N_14188,N_10437,N_11095);
and U14189 (N_14189,N_11525,N_11090);
or U14190 (N_14190,N_9160,N_11919);
and U14191 (N_14191,N_11612,N_9181);
xnor U14192 (N_14192,N_11963,N_9133);
or U14193 (N_14193,N_9285,N_11509);
nand U14194 (N_14194,N_11740,N_10906);
and U14195 (N_14195,N_10294,N_10755);
nand U14196 (N_14196,N_10201,N_9563);
and U14197 (N_14197,N_10245,N_10791);
xor U14198 (N_14198,N_11204,N_9745);
and U14199 (N_14199,N_10233,N_9692);
nand U14200 (N_14200,N_9611,N_9383);
nand U14201 (N_14201,N_11632,N_10438);
nand U14202 (N_14202,N_10205,N_9996);
xor U14203 (N_14203,N_9568,N_9664);
xnor U14204 (N_14204,N_10309,N_10020);
or U14205 (N_14205,N_10068,N_11746);
xor U14206 (N_14206,N_11218,N_9005);
or U14207 (N_14207,N_10207,N_10867);
and U14208 (N_14208,N_11412,N_10271);
or U14209 (N_14209,N_9101,N_11573);
or U14210 (N_14210,N_9166,N_10021);
nand U14211 (N_14211,N_11956,N_11683);
xor U14212 (N_14212,N_10860,N_9316);
nor U14213 (N_14213,N_11991,N_9825);
or U14214 (N_14214,N_9893,N_11016);
nand U14215 (N_14215,N_11476,N_11337);
or U14216 (N_14216,N_9709,N_11581);
and U14217 (N_14217,N_11976,N_11506);
nand U14218 (N_14218,N_10988,N_11214);
xnor U14219 (N_14219,N_11580,N_10056);
xnor U14220 (N_14220,N_9015,N_11343);
nor U14221 (N_14221,N_10083,N_11380);
and U14222 (N_14222,N_10473,N_10710);
or U14223 (N_14223,N_10547,N_11107);
nand U14224 (N_14224,N_9612,N_11754);
xnor U14225 (N_14225,N_10789,N_10189);
nor U14226 (N_14226,N_9592,N_11144);
nor U14227 (N_14227,N_11508,N_10459);
nor U14228 (N_14228,N_9224,N_9184);
and U14229 (N_14229,N_9687,N_11007);
or U14230 (N_14230,N_11796,N_11945);
or U14231 (N_14231,N_11343,N_10067);
nand U14232 (N_14232,N_9476,N_9380);
xor U14233 (N_14233,N_10384,N_11421);
and U14234 (N_14234,N_10315,N_9636);
nor U14235 (N_14235,N_10471,N_10009);
xnor U14236 (N_14236,N_10084,N_10359);
or U14237 (N_14237,N_9567,N_11429);
nor U14238 (N_14238,N_9107,N_11741);
xor U14239 (N_14239,N_10249,N_9504);
and U14240 (N_14240,N_10275,N_11259);
nand U14241 (N_14241,N_11291,N_11290);
xor U14242 (N_14242,N_9026,N_9668);
nand U14243 (N_14243,N_9455,N_11057);
and U14244 (N_14244,N_11318,N_11351);
nor U14245 (N_14245,N_10496,N_11499);
and U14246 (N_14246,N_10685,N_10119);
xnor U14247 (N_14247,N_9405,N_10312);
or U14248 (N_14248,N_9133,N_11942);
and U14249 (N_14249,N_11506,N_9684);
xnor U14250 (N_14250,N_9352,N_9163);
nor U14251 (N_14251,N_9701,N_10550);
nand U14252 (N_14252,N_11213,N_9235);
xnor U14253 (N_14253,N_10307,N_11530);
nor U14254 (N_14254,N_9447,N_11708);
or U14255 (N_14255,N_11359,N_9284);
nand U14256 (N_14256,N_11088,N_10881);
nand U14257 (N_14257,N_11533,N_11026);
or U14258 (N_14258,N_9452,N_10788);
nor U14259 (N_14259,N_10427,N_10766);
nor U14260 (N_14260,N_11494,N_10753);
and U14261 (N_14261,N_11982,N_11421);
nor U14262 (N_14262,N_9768,N_9536);
and U14263 (N_14263,N_9854,N_11067);
nor U14264 (N_14264,N_10844,N_9331);
nor U14265 (N_14265,N_11582,N_9647);
nand U14266 (N_14266,N_10676,N_11776);
xor U14267 (N_14267,N_10519,N_9118);
and U14268 (N_14268,N_10068,N_9906);
nand U14269 (N_14269,N_10326,N_11440);
xor U14270 (N_14270,N_10421,N_9849);
xor U14271 (N_14271,N_11652,N_11492);
xor U14272 (N_14272,N_10783,N_10013);
nand U14273 (N_14273,N_9817,N_11251);
nand U14274 (N_14274,N_9374,N_9141);
and U14275 (N_14275,N_11230,N_10069);
or U14276 (N_14276,N_11406,N_10212);
nor U14277 (N_14277,N_11698,N_11259);
nand U14278 (N_14278,N_10175,N_11665);
nor U14279 (N_14279,N_10994,N_10387);
nand U14280 (N_14280,N_11603,N_10976);
xor U14281 (N_14281,N_11560,N_11367);
nor U14282 (N_14282,N_11328,N_10887);
or U14283 (N_14283,N_10011,N_9531);
nand U14284 (N_14284,N_10164,N_11092);
or U14285 (N_14285,N_9914,N_10533);
xor U14286 (N_14286,N_9329,N_11279);
nor U14287 (N_14287,N_9411,N_11472);
nor U14288 (N_14288,N_9204,N_10509);
nand U14289 (N_14289,N_11732,N_10670);
nor U14290 (N_14290,N_9210,N_9995);
or U14291 (N_14291,N_10080,N_11722);
and U14292 (N_14292,N_9728,N_9039);
or U14293 (N_14293,N_9816,N_11195);
nand U14294 (N_14294,N_9373,N_10962);
and U14295 (N_14295,N_10435,N_9344);
nor U14296 (N_14296,N_9180,N_10547);
or U14297 (N_14297,N_9897,N_11053);
or U14298 (N_14298,N_9635,N_11015);
xor U14299 (N_14299,N_10979,N_9959);
xor U14300 (N_14300,N_10571,N_10715);
nor U14301 (N_14301,N_9069,N_9176);
xor U14302 (N_14302,N_11816,N_11767);
or U14303 (N_14303,N_10220,N_9718);
xor U14304 (N_14304,N_9601,N_9332);
nor U14305 (N_14305,N_11236,N_11857);
or U14306 (N_14306,N_10221,N_9224);
nand U14307 (N_14307,N_9979,N_9658);
and U14308 (N_14308,N_9612,N_9216);
nor U14309 (N_14309,N_10094,N_10166);
or U14310 (N_14310,N_11036,N_9772);
nor U14311 (N_14311,N_11184,N_11527);
xnor U14312 (N_14312,N_10174,N_11416);
xor U14313 (N_14313,N_10389,N_10918);
nand U14314 (N_14314,N_11496,N_10711);
xor U14315 (N_14315,N_9254,N_11875);
nand U14316 (N_14316,N_11252,N_11051);
and U14317 (N_14317,N_9932,N_11913);
nand U14318 (N_14318,N_9411,N_11614);
nand U14319 (N_14319,N_10353,N_10899);
and U14320 (N_14320,N_11460,N_9330);
and U14321 (N_14321,N_11135,N_9668);
or U14322 (N_14322,N_11229,N_11335);
nand U14323 (N_14323,N_10094,N_10031);
or U14324 (N_14324,N_10444,N_10767);
xor U14325 (N_14325,N_9078,N_11530);
nand U14326 (N_14326,N_11001,N_9418);
nor U14327 (N_14327,N_11281,N_10107);
xnor U14328 (N_14328,N_11707,N_11879);
nor U14329 (N_14329,N_11986,N_9382);
nand U14330 (N_14330,N_10448,N_9190);
nor U14331 (N_14331,N_11912,N_9108);
or U14332 (N_14332,N_9691,N_11219);
and U14333 (N_14333,N_9997,N_11710);
nor U14334 (N_14334,N_9637,N_11581);
nor U14335 (N_14335,N_9416,N_10541);
xor U14336 (N_14336,N_10924,N_9133);
or U14337 (N_14337,N_10374,N_9265);
or U14338 (N_14338,N_9252,N_11505);
or U14339 (N_14339,N_11341,N_9024);
and U14340 (N_14340,N_9881,N_10253);
nand U14341 (N_14341,N_9467,N_10973);
and U14342 (N_14342,N_11964,N_10736);
and U14343 (N_14343,N_9000,N_10358);
or U14344 (N_14344,N_9533,N_11121);
xnor U14345 (N_14345,N_11357,N_9359);
or U14346 (N_14346,N_10554,N_10818);
nand U14347 (N_14347,N_10590,N_11391);
or U14348 (N_14348,N_11695,N_11106);
xnor U14349 (N_14349,N_9883,N_10292);
or U14350 (N_14350,N_11147,N_10822);
and U14351 (N_14351,N_9184,N_9220);
and U14352 (N_14352,N_10364,N_9846);
nand U14353 (N_14353,N_9456,N_10676);
nand U14354 (N_14354,N_10810,N_9541);
or U14355 (N_14355,N_11954,N_9968);
nand U14356 (N_14356,N_11345,N_9855);
and U14357 (N_14357,N_9231,N_9983);
xnor U14358 (N_14358,N_9529,N_9990);
nor U14359 (N_14359,N_11155,N_11696);
nor U14360 (N_14360,N_11549,N_10636);
xnor U14361 (N_14361,N_9360,N_9265);
nand U14362 (N_14362,N_11078,N_10690);
or U14363 (N_14363,N_9160,N_11708);
or U14364 (N_14364,N_9573,N_10934);
or U14365 (N_14365,N_11205,N_10225);
and U14366 (N_14366,N_10281,N_10750);
nand U14367 (N_14367,N_11409,N_10239);
or U14368 (N_14368,N_10677,N_10858);
nor U14369 (N_14369,N_10752,N_10615);
nor U14370 (N_14370,N_9922,N_11215);
and U14371 (N_14371,N_10936,N_11844);
or U14372 (N_14372,N_10058,N_9525);
and U14373 (N_14373,N_11881,N_9493);
xor U14374 (N_14374,N_9951,N_10278);
nor U14375 (N_14375,N_11401,N_11112);
and U14376 (N_14376,N_11342,N_11984);
or U14377 (N_14377,N_9446,N_10425);
nand U14378 (N_14378,N_9332,N_10047);
and U14379 (N_14379,N_10690,N_11508);
and U14380 (N_14380,N_11766,N_9991);
xnor U14381 (N_14381,N_11439,N_9731);
or U14382 (N_14382,N_11127,N_10920);
and U14383 (N_14383,N_9889,N_11389);
and U14384 (N_14384,N_11949,N_11769);
nand U14385 (N_14385,N_9377,N_11749);
xnor U14386 (N_14386,N_10448,N_11925);
and U14387 (N_14387,N_10980,N_11727);
xor U14388 (N_14388,N_11266,N_10970);
xor U14389 (N_14389,N_9565,N_11648);
and U14390 (N_14390,N_10746,N_11110);
and U14391 (N_14391,N_11276,N_10015);
or U14392 (N_14392,N_9903,N_10191);
and U14393 (N_14393,N_11551,N_9055);
xor U14394 (N_14394,N_9481,N_11678);
nor U14395 (N_14395,N_9392,N_10414);
nand U14396 (N_14396,N_9159,N_10276);
or U14397 (N_14397,N_11301,N_11094);
nand U14398 (N_14398,N_10431,N_10032);
nor U14399 (N_14399,N_10915,N_11019);
nand U14400 (N_14400,N_11323,N_11877);
or U14401 (N_14401,N_11619,N_11693);
xor U14402 (N_14402,N_11593,N_10008);
nand U14403 (N_14403,N_9422,N_10272);
nor U14404 (N_14404,N_9583,N_11792);
xnor U14405 (N_14405,N_9495,N_10119);
nand U14406 (N_14406,N_9242,N_9781);
nor U14407 (N_14407,N_11633,N_11784);
xnor U14408 (N_14408,N_9945,N_11885);
nor U14409 (N_14409,N_9107,N_10087);
nor U14410 (N_14410,N_10328,N_9028);
nor U14411 (N_14411,N_9591,N_9754);
or U14412 (N_14412,N_11356,N_10596);
and U14413 (N_14413,N_9996,N_11152);
nor U14414 (N_14414,N_9408,N_11995);
or U14415 (N_14415,N_11197,N_10255);
or U14416 (N_14416,N_10664,N_10759);
or U14417 (N_14417,N_9211,N_9981);
and U14418 (N_14418,N_11353,N_9519);
nor U14419 (N_14419,N_10625,N_10822);
and U14420 (N_14420,N_10854,N_11985);
nor U14421 (N_14421,N_9856,N_10025);
xor U14422 (N_14422,N_9835,N_11030);
nor U14423 (N_14423,N_10339,N_11268);
or U14424 (N_14424,N_9822,N_11550);
or U14425 (N_14425,N_10616,N_9146);
or U14426 (N_14426,N_9561,N_9975);
nor U14427 (N_14427,N_10810,N_11853);
and U14428 (N_14428,N_10696,N_9019);
xor U14429 (N_14429,N_11252,N_9059);
xnor U14430 (N_14430,N_9764,N_10590);
nor U14431 (N_14431,N_9961,N_10688);
and U14432 (N_14432,N_10874,N_9193);
and U14433 (N_14433,N_11999,N_10216);
xnor U14434 (N_14434,N_11396,N_9354);
xnor U14435 (N_14435,N_10572,N_9346);
and U14436 (N_14436,N_10728,N_11583);
or U14437 (N_14437,N_10688,N_9269);
and U14438 (N_14438,N_11982,N_11291);
nand U14439 (N_14439,N_10627,N_10557);
and U14440 (N_14440,N_10628,N_11132);
nand U14441 (N_14441,N_11952,N_9786);
nand U14442 (N_14442,N_10943,N_11822);
or U14443 (N_14443,N_9096,N_9629);
and U14444 (N_14444,N_10457,N_9905);
xor U14445 (N_14445,N_10473,N_10931);
nand U14446 (N_14446,N_11227,N_10733);
xor U14447 (N_14447,N_9954,N_9361);
nand U14448 (N_14448,N_11116,N_11128);
or U14449 (N_14449,N_10181,N_11069);
nor U14450 (N_14450,N_11577,N_9999);
nor U14451 (N_14451,N_10421,N_10089);
or U14452 (N_14452,N_9599,N_11790);
or U14453 (N_14453,N_11215,N_10259);
or U14454 (N_14454,N_11899,N_10136);
or U14455 (N_14455,N_11075,N_11354);
or U14456 (N_14456,N_11669,N_10962);
and U14457 (N_14457,N_9774,N_11827);
nor U14458 (N_14458,N_11218,N_10695);
nand U14459 (N_14459,N_10165,N_10221);
nand U14460 (N_14460,N_11894,N_11431);
xnor U14461 (N_14461,N_10236,N_9689);
nand U14462 (N_14462,N_11609,N_10684);
and U14463 (N_14463,N_10940,N_11928);
nor U14464 (N_14464,N_11218,N_9119);
xnor U14465 (N_14465,N_11329,N_9577);
nor U14466 (N_14466,N_9164,N_10356);
nor U14467 (N_14467,N_11882,N_9466);
nand U14468 (N_14468,N_9241,N_11426);
nand U14469 (N_14469,N_10442,N_10803);
nor U14470 (N_14470,N_10937,N_11038);
or U14471 (N_14471,N_9894,N_11357);
or U14472 (N_14472,N_10295,N_10649);
xor U14473 (N_14473,N_9848,N_10818);
xor U14474 (N_14474,N_9961,N_11003);
and U14475 (N_14475,N_11451,N_9546);
nand U14476 (N_14476,N_11064,N_10143);
nand U14477 (N_14477,N_10646,N_10355);
xnor U14478 (N_14478,N_11050,N_9529);
or U14479 (N_14479,N_10795,N_10195);
or U14480 (N_14480,N_9241,N_11154);
nor U14481 (N_14481,N_10187,N_10313);
and U14482 (N_14482,N_10883,N_9365);
xor U14483 (N_14483,N_10115,N_9490);
and U14484 (N_14484,N_9886,N_9570);
nor U14485 (N_14485,N_11541,N_10539);
xnor U14486 (N_14486,N_9407,N_9935);
nand U14487 (N_14487,N_9134,N_10227);
and U14488 (N_14488,N_9138,N_10362);
and U14489 (N_14489,N_9531,N_9614);
nor U14490 (N_14490,N_11734,N_10411);
nor U14491 (N_14491,N_9665,N_9437);
and U14492 (N_14492,N_10579,N_10668);
or U14493 (N_14493,N_10256,N_10878);
and U14494 (N_14494,N_9189,N_10707);
or U14495 (N_14495,N_11061,N_11237);
nand U14496 (N_14496,N_9621,N_11473);
or U14497 (N_14497,N_10245,N_10288);
nand U14498 (N_14498,N_10698,N_9892);
nor U14499 (N_14499,N_11197,N_10620);
nand U14500 (N_14500,N_10119,N_11941);
xor U14501 (N_14501,N_9716,N_10084);
nand U14502 (N_14502,N_9552,N_11803);
xnor U14503 (N_14503,N_11788,N_10044);
xnor U14504 (N_14504,N_10502,N_11057);
nor U14505 (N_14505,N_9560,N_9796);
nor U14506 (N_14506,N_11632,N_9256);
and U14507 (N_14507,N_11272,N_11819);
nand U14508 (N_14508,N_11822,N_9638);
and U14509 (N_14509,N_9706,N_11898);
and U14510 (N_14510,N_11415,N_9898);
and U14511 (N_14511,N_11720,N_10524);
xor U14512 (N_14512,N_9511,N_9740);
or U14513 (N_14513,N_9028,N_10512);
xnor U14514 (N_14514,N_11669,N_10321);
or U14515 (N_14515,N_10058,N_11281);
and U14516 (N_14516,N_9747,N_10725);
nor U14517 (N_14517,N_10812,N_9951);
or U14518 (N_14518,N_9760,N_9202);
xnor U14519 (N_14519,N_9451,N_11693);
and U14520 (N_14520,N_10416,N_10828);
nor U14521 (N_14521,N_10532,N_10921);
nand U14522 (N_14522,N_10176,N_9712);
xor U14523 (N_14523,N_9501,N_11475);
or U14524 (N_14524,N_11884,N_9959);
nand U14525 (N_14525,N_10747,N_10972);
or U14526 (N_14526,N_11129,N_11307);
xor U14527 (N_14527,N_10805,N_11403);
nand U14528 (N_14528,N_9765,N_10923);
nor U14529 (N_14529,N_10101,N_11097);
nand U14530 (N_14530,N_11756,N_9738);
xnor U14531 (N_14531,N_11292,N_9480);
xnor U14532 (N_14532,N_11648,N_11989);
nand U14533 (N_14533,N_9622,N_10097);
xnor U14534 (N_14534,N_11502,N_10798);
and U14535 (N_14535,N_11633,N_9081);
xnor U14536 (N_14536,N_11480,N_10337);
xnor U14537 (N_14537,N_11725,N_9050);
nand U14538 (N_14538,N_10075,N_10825);
and U14539 (N_14539,N_10600,N_10954);
xor U14540 (N_14540,N_9134,N_10057);
and U14541 (N_14541,N_11747,N_9153);
xor U14542 (N_14542,N_11252,N_10583);
and U14543 (N_14543,N_10651,N_9080);
or U14544 (N_14544,N_10347,N_9571);
xnor U14545 (N_14545,N_10060,N_11229);
and U14546 (N_14546,N_11795,N_11283);
or U14547 (N_14547,N_10701,N_10239);
nor U14548 (N_14548,N_11628,N_9254);
nor U14549 (N_14549,N_11294,N_9706);
or U14550 (N_14550,N_9693,N_9023);
or U14551 (N_14551,N_10353,N_11747);
or U14552 (N_14552,N_10797,N_9978);
nor U14553 (N_14553,N_11970,N_10465);
xnor U14554 (N_14554,N_11748,N_10187);
nand U14555 (N_14555,N_10074,N_10072);
or U14556 (N_14556,N_10248,N_11382);
and U14557 (N_14557,N_11692,N_10762);
and U14558 (N_14558,N_9174,N_9355);
nor U14559 (N_14559,N_10336,N_11264);
nor U14560 (N_14560,N_11396,N_9052);
nand U14561 (N_14561,N_10259,N_10783);
and U14562 (N_14562,N_11715,N_10140);
and U14563 (N_14563,N_10943,N_10485);
nor U14564 (N_14564,N_9108,N_9967);
or U14565 (N_14565,N_11625,N_9635);
xor U14566 (N_14566,N_11837,N_10200);
xnor U14567 (N_14567,N_11492,N_11774);
and U14568 (N_14568,N_10389,N_11908);
or U14569 (N_14569,N_9957,N_10115);
nand U14570 (N_14570,N_9973,N_11004);
xor U14571 (N_14571,N_9336,N_9596);
nor U14572 (N_14572,N_9047,N_10394);
nand U14573 (N_14573,N_9653,N_11066);
and U14574 (N_14574,N_11112,N_10783);
and U14575 (N_14575,N_11706,N_10158);
and U14576 (N_14576,N_9451,N_10648);
and U14577 (N_14577,N_10761,N_10091);
nor U14578 (N_14578,N_11944,N_9838);
xnor U14579 (N_14579,N_10653,N_9319);
nand U14580 (N_14580,N_11671,N_9361);
or U14581 (N_14581,N_11463,N_9587);
xnor U14582 (N_14582,N_11765,N_9424);
nand U14583 (N_14583,N_11208,N_10581);
and U14584 (N_14584,N_9783,N_11010);
or U14585 (N_14585,N_10635,N_9241);
or U14586 (N_14586,N_10879,N_11544);
xor U14587 (N_14587,N_11948,N_9136);
and U14588 (N_14588,N_10992,N_11921);
nand U14589 (N_14589,N_11563,N_10037);
and U14590 (N_14590,N_9803,N_10705);
and U14591 (N_14591,N_11707,N_10317);
or U14592 (N_14592,N_9928,N_9323);
or U14593 (N_14593,N_11803,N_9595);
xnor U14594 (N_14594,N_11908,N_9937);
nor U14595 (N_14595,N_9706,N_11880);
or U14596 (N_14596,N_11758,N_11021);
xor U14597 (N_14597,N_11145,N_9276);
nand U14598 (N_14598,N_11076,N_11444);
xnor U14599 (N_14599,N_9352,N_11949);
and U14600 (N_14600,N_9247,N_10596);
and U14601 (N_14601,N_9154,N_10193);
nand U14602 (N_14602,N_11201,N_10239);
nand U14603 (N_14603,N_11241,N_10626);
and U14604 (N_14604,N_11182,N_11798);
xor U14605 (N_14605,N_9305,N_10049);
and U14606 (N_14606,N_10994,N_9794);
nand U14607 (N_14607,N_11994,N_11090);
xor U14608 (N_14608,N_11892,N_10821);
xnor U14609 (N_14609,N_9169,N_10378);
or U14610 (N_14610,N_11383,N_9667);
or U14611 (N_14611,N_9369,N_10177);
nor U14612 (N_14612,N_10596,N_10765);
or U14613 (N_14613,N_9284,N_10863);
or U14614 (N_14614,N_9801,N_10436);
nor U14615 (N_14615,N_11274,N_11224);
nor U14616 (N_14616,N_9894,N_11332);
nor U14617 (N_14617,N_9668,N_10261);
nor U14618 (N_14618,N_10785,N_11524);
nor U14619 (N_14619,N_11028,N_9570);
and U14620 (N_14620,N_11880,N_10411);
or U14621 (N_14621,N_9081,N_9121);
or U14622 (N_14622,N_10020,N_10522);
or U14623 (N_14623,N_11665,N_9682);
nand U14624 (N_14624,N_9158,N_9385);
nand U14625 (N_14625,N_10595,N_10621);
nand U14626 (N_14626,N_10871,N_10128);
and U14627 (N_14627,N_10105,N_9209);
xor U14628 (N_14628,N_11218,N_10777);
and U14629 (N_14629,N_11535,N_9619);
nor U14630 (N_14630,N_9080,N_9883);
or U14631 (N_14631,N_11611,N_9178);
and U14632 (N_14632,N_9304,N_11622);
xnor U14633 (N_14633,N_10432,N_9375);
nand U14634 (N_14634,N_10816,N_11511);
nand U14635 (N_14635,N_10222,N_10958);
nand U14636 (N_14636,N_11425,N_11237);
xor U14637 (N_14637,N_11815,N_10041);
nand U14638 (N_14638,N_9731,N_11251);
and U14639 (N_14639,N_10392,N_9209);
and U14640 (N_14640,N_10325,N_9695);
xor U14641 (N_14641,N_9567,N_11712);
and U14642 (N_14642,N_9983,N_11994);
nand U14643 (N_14643,N_10542,N_10261);
and U14644 (N_14644,N_10087,N_9618);
nor U14645 (N_14645,N_11396,N_10079);
nand U14646 (N_14646,N_11528,N_9744);
xor U14647 (N_14647,N_9642,N_11738);
and U14648 (N_14648,N_9096,N_10391);
xor U14649 (N_14649,N_9799,N_11060);
xor U14650 (N_14650,N_9163,N_9612);
nand U14651 (N_14651,N_9069,N_10642);
nor U14652 (N_14652,N_9174,N_9433);
nor U14653 (N_14653,N_11325,N_9161);
nor U14654 (N_14654,N_9263,N_11570);
xor U14655 (N_14655,N_11092,N_9092);
nand U14656 (N_14656,N_9742,N_10624);
nand U14657 (N_14657,N_10228,N_10178);
xor U14658 (N_14658,N_11872,N_9648);
and U14659 (N_14659,N_10497,N_10054);
xor U14660 (N_14660,N_10865,N_10460);
and U14661 (N_14661,N_11600,N_9224);
nand U14662 (N_14662,N_9877,N_9465);
and U14663 (N_14663,N_11336,N_10098);
and U14664 (N_14664,N_9987,N_11842);
nand U14665 (N_14665,N_10111,N_9659);
nor U14666 (N_14666,N_10411,N_9114);
or U14667 (N_14667,N_10770,N_11474);
or U14668 (N_14668,N_9168,N_9678);
xnor U14669 (N_14669,N_9764,N_10022);
and U14670 (N_14670,N_9680,N_11134);
and U14671 (N_14671,N_9314,N_11117);
nor U14672 (N_14672,N_9824,N_10876);
or U14673 (N_14673,N_10711,N_11118);
nand U14674 (N_14674,N_9914,N_11237);
nand U14675 (N_14675,N_9867,N_11784);
and U14676 (N_14676,N_11015,N_11449);
nor U14677 (N_14677,N_9922,N_10417);
nand U14678 (N_14678,N_9936,N_11753);
nor U14679 (N_14679,N_10910,N_9593);
nor U14680 (N_14680,N_11941,N_9477);
or U14681 (N_14681,N_9372,N_11263);
nor U14682 (N_14682,N_9160,N_10373);
nor U14683 (N_14683,N_11310,N_9159);
xor U14684 (N_14684,N_11274,N_9202);
nor U14685 (N_14685,N_9394,N_11683);
xor U14686 (N_14686,N_9369,N_10562);
nor U14687 (N_14687,N_10346,N_10083);
nor U14688 (N_14688,N_10083,N_9138);
and U14689 (N_14689,N_10021,N_11444);
nand U14690 (N_14690,N_11895,N_10758);
xor U14691 (N_14691,N_10379,N_9831);
or U14692 (N_14692,N_9670,N_11309);
nand U14693 (N_14693,N_11329,N_9817);
xnor U14694 (N_14694,N_9819,N_10438);
and U14695 (N_14695,N_9953,N_11032);
and U14696 (N_14696,N_11481,N_9173);
and U14697 (N_14697,N_11464,N_9596);
and U14698 (N_14698,N_9380,N_10724);
xnor U14699 (N_14699,N_11059,N_9799);
xor U14700 (N_14700,N_10831,N_11784);
nor U14701 (N_14701,N_10123,N_10963);
nand U14702 (N_14702,N_10617,N_11375);
nor U14703 (N_14703,N_10974,N_9113);
xor U14704 (N_14704,N_9490,N_10864);
nor U14705 (N_14705,N_10666,N_11796);
and U14706 (N_14706,N_10940,N_11729);
or U14707 (N_14707,N_9652,N_10450);
or U14708 (N_14708,N_10485,N_10502);
nor U14709 (N_14709,N_11921,N_9540);
and U14710 (N_14710,N_11775,N_9395);
nor U14711 (N_14711,N_10128,N_11376);
nor U14712 (N_14712,N_10013,N_10591);
or U14713 (N_14713,N_11410,N_10614);
nor U14714 (N_14714,N_11522,N_11897);
and U14715 (N_14715,N_9598,N_11076);
and U14716 (N_14716,N_11171,N_9962);
xor U14717 (N_14717,N_10996,N_10036);
nor U14718 (N_14718,N_10688,N_9247);
or U14719 (N_14719,N_11457,N_11841);
nand U14720 (N_14720,N_11034,N_9765);
xnor U14721 (N_14721,N_9921,N_10317);
or U14722 (N_14722,N_10897,N_11770);
or U14723 (N_14723,N_11151,N_11175);
xor U14724 (N_14724,N_10692,N_11448);
and U14725 (N_14725,N_9286,N_9452);
or U14726 (N_14726,N_11245,N_9581);
and U14727 (N_14727,N_9928,N_10293);
nor U14728 (N_14728,N_9783,N_9977);
nor U14729 (N_14729,N_11548,N_11008);
and U14730 (N_14730,N_10481,N_11446);
or U14731 (N_14731,N_11199,N_10373);
xor U14732 (N_14732,N_11835,N_11883);
nand U14733 (N_14733,N_9196,N_9635);
nor U14734 (N_14734,N_9934,N_11733);
or U14735 (N_14735,N_9952,N_11421);
nand U14736 (N_14736,N_11390,N_10103);
nand U14737 (N_14737,N_9682,N_11939);
xor U14738 (N_14738,N_11763,N_10917);
or U14739 (N_14739,N_9413,N_11799);
nor U14740 (N_14740,N_11107,N_9696);
nor U14741 (N_14741,N_11336,N_11189);
xnor U14742 (N_14742,N_11394,N_11170);
and U14743 (N_14743,N_9904,N_9339);
and U14744 (N_14744,N_10105,N_11621);
xnor U14745 (N_14745,N_11966,N_10238);
nand U14746 (N_14746,N_9715,N_11876);
or U14747 (N_14747,N_11306,N_9924);
nor U14748 (N_14748,N_11218,N_11846);
nand U14749 (N_14749,N_10042,N_11870);
nand U14750 (N_14750,N_10078,N_10080);
and U14751 (N_14751,N_10306,N_11238);
nor U14752 (N_14752,N_11940,N_10043);
xnor U14753 (N_14753,N_11178,N_11016);
or U14754 (N_14754,N_9068,N_11889);
xor U14755 (N_14755,N_11301,N_11020);
nand U14756 (N_14756,N_10553,N_9291);
and U14757 (N_14757,N_9391,N_11086);
and U14758 (N_14758,N_9177,N_11289);
and U14759 (N_14759,N_11984,N_9247);
nand U14760 (N_14760,N_9672,N_9869);
nand U14761 (N_14761,N_11804,N_9778);
nand U14762 (N_14762,N_10784,N_10263);
nand U14763 (N_14763,N_11164,N_11805);
or U14764 (N_14764,N_11357,N_11287);
nand U14765 (N_14765,N_11933,N_10860);
nand U14766 (N_14766,N_10775,N_11204);
and U14767 (N_14767,N_10991,N_10309);
xnor U14768 (N_14768,N_11367,N_10499);
xor U14769 (N_14769,N_11546,N_11251);
nor U14770 (N_14770,N_9759,N_11061);
nor U14771 (N_14771,N_10746,N_9764);
nand U14772 (N_14772,N_11046,N_9756);
xor U14773 (N_14773,N_10107,N_10995);
and U14774 (N_14774,N_10349,N_9190);
and U14775 (N_14775,N_11568,N_9566);
nor U14776 (N_14776,N_11660,N_10110);
or U14777 (N_14777,N_10593,N_10749);
nor U14778 (N_14778,N_9779,N_10050);
xnor U14779 (N_14779,N_10745,N_10863);
nand U14780 (N_14780,N_9465,N_10899);
nand U14781 (N_14781,N_10966,N_10157);
nor U14782 (N_14782,N_10383,N_9120);
and U14783 (N_14783,N_11133,N_10999);
and U14784 (N_14784,N_11995,N_11949);
nor U14785 (N_14785,N_10714,N_9902);
nor U14786 (N_14786,N_9280,N_10630);
and U14787 (N_14787,N_9873,N_10774);
xor U14788 (N_14788,N_10371,N_9207);
xor U14789 (N_14789,N_9508,N_11261);
and U14790 (N_14790,N_10593,N_9230);
or U14791 (N_14791,N_11766,N_9696);
and U14792 (N_14792,N_10376,N_10039);
or U14793 (N_14793,N_11902,N_10135);
nand U14794 (N_14794,N_11664,N_10271);
nor U14795 (N_14795,N_10265,N_9689);
xnor U14796 (N_14796,N_10860,N_10946);
xor U14797 (N_14797,N_11384,N_9087);
xnor U14798 (N_14798,N_10016,N_11122);
nor U14799 (N_14799,N_11433,N_10484);
and U14800 (N_14800,N_11949,N_11826);
nor U14801 (N_14801,N_11166,N_9154);
nand U14802 (N_14802,N_9840,N_9278);
nor U14803 (N_14803,N_9244,N_9014);
or U14804 (N_14804,N_10677,N_9586);
xnor U14805 (N_14805,N_11063,N_10589);
nor U14806 (N_14806,N_11085,N_9951);
nand U14807 (N_14807,N_9527,N_9365);
xnor U14808 (N_14808,N_10469,N_10104);
and U14809 (N_14809,N_10007,N_11979);
xnor U14810 (N_14810,N_9921,N_11844);
or U14811 (N_14811,N_11820,N_9645);
or U14812 (N_14812,N_9808,N_10424);
and U14813 (N_14813,N_9736,N_11540);
and U14814 (N_14814,N_9054,N_11893);
nor U14815 (N_14815,N_9142,N_11947);
nor U14816 (N_14816,N_10719,N_9371);
xnor U14817 (N_14817,N_10296,N_11217);
xor U14818 (N_14818,N_9698,N_9109);
nand U14819 (N_14819,N_11253,N_11013);
nor U14820 (N_14820,N_11006,N_11885);
or U14821 (N_14821,N_10739,N_10348);
or U14822 (N_14822,N_11544,N_9929);
and U14823 (N_14823,N_9330,N_10508);
nor U14824 (N_14824,N_10855,N_10376);
nor U14825 (N_14825,N_9638,N_9539);
or U14826 (N_14826,N_10551,N_9498);
or U14827 (N_14827,N_10064,N_10338);
or U14828 (N_14828,N_10703,N_11701);
xor U14829 (N_14829,N_9245,N_9583);
nor U14830 (N_14830,N_9290,N_10942);
nor U14831 (N_14831,N_10769,N_9744);
and U14832 (N_14832,N_9370,N_11187);
xnor U14833 (N_14833,N_9010,N_9112);
nor U14834 (N_14834,N_11369,N_10772);
nor U14835 (N_14835,N_10379,N_10174);
or U14836 (N_14836,N_10190,N_10336);
and U14837 (N_14837,N_11966,N_10445);
and U14838 (N_14838,N_9350,N_9208);
nor U14839 (N_14839,N_10379,N_9218);
xor U14840 (N_14840,N_10017,N_10464);
xnor U14841 (N_14841,N_9516,N_10884);
xnor U14842 (N_14842,N_10667,N_10967);
and U14843 (N_14843,N_9347,N_9371);
nand U14844 (N_14844,N_11866,N_9281);
xor U14845 (N_14845,N_10013,N_10440);
nor U14846 (N_14846,N_11307,N_11949);
or U14847 (N_14847,N_11848,N_11331);
or U14848 (N_14848,N_10360,N_10618);
nand U14849 (N_14849,N_11534,N_10372);
nand U14850 (N_14850,N_9604,N_9364);
nand U14851 (N_14851,N_11799,N_10142);
nor U14852 (N_14852,N_9905,N_10658);
xor U14853 (N_14853,N_10557,N_10957);
nand U14854 (N_14854,N_9788,N_11850);
nor U14855 (N_14855,N_9485,N_10608);
and U14856 (N_14856,N_9678,N_10713);
and U14857 (N_14857,N_11581,N_11612);
nand U14858 (N_14858,N_11165,N_11736);
xor U14859 (N_14859,N_9406,N_11860);
and U14860 (N_14860,N_11488,N_9472);
nor U14861 (N_14861,N_10889,N_11298);
or U14862 (N_14862,N_10041,N_11274);
nand U14863 (N_14863,N_9366,N_11963);
and U14864 (N_14864,N_11129,N_11805);
nand U14865 (N_14865,N_11720,N_11272);
xor U14866 (N_14866,N_11372,N_10467);
and U14867 (N_14867,N_9683,N_10774);
xor U14868 (N_14868,N_10777,N_11390);
and U14869 (N_14869,N_9837,N_11902);
xor U14870 (N_14870,N_10638,N_10686);
xnor U14871 (N_14871,N_11167,N_10033);
xor U14872 (N_14872,N_9474,N_9515);
nor U14873 (N_14873,N_9098,N_10519);
nor U14874 (N_14874,N_9112,N_9453);
xnor U14875 (N_14875,N_10107,N_10917);
xnor U14876 (N_14876,N_10098,N_9566);
and U14877 (N_14877,N_9471,N_9407);
xor U14878 (N_14878,N_11707,N_10588);
xor U14879 (N_14879,N_10855,N_10915);
xor U14880 (N_14880,N_11407,N_9555);
xor U14881 (N_14881,N_10312,N_9449);
xnor U14882 (N_14882,N_11947,N_11517);
or U14883 (N_14883,N_10345,N_10544);
nor U14884 (N_14884,N_11585,N_9669);
nor U14885 (N_14885,N_9826,N_10554);
nand U14886 (N_14886,N_9789,N_10832);
and U14887 (N_14887,N_10566,N_9406);
or U14888 (N_14888,N_10927,N_10617);
or U14889 (N_14889,N_9017,N_9770);
and U14890 (N_14890,N_10626,N_10291);
xnor U14891 (N_14891,N_10861,N_11846);
xor U14892 (N_14892,N_9650,N_10240);
nand U14893 (N_14893,N_11673,N_11461);
and U14894 (N_14894,N_10804,N_10193);
xor U14895 (N_14895,N_10113,N_9487);
and U14896 (N_14896,N_11078,N_11050);
nor U14897 (N_14897,N_9447,N_10078);
or U14898 (N_14898,N_11166,N_10234);
or U14899 (N_14899,N_11997,N_11077);
and U14900 (N_14900,N_10241,N_11986);
nor U14901 (N_14901,N_11350,N_9205);
nand U14902 (N_14902,N_10846,N_9958);
xor U14903 (N_14903,N_11078,N_9550);
nor U14904 (N_14904,N_9514,N_11654);
or U14905 (N_14905,N_11061,N_10694);
xnor U14906 (N_14906,N_9946,N_9185);
nand U14907 (N_14907,N_11659,N_11231);
or U14908 (N_14908,N_9945,N_10975);
and U14909 (N_14909,N_10955,N_10471);
xor U14910 (N_14910,N_10113,N_9952);
nor U14911 (N_14911,N_10163,N_11139);
xor U14912 (N_14912,N_10191,N_11177);
and U14913 (N_14913,N_10564,N_9781);
nor U14914 (N_14914,N_10024,N_9230);
nor U14915 (N_14915,N_10978,N_9691);
and U14916 (N_14916,N_11125,N_11572);
or U14917 (N_14917,N_10706,N_9801);
nor U14918 (N_14918,N_11846,N_9980);
and U14919 (N_14919,N_10485,N_10748);
nand U14920 (N_14920,N_11448,N_9380);
xor U14921 (N_14921,N_10809,N_10242);
and U14922 (N_14922,N_9361,N_11447);
and U14923 (N_14923,N_11085,N_9277);
nor U14924 (N_14924,N_11882,N_11484);
xor U14925 (N_14925,N_9847,N_11645);
xnor U14926 (N_14926,N_11781,N_11384);
and U14927 (N_14927,N_10391,N_9927);
and U14928 (N_14928,N_11848,N_10345);
and U14929 (N_14929,N_10397,N_11217);
and U14930 (N_14930,N_9636,N_11472);
nand U14931 (N_14931,N_9122,N_10068);
nand U14932 (N_14932,N_10516,N_11456);
or U14933 (N_14933,N_9213,N_11740);
or U14934 (N_14934,N_9889,N_9846);
nand U14935 (N_14935,N_10405,N_11387);
or U14936 (N_14936,N_11314,N_10662);
and U14937 (N_14937,N_10501,N_10879);
nor U14938 (N_14938,N_11009,N_9161);
and U14939 (N_14939,N_9876,N_10630);
xnor U14940 (N_14940,N_11178,N_11577);
nor U14941 (N_14941,N_11830,N_10674);
nand U14942 (N_14942,N_11539,N_11638);
nand U14943 (N_14943,N_9992,N_11307);
xnor U14944 (N_14944,N_9321,N_10182);
and U14945 (N_14945,N_10989,N_9645);
nand U14946 (N_14946,N_9854,N_11029);
or U14947 (N_14947,N_9762,N_11464);
or U14948 (N_14948,N_9124,N_11467);
or U14949 (N_14949,N_10406,N_11624);
and U14950 (N_14950,N_9752,N_10256);
xor U14951 (N_14951,N_9234,N_11777);
or U14952 (N_14952,N_9209,N_9007);
or U14953 (N_14953,N_11232,N_10395);
and U14954 (N_14954,N_9342,N_10329);
nand U14955 (N_14955,N_10113,N_11075);
or U14956 (N_14956,N_10518,N_9550);
nand U14957 (N_14957,N_9096,N_9592);
nand U14958 (N_14958,N_10464,N_9744);
or U14959 (N_14959,N_10531,N_10482);
or U14960 (N_14960,N_11766,N_9572);
nand U14961 (N_14961,N_11184,N_10616);
nor U14962 (N_14962,N_10327,N_10264);
xor U14963 (N_14963,N_9376,N_11127);
or U14964 (N_14964,N_10181,N_11606);
and U14965 (N_14965,N_9666,N_10784);
nor U14966 (N_14966,N_11866,N_11978);
nand U14967 (N_14967,N_10324,N_9816);
nand U14968 (N_14968,N_10988,N_11992);
nand U14969 (N_14969,N_9141,N_11387);
and U14970 (N_14970,N_10050,N_11327);
nand U14971 (N_14971,N_10341,N_10352);
xor U14972 (N_14972,N_9993,N_11110);
or U14973 (N_14973,N_10719,N_11158);
or U14974 (N_14974,N_10109,N_11752);
nand U14975 (N_14975,N_11461,N_11721);
or U14976 (N_14976,N_11099,N_9992);
nand U14977 (N_14977,N_9394,N_9824);
or U14978 (N_14978,N_10532,N_11427);
and U14979 (N_14979,N_11691,N_10772);
nor U14980 (N_14980,N_9279,N_10124);
nand U14981 (N_14981,N_10877,N_11161);
or U14982 (N_14982,N_11879,N_10140);
or U14983 (N_14983,N_10301,N_10793);
xnor U14984 (N_14984,N_10261,N_11946);
nor U14985 (N_14985,N_11435,N_9502);
nand U14986 (N_14986,N_11398,N_11619);
and U14987 (N_14987,N_10158,N_10330);
or U14988 (N_14988,N_9990,N_9134);
nor U14989 (N_14989,N_9991,N_9166);
nand U14990 (N_14990,N_10165,N_9818);
or U14991 (N_14991,N_10159,N_10550);
nor U14992 (N_14992,N_11544,N_10686);
or U14993 (N_14993,N_11632,N_10124);
nand U14994 (N_14994,N_10320,N_11321);
or U14995 (N_14995,N_11686,N_10398);
xnor U14996 (N_14996,N_9711,N_9308);
nand U14997 (N_14997,N_10458,N_11956);
and U14998 (N_14998,N_9376,N_9510);
nor U14999 (N_14999,N_9931,N_11251);
or UO_0 (O_0,N_14248,N_12004);
nor UO_1 (O_1,N_13942,N_13758);
nand UO_2 (O_2,N_14371,N_14516);
or UO_3 (O_3,N_13209,N_14438);
or UO_4 (O_4,N_14720,N_14092);
and UO_5 (O_5,N_13249,N_14868);
xnor UO_6 (O_6,N_13029,N_12884);
xor UO_7 (O_7,N_12044,N_13906);
xor UO_8 (O_8,N_13581,N_14779);
nand UO_9 (O_9,N_14508,N_14096);
nand UO_10 (O_10,N_14550,N_13287);
and UO_11 (O_11,N_12805,N_12904);
nand UO_12 (O_12,N_12114,N_13233);
and UO_13 (O_13,N_14917,N_13598);
nor UO_14 (O_14,N_13722,N_12619);
nor UO_15 (O_15,N_14826,N_12618);
and UO_16 (O_16,N_14206,N_12738);
and UO_17 (O_17,N_12636,N_14789);
or UO_18 (O_18,N_14003,N_12871);
nand UO_19 (O_19,N_12315,N_13297);
xor UO_20 (O_20,N_12918,N_12401);
or UO_21 (O_21,N_12051,N_13450);
nand UO_22 (O_22,N_14776,N_14325);
or UO_23 (O_23,N_13790,N_14062);
nor UO_24 (O_24,N_13939,N_13898);
or UO_25 (O_25,N_13313,N_14835);
or UO_26 (O_26,N_13320,N_13378);
or UO_27 (O_27,N_14485,N_12715);
nor UO_28 (O_28,N_12100,N_14635);
xnor UO_29 (O_29,N_14945,N_14382);
nor UO_30 (O_30,N_12843,N_14319);
nor UO_31 (O_31,N_12197,N_12784);
xnor UO_32 (O_32,N_14712,N_14671);
nor UO_33 (O_33,N_12142,N_13867);
nand UO_34 (O_34,N_14555,N_14925);
and UO_35 (O_35,N_13031,N_14342);
nor UO_36 (O_36,N_13871,N_14472);
and UO_37 (O_37,N_12126,N_12534);
nand UO_38 (O_38,N_13769,N_14468);
or UO_39 (O_39,N_14402,N_12926);
nor UO_40 (O_40,N_13434,N_13159);
nand UO_41 (O_41,N_13030,N_12400);
nand UO_42 (O_42,N_13234,N_12943);
or UO_43 (O_43,N_14081,N_12091);
nor UO_44 (O_44,N_14164,N_14245);
nor UO_45 (O_45,N_12722,N_13724);
or UO_46 (O_46,N_14697,N_12644);
nand UO_47 (O_47,N_12087,N_13833);
and UO_48 (O_48,N_13124,N_14410);
nand UO_49 (O_49,N_13370,N_12676);
xor UO_50 (O_50,N_13281,N_13654);
and UO_51 (O_51,N_14037,N_13520);
xor UO_52 (O_52,N_14763,N_12081);
nor UO_53 (O_53,N_12632,N_14023);
or UO_54 (O_54,N_12421,N_13621);
or UO_55 (O_55,N_13932,N_14397);
xor UO_56 (O_56,N_12076,N_14258);
xor UO_57 (O_57,N_13256,N_12558);
or UO_58 (O_58,N_13967,N_14506);
nand UO_59 (O_59,N_13717,N_13672);
or UO_60 (O_60,N_14277,N_14218);
xor UO_61 (O_61,N_14788,N_13341);
or UO_62 (O_62,N_14955,N_13262);
nor UO_63 (O_63,N_14931,N_14898);
and UO_64 (O_64,N_13919,N_13042);
xor UO_65 (O_65,N_12121,N_14842);
nand UO_66 (O_66,N_14899,N_13106);
nor UO_67 (O_67,N_14591,N_14243);
and UO_68 (O_68,N_14974,N_14376);
nor UO_69 (O_69,N_12058,N_13893);
and UO_70 (O_70,N_13109,N_13447);
nand UO_71 (O_71,N_14230,N_13868);
xnor UO_72 (O_72,N_13556,N_12679);
xnor UO_73 (O_73,N_12913,N_12077);
or UO_74 (O_74,N_14878,N_12308);
and UO_75 (O_75,N_12690,N_13528);
xnor UO_76 (O_76,N_12949,N_12161);
xor UO_77 (O_77,N_12099,N_12356);
nor UO_78 (O_78,N_14991,N_13546);
or UO_79 (O_79,N_12245,N_13478);
and UO_80 (O_80,N_12007,N_12425);
nand UO_81 (O_81,N_14777,N_14191);
nor UO_82 (O_82,N_13537,N_14540);
nor UO_83 (O_83,N_13335,N_12958);
nor UO_84 (O_84,N_13795,N_14068);
and UO_85 (O_85,N_14006,N_14745);
nand UO_86 (O_86,N_14098,N_12916);
or UO_87 (O_87,N_14662,N_12629);
xnor UO_88 (O_88,N_12553,N_13436);
xor UO_89 (O_89,N_12300,N_13255);
or UO_90 (O_90,N_14348,N_14474);
nand UO_91 (O_91,N_14304,N_14874);
or UO_92 (O_92,N_13318,N_12964);
and UO_93 (O_93,N_12422,N_14061);
xnor UO_94 (O_94,N_14856,N_14774);
xor UO_95 (O_95,N_13583,N_12668);
nor UO_96 (O_96,N_12192,N_12413);
xor UO_97 (O_97,N_13702,N_14565);
and UO_98 (O_98,N_13531,N_13164);
and UO_99 (O_99,N_12180,N_12033);
nand UO_100 (O_100,N_13943,N_14606);
and UO_101 (O_101,N_13965,N_12117);
nor UO_102 (O_102,N_13259,N_12224);
or UO_103 (O_103,N_14205,N_12022);
nor UO_104 (O_104,N_12344,N_12795);
nor UO_105 (O_105,N_12677,N_12663);
nor UO_106 (O_106,N_14271,N_14155);
xor UO_107 (O_107,N_14244,N_12490);
or UO_108 (O_108,N_13728,N_13153);
nor UO_109 (O_109,N_13093,N_12439);
and UO_110 (O_110,N_12823,N_13477);
nand UO_111 (O_111,N_13529,N_12818);
nand UO_112 (O_112,N_14993,N_13397);
nor UO_113 (O_113,N_13718,N_12230);
nand UO_114 (O_114,N_13146,N_13078);
nand UO_115 (O_115,N_12900,N_14186);
or UO_116 (O_116,N_13165,N_14869);
xnor UO_117 (O_117,N_13211,N_12647);
xor UO_118 (O_118,N_14538,N_13612);
and UO_119 (O_119,N_13899,N_13482);
or UO_120 (O_120,N_12342,N_14743);
nor UO_121 (O_121,N_13483,N_13243);
nor UO_122 (O_122,N_14142,N_12516);
or UO_123 (O_123,N_14741,N_13872);
nand UO_124 (O_124,N_14957,N_14701);
and UO_125 (O_125,N_13316,N_12732);
nor UO_126 (O_126,N_13437,N_13996);
and UO_127 (O_127,N_13847,N_12312);
nor UO_128 (O_128,N_13055,N_12491);
or UO_129 (O_129,N_13610,N_13499);
nor UO_130 (O_130,N_12651,N_13552);
or UO_131 (O_131,N_12797,N_13570);
or UO_132 (O_132,N_13653,N_14041);
and UO_133 (O_133,N_12810,N_12469);
xor UO_134 (O_134,N_13665,N_14052);
xnor UO_135 (O_135,N_12073,N_12195);
nand UO_136 (O_136,N_12821,N_13559);
nor UO_137 (O_137,N_12997,N_12538);
xnor UO_138 (O_138,N_13513,N_13676);
and UO_139 (O_139,N_13380,N_14548);
xnor UO_140 (O_140,N_14350,N_13937);
xor UO_141 (O_141,N_12360,N_12567);
or UO_142 (O_142,N_12443,N_13538);
or UO_143 (O_143,N_13792,N_14463);
xor UO_144 (O_144,N_13971,N_12666);
and UO_145 (O_145,N_12637,N_13202);
nor UO_146 (O_146,N_12254,N_12890);
and UO_147 (O_147,N_12232,N_13726);
and UO_148 (O_148,N_13629,N_14707);
and UO_149 (O_149,N_13830,N_13772);
nand UO_150 (O_150,N_13801,N_14407);
and UO_151 (O_151,N_12447,N_14612);
xnor UO_152 (O_152,N_13828,N_12115);
or UO_153 (O_153,N_14769,N_14302);
xnor UO_154 (O_154,N_12909,N_13577);
xor UO_155 (O_155,N_12247,N_13983);
nor UO_156 (O_156,N_14781,N_13487);
nand UO_157 (O_157,N_13405,N_14306);
and UO_158 (O_158,N_13843,N_14074);
or UO_159 (O_159,N_12053,N_12525);
or UO_160 (O_160,N_13170,N_12955);
nor UO_161 (O_161,N_14631,N_13931);
nand UO_162 (O_162,N_12646,N_12454);
nand UO_163 (O_163,N_13574,N_13492);
or UO_164 (O_164,N_13825,N_13885);
or UO_165 (O_165,N_13310,N_13375);
or UO_166 (O_166,N_13043,N_14956);
xor UO_167 (O_167,N_13714,N_14927);
xor UO_168 (O_168,N_12207,N_12886);
and UO_169 (O_169,N_12063,N_14283);
and UO_170 (O_170,N_14887,N_14623);
xor UO_171 (O_171,N_12107,N_13144);
nor UO_172 (O_172,N_12354,N_14311);
nand UO_173 (O_173,N_12119,N_12075);
nor UO_174 (O_174,N_12580,N_13956);
or UO_175 (O_175,N_12378,N_14406);
or UO_176 (O_176,N_13275,N_13107);
nor UO_177 (O_177,N_13488,N_13486);
and UO_178 (O_178,N_14380,N_12640);
nor UO_179 (O_179,N_14080,N_14487);
xnor UO_180 (O_180,N_13510,N_12206);
nor UO_181 (O_181,N_14702,N_14175);
xnor UO_182 (O_182,N_13675,N_14816);
nand UO_183 (O_183,N_14532,N_12790);
nor UO_184 (O_184,N_12683,N_13567);
and UO_185 (O_185,N_14112,N_12578);
nor UO_186 (O_186,N_13926,N_12872);
or UO_187 (O_187,N_14576,N_13069);
nor UO_188 (O_188,N_12962,N_14423);
and UO_189 (O_189,N_14130,N_13196);
nor UO_190 (O_190,N_14113,N_13303);
nor UO_191 (O_191,N_13417,N_14111);
nand UO_192 (O_192,N_14054,N_12947);
and UO_193 (O_193,N_14568,N_13445);
and UO_194 (O_194,N_13362,N_14585);
nor UO_195 (O_195,N_12763,N_13184);
and UO_196 (O_196,N_14699,N_13509);
nor UO_197 (O_197,N_12485,N_12280);
nor UO_198 (O_198,N_12819,N_14169);
nor UO_199 (O_199,N_14501,N_13810);
nand UO_200 (O_200,N_14073,N_12084);
or UO_201 (O_201,N_12339,N_14024);
or UO_202 (O_202,N_13684,N_13814);
xnor UO_203 (O_203,N_14676,N_13511);
nand UO_204 (O_204,N_12542,N_14457);
nand UO_205 (O_205,N_12160,N_14910);
and UO_206 (O_206,N_12170,N_12950);
nand UO_207 (O_207,N_12513,N_14324);
nor UO_208 (O_208,N_12338,N_12687);
and UO_209 (O_209,N_14921,N_14126);
xor UO_210 (O_210,N_12524,N_14754);
nor UO_211 (O_211,N_13194,N_13517);
nand UO_212 (O_212,N_14195,N_12437);
nor UO_213 (O_213,N_12658,N_14920);
or UO_214 (O_214,N_12734,N_13875);
nor UO_215 (O_215,N_12768,N_12320);
or UO_216 (O_216,N_12585,N_12655);
nor UO_217 (O_217,N_13079,N_12220);
xnor UO_218 (O_218,N_14711,N_14505);
nor UO_219 (O_219,N_13803,N_13744);
or UO_220 (O_220,N_12435,N_13916);
or UO_221 (O_221,N_12897,N_12601);
and UO_222 (O_222,N_14251,N_14451);
xor UO_223 (O_223,N_13630,N_13306);
and UO_224 (O_224,N_12255,N_14780);
and UO_225 (O_225,N_14543,N_14851);
xor UO_226 (O_226,N_13688,N_14675);
and UO_227 (O_227,N_14043,N_12591);
xnor UO_228 (O_228,N_14118,N_13985);
and UO_229 (O_229,N_14886,N_14456);
xor UO_230 (O_230,N_14431,N_12630);
and UO_231 (O_231,N_14066,N_12019);
nand UO_232 (O_232,N_13840,N_13948);
and UO_233 (O_233,N_12587,N_13788);
nor UO_234 (O_234,N_13317,N_13323);
nor UO_235 (O_235,N_14286,N_14393);
nand UO_236 (O_236,N_13394,N_12132);
or UO_237 (O_237,N_12796,N_14400);
or UO_238 (O_238,N_13218,N_14018);
nor UO_239 (O_239,N_13749,N_12945);
nor UO_240 (O_240,N_14419,N_14137);
and UO_241 (O_241,N_12590,N_14087);
and UO_242 (O_242,N_13090,N_12480);
nand UO_243 (O_243,N_13992,N_14655);
nor UO_244 (O_244,N_14524,N_13009);
xor UO_245 (O_245,N_13530,N_12728);
nand UO_246 (O_246,N_12939,N_13314);
xor UO_247 (O_247,N_14071,N_13041);
nand UO_248 (O_248,N_14637,N_12592);
nand UO_249 (O_249,N_14978,N_12292);
nand UO_250 (O_250,N_13080,N_13823);
nor UO_251 (O_251,N_12769,N_13783);
nand UO_252 (O_252,N_12365,N_12062);
or UO_253 (O_253,N_13922,N_14847);
xor UO_254 (O_254,N_12282,N_12863);
xnor UO_255 (O_255,N_14625,N_13013);
and UO_256 (O_256,N_12102,N_12817);
nor UO_257 (O_257,N_12833,N_13426);
nor UO_258 (O_258,N_14417,N_14226);
xor UO_259 (O_259,N_12678,N_14272);
nor UO_260 (O_260,N_13748,N_13774);
nand UO_261 (O_261,N_13237,N_13099);
nand UO_262 (O_262,N_14976,N_13934);
or UO_263 (O_263,N_12698,N_12596);
or UO_264 (O_264,N_14904,N_13439);
xnor UO_265 (O_265,N_12188,N_14782);
or UO_266 (O_266,N_12340,N_13189);
or UO_267 (O_267,N_12462,N_12412);
xnor UO_268 (O_268,N_13293,N_13860);
and UO_269 (O_269,N_12731,N_12508);
and UO_270 (O_270,N_12605,N_14141);
xnor UO_271 (O_271,N_12735,N_14047);
or UO_272 (O_272,N_13601,N_14691);
xor UO_273 (O_273,N_14845,N_13897);
xor UO_274 (O_274,N_13096,N_14359);
and UO_275 (O_275,N_14048,N_12688);
or UO_276 (O_276,N_13644,N_14703);
nand UO_277 (O_277,N_13061,N_12070);
or UO_278 (O_278,N_13761,N_14704);
xnor UO_279 (O_279,N_12353,N_14039);
nand UO_280 (O_280,N_13851,N_14775);
and UO_281 (O_281,N_14454,N_14131);
xnor UO_282 (O_282,N_12749,N_13108);
nor UO_283 (O_283,N_14525,N_13576);
nand UO_284 (O_284,N_14409,N_12569);
nand UO_285 (O_285,N_12536,N_12438);
or UO_286 (O_286,N_14268,N_13207);
nand UO_287 (O_287,N_12766,N_14210);
nand UO_288 (O_288,N_14441,N_14069);
nand UO_289 (O_289,N_12093,N_13782);
and UO_290 (O_290,N_12992,N_13308);
xor UO_291 (O_291,N_14617,N_12083);
and UO_292 (O_292,N_14561,N_12330);
nand UO_293 (O_293,N_13890,N_14966);
nand UO_294 (O_294,N_13796,N_13444);
and UO_295 (O_295,N_13910,N_13565);
and UO_296 (O_296,N_14725,N_14193);
and UO_297 (O_297,N_14687,N_13240);
or UO_298 (O_298,N_13568,N_13283);
xnor UO_299 (O_299,N_12989,N_12164);
nand UO_300 (O_300,N_14385,N_13869);
or UO_301 (O_301,N_14837,N_14370);
nand UO_302 (O_302,N_14153,N_12429);
xnor UO_303 (O_303,N_12978,N_13590);
or UO_304 (O_304,N_14197,N_14345);
nand UO_305 (O_305,N_14426,N_13355);
xnor UO_306 (O_306,N_13519,N_14592);
or UO_307 (O_307,N_13642,N_14929);
xor UO_308 (O_308,N_14204,N_12285);
and UO_309 (O_309,N_12975,N_12377);
nand UO_310 (O_310,N_14822,N_13924);
nor UO_311 (O_311,N_12436,N_12082);
xnor UO_312 (O_312,N_14165,N_14187);
or UO_313 (O_313,N_12924,N_12737);
xnor UO_314 (O_314,N_12009,N_14852);
or UO_315 (O_315,N_12394,N_14241);
nand UO_316 (O_316,N_13637,N_14147);
and UO_317 (O_317,N_14088,N_12849);
and UO_318 (O_318,N_12951,N_13126);
nor UO_319 (O_319,N_14857,N_12139);
nor UO_320 (O_320,N_12969,N_12654);
nor UO_321 (O_321,N_14217,N_14751);
nand UO_322 (O_322,N_13682,N_13072);
nand UO_323 (O_323,N_13850,N_14573);
and UO_324 (O_324,N_13130,N_14876);
xnor UO_325 (O_325,N_14649,N_13379);
nor UO_326 (O_326,N_14049,N_14188);
or UO_327 (O_327,N_14101,N_13760);
and UO_328 (O_328,N_14808,N_13000);
nand UO_329 (O_329,N_13859,N_13549);
and UO_330 (O_330,N_12211,N_13414);
and UO_331 (O_331,N_14343,N_14552);
and UO_332 (O_332,N_13457,N_12457);
nor UO_333 (O_333,N_13994,N_13734);
or UO_334 (O_334,N_13648,N_14959);
nand UO_335 (O_335,N_14680,N_14354);
and UO_336 (O_336,N_13945,N_13589);
nand UO_337 (O_337,N_12675,N_14194);
and UO_338 (O_338,N_14850,N_12708);
nand UO_339 (O_339,N_12674,N_14365);
and UO_340 (O_340,N_14479,N_12294);
xnor UO_341 (O_341,N_13960,N_13753);
nand UO_342 (O_342,N_14526,N_14972);
nor UO_343 (O_343,N_13599,N_14174);
or UO_344 (O_344,N_13951,N_12550);
xor UO_345 (O_345,N_14378,N_13077);
nand UO_346 (O_346,N_13911,N_12695);
and UO_347 (O_347,N_12673,N_14119);
or UO_348 (O_348,N_12461,N_12561);
or UO_349 (O_349,N_14651,N_14519);
xnor UO_350 (O_350,N_14836,N_13349);
xor UO_351 (O_351,N_13606,N_13161);
or UO_352 (O_352,N_14867,N_14705);
nand UO_353 (O_353,N_12702,N_13004);
and UO_354 (O_354,N_13026,N_13972);
xor UO_355 (O_355,N_13770,N_14969);
or UO_356 (O_356,N_12466,N_12276);
or UO_357 (O_357,N_12216,N_13101);
nand UO_358 (O_358,N_13609,N_14148);
or UO_359 (O_359,N_12384,N_12842);
and UO_360 (O_360,N_13778,N_14323);
nand UO_361 (O_361,N_14284,N_12925);
nand UO_362 (O_362,N_13127,N_13432);
nor UO_363 (O_363,N_12523,N_12707);
and UO_364 (O_364,N_13266,N_12921);
and UO_365 (O_365,N_14854,N_12297);
nand UO_366 (O_366,N_12444,N_13175);
nand UO_367 (O_367,N_12003,N_13430);
xor UO_368 (O_368,N_12337,N_13908);
nor UO_369 (O_369,N_12193,N_13914);
and UO_370 (O_370,N_14677,N_12249);
nor UO_371 (O_371,N_14185,N_13640);
nand UO_372 (O_372,N_14333,N_13200);
and UO_373 (O_373,N_14178,N_14667);
nor UO_374 (O_374,N_14360,N_12816);
xnor UO_375 (O_375,N_13268,N_12392);
or UO_376 (O_376,N_14114,N_14940);
and UO_377 (O_377,N_12672,N_14733);
or UO_378 (O_378,N_14143,N_14716);
xor UO_379 (O_379,N_14880,N_14843);
and UO_380 (O_380,N_14428,N_12946);
nand UO_381 (O_381,N_14414,N_13846);
xnor UO_382 (O_382,N_14740,N_13856);
and UO_383 (O_383,N_12696,N_12803);
nand UO_384 (O_384,N_14465,N_14738);
nand UO_385 (O_385,N_12899,N_13928);
xor UO_386 (O_386,N_14918,N_12667);
and UO_387 (O_387,N_12028,N_13829);
or UO_388 (O_388,N_14575,N_12068);
nand UO_389 (O_389,N_13238,N_13618);
and UO_390 (O_390,N_14624,N_14116);
nand UO_391 (O_391,N_13235,N_12552);
nand UO_392 (O_392,N_13588,N_14714);
and UO_393 (O_393,N_12652,N_12915);
nand UO_394 (O_394,N_14427,N_12047);
nor UO_395 (O_395,N_13250,N_12465);
nand UO_396 (O_396,N_14085,N_14404);
or UO_397 (O_397,N_13876,N_14636);
and UO_398 (O_398,N_13001,N_14179);
or UO_399 (O_399,N_12256,N_14715);
and UO_400 (O_400,N_13604,N_12258);
nor UO_401 (O_401,N_13522,N_14466);
nor UO_402 (O_402,N_14616,N_14578);
xor UO_403 (O_403,N_14224,N_14100);
xor UO_404 (O_404,N_12172,N_13553);
nand UO_405 (O_405,N_13635,N_12775);
nand UO_406 (O_406,N_13157,N_14344);
nor UO_407 (O_407,N_12061,N_12124);
or UO_408 (O_408,N_13404,N_13221);
and UO_409 (O_409,N_12794,N_13961);
nor UO_410 (O_410,N_12554,N_14692);
nand UO_411 (O_411,N_13877,N_13952);
nor UO_412 (O_412,N_12684,N_12011);
and UO_413 (O_413,N_13424,N_14027);
nor UO_414 (O_414,N_13465,N_12039);
xor UO_415 (O_415,N_12638,N_12110);
nand UO_416 (O_416,N_12390,N_13594);
xnor UO_417 (O_417,N_14500,N_12246);
nand UO_418 (O_418,N_14828,N_14013);
or UO_419 (O_419,N_14234,N_12759);
xnor UO_420 (O_420,N_13946,N_14225);
nor UO_421 (O_421,N_14663,N_13578);
or UO_422 (O_422,N_13789,N_12577);
and UO_423 (O_423,N_12893,N_14388);
nor UO_424 (O_424,N_14864,N_14444);
and UO_425 (O_425,N_12458,N_14793);
xnor UO_426 (O_426,N_13712,N_12854);
and UO_427 (O_427,N_13651,N_13348);
nand UO_428 (O_428,N_14672,N_12807);
or UO_429 (O_429,N_12857,N_14510);
nor UO_430 (O_430,N_13120,N_14784);
or UO_431 (O_431,N_14522,N_13639);
or UO_432 (O_432,N_12791,N_12982);
nor UO_433 (O_433,N_12834,N_12518);
xnor UO_434 (O_434,N_14572,N_12289);
nand UO_435 (O_435,N_13862,N_13981);
nor UO_436 (O_436,N_14834,N_14229);
or UO_437 (O_437,N_14034,N_14176);
and UO_438 (O_438,N_13793,N_12034);
or UO_439 (O_439,N_13839,N_13536);
and UO_440 (O_440,N_12223,N_12616);
xnor UO_441 (O_441,N_12017,N_12574);
xor UO_442 (O_442,N_14610,N_12395);
nand UO_443 (O_443,N_13188,N_14737);
or UO_444 (O_444,N_12079,N_13681);
nand UO_445 (O_445,N_12944,N_14762);
and UO_446 (O_446,N_14798,N_14570);
nor UO_447 (O_447,N_14628,N_13959);
nand UO_448 (O_448,N_12650,N_14213);
and UO_449 (O_449,N_13707,N_14961);
nor UO_450 (O_450,N_13421,N_13678);
xor UO_451 (O_451,N_13446,N_13927);
nand UO_452 (O_452,N_14932,N_12305);
xnor UO_453 (O_453,N_13239,N_14936);
nand UO_454 (O_454,N_14795,N_12510);
xor UO_455 (O_455,N_13878,N_12937);
and UO_456 (O_456,N_12275,N_12877);
xnor UO_457 (O_457,N_14420,N_13371);
xnor UO_458 (O_458,N_13286,N_12136);
or UO_459 (O_459,N_14433,N_14012);
or UO_460 (O_460,N_12293,N_13141);
and UO_461 (O_461,N_14390,N_14266);
and UO_462 (O_462,N_12409,N_14689);
xnor UO_463 (O_463,N_12086,N_13560);
xor UO_464 (O_464,N_13067,N_13671);
and UO_465 (O_465,N_13708,N_14352);
or UO_466 (O_466,N_12729,N_13007);
nand UO_467 (O_467,N_12369,N_14764);
and UO_468 (O_468,N_13929,N_12383);
and UO_469 (O_469,N_13970,N_12482);
nor UO_470 (O_470,N_14660,N_14392);
or UO_471 (O_471,N_14829,N_14838);
or UO_472 (O_472,N_14813,N_12799);
nand UO_473 (O_473,N_12862,N_12993);
nand UO_474 (O_474,N_13245,N_14338);
or UO_475 (O_475,N_13251,N_14154);
and UO_476 (O_476,N_14440,N_14987);
xor UO_477 (O_477,N_13301,N_12311);
xnor UO_478 (O_478,N_14489,N_13427);
xnor UO_479 (O_479,N_12329,N_12196);
or UO_480 (O_480,N_14497,N_14952);
nor UO_481 (O_481,N_14462,N_12757);
nor UO_482 (O_482,N_13066,N_14491);
nor UO_483 (O_483,N_13525,N_13881);
xor UO_484 (O_484,N_13040,N_12645);
xor UO_485 (O_485,N_12270,N_12876);
nor UO_486 (O_486,N_12547,N_12097);
nand UO_487 (O_487,N_14328,N_14051);
nand UO_488 (O_488,N_14124,N_13035);
or UO_489 (O_489,N_14482,N_13302);
or UO_490 (O_490,N_12568,N_14391);
xor UO_491 (O_491,N_13294,N_13706);
xnor UO_492 (O_492,N_13279,N_12212);
or UO_493 (O_493,N_13091,N_14502);
and UO_494 (O_494,N_13563,N_13137);
nand UO_495 (O_495,N_13299,N_13889);
or UO_496 (O_496,N_14121,N_12328);
or UO_497 (O_497,N_13521,N_13181);
and UO_498 (O_498,N_13669,N_14220);
xnor UO_499 (O_499,N_14040,N_12231);
or UO_500 (O_500,N_13329,N_12050);
nor UO_501 (O_501,N_13385,N_12595);
or UO_502 (O_502,N_14953,N_14520);
nand UO_503 (O_503,N_12159,N_13305);
or UO_504 (O_504,N_12399,N_12244);
and UO_505 (O_505,N_13920,N_14928);
or UO_506 (O_506,N_14301,N_14812);
and UO_507 (O_507,N_14166,N_14412);
and UO_508 (O_508,N_14588,N_12856);
nand UO_509 (O_509,N_12938,N_14416);
or UO_510 (O_510,N_12357,N_12194);
nand UO_511 (O_511,N_13879,N_12131);
or UO_512 (O_512,N_13395,N_14010);
nor UO_513 (O_513,N_12200,N_13118);
nor UO_514 (O_514,N_12286,N_13811);
and UO_515 (O_515,N_13086,N_14718);
or UO_516 (O_516,N_14160,N_14846);
xnor UO_517 (O_517,N_13393,N_13296);
nor UO_518 (O_518,N_14364,N_12956);
nor UO_519 (O_519,N_14368,N_13232);
nand UO_520 (O_520,N_13062,N_13668);
and UO_521 (O_521,N_12977,N_12171);
nand UO_522 (O_522,N_13955,N_14923);
or UO_523 (O_523,N_13475,N_12999);
nand UO_524 (O_524,N_13364,N_14884);
or UO_525 (O_525,N_13277,N_14014);
or UO_526 (O_526,N_12191,N_12903);
nor UO_527 (O_527,N_13185,N_12971);
and UO_528 (O_528,N_14381,N_14076);
nor UO_529 (O_529,N_12895,N_14621);
or UO_530 (O_530,N_12317,N_12515);
nand UO_531 (O_531,N_13991,N_13622);
or UO_532 (O_532,N_14787,N_13183);
nor UO_533 (O_533,N_14123,N_13656);
and UO_534 (O_534,N_12622,N_13561);
nand UO_535 (O_535,N_14608,N_13799);
xnor UO_536 (O_536,N_12210,N_13800);
and UO_537 (O_537,N_13178,N_13104);
and UO_538 (O_538,N_14261,N_14021);
or UO_539 (O_539,N_13685,N_14279);
or UO_540 (O_540,N_12889,N_13613);
xor UO_541 (O_541,N_12049,N_13710);
or UO_542 (O_542,N_12815,N_12836);
and UO_543 (O_543,N_12880,N_14086);
or UO_544 (O_544,N_13659,N_14192);
nand UO_545 (O_545,N_13892,N_14478);
and UO_546 (O_546,N_12069,N_14529);
and UO_547 (O_547,N_13704,N_12549);
xor UO_548 (O_548,N_14445,N_13059);
nand UO_549 (O_549,N_13187,N_12301);
xor UO_550 (O_550,N_12464,N_14801);
nor UO_551 (O_551,N_14029,N_14558);
and UO_552 (O_552,N_12846,N_14989);
and UO_553 (O_553,N_14665,N_14181);
xnor UO_554 (O_554,N_14933,N_12844);
nor UO_555 (O_555,N_14227,N_14650);
and UO_556 (O_556,N_12288,N_13818);
xor UO_557 (O_557,N_14140,N_13870);
or UO_558 (O_558,N_13267,N_14819);
nand UO_559 (O_559,N_12106,N_12243);
and UO_560 (O_560,N_12907,N_14253);
nor UO_561 (O_561,N_12533,N_12064);
nand UO_562 (O_562,N_13735,N_12374);
nor UO_563 (O_563,N_13151,N_12426);
or UO_564 (O_564,N_12204,N_12333);
and UO_565 (O_565,N_13186,N_12038);
nor UO_566 (O_566,N_14150,N_12366);
and UO_567 (O_567,N_14581,N_13114);
or UO_568 (O_568,N_13337,N_13212);
or UO_569 (O_569,N_13095,N_13192);
nand UO_570 (O_570,N_12861,N_13498);
nand UO_571 (O_571,N_12748,N_14547);
nor UO_572 (O_572,N_13129,N_12407);
or UO_573 (O_573,N_13065,N_14903);
xnor UO_574 (O_574,N_12190,N_14282);
nor UO_575 (O_575,N_14639,N_12661);
and UO_576 (O_576,N_14128,N_14633);
and UO_577 (O_577,N_12229,N_13901);
xnor UO_578 (O_578,N_13731,N_13691);
xnor UO_579 (O_579,N_12140,N_12237);
and UO_580 (O_580,N_13696,N_14644);
nand UO_581 (O_581,N_12583,N_12347);
or UO_582 (O_582,N_13122,N_13057);
or UO_583 (O_583,N_12537,N_12382);
or UO_584 (O_584,N_13402,N_13806);
nand UO_585 (O_585,N_12316,N_13449);
and UO_586 (O_586,N_13584,N_12016);
or UO_587 (O_587,N_14536,N_12988);
nor UO_588 (O_588,N_13260,N_14270);
nand UO_589 (O_589,N_14577,N_13935);
nor UO_590 (O_590,N_14495,N_14563);
nor UO_591 (O_591,N_12700,N_13128);
nand UO_592 (O_592,N_12314,N_13431);
xor UO_593 (O_593,N_13649,N_13480);
or UO_594 (O_594,N_13587,N_13854);
nor UO_595 (O_595,N_13887,N_12631);
xor UO_596 (O_596,N_13372,N_14604);
nor UO_597 (O_597,N_12072,N_13933);
and UO_598 (O_598,N_13094,N_12548);
xor UO_599 (O_599,N_13285,N_13698);
nand UO_600 (O_600,N_14332,N_14807);
or UO_601 (O_601,N_12528,N_12752);
nand UO_602 (O_602,N_12801,N_13073);
xor UO_603 (O_603,N_12837,N_14814);
xor UO_604 (O_604,N_12624,N_12575);
nor UO_605 (O_605,N_14256,N_14435);
nand UO_606 (O_606,N_14240,N_13198);
nand UO_607 (O_607,N_14710,N_13028);
nor UO_608 (O_608,N_13990,N_13179);
nand UO_609 (O_609,N_14997,N_12671);
or UO_610 (O_610,N_13716,N_14984);
nor UO_611 (O_611,N_12570,N_14223);
or UO_612 (O_612,N_12104,N_13386);
or UO_613 (O_613,N_12074,N_14046);
or UO_614 (O_614,N_13116,N_12123);
nand UO_615 (O_615,N_14336,N_12265);
nand UO_616 (O_616,N_14449,N_12612);
and UO_617 (O_617,N_14168,N_12295);
xor UO_618 (O_618,N_13721,N_13176);
nand UO_619 (O_619,N_13205,N_13321);
xor UO_620 (O_620,N_14962,N_12056);
xnor UO_621 (O_621,N_13354,N_12980);
or UO_622 (O_622,N_12448,N_12633);
or UO_623 (O_623,N_12743,N_12642);
nor UO_624 (O_624,N_13220,N_13110);
and UO_625 (O_625,N_14896,N_14890);
xor UO_626 (O_626,N_13729,N_13248);
xnor UO_627 (O_627,N_12066,N_12754);
xor UO_628 (O_628,N_13039,N_14107);
xnor UO_629 (O_629,N_14470,N_13309);
xor UO_630 (O_630,N_14309,N_14724);
or UO_631 (O_631,N_13507,N_12770);
nor UO_632 (O_632,N_14432,N_14170);
or UO_633 (O_633,N_14411,N_14448);
xor UO_634 (O_634,N_14139,N_14603);
or UO_635 (O_635,N_12041,N_14642);
xnor UO_636 (O_636,N_13340,N_13155);
nor UO_637 (O_637,N_12878,N_12322);
xnor UO_638 (O_638,N_13473,N_12359);
or UO_639 (O_639,N_14221,N_14648);
or UO_640 (O_640,N_14646,N_14257);
xnor UO_641 (O_641,N_12455,N_13489);
or UO_642 (O_642,N_12419,N_12984);
nor UO_643 (O_643,N_13254,N_14653);
and UO_644 (O_644,N_12717,N_14252);
or UO_645 (O_645,N_14872,N_12917);
xor UO_646 (O_646,N_14157,N_13514);
and UO_647 (O_647,N_14439,N_13274);
and UO_648 (O_648,N_12213,N_13780);
nand UO_649 (O_649,N_13705,N_13280);
and UO_650 (O_650,N_13396,N_13481);
and UO_651 (O_651,N_13909,N_12539);
or UO_652 (O_652,N_14509,N_12726);
or UO_653 (O_653,N_13311,N_14207);
and UO_654 (O_654,N_12725,N_12681);
or UO_655 (O_655,N_13087,N_14512);
and UO_656 (O_656,N_14611,N_14494);
nand UO_657 (O_657,N_14654,N_14670);
and UO_658 (O_658,N_13425,N_12209);
and UO_659 (O_659,N_14326,N_12484);
or UO_660 (O_660,N_14973,N_12396);
nand UO_661 (O_661,N_12025,N_14216);
and UO_662 (O_662,N_13258,N_14916);
nor UO_663 (O_663,N_13365,N_12562);
nand UO_664 (O_664,N_14690,N_14693);
xor UO_665 (O_665,N_13428,N_13756);
xnor UO_666 (O_666,N_13504,N_12691);
nand UO_667 (O_667,N_13023,N_14467);
nor UO_668 (O_668,N_12736,N_14750);
nand UO_669 (O_669,N_13886,N_13036);
nand UO_670 (O_670,N_12670,N_13562);
or UO_671 (O_671,N_12589,N_13607);
xor UO_672 (O_672,N_14138,N_13557);
nand UO_673 (O_673,N_12983,N_14016);
xnor UO_674 (O_674,N_12839,N_12685);
nor UO_675 (O_675,N_13411,N_14477);
xor UO_676 (O_676,N_14627,N_13214);
xor UO_677 (O_677,N_13921,N_13253);
xnor UO_678 (O_678,N_13670,N_13980);
or UO_679 (O_679,N_14077,N_12427);
nor UO_680 (O_680,N_12236,N_14015);
or UO_681 (O_681,N_12036,N_12189);
xor UO_682 (O_682,N_13410,N_13471);
xor UO_683 (O_683,N_13468,N_14678);
and UO_684 (O_684,N_14228,N_14666);
xor UO_685 (O_685,N_13006,N_13138);
xnor UO_686 (O_686,N_14546,N_13938);
nor UO_687 (O_687,N_13742,N_12303);
nand UO_688 (O_688,N_13049,N_12767);
and UO_689 (O_689,N_14222,N_12781);
nor UO_690 (O_690,N_14935,N_12376);
or UO_691 (O_691,N_14602,N_13611);
nor UO_692 (O_692,N_13494,N_14236);
and UO_693 (O_693,N_14249,N_14695);
xor UO_694 (O_694,N_13540,N_13863);
xor UO_695 (O_695,N_12892,N_13284);
and UO_696 (O_696,N_14894,N_14749);
nor UO_697 (O_697,N_13794,N_12919);
nor UO_698 (O_698,N_14996,N_14316);
xor UO_699 (O_699,N_14356,N_13092);
nor UO_700 (O_700,N_14209,N_13051);
xor UO_701 (O_701,N_12764,N_12178);
nor UO_702 (O_702,N_13575,N_12067);
nor UO_703 (O_703,N_14329,N_13454);
or UO_704 (O_704,N_14944,N_14313);
nor UO_705 (O_705,N_14493,N_12222);
xnor UO_706 (O_706,N_12325,N_12348);
and UO_707 (O_707,N_14263,N_12942);
or UO_708 (O_708,N_12450,N_13845);
nand UO_709 (O_709,N_12141,N_13336);
and UO_710 (O_710,N_14308,N_14726);
xnor UO_711 (O_711,N_12792,N_13330);
nand UO_712 (O_712,N_13736,N_13779);
nor UO_713 (O_713,N_14199,N_13459);
xnor UO_714 (O_714,N_12018,N_12015);
xor UO_715 (O_715,N_14598,N_13673);
xnor UO_716 (O_716,N_12617,N_12755);
and UO_717 (O_717,N_13407,N_12742);
or UO_718 (O_718,N_14533,N_12380);
or UO_719 (O_719,N_12405,N_12446);
and UO_720 (O_720,N_12762,N_13203);
nor UO_721 (O_721,N_13491,N_12433);
nor UO_722 (O_722,N_12615,N_12156);
xnor UO_723 (O_723,N_13571,N_14219);
or UO_724 (O_724,N_14579,N_13663);
or UO_725 (O_725,N_13645,N_12827);
nor UO_726 (O_726,N_13527,N_14986);
and UO_727 (O_727,N_14958,N_12634);
nand UO_728 (O_728,N_14399,N_14492);
nand UO_729 (O_729,N_12987,N_14647);
and UO_730 (O_730,N_13484,N_12005);
and UO_731 (O_731,N_12535,N_14645);
or UO_732 (O_732,N_12719,N_14357);
nand UO_733 (O_733,N_13746,N_13787);
xnor UO_734 (O_734,N_14453,N_12598);
nor UO_735 (O_735,N_14802,N_12777);
xor UO_736 (O_736,N_13216,N_12478);
xnor UO_737 (O_737,N_12714,N_13230);
and UO_738 (O_738,N_14437,N_14208);
or UO_739 (O_739,N_13182,N_14900);
and UO_740 (O_740,N_14528,N_12253);
xnor UO_741 (O_741,N_13282,N_12682);
or UO_742 (O_742,N_12864,N_14202);
nor UO_743 (O_743,N_14870,N_13460);
xor UO_744 (O_744,N_12185,N_14099);
nor UO_745 (O_745,N_13304,N_14450);
nand UO_746 (O_746,N_13827,N_14883);
nor UO_747 (O_747,N_12239,N_14375);
xor UO_748 (O_748,N_12162,N_14171);
xnor UO_749 (O_749,N_14609,N_12641);
and UO_750 (O_750,N_13986,N_14875);
and UO_751 (O_751,N_12745,N_12505);
xor UO_752 (O_752,N_14937,N_12832);
nand UO_753 (O_753,N_14036,N_13711);
or UO_754 (O_754,N_14799,N_13322);
nand UO_755 (O_755,N_12135,N_12122);
nor UO_756 (O_756,N_13231,N_14708);
or UO_757 (O_757,N_14173,N_12785);
or UO_758 (O_758,N_12154,N_12299);
nand UO_759 (O_759,N_14369,N_12321);
and UO_760 (O_760,N_14044,N_13631);
xnor UO_761 (O_761,N_12351,N_12808);
or UO_762 (O_762,N_14395,N_13014);
or UO_763 (O_763,N_14753,N_14351);
or UO_764 (O_764,N_12867,N_12765);
xor UO_765 (O_765,N_13894,N_13834);
nand UO_766 (O_766,N_13797,N_13953);
or UO_767 (O_767,N_12125,N_12653);
or UO_768 (O_768,N_12221,N_12032);
nand UO_769 (O_769,N_12825,N_12071);
nand UO_770 (O_770,N_13852,N_13974);
and UO_771 (O_771,N_12665,N_13263);
and UO_772 (O_772,N_12309,N_13874);
nor UO_773 (O_773,N_13246,N_14861);
nor UO_774 (O_774,N_13333,N_13777);
or UO_775 (O_775,N_14167,N_13261);
nor UO_776 (O_776,N_13204,N_13750);
xnor UO_777 (O_777,N_13213,N_12248);
and UO_778 (O_778,N_14273,N_12198);
xor UO_779 (O_779,N_14698,N_14094);
or UO_780 (O_780,N_12506,N_13493);
and UO_781 (O_781,N_13052,N_12704);
xnor UO_782 (O_782,N_13347,N_12355);
and UO_783 (O_783,N_14688,N_13384);
or UO_784 (O_784,N_12559,N_13377);
nor UO_785 (O_785,N_13884,N_14067);
xnor UO_786 (O_786,N_13463,N_14535);
xor UO_787 (O_787,N_12403,N_13360);
nand UO_788 (O_788,N_14907,N_12588);
nand UO_789 (O_789,N_12474,N_14151);
and UO_790 (O_790,N_12440,N_12218);
and UO_791 (O_791,N_14290,N_12291);
nor UO_792 (O_792,N_12103,N_14362);
nand UO_793 (O_793,N_13627,N_13689);
nor UO_794 (O_794,N_12235,N_12411);
or UO_795 (O_795,N_12934,N_12787);
or UO_796 (O_796,N_14748,N_12471);
nand UO_797 (O_797,N_12363,N_12802);
nand UO_798 (O_798,N_14567,N_13923);
nand UO_799 (O_799,N_14664,N_14946);
and UO_800 (O_800,N_14490,N_14965);
nand UO_801 (O_801,N_14618,N_12532);
and UO_802 (O_802,N_14574,N_14817);
or UO_803 (O_803,N_14035,N_14736);
nor UO_804 (O_804,N_13617,N_13389);
nor UO_805 (O_805,N_13121,N_13667);
xor UO_806 (O_806,N_12467,N_13350);
nor UO_807 (O_807,N_12148,N_13105);
or UO_808 (O_808,N_12472,N_13591);
nor UO_809 (O_809,N_14215,N_12459);
or UO_810 (O_810,N_13154,N_13968);
nor UO_811 (O_811,N_13353,N_12875);
or UO_812 (O_812,N_12961,N_14394);
xor UO_813 (O_813,N_12774,N_13063);
nand UO_814 (O_814,N_13661,N_14366);
and UO_815 (O_815,N_12882,N_14805);
or UO_816 (O_816,N_12840,N_12397);
xnor UO_817 (O_817,N_14723,N_12381);
nand UO_818 (O_818,N_12606,N_12908);
nand UO_819 (O_819,N_13497,N_12176);
nand UO_820 (O_820,N_14582,N_12442);
nor UO_821 (O_821,N_13623,N_13602);
nor UO_822 (O_822,N_12416,N_13168);
xnor UO_823 (O_823,N_12522,N_13976);
xor UO_824 (O_824,N_14685,N_14291);
nand UO_825 (O_825,N_13423,N_12620);
xor UO_826 (O_826,N_14127,N_12800);
nor UO_827 (O_827,N_14082,N_12109);
nand UO_828 (O_828,N_12870,N_13060);
nand UO_829 (O_829,N_13915,N_14177);
xnor UO_830 (O_830,N_14310,N_14683);
nor UO_831 (O_831,N_12080,N_13677);
nor UO_832 (O_832,N_13033,N_14498);
and UO_833 (O_833,N_14760,N_13719);
nand UO_834 (O_834,N_14161,N_12307);
nor UO_835 (O_835,N_14815,N_14349);
nand UO_836 (O_836,N_12701,N_14521);
or UO_837 (O_837,N_14408,N_14607);
and UO_838 (O_838,N_13784,N_13808);
or UO_839 (O_839,N_14429,N_13543);
nand UO_840 (O_840,N_14305,N_12780);
and UO_841 (O_841,N_13429,N_12281);
nor UO_842 (O_842,N_13381,N_13495);
and UO_843 (O_843,N_12251,N_12565);
or UO_844 (O_844,N_12858,N_12501);
nand UO_845 (O_845,N_12252,N_12389);
nor UO_846 (O_846,N_13100,N_13145);
nor UO_847 (O_847,N_13135,N_14951);
nor UO_848 (O_848,N_14254,N_13500);
xnor UO_849 (O_849,N_13332,N_13741);
or UO_850 (O_850,N_13215,N_14544);
or UO_851 (O_851,N_14200,N_12199);
xnor UO_852 (O_852,N_12120,N_12557);
nor UO_853 (O_853,N_12225,N_14095);
or UO_854 (O_854,N_14596,N_13466);
nor UO_855 (O_855,N_14771,N_14990);
and UO_856 (O_856,N_13102,N_12563);
or UO_857 (O_857,N_14770,N_12709);
xor UO_858 (O_858,N_12147,N_13307);
xnor UO_859 (O_859,N_13097,N_12181);
or UO_860 (O_860,N_12756,N_14511);
nand UO_861 (O_861,N_12417,N_14564);
nand UO_862 (O_862,N_14963,N_12367);
nor UO_863 (O_863,N_12456,N_14700);
or UO_864 (O_864,N_13140,N_12259);
xnor UO_865 (O_865,N_13406,N_14979);
or UO_866 (O_866,N_14614,N_12694);
xnor UO_867 (O_867,N_13298,N_14706);
and UO_868 (O_868,N_13807,N_13047);
or UO_869 (O_869,N_12208,N_12489);
nand UO_870 (O_870,N_14971,N_12000);
and UO_871 (O_871,N_12452,N_14593);
nor UO_872 (O_872,N_14278,N_14436);
nor UO_873 (O_873,N_12930,N_13420);
xor UO_874 (O_874,N_14084,N_12773);
xor UO_875 (O_875,N_12976,N_13264);
xor UO_876 (O_876,N_14264,N_14943);
and UO_877 (O_877,N_13680,N_12529);
or UO_878 (O_878,N_12657,N_14237);
nand UO_879 (O_879,N_14732,N_12814);
xnor UO_880 (O_880,N_12820,N_12954);
and UO_881 (O_881,N_13658,N_14260);
xor UO_882 (O_882,N_14717,N_12920);
xor UO_883 (O_883,N_13312,N_14386);
and UO_884 (O_884,N_13995,N_13505);
nor UO_885 (O_885,N_13443,N_14327);
xor UO_886 (O_886,N_12798,N_13842);
nor UO_887 (O_887,N_14473,N_14559);
nor UO_888 (O_888,N_12346,N_14307);
or UO_889 (O_889,N_14599,N_12052);
xnor UO_890 (O_890,N_14825,N_14022);
and UO_891 (O_891,N_12133,N_14939);
nand UO_892 (O_892,N_13012,N_14792);
or UO_893 (O_893,N_13913,N_12973);
nor UO_894 (O_894,N_14486,N_14866);
nand UO_895 (O_895,N_14353,N_12788);
xnor UO_896 (O_896,N_13024,N_13666);
xor UO_897 (O_897,N_14267,N_14019);
nor UO_898 (O_898,N_14059,N_12431);
nand UO_899 (O_899,N_14605,N_13695);
and UO_900 (O_900,N_13008,N_14053);
xnor UO_901 (O_901,N_12334,N_12689);
and UO_902 (O_902,N_14523,N_12560);
nor UO_903 (O_903,N_14830,N_12970);
or UO_904 (O_904,N_14885,N_12628);
xor UO_905 (O_905,N_12186,N_12098);
xor UO_906 (O_906,N_13193,N_13117);
or UO_907 (O_907,N_12531,N_12789);
xor UO_908 (O_908,N_14183,N_14686);
xnor UO_909 (O_909,N_13614,N_13242);
and UO_910 (O_910,N_12520,N_12335);
nand UO_911 (O_911,N_13699,N_12906);
nor UO_912 (O_912,N_12094,N_13376);
xnor UO_913 (O_913,N_12613,N_14109);
and UO_914 (O_914,N_13327,N_12873);
nand UO_915 (O_915,N_13616,N_13743);
nand UO_916 (O_916,N_13442,N_14287);
or UO_917 (O_917,N_12497,N_13725);
xor UO_918 (O_918,N_14152,N_14281);
or UO_919 (O_919,N_14791,N_14129);
xnor UO_920 (O_920,N_13679,N_13973);
and UO_921 (O_921,N_14981,N_13542);
nor UO_922 (O_922,N_13819,N_14265);
or UO_923 (O_923,N_13941,N_13762);
and UO_924 (O_924,N_14734,N_14982);
nand UO_925 (O_925,N_12968,N_13025);
or UO_926 (O_926,N_14093,N_13858);
or UO_927 (O_927,N_14773,N_12241);
nand UO_928 (O_928,N_14657,N_13344);
xnor UO_929 (O_929,N_13315,N_12278);
nand UO_930 (O_930,N_13958,N_13342);
nand UO_931 (O_931,N_13132,N_12173);
and UO_932 (O_932,N_13324,N_12205);
nand UO_933 (O_933,N_12985,N_13413);
xor UO_934 (O_934,N_12931,N_12430);
nor UO_935 (O_935,N_14768,N_14079);
nand UO_936 (O_936,N_13496,N_13195);
xnor UO_937 (O_937,N_14484,N_12627);
nand UO_938 (O_938,N_14730,N_12020);
xor UO_939 (O_939,N_13390,N_12313);
nor UO_940 (O_940,N_13044,N_13226);
nor UO_941 (O_941,N_14571,N_13686);
and UO_942 (O_942,N_13628,N_12804);
nand UO_943 (O_943,N_13861,N_12498);
nor UO_944 (O_944,N_13608,N_12350);
or UO_945 (O_945,N_12914,N_14443);
nor UO_946 (O_946,N_13524,N_12996);
and UO_947 (O_947,N_14967,N_14877);
or UO_948 (O_948,N_13343,N_13334);
or UO_949 (O_949,N_13422,N_13056);
xnor UO_950 (O_950,N_14042,N_13755);
or UO_951 (O_951,N_14831,N_14430);
or UO_952 (O_952,N_13502,N_12543);
xnor UO_953 (O_953,N_12290,N_13300);
and UO_954 (O_954,N_12152,N_12262);
nor UO_955 (O_955,N_12492,N_14778);
nand UO_956 (O_956,N_12341,N_12847);
and UO_957 (O_957,N_13545,N_14070);
nor UO_958 (O_958,N_12868,N_14844);
or UO_959 (O_959,N_14507,N_14809);
and UO_960 (O_960,N_14772,N_13368);
nand UO_961 (O_961,N_12519,N_13366);
xor UO_962 (O_962,N_13766,N_14994);
and UO_963 (O_963,N_14026,N_13768);
nand UO_964 (O_964,N_14330,N_13815);
xor UO_965 (O_965,N_14295,N_14358);
nor UO_966 (O_966,N_13083,N_12593);
and UO_967 (O_967,N_14106,N_13148);
and UO_968 (O_968,N_12739,N_13358);
xnor UO_969 (O_969,N_13359,N_12226);
xor UO_970 (O_970,N_12928,N_14089);
or UO_971 (O_971,N_14597,N_12349);
or UO_972 (O_972,N_14065,N_13821);
xnor UO_973 (O_973,N_14800,N_13620);
and UO_974 (O_974,N_13015,N_12323);
xnor UO_975 (O_975,N_12546,N_13902);
xor UO_976 (O_976,N_12393,N_14985);
nor UO_977 (O_977,N_14679,N_12604);
nor UO_978 (O_978,N_12138,N_13352);
nand UO_979 (O_979,N_13539,N_14634);
nand UO_980 (O_980,N_14919,N_12151);
xor UO_981 (O_981,N_14804,N_12656);
or UO_982 (O_982,N_14515,N_12896);
nor UO_983 (O_983,N_13415,N_13745);
nor UO_984 (O_984,N_14001,N_14398);
or UO_985 (O_985,N_13723,N_12273);
xor UO_986 (O_986,N_14211,N_12108);
nor UO_987 (O_987,N_12240,N_12850);
nand UO_988 (O_988,N_13374,N_13224);
and UO_989 (O_989,N_12812,N_12610);
xnor UO_990 (O_990,N_13270,N_14103);
or UO_991 (O_991,N_13022,N_13002);
nand UO_992 (O_992,N_13526,N_13569);
nor UO_993 (O_993,N_12597,N_14480);
nor UO_994 (O_994,N_13554,N_12990);
nor UO_995 (O_995,N_14820,N_14613);
and UO_996 (O_996,N_13088,N_12163);
xnor UO_997 (O_997,N_14214,N_14580);
xnor UO_998 (O_998,N_13085,N_12324);
nand UO_999 (O_999,N_14823,N_14425);
or UO_1000 (O_1000,N_12527,N_13201);
xor UO_1001 (O_1001,N_14401,N_14909);
and UO_1002 (O_1002,N_12626,N_14496);
nand UO_1003 (O_1003,N_13119,N_14942);
nand UO_1004 (O_1004,N_14058,N_14948);
nand UO_1005 (O_1005,N_14363,N_13977);
or UO_1006 (O_1006,N_13555,N_13048);
and UO_1007 (O_1007,N_12112,N_12703);
and UO_1008 (O_1008,N_12470,N_13461);
or UO_1009 (O_1009,N_13011,N_14853);
and UO_1010 (O_1010,N_13882,N_12571);
nor UO_1011 (O_1011,N_12364,N_12137);
and UO_1012 (O_1012,N_13156,N_14105);
xor UO_1013 (O_1013,N_12116,N_13896);
nand UO_1014 (O_1014,N_12388,N_14145);
or UO_1015 (O_1015,N_14911,N_12361);
nor UO_1016 (O_1016,N_13173,N_14902);
xor UO_1017 (O_1017,N_12952,N_13177);
nand UO_1018 (O_1018,N_13751,N_12783);
and UO_1019 (O_1019,N_14590,N_14924);
nor UO_1020 (O_1020,N_12545,N_14004);
nor UO_1021 (O_1021,N_12238,N_12408);
and UO_1022 (O_1022,N_12723,N_14134);
and UO_1023 (O_1023,N_13081,N_12509);
or UO_1024 (O_1024,N_14233,N_13357);
or UO_1025 (O_1025,N_12166,N_13167);
nand UO_1026 (O_1026,N_12445,N_12932);
and UO_1027 (O_1027,N_12760,N_12806);
and UO_1028 (O_1028,N_14367,N_14008);
nor UO_1029 (O_1029,N_13573,N_13998);
or UO_1030 (O_1030,N_14652,N_13664);
xnor UO_1031 (O_1031,N_12564,N_12250);
or UO_1032 (O_1032,N_12879,N_14274);
and UO_1033 (O_1033,N_12706,N_12424);
and UO_1034 (O_1034,N_13786,N_12746);
xnor UO_1035 (O_1035,N_14339,N_12933);
xor UO_1036 (O_1036,N_14102,N_12234);
nand UO_1037 (O_1037,N_13966,N_12811);
nor UO_1038 (O_1038,N_13925,N_13210);
or UO_1039 (O_1039,N_13512,N_13223);
nor UO_1040 (O_1040,N_12566,N_14045);
or UO_1041 (O_1041,N_13626,N_13978);
nand UO_1042 (O_1042,N_14235,N_12782);
xor UO_1043 (O_1043,N_13291,N_14794);
xor UO_1044 (O_1044,N_13027,N_12831);
xnor UO_1045 (O_1045,N_13162,N_12130);
and UO_1046 (O_1046,N_13433,N_14159);
nand UO_1047 (O_1047,N_13988,N_12608);
nand UO_1048 (O_1048,N_13709,N_13038);
nand UO_1049 (O_1049,N_13150,N_13172);
nand UO_1050 (O_1050,N_14954,N_13021);
and UO_1051 (O_1051,N_14072,N_14063);
nor UO_1052 (O_1052,N_12128,N_12511);
or UO_1053 (O_1053,N_13400,N_14396);
or UO_1054 (O_1054,N_12586,N_13070);
and UO_1055 (O_1055,N_12948,N_12368);
xor UO_1056 (O_1056,N_14584,N_13435);
nor UO_1057 (O_1057,N_13771,N_14641);
nand UO_1058 (O_1058,N_13848,N_13276);
nor UO_1059 (O_1059,N_13523,N_14761);
and UO_1060 (O_1060,N_14011,N_12261);
or UO_1061 (O_1061,N_14684,N_14031);
nor UO_1062 (O_1062,N_13633,N_14541);
and UO_1063 (O_1063,N_13596,N_14818);
and UO_1064 (O_1064,N_12991,N_12113);
nand UO_1065 (O_1065,N_13816,N_12826);
nor UO_1066 (O_1066,N_13190,N_14858);
xor UO_1067 (O_1067,N_14461,N_14747);
nor UO_1068 (O_1068,N_14146,N_14259);
or UO_1069 (O_1069,N_13764,N_14594);
or UO_1070 (O_1070,N_12182,N_13269);
and UO_1071 (O_1071,N_12143,N_14901);
and UO_1072 (O_1072,N_14839,N_13046);
or UO_1073 (O_1073,N_14180,N_12848);
and UO_1074 (O_1074,N_14299,N_14009);
nor UO_1075 (O_1075,N_14905,N_12874);
nor UO_1076 (O_1076,N_12555,N_12242);
or UO_1077 (O_1077,N_13288,N_14293);
nand UO_1078 (O_1078,N_13662,N_12935);
and UO_1079 (O_1079,N_14231,N_14452);
and UO_1080 (O_1080,N_13826,N_13133);
and UO_1081 (O_1081,N_14156,N_14162);
or UO_1082 (O_1082,N_12887,N_13657);
nand UO_1083 (O_1083,N_13836,N_14097);
and UO_1084 (O_1084,N_12486,N_12055);
nand UO_1085 (O_1085,N_12214,N_13273);
and UO_1086 (O_1086,N_14755,N_12727);
and UO_1087 (O_1087,N_13975,N_12495);
nor UO_1088 (O_1088,N_14569,N_14891);
xnor UO_1089 (O_1089,N_14586,N_12852);
or UO_1090 (O_1090,N_14314,N_14560);
or UO_1091 (O_1091,N_12502,N_13409);
nor UO_1092 (O_1092,N_12434,N_12972);
or UO_1093 (O_1093,N_14122,N_13638);
nand UO_1094 (O_1094,N_14000,N_13715);
or UO_1095 (O_1095,N_14163,N_13603);
nor UO_1096 (O_1096,N_13652,N_13440);
xnor UO_1097 (O_1097,N_14504,N_12713);
nand UO_1098 (O_1098,N_12953,N_13804);
and UO_1099 (O_1099,N_14488,N_13257);
xor UO_1100 (O_1100,N_12277,N_13962);
or UO_1101 (O_1101,N_12526,N_14995);
or UO_1102 (O_1102,N_14849,N_13544);
and UO_1103 (O_1103,N_14889,N_14032);
xor UO_1104 (O_1104,N_13999,N_12866);
or UO_1105 (O_1105,N_12127,N_13982);
nor UO_1106 (O_1106,N_14442,N_14539);
nand UO_1107 (O_1107,N_13050,N_13624);
nor UO_1108 (O_1108,N_14198,N_12860);
or UO_1109 (O_1109,N_14553,N_12183);
nor UO_1110 (O_1110,N_12008,N_14172);
or UO_1111 (O_1111,N_12974,N_12168);
nand UO_1112 (O_1112,N_12035,N_12995);
nor UO_1113 (O_1113,N_14721,N_14212);
nand UO_1114 (O_1114,N_13905,N_12331);
nand UO_1115 (O_1115,N_12960,N_12415);
or UO_1116 (O_1116,N_14873,N_13551);
and UO_1117 (O_1117,N_13740,N_14656);
or UO_1118 (O_1118,N_12203,N_12406);
or UO_1119 (O_1119,N_14335,N_14731);
nor UO_1120 (O_1120,N_12838,N_14970);
nand UO_1121 (O_1121,N_12105,N_13319);
or UO_1122 (O_1122,N_14514,N_14537);
nor UO_1123 (O_1123,N_14673,N_13798);
nor UO_1124 (O_1124,N_12556,N_12059);
nor UO_1125 (O_1125,N_12268,N_14292);
xnor UO_1126 (O_1126,N_13018,N_13388);
xor UO_1127 (O_1127,N_13053,N_14530);
and UO_1128 (O_1128,N_13016,N_14483);
xnor UO_1129 (O_1129,N_14373,N_13767);
nor UO_1130 (O_1130,N_13247,N_14947);
xor UO_1131 (O_1131,N_13169,N_13082);
and UO_1132 (O_1132,N_13533,N_14934);
or UO_1133 (O_1133,N_12027,N_12697);
or UO_1134 (O_1134,N_12386,N_12149);
nor UO_1135 (O_1135,N_14133,N_14296);
nand UO_1136 (O_1136,N_13289,N_12664);
nor UO_1137 (O_1137,N_12283,N_14557);
and UO_1138 (O_1138,N_12012,N_13775);
and UO_1139 (O_1139,N_14895,N_12998);
or UO_1140 (O_1140,N_14811,N_14346);
or UO_1141 (O_1141,N_12581,N_12144);
nand UO_1142 (O_1142,N_14104,N_12089);
nor UO_1143 (O_1143,N_14796,N_13582);
or UO_1144 (O_1144,N_12753,N_12319);
xor UO_1145 (O_1145,N_12145,N_14025);
nor UO_1146 (O_1146,N_12940,N_12287);
and UO_1147 (O_1147,N_12432,N_13690);
and UO_1148 (O_1148,N_13865,N_13813);
and UO_1149 (O_1149,N_14334,N_12219);
and UO_1150 (O_1150,N_14638,N_12822);
nor UO_1151 (O_1151,N_13241,N_12101);
xor UO_1152 (O_1152,N_14832,N_12362);
and UO_1153 (O_1153,N_13418,N_14285);
or UO_1154 (O_1154,N_12750,N_14766);
nor UO_1155 (O_1155,N_13625,N_13401);
or UO_1156 (O_1156,N_14262,N_13832);
nor UO_1157 (O_1157,N_13883,N_12398);
and UO_1158 (O_1158,N_14298,N_13139);
and UO_1159 (O_1159,N_13820,N_13534);
nor UO_1160 (O_1160,N_13074,N_12090);
xnor UO_1161 (O_1161,N_12635,N_14744);
nand UO_1162 (O_1162,N_14999,N_14056);
xor UO_1163 (O_1163,N_14643,N_13438);
or UO_1164 (O_1164,N_13501,N_13700);
xor UO_1165 (O_1165,N_14297,N_14742);
nand UO_1166 (O_1166,N_12054,N_13730);
or UO_1167 (O_1167,N_12521,N_12648);
nand UO_1168 (O_1168,N_12479,N_14549);
xor UO_1169 (O_1169,N_12504,N_14661);
xor UO_1170 (O_1170,N_12751,N_13619);
nand UO_1171 (O_1171,N_14403,N_14735);
or UO_1172 (O_1172,N_14865,N_13328);
and UO_1173 (O_1173,N_13032,N_14545);
or UO_1174 (O_1174,N_12318,N_12551);
nor UO_1175 (O_1175,N_14998,N_12088);
or UO_1176 (O_1176,N_12451,N_14786);
nand UO_1177 (O_1177,N_12343,N_14132);
nand UO_1178 (O_1178,N_13111,N_13142);
xor UO_1179 (O_1179,N_14476,N_12306);
nand UO_1180 (O_1180,N_13076,N_12336);
xnor UO_1181 (O_1181,N_12579,N_12046);
or UO_1182 (O_1182,N_12488,N_14387);
xor UO_1183 (O_1183,N_14632,N_13034);
and UO_1184 (O_1184,N_14908,N_12352);
xnor UO_1185 (O_1185,N_13338,N_14158);
xnor UO_1186 (O_1186,N_13687,N_12639);
xnor UO_1187 (O_1187,N_13558,N_13351);
and UO_1188 (O_1188,N_13660,N_13399);
nand UO_1189 (O_1189,N_13453,N_14988);
nor UO_1190 (O_1190,N_13936,N_14002);
xor UO_1191 (O_1191,N_13532,N_12923);
or UO_1192 (O_1192,N_14418,N_12659);
xor UO_1193 (O_1193,N_12517,N_14746);
xor UO_1194 (O_1194,N_14057,N_14658);
nand UO_1195 (O_1195,N_12941,N_12881);
and UO_1196 (O_1196,N_12721,N_14583);
or UO_1197 (O_1197,N_13382,N_12410);
nor UO_1198 (O_1198,N_14629,N_14806);
or UO_1199 (O_1199,N_13115,N_14960);
or UO_1200 (O_1200,N_12187,N_12594);
or UO_1201 (O_1201,N_14320,N_12026);
or UO_1202 (O_1202,N_13003,N_12201);
or UO_1203 (O_1203,N_14203,N_14144);
nor UO_1204 (O_1204,N_13005,N_13547);
or UO_1205 (O_1205,N_12599,N_13701);
nand UO_1206 (O_1206,N_14331,N_14424);
or UO_1207 (O_1207,N_14078,N_14765);
and UO_1208 (O_1208,N_13646,N_13855);
and UO_1209 (O_1209,N_14110,N_12660);
or UO_1210 (O_1210,N_12830,N_12582);
xor UO_1211 (O_1211,N_13451,N_13416);
nor UO_1212 (O_1212,N_14992,N_13112);
nand UO_1213 (O_1213,N_12922,N_12959);
nor UO_1214 (O_1214,N_12986,N_14860);
xnor UO_1215 (O_1215,N_12600,N_13954);
and UO_1216 (O_1216,N_12607,N_12169);
and UO_1217 (O_1217,N_12001,N_12228);
nand UO_1218 (O_1218,N_12625,N_12649);
nor UO_1219 (O_1219,N_14091,N_13697);
nor UO_1220 (O_1220,N_12494,N_12428);
and UO_1221 (O_1221,N_13113,N_13947);
and UO_1222 (O_1222,N_14255,N_13479);
xor UO_1223 (O_1223,N_13809,N_12888);
or UO_1224 (O_1224,N_14460,N_14915);
nor UO_1225 (O_1225,N_13738,N_13949);
or UO_1226 (O_1226,N_13548,N_12037);
nor UO_1227 (O_1227,N_14189,N_14855);
or UO_1228 (O_1228,N_14455,N_13773);
nand UO_1229 (O_1229,N_12724,N_14848);
nand UO_1230 (O_1230,N_13217,N_14681);
xor UO_1231 (O_1231,N_14601,N_14983);
and UO_1232 (O_1232,N_14615,N_12423);
nor UO_1233 (O_1233,N_12835,N_14347);
or UO_1234 (O_1234,N_13831,N_14620);
nor UO_1235 (O_1235,N_14682,N_12449);
xnor UO_1236 (O_1236,N_12379,N_13837);
xor UO_1237 (O_1237,N_13964,N_12692);
nor UO_1238 (O_1238,N_12095,N_13641);
nand UO_1239 (O_1239,N_12503,N_12898);
xor UO_1240 (O_1240,N_14783,N_14475);
or UO_1241 (O_1241,N_13595,N_14600);
xnor UO_1242 (O_1242,N_12643,N_12177);
and UO_1243 (O_1243,N_14810,N_14803);
and UO_1244 (O_1244,N_13391,N_14595);
xor UO_1245 (O_1245,N_12264,N_14863);
nor UO_1246 (O_1246,N_14912,N_13817);
or UO_1247 (O_1247,N_13470,N_13398);
nor UO_1248 (O_1248,N_14276,N_12883);
and UO_1249 (O_1249,N_13580,N_13252);
and UO_1250 (O_1250,N_12475,N_14300);
and UO_1251 (O_1251,N_14242,N_14005);
or UO_1252 (O_1252,N_13747,N_13448);
and UO_1253 (O_1253,N_13472,N_13222);
nand UO_1254 (O_1254,N_13010,N_12021);
or UO_1255 (O_1255,N_12263,N_12621);
xor UO_1256 (O_1256,N_14115,N_14017);
or UO_1257 (O_1257,N_12092,N_13737);
or UO_1258 (O_1258,N_12891,N_13597);
nand UO_1259 (O_1259,N_12693,N_13880);
nand UO_1260 (O_1260,N_13292,N_12758);
and UO_1261 (O_1261,N_13752,N_13841);
nand UO_1262 (O_1262,N_14881,N_12741);
xor UO_1263 (O_1263,N_14882,N_12514);
xnor UO_1264 (O_1264,N_12391,N_12902);
nand UO_1265 (O_1265,N_13089,N_12129);
or UO_1266 (O_1266,N_14246,N_13197);
nand UO_1267 (O_1267,N_12460,N_12267);
nand UO_1268 (O_1268,N_12387,N_14108);
or UO_1269 (O_1269,N_13634,N_12304);
nand UO_1270 (O_1270,N_14238,N_14384);
and UO_1271 (O_1271,N_12609,N_12859);
xor UO_1272 (O_1272,N_13045,N_12441);
and UO_1273 (O_1273,N_12085,N_12463);
and UO_1274 (O_1274,N_14269,N_13506);
or UO_1275 (O_1275,N_14247,N_14696);
and UO_1276 (O_1276,N_13857,N_14551);
or UO_1277 (O_1277,N_13888,N_12905);
and UO_1278 (O_1278,N_13064,N_14879);
nand UO_1279 (O_1279,N_12855,N_12911);
or UO_1280 (O_1280,N_14315,N_14922);
and UO_1281 (O_1281,N_13326,N_13084);
or UO_1282 (O_1282,N_13290,N_12584);
and UO_1283 (O_1283,N_12711,N_12994);
nor UO_1284 (O_1284,N_13989,N_12912);
nand UO_1285 (O_1285,N_14372,N_14930);
nand UO_1286 (O_1286,N_12869,N_13361);
xnor UO_1287 (O_1287,N_14566,N_12060);
or UO_1288 (O_1288,N_12761,N_13191);
nor UO_1289 (O_1289,N_12468,N_14824);
nor UO_1290 (O_1290,N_14321,N_14503);
nor UO_1291 (O_1291,N_13900,N_14383);
or UO_1292 (O_1292,N_12266,N_13383);
or UO_1293 (O_1293,N_13944,N_12284);
or UO_1294 (O_1294,N_13208,N_12158);
nand UO_1295 (O_1295,N_12157,N_14413);
and UO_1296 (O_1296,N_13727,N_13508);
nand UO_1297 (O_1297,N_12669,N_12712);
nand UO_1298 (O_1298,N_12227,N_13593);
xnor UO_1299 (O_1299,N_13346,N_12134);
or UO_1300 (O_1300,N_12184,N_12029);
nand UO_1301 (O_1301,N_12981,N_13592);
and UO_1302 (O_1302,N_13503,N_12372);
xnor UO_1303 (O_1303,N_13822,N_13541);
xor UO_1304 (O_1304,N_12345,N_13732);
xor UO_1305 (O_1305,N_12483,N_12786);
nand UO_1306 (O_1306,N_12260,N_12175);
nand UO_1307 (O_1307,N_14759,N_13776);
and UO_1308 (O_1308,N_13103,N_14713);
or UO_1309 (O_1309,N_14694,N_14028);
or UO_1310 (O_1310,N_12865,N_12078);
nor UO_1311 (O_1311,N_12740,N_14821);
or UO_1312 (O_1312,N_14446,N_14064);
xor UO_1313 (O_1313,N_12965,N_12048);
nor UO_1314 (O_1314,N_14125,N_13518);
nor UO_1315 (O_1315,N_12813,N_13987);
nand UO_1316 (O_1316,N_13957,N_14728);
or UO_1317 (O_1317,N_13997,N_13791);
and UO_1318 (O_1318,N_13058,N_12414);
nand UO_1319 (O_1319,N_14337,N_14379);
nor UO_1320 (O_1320,N_13891,N_12174);
or UO_1321 (O_1321,N_13441,N_13586);
nand UO_1322 (O_1322,N_12611,N_13408);
nand UO_1323 (O_1323,N_13019,N_12512);
and UO_1324 (O_1324,N_13136,N_12507);
xnor UO_1325 (O_1325,N_14294,N_13765);
nand UO_1326 (O_1326,N_14840,N_13585);
nor UO_1327 (O_1327,N_14841,N_12002);
nor UO_1328 (O_1328,N_12779,N_12680);
xnor UO_1329 (O_1329,N_13904,N_13265);
xnor UO_1330 (O_1330,N_12771,N_13278);
and UO_1331 (O_1331,N_12371,N_13550);
or UO_1332 (O_1332,N_13918,N_12065);
nor UO_1333 (O_1333,N_13647,N_13469);
nand UO_1334 (O_1334,N_13225,N_12013);
or UO_1335 (O_1335,N_12358,N_14893);
nor UO_1336 (O_1336,N_12686,N_13158);
or UO_1337 (O_1337,N_13516,N_12851);
xnor UO_1338 (O_1338,N_12057,N_13853);
and UO_1339 (O_1339,N_12370,N_14968);
and UO_1340 (O_1340,N_13713,N_12540);
or UO_1341 (O_1341,N_12024,N_13844);
nor UO_1342 (O_1342,N_14075,N_14182);
or UO_1343 (O_1343,N_14464,N_13849);
or UO_1344 (O_1344,N_12500,N_12699);
nor UO_1345 (O_1345,N_14083,N_13467);
nor UO_1346 (O_1346,N_12576,N_14674);
or UO_1347 (O_1347,N_14318,N_14626);
and UO_1348 (O_1348,N_14587,N_14060);
nor UO_1349 (O_1349,N_14622,N_13674);
nand UO_1350 (O_1350,N_13979,N_14120);
and UO_1351 (O_1351,N_14459,N_12927);
nor UO_1352 (O_1352,N_13535,N_12385);
or UO_1353 (O_1353,N_12274,N_13757);
nor UO_1354 (O_1354,N_14964,N_13692);
nor UO_1355 (O_1355,N_12279,N_14729);
and UO_1356 (O_1356,N_14136,N_13166);
nor UO_1357 (O_1357,N_14562,N_13605);
or UO_1358 (O_1358,N_13969,N_12326);
or UO_1359 (O_1359,N_14554,N_12966);
xor UO_1360 (O_1360,N_14341,N_14669);
or UO_1361 (O_1361,N_12118,N_14469);
and UO_1362 (O_1362,N_13917,N_12023);
nor UO_1363 (O_1363,N_13632,N_14038);
and UO_1364 (O_1364,N_14977,N_14790);
and UO_1365 (O_1365,N_14030,N_13733);
nor UO_1366 (O_1366,N_13452,N_13174);
or UO_1367 (O_1367,N_12030,N_12705);
nor UO_1368 (O_1368,N_12179,N_13229);
nor UO_1369 (O_1369,N_13228,N_14859);
or UO_1370 (O_1370,N_14196,N_13054);
and UO_1371 (O_1371,N_13295,N_13835);
or UO_1372 (O_1372,N_13993,N_12623);
xnor UO_1373 (O_1373,N_12845,N_13131);
nor UO_1374 (O_1374,N_14926,N_14719);
or UO_1375 (O_1375,N_12894,N_12718);
and UO_1376 (O_1376,N_13643,N_13940);
and UO_1377 (O_1377,N_12499,N_14767);
nand UO_1378 (O_1378,N_12829,N_12487);
nand UO_1379 (O_1379,N_13458,N_14556);
nor UO_1380 (O_1380,N_12146,N_12614);
nor UO_1381 (O_1381,N_13455,N_12901);
xnor UO_1382 (O_1382,N_13693,N_14827);
nor UO_1383 (O_1383,N_13485,N_12747);
or UO_1384 (O_1384,N_14322,N_13636);
xnor UO_1385 (O_1385,N_13419,N_13134);
nand UO_1386 (O_1386,N_14317,N_13236);
or UO_1387 (O_1387,N_14513,N_13963);
xor UO_1388 (O_1388,N_14630,N_12662);
xnor UO_1389 (O_1389,N_12929,N_13412);
and UO_1390 (O_1390,N_13075,N_12809);
and UO_1391 (O_1391,N_14757,N_13367);
xnor UO_1392 (O_1392,N_13271,N_12710);
nand UO_1393 (O_1393,N_14447,N_12327);
nand UO_1394 (O_1394,N_14374,N_12476);
nand UO_1395 (O_1395,N_14980,N_12153);
xor UO_1396 (O_1396,N_13392,N_13369);
nor UO_1397 (O_1397,N_13272,N_14913);
or UO_1398 (O_1398,N_14531,N_13476);
xor UO_1399 (O_1399,N_12477,N_12824);
nand UO_1400 (O_1400,N_14542,N_12014);
xor UO_1401 (O_1401,N_14275,N_12418);
and UO_1402 (O_1402,N_13907,N_14897);
xnor UO_1403 (O_1403,N_14619,N_13147);
nand UO_1404 (O_1404,N_12006,N_12573);
nand UO_1405 (O_1405,N_13125,N_14055);
nand UO_1406 (O_1406,N_13160,N_12215);
or UO_1407 (O_1407,N_12404,N_13171);
or UO_1408 (O_1408,N_13703,N_12853);
xnor UO_1409 (O_1409,N_13930,N_14361);
or UO_1410 (O_1410,N_14871,N_13566);
xor UO_1411 (O_1411,N_14421,N_13227);
or UO_1412 (O_1412,N_14020,N_13802);
nand UO_1413 (O_1413,N_12776,N_12269);
xnor UO_1414 (O_1414,N_13683,N_14938);
xor UO_1415 (O_1415,N_13403,N_14727);
nor UO_1416 (O_1416,N_13017,N_14797);
nand UO_1417 (O_1417,N_14135,N_12031);
nor UO_1418 (O_1418,N_12310,N_12603);
nand UO_1419 (O_1419,N_14941,N_12298);
or UO_1420 (O_1420,N_12716,N_14184);
and UO_1421 (O_1421,N_13781,N_13345);
nor UO_1422 (O_1422,N_13615,N_14471);
nand UO_1423 (O_1423,N_12957,N_13655);
xnor UO_1424 (O_1424,N_13462,N_13325);
or UO_1425 (O_1425,N_12841,N_14250);
or UO_1426 (O_1426,N_13564,N_13363);
xnor UO_1427 (O_1427,N_13339,N_14975);
nor UO_1428 (O_1428,N_12473,N_12217);
and UO_1429 (O_1429,N_13515,N_14340);
xnor UO_1430 (O_1430,N_14892,N_12979);
or UO_1431 (O_1431,N_12375,N_12963);
xnor UO_1432 (O_1432,N_13600,N_13244);
xor UO_1433 (O_1433,N_13824,N_12420);
nor UO_1434 (O_1434,N_13739,N_13199);
xor UO_1435 (O_1435,N_14517,N_13020);
xor UO_1436 (O_1436,N_13387,N_12493);
nand UO_1437 (O_1437,N_14758,N_14289);
nand UO_1438 (O_1438,N_14312,N_12572);
and UO_1439 (O_1439,N_12828,N_14201);
or UO_1440 (O_1440,N_12402,N_13474);
and UO_1441 (O_1441,N_12373,N_12910);
and UO_1442 (O_1442,N_12155,N_14007);
or UO_1443 (O_1443,N_13950,N_12793);
xnor UO_1444 (O_1444,N_14668,N_13163);
nand UO_1445 (O_1445,N_12010,N_14239);
xor UO_1446 (O_1446,N_13152,N_14589);
or UO_1447 (O_1447,N_14785,N_12481);
nand UO_1448 (O_1448,N_12165,N_13206);
nand UO_1449 (O_1449,N_13149,N_13812);
nor UO_1450 (O_1450,N_12936,N_14090);
or UO_1451 (O_1451,N_12544,N_14659);
nor UO_1452 (O_1452,N_13895,N_14033);
or UO_1453 (O_1453,N_13098,N_13694);
and UO_1454 (O_1454,N_14906,N_14914);
and UO_1455 (O_1455,N_14534,N_12045);
nand UO_1456 (O_1456,N_14117,N_14422);
or UO_1457 (O_1457,N_13071,N_12730);
xnor UO_1458 (O_1458,N_12111,N_12040);
xnor UO_1459 (O_1459,N_12167,N_12043);
xor UO_1460 (O_1460,N_13805,N_14527);
or UO_1461 (O_1461,N_12720,N_13759);
and UO_1462 (O_1462,N_14499,N_13903);
and UO_1463 (O_1463,N_13219,N_14458);
and UO_1464 (O_1464,N_14640,N_13763);
nor UO_1465 (O_1465,N_12257,N_14888);
xor UO_1466 (O_1466,N_13866,N_12541);
and UO_1467 (O_1467,N_13356,N_12496);
xnor UO_1468 (O_1468,N_12885,N_12744);
nand UO_1469 (O_1469,N_12150,N_14303);
nor UO_1470 (O_1470,N_12096,N_13572);
nand UO_1471 (O_1471,N_14190,N_13912);
or UO_1472 (O_1472,N_13464,N_14389);
nand UO_1473 (O_1473,N_12042,N_12271);
and UO_1474 (O_1474,N_12967,N_12772);
or UO_1475 (O_1475,N_14722,N_14050);
or UO_1476 (O_1476,N_14149,N_14756);
nor UO_1477 (O_1477,N_14405,N_13456);
xnor UO_1478 (O_1478,N_13123,N_14280);
xnor UO_1479 (O_1479,N_12453,N_13579);
nand UO_1480 (O_1480,N_13373,N_13864);
xnor UO_1481 (O_1481,N_12733,N_14833);
xor UO_1482 (O_1482,N_12202,N_13068);
and UO_1483 (O_1483,N_13143,N_14862);
or UO_1484 (O_1484,N_14232,N_12272);
nand UO_1485 (O_1485,N_14355,N_14752);
and UO_1486 (O_1486,N_12778,N_13037);
nand UO_1487 (O_1487,N_14288,N_14481);
or UO_1488 (O_1488,N_13331,N_13650);
xnor UO_1489 (O_1489,N_14518,N_13838);
and UO_1490 (O_1490,N_13720,N_12296);
nand UO_1491 (O_1491,N_13180,N_13785);
or UO_1492 (O_1492,N_12302,N_14377);
nor UO_1493 (O_1493,N_12602,N_14434);
nor UO_1494 (O_1494,N_12332,N_13984);
nand UO_1495 (O_1495,N_14739,N_14415);
or UO_1496 (O_1496,N_13754,N_14950);
nor UO_1497 (O_1497,N_12530,N_13873);
or UO_1498 (O_1498,N_14709,N_13490);
xnor UO_1499 (O_1499,N_14949,N_12233);
nor UO_1500 (O_1500,N_12331,N_12868);
nor UO_1501 (O_1501,N_12177,N_12927);
xnor UO_1502 (O_1502,N_14017,N_13943);
nor UO_1503 (O_1503,N_13022,N_12177);
nand UO_1504 (O_1504,N_14971,N_12483);
xor UO_1505 (O_1505,N_12469,N_12059);
nand UO_1506 (O_1506,N_12235,N_12234);
or UO_1507 (O_1507,N_12355,N_13471);
and UO_1508 (O_1508,N_13313,N_12075);
nand UO_1509 (O_1509,N_14893,N_13556);
nand UO_1510 (O_1510,N_14532,N_14128);
xor UO_1511 (O_1511,N_12069,N_12585);
nand UO_1512 (O_1512,N_14862,N_13357);
xnor UO_1513 (O_1513,N_12182,N_14556);
nor UO_1514 (O_1514,N_13971,N_13502);
nor UO_1515 (O_1515,N_13690,N_12151);
nor UO_1516 (O_1516,N_14045,N_14409);
nor UO_1517 (O_1517,N_13358,N_14418);
or UO_1518 (O_1518,N_13967,N_12123);
nand UO_1519 (O_1519,N_13848,N_14957);
nor UO_1520 (O_1520,N_14468,N_14841);
nand UO_1521 (O_1521,N_12488,N_13755);
nor UO_1522 (O_1522,N_12727,N_13888);
or UO_1523 (O_1523,N_12157,N_12017);
nor UO_1524 (O_1524,N_12389,N_14858);
nor UO_1525 (O_1525,N_12547,N_13933);
or UO_1526 (O_1526,N_13022,N_13416);
and UO_1527 (O_1527,N_13559,N_13798);
xnor UO_1528 (O_1528,N_14362,N_13159);
or UO_1529 (O_1529,N_12657,N_12662);
or UO_1530 (O_1530,N_12372,N_13280);
and UO_1531 (O_1531,N_12114,N_12327);
nor UO_1532 (O_1532,N_13245,N_14311);
nand UO_1533 (O_1533,N_14043,N_12956);
nor UO_1534 (O_1534,N_14683,N_13176);
xor UO_1535 (O_1535,N_14835,N_14305);
and UO_1536 (O_1536,N_13275,N_14497);
xnor UO_1537 (O_1537,N_14366,N_14078);
and UO_1538 (O_1538,N_12322,N_13109);
and UO_1539 (O_1539,N_14646,N_14270);
nand UO_1540 (O_1540,N_12133,N_14827);
or UO_1541 (O_1541,N_12604,N_13020);
nand UO_1542 (O_1542,N_13403,N_13217);
or UO_1543 (O_1543,N_14242,N_13415);
nand UO_1544 (O_1544,N_13744,N_14020);
and UO_1545 (O_1545,N_14097,N_12969);
nand UO_1546 (O_1546,N_14183,N_14697);
or UO_1547 (O_1547,N_13812,N_13366);
or UO_1548 (O_1548,N_13343,N_14664);
xnor UO_1549 (O_1549,N_13593,N_12108);
and UO_1550 (O_1550,N_13773,N_13343);
nand UO_1551 (O_1551,N_13365,N_13923);
xnor UO_1552 (O_1552,N_14443,N_13105);
nor UO_1553 (O_1553,N_14063,N_13449);
nand UO_1554 (O_1554,N_13066,N_13854);
nor UO_1555 (O_1555,N_14143,N_13854);
nand UO_1556 (O_1556,N_14251,N_12172);
nand UO_1557 (O_1557,N_12022,N_14309);
nand UO_1558 (O_1558,N_12871,N_12537);
nor UO_1559 (O_1559,N_13786,N_13663);
xor UO_1560 (O_1560,N_13214,N_13083);
and UO_1561 (O_1561,N_13254,N_14299);
or UO_1562 (O_1562,N_14726,N_14364);
xnor UO_1563 (O_1563,N_13901,N_14398);
or UO_1564 (O_1564,N_12788,N_14123);
nand UO_1565 (O_1565,N_12663,N_12239);
or UO_1566 (O_1566,N_14021,N_12085);
nand UO_1567 (O_1567,N_13893,N_13248);
nor UO_1568 (O_1568,N_14321,N_13239);
and UO_1569 (O_1569,N_14269,N_13683);
nor UO_1570 (O_1570,N_12322,N_12848);
or UO_1571 (O_1571,N_13458,N_12642);
nand UO_1572 (O_1572,N_14303,N_12196);
nand UO_1573 (O_1573,N_14931,N_14364);
nand UO_1574 (O_1574,N_12882,N_12818);
nand UO_1575 (O_1575,N_12700,N_13469);
or UO_1576 (O_1576,N_12106,N_13352);
nand UO_1577 (O_1577,N_12046,N_12558);
and UO_1578 (O_1578,N_12088,N_12469);
nand UO_1579 (O_1579,N_14730,N_13907);
nor UO_1580 (O_1580,N_14459,N_14848);
nor UO_1581 (O_1581,N_12436,N_14915);
nand UO_1582 (O_1582,N_12022,N_12574);
nor UO_1583 (O_1583,N_14449,N_12687);
nand UO_1584 (O_1584,N_12330,N_14445);
or UO_1585 (O_1585,N_14927,N_14190);
or UO_1586 (O_1586,N_12510,N_12386);
nor UO_1587 (O_1587,N_13440,N_14749);
xor UO_1588 (O_1588,N_14163,N_13172);
nand UO_1589 (O_1589,N_13086,N_14044);
and UO_1590 (O_1590,N_13852,N_14903);
and UO_1591 (O_1591,N_14956,N_13869);
and UO_1592 (O_1592,N_14799,N_12485);
and UO_1593 (O_1593,N_12969,N_13430);
and UO_1594 (O_1594,N_12749,N_14459);
and UO_1595 (O_1595,N_14390,N_12404);
nand UO_1596 (O_1596,N_12418,N_14849);
nand UO_1597 (O_1597,N_13090,N_13710);
xnor UO_1598 (O_1598,N_14477,N_14746);
or UO_1599 (O_1599,N_12484,N_14646);
or UO_1600 (O_1600,N_12261,N_13000);
xor UO_1601 (O_1601,N_13213,N_13004);
xnor UO_1602 (O_1602,N_13326,N_14647);
xnor UO_1603 (O_1603,N_12100,N_14366);
nor UO_1604 (O_1604,N_12427,N_14281);
or UO_1605 (O_1605,N_14426,N_13479);
nand UO_1606 (O_1606,N_13617,N_14302);
xnor UO_1607 (O_1607,N_13409,N_13534);
and UO_1608 (O_1608,N_14542,N_13106);
and UO_1609 (O_1609,N_13879,N_13647);
and UO_1610 (O_1610,N_13365,N_12989);
xor UO_1611 (O_1611,N_13782,N_12769);
nand UO_1612 (O_1612,N_13254,N_13297);
nor UO_1613 (O_1613,N_12554,N_13398);
nand UO_1614 (O_1614,N_12486,N_14984);
xnor UO_1615 (O_1615,N_13911,N_13099);
nor UO_1616 (O_1616,N_13492,N_13931);
nand UO_1617 (O_1617,N_14596,N_13527);
and UO_1618 (O_1618,N_14060,N_14663);
nand UO_1619 (O_1619,N_14458,N_13509);
and UO_1620 (O_1620,N_12095,N_13522);
or UO_1621 (O_1621,N_13106,N_13129);
xnor UO_1622 (O_1622,N_14727,N_12192);
nor UO_1623 (O_1623,N_14174,N_14586);
xnor UO_1624 (O_1624,N_14138,N_12580);
or UO_1625 (O_1625,N_13446,N_13627);
xor UO_1626 (O_1626,N_13970,N_14785);
or UO_1627 (O_1627,N_14443,N_13869);
xor UO_1628 (O_1628,N_13221,N_14447);
nand UO_1629 (O_1629,N_12602,N_13702);
nor UO_1630 (O_1630,N_13081,N_14636);
xnor UO_1631 (O_1631,N_12394,N_14165);
and UO_1632 (O_1632,N_13522,N_13810);
or UO_1633 (O_1633,N_12962,N_12307);
xnor UO_1634 (O_1634,N_14372,N_14877);
nand UO_1635 (O_1635,N_12173,N_14846);
nor UO_1636 (O_1636,N_13609,N_12199);
or UO_1637 (O_1637,N_14487,N_13155);
nor UO_1638 (O_1638,N_13965,N_12383);
nand UO_1639 (O_1639,N_14861,N_13705);
or UO_1640 (O_1640,N_13626,N_13607);
xor UO_1641 (O_1641,N_13340,N_12696);
or UO_1642 (O_1642,N_14738,N_12024);
nor UO_1643 (O_1643,N_14607,N_12155);
nand UO_1644 (O_1644,N_12358,N_12930);
nor UO_1645 (O_1645,N_12432,N_14412);
xnor UO_1646 (O_1646,N_14880,N_14680);
or UO_1647 (O_1647,N_14243,N_12968);
nor UO_1648 (O_1648,N_13324,N_13819);
nand UO_1649 (O_1649,N_14571,N_12051);
or UO_1650 (O_1650,N_13134,N_13441);
or UO_1651 (O_1651,N_13453,N_13368);
xnor UO_1652 (O_1652,N_12222,N_14125);
or UO_1653 (O_1653,N_14633,N_14402);
nand UO_1654 (O_1654,N_14945,N_12022);
and UO_1655 (O_1655,N_14832,N_13233);
nor UO_1656 (O_1656,N_13247,N_14232);
or UO_1657 (O_1657,N_12806,N_13507);
nand UO_1658 (O_1658,N_12859,N_13014);
nand UO_1659 (O_1659,N_13433,N_14522);
xnor UO_1660 (O_1660,N_13128,N_14383);
xor UO_1661 (O_1661,N_13806,N_12677);
or UO_1662 (O_1662,N_12710,N_12149);
nor UO_1663 (O_1663,N_14360,N_12416);
xnor UO_1664 (O_1664,N_12706,N_14821);
nand UO_1665 (O_1665,N_12310,N_12605);
or UO_1666 (O_1666,N_13044,N_12597);
nor UO_1667 (O_1667,N_14632,N_14526);
nand UO_1668 (O_1668,N_14470,N_12745);
or UO_1669 (O_1669,N_14282,N_12294);
xnor UO_1670 (O_1670,N_14371,N_13719);
nor UO_1671 (O_1671,N_14693,N_13735);
xor UO_1672 (O_1672,N_13530,N_13451);
and UO_1673 (O_1673,N_13010,N_12539);
nor UO_1674 (O_1674,N_12471,N_12478);
and UO_1675 (O_1675,N_12452,N_13017);
and UO_1676 (O_1676,N_12857,N_12366);
xnor UO_1677 (O_1677,N_13816,N_14430);
xor UO_1678 (O_1678,N_14959,N_12910);
nor UO_1679 (O_1679,N_13622,N_13733);
and UO_1680 (O_1680,N_12305,N_12814);
or UO_1681 (O_1681,N_14540,N_13458);
nand UO_1682 (O_1682,N_14208,N_13604);
or UO_1683 (O_1683,N_13482,N_14846);
or UO_1684 (O_1684,N_13060,N_12722);
or UO_1685 (O_1685,N_13410,N_13920);
nand UO_1686 (O_1686,N_12186,N_14965);
and UO_1687 (O_1687,N_13126,N_13227);
nor UO_1688 (O_1688,N_12762,N_14840);
and UO_1689 (O_1689,N_12574,N_12496);
or UO_1690 (O_1690,N_13428,N_13337);
or UO_1691 (O_1691,N_13578,N_14870);
xor UO_1692 (O_1692,N_13558,N_12453);
or UO_1693 (O_1693,N_14072,N_12771);
and UO_1694 (O_1694,N_12363,N_12010);
or UO_1695 (O_1695,N_13593,N_14195);
and UO_1696 (O_1696,N_14121,N_13796);
xnor UO_1697 (O_1697,N_14910,N_12252);
nand UO_1698 (O_1698,N_14647,N_14188);
and UO_1699 (O_1699,N_14584,N_12267);
nand UO_1700 (O_1700,N_12299,N_14134);
and UO_1701 (O_1701,N_12272,N_14443);
and UO_1702 (O_1702,N_12533,N_12354);
and UO_1703 (O_1703,N_12340,N_13390);
and UO_1704 (O_1704,N_14758,N_14678);
or UO_1705 (O_1705,N_13159,N_14752);
xor UO_1706 (O_1706,N_14027,N_12738);
nor UO_1707 (O_1707,N_12056,N_12728);
nand UO_1708 (O_1708,N_12471,N_13174);
or UO_1709 (O_1709,N_14204,N_13409);
xor UO_1710 (O_1710,N_12765,N_14324);
or UO_1711 (O_1711,N_14341,N_13473);
xnor UO_1712 (O_1712,N_14363,N_12946);
xnor UO_1713 (O_1713,N_14826,N_14212);
or UO_1714 (O_1714,N_13994,N_14859);
nor UO_1715 (O_1715,N_14780,N_14025);
xor UO_1716 (O_1716,N_12226,N_12453);
nor UO_1717 (O_1717,N_12519,N_14913);
nor UO_1718 (O_1718,N_12273,N_12333);
or UO_1719 (O_1719,N_13260,N_14737);
nand UO_1720 (O_1720,N_14793,N_14178);
nand UO_1721 (O_1721,N_14138,N_12345);
nor UO_1722 (O_1722,N_13656,N_13197);
or UO_1723 (O_1723,N_12556,N_12330);
nand UO_1724 (O_1724,N_14206,N_14109);
nand UO_1725 (O_1725,N_12827,N_12545);
or UO_1726 (O_1726,N_13186,N_12991);
nand UO_1727 (O_1727,N_14981,N_12180);
or UO_1728 (O_1728,N_12644,N_12655);
and UO_1729 (O_1729,N_12216,N_12775);
or UO_1730 (O_1730,N_13989,N_14239);
or UO_1731 (O_1731,N_14328,N_14837);
nand UO_1732 (O_1732,N_12901,N_14476);
nand UO_1733 (O_1733,N_13273,N_12711);
nand UO_1734 (O_1734,N_13688,N_14985);
or UO_1735 (O_1735,N_12989,N_14290);
nor UO_1736 (O_1736,N_13090,N_14194);
and UO_1737 (O_1737,N_13696,N_14771);
xnor UO_1738 (O_1738,N_12965,N_13603);
and UO_1739 (O_1739,N_12852,N_13008);
nor UO_1740 (O_1740,N_12986,N_14614);
nand UO_1741 (O_1741,N_12295,N_14176);
nand UO_1742 (O_1742,N_13494,N_12735);
and UO_1743 (O_1743,N_12364,N_13098);
or UO_1744 (O_1744,N_12071,N_13763);
xor UO_1745 (O_1745,N_12689,N_12594);
nand UO_1746 (O_1746,N_14891,N_12856);
xor UO_1747 (O_1747,N_14254,N_13698);
and UO_1748 (O_1748,N_12395,N_14988);
nor UO_1749 (O_1749,N_14747,N_13261);
and UO_1750 (O_1750,N_13537,N_13150);
nor UO_1751 (O_1751,N_14202,N_13834);
or UO_1752 (O_1752,N_14204,N_12280);
xnor UO_1753 (O_1753,N_14909,N_14231);
and UO_1754 (O_1754,N_12510,N_12087);
and UO_1755 (O_1755,N_13949,N_12305);
nor UO_1756 (O_1756,N_13399,N_13166);
or UO_1757 (O_1757,N_14998,N_14301);
xor UO_1758 (O_1758,N_14487,N_14377);
xor UO_1759 (O_1759,N_14360,N_12862);
or UO_1760 (O_1760,N_13881,N_12631);
and UO_1761 (O_1761,N_12067,N_12500);
nor UO_1762 (O_1762,N_12935,N_13001);
nor UO_1763 (O_1763,N_14894,N_13061);
or UO_1764 (O_1764,N_14059,N_13934);
or UO_1765 (O_1765,N_14728,N_14559);
nand UO_1766 (O_1766,N_14023,N_14719);
or UO_1767 (O_1767,N_12168,N_12473);
xnor UO_1768 (O_1768,N_13887,N_12301);
nand UO_1769 (O_1769,N_12596,N_13238);
or UO_1770 (O_1770,N_14631,N_13909);
nor UO_1771 (O_1771,N_13991,N_13821);
nand UO_1772 (O_1772,N_12956,N_13843);
xor UO_1773 (O_1773,N_13104,N_14725);
nor UO_1774 (O_1774,N_12725,N_13257);
and UO_1775 (O_1775,N_12001,N_12273);
or UO_1776 (O_1776,N_14311,N_12623);
nand UO_1777 (O_1777,N_12091,N_14679);
and UO_1778 (O_1778,N_14673,N_14803);
and UO_1779 (O_1779,N_12882,N_14445);
nand UO_1780 (O_1780,N_12358,N_14002);
xor UO_1781 (O_1781,N_12190,N_13968);
or UO_1782 (O_1782,N_13188,N_13895);
and UO_1783 (O_1783,N_12095,N_13079);
nor UO_1784 (O_1784,N_12842,N_12285);
nand UO_1785 (O_1785,N_12455,N_12484);
or UO_1786 (O_1786,N_12125,N_12401);
nand UO_1787 (O_1787,N_14442,N_14478);
xor UO_1788 (O_1788,N_13767,N_14550);
and UO_1789 (O_1789,N_13780,N_13228);
nor UO_1790 (O_1790,N_13983,N_14734);
and UO_1791 (O_1791,N_12281,N_13151);
or UO_1792 (O_1792,N_12398,N_13794);
or UO_1793 (O_1793,N_13760,N_12989);
and UO_1794 (O_1794,N_12802,N_13064);
xor UO_1795 (O_1795,N_12710,N_14219);
and UO_1796 (O_1796,N_14877,N_13725);
or UO_1797 (O_1797,N_13397,N_12496);
nand UO_1798 (O_1798,N_12411,N_13738);
nand UO_1799 (O_1799,N_12403,N_13822);
nand UO_1800 (O_1800,N_12791,N_13009);
xor UO_1801 (O_1801,N_14342,N_14504);
and UO_1802 (O_1802,N_14567,N_12820);
nor UO_1803 (O_1803,N_12944,N_14260);
or UO_1804 (O_1804,N_12003,N_14177);
nor UO_1805 (O_1805,N_13938,N_13528);
and UO_1806 (O_1806,N_13804,N_14712);
or UO_1807 (O_1807,N_12016,N_14942);
nand UO_1808 (O_1808,N_14398,N_13766);
nand UO_1809 (O_1809,N_13740,N_12196);
xor UO_1810 (O_1810,N_13036,N_13170);
or UO_1811 (O_1811,N_12438,N_12708);
xnor UO_1812 (O_1812,N_13917,N_13898);
nor UO_1813 (O_1813,N_13698,N_14748);
nor UO_1814 (O_1814,N_12323,N_12897);
or UO_1815 (O_1815,N_13787,N_14121);
xnor UO_1816 (O_1816,N_14712,N_14523);
nand UO_1817 (O_1817,N_13908,N_12518);
nand UO_1818 (O_1818,N_14487,N_12057);
xor UO_1819 (O_1819,N_14015,N_14901);
xnor UO_1820 (O_1820,N_12482,N_12836);
nand UO_1821 (O_1821,N_13747,N_14276);
xor UO_1822 (O_1822,N_12149,N_12646);
xnor UO_1823 (O_1823,N_14215,N_12611);
nand UO_1824 (O_1824,N_14567,N_13488);
xor UO_1825 (O_1825,N_13315,N_13194);
xor UO_1826 (O_1826,N_14051,N_12452);
xnor UO_1827 (O_1827,N_14578,N_13971);
or UO_1828 (O_1828,N_12980,N_13580);
nor UO_1829 (O_1829,N_14287,N_14637);
nor UO_1830 (O_1830,N_13878,N_13123);
or UO_1831 (O_1831,N_13857,N_14175);
xor UO_1832 (O_1832,N_14802,N_14837);
xnor UO_1833 (O_1833,N_14598,N_14536);
nand UO_1834 (O_1834,N_14834,N_13629);
or UO_1835 (O_1835,N_12256,N_13937);
or UO_1836 (O_1836,N_13310,N_13138);
or UO_1837 (O_1837,N_14775,N_14503);
nor UO_1838 (O_1838,N_14513,N_12420);
nor UO_1839 (O_1839,N_14767,N_13936);
or UO_1840 (O_1840,N_12785,N_12143);
xnor UO_1841 (O_1841,N_12712,N_14932);
and UO_1842 (O_1842,N_12625,N_13527);
or UO_1843 (O_1843,N_13473,N_13513);
nand UO_1844 (O_1844,N_12228,N_12306);
nor UO_1845 (O_1845,N_14088,N_12103);
xnor UO_1846 (O_1846,N_14215,N_12419);
and UO_1847 (O_1847,N_14957,N_14597);
nor UO_1848 (O_1848,N_13995,N_13590);
nor UO_1849 (O_1849,N_13294,N_13119);
nor UO_1850 (O_1850,N_14899,N_12160);
nand UO_1851 (O_1851,N_12969,N_12959);
xnor UO_1852 (O_1852,N_13859,N_14199);
nor UO_1853 (O_1853,N_14366,N_13738);
or UO_1854 (O_1854,N_12765,N_12763);
and UO_1855 (O_1855,N_13851,N_12313);
nor UO_1856 (O_1856,N_14451,N_12923);
or UO_1857 (O_1857,N_12999,N_12559);
nand UO_1858 (O_1858,N_14098,N_14798);
nor UO_1859 (O_1859,N_14742,N_12715);
xor UO_1860 (O_1860,N_12164,N_12680);
and UO_1861 (O_1861,N_12152,N_12755);
or UO_1862 (O_1862,N_13897,N_12816);
nor UO_1863 (O_1863,N_14767,N_12562);
nand UO_1864 (O_1864,N_13461,N_12379);
and UO_1865 (O_1865,N_12016,N_14442);
nand UO_1866 (O_1866,N_12280,N_12100);
nand UO_1867 (O_1867,N_14681,N_14588);
xor UO_1868 (O_1868,N_12729,N_12322);
and UO_1869 (O_1869,N_13875,N_12143);
xnor UO_1870 (O_1870,N_14257,N_13138);
and UO_1871 (O_1871,N_13533,N_14702);
nand UO_1872 (O_1872,N_12699,N_13478);
nor UO_1873 (O_1873,N_12414,N_14551);
or UO_1874 (O_1874,N_12064,N_12136);
nand UO_1875 (O_1875,N_13986,N_12000);
nand UO_1876 (O_1876,N_14339,N_12656);
nor UO_1877 (O_1877,N_12015,N_12661);
or UO_1878 (O_1878,N_13276,N_12166);
xnor UO_1879 (O_1879,N_13815,N_12466);
and UO_1880 (O_1880,N_12944,N_12874);
or UO_1881 (O_1881,N_14654,N_14594);
nand UO_1882 (O_1882,N_13874,N_14046);
xnor UO_1883 (O_1883,N_13791,N_12740);
xnor UO_1884 (O_1884,N_12395,N_12625);
xor UO_1885 (O_1885,N_12415,N_14381);
xor UO_1886 (O_1886,N_12468,N_14657);
and UO_1887 (O_1887,N_14541,N_12527);
or UO_1888 (O_1888,N_14424,N_13649);
nand UO_1889 (O_1889,N_14322,N_13659);
nand UO_1890 (O_1890,N_12283,N_14028);
and UO_1891 (O_1891,N_13800,N_12701);
nor UO_1892 (O_1892,N_12023,N_13761);
and UO_1893 (O_1893,N_12435,N_12585);
or UO_1894 (O_1894,N_12170,N_12717);
nand UO_1895 (O_1895,N_13117,N_14863);
xor UO_1896 (O_1896,N_12082,N_14154);
xor UO_1897 (O_1897,N_14099,N_12305);
and UO_1898 (O_1898,N_12390,N_12590);
and UO_1899 (O_1899,N_14370,N_13108);
nor UO_1900 (O_1900,N_14645,N_13641);
nor UO_1901 (O_1901,N_14312,N_14497);
nand UO_1902 (O_1902,N_13300,N_13260);
xnor UO_1903 (O_1903,N_12828,N_14083);
nor UO_1904 (O_1904,N_14211,N_12353);
and UO_1905 (O_1905,N_14633,N_14784);
xnor UO_1906 (O_1906,N_13546,N_13244);
xnor UO_1907 (O_1907,N_13888,N_12922);
or UO_1908 (O_1908,N_12628,N_14449);
nand UO_1909 (O_1909,N_13754,N_14462);
nor UO_1910 (O_1910,N_13940,N_12028);
and UO_1911 (O_1911,N_14216,N_13465);
or UO_1912 (O_1912,N_13189,N_13198);
xnor UO_1913 (O_1913,N_14098,N_13574);
nor UO_1914 (O_1914,N_13883,N_12989);
and UO_1915 (O_1915,N_13236,N_12347);
and UO_1916 (O_1916,N_14448,N_13488);
nand UO_1917 (O_1917,N_12818,N_13017);
nor UO_1918 (O_1918,N_13830,N_14981);
or UO_1919 (O_1919,N_13219,N_12197);
xor UO_1920 (O_1920,N_12316,N_13273);
or UO_1921 (O_1921,N_13186,N_12669);
and UO_1922 (O_1922,N_12541,N_14365);
and UO_1923 (O_1923,N_13087,N_14469);
xor UO_1924 (O_1924,N_14688,N_12609);
or UO_1925 (O_1925,N_14520,N_14268);
and UO_1926 (O_1926,N_12618,N_13155);
and UO_1927 (O_1927,N_14258,N_13835);
nand UO_1928 (O_1928,N_12828,N_13297);
or UO_1929 (O_1929,N_14096,N_14961);
or UO_1930 (O_1930,N_14007,N_13971);
or UO_1931 (O_1931,N_12932,N_13507);
nand UO_1932 (O_1932,N_14097,N_14669);
or UO_1933 (O_1933,N_13301,N_14725);
and UO_1934 (O_1934,N_13757,N_13242);
nor UO_1935 (O_1935,N_12719,N_13165);
nor UO_1936 (O_1936,N_14234,N_12396);
nor UO_1937 (O_1937,N_14241,N_14985);
nor UO_1938 (O_1938,N_14067,N_12131);
and UO_1939 (O_1939,N_12460,N_12956);
or UO_1940 (O_1940,N_14433,N_12898);
nor UO_1941 (O_1941,N_14179,N_12358);
and UO_1942 (O_1942,N_14805,N_13959);
or UO_1943 (O_1943,N_12053,N_14775);
xor UO_1944 (O_1944,N_13201,N_14735);
or UO_1945 (O_1945,N_13171,N_14165);
nand UO_1946 (O_1946,N_13685,N_12926);
and UO_1947 (O_1947,N_14678,N_12355);
nand UO_1948 (O_1948,N_14640,N_12403);
xor UO_1949 (O_1949,N_14684,N_13733);
and UO_1950 (O_1950,N_14898,N_13452);
and UO_1951 (O_1951,N_14907,N_14934);
nor UO_1952 (O_1952,N_12345,N_14314);
and UO_1953 (O_1953,N_14405,N_13555);
and UO_1954 (O_1954,N_13440,N_14102);
nor UO_1955 (O_1955,N_13095,N_14521);
nand UO_1956 (O_1956,N_13292,N_13275);
xor UO_1957 (O_1957,N_13223,N_13932);
nor UO_1958 (O_1958,N_14073,N_13188);
or UO_1959 (O_1959,N_13119,N_12731);
and UO_1960 (O_1960,N_12221,N_14042);
xor UO_1961 (O_1961,N_12975,N_12574);
xor UO_1962 (O_1962,N_13120,N_14002);
nand UO_1963 (O_1963,N_13475,N_12983);
or UO_1964 (O_1964,N_14825,N_14208);
or UO_1965 (O_1965,N_13801,N_14827);
nor UO_1966 (O_1966,N_14903,N_12833);
nor UO_1967 (O_1967,N_12863,N_12401);
nor UO_1968 (O_1968,N_14301,N_14549);
nor UO_1969 (O_1969,N_12715,N_14667);
nand UO_1970 (O_1970,N_13302,N_13097);
xor UO_1971 (O_1971,N_13137,N_12164);
xor UO_1972 (O_1972,N_13216,N_14403);
or UO_1973 (O_1973,N_12340,N_14560);
nor UO_1974 (O_1974,N_14469,N_13899);
nor UO_1975 (O_1975,N_13066,N_12522);
nor UO_1976 (O_1976,N_14732,N_12089);
and UO_1977 (O_1977,N_12946,N_12215);
or UO_1978 (O_1978,N_13432,N_12007);
or UO_1979 (O_1979,N_13530,N_14216);
nor UO_1980 (O_1980,N_14016,N_14306);
nor UO_1981 (O_1981,N_13750,N_13168);
and UO_1982 (O_1982,N_12454,N_12601);
and UO_1983 (O_1983,N_14652,N_13086);
xnor UO_1984 (O_1984,N_12521,N_13440);
and UO_1985 (O_1985,N_12083,N_14526);
nand UO_1986 (O_1986,N_13132,N_12660);
xor UO_1987 (O_1987,N_12822,N_13334);
nor UO_1988 (O_1988,N_13713,N_13573);
nor UO_1989 (O_1989,N_12360,N_14357);
nand UO_1990 (O_1990,N_13161,N_13538);
nand UO_1991 (O_1991,N_14591,N_12340);
and UO_1992 (O_1992,N_13140,N_14916);
nor UO_1993 (O_1993,N_14745,N_12371);
or UO_1994 (O_1994,N_14001,N_13270);
nor UO_1995 (O_1995,N_12482,N_12543);
xor UO_1996 (O_1996,N_14371,N_12289);
xnor UO_1997 (O_1997,N_13055,N_14523);
or UO_1998 (O_1998,N_12076,N_12912);
and UO_1999 (O_1999,N_12918,N_14916);
endmodule