module basic_500_3000_500_15_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_266,In_201);
and U1 (N_1,In_339,In_492);
nor U2 (N_2,In_182,In_471);
nand U3 (N_3,In_64,In_276);
or U4 (N_4,In_119,In_352);
nand U5 (N_5,In_149,In_204);
and U6 (N_6,In_130,In_245);
nor U7 (N_7,In_9,In_242);
and U8 (N_8,In_141,In_158);
nor U9 (N_9,In_137,In_333);
and U10 (N_10,In_95,In_486);
and U11 (N_11,In_224,In_360);
nor U12 (N_12,In_319,In_332);
and U13 (N_13,In_7,In_381);
and U14 (N_14,In_343,In_449);
and U15 (N_15,In_498,In_465);
nor U16 (N_16,In_177,In_372);
and U17 (N_17,In_226,In_402);
nand U18 (N_18,In_363,In_349);
nand U19 (N_19,In_356,In_35);
and U20 (N_20,In_416,In_52);
nand U21 (N_21,In_404,In_344);
nor U22 (N_22,In_112,In_12);
nand U23 (N_23,In_274,In_209);
and U24 (N_24,In_418,In_308);
or U25 (N_25,In_213,In_70);
or U26 (N_26,In_268,In_73);
nor U27 (N_27,In_161,In_239);
or U28 (N_28,In_490,In_215);
nand U29 (N_29,In_179,In_432);
or U30 (N_30,In_54,In_63);
and U31 (N_31,In_85,In_285);
or U32 (N_32,In_246,In_310);
or U33 (N_33,In_167,In_21);
nand U34 (N_34,In_19,In_173);
and U35 (N_35,In_292,In_263);
nand U36 (N_36,In_261,In_45);
nand U37 (N_37,In_106,In_10);
or U38 (N_38,In_155,In_89);
and U39 (N_39,In_484,In_313);
or U40 (N_40,In_474,In_190);
and U41 (N_41,In_244,In_34);
or U42 (N_42,In_176,In_139);
nand U43 (N_43,In_377,In_168);
nand U44 (N_44,In_369,In_468);
nor U45 (N_45,In_279,In_16);
nand U46 (N_46,In_288,In_162);
or U47 (N_47,In_87,In_307);
nor U48 (N_48,In_271,In_116);
or U49 (N_49,In_304,In_39);
and U50 (N_50,In_75,In_353);
and U51 (N_51,In_227,In_248);
and U52 (N_52,In_145,In_278);
or U53 (N_53,In_23,In_11);
nor U54 (N_54,In_380,In_131);
nor U55 (N_55,In_294,In_76);
or U56 (N_56,In_488,In_305);
and U57 (N_57,In_107,In_154);
nor U58 (N_58,In_97,In_440);
nand U59 (N_59,In_121,In_125);
nand U60 (N_60,In_118,In_36);
nor U61 (N_61,In_122,In_96);
nand U62 (N_62,In_153,In_311);
and U63 (N_63,In_175,In_126);
nand U64 (N_64,In_216,In_20);
or U65 (N_65,In_152,In_303);
nand U66 (N_66,In_456,In_479);
nand U67 (N_67,In_495,In_299);
or U68 (N_68,In_229,In_396);
or U69 (N_69,In_291,In_234);
nor U70 (N_70,In_384,In_426);
or U71 (N_71,In_337,In_79);
or U72 (N_72,In_267,In_264);
or U73 (N_73,In_389,In_413);
nand U74 (N_74,In_14,In_6);
nor U75 (N_75,In_25,In_351);
nand U76 (N_76,In_364,In_58);
and U77 (N_77,In_342,In_482);
and U78 (N_78,In_188,In_448);
nor U79 (N_79,In_71,In_287);
or U80 (N_80,In_217,In_200);
nand U81 (N_81,In_487,In_460);
nor U82 (N_82,In_24,In_198);
nand U83 (N_83,In_346,In_15);
nand U84 (N_84,In_83,In_476);
nor U85 (N_85,In_38,In_373);
or U86 (N_86,In_314,In_454);
or U87 (N_87,In_408,In_0);
or U88 (N_88,In_262,In_214);
and U89 (N_89,In_283,In_273);
and U90 (N_90,In_133,In_235);
and U91 (N_91,In_388,In_443);
and U92 (N_92,In_336,In_140);
and U93 (N_93,In_221,In_124);
or U94 (N_94,In_48,In_347);
and U95 (N_95,In_420,In_123);
and U96 (N_96,In_453,In_27);
nand U97 (N_97,In_113,In_406);
nor U98 (N_98,In_499,In_483);
and U99 (N_99,In_382,In_451);
nand U100 (N_100,In_378,In_357);
and U101 (N_101,In_407,In_47);
nor U102 (N_102,In_324,In_435);
nand U103 (N_103,In_187,In_361);
and U104 (N_104,In_370,In_400);
nor U105 (N_105,In_391,In_290);
and U106 (N_106,In_318,In_461);
nand U107 (N_107,In_22,In_60);
and U108 (N_108,In_441,In_386);
or U109 (N_109,In_192,In_210);
or U110 (N_110,In_289,In_183);
nor U111 (N_111,In_421,In_172);
or U112 (N_112,In_86,In_222);
and U113 (N_113,In_136,In_1);
nand U114 (N_114,In_254,In_419);
nor U115 (N_115,In_296,In_259);
and U116 (N_116,In_350,In_497);
or U117 (N_117,In_148,In_41);
or U118 (N_118,In_160,In_80);
nor U119 (N_119,In_258,In_146);
and U120 (N_120,In_240,In_120);
nor U121 (N_121,In_69,In_417);
and U122 (N_122,In_321,In_30);
nor U123 (N_123,In_8,In_84);
and U124 (N_124,In_197,In_395);
and U125 (N_125,In_171,In_341);
nor U126 (N_126,In_338,In_412);
nor U127 (N_127,In_206,In_286);
or U128 (N_128,In_99,In_472);
or U129 (N_129,In_67,In_383);
nor U130 (N_130,In_223,In_108);
nor U131 (N_131,In_434,In_301);
and U132 (N_132,In_142,In_496);
or U133 (N_133,In_205,In_243);
nand U134 (N_134,In_29,In_128);
or U135 (N_135,In_322,In_359);
nor U136 (N_136,In_265,In_485);
nand U137 (N_137,In_98,In_94);
or U138 (N_138,In_439,In_379);
or U139 (N_139,In_191,In_480);
nand U140 (N_140,In_320,In_316);
and U141 (N_141,In_376,In_132);
or U142 (N_142,In_13,In_199);
nor U143 (N_143,In_65,In_457);
nor U144 (N_144,In_51,In_50);
nor U145 (N_145,In_452,In_428);
and U146 (N_146,In_230,In_427);
nor U147 (N_147,In_280,In_170);
and U148 (N_148,In_101,In_247);
nor U149 (N_149,In_77,In_117);
nor U150 (N_150,In_163,In_255);
nor U151 (N_151,In_411,In_478);
nand U152 (N_152,In_257,In_473);
nand U153 (N_153,In_270,In_447);
nor U154 (N_154,In_241,In_423);
nand U155 (N_155,In_57,In_147);
or U156 (N_156,In_277,In_127);
nor U157 (N_157,In_340,In_202);
nand U158 (N_158,In_88,In_165);
and U159 (N_159,In_459,In_367);
and U160 (N_160,In_32,In_387);
or U161 (N_161,In_348,In_256);
nand U162 (N_162,In_401,In_103);
nand U163 (N_163,In_82,In_233);
nor U164 (N_164,In_220,In_463);
nor U165 (N_165,In_135,In_178);
and U166 (N_166,In_462,In_18);
nand U167 (N_167,In_231,In_138);
or U168 (N_168,In_225,In_374);
nand U169 (N_169,In_104,In_92);
nand U170 (N_170,In_150,In_253);
or U171 (N_171,In_212,In_385);
and U172 (N_172,In_298,In_46);
nor U173 (N_173,In_437,In_72);
or U174 (N_174,In_325,In_189);
nor U175 (N_175,In_129,In_393);
or U176 (N_176,In_477,In_66);
or U177 (N_177,In_424,In_326);
or U178 (N_178,In_442,In_328);
nor U179 (N_179,In_260,In_309);
nor U180 (N_180,In_284,In_470);
or U181 (N_181,In_110,In_429);
nor U182 (N_182,In_371,In_269);
nand U183 (N_183,In_203,In_114);
or U184 (N_184,In_466,In_446);
or U185 (N_185,In_157,In_397);
nor U186 (N_186,In_93,In_185);
nand U187 (N_187,In_293,In_390);
or U188 (N_188,In_433,In_81);
and U189 (N_189,In_151,In_315);
and U190 (N_190,In_394,In_4);
nor U191 (N_191,In_491,In_272);
and U192 (N_192,In_102,In_415);
and U193 (N_193,In_392,In_2);
or U194 (N_194,In_410,In_481);
or U195 (N_195,In_414,In_55);
or U196 (N_196,In_458,In_232);
nand U197 (N_197,In_475,In_174);
nor U198 (N_198,In_180,In_317);
nand U199 (N_199,In_219,In_399);
nand U200 (N_200,In_143,In_375);
xor U201 (N_201,N_40,N_61);
or U202 (N_202,In_444,In_78);
nor U203 (N_203,N_96,In_31);
and U204 (N_204,N_84,N_182);
and U205 (N_205,N_21,In_252);
or U206 (N_206,N_122,N_11);
or U207 (N_207,In_464,N_48);
nand U208 (N_208,N_116,In_105);
nor U209 (N_209,N_136,In_207);
nor U210 (N_210,N_16,In_494);
nand U211 (N_211,In_33,In_403);
or U212 (N_212,N_4,N_89);
or U213 (N_213,N_197,In_312);
or U214 (N_214,In_144,N_8);
and U215 (N_215,In_345,In_302);
or U216 (N_216,N_105,N_106);
nor U217 (N_217,In_208,In_237);
and U218 (N_218,N_100,N_99);
or U219 (N_219,N_173,In_489);
and U220 (N_220,In_430,N_74);
or U221 (N_221,N_193,N_162);
or U222 (N_222,N_196,In_450);
xnor U223 (N_223,N_157,N_109);
or U224 (N_224,N_194,N_160);
or U225 (N_225,N_169,N_185);
or U226 (N_226,N_0,N_86);
nor U227 (N_227,N_101,N_124);
and U228 (N_228,N_198,In_368);
and U229 (N_229,In_354,In_398);
nor U230 (N_230,N_90,In_250);
or U231 (N_231,In_211,In_295);
and U232 (N_232,N_46,In_335);
and U233 (N_233,N_85,In_358);
nand U234 (N_234,In_61,In_37);
and U235 (N_235,N_186,N_195);
or U236 (N_236,N_123,N_117);
nand U237 (N_237,N_143,In_196);
or U238 (N_238,In_228,In_44);
and U239 (N_239,In_329,N_161);
nor U240 (N_240,N_130,N_95);
nor U241 (N_241,In_445,N_28);
or U242 (N_242,N_43,N_175);
nor U243 (N_243,N_37,In_366);
nand U244 (N_244,N_35,N_171);
nand U245 (N_245,N_149,N_66);
or U246 (N_246,N_180,In_181);
nor U247 (N_247,In_467,In_282);
and U248 (N_248,N_57,N_164);
nor U249 (N_249,N_159,N_153);
or U250 (N_250,In_323,N_49);
or U251 (N_251,N_55,N_148);
nor U252 (N_252,In_238,N_73);
or U253 (N_253,N_77,N_140);
nor U254 (N_254,N_1,N_27);
nand U255 (N_255,In_109,In_431);
and U256 (N_256,N_44,N_151);
nand U257 (N_257,In_195,N_62);
or U258 (N_258,N_165,N_115);
and U259 (N_259,In_43,N_154);
or U260 (N_260,N_181,In_194);
nor U261 (N_261,In_331,In_281);
and U262 (N_262,In_455,N_91);
and U263 (N_263,In_59,In_355);
nor U264 (N_264,N_125,N_80);
nor U265 (N_265,N_63,N_126);
nor U266 (N_266,In_17,N_15);
nor U267 (N_267,N_7,In_362);
nor U268 (N_268,N_150,N_104);
nor U269 (N_269,In_306,N_59);
nor U270 (N_270,In_251,N_79);
or U271 (N_271,N_112,N_179);
or U272 (N_272,N_70,N_135);
and U273 (N_273,N_120,N_18);
and U274 (N_274,N_17,N_199);
or U275 (N_275,N_118,N_137);
and U276 (N_276,N_19,N_92);
and U277 (N_277,N_107,N_142);
or U278 (N_278,N_158,N_52);
nor U279 (N_279,In_425,In_236);
nor U280 (N_280,N_111,N_178);
nor U281 (N_281,N_75,N_114);
nor U282 (N_282,In_438,N_108);
or U283 (N_283,In_164,In_184);
nand U284 (N_284,N_53,N_183);
and U285 (N_285,In_193,N_192);
nor U286 (N_286,N_139,N_129);
and U287 (N_287,In_365,In_28);
nor U288 (N_288,N_134,N_132);
and U289 (N_289,N_94,N_56);
nor U290 (N_290,In_469,In_186);
nand U291 (N_291,N_10,N_22);
nor U292 (N_292,In_111,N_102);
nand U293 (N_293,N_172,In_330);
and U294 (N_294,In_493,N_23);
nand U295 (N_295,N_50,N_38);
nand U296 (N_296,N_36,N_6);
nand U297 (N_297,N_131,N_128);
nand U298 (N_298,N_88,N_145);
nand U299 (N_299,N_42,N_127);
nor U300 (N_300,N_144,N_146);
nand U301 (N_301,N_163,N_110);
nand U302 (N_302,N_152,N_168);
nand U303 (N_303,N_51,N_174);
nand U304 (N_304,N_47,N_26);
or U305 (N_305,N_54,N_147);
or U306 (N_306,N_176,N_20);
nand U307 (N_307,In_40,N_58);
and U308 (N_308,N_121,N_5);
nor U309 (N_309,In_56,In_275);
or U310 (N_310,N_113,In_90);
nor U311 (N_311,N_76,N_93);
or U312 (N_312,In_405,In_3);
and U313 (N_313,N_2,In_169);
and U314 (N_314,N_82,N_103);
or U315 (N_315,N_29,N_14);
nand U316 (N_316,In_134,In_218);
nor U317 (N_317,N_87,N_177);
or U318 (N_318,N_81,N_187);
and U319 (N_319,In_91,In_115);
nor U320 (N_320,N_3,N_71);
nand U321 (N_321,N_69,N_65);
nor U322 (N_322,N_119,N_138);
and U323 (N_323,N_24,In_159);
and U324 (N_324,N_68,N_67);
or U325 (N_325,N_155,N_133);
and U326 (N_326,N_184,N_83);
nor U327 (N_327,N_9,N_31);
or U328 (N_328,N_190,N_72);
and U329 (N_329,N_32,In_297);
nand U330 (N_330,N_41,In_166);
or U331 (N_331,N_13,In_5);
nor U332 (N_332,N_30,In_249);
nor U333 (N_333,In_334,N_78);
or U334 (N_334,N_34,N_170);
or U335 (N_335,N_156,N_64);
or U336 (N_336,N_12,In_327);
nand U337 (N_337,In_26,N_97);
nand U338 (N_338,N_33,N_167);
nor U339 (N_339,In_42,In_436);
or U340 (N_340,In_100,In_74);
and U341 (N_341,N_166,In_53);
nor U342 (N_342,N_188,In_422);
and U343 (N_343,N_98,In_49);
nand U344 (N_344,In_409,In_62);
nor U345 (N_345,N_189,N_191);
nor U346 (N_346,N_60,N_45);
nor U347 (N_347,In_300,In_156);
nor U348 (N_348,N_25,N_141);
or U349 (N_349,In_68,N_39);
nand U350 (N_350,In_186,N_42);
or U351 (N_351,In_323,N_23);
nor U352 (N_352,N_179,N_20);
or U353 (N_353,N_153,N_105);
nor U354 (N_354,N_63,In_282);
or U355 (N_355,N_134,N_169);
nor U356 (N_356,N_176,N_141);
or U357 (N_357,N_107,In_17);
nor U358 (N_358,In_181,N_94);
nand U359 (N_359,N_103,In_403);
or U360 (N_360,In_297,In_166);
nand U361 (N_361,N_157,N_60);
or U362 (N_362,N_61,N_123);
nor U363 (N_363,N_174,In_156);
or U364 (N_364,In_405,N_196);
or U365 (N_365,N_9,N_173);
xnor U366 (N_366,N_187,N_58);
nor U367 (N_367,In_422,N_8);
and U368 (N_368,N_125,In_42);
or U369 (N_369,N_123,N_151);
nand U370 (N_370,In_237,N_32);
nor U371 (N_371,In_334,N_47);
nand U372 (N_372,N_182,N_150);
or U373 (N_373,In_194,In_62);
nand U374 (N_374,In_105,In_115);
and U375 (N_375,N_148,In_49);
or U376 (N_376,In_78,N_6);
or U377 (N_377,N_10,In_431);
or U378 (N_378,N_30,N_167);
and U379 (N_379,N_10,N_119);
or U380 (N_380,In_90,In_44);
and U381 (N_381,N_144,N_158);
nand U382 (N_382,N_22,In_281);
or U383 (N_383,N_10,In_455);
or U384 (N_384,N_171,In_275);
or U385 (N_385,N_139,N_53);
or U386 (N_386,N_27,N_103);
and U387 (N_387,N_181,N_86);
xor U388 (N_388,In_74,N_162);
and U389 (N_389,In_455,N_188);
and U390 (N_390,N_191,N_47);
or U391 (N_391,N_80,N_83);
and U392 (N_392,In_43,N_116);
and U393 (N_393,N_130,N_60);
and U394 (N_394,N_196,N_189);
and U395 (N_395,N_188,N_18);
nand U396 (N_396,N_130,N_42);
nor U397 (N_397,In_375,N_13);
nor U398 (N_398,N_70,N_141);
and U399 (N_399,N_79,N_183);
and U400 (N_400,N_270,N_237);
nand U401 (N_401,N_348,N_368);
nand U402 (N_402,N_371,N_232);
and U403 (N_403,N_291,N_255);
nor U404 (N_404,N_385,N_256);
nor U405 (N_405,N_326,N_327);
nor U406 (N_406,N_307,N_365);
nor U407 (N_407,N_369,N_222);
nand U408 (N_408,N_393,N_304);
and U409 (N_409,N_322,N_280);
and U410 (N_410,N_357,N_258);
and U411 (N_411,N_221,N_331);
nor U412 (N_412,N_275,N_272);
or U413 (N_413,N_363,N_396);
and U414 (N_414,N_208,N_314);
and U415 (N_415,N_305,N_204);
or U416 (N_416,N_281,N_273);
or U417 (N_417,N_338,N_243);
nor U418 (N_418,N_343,N_379);
xnor U419 (N_419,N_381,N_228);
nor U420 (N_420,N_238,N_374);
and U421 (N_421,N_346,N_210);
and U422 (N_422,N_205,N_292);
nor U423 (N_423,N_220,N_310);
and U424 (N_424,N_392,N_398);
or U425 (N_425,N_341,N_278);
nand U426 (N_426,N_344,N_260);
nor U427 (N_427,N_382,N_376);
or U428 (N_428,N_325,N_388);
and U429 (N_429,N_264,N_332);
nand U430 (N_430,N_216,N_252);
or U431 (N_431,N_277,N_309);
nand U432 (N_432,N_279,N_257);
nor U433 (N_433,N_328,N_318);
nor U434 (N_434,N_362,N_370);
nor U435 (N_435,N_384,N_316);
nor U436 (N_436,N_395,N_231);
and U437 (N_437,N_321,N_387);
nand U438 (N_438,N_315,N_271);
and U439 (N_439,N_212,N_337);
nand U440 (N_440,N_364,N_367);
or U441 (N_441,N_233,N_224);
nand U442 (N_442,N_313,N_267);
or U443 (N_443,N_345,N_334);
nor U444 (N_444,N_342,N_246);
and U445 (N_445,N_223,N_356);
or U446 (N_446,N_361,N_306);
nor U447 (N_447,N_351,N_375);
nor U448 (N_448,N_300,N_248);
and U449 (N_449,N_225,N_383);
nand U450 (N_450,N_296,N_336);
nor U451 (N_451,N_299,N_399);
nor U452 (N_452,N_389,N_354);
nand U453 (N_453,N_289,N_203);
and U454 (N_454,N_377,N_261);
or U455 (N_455,N_349,N_311);
nand U456 (N_456,N_262,N_229);
nor U457 (N_457,N_380,N_303);
nor U458 (N_458,N_219,N_214);
nor U459 (N_459,N_353,N_266);
xnor U460 (N_460,N_236,N_276);
nor U461 (N_461,N_394,N_268);
nor U462 (N_462,N_359,N_298);
and U463 (N_463,N_397,N_358);
and U464 (N_464,N_373,N_372);
nand U465 (N_465,N_386,N_317);
and U466 (N_466,N_250,N_240);
and U467 (N_467,N_265,N_207);
nand U468 (N_468,N_269,N_263);
nor U469 (N_469,N_200,N_335);
and U470 (N_470,N_217,N_254);
nand U471 (N_471,N_293,N_287);
nor U472 (N_472,N_294,N_378);
and U473 (N_473,N_312,N_234);
nand U474 (N_474,N_206,N_284);
nor U475 (N_475,N_213,N_288);
or U476 (N_476,N_226,N_333);
nor U477 (N_477,N_329,N_282);
nor U478 (N_478,N_201,N_352);
nand U479 (N_479,N_259,N_347);
and U480 (N_480,N_285,N_209);
xnor U481 (N_481,N_274,N_339);
or U482 (N_482,N_290,N_320);
nor U483 (N_483,N_366,N_202);
nand U484 (N_484,N_324,N_301);
and U485 (N_485,N_245,N_355);
nand U486 (N_486,N_319,N_242);
and U487 (N_487,N_323,N_302);
nor U488 (N_488,N_295,N_211);
and U489 (N_489,N_235,N_391);
nor U490 (N_490,N_215,N_253);
nor U491 (N_491,N_308,N_230);
nand U492 (N_492,N_249,N_390);
or U493 (N_493,N_297,N_241);
and U494 (N_494,N_283,N_251);
and U495 (N_495,N_350,N_244);
nor U496 (N_496,N_330,N_286);
or U497 (N_497,N_227,N_360);
and U498 (N_498,N_340,N_218);
or U499 (N_499,N_247,N_239);
or U500 (N_500,N_206,N_257);
nand U501 (N_501,N_266,N_217);
nand U502 (N_502,N_291,N_315);
or U503 (N_503,N_330,N_250);
nand U504 (N_504,N_326,N_306);
nand U505 (N_505,N_353,N_304);
nor U506 (N_506,N_321,N_229);
and U507 (N_507,N_219,N_284);
and U508 (N_508,N_336,N_377);
nand U509 (N_509,N_256,N_282);
and U510 (N_510,N_218,N_390);
nor U511 (N_511,N_391,N_227);
nor U512 (N_512,N_217,N_207);
nor U513 (N_513,N_340,N_377);
or U514 (N_514,N_376,N_339);
or U515 (N_515,N_224,N_341);
nand U516 (N_516,N_262,N_320);
nand U517 (N_517,N_208,N_336);
nand U518 (N_518,N_226,N_362);
nor U519 (N_519,N_340,N_378);
and U520 (N_520,N_334,N_399);
nand U521 (N_521,N_398,N_334);
nor U522 (N_522,N_369,N_218);
nand U523 (N_523,N_256,N_382);
and U524 (N_524,N_292,N_218);
nand U525 (N_525,N_200,N_267);
xor U526 (N_526,N_261,N_290);
and U527 (N_527,N_221,N_353);
nand U528 (N_528,N_397,N_223);
or U529 (N_529,N_248,N_360);
or U530 (N_530,N_243,N_229);
or U531 (N_531,N_282,N_389);
and U532 (N_532,N_313,N_310);
or U533 (N_533,N_306,N_266);
or U534 (N_534,N_305,N_390);
and U535 (N_535,N_231,N_378);
and U536 (N_536,N_284,N_245);
nor U537 (N_537,N_365,N_247);
and U538 (N_538,N_385,N_302);
or U539 (N_539,N_308,N_270);
or U540 (N_540,N_303,N_274);
nand U541 (N_541,N_391,N_335);
nor U542 (N_542,N_376,N_340);
or U543 (N_543,N_205,N_322);
nor U544 (N_544,N_230,N_235);
nor U545 (N_545,N_391,N_211);
and U546 (N_546,N_360,N_390);
or U547 (N_547,N_345,N_206);
nand U548 (N_548,N_362,N_365);
and U549 (N_549,N_373,N_332);
and U550 (N_550,N_339,N_221);
nor U551 (N_551,N_340,N_309);
and U552 (N_552,N_230,N_392);
or U553 (N_553,N_296,N_358);
or U554 (N_554,N_200,N_248);
or U555 (N_555,N_324,N_304);
or U556 (N_556,N_220,N_273);
nor U557 (N_557,N_362,N_229);
and U558 (N_558,N_358,N_383);
nor U559 (N_559,N_218,N_228);
and U560 (N_560,N_367,N_273);
and U561 (N_561,N_322,N_281);
and U562 (N_562,N_320,N_232);
and U563 (N_563,N_279,N_325);
xor U564 (N_564,N_222,N_225);
nor U565 (N_565,N_364,N_318);
or U566 (N_566,N_281,N_249);
nand U567 (N_567,N_290,N_213);
nand U568 (N_568,N_275,N_318);
and U569 (N_569,N_348,N_261);
nor U570 (N_570,N_313,N_260);
and U571 (N_571,N_201,N_392);
nor U572 (N_572,N_392,N_298);
and U573 (N_573,N_366,N_226);
or U574 (N_574,N_364,N_268);
nor U575 (N_575,N_254,N_309);
or U576 (N_576,N_289,N_374);
nor U577 (N_577,N_249,N_225);
and U578 (N_578,N_328,N_305);
nor U579 (N_579,N_318,N_383);
or U580 (N_580,N_301,N_318);
nand U581 (N_581,N_397,N_236);
and U582 (N_582,N_379,N_228);
xnor U583 (N_583,N_282,N_310);
and U584 (N_584,N_263,N_255);
or U585 (N_585,N_355,N_331);
nor U586 (N_586,N_342,N_347);
nand U587 (N_587,N_248,N_277);
and U588 (N_588,N_271,N_368);
or U589 (N_589,N_225,N_393);
and U590 (N_590,N_398,N_386);
or U591 (N_591,N_277,N_274);
or U592 (N_592,N_386,N_388);
nand U593 (N_593,N_390,N_278);
and U594 (N_594,N_237,N_343);
or U595 (N_595,N_239,N_221);
or U596 (N_596,N_315,N_254);
and U597 (N_597,N_383,N_381);
nor U598 (N_598,N_358,N_331);
nand U599 (N_599,N_297,N_359);
or U600 (N_600,N_417,N_421);
nand U601 (N_601,N_592,N_545);
xor U602 (N_602,N_454,N_532);
and U603 (N_603,N_449,N_442);
nand U604 (N_604,N_461,N_511);
and U605 (N_605,N_577,N_565);
and U606 (N_606,N_587,N_572);
nand U607 (N_607,N_526,N_510);
nor U608 (N_608,N_594,N_440);
and U609 (N_609,N_401,N_561);
nor U610 (N_610,N_582,N_583);
nor U611 (N_611,N_414,N_500);
and U612 (N_612,N_405,N_567);
and U613 (N_613,N_434,N_413);
and U614 (N_614,N_408,N_426);
or U615 (N_615,N_574,N_538);
or U616 (N_616,N_578,N_451);
or U617 (N_617,N_444,N_455);
nor U618 (N_618,N_430,N_513);
or U619 (N_619,N_458,N_445);
and U620 (N_620,N_447,N_537);
nor U621 (N_621,N_584,N_424);
nand U622 (N_622,N_552,N_585);
nand U623 (N_623,N_409,N_546);
nor U624 (N_624,N_425,N_403);
nand U625 (N_625,N_496,N_450);
nor U626 (N_626,N_539,N_566);
nor U627 (N_627,N_469,N_512);
or U628 (N_628,N_576,N_488);
nor U629 (N_629,N_483,N_505);
and U630 (N_630,N_508,N_431);
and U631 (N_631,N_479,N_599);
or U632 (N_632,N_590,N_460);
nand U633 (N_633,N_453,N_547);
nand U634 (N_634,N_507,N_400);
nand U635 (N_635,N_486,N_573);
nand U636 (N_636,N_558,N_516);
nor U637 (N_637,N_501,N_553);
nor U638 (N_638,N_543,N_457);
or U639 (N_639,N_477,N_588);
nor U640 (N_640,N_465,N_517);
nand U641 (N_641,N_544,N_474);
nor U642 (N_642,N_593,N_436);
and U643 (N_643,N_597,N_491);
and U644 (N_644,N_560,N_559);
and U645 (N_645,N_522,N_598);
and U646 (N_646,N_528,N_489);
nor U647 (N_647,N_595,N_433);
or U648 (N_648,N_551,N_506);
nor U649 (N_649,N_467,N_525);
nand U650 (N_650,N_407,N_415);
nor U651 (N_651,N_523,N_487);
nor U652 (N_652,N_596,N_535);
nor U653 (N_653,N_556,N_518);
nand U654 (N_654,N_564,N_498);
or U655 (N_655,N_557,N_527);
and U656 (N_656,N_412,N_411);
or U657 (N_657,N_448,N_422);
nand U658 (N_658,N_530,N_563);
nor U659 (N_659,N_482,N_549);
and U660 (N_660,N_439,N_502);
and U661 (N_661,N_468,N_504);
or U662 (N_662,N_462,N_569);
or U663 (N_663,N_581,N_478);
nor U664 (N_664,N_446,N_438);
and U665 (N_665,N_420,N_509);
or U666 (N_666,N_463,N_586);
nor U667 (N_667,N_562,N_503);
and U668 (N_668,N_499,N_514);
nor U669 (N_669,N_437,N_418);
nand U670 (N_670,N_475,N_419);
nor U671 (N_671,N_428,N_591);
nor U672 (N_672,N_481,N_533);
or U673 (N_673,N_473,N_484);
and U674 (N_674,N_441,N_579);
or U675 (N_675,N_410,N_519);
and U676 (N_676,N_497,N_536);
and U677 (N_677,N_471,N_531);
nor U678 (N_678,N_555,N_575);
and U679 (N_679,N_520,N_541);
and U680 (N_680,N_571,N_459);
nor U681 (N_681,N_416,N_570);
or U682 (N_682,N_435,N_432);
xnor U683 (N_683,N_548,N_402);
nand U684 (N_684,N_423,N_492);
nor U685 (N_685,N_485,N_554);
and U686 (N_686,N_406,N_452);
xor U687 (N_687,N_429,N_568);
nand U688 (N_688,N_404,N_472);
and U689 (N_689,N_589,N_466);
or U690 (N_690,N_476,N_495);
nand U691 (N_691,N_550,N_480);
or U692 (N_692,N_464,N_580);
or U693 (N_693,N_529,N_443);
nor U694 (N_694,N_540,N_470);
and U695 (N_695,N_524,N_542);
or U696 (N_696,N_493,N_494);
nand U697 (N_697,N_490,N_515);
nand U698 (N_698,N_456,N_427);
nor U699 (N_699,N_534,N_521);
nor U700 (N_700,N_556,N_514);
nand U701 (N_701,N_506,N_575);
nand U702 (N_702,N_459,N_424);
xnor U703 (N_703,N_454,N_541);
and U704 (N_704,N_485,N_436);
nand U705 (N_705,N_482,N_557);
and U706 (N_706,N_505,N_434);
and U707 (N_707,N_527,N_490);
and U708 (N_708,N_554,N_458);
or U709 (N_709,N_583,N_440);
and U710 (N_710,N_482,N_426);
and U711 (N_711,N_574,N_528);
and U712 (N_712,N_503,N_450);
nand U713 (N_713,N_492,N_574);
and U714 (N_714,N_508,N_546);
nor U715 (N_715,N_405,N_562);
nand U716 (N_716,N_493,N_551);
nor U717 (N_717,N_494,N_563);
and U718 (N_718,N_405,N_443);
and U719 (N_719,N_427,N_559);
or U720 (N_720,N_531,N_566);
or U721 (N_721,N_467,N_536);
and U722 (N_722,N_528,N_592);
nand U723 (N_723,N_451,N_560);
nand U724 (N_724,N_559,N_582);
or U725 (N_725,N_581,N_527);
nand U726 (N_726,N_403,N_404);
nor U727 (N_727,N_511,N_498);
and U728 (N_728,N_428,N_526);
or U729 (N_729,N_595,N_448);
nand U730 (N_730,N_469,N_574);
nor U731 (N_731,N_439,N_426);
or U732 (N_732,N_435,N_550);
and U733 (N_733,N_546,N_570);
and U734 (N_734,N_458,N_433);
and U735 (N_735,N_417,N_535);
nand U736 (N_736,N_551,N_460);
or U737 (N_737,N_504,N_540);
and U738 (N_738,N_507,N_456);
or U739 (N_739,N_442,N_502);
nor U740 (N_740,N_539,N_423);
nor U741 (N_741,N_572,N_445);
nand U742 (N_742,N_525,N_557);
nand U743 (N_743,N_545,N_597);
nand U744 (N_744,N_495,N_515);
nand U745 (N_745,N_427,N_474);
nor U746 (N_746,N_465,N_433);
and U747 (N_747,N_408,N_412);
and U748 (N_748,N_563,N_517);
or U749 (N_749,N_423,N_529);
and U750 (N_750,N_418,N_524);
nor U751 (N_751,N_441,N_556);
nand U752 (N_752,N_491,N_490);
and U753 (N_753,N_442,N_577);
or U754 (N_754,N_493,N_451);
nand U755 (N_755,N_477,N_471);
nor U756 (N_756,N_501,N_450);
or U757 (N_757,N_431,N_529);
or U758 (N_758,N_472,N_460);
nand U759 (N_759,N_599,N_453);
or U760 (N_760,N_523,N_515);
nor U761 (N_761,N_514,N_488);
or U762 (N_762,N_568,N_577);
nand U763 (N_763,N_452,N_510);
nand U764 (N_764,N_586,N_429);
or U765 (N_765,N_402,N_421);
xnor U766 (N_766,N_480,N_531);
or U767 (N_767,N_524,N_582);
and U768 (N_768,N_593,N_519);
or U769 (N_769,N_597,N_500);
and U770 (N_770,N_554,N_470);
and U771 (N_771,N_460,N_566);
and U772 (N_772,N_589,N_432);
nand U773 (N_773,N_411,N_553);
nand U774 (N_774,N_464,N_579);
or U775 (N_775,N_512,N_400);
nor U776 (N_776,N_452,N_416);
nand U777 (N_777,N_581,N_453);
or U778 (N_778,N_548,N_432);
nand U779 (N_779,N_477,N_468);
and U780 (N_780,N_544,N_556);
or U781 (N_781,N_519,N_573);
nand U782 (N_782,N_539,N_473);
nor U783 (N_783,N_430,N_583);
nand U784 (N_784,N_529,N_561);
nor U785 (N_785,N_549,N_565);
nor U786 (N_786,N_557,N_438);
nor U787 (N_787,N_493,N_437);
or U788 (N_788,N_486,N_567);
or U789 (N_789,N_547,N_480);
and U790 (N_790,N_528,N_460);
nand U791 (N_791,N_459,N_483);
nand U792 (N_792,N_420,N_597);
and U793 (N_793,N_507,N_553);
and U794 (N_794,N_555,N_498);
xor U795 (N_795,N_597,N_596);
nand U796 (N_796,N_475,N_593);
nor U797 (N_797,N_480,N_433);
nor U798 (N_798,N_539,N_418);
nor U799 (N_799,N_533,N_546);
and U800 (N_800,N_676,N_657);
nor U801 (N_801,N_655,N_648);
nand U802 (N_802,N_663,N_662);
nor U803 (N_803,N_736,N_686);
nor U804 (N_804,N_794,N_684);
or U805 (N_805,N_720,N_704);
or U806 (N_806,N_692,N_630);
nand U807 (N_807,N_632,N_740);
or U808 (N_808,N_798,N_633);
nor U809 (N_809,N_641,N_709);
nor U810 (N_810,N_666,N_726);
and U811 (N_811,N_619,N_601);
nor U812 (N_812,N_696,N_661);
and U813 (N_813,N_734,N_658);
nor U814 (N_814,N_725,N_617);
nor U815 (N_815,N_722,N_756);
nand U816 (N_816,N_625,N_714);
nand U817 (N_817,N_644,N_693);
or U818 (N_818,N_691,N_745);
nand U819 (N_819,N_622,N_674);
nand U820 (N_820,N_653,N_636);
xor U821 (N_821,N_694,N_721);
and U822 (N_822,N_631,N_628);
or U823 (N_823,N_642,N_713);
or U824 (N_824,N_705,N_789);
and U825 (N_825,N_609,N_729);
and U826 (N_826,N_646,N_790);
or U827 (N_827,N_607,N_793);
nand U828 (N_828,N_784,N_749);
or U829 (N_829,N_618,N_690);
nand U830 (N_830,N_796,N_620);
nor U831 (N_831,N_748,N_774);
nor U832 (N_832,N_717,N_671);
nor U833 (N_833,N_652,N_660);
nor U834 (N_834,N_687,N_771);
or U835 (N_835,N_742,N_754);
nor U836 (N_836,N_635,N_664);
nand U837 (N_837,N_712,N_697);
and U838 (N_838,N_672,N_730);
nor U839 (N_839,N_627,N_768);
nand U840 (N_840,N_639,N_682);
or U841 (N_841,N_761,N_751);
or U842 (N_842,N_605,N_624);
and U843 (N_843,N_703,N_741);
or U844 (N_844,N_723,N_737);
nor U845 (N_845,N_689,N_600);
nand U846 (N_846,N_795,N_702);
nand U847 (N_847,N_763,N_728);
or U848 (N_848,N_647,N_743);
nor U849 (N_849,N_777,N_780);
and U850 (N_850,N_779,N_615);
or U851 (N_851,N_765,N_665);
nor U852 (N_852,N_782,N_602);
and U853 (N_853,N_680,N_738);
and U854 (N_854,N_612,N_699);
nor U855 (N_855,N_669,N_643);
and U856 (N_856,N_750,N_629);
nand U857 (N_857,N_711,N_688);
and U858 (N_858,N_746,N_772);
nand U859 (N_859,N_766,N_758);
and U860 (N_860,N_708,N_727);
and U861 (N_861,N_613,N_603);
nor U862 (N_862,N_606,N_659);
and U863 (N_863,N_785,N_797);
or U864 (N_864,N_753,N_733);
nor U865 (N_865,N_757,N_604);
nand U866 (N_866,N_656,N_791);
nand U867 (N_867,N_640,N_623);
and U868 (N_868,N_781,N_732);
nand U869 (N_869,N_654,N_679);
or U870 (N_870,N_770,N_773);
nand U871 (N_871,N_762,N_799);
and U872 (N_872,N_710,N_649);
nand U873 (N_873,N_616,N_621);
and U874 (N_874,N_626,N_610);
nand U875 (N_875,N_645,N_683);
or U876 (N_876,N_744,N_675);
or U877 (N_877,N_724,N_792);
and U878 (N_878,N_707,N_752);
or U879 (N_879,N_608,N_719);
and U880 (N_880,N_706,N_767);
nand U881 (N_881,N_695,N_678);
or U882 (N_882,N_685,N_716);
nor U883 (N_883,N_755,N_667);
nand U884 (N_884,N_637,N_611);
or U885 (N_885,N_759,N_787);
nor U886 (N_886,N_718,N_764);
and U887 (N_887,N_681,N_776);
and U888 (N_888,N_701,N_760);
and U889 (N_889,N_650,N_614);
or U890 (N_890,N_788,N_715);
and U891 (N_891,N_786,N_673);
or U892 (N_892,N_731,N_700);
or U893 (N_893,N_775,N_747);
nand U894 (N_894,N_769,N_634);
nor U895 (N_895,N_778,N_668);
nor U896 (N_896,N_638,N_698);
and U897 (N_897,N_651,N_739);
nand U898 (N_898,N_670,N_735);
and U899 (N_899,N_783,N_677);
nand U900 (N_900,N_721,N_673);
and U901 (N_901,N_766,N_724);
nand U902 (N_902,N_626,N_678);
nor U903 (N_903,N_650,N_675);
nor U904 (N_904,N_702,N_737);
or U905 (N_905,N_614,N_755);
or U906 (N_906,N_653,N_605);
and U907 (N_907,N_665,N_776);
or U908 (N_908,N_650,N_657);
nor U909 (N_909,N_760,N_737);
and U910 (N_910,N_641,N_607);
nor U911 (N_911,N_735,N_618);
nor U912 (N_912,N_777,N_766);
nor U913 (N_913,N_678,N_787);
nand U914 (N_914,N_607,N_650);
nor U915 (N_915,N_761,N_742);
nand U916 (N_916,N_660,N_619);
nor U917 (N_917,N_700,N_666);
nor U918 (N_918,N_799,N_606);
and U919 (N_919,N_709,N_619);
nor U920 (N_920,N_758,N_789);
or U921 (N_921,N_780,N_706);
nand U922 (N_922,N_765,N_773);
and U923 (N_923,N_783,N_700);
and U924 (N_924,N_718,N_665);
or U925 (N_925,N_786,N_707);
nand U926 (N_926,N_723,N_767);
nor U927 (N_927,N_604,N_663);
nand U928 (N_928,N_746,N_670);
and U929 (N_929,N_741,N_685);
xnor U930 (N_930,N_652,N_665);
nand U931 (N_931,N_754,N_746);
nor U932 (N_932,N_622,N_661);
nor U933 (N_933,N_739,N_747);
and U934 (N_934,N_631,N_677);
or U935 (N_935,N_771,N_602);
nand U936 (N_936,N_602,N_612);
and U937 (N_937,N_777,N_725);
and U938 (N_938,N_736,N_731);
nor U939 (N_939,N_745,N_799);
and U940 (N_940,N_711,N_736);
and U941 (N_941,N_785,N_700);
or U942 (N_942,N_700,N_649);
and U943 (N_943,N_729,N_615);
nand U944 (N_944,N_788,N_674);
or U945 (N_945,N_627,N_775);
nand U946 (N_946,N_751,N_757);
or U947 (N_947,N_687,N_793);
nand U948 (N_948,N_616,N_769);
and U949 (N_949,N_684,N_709);
or U950 (N_950,N_617,N_731);
and U951 (N_951,N_635,N_707);
and U952 (N_952,N_730,N_770);
nand U953 (N_953,N_758,N_642);
nor U954 (N_954,N_779,N_777);
and U955 (N_955,N_608,N_727);
or U956 (N_956,N_773,N_618);
or U957 (N_957,N_775,N_600);
nor U958 (N_958,N_790,N_659);
nand U959 (N_959,N_734,N_661);
and U960 (N_960,N_740,N_631);
or U961 (N_961,N_709,N_788);
or U962 (N_962,N_732,N_774);
or U963 (N_963,N_613,N_696);
nor U964 (N_964,N_798,N_728);
nor U965 (N_965,N_655,N_712);
and U966 (N_966,N_755,N_707);
or U967 (N_967,N_642,N_753);
nand U968 (N_968,N_653,N_641);
or U969 (N_969,N_617,N_757);
nand U970 (N_970,N_733,N_684);
nor U971 (N_971,N_780,N_631);
nor U972 (N_972,N_676,N_784);
nand U973 (N_973,N_731,N_798);
and U974 (N_974,N_745,N_648);
nand U975 (N_975,N_771,N_642);
and U976 (N_976,N_741,N_657);
nand U977 (N_977,N_690,N_759);
or U978 (N_978,N_712,N_680);
or U979 (N_979,N_790,N_604);
nand U980 (N_980,N_626,N_777);
nand U981 (N_981,N_676,N_656);
or U982 (N_982,N_637,N_658);
nor U983 (N_983,N_685,N_739);
and U984 (N_984,N_613,N_702);
nand U985 (N_985,N_754,N_748);
nor U986 (N_986,N_744,N_715);
and U987 (N_987,N_708,N_653);
or U988 (N_988,N_641,N_633);
xor U989 (N_989,N_776,N_784);
or U990 (N_990,N_710,N_776);
nand U991 (N_991,N_739,N_608);
nor U992 (N_992,N_715,N_683);
or U993 (N_993,N_687,N_646);
or U994 (N_994,N_678,N_730);
and U995 (N_995,N_744,N_733);
or U996 (N_996,N_691,N_736);
nor U997 (N_997,N_736,N_718);
nor U998 (N_998,N_670,N_703);
nand U999 (N_999,N_799,N_731);
or U1000 (N_1000,N_848,N_984);
nand U1001 (N_1001,N_859,N_822);
nor U1002 (N_1002,N_865,N_960);
nand U1003 (N_1003,N_947,N_910);
and U1004 (N_1004,N_810,N_897);
nor U1005 (N_1005,N_890,N_878);
and U1006 (N_1006,N_916,N_999);
or U1007 (N_1007,N_800,N_934);
nand U1008 (N_1008,N_904,N_908);
and U1009 (N_1009,N_873,N_978);
nor U1010 (N_1010,N_813,N_828);
nand U1011 (N_1011,N_922,N_926);
nand U1012 (N_1012,N_811,N_841);
nand U1013 (N_1013,N_931,N_876);
nor U1014 (N_1014,N_830,N_961);
nor U1015 (N_1015,N_935,N_900);
and U1016 (N_1016,N_942,N_893);
and U1017 (N_1017,N_937,N_808);
nor U1018 (N_1018,N_905,N_872);
or U1019 (N_1019,N_857,N_913);
nand U1020 (N_1020,N_879,N_918);
nor U1021 (N_1021,N_985,N_815);
or U1022 (N_1022,N_964,N_842);
nor U1023 (N_1023,N_962,N_899);
nand U1024 (N_1024,N_892,N_887);
nor U1025 (N_1025,N_932,N_854);
nor U1026 (N_1026,N_888,N_834);
or U1027 (N_1027,N_987,N_924);
and U1028 (N_1028,N_869,N_901);
nor U1029 (N_1029,N_967,N_807);
nor U1030 (N_1030,N_805,N_921);
nor U1031 (N_1031,N_944,N_812);
and U1032 (N_1032,N_886,N_955);
nor U1033 (N_1033,N_816,N_824);
nor U1034 (N_1034,N_866,N_909);
nor U1035 (N_1035,N_957,N_976);
or U1036 (N_1036,N_914,N_829);
or U1037 (N_1037,N_991,N_871);
nand U1038 (N_1038,N_835,N_839);
nor U1039 (N_1039,N_954,N_802);
nand U1040 (N_1040,N_983,N_875);
nand U1041 (N_1041,N_884,N_974);
nand U1042 (N_1042,N_855,N_838);
and U1043 (N_1043,N_868,N_948);
nand U1044 (N_1044,N_950,N_971);
nand U1045 (N_1045,N_966,N_864);
or U1046 (N_1046,N_993,N_826);
nor U1047 (N_1047,N_936,N_858);
nor U1048 (N_1048,N_970,N_989);
and U1049 (N_1049,N_862,N_856);
and U1050 (N_1050,N_982,N_851);
and U1051 (N_1051,N_889,N_867);
or U1052 (N_1052,N_827,N_911);
and U1053 (N_1053,N_981,N_920);
or U1054 (N_1054,N_939,N_846);
nand U1055 (N_1055,N_881,N_959);
or U1056 (N_1056,N_946,N_997);
and U1057 (N_1057,N_820,N_992);
or U1058 (N_1058,N_930,N_977);
or U1059 (N_1059,N_801,N_953);
and U1060 (N_1060,N_877,N_831);
and U1061 (N_1061,N_965,N_995);
nand U1062 (N_1062,N_833,N_912);
or U1063 (N_1063,N_863,N_844);
nor U1064 (N_1064,N_990,N_885);
and U1065 (N_1065,N_949,N_845);
and U1066 (N_1066,N_819,N_907);
nand U1067 (N_1067,N_804,N_906);
nor U1068 (N_1068,N_823,N_860);
nand U1069 (N_1069,N_986,N_994);
and U1070 (N_1070,N_973,N_832);
or U1071 (N_1071,N_928,N_903);
and U1072 (N_1072,N_963,N_883);
and U1073 (N_1073,N_975,N_874);
nor U1074 (N_1074,N_882,N_896);
nor U1075 (N_1075,N_809,N_891);
or U1076 (N_1076,N_941,N_843);
nand U1077 (N_1077,N_847,N_933);
and U1078 (N_1078,N_825,N_943);
or U1079 (N_1079,N_853,N_898);
or U1080 (N_1080,N_969,N_979);
nand U1081 (N_1081,N_852,N_980);
and U1082 (N_1082,N_915,N_894);
nor U1083 (N_1083,N_817,N_940);
and U1084 (N_1084,N_996,N_880);
nand U1085 (N_1085,N_958,N_814);
and U1086 (N_1086,N_836,N_923);
and U1087 (N_1087,N_837,N_972);
xnor U1088 (N_1088,N_929,N_927);
nor U1089 (N_1089,N_952,N_850);
and U1090 (N_1090,N_840,N_919);
nor U1091 (N_1091,N_849,N_895);
or U1092 (N_1092,N_925,N_861);
nor U1093 (N_1093,N_998,N_956);
or U1094 (N_1094,N_870,N_917);
and U1095 (N_1095,N_902,N_938);
or U1096 (N_1096,N_988,N_968);
nor U1097 (N_1097,N_803,N_951);
or U1098 (N_1098,N_806,N_818);
and U1099 (N_1099,N_945,N_821);
nor U1100 (N_1100,N_875,N_918);
nand U1101 (N_1101,N_926,N_898);
or U1102 (N_1102,N_951,N_954);
and U1103 (N_1103,N_938,N_894);
or U1104 (N_1104,N_927,N_854);
nor U1105 (N_1105,N_868,N_832);
or U1106 (N_1106,N_802,N_910);
nand U1107 (N_1107,N_847,N_832);
nand U1108 (N_1108,N_925,N_963);
or U1109 (N_1109,N_923,N_961);
and U1110 (N_1110,N_847,N_884);
and U1111 (N_1111,N_814,N_947);
and U1112 (N_1112,N_883,N_955);
or U1113 (N_1113,N_860,N_999);
nor U1114 (N_1114,N_860,N_851);
nor U1115 (N_1115,N_963,N_940);
and U1116 (N_1116,N_917,N_890);
nand U1117 (N_1117,N_933,N_805);
and U1118 (N_1118,N_866,N_877);
or U1119 (N_1119,N_913,N_803);
or U1120 (N_1120,N_910,N_886);
and U1121 (N_1121,N_928,N_965);
and U1122 (N_1122,N_908,N_975);
and U1123 (N_1123,N_947,N_876);
or U1124 (N_1124,N_844,N_805);
and U1125 (N_1125,N_861,N_967);
nor U1126 (N_1126,N_970,N_996);
nand U1127 (N_1127,N_860,N_829);
nand U1128 (N_1128,N_952,N_969);
nor U1129 (N_1129,N_823,N_834);
nor U1130 (N_1130,N_854,N_851);
or U1131 (N_1131,N_835,N_972);
nand U1132 (N_1132,N_998,N_881);
and U1133 (N_1133,N_962,N_985);
or U1134 (N_1134,N_903,N_832);
nor U1135 (N_1135,N_889,N_996);
and U1136 (N_1136,N_842,N_893);
xor U1137 (N_1137,N_926,N_819);
nor U1138 (N_1138,N_862,N_850);
and U1139 (N_1139,N_858,N_818);
nor U1140 (N_1140,N_880,N_877);
nand U1141 (N_1141,N_912,N_852);
nand U1142 (N_1142,N_844,N_936);
nand U1143 (N_1143,N_835,N_997);
or U1144 (N_1144,N_893,N_977);
xor U1145 (N_1145,N_909,N_991);
and U1146 (N_1146,N_945,N_840);
nand U1147 (N_1147,N_889,N_869);
nor U1148 (N_1148,N_908,N_923);
and U1149 (N_1149,N_927,N_874);
and U1150 (N_1150,N_906,N_832);
and U1151 (N_1151,N_843,N_965);
and U1152 (N_1152,N_978,N_970);
nand U1153 (N_1153,N_837,N_802);
or U1154 (N_1154,N_958,N_951);
nor U1155 (N_1155,N_808,N_947);
nand U1156 (N_1156,N_830,N_891);
nor U1157 (N_1157,N_859,N_986);
or U1158 (N_1158,N_812,N_999);
nor U1159 (N_1159,N_801,N_882);
and U1160 (N_1160,N_881,N_874);
nor U1161 (N_1161,N_840,N_972);
and U1162 (N_1162,N_949,N_964);
nor U1163 (N_1163,N_917,N_878);
or U1164 (N_1164,N_876,N_951);
or U1165 (N_1165,N_867,N_861);
nand U1166 (N_1166,N_952,N_867);
or U1167 (N_1167,N_938,N_960);
nand U1168 (N_1168,N_889,N_975);
and U1169 (N_1169,N_959,N_823);
nor U1170 (N_1170,N_806,N_830);
and U1171 (N_1171,N_914,N_843);
or U1172 (N_1172,N_945,N_827);
nand U1173 (N_1173,N_983,N_923);
or U1174 (N_1174,N_824,N_985);
nor U1175 (N_1175,N_960,N_909);
or U1176 (N_1176,N_891,N_938);
or U1177 (N_1177,N_937,N_980);
nor U1178 (N_1178,N_992,N_824);
nand U1179 (N_1179,N_911,N_834);
nand U1180 (N_1180,N_997,N_908);
or U1181 (N_1181,N_901,N_848);
nand U1182 (N_1182,N_897,N_911);
or U1183 (N_1183,N_923,N_806);
or U1184 (N_1184,N_901,N_986);
or U1185 (N_1185,N_934,N_857);
nor U1186 (N_1186,N_804,N_875);
and U1187 (N_1187,N_986,N_964);
nor U1188 (N_1188,N_969,N_913);
nor U1189 (N_1189,N_819,N_942);
nand U1190 (N_1190,N_945,N_844);
or U1191 (N_1191,N_983,N_820);
nand U1192 (N_1192,N_944,N_913);
and U1193 (N_1193,N_908,N_839);
nand U1194 (N_1194,N_883,N_839);
and U1195 (N_1195,N_815,N_958);
and U1196 (N_1196,N_864,N_950);
nand U1197 (N_1197,N_945,N_814);
nand U1198 (N_1198,N_853,N_899);
nand U1199 (N_1199,N_922,N_873);
nor U1200 (N_1200,N_1184,N_1059);
nor U1201 (N_1201,N_1037,N_1023);
nand U1202 (N_1202,N_1033,N_1139);
and U1203 (N_1203,N_1015,N_1197);
and U1204 (N_1204,N_1077,N_1128);
or U1205 (N_1205,N_1048,N_1032);
nor U1206 (N_1206,N_1009,N_1165);
and U1207 (N_1207,N_1018,N_1195);
nand U1208 (N_1208,N_1011,N_1140);
nor U1209 (N_1209,N_1111,N_1024);
nor U1210 (N_1210,N_1188,N_1153);
and U1211 (N_1211,N_1066,N_1148);
or U1212 (N_1212,N_1081,N_1105);
and U1213 (N_1213,N_1088,N_1110);
or U1214 (N_1214,N_1064,N_1054);
nand U1215 (N_1215,N_1145,N_1118);
nand U1216 (N_1216,N_1181,N_1055);
or U1217 (N_1217,N_1103,N_1121);
or U1218 (N_1218,N_1030,N_1102);
nor U1219 (N_1219,N_1127,N_1007);
nand U1220 (N_1220,N_1194,N_1065);
or U1221 (N_1221,N_1095,N_1146);
or U1222 (N_1222,N_1176,N_1096);
and U1223 (N_1223,N_1014,N_1017);
and U1224 (N_1224,N_1010,N_1090);
or U1225 (N_1225,N_1164,N_1160);
or U1226 (N_1226,N_1039,N_1013);
nor U1227 (N_1227,N_1152,N_1004);
nor U1228 (N_1228,N_1162,N_1143);
nand U1229 (N_1229,N_1047,N_1022);
nand U1230 (N_1230,N_1051,N_1183);
nor U1231 (N_1231,N_1092,N_1142);
or U1232 (N_1232,N_1167,N_1124);
nor U1233 (N_1233,N_1166,N_1057);
or U1234 (N_1234,N_1122,N_1191);
nand U1235 (N_1235,N_1170,N_1120);
nor U1236 (N_1236,N_1116,N_1106);
nand U1237 (N_1237,N_1001,N_1151);
nor U1238 (N_1238,N_1028,N_1182);
nor U1239 (N_1239,N_1008,N_1071);
nor U1240 (N_1240,N_1156,N_1006);
or U1241 (N_1241,N_1114,N_1137);
and U1242 (N_1242,N_1060,N_1169);
nor U1243 (N_1243,N_1187,N_1198);
nand U1244 (N_1244,N_1021,N_1079);
nand U1245 (N_1245,N_1125,N_1147);
or U1246 (N_1246,N_1173,N_1135);
nor U1247 (N_1247,N_1113,N_1005);
nor U1248 (N_1248,N_1083,N_1029);
nand U1249 (N_1249,N_1168,N_1100);
nand U1250 (N_1250,N_1178,N_1080);
or U1251 (N_1251,N_1063,N_1097);
and U1252 (N_1252,N_1089,N_1074);
nand U1253 (N_1253,N_1036,N_1072);
nand U1254 (N_1254,N_1175,N_1049);
or U1255 (N_1255,N_1034,N_1185);
nor U1256 (N_1256,N_1085,N_1109);
nor U1257 (N_1257,N_1069,N_1192);
nor U1258 (N_1258,N_1180,N_1115);
and U1259 (N_1259,N_1099,N_1019);
or U1260 (N_1260,N_1130,N_1094);
or U1261 (N_1261,N_1150,N_1087);
nand U1262 (N_1262,N_1131,N_1025);
nand U1263 (N_1263,N_1112,N_1199);
or U1264 (N_1264,N_1177,N_1123);
or U1265 (N_1265,N_1107,N_1108);
and U1266 (N_1266,N_1141,N_1155);
or U1267 (N_1267,N_1038,N_1134);
or U1268 (N_1268,N_1174,N_1126);
xnor U1269 (N_1269,N_1138,N_1093);
nand U1270 (N_1270,N_1073,N_1067);
nand U1271 (N_1271,N_1172,N_1091);
nor U1272 (N_1272,N_1104,N_1171);
nor U1273 (N_1273,N_1020,N_1129);
nand U1274 (N_1274,N_1084,N_1149);
nand U1275 (N_1275,N_1119,N_1027);
nand U1276 (N_1276,N_1040,N_1132);
and U1277 (N_1277,N_1053,N_1098);
or U1278 (N_1278,N_1035,N_1136);
nand U1279 (N_1279,N_1161,N_1026);
or U1280 (N_1280,N_1031,N_1163);
and U1281 (N_1281,N_1016,N_1159);
nor U1282 (N_1282,N_1000,N_1041);
and U1283 (N_1283,N_1179,N_1056);
and U1284 (N_1284,N_1045,N_1002);
and U1285 (N_1285,N_1082,N_1044);
nor U1286 (N_1286,N_1042,N_1078);
nand U1287 (N_1287,N_1193,N_1157);
or U1288 (N_1288,N_1075,N_1101);
nand U1289 (N_1289,N_1012,N_1196);
nand U1290 (N_1290,N_1190,N_1189);
nor U1291 (N_1291,N_1043,N_1058);
nand U1292 (N_1292,N_1117,N_1061);
or U1293 (N_1293,N_1154,N_1133);
or U1294 (N_1294,N_1068,N_1062);
nor U1295 (N_1295,N_1076,N_1186);
nand U1296 (N_1296,N_1144,N_1086);
or U1297 (N_1297,N_1003,N_1046);
nor U1298 (N_1298,N_1070,N_1158);
nor U1299 (N_1299,N_1052,N_1050);
nor U1300 (N_1300,N_1127,N_1065);
or U1301 (N_1301,N_1192,N_1042);
and U1302 (N_1302,N_1160,N_1051);
nor U1303 (N_1303,N_1133,N_1169);
or U1304 (N_1304,N_1048,N_1007);
and U1305 (N_1305,N_1092,N_1139);
or U1306 (N_1306,N_1172,N_1180);
and U1307 (N_1307,N_1059,N_1108);
or U1308 (N_1308,N_1137,N_1193);
nand U1309 (N_1309,N_1182,N_1017);
nor U1310 (N_1310,N_1083,N_1040);
nor U1311 (N_1311,N_1199,N_1193);
nor U1312 (N_1312,N_1041,N_1104);
or U1313 (N_1313,N_1127,N_1181);
or U1314 (N_1314,N_1152,N_1153);
nor U1315 (N_1315,N_1026,N_1036);
nor U1316 (N_1316,N_1012,N_1113);
and U1317 (N_1317,N_1146,N_1185);
nand U1318 (N_1318,N_1091,N_1076);
and U1319 (N_1319,N_1010,N_1034);
nor U1320 (N_1320,N_1015,N_1127);
nor U1321 (N_1321,N_1045,N_1194);
nand U1322 (N_1322,N_1104,N_1186);
or U1323 (N_1323,N_1187,N_1133);
and U1324 (N_1324,N_1099,N_1189);
or U1325 (N_1325,N_1087,N_1040);
or U1326 (N_1326,N_1189,N_1170);
or U1327 (N_1327,N_1154,N_1069);
nor U1328 (N_1328,N_1183,N_1129);
and U1329 (N_1329,N_1013,N_1071);
or U1330 (N_1330,N_1157,N_1007);
or U1331 (N_1331,N_1019,N_1082);
nand U1332 (N_1332,N_1134,N_1100);
nor U1333 (N_1333,N_1105,N_1054);
nor U1334 (N_1334,N_1055,N_1048);
and U1335 (N_1335,N_1184,N_1094);
nor U1336 (N_1336,N_1061,N_1006);
or U1337 (N_1337,N_1074,N_1167);
and U1338 (N_1338,N_1191,N_1193);
nand U1339 (N_1339,N_1165,N_1124);
nor U1340 (N_1340,N_1072,N_1033);
and U1341 (N_1341,N_1127,N_1002);
and U1342 (N_1342,N_1000,N_1019);
nand U1343 (N_1343,N_1003,N_1146);
nand U1344 (N_1344,N_1127,N_1064);
nor U1345 (N_1345,N_1056,N_1126);
nor U1346 (N_1346,N_1057,N_1054);
nor U1347 (N_1347,N_1118,N_1192);
nor U1348 (N_1348,N_1190,N_1042);
and U1349 (N_1349,N_1193,N_1021);
nand U1350 (N_1350,N_1065,N_1012);
or U1351 (N_1351,N_1040,N_1029);
nor U1352 (N_1352,N_1165,N_1123);
nand U1353 (N_1353,N_1025,N_1031);
nor U1354 (N_1354,N_1150,N_1091);
and U1355 (N_1355,N_1110,N_1155);
nand U1356 (N_1356,N_1050,N_1018);
and U1357 (N_1357,N_1177,N_1179);
and U1358 (N_1358,N_1014,N_1078);
and U1359 (N_1359,N_1030,N_1139);
and U1360 (N_1360,N_1148,N_1094);
and U1361 (N_1361,N_1184,N_1003);
and U1362 (N_1362,N_1014,N_1065);
nand U1363 (N_1363,N_1196,N_1036);
or U1364 (N_1364,N_1140,N_1047);
nand U1365 (N_1365,N_1194,N_1090);
or U1366 (N_1366,N_1163,N_1004);
nand U1367 (N_1367,N_1079,N_1070);
or U1368 (N_1368,N_1141,N_1184);
nand U1369 (N_1369,N_1076,N_1183);
nand U1370 (N_1370,N_1012,N_1018);
or U1371 (N_1371,N_1199,N_1032);
and U1372 (N_1372,N_1132,N_1188);
nor U1373 (N_1373,N_1052,N_1066);
nor U1374 (N_1374,N_1025,N_1040);
nand U1375 (N_1375,N_1149,N_1143);
and U1376 (N_1376,N_1053,N_1007);
nand U1377 (N_1377,N_1087,N_1045);
and U1378 (N_1378,N_1007,N_1026);
nor U1379 (N_1379,N_1088,N_1196);
or U1380 (N_1380,N_1194,N_1019);
or U1381 (N_1381,N_1122,N_1079);
and U1382 (N_1382,N_1032,N_1098);
xnor U1383 (N_1383,N_1057,N_1105);
or U1384 (N_1384,N_1154,N_1013);
or U1385 (N_1385,N_1180,N_1175);
or U1386 (N_1386,N_1092,N_1049);
nand U1387 (N_1387,N_1022,N_1125);
nand U1388 (N_1388,N_1000,N_1187);
or U1389 (N_1389,N_1146,N_1063);
nand U1390 (N_1390,N_1017,N_1102);
xor U1391 (N_1391,N_1147,N_1175);
or U1392 (N_1392,N_1081,N_1156);
nor U1393 (N_1393,N_1143,N_1181);
nor U1394 (N_1394,N_1110,N_1030);
nand U1395 (N_1395,N_1112,N_1145);
and U1396 (N_1396,N_1146,N_1096);
and U1397 (N_1397,N_1198,N_1161);
or U1398 (N_1398,N_1147,N_1165);
nor U1399 (N_1399,N_1010,N_1155);
nor U1400 (N_1400,N_1217,N_1330);
nand U1401 (N_1401,N_1352,N_1338);
or U1402 (N_1402,N_1298,N_1392);
nand U1403 (N_1403,N_1220,N_1251);
nand U1404 (N_1404,N_1268,N_1216);
nor U1405 (N_1405,N_1332,N_1283);
and U1406 (N_1406,N_1316,N_1257);
nor U1407 (N_1407,N_1269,N_1231);
or U1408 (N_1408,N_1219,N_1333);
and U1409 (N_1409,N_1303,N_1385);
or U1410 (N_1410,N_1275,N_1288);
or U1411 (N_1411,N_1238,N_1373);
or U1412 (N_1412,N_1278,N_1313);
nand U1413 (N_1413,N_1314,N_1381);
or U1414 (N_1414,N_1261,N_1299);
nor U1415 (N_1415,N_1293,N_1372);
or U1416 (N_1416,N_1256,N_1201);
nor U1417 (N_1417,N_1344,N_1259);
and U1418 (N_1418,N_1252,N_1311);
nor U1419 (N_1419,N_1263,N_1368);
nor U1420 (N_1420,N_1272,N_1226);
or U1421 (N_1421,N_1273,N_1355);
or U1422 (N_1422,N_1215,N_1205);
nand U1423 (N_1423,N_1235,N_1397);
nor U1424 (N_1424,N_1221,N_1237);
and U1425 (N_1425,N_1229,N_1258);
or U1426 (N_1426,N_1391,N_1315);
nand U1427 (N_1427,N_1339,N_1354);
nor U1428 (N_1428,N_1208,N_1209);
or U1429 (N_1429,N_1342,N_1271);
and U1430 (N_1430,N_1395,N_1239);
nand U1431 (N_1431,N_1324,N_1270);
and U1432 (N_1432,N_1227,N_1294);
nand U1433 (N_1433,N_1246,N_1331);
nor U1434 (N_1434,N_1399,N_1377);
nand U1435 (N_1435,N_1267,N_1379);
nand U1436 (N_1436,N_1264,N_1281);
nand U1437 (N_1437,N_1382,N_1383);
and U1438 (N_1438,N_1370,N_1244);
nand U1439 (N_1439,N_1389,N_1224);
nor U1440 (N_1440,N_1203,N_1353);
or U1441 (N_1441,N_1343,N_1253);
nand U1442 (N_1442,N_1341,N_1326);
nand U1443 (N_1443,N_1320,N_1290);
and U1444 (N_1444,N_1384,N_1211);
nand U1445 (N_1445,N_1374,N_1212);
or U1446 (N_1446,N_1286,N_1297);
and U1447 (N_1447,N_1300,N_1348);
nor U1448 (N_1448,N_1365,N_1317);
and U1449 (N_1449,N_1260,N_1213);
nor U1450 (N_1450,N_1302,N_1388);
nor U1451 (N_1451,N_1349,N_1265);
and U1452 (N_1452,N_1361,N_1301);
nand U1453 (N_1453,N_1277,N_1318);
nor U1454 (N_1454,N_1360,N_1367);
or U1455 (N_1455,N_1262,N_1323);
nor U1456 (N_1456,N_1319,N_1312);
nor U1457 (N_1457,N_1223,N_1328);
nand U1458 (N_1458,N_1366,N_1375);
nor U1459 (N_1459,N_1228,N_1254);
or U1460 (N_1460,N_1266,N_1234);
or U1461 (N_1461,N_1327,N_1296);
nand U1462 (N_1462,N_1322,N_1335);
and U1463 (N_1463,N_1369,N_1340);
and U1464 (N_1464,N_1210,N_1247);
nor U1465 (N_1465,N_1248,N_1345);
nor U1466 (N_1466,N_1274,N_1292);
and U1467 (N_1467,N_1255,N_1337);
nand U1468 (N_1468,N_1222,N_1356);
or U1469 (N_1469,N_1276,N_1280);
nand U1470 (N_1470,N_1207,N_1243);
nand U1471 (N_1471,N_1350,N_1346);
nor U1472 (N_1472,N_1329,N_1206);
or U1473 (N_1473,N_1362,N_1305);
or U1474 (N_1474,N_1394,N_1359);
or U1475 (N_1475,N_1351,N_1202);
nand U1476 (N_1476,N_1334,N_1347);
and U1477 (N_1477,N_1236,N_1245);
nand U1478 (N_1478,N_1398,N_1364);
nand U1479 (N_1479,N_1289,N_1304);
nand U1480 (N_1480,N_1282,N_1358);
or U1481 (N_1481,N_1307,N_1308);
or U1482 (N_1482,N_1230,N_1250);
or U1483 (N_1483,N_1249,N_1309);
nor U1484 (N_1484,N_1285,N_1390);
nand U1485 (N_1485,N_1214,N_1396);
nor U1486 (N_1486,N_1279,N_1386);
nor U1487 (N_1487,N_1232,N_1240);
or U1488 (N_1488,N_1291,N_1357);
or U1489 (N_1489,N_1325,N_1295);
and U1490 (N_1490,N_1310,N_1387);
nor U1491 (N_1491,N_1241,N_1204);
and U1492 (N_1492,N_1371,N_1233);
or U1493 (N_1493,N_1393,N_1363);
nand U1494 (N_1494,N_1284,N_1336);
or U1495 (N_1495,N_1225,N_1321);
nor U1496 (N_1496,N_1242,N_1376);
and U1497 (N_1497,N_1218,N_1378);
or U1498 (N_1498,N_1200,N_1380);
and U1499 (N_1499,N_1287,N_1306);
nand U1500 (N_1500,N_1389,N_1312);
or U1501 (N_1501,N_1317,N_1201);
and U1502 (N_1502,N_1378,N_1335);
nor U1503 (N_1503,N_1279,N_1307);
or U1504 (N_1504,N_1265,N_1213);
and U1505 (N_1505,N_1320,N_1249);
nand U1506 (N_1506,N_1244,N_1289);
nor U1507 (N_1507,N_1209,N_1201);
or U1508 (N_1508,N_1268,N_1235);
and U1509 (N_1509,N_1243,N_1288);
nor U1510 (N_1510,N_1360,N_1330);
and U1511 (N_1511,N_1313,N_1316);
nand U1512 (N_1512,N_1258,N_1349);
and U1513 (N_1513,N_1350,N_1273);
nand U1514 (N_1514,N_1344,N_1230);
nand U1515 (N_1515,N_1218,N_1382);
or U1516 (N_1516,N_1349,N_1322);
nand U1517 (N_1517,N_1397,N_1360);
nor U1518 (N_1518,N_1371,N_1315);
nand U1519 (N_1519,N_1367,N_1245);
and U1520 (N_1520,N_1340,N_1373);
and U1521 (N_1521,N_1281,N_1215);
and U1522 (N_1522,N_1202,N_1312);
or U1523 (N_1523,N_1307,N_1288);
nor U1524 (N_1524,N_1371,N_1311);
nor U1525 (N_1525,N_1315,N_1248);
xnor U1526 (N_1526,N_1354,N_1231);
and U1527 (N_1527,N_1209,N_1232);
and U1528 (N_1528,N_1251,N_1376);
nor U1529 (N_1529,N_1276,N_1286);
nor U1530 (N_1530,N_1285,N_1394);
or U1531 (N_1531,N_1262,N_1282);
nor U1532 (N_1532,N_1247,N_1389);
and U1533 (N_1533,N_1244,N_1333);
nor U1534 (N_1534,N_1373,N_1221);
nor U1535 (N_1535,N_1274,N_1268);
and U1536 (N_1536,N_1218,N_1252);
nor U1537 (N_1537,N_1372,N_1287);
nor U1538 (N_1538,N_1203,N_1289);
nor U1539 (N_1539,N_1221,N_1389);
or U1540 (N_1540,N_1256,N_1218);
nor U1541 (N_1541,N_1252,N_1365);
nor U1542 (N_1542,N_1274,N_1230);
or U1543 (N_1543,N_1250,N_1286);
and U1544 (N_1544,N_1205,N_1273);
nor U1545 (N_1545,N_1367,N_1351);
and U1546 (N_1546,N_1327,N_1300);
nor U1547 (N_1547,N_1326,N_1203);
nand U1548 (N_1548,N_1338,N_1364);
or U1549 (N_1549,N_1307,N_1349);
or U1550 (N_1550,N_1367,N_1304);
xor U1551 (N_1551,N_1354,N_1352);
and U1552 (N_1552,N_1397,N_1248);
or U1553 (N_1553,N_1376,N_1340);
nand U1554 (N_1554,N_1290,N_1241);
nand U1555 (N_1555,N_1359,N_1385);
and U1556 (N_1556,N_1392,N_1320);
or U1557 (N_1557,N_1389,N_1200);
nor U1558 (N_1558,N_1206,N_1245);
nand U1559 (N_1559,N_1361,N_1344);
or U1560 (N_1560,N_1295,N_1221);
nor U1561 (N_1561,N_1364,N_1254);
or U1562 (N_1562,N_1239,N_1211);
nand U1563 (N_1563,N_1300,N_1331);
nand U1564 (N_1564,N_1276,N_1392);
nor U1565 (N_1565,N_1340,N_1364);
nor U1566 (N_1566,N_1382,N_1248);
nor U1567 (N_1567,N_1359,N_1255);
and U1568 (N_1568,N_1362,N_1286);
or U1569 (N_1569,N_1203,N_1313);
nand U1570 (N_1570,N_1214,N_1318);
and U1571 (N_1571,N_1376,N_1378);
nand U1572 (N_1572,N_1251,N_1238);
and U1573 (N_1573,N_1245,N_1375);
nand U1574 (N_1574,N_1304,N_1390);
nand U1575 (N_1575,N_1226,N_1246);
and U1576 (N_1576,N_1395,N_1278);
and U1577 (N_1577,N_1382,N_1360);
and U1578 (N_1578,N_1284,N_1331);
and U1579 (N_1579,N_1379,N_1296);
nor U1580 (N_1580,N_1288,N_1305);
nor U1581 (N_1581,N_1230,N_1266);
or U1582 (N_1582,N_1378,N_1213);
nand U1583 (N_1583,N_1204,N_1360);
nand U1584 (N_1584,N_1277,N_1355);
or U1585 (N_1585,N_1227,N_1251);
nor U1586 (N_1586,N_1280,N_1258);
or U1587 (N_1587,N_1316,N_1288);
and U1588 (N_1588,N_1366,N_1239);
and U1589 (N_1589,N_1392,N_1261);
or U1590 (N_1590,N_1262,N_1376);
nand U1591 (N_1591,N_1294,N_1270);
and U1592 (N_1592,N_1240,N_1316);
and U1593 (N_1593,N_1283,N_1240);
or U1594 (N_1594,N_1349,N_1213);
nand U1595 (N_1595,N_1220,N_1211);
nand U1596 (N_1596,N_1255,N_1202);
and U1597 (N_1597,N_1336,N_1382);
and U1598 (N_1598,N_1338,N_1230);
and U1599 (N_1599,N_1328,N_1333);
and U1600 (N_1600,N_1466,N_1496);
nand U1601 (N_1601,N_1432,N_1417);
or U1602 (N_1602,N_1589,N_1596);
nor U1603 (N_1603,N_1464,N_1439);
nor U1604 (N_1604,N_1414,N_1551);
nor U1605 (N_1605,N_1401,N_1467);
nand U1606 (N_1606,N_1489,N_1509);
or U1607 (N_1607,N_1549,N_1402);
nand U1608 (N_1608,N_1488,N_1456);
nand U1609 (N_1609,N_1514,N_1420);
nand U1610 (N_1610,N_1582,N_1538);
nand U1611 (N_1611,N_1480,N_1500);
nand U1612 (N_1612,N_1460,N_1434);
and U1613 (N_1613,N_1413,N_1447);
nor U1614 (N_1614,N_1555,N_1592);
or U1615 (N_1615,N_1587,N_1491);
and U1616 (N_1616,N_1476,N_1527);
or U1617 (N_1617,N_1498,N_1481);
and U1618 (N_1618,N_1553,N_1449);
or U1619 (N_1619,N_1594,N_1451);
and U1620 (N_1620,N_1559,N_1580);
and U1621 (N_1621,N_1463,N_1472);
nand U1622 (N_1622,N_1428,N_1517);
nand U1623 (N_1623,N_1520,N_1506);
and U1624 (N_1624,N_1407,N_1550);
or U1625 (N_1625,N_1547,N_1571);
nor U1626 (N_1626,N_1415,N_1597);
nand U1627 (N_1627,N_1530,N_1442);
and U1628 (N_1628,N_1518,N_1411);
and U1629 (N_1629,N_1431,N_1532);
nor U1630 (N_1630,N_1543,N_1444);
nor U1631 (N_1631,N_1537,N_1536);
and U1632 (N_1632,N_1535,N_1574);
nand U1633 (N_1633,N_1531,N_1521);
or U1634 (N_1634,N_1523,N_1577);
nand U1635 (N_1635,N_1408,N_1598);
nor U1636 (N_1636,N_1557,N_1525);
or U1637 (N_1637,N_1583,N_1516);
nor U1638 (N_1638,N_1418,N_1524);
or U1639 (N_1639,N_1503,N_1507);
nor U1640 (N_1640,N_1505,N_1400);
nand U1641 (N_1641,N_1484,N_1446);
and U1642 (N_1642,N_1425,N_1542);
or U1643 (N_1643,N_1435,N_1522);
nand U1644 (N_1644,N_1437,N_1526);
or U1645 (N_1645,N_1424,N_1479);
nand U1646 (N_1646,N_1490,N_1492);
nand U1647 (N_1647,N_1461,N_1548);
or U1648 (N_1648,N_1416,N_1445);
or U1649 (N_1649,N_1430,N_1495);
nand U1650 (N_1650,N_1477,N_1405);
and U1651 (N_1651,N_1469,N_1519);
xnor U1652 (N_1652,N_1534,N_1504);
and U1653 (N_1653,N_1513,N_1515);
or U1654 (N_1654,N_1443,N_1568);
nor U1655 (N_1655,N_1468,N_1508);
and U1656 (N_1656,N_1438,N_1561);
and U1657 (N_1657,N_1455,N_1575);
and U1658 (N_1658,N_1485,N_1433);
nor U1659 (N_1659,N_1459,N_1539);
nor U1660 (N_1660,N_1448,N_1569);
nand U1661 (N_1661,N_1578,N_1478);
or U1662 (N_1662,N_1493,N_1454);
or U1663 (N_1663,N_1593,N_1556);
or U1664 (N_1664,N_1404,N_1426);
or U1665 (N_1665,N_1423,N_1588);
and U1666 (N_1666,N_1483,N_1465);
nand U1667 (N_1667,N_1560,N_1554);
and U1668 (N_1668,N_1501,N_1473);
nand U1669 (N_1669,N_1497,N_1591);
and U1670 (N_1670,N_1595,N_1471);
nand U1671 (N_1671,N_1462,N_1458);
or U1672 (N_1672,N_1567,N_1566);
xor U1673 (N_1673,N_1494,N_1576);
nor U1674 (N_1674,N_1406,N_1427);
nor U1675 (N_1675,N_1586,N_1544);
nand U1676 (N_1676,N_1572,N_1590);
xor U1677 (N_1677,N_1545,N_1441);
nand U1678 (N_1678,N_1540,N_1470);
nor U1679 (N_1679,N_1412,N_1584);
nand U1680 (N_1680,N_1563,N_1453);
and U1681 (N_1681,N_1541,N_1564);
and U1682 (N_1682,N_1429,N_1450);
nand U1683 (N_1683,N_1502,N_1452);
nor U1684 (N_1684,N_1440,N_1486);
nand U1685 (N_1685,N_1529,N_1457);
nor U1686 (N_1686,N_1565,N_1570);
and U1687 (N_1687,N_1510,N_1581);
or U1688 (N_1688,N_1528,N_1421);
nand U1689 (N_1689,N_1403,N_1558);
and U1690 (N_1690,N_1410,N_1487);
and U1691 (N_1691,N_1533,N_1499);
nand U1692 (N_1692,N_1436,N_1474);
and U1693 (N_1693,N_1573,N_1419);
xor U1694 (N_1694,N_1512,N_1482);
or U1695 (N_1695,N_1422,N_1579);
or U1696 (N_1696,N_1409,N_1599);
or U1697 (N_1697,N_1511,N_1546);
or U1698 (N_1698,N_1562,N_1585);
or U1699 (N_1699,N_1552,N_1475);
or U1700 (N_1700,N_1431,N_1468);
and U1701 (N_1701,N_1517,N_1491);
nand U1702 (N_1702,N_1421,N_1555);
nand U1703 (N_1703,N_1471,N_1546);
or U1704 (N_1704,N_1419,N_1452);
nand U1705 (N_1705,N_1469,N_1548);
nor U1706 (N_1706,N_1592,N_1508);
or U1707 (N_1707,N_1546,N_1541);
or U1708 (N_1708,N_1437,N_1447);
nor U1709 (N_1709,N_1484,N_1455);
or U1710 (N_1710,N_1599,N_1568);
nor U1711 (N_1711,N_1476,N_1534);
nor U1712 (N_1712,N_1484,N_1568);
nor U1713 (N_1713,N_1539,N_1545);
nor U1714 (N_1714,N_1541,N_1455);
xnor U1715 (N_1715,N_1477,N_1587);
or U1716 (N_1716,N_1589,N_1555);
and U1717 (N_1717,N_1520,N_1570);
and U1718 (N_1718,N_1456,N_1474);
nand U1719 (N_1719,N_1581,N_1402);
nand U1720 (N_1720,N_1541,N_1443);
and U1721 (N_1721,N_1595,N_1565);
and U1722 (N_1722,N_1556,N_1525);
or U1723 (N_1723,N_1487,N_1513);
nor U1724 (N_1724,N_1548,N_1555);
nor U1725 (N_1725,N_1503,N_1496);
and U1726 (N_1726,N_1592,N_1437);
or U1727 (N_1727,N_1578,N_1550);
or U1728 (N_1728,N_1548,N_1493);
and U1729 (N_1729,N_1512,N_1472);
or U1730 (N_1730,N_1494,N_1546);
nor U1731 (N_1731,N_1489,N_1567);
nor U1732 (N_1732,N_1559,N_1432);
nand U1733 (N_1733,N_1586,N_1443);
and U1734 (N_1734,N_1431,N_1542);
or U1735 (N_1735,N_1416,N_1596);
nand U1736 (N_1736,N_1474,N_1556);
or U1737 (N_1737,N_1579,N_1547);
nand U1738 (N_1738,N_1565,N_1550);
nand U1739 (N_1739,N_1500,N_1559);
nand U1740 (N_1740,N_1463,N_1493);
or U1741 (N_1741,N_1591,N_1552);
nand U1742 (N_1742,N_1416,N_1447);
nor U1743 (N_1743,N_1432,N_1520);
and U1744 (N_1744,N_1479,N_1543);
nor U1745 (N_1745,N_1550,N_1485);
nand U1746 (N_1746,N_1405,N_1414);
or U1747 (N_1747,N_1403,N_1441);
and U1748 (N_1748,N_1557,N_1470);
and U1749 (N_1749,N_1557,N_1553);
nand U1750 (N_1750,N_1528,N_1535);
nand U1751 (N_1751,N_1438,N_1416);
or U1752 (N_1752,N_1547,N_1463);
and U1753 (N_1753,N_1417,N_1463);
and U1754 (N_1754,N_1481,N_1444);
and U1755 (N_1755,N_1577,N_1548);
and U1756 (N_1756,N_1482,N_1503);
or U1757 (N_1757,N_1568,N_1516);
and U1758 (N_1758,N_1435,N_1557);
and U1759 (N_1759,N_1574,N_1524);
and U1760 (N_1760,N_1590,N_1570);
and U1761 (N_1761,N_1408,N_1464);
nor U1762 (N_1762,N_1453,N_1561);
nor U1763 (N_1763,N_1411,N_1431);
nand U1764 (N_1764,N_1502,N_1529);
and U1765 (N_1765,N_1515,N_1547);
nor U1766 (N_1766,N_1429,N_1474);
nand U1767 (N_1767,N_1590,N_1520);
nand U1768 (N_1768,N_1476,N_1496);
nand U1769 (N_1769,N_1463,N_1416);
nor U1770 (N_1770,N_1562,N_1405);
or U1771 (N_1771,N_1549,N_1539);
and U1772 (N_1772,N_1503,N_1444);
and U1773 (N_1773,N_1497,N_1558);
nand U1774 (N_1774,N_1529,N_1411);
or U1775 (N_1775,N_1527,N_1410);
nor U1776 (N_1776,N_1439,N_1514);
nand U1777 (N_1777,N_1512,N_1458);
or U1778 (N_1778,N_1450,N_1458);
nor U1779 (N_1779,N_1562,N_1409);
or U1780 (N_1780,N_1528,N_1507);
nor U1781 (N_1781,N_1529,N_1453);
nor U1782 (N_1782,N_1518,N_1455);
or U1783 (N_1783,N_1456,N_1526);
xnor U1784 (N_1784,N_1578,N_1539);
or U1785 (N_1785,N_1450,N_1545);
xnor U1786 (N_1786,N_1509,N_1470);
nor U1787 (N_1787,N_1465,N_1471);
and U1788 (N_1788,N_1449,N_1436);
or U1789 (N_1789,N_1401,N_1549);
and U1790 (N_1790,N_1440,N_1458);
nor U1791 (N_1791,N_1592,N_1438);
nand U1792 (N_1792,N_1422,N_1509);
nor U1793 (N_1793,N_1532,N_1509);
nor U1794 (N_1794,N_1595,N_1558);
nor U1795 (N_1795,N_1536,N_1511);
and U1796 (N_1796,N_1565,N_1592);
nand U1797 (N_1797,N_1515,N_1449);
and U1798 (N_1798,N_1548,N_1560);
and U1799 (N_1799,N_1559,N_1441);
and U1800 (N_1800,N_1608,N_1605);
and U1801 (N_1801,N_1745,N_1723);
and U1802 (N_1802,N_1786,N_1630);
nand U1803 (N_1803,N_1639,N_1730);
or U1804 (N_1804,N_1758,N_1751);
nand U1805 (N_1805,N_1783,N_1683);
or U1806 (N_1806,N_1789,N_1689);
and U1807 (N_1807,N_1696,N_1648);
nand U1808 (N_1808,N_1795,N_1729);
nor U1809 (N_1809,N_1688,N_1618);
nor U1810 (N_1810,N_1661,N_1773);
nand U1811 (N_1811,N_1788,N_1752);
nor U1812 (N_1812,N_1685,N_1679);
or U1813 (N_1813,N_1771,N_1719);
nand U1814 (N_1814,N_1657,N_1669);
and U1815 (N_1815,N_1663,N_1700);
and U1816 (N_1816,N_1623,N_1655);
nor U1817 (N_1817,N_1770,N_1701);
and U1818 (N_1818,N_1732,N_1603);
nand U1819 (N_1819,N_1746,N_1767);
and U1820 (N_1820,N_1613,N_1627);
and U1821 (N_1821,N_1607,N_1601);
nand U1822 (N_1822,N_1763,N_1687);
nand U1823 (N_1823,N_1791,N_1785);
nor U1824 (N_1824,N_1602,N_1684);
nand U1825 (N_1825,N_1711,N_1634);
nor U1826 (N_1826,N_1664,N_1738);
or U1827 (N_1827,N_1726,N_1673);
nand U1828 (N_1828,N_1671,N_1675);
nor U1829 (N_1829,N_1635,N_1604);
nand U1830 (N_1830,N_1762,N_1660);
nand U1831 (N_1831,N_1695,N_1713);
nor U1832 (N_1832,N_1764,N_1631);
nand U1833 (N_1833,N_1744,N_1677);
xor U1834 (N_1834,N_1780,N_1728);
or U1835 (N_1835,N_1702,N_1636);
nor U1836 (N_1836,N_1778,N_1667);
nand U1837 (N_1837,N_1756,N_1697);
nand U1838 (N_1838,N_1735,N_1686);
or U1839 (N_1839,N_1644,N_1624);
nand U1840 (N_1840,N_1694,N_1658);
and U1841 (N_1841,N_1692,N_1761);
and U1842 (N_1842,N_1610,N_1676);
nand U1843 (N_1843,N_1725,N_1681);
nor U1844 (N_1844,N_1739,N_1733);
or U1845 (N_1845,N_1731,N_1779);
and U1846 (N_1846,N_1775,N_1665);
nand U1847 (N_1847,N_1653,N_1654);
or U1848 (N_1848,N_1629,N_1650);
nand U1849 (N_1849,N_1748,N_1724);
nand U1850 (N_1850,N_1600,N_1718);
nor U1851 (N_1851,N_1798,N_1737);
and U1852 (N_1852,N_1776,N_1643);
nand U1853 (N_1853,N_1668,N_1768);
nand U1854 (N_1854,N_1666,N_1609);
xnor U1855 (N_1855,N_1714,N_1766);
nand U1856 (N_1856,N_1637,N_1790);
nor U1857 (N_1857,N_1799,N_1670);
or U1858 (N_1858,N_1651,N_1727);
and U1859 (N_1859,N_1774,N_1740);
and U1860 (N_1860,N_1793,N_1721);
nand U1861 (N_1861,N_1656,N_1716);
or U1862 (N_1862,N_1645,N_1715);
nand U1863 (N_1863,N_1743,N_1617);
nor U1864 (N_1864,N_1753,N_1757);
or U1865 (N_1865,N_1772,N_1720);
nor U1866 (N_1866,N_1703,N_1792);
or U1867 (N_1867,N_1659,N_1641);
nor U1868 (N_1868,N_1698,N_1680);
nor U1869 (N_1869,N_1632,N_1704);
nand U1870 (N_1870,N_1707,N_1777);
nor U1871 (N_1871,N_1621,N_1736);
nand U1872 (N_1872,N_1796,N_1620);
or U1873 (N_1873,N_1682,N_1611);
or U1874 (N_1874,N_1642,N_1722);
nor U1875 (N_1875,N_1760,N_1672);
nand U1876 (N_1876,N_1706,N_1712);
or U1877 (N_1877,N_1612,N_1662);
or U1878 (N_1878,N_1765,N_1754);
nand U1879 (N_1879,N_1690,N_1615);
nand U1880 (N_1880,N_1749,N_1699);
nor U1881 (N_1881,N_1741,N_1633);
or U1882 (N_1882,N_1755,N_1750);
nand U1883 (N_1883,N_1646,N_1614);
and U1884 (N_1884,N_1769,N_1717);
nor U1885 (N_1885,N_1734,N_1759);
nor U1886 (N_1886,N_1626,N_1647);
and U1887 (N_1887,N_1622,N_1709);
nor U1888 (N_1888,N_1640,N_1782);
nand U1889 (N_1889,N_1797,N_1674);
and U1890 (N_1890,N_1652,N_1742);
nand U1891 (N_1891,N_1678,N_1710);
nor U1892 (N_1892,N_1787,N_1691);
or U1893 (N_1893,N_1649,N_1619);
and U1894 (N_1894,N_1638,N_1794);
or U1895 (N_1895,N_1625,N_1747);
nor U1896 (N_1896,N_1781,N_1784);
or U1897 (N_1897,N_1616,N_1606);
and U1898 (N_1898,N_1693,N_1708);
and U1899 (N_1899,N_1628,N_1705);
nor U1900 (N_1900,N_1794,N_1793);
and U1901 (N_1901,N_1618,N_1665);
nand U1902 (N_1902,N_1674,N_1662);
and U1903 (N_1903,N_1688,N_1707);
nor U1904 (N_1904,N_1742,N_1626);
or U1905 (N_1905,N_1706,N_1663);
nor U1906 (N_1906,N_1781,N_1795);
nand U1907 (N_1907,N_1777,N_1688);
nand U1908 (N_1908,N_1625,N_1716);
or U1909 (N_1909,N_1645,N_1781);
nor U1910 (N_1910,N_1620,N_1723);
and U1911 (N_1911,N_1752,N_1621);
and U1912 (N_1912,N_1708,N_1722);
nor U1913 (N_1913,N_1724,N_1796);
nand U1914 (N_1914,N_1765,N_1646);
nor U1915 (N_1915,N_1623,N_1617);
and U1916 (N_1916,N_1741,N_1668);
or U1917 (N_1917,N_1601,N_1773);
and U1918 (N_1918,N_1602,N_1676);
nand U1919 (N_1919,N_1611,N_1639);
nor U1920 (N_1920,N_1690,N_1631);
nor U1921 (N_1921,N_1695,N_1719);
and U1922 (N_1922,N_1769,N_1760);
or U1923 (N_1923,N_1622,N_1680);
and U1924 (N_1924,N_1713,N_1669);
or U1925 (N_1925,N_1729,N_1606);
or U1926 (N_1926,N_1718,N_1762);
nand U1927 (N_1927,N_1724,N_1688);
nand U1928 (N_1928,N_1782,N_1698);
nand U1929 (N_1929,N_1675,N_1604);
nor U1930 (N_1930,N_1631,N_1798);
nor U1931 (N_1931,N_1657,N_1662);
nand U1932 (N_1932,N_1608,N_1731);
nor U1933 (N_1933,N_1711,N_1705);
nand U1934 (N_1934,N_1717,N_1719);
nor U1935 (N_1935,N_1626,N_1787);
nand U1936 (N_1936,N_1656,N_1660);
nand U1937 (N_1937,N_1702,N_1790);
and U1938 (N_1938,N_1713,N_1761);
nor U1939 (N_1939,N_1629,N_1790);
or U1940 (N_1940,N_1600,N_1660);
nand U1941 (N_1941,N_1763,N_1788);
or U1942 (N_1942,N_1729,N_1675);
or U1943 (N_1943,N_1660,N_1608);
nand U1944 (N_1944,N_1622,N_1739);
nor U1945 (N_1945,N_1665,N_1695);
or U1946 (N_1946,N_1781,N_1726);
or U1947 (N_1947,N_1688,N_1721);
xnor U1948 (N_1948,N_1773,N_1762);
nand U1949 (N_1949,N_1655,N_1789);
and U1950 (N_1950,N_1775,N_1621);
nor U1951 (N_1951,N_1666,N_1657);
or U1952 (N_1952,N_1730,N_1763);
nand U1953 (N_1953,N_1687,N_1768);
nand U1954 (N_1954,N_1762,N_1602);
nor U1955 (N_1955,N_1627,N_1711);
or U1956 (N_1956,N_1666,N_1782);
nor U1957 (N_1957,N_1601,N_1656);
or U1958 (N_1958,N_1712,N_1614);
nand U1959 (N_1959,N_1680,N_1796);
nor U1960 (N_1960,N_1644,N_1652);
nand U1961 (N_1961,N_1623,N_1681);
nor U1962 (N_1962,N_1773,N_1606);
and U1963 (N_1963,N_1762,N_1742);
nor U1964 (N_1964,N_1683,N_1785);
nand U1965 (N_1965,N_1625,N_1717);
nand U1966 (N_1966,N_1642,N_1633);
or U1967 (N_1967,N_1625,N_1692);
nor U1968 (N_1968,N_1733,N_1648);
nor U1969 (N_1969,N_1738,N_1665);
nor U1970 (N_1970,N_1756,N_1753);
and U1971 (N_1971,N_1640,N_1725);
or U1972 (N_1972,N_1637,N_1705);
nor U1973 (N_1973,N_1737,N_1732);
nor U1974 (N_1974,N_1730,N_1729);
nand U1975 (N_1975,N_1706,N_1722);
nand U1976 (N_1976,N_1628,N_1617);
nor U1977 (N_1977,N_1701,N_1714);
nor U1978 (N_1978,N_1668,N_1712);
nor U1979 (N_1979,N_1604,N_1735);
nor U1980 (N_1980,N_1693,N_1772);
or U1981 (N_1981,N_1656,N_1715);
nor U1982 (N_1982,N_1670,N_1610);
nand U1983 (N_1983,N_1728,N_1629);
or U1984 (N_1984,N_1709,N_1726);
or U1985 (N_1985,N_1757,N_1726);
nand U1986 (N_1986,N_1731,N_1670);
nand U1987 (N_1987,N_1725,N_1615);
and U1988 (N_1988,N_1763,N_1683);
nor U1989 (N_1989,N_1627,N_1771);
nand U1990 (N_1990,N_1667,N_1614);
nand U1991 (N_1991,N_1636,N_1784);
nand U1992 (N_1992,N_1633,N_1605);
or U1993 (N_1993,N_1619,N_1621);
and U1994 (N_1994,N_1631,N_1726);
nor U1995 (N_1995,N_1740,N_1666);
nand U1996 (N_1996,N_1644,N_1705);
and U1997 (N_1997,N_1763,N_1700);
and U1998 (N_1998,N_1692,N_1683);
nand U1999 (N_1999,N_1603,N_1740);
nand U2000 (N_2000,N_1847,N_1821);
or U2001 (N_2001,N_1845,N_1964);
nand U2002 (N_2002,N_1841,N_1862);
nor U2003 (N_2003,N_1989,N_1979);
and U2004 (N_2004,N_1991,N_1816);
and U2005 (N_2005,N_1888,N_1887);
and U2006 (N_2006,N_1925,N_1891);
nor U2007 (N_2007,N_1952,N_1894);
nand U2008 (N_2008,N_1954,N_1871);
or U2009 (N_2009,N_1968,N_1992);
nor U2010 (N_2010,N_1839,N_1844);
nand U2011 (N_2011,N_1801,N_1958);
and U2012 (N_2012,N_1805,N_1988);
nand U2013 (N_2013,N_1961,N_1955);
nor U2014 (N_2014,N_1935,N_1865);
nand U2015 (N_2015,N_1949,N_1900);
or U2016 (N_2016,N_1851,N_1944);
nand U2017 (N_2017,N_1999,N_1902);
or U2018 (N_2018,N_1860,N_1885);
or U2019 (N_2019,N_1904,N_1922);
nand U2020 (N_2020,N_1933,N_1828);
or U2021 (N_2021,N_1923,N_1893);
nor U2022 (N_2022,N_1895,N_1946);
and U2023 (N_2023,N_1833,N_1863);
or U2024 (N_2024,N_1937,N_1882);
or U2025 (N_2025,N_1974,N_1864);
or U2026 (N_2026,N_1912,N_1875);
nor U2027 (N_2027,N_1826,N_1899);
nand U2028 (N_2028,N_1994,N_1921);
nand U2029 (N_2029,N_1982,N_1905);
or U2030 (N_2030,N_1919,N_1832);
and U2031 (N_2031,N_1971,N_1840);
nor U2032 (N_2032,N_1884,N_1890);
nand U2033 (N_2033,N_1948,N_1931);
or U2034 (N_2034,N_1854,N_1995);
nand U2035 (N_2035,N_1837,N_1870);
or U2036 (N_2036,N_1966,N_1858);
or U2037 (N_2037,N_1881,N_1872);
nor U2038 (N_2038,N_1812,N_1836);
nand U2039 (N_2039,N_1908,N_1956);
or U2040 (N_2040,N_1917,N_1907);
nand U2041 (N_2041,N_1803,N_1850);
and U2042 (N_2042,N_1848,N_1835);
nor U2043 (N_2043,N_1996,N_1975);
nand U2044 (N_2044,N_1957,N_1825);
or U2045 (N_2045,N_1943,N_1969);
and U2046 (N_2046,N_1879,N_1810);
nand U2047 (N_2047,N_1831,N_1906);
and U2048 (N_2048,N_1967,N_1852);
nand U2049 (N_2049,N_1874,N_1983);
nor U2050 (N_2050,N_1898,N_1834);
nor U2051 (N_2051,N_1903,N_1813);
nand U2052 (N_2052,N_1945,N_1824);
nand U2053 (N_2053,N_1911,N_1932);
nor U2054 (N_2054,N_1918,N_1978);
or U2055 (N_2055,N_1901,N_1942);
nor U2056 (N_2056,N_1953,N_1960);
nor U2057 (N_2057,N_1869,N_1827);
nor U2058 (N_2058,N_1990,N_1973);
nand U2059 (N_2059,N_1838,N_1986);
nand U2060 (N_2060,N_1926,N_1855);
or U2061 (N_2061,N_1897,N_1818);
nor U2062 (N_2062,N_1873,N_1963);
nor U2063 (N_2063,N_1846,N_1815);
and U2064 (N_2064,N_1814,N_1819);
and U2065 (N_2065,N_1951,N_1980);
and U2066 (N_2066,N_1843,N_1866);
nand U2067 (N_2067,N_1976,N_1886);
and U2068 (N_2068,N_1853,N_1861);
nor U2069 (N_2069,N_1808,N_1984);
and U2070 (N_2070,N_1962,N_1950);
nor U2071 (N_2071,N_1868,N_1823);
nor U2072 (N_2072,N_1941,N_1804);
and U2073 (N_2073,N_1809,N_1939);
or U2074 (N_2074,N_1830,N_1920);
nand U2075 (N_2075,N_1822,N_1889);
or U2076 (N_2076,N_1970,N_1998);
nor U2077 (N_2077,N_1820,N_1938);
or U2078 (N_2078,N_1997,N_1929);
or U2079 (N_2079,N_1806,N_1880);
nor U2080 (N_2080,N_1972,N_1977);
nor U2081 (N_2081,N_1981,N_1930);
or U2082 (N_2082,N_1924,N_1856);
and U2083 (N_2083,N_1892,N_1947);
nor U2084 (N_2084,N_1857,N_1910);
nor U2085 (N_2085,N_1987,N_1878);
and U2086 (N_2086,N_1940,N_1800);
and U2087 (N_2087,N_1993,N_1807);
nor U2088 (N_2088,N_1842,N_1909);
nand U2089 (N_2089,N_1934,N_1877);
nor U2090 (N_2090,N_1867,N_1916);
nor U2091 (N_2091,N_1829,N_1927);
or U2092 (N_2092,N_1883,N_1811);
or U2093 (N_2093,N_1985,N_1859);
nand U2094 (N_2094,N_1896,N_1876);
or U2095 (N_2095,N_1914,N_1936);
or U2096 (N_2096,N_1959,N_1913);
and U2097 (N_2097,N_1915,N_1849);
and U2098 (N_2098,N_1928,N_1802);
xnor U2099 (N_2099,N_1817,N_1965);
nand U2100 (N_2100,N_1849,N_1847);
nor U2101 (N_2101,N_1974,N_1928);
nor U2102 (N_2102,N_1854,N_1856);
and U2103 (N_2103,N_1993,N_1991);
or U2104 (N_2104,N_1833,N_1932);
and U2105 (N_2105,N_1929,N_1849);
and U2106 (N_2106,N_1903,N_1963);
nand U2107 (N_2107,N_1835,N_1958);
or U2108 (N_2108,N_1838,N_1957);
or U2109 (N_2109,N_1865,N_1879);
nand U2110 (N_2110,N_1859,N_1966);
and U2111 (N_2111,N_1978,N_1856);
nor U2112 (N_2112,N_1991,N_1810);
or U2113 (N_2113,N_1812,N_1973);
or U2114 (N_2114,N_1807,N_1871);
nand U2115 (N_2115,N_1902,N_1890);
and U2116 (N_2116,N_1875,N_1919);
nand U2117 (N_2117,N_1931,N_1995);
nor U2118 (N_2118,N_1822,N_1816);
nand U2119 (N_2119,N_1949,N_1807);
nor U2120 (N_2120,N_1852,N_1819);
and U2121 (N_2121,N_1826,N_1806);
nor U2122 (N_2122,N_1886,N_1848);
nor U2123 (N_2123,N_1871,N_1934);
nand U2124 (N_2124,N_1889,N_1838);
or U2125 (N_2125,N_1995,N_1901);
and U2126 (N_2126,N_1961,N_1883);
and U2127 (N_2127,N_1965,N_1904);
and U2128 (N_2128,N_1953,N_1966);
or U2129 (N_2129,N_1902,N_1985);
or U2130 (N_2130,N_1930,N_1887);
nand U2131 (N_2131,N_1819,N_1868);
and U2132 (N_2132,N_1904,N_1837);
nor U2133 (N_2133,N_1966,N_1838);
and U2134 (N_2134,N_1923,N_1826);
or U2135 (N_2135,N_1843,N_1932);
and U2136 (N_2136,N_1864,N_1807);
nor U2137 (N_2137,N_1829,N_1824);
or U2138 (N_2138,N_1839,N_1928);
and U2139 (N_2139,N_1954,N_1814);
or U2140 (N_2140,N_1831,N_1841);
or U2141 (N_2141,N_1844,N_1879);
nand U2142 (N_2142,N_1833,N_1866);
nand U2143 (N_2143,N_1914,N_1945);
nor U2144 (N_2144,N_1838,N_1813);
nor U2145 (N_2145,N_1805,N_1857);
nor U2146 (N_2146,N_1866,N_1948);
and U2147 (N_2147,N_1932,N_1944);
nand U2148 (N_2148,N_1829,N_1942);
nand U2149 (N_2149,N_1899,N_1948);
nand U2150 (N_2150,N_1960,N_1823);
nor U2151 (N_2151,N_1940,N_1805);
or U2152 (N_2152,N_1919,N_1819);
and U2153 (N_2153,N_1899,N_1846);
nor U2154 (N_2154,N_1871,N_1935);
or U2155 (N_2155,N_1908,N_1971);
nor U2156 (N_2156,N_1986,N_1969);
or U2157 (N_2157,N_1942,N_1918);
and U2158 (N_2158,N_1840,N_1808);
or U2159 (N_2159,N_1803,N_1835);
or U2160 (N_2160,N_1893,N_1874);
nand U2161 (N_2161,N_1894,N_1980);
nor U2162 (N_2162,N_1901,N_1994);
or U2163 (N_2163,N_1975,N_1847);
xor U2164 (N_2164,N_1934,N_1942);
or U2165 (N_2165,N_1847,N_1995);
nor U2166 (N_2166,N_1825,N_1895);
and U2167 (N_2167,N_1820,N_1933);
nand U2168 (N_2168,N_1909,N_1874);
nor U2169 (N_2169,N_1865,N_1902);
nand U2170 (N_2170,N_1948,N_1831);
nor U2171 (N_2171,N_1808,N_1852);
nand U2172 (N_2172,N_1851,N_1930);
and U2173 (N_2173,N_1925,N_1991);
nor U2174 (N_2174,N_1949,N_1874);
or U2175 (N_2175,N_1927,N_1807);
nand U2176 (N_2176,N_1901,N_1922);
nor U2177 (N_2177,N_1905,N_1872);
nand U2178 (N_2178,N_1992,N_1961);
nor U2179 (N_2179,N_1979,N_1904);
nor U2180 (N_2180,N_1892,N_1845);
nand U2181 (N_2181,N_1876,N_1850);
or U2182 (N_2182,N_1998,N_1905);
nand U2183 (N_2183,N_1836,N_1908);
nor U2184 (N_2184,N_1920,N_1894);
xor U2185 (N_2185,N_1966,N_1964);
or U2186 (N_2186,N_1901,N_1887);
nand U2187 (N_2187,N_1898,N_1922);
nor U2188 (N_2188,N_1944,N_1961);
or U2189 (N_2189,N_1905,N_1980);
or U2190 (N_2190,N_1861,N_1900);
or U2191 (N_2191,N_1857,N_1875);
nor U2192 (N_2192,N_1818,N_1876);
nor U2193 (N_2193,N_1991,N_1934);
and U2194 (N_2194,N_1904,N_1853);
and U2195 (N_2195,N_1976,N_1985);
nand U2196 (N_2196,N_1828,N_1974);
nand U2197 (N_2197,N_1840,N_1861);
or U2198 (N_2198,N_1945,N_1858);
nand U2199 (N_2199,N_1965,N_1892);
or U2200 (N_2200,N_2080,N_2046);
or U2201 (N_2201,N_2115,N_2096);
nor U2202 (N_2202,N_2154,N_2091);
nor U2203 (N_2203,N_2076,N_2001);
and U2204 (N_2204,N_2053,N_2125);
and U2205 (N_2205,N_2108,N_2127);
or U2206 (N_2206,N_2140,N_2195);
nand U2207 (N_2207,N_2089,N_2132);
nor U2208 (N_2208,N_2134,N_2184);
nor U2209 (N_2209,N_2114,N_2094);
or U2210 (N_2210,N_2043,N_2121);
nand U2211 (N_2211,N_2181,N_2050);
or U2212 (N_2212,N_2088,N_2017);
or U2213 (N_2213,N_2015,N_2042);
or U2214 (N_2214,N_2104,N_2130);
xor U2215 (N_2215,N_2009,N_2155);
nor U2216 (N_2216,N_2179,N_2090);
and U2217 (N_2217,N_2072,N_2193);
or U2218 (N_2218,N_2049,N_2145);
or U2219 (N_2219,N_2185,N_2178);
nand U2220 (N_2220,N_2141,N_2086);
or U2221 (N_2221,N_2191,N_2031);
nand U2222 (N_2222,N_2033,N_2014);
or U2223 (N_2223,N_2190,N_2167);
nand U2224 (N_2224,N_2133,N_2016);
and U2225 (N_2225,N_2162,N_2047);
and U2226 (N_2226,N_2028,N_2002);
nand U2227 (N_2227,N_2194,N_2171);
nor U2228 (N_2228,N_2095,N_2135);
nor U2229 (N_2229,N_2119,N_2146);
or U2230 (N_2230,N_2112,N_2144);
nand U2231 (N_2231,N_2077,N_2150);
and U2232 (N_2232,N_2105,N_2153);
or U2233 (N_2233,N_2111,N_2169);
nor U2234 (N_2234,N_2055,N_2142);
nor U2235 (N_2235,N_2052,N_2018);
or U2236 (N_2236,N_2068,N_2092);
or U2237 (N_2237,N_2093,N_2000);
and U2238 (N_2238,N_2138,N_2157);
nand U2239 (N_2239,N_2098,N_2066);
nor U2240 (N_2240,N_2174,N_2177);
nand U2241 (N_2241,N_2054,N_2026);
nor U2242 (N_2242,N_2180,N_2136);
nand U2243 (N_2243,N_2170,N_2041);
nor U2244 (N_2244,N_2034,N_2152);
nand U2245 (N_2245,N_2126,N_2020);
and U2246 (N_2246,N_2165,N_2058);
and U2247 (N_2247,N_2023,N_2060);
and U2248 (N_2248,N_2074,N_2101);
nor U2249 (N_2249,N_2137,N_2122);
or U2250 (N_2250,N_2045,N_2061);
nor U2251 (N_2251,N_2097,N_2063);
or U2252 (N_2252,N_2004,N_2024);
and U2253 (N_2253,N_2118,N_2128);
nor U2254 (N_2254,N_2120,N_2083);
and U2255 (N_2255,N_2071,N_2005);
nor U2256 (N_2256,N_2164,N_2019);
nor U2257 (N_2257,N_2188,N_2069);
nand U2258 (N_2258,N_2064,N_2021);
or U2259 (N_2259,N_2149,N_2187);
and U2260 (N_2260,N_2124,N_2100);
or U2261 (N_2261,N_2166,N_2197);
and U2262 (N_2262,N_2196,N_2029);
nand U2263 (N_2263,N_2182,N_2078);
nand U2264 (N_2264,N_2160,N_2148);
or U2265 (N_2265,N_2139,N_2102);
and U2266 (N_2266,N_2051,N_2147);
or U2267 (N_2267,N_2082,N_2107);
nor U2268 (N_2268,N_2032,N_2013);
and U2269 (N_2269,N_2070,N_2109);
or U2270 (N_2270,N_2151,N_2073);
nand U2271 (N_2271,N_2106,N_2161);
nor U2272 (N_2272,N_2159,N_2006);
nor U2273 (N_2273,N_2065,N_2036);
and U2274 (N_2274,N_2199,N_2099);
nor U2275 (N_2275,N_2123,N_2173);
nand U2276 (N_2276,N_2044,N_2131);
and U2277 (N_2277,N_2116,N_2038);
nand U2278 (N_2278,N_2183,N_2030);
and U2279 (N_2279,N_2010,N_2176);
nor U2280 (N_2280,N_2039,N_2012);
or U2281 (N_2281,N_2156,N_2084);
and U2282 (N_2282,N_2056,N_2113);
nand U2283 (N_2283,N_2025,N_2067);
xor U2284 (N_2284,N_2003,N_2079);
nand U2285 (N_2285,N_2168,N_2037);
xnor U2286 (N_2286,N_2163,N_2008);
nand U2287 (N_2287,N_2129,N_2007);
nor U2288 (N_2288,N_2035,N_2198);
and U2289 (N_2289,N_2175,N_2040);
nand U2290 (N_2290,N_2075,N_2103);
and U2291 (N_2291,N_2057,N_2027);
and U2292 (N_2292,N_2081,N_2110);
and U2293 (N_2293,N_2117,N_2059);
and U2294 (N_2294,N_2048,N_2085);
nand U2295 (N_2295,N_2011,N_2186);
nand U2296 (N_2296,N_2022,N_2143);
or U2297 (N_2297,N_2172,N_2189);
nor U2298 (N_2298,N_2158,N_2087);
nor U2299 (N_2299,N_2192,N_2062);
xor U2300 (N_2300,N_2083,N_2140);
nor U2301 (N_2301,N_2039,N_2069);
or U2302 (N_2302,N_2000,N_2047);
and U2303 (N_2303,N_2047,N_2036);
nor U2304 (N_2304,N_2116,N_2027);
and U2305 (N_2305,N_2066,N_2190);
nor U2306 (N_2306,N_2120,N_2096);
or U2307 (N_2307,N_2090,N_2125);
or U2308 (N_2308,N_2146,N_2133);
nand U2309 (N_2309,N_2002,N_2095);
nor U2310 (N_2310,N_2059,N_2165);
or U2311 (N_2311,N_2130,N_2119);
and U2312 (N_2312,N_2094,N_2035);
nor U2313 (N_2313,N_2109,N_2055);
nand U2314 (N_2314,N_2122,N_2140);
nand U2315 (N_2315,N_2191,N_2030);
or U2316 (N_2316,N_2188,N_2181);
nor U2317 (N_2317,N_2055,N_2077);
or U2318 (N_2318,N_2096,N_2124);
nor U2319 (N_2319,N_2126,N_2059);
or U2320 (N_2320,N_2198,N_2038);
nor U2321 (N_2321,N_2051,N_2115);
and U2322 (N_2322,N_2172,N_2099);
nand U2323 (N_2323,N_2127,N_2088);
nor U2324 (N_2324,N_2012,N_2026);
nor U2325 (N_2325,N_2011,N_2058);
or U2326 (N_2326,N_2020,N_2012);
nor U2327 (N_2327,N_2151,N_2022);
and U2328 (N_2328,N_2066,N_2062);
or U2329 (N_2329,N_2142,N_2002);
nor U2330 (N_2330,N_2169,N_2020);
or U2331 (N_2331,N_2091,N_2123);
and U2332 (N_2332,N_2006,N_2136);
nand U2333 (N_2333,N_2033,N_2192);
nor U2334 (N_2334,N_2122,N_2067);
or U2335 (N_2335,N_2050,N_2164);
or U2336 (N_2336,N_2018,N_2105);
or U2337 (N_2337,N_2082,N_2043);
and U2338 (N_2338,N_2063,N_2002);
xnor U2339 (N_2339,N_2167,N_2120);
nor U2340 (N_2340,N_2039,N_2022);
nor U2341 (N_2341,N_2100,N_2000);
or U2342 (N_2342,N_2072,N_2079);
nand U2343 (N_2343,N_2141,N_2150);
and U2344 (N_2344,N_2197,N_2008);
or U2345 (N_2345,N_2045,N_2003);
nor U2346 (N_2346,N_2169,N_2178);
nor U2347 (N_2347,N_2153,N_2096);
and U2348 (N_2348,N_2042,N_2117);
nand U2349 (N_2349,N_2077,N_2146);
and U2350 (N_2350,N_2036,N_2117);
and U2351 (N_2351,N_2104,N_2180);
or U2352 (N_2352,N_2097,N_2109);
and U2353 (N_2353,N_2115,N_2183);
and U2354 (N_2354,N_2044,N_2165);
nand U2355 (N_2355,N_2155,N_2007);
or U2356 (N_2356,N_2113,N_2024);
nand U2357 (N_2357,N_2025,N_2007);
and U2358 (N_2358,N_2063,N_2102);
nor U2359 (N_2359,N_2177,N_2028);
and U2360 (N_2360,N_2055,N_2108);
nand U2361 (N_2361,N_2110,N_2018);
and U2362 (N_2362,N_2059,N_2047);
nor U2363 (N_2363,N_2170,N_2115);
or U2364 (N_2364,N_2062,N_2103);
and U2365 (N_2365,N_2153,N_2091);
and U2366 (N_2366,N_2182,N_2095);
and U2367 (N_2367,N_2100,N_2120);
nor U2368 (N_2368,N_2153,N_2115);
and U2369 (N_2369,N_2108,N_2185);
or U2370 (N_2370,N_2030,N_2037);
nor U2371 (N_2371,N_2104,N_2115);
nand U2372 (N_2372,N_2178,N_2189);
nor U2373 (N_2373,N_2082,N_2115);
nor U2374 (N_2374,N_2139,N_2002);
and U2375 (N_2375,N_2140,N_2044);
and U2376 (N_2376,N_2175,N_2019);
or U2377 (N_2377,N_2084,N_2146);
and U2378 (N_2378,N_2102,N_2045);
or U2379 (N_2379,N_2108,N_2085);
nand U2380 (N_2380,N_2198,N_2192);
nor U2381 (N_2381,N_2092,N_2184);
nor U2382 (N_2382,N_2016,N_2127);
nor U2383 (N_2383,N_2161,N_2170);
and U2384 (N_2384,N_2043,N_2164);
and U2385 (N_2385,N_2118,N_2081);
and U2386 (N_2386,N_2076,N_2158);
or U2387 (N_2387,N_2050,N_2026);
nor U2388 (N_2388,N_2082,N_2076);
and U2389 (N_2389,N_2082,N_2124);
nand U2390 (N_2390,N_2016,N_2001);
nor U2391 (N_2391,N_2151,N_2039);
nand U2392 (N_2392,N_2158,N_2081);
nor U2393 (N_2393,N_2068,N_2189);
nand U2394 (N_2394,N_2135,N_2171);
nand U2395 (N_2395,N_2073,N_2024);
and U2396 (N_2396,N_2157,N_2137);
nand U2397 (N_2397,N_2199,N_2159);
and U2398 (N_2398,N_2080,N_2054);
nor U2399 (N_2399,N_2028,N_2064);
or U2400 (N_2400,N_2221,N_2390);
nand U2401 (N_2401,N_2245,N_2317);
nor U2402 (N_2402,N_2273,N_2217);
nor U2403 (N_2403,N_2363,N_2206);
or U2404 (N_2404,N_2235,N_2391);
xnor U2405 (N_2405,N_2253,N_2200);
nor U2406 (N_2406,N_2352,N_2241);
nand U2407 (N_2407,N_2215,N_2214);
nor U2408 (N_2408,N_2308,N_2236);
or U2409 (N_2409,N_2271,N_2355);
nand U2410 (N_2410,N_2329,N_2290);
or U2411 (N_2411,N_2367,N_2321);
nand U2412 (N_2412,N_2396,N_2387);
nand U2413 (N_2413,N_2399,N_2263);
or U2414 (N_2414,N_2294,N_2288);
nand U2415 (N_2415,N_2371,N_2335);
or U2416 (N_2416,N_2356,N_2372);
nor U2417 (N_2417,N_2219,N_2323);
nor U2418 (N_2418,N_2347,N_2333);
nand U2419 (N_2419,N_2257,N_2362);
and U2420 (N_2420,N_2346,N_2305);
and U2421 (N_2421,N_2260,N_2315);
and U2422 (N_2422,N_2274,N_2278);
nor U2423 (N_2423,N_2327,N_2303);
nor U2424 (N_2424,N_2341,N_2351);
nor U2425 (N_2425,N_2208,N_2272);
and U2426 (N_2426,N_2311,N_2330);
and U2427 (N_2427,N_2234,N_2336);
and U2428 (N_2428,N_2345,N_2324);
nand U2429 (N_2429,N_2384,N_2275);
or U2430 (N_2430,N_2220,N_2310);
or U2431 (N_2431,N_2285,N_2366);
nor U2432 (N_2432,N_2360,N_2226);
or U2433 (N_2433,N_2368,N_2279);
nand U2434 (N_2434,N_2377,N_2261);
nor U2435 (N_2435,N_2250,N_2344);
nor U2436 (N_2436,N_2238,N_2232);
and U2437 (N_2437,N_2316,N_2291);
nand U2438 (N_2438,N_2281,N_2201);
nand U2439 (N_2439,N_2223,N_2301);
nand U2440 (N_2440,N_2252,N_2216);
and U2441 (N_2441,N_2386,N_2332);
nand U2442 (N_2442,N_2262,N_2202);
or U2443 (N_2443,N_2348,N_2313);
and U2444 (N_2444,N_2296,N_2394);
and U2445 (N_2445,N_2339,N_2358);
nor U2446 (N_2446,N_2342,N_2318);
nand U2447 (N_2447,N_2211,N_2283);
nor U2448 (N_2448,N_2375,N_2205);
nor U2449 (N_2449,N_2293,N_2269);
nor U2450 (N_2450,N_2383,N_2388);
nand U2451 (N_2451,N_2210,N_2298);
nand U2452 (N_2452,N_2254,N_2282);
and U2453 (N_2453,N_2304,N_2231);
nand U2454 (N_2454,N_2277,N_2230);
nor U2455 (N_2455,N_2349,N_2343);
nor U2456 (N_2456,N_2379,N_2292);
and U2457 (N_2457,N_2338,N_2392);
or U2458 (N_2458,N_2328,N_2256);
nor U2459 (N_2459,N_2204,N_2381);
nand U2460 (N_2460,N_2228,N_2354);
or U2461 (N_2461,N_2237,N_2264);
nand U2462 (N_2462,N_2255,N_2259);
or U2463 (N_2463,N_2306,N_2370);
and U2464 (N_2464,N_2307,N_2244);
nor U2465 (N_2465,N_2326,N_2225);
nor U2466 (N_2466,N_2287,N_2337);
nor U2467 (N_2467,N_2268,N_2276);
and U2468 (N_2468,N_2364,N_2212);
or U2469 (N_2469,N_2209,N_2251);
or U2470 (N_2470,N_2397,N_2249);
nor U2471 (N_2471,N_2395,N_2295);
or U2472 (N_2472,N_2340,N_2243);
or U2473 (N_2473,N_2297,N_2203);
nor U2474 (N_2474,N_2289,N_2380);
and U2475 (N_2475,N_2258,N_2227);
nor U2476 (N_2476,N_2247,N_2365);
nor U2477 (N_2477,N_2229,N_2331);
and U2478 (N_2478,N_2334,N_2312);
and U2479 (N_2479,N_2361,N_2300);
nor U2480 (N_2480,N_2314,N_2373);
nand U2481 (N_2481,N_2302,N_2393);
and U2482 (N_2482,N_2246,N_2322);
or U2483 (N_2483,N_2248,N_2218);
nand U2484 (N_2484,N_2378,N_2350);
or U2485 (N_2485,N_2239,N_2374);
nand U2486 (N_2486,N_2398,N_2266);
nor U2487 (N_2487,N_2286,N_2207);
nand U2488 (N_2488,N_2357,N_2382);
nor U2489 (N_2489,N_2222,N_2325);
nor U2490 (N_2490,N_2242,N_2280);
nand U2491 (N_2491,N_2240,N_2284);
and U2492 (N_2492,N_2389,N_2385);
and U2493 (N_2493,N_2213,N_2376);
or U2494 (N_2494,N_2319,N_2265);
nor U2495 (N_2495,N_2224,N_2320);
nor U2496 (N_2496,N_2267,N_2299);
nor U2497 (N_2497,N_2353,N_2309);
nor U2498 (N_2498,N_2359,N_2369);
or U2499 (N_2499,N_2233,N_2270);
nor U2500 (N_2500,N_2322,N_2282);
nand U2501 (N_2501,N_2239,N_2294);
and U2502 (N_2502,N_2246,N_2218);
or U2503 (N_2503,N_2335,N_2316);
or U2504 (N_2504,N_2222,N_2200);
and U2505 (N_2505,N_2267,N_2224);
and U2506 (N_2506,N_2379,N_2394);
and U2507 (N_2507,N_2274,N_2349);
nand U2508 (N_2508,N_2394,N_2362);
and U2509 (N_2509,N_2378,N_2365);
nand U2510 (N_2510,N_2376,N_2311);
or U2511 (N_2511,N_2288,N_2303);
and U2512 (N_2512,N_2240,N_2204);
and U2513 (N_2513,N_2260,N_2294);
nand U2514 (N_2514,N_2293,N_2317);
and U2515 (N_2515,N_2240,N_2273);
nand U2516 (N_2516,N_2391,N_2378);
or U2517 (N_2517,N_2312,N_2226);
nand U2518 (N_2518,N_2318,N_2385);
nor U2519 (N_2519,N_2301,N_2381);
and U2520 (N_2520,N_2214,N_2229);
nand U2521 (N_2521,N_2363,N_2343);
nand U2522 (N_2522,N_2220,N_2337);
or U2523 (N_2523,N_2279,N_2260);
nor U2524 (N_2524,N_2258,N_2344);
nor U2525 (N_2525,N_2222,N_2249);
nand U2526 (N_2526,N_2387,N_2283);
nor U2527 (N_2527,N_2309,N_2362);
nor U2528 (N_2528,N_2308,N_2328);
nor U2529 (N_2529,N_2315,N_2326);
and U2530 (N_2530,N_2220,N_2383);
nor U2531 (N_2531,N_2249,N_2235);
and U2532 (N_2532,N_2221,N_2306);
or U2533 (N_2533,N_2292,N_2294);
and U2534 (N_2534,N_2308,N_2348);
and U2535 (N_2535,N_2382,N_2269);
or U2536 (N_2536,N_2309,N_2371);
and U2537 (N_2537,N_2312,N_2278);
and U2538 (N_2538,N_2202,N_2387);
and U2539 (N_2539,N_2333,N_2308);
nand U2540 (N_2540,N_2335,N_2363);
and U2541 (N_2541,N_2326,N_2324);
or U2542 (N_2542,N_2273,N_2225);
or U2543 (N_2543,N_2264,N_2236);
nor U2544 (N_2544,N_2386,N_2227);
and U2545 (N_2545,N_2292,N_2284);
nand U2546 (N_2546,N_2263,N_2364);
or U2547 (N_2547,N_2200,N_2391);
nor U2548 (N_2548,N_2276,N_2377);
nand U2549 (N_2549,N_2206,N_2310);
nor U2550 (N_2550,N_2274,N_2231);
nor U2551 (N_2551,N_2382,N_2347);
nor U2552 (N_2552,N_2350,N_2302);
or U2553 (N_2553,N_2281,N_2230);
nand U2554 (N_2554,N_2335,N_2391);
or U2555 (N_2555,N_2261,N_2220);
nor U2556 (N_2556,N_2277,N_2395);
and U2557 (N_2557,N_2303,N_2252);
and U2558 (N_2558,N_2260,N_2320);
nand U2559 (N_2559,N_2310,N_2271);
and U2560 (N_2560,N_2383,N_2267);
nand U2561 (N_2561,N_2324,N_2256);
nand U2562 (N_2562,N_2207,N_2365);
or U2563 (N_2563,N_2262,N_2272);
or U2564 (N_2564,N_2290,N_2340);
xor U2565 (N_2565,N_2315,N_2374);
or U2566 (N_2566,N_2282,N_2210);
xor U2567 (N_2567,N_2345,N_2344);
nor U2568 (N_2568,N_2306,N_2373);
and U2569 (N_2569,N_2245,N_2251);
nor U2570 (N_2570,N_2212,N_2355);
or U2571 (N_2571,N_2220,N_2222);
or U2572 (N_2572,N_2347,N_2201);
and U2573 (N_2573,N_2202,N_2383);
or U2574 (N_2574,N_2393,N_2297);
or U2575 (N_2575,N_2253,N_2297);
nand U2576 (N_2576,N_2397,N_2272);
nand U2577 (N_2577,N_2209,N_2243);
nand U2578 (N_2578,N_2346,N_2292);
or U2579 (N_2579,N_2218,N_2331);
and U2580 (N_2580,N_2203,N_2367);
nor U2581 (N_2581,N_2325,N_2341);
nor U2582 (N_2582,N_2333,N_2221);
or U2583 (N_2583,N_2316,N_2211);
and U2584 (N_2584,N_2381,N_2231);
nand U2585 (N_2585,N_2261,N_2212);
and U2586 (N_2586,N_2338,N_2232);
nor U2587 (N_2587,N_2206,N_2341);
and U2588 (N_2588,N_2214,N_2294);
nor U2589 (N_2589,N_2224,N_2246);
or U2590 (N_2590,N_2355,N_2334);
and U2591 (N_2591,N_2365,N_2238);
or U2592 (N_2592,N_2371,N_2397);
nor U2593 (N_2593,N_2212,N_2385);
xnor U2594 (N_2594,N_2253,N_2266);
and U2595 (N_2595,N_2321,N_2338);
and U2596 (N_2596,N_2257,N_2370);
or U2597 (N_2597,N_2246,N_2200);
nor U2598 (N_2598,N_2289,N_2286);
and U2599 (N_2599,N_2271,N_2354);
and U2600 (N_2600,N_2585,N_2562);
nand U2601 (N_2601,N_2404,N_2432);
or U2602 (N_2602,N_2401,N_2575);
and U2603 (N_2603,N_2477,N_2516);
nand U2604 (N_2604,N_2539,N_2545);
and U2605 (N_2605,N_2510,N_2424);
nor U2606 (N_2606,N_2472,N_2578);
and U2607 (N_2607,N_2487,N_2568);
and U2608 (N_2608,N_2534,N_2447);
and U2609 (N_2609,N_2513,N_2490);
and U2610 (N_2610,N_2553,N_2485);
and U2611 (N_2611,N_2451,N_2535);
nor U2612 (N_2612,N_2426,N_2584);
nor U2613 (N_2613,N_2457,N_2446);
nand U2614 (N_2614,N_2528,N_2467);
nand U2615 (N_2615,N_2583,N_2420);
nand U2616 (N_2616,N_2500,N_2549);
or U2617 (N_2617,N_2461,N_2517);
xor U2618 (N_2618,N_2544,N_2418);
or U2619 (N_2619,N_2499,N_2514);
nor U2620 (N_2620,N_2559,N_2589);
nand U2621 (N_2621,N_2430,N_2458);
nor U2622 (N_2622,N_2492,N_2483);
nand U2623 (N_2623,N_2577,N_2591);
and U2624 (N_2624,N_2557,N_2422);
and U2625 (N_2625,N_2501,N_2419);
nand U2626 (N_2626,N_2541,N_2521);
nor U2627 (N_2627,N_2507,N_2470);
xor U2628 (N_2628,N_2405,N_2596);
nand U2629 (N_2629,N_2561,N_2480);
or U2630 (N_2630,N_2569,N_2427);
and U2631 (N_2631,N_2506,N_2538);
nand U2632 (N_2632,N_2403,N_2491);
nand U2633 (N_2633,N_2504,N_2524);
or U2634 (N_2634,N_2421,N_2548);
nand U2635 (N_2635,N_2408,N_2508);
or U2636 (N_2636,N_2522,N_2592);
nor U2637 (N_2637,N_2416,N_2540);
or U2638 (N_2638,N_2462,N_2448);
or U2639 (N_2639,N_2465,N_2529);
nor U2640 (N_2640,N_2429,N_2414);
nor U2641 (N_2641,N_2460,N_2512);
and U2642 (N_2642,N_2459,N_2594);
or U2643 (N_2643,N_2558,N_2597);
nor U2644 (N_2644,N_2590,N_2471);
nand U2645 (N_2645,N_2431,N_2527);
or U2646 (N_2646,N_2482,N_2413);
nand U2647 (N_2647,N_2473,N_2515);
and U2648 (N_2648,N_2475,N_2518);
and U2649 (N_2649,N_2536,N_2478);
and U2650 (N_2650,N_2556,N_2481);
or U2651 (N_2651,N_2574,N_2455);
or U2652 (N_2652,N_2464,N_2417);
and U2653 (N_2653,N_2494,N_2571);
or U2654 (N_2654,N_2407,N_2443);
nor U2655 (N_2655,N_2402,N_2442);
nor U2656 (N_2656,N_2488,N_2511);
and U2657 (N_2657,N_2463,N_2576);
nand U2658 (N_2658,N_2554,N_2573);
or U2659 (N_2659,N_2476,N_2532);
xor U2660 (N_2660,N_2452,N_2587);
nor U2661 (N_2661,N_2555,N_2497);
nand U2662 (N_2662,N_2546,N_2474);
or U2663 (N_2663,N_2599,N_2437);
and U2664 (N_2664,N_2531,N_2560);
and U2665 (N_2665,N_2469,N_2406);
nand U2666 (N_2666,N_2409,N_2533);
or U2667 (N_2667,N_2410,N_2543);
nand U2668 (N_2668,N_2412,N_2493);
nor U2669 (N_2669,N_2439,N_2440);
and U2670 (N_2670,N_2550,N_2456);
nand U2671 (N_2671,N_2595,N_2593);
nand U2672 (N_2672,N_2503,N_2566);
nor U2673 (N_2673,N_2441,N_2580);
or U2674 (N_2674,N_2425,N_2423);
or U2675 (N_2675,N_2509,N_2411);
or U2676 (N_2676,N_2453,N_2496);
nor U2677 (N_2677,N_2454,N_2530);
nand U2678 (N_2678,N_2433,N_2435);
nand U2679 (N_2679,N_2498,N_2449);
and U2680 (N_2680,N_2466,N_2495);
and U2681 (N_2681,N_2434,N_2523);
nand U2682 (N_2682,N_2547,N_2598);
nand U2683 (N_2683,N_2563,N_2525);
nand U2684 (N_2684,N_2486,N_2520);
nor U2685 (N_2685,N_2570,N_2551);
or U2686 (N_2686,N_2586,N_2489);
and U2687 (N_2687,N_2502,N_2505);
or U2688 (N_2688,N_2400,N_2519);
nor U2689 (N_2689,N_2436,N_2415);
or U2690 (N_2690,N_2450,N_2428);
nor U2691 (N_2691,N_2572,N_2542);
nor U2692 (N_2692,N_2484,N_2588);
nand U2693 (N_2693,N_2445,N_2438);
nor U2694 (N_2694,N_2567,N_2552);
or U2695 (N_2695,N_2581,N_2526);
and U2696 (N_2696,N_2468,N_2564);
nand U2697 (N_2697,N_2565,N_2582);
nor U2698 (N_2698,N_2479,N_2537);
or U2699 (N_2699,N_2579,N_2444);
and U2700 (N_2700,N_2506,N_2576);
nand U2701 (N_2701,N_2483,N_2434);
nand U2702 (N_2702,N_2579,N_2536);
nand U2703 (N_2703,N_2534,N_2564);
nor U2704 (N_2704,N_2495,N_2585);
or U2705 (N_2705,N_2594,N_2581);
nand U2706 (N_2706,N_2492,N_2498);
or U2707 (N_2707,N_2454,N_2521);
nand U2708 (N_2708,N_2481,N_2577);
nor U2709 (N_2709,N_2555,N_2469);
or U2710 (N_2710,N_2555,N_2482);
nor U2711 (N_2711,N_2409,N_2413);
or U2712 (N_2712,N_2443,N_2402);
or U2713 (N_2713,N_2522,N_2428);
nand U2714 (N_2714,N_2566,N_2587);
nor U2715 (N_2715,N_2494,N_2596);
nand U2716 (N_2716,N_2426,N_2506);
nor U2717 (N_2717,N_2551,N_2504);
xor U2718 (N_2718,N_2547,N_2456);
and U2719 (N_2719,N_2460,N_2430);
nand U2720 (N_2720,N_2475,N_2598);
nor U2721 (N_2721,N_2456,N_2421);
nor U2722 (N_2722,N_2535,N_2522);
or U2723 (N_2723,N_2516,N_2424);
and U2724 (N_2724,N_2537,N_2554);
nor U2725 (N_2725,N_2447,N_2491);
and U2726 (N_2726,N_2426,N_2421);
nor U2727 (N_2727,N_2585,N_2450);
nand U2728 (N_2728,N_2558,N_2427);
nor U2729 (N_2729,N_2519,N_2441);
or U2730 (N_2730,N_2522,N_2550);
or U2731 (N_2731,N_2530,N_2574);
or U2732 (N_2732,N_2547,N_2481);
and U2733 (N_2733,N_2506,N_2479);
nand U2734 (N_2734,N_2469,N_2552);
and U2735 (N_2735,N_2516,N_2489);
nor U2736 (N_2736,N_2481,N_2434);
nor U2737 (N_2737,N_2442,N_2423);
or U2738 (N_2738,N_2560,N_2407);
and U2739 (N_2739,N_2408,N_2584);
nor U2740 (N_2740,N_2437,N_2548);
nor U2741 (N_2741,N_2411,N_2534);
or U2742 (N_2742,N_2529,N_2536);
nand U2743 (N_2743,N_2449,N_2430);
nand U2744 (N_2744,N_2474,N_2431);
and U2745 (N_2745,N_2593,N_2470);
nor U2746 (N_2746,N_2568,N_2452);
and U2747 (N_2747,N_2409,N_2461);
nand U2748 (N_2748,N_2569,N_2424);
nor U2749 (N_2749,N_2502,N_2570);
nand U2750 (N_2750,N_2497,N_2589);
or U2751 (N_2751,N_2409,N_2452);
nor U2752 (N_2752,N_2412,N_2463);
or U2753 (N_2753,N_2460,N_2486);
nor U2754 (N_2754,N_2444,N_2466);
and U2755 (N_2755,N_2501,N_2462);
nand U2756 (N_2756,N_2477,N_2569);
and U2757 (N_2757,N_2536,N_2493);
and U2758 (N_2758,N_2473,N_2537);
or U2759 (N_2759,N_2471,N_2512);
nor U2760 (N_2760,N_2595,N_2479);
nand U2761 (N_2761,N_2443,N_2560);
and U2762 (N_2762,N_2478,N_2544);
and U2763 (N_2763,N_2530,N_2491);
nor U2764 (N_2764,N_2495,N_2584);
or U2765 (N_2765,N_2483,N_2510);
and U2766 (N_2766,N_2476,N_2400);
nor U2767 (N_2767,N_2560,N_2500);
nor U2768 (N_2768,N_2489,N_2569);
and U2769 (N_2769,N_2490,N_2594);
or U2770 (N_2770,N_2499,N_2442);
or U2771 (N_2771,N_2535,N_2532);
nand U2772 (N_2772,N_2467,N_2445);
nand U2773 (N_2773,N_2556,N_2523);
and U2774 (N_2774,N_2584,N_2436);
and U2775 (N_2775,N_2481,N_2591);
xor U2776 (N_2776,N_2524,N_2480);
or U2777 (N_2777,N_2558,N_2570);
nand U2778 (N_2778,N_2496,N_2533);
and U2779 (N_2779,N_2474,N_2536);
nand U2780 (N_2780,N_2531,N_2586);
nand U2781 (N_2781,N_2526,N_2458);
or U2782 (N_2782,N_2406,N_2571);
or U2783 (N_2783,N_2586,N_2444);
and U2784 (N_2784,N_2571,N_2557);
nand U2785 (N_2785,N_2463,N_2555);
and U2786 (N_2786,N_2436,N_2595);
nor U2787 (N_2787,N_2443,N_2425);
and U2788 (N_2788,N_2572,N_2538);
nand U2789 (N_2789,N_2412,N_2445);
and U2790 (N_2790,N_2461,N_2542);
nor U2791 (N_2791,N_2429,N_2431);
or U2792 (N_2792,N_2412,N_2415);
and U2793 (N_2793,N_2512,N_2502);
nand U2794 (N_2794,N_2593,N_2437);
nor U2795 (N_2795,N_2466,N_2525);
nor U2796 (N_2796,N_2491,N_2534);
nor U2797 (N_2797,N_2515,N_2571);
and U2798 (N_2798,N_2580,N_2489);
or U2799 (N_2799,N_2580,N_2494);
nand U2800 (N_2800,N_2791,N_2737);
nor U2801 (N_2801,N_2674,N_2738);
xnor U2802 (N_2802,N_2656,N_2788);
and U2803 (N_2803,N_2729,N_2694);
or U2804 (N_2804,N_2723,N_2635);
nor U2805 (N_2805,N_2797,N_2643);
nor U2806 (N_2806,N_2762,N_2733);
nor U2807 (N_2807,N_2639,N_2756);
nor U2808 (N_2808,N_2721,N_2611);
nor U2809 (N_2809,N_2712,N_2795);
and U2810 (N_2810,N_2641,N_2637);
and U2811 (N_2811,N_2632,N_2730);
and U2812 (N_2812,N_2612,N_2638);
nor U2813 (N_2813,N_2703,N_2681);
or U2814 (N_2814,N_2680,N_2649);
nor U2815 (N_2815,N_2731,N_2710);
nor U2816 (N_2816,N_2604,N_2758);
or U2817 (N_2817,N_2700,N_2627);
nand U2818 (N_2818,N_2636,N_2744);
nor U2819 (N_2819,N_2622,N_2769);
or U2820 (N_2820,N_2796,N_2662);
nand U2821 (N_2821,N_2655,N_2706);
nor U2822 (N_2822,N_2682,N_2666);
or U2823 (N_2823,N_2647,N_2701);
or U2824 (N_2824,N_2614,N_2619);
nand U2825 (N_2825,N_2657,N_2754);
nand U2826 (N_2826,N_2794,N_2789);
nand U2827 (N_2827,N_2772,N_2739);
nand U2828 (N_2828,N_2601,N_2617);
nand U2829 (N_2829,N_2652,N_2709);
and U2830 (N_2830,N_2751,N_2654);
and U2831 (N_2831,N_2667,N_2623);
nor U2832 (N_2832,N_2644,N_2671);
and U2833 (N_2833,N_2640,N_2745);
nor U2834 (N_2834,N_2678,N_2683);
nand U2835 (N_2835,N_2621,N_2626);
and U2836 (N_2836,N_2741,N_2602);
and U2837 (N_2837,N_2668,N_2699);
nand U2838 (N_2838,N_2784,N_2697);
nand U2839 (N_2839,N_2625,N_2673);
nand U2840 (N_2840,N_2669,N_2757);
or U2841 (N_2841,N_2761,N_2716);
nor U2842 (N_2842,N_2628,N_2743);
nand U2843 (N_2843,N_2735,N_2686);
and U2844 (N_2844,N_2613,N_2750);
nand U2845 (N_2845,N_2675,N_2642);
and U2846 (N_2846,N_2693,N_2771);
or U2847 (N_2847,N_2755,N_2661);
and U2848 (N_2848,N_2663,N_2798);
nor U2849 (N_2849,N_2624,N_2764);
or U2850 (N_2850,N_2692,N_2748);
nor U2851 (N_2851,N_2610,N_2773);
nor U2852 (N_2852,N_2608,N_2620);
nor U2853 (N_2853,N_2783,N_2672);
or U2854 (N_2854,N_2793,N_2770);
and U2855 (N_2855,N_2724,N_2600);
and U2856 (N_2856,N_2607,N_2776);
nor U2857 (N_2857,N_2696,N_2646);
nor U2858 (N_2858,N_2631,N_2629);
and U2859 (N_2859,N_2752,N_2702);
nand U2860 (N_2860,N_2688,N_2695);
and U2861 (N_2861,N_2799,N_2782);
and U2862 (N_2862,N_2634,N_2713);
nor U2863 (N_2863,N_2616,N_2777);
and U2864 (N_2864,N_2650,N_2633);
or U2865 (N_2865,N_2725,N_2722);
nor U2866 (N_2866,N_2690,N_2685);
nor U2867 (N_2867,N_2753,N_2727);
or U2868 (N_2868,N_2645,N_2714);
nand U2869 (N_2869,N_2670,N_2687);
or U2870 (N_2870,N_2774,N_2658);
and U2871 (N_2871,N_2718,N_2781);
nand U2872 (N_2872,N_2715,N_2677);
and U2873 (N_2873,N_2787,N_2653);
nand U2874 (N_2874,N_2792,N_2780);
nand U2875 (N_2875,N_2665,N_2747);
nand U2876 (N_2876,N_2720,N_2785);
nor U2877 (N_2877,N_2778,N_2736);
and U2878 (N_2878,N_2684,N_2606);
or U2879 (N_2879,N_2719,N_2779);
and U2880 (N_2880,N_2603,N_2790);
nand U2881 (N_2881,N_2651,N_2726);
nor U2882 (N_2882,N_2630,N_2746);
and U2883 (N_2883,N_2749,N_2768);
nand U2884 (N_2884,N_2732,N_2664);
or U2885 (N_2885,N_2767,N_2711);
nor U2886 (N_2886,N_2704,N_2734);
nor U2887 (N_2887,N_2659,N_2615);
and U2888 (N_2888,N_2742,N_2689);
or U2889 (N_2889,N_2728,N_2708);
nand U2890 (N_2890,N_2775,N_2707);
and U2891 (N_2891,N_2605,N_2705);
or U2892 (N_2892,N_2609,N_2679);
and U2893 (N_2893,N_2759,N_2676);
nand U2894 (N_2894,N_2717,N_2763);
nand U2895 (N_2895,N_2766,N_2760);
and U2896 (N_2896,N_2765,N_2698);
nor U2897 (N_2897,N_2740,N_2618);
nor U2898 (N_2898,N_2648,N_2660);
nand U2899 (N_2899,N_2786,N_2691);
and U2900 (N_2900,N_2601,N_2731);
or U2901 (N_2901,N_2747,N_2774);
nand U2902 (N_2902,N_2641,N_2695);
nand U2903 (N_2903,N_2755,N_2635);
nor U2904 (N_2904,N_2694,N_2780);
and U2905 (N_2905,N_2628,N_2636);
or U2906 (N_2906,N_2647,N_2619);
and U2907 (N_2907,N_2751,N_2773);
or U2908 (N_2908,N_2693,N_2687);
or U2909 (N_2909,N_2613,N_2728);
or U2910 (N_2910,N_2666,N_2653);
nand U2911 (N_2911,N_2720,N_2674);
nand U2912 (N_2912,N_2728,N_2719);
and U2913 (N_2913,N_2786,N_2789);
nor U2914 (N_2914,N_2642,N_2603);
or U2915 (N_2915,N_2673,N_2725);
or U2916 (N_2916,N_2645,N_2735);
or U2917 (N_2917,N_2673,N_2755);
nand U2918 (N_2918,N_2651,N_2705);
or U2919 (N_2919,N_2745,N_2685);
and U2920 (N_2920,N_2731,N_2692);
nand U2921 (N_2921,N_2684,N_2730);
or U2922 (N_2922,N_2744,N_2784);
nand U2923 (N_2923,N_2746,N_2600);
and U2924 (N_2924,N_2774,N_2759);
or U2925 (N_2925,N_2666,N_2650);
nand U2926 (N_2926,N_2730,N_2626);
nor U2927 (N_2927,N_2728,N_2642);
nor U2928 (N_2928,N_2753,N_2664);
nand U2929 (N_2929,N_2669,N_2749);
nor U2930 (N_2930,N_2694,N_2608);
nor U2931 (N_2931,N_2687,N_2721);
nor U2932 (N_2932,N_2684,N_2788);
nor U2933 (N_2933,N_2645,N_2742);
and U2934 (N_2934,N_2640,N_2648);
or U2935 (N_2935,N_2738,N_2761);
nor U2936 (N_2936,N_2630,N_2706);
nand U2937 (N_2937,N_2773,N_2603);
and U2938 (N_2938,N_2688,N_2749);
and U2939 (N_2939,N_2664,N_2610);
nor U2940 (N_2940,N_2748,N_2653);
or U2941 (N_2941,N_2741,N_2712);
xnor U2942 (N_2942,N_2791,N_2713);
nand U2943 (N_2943,N_2668,N_2618);
nand U2944 (N_2944,N_2753,N_2735);
nor U2945 (N_2945,N_2740,N_2774);
or U2946 (N_2946,N_2641,N_2709);
or U2947 (N_2947,N_2697,N_2760);
xor U2948 (N_2948,N_2766,N_2660);
nor U2949 (N_2949,N_2632,N_2662);
nor U2950 (N_2950,N_2638,N_2652);
or U2951 (N_2951,N_2793,N_2673);
or U2952 (N_2952,N_2764,N_2714);
and U2953 (N_2953,N_2763,N_2732);
and U2954 (N_2954,N_2779,N_2679);
or U2955 (N_2955,N_2767,N_2649);
and U2956 (N_2956,N_2632,N_2626);
nand U2957 (N_2957,N_2785,N_2694);
and U2958 (N_2958,N_2759,N_2738);
nand U2959 (N_2959,N_2749,N_2675);
nand U2960 (N_2960,N_2784,N_2687);
nor U2961 (N_2961,N_2609,N_2671);
and U2962 (N_2962,N_2600,N_2708);
and U2963 (N_2963,N_2676,N_2677);
xnor U2964 (N_2964,N_2760,N_2780);
and U2965 (N_2965,N_2664,N_2668);
nor U2966 (N_2966,N_2761,N_2778);
and U2967 (N_2967,N_2638,N_2776);
nand U2968 (N_2968,N_2783,N_2686);
or U2969 (N_2969,N_2728,N_2786);
or U2970 (N_2970,N_2721,N_2785);
nand U2971 (N_2971,N_2772,N_2715);
nand U2972 (N_2972,N_2610,N_2684);
nor U2973 (N_2973,N_2726,N_2687);
or U2974 (N_2974,N_2608,N_2670);
and U2975 (N_2975,N_2757,N_2650);
nand U2976 (N_2976,N_2684,N_2748);
and U2977 (N_2977,N_2643,N_2737);
nand U2978 (N_2978,N_2702,N_2732);
nor U2979 (N_2979,N_2772,N_2796);
and U2980 (N_2980,N_2719,N_2613);
or U2981 (N_2981,N_2639,N_2728);
nor U2982 (N_2982,N_2754,N_2715);
or U2983 (N_2983,N_2635,N_2793);
nand U2984 (N_2984,N_2661,N_2751);
and U2985 (N_2985,N_2717,N_2751);
nor U2986 (N_2986,N_2745,N_2773);
nand U2987 (N_2987,N_2687,N_2616);
nor U2988 (N_2988,N_2792,N_2730);
or U2989 (N_2989,N_2672,N_2787);
nand U2990 (N_2990,N_2622,N_2630);
and U2991 (N_2991,N_2739,N_2619);
and U2992 (N_2992,N_2785,N_2606);
nand U2993 (N_2993,N_2662,N_2628);
nand U2994 (N_2994,N_2640,N_2604);
nor U2995 (N_2995,N_2670,N_2643);
nand U2996 (N_2996,N_2717,N_2757);
or U2997 (N_2997,N_2600,N_2659);
and U2998 (N_2998,N_2611,N_2743);
and U2999 (N_2999,N_2641,N_2728);
or UO_0 (O_0,N_2819,N_2863);
nor UO_1 (O_1,N_2992,N_2952);
nor UO_2 (O_2,N_2960,N_2826);
nor UO_3 (O_3,N_2931,N_2953);
nand UO_4 (O_4,N_2964,N_2875);
and UO_5 (O_5,N_2905,N_2965);
xor UO_6 (O_6,N_2856,N_2828);
nor UO_7 (O_7,N_2838,N_2911);
nand UO_8 (O_8,N_2831,N_2842);
nand UO_9 (O_9,N_2805,N_2809);
nor UO_10 (O_10,N_2873,N_2942);
and UO_11 (O_11,N_2937,N_2966);
nand UO_12 (O_12,N_2973,N_2804);
nor UO_13 (O_13,N_2907,N_2812);
nand UO_14 (O_14,N_2957,N_2853);
nand UO_15 (O_15,N_2827,N_2886);
and UO_16 (O_16,N_2896,N_2803);
nor UO_17 (O_17,N_2921,N_2975);
nand UO_18 (O_18,N_2903,N_2970);
or UO_19 (O_19,N_2870,N_2800);
nor UO_20 (O_20,N_2949,N_2845);
nand UO_21 (O_21,N_2833,N_2945);
and UO_22 (O_22,N_2976,N_2859);
and UO_23 (O_23,N_2988,N_2948);
nand UO_24 (O_24,N_2815,N_2802);
nor UO_25 (O_25,N_2829,N_2925);
nor UO_26 (O_26,N_2995,N_2862);
nor UO_27 (O_27,N_2820,N_2874);
and UO_28 (O_28,N_2987,N_2861);
nand UO_29 (O_29,N_2824,N_2951);
or UO_30 (O_30,N_2985,N_2923);
or UO_31 (O_31,N_2898,N_2916);
and UO_32 (O_32,N_2865,N_2927);
or UO_33 (O_33,N_2940,N_2852);
and UO_34 (O_34,N_2872,N_2825);
nand UO_35 (O_35,N_2847,N_2986);
nand UO_36 (O_36,N_2946,N_2933);
and UO_37 (O_37,N_2991,N_2947);
and UO_38 (O_38,N_2854,N_2971);
or UO_39 (O_39,N_2883,N_2881);
or UO_40 (O_40,N_2936,N_2901);
or UO_41 (O_41,N_2899,N_2908);
and UO_42 (O_42,N_2906,N_2962);
nor UO_43 (O_43,N_2846,N_2918);
nand UO_44 (O_44,N_2938,N_2851);
or UO_45 (O_45,N_2902,N_2989);
and UO_46 (O_46,N_2910,N_2849);
and UO_47 (O_47,N_2891,N_2996);
and UO_48 (O_48,N_2994,N_2928);
nand UO_49 (O_49,N_2926,N_2884);
nand UO_50 (O_50,N_2968,N_2888);
nand UO_51 (O_51,N_2832,N_2839);
and UO_52 (O_52,N_2848,N_2864);
or UO_53 (O_53,N_2808,N_2879);
or UO_54 (O_54,N_2932,N_2956);
nand UO_55 (O_55,N_2924,N_2816);
or UO_56 (O_56,N_2857,N_2941);
nor UO_57 (O_57,N_2979,N_2963);
and UO_58 (O_58,N_2944,N_2929);
and UO_59 (O_59,N_2990,N_2977);
or UO_60 (O_60,N_2961,N_2871);
nand UO_61 (O_61,N_2893,N_2959);
and UO_62 (O_62,N_2840,N_2913);
nand UO_63 (O_63,N_2972,N_2998);
nand UO_64 (O_64,N_2984,N_2867);
nor UO_65 (O_65,N_2860,N_2887);
nor UO_66 (O_66,N_2890,N_2837);
or UO_67 (O_67,N_2813,N_2878);
or UO_68 (O_68,N_2997,N_2978);
nand UO_69 (O_69,N_2895,N_2980);
and UO_70 (O_70,N_2894,N_2868);
and UO_71 (O_71,N_2909,N_2955);
and UO_72 (O_72,N_2914,N_2877);
nand UO_73 (O_73,N_2993,N_2814);
nand UO_74 (O_74,N_2930,N_2811);
nor UO_75 (O_75,N_2869,N_2850);
or UO_76 (O_76,N_2843,N_2919);
nor UO_77 (O_77,N_2912,N_2967);
xor UO_78 (O_78,N_2915,N_2834);
nand UO_79 (O_79,N_2835,N_2920);
or UO_80 (O_80,N_2900,N_2969);
or UO_81 (O_81,N_2841,N_2807);
nand UO_82 (O_82,N_2922,N_2999);
nor UO_83 (O_83,N_2935,N_2880);
and UO_84 (O_84,N_2904,N_2950);
nand UO_85 (O_85,N_2981,N_2958);
or UO_86 (O_86,N_2982,N_2806);
or UO_87 (O_87,N_2844,N_2876);
nand UO_88 (O_88,N_2983,N_2823);
and UO_89 (O_89,N_2810,N_2954);
nand UO_90 (O_90,N_2866,N_2974);
nor UO_91 (O_91,N_2897,N_2917);
nand UO_92 (O_92,N_2822,N_2882);
xor UO_93 (O_93,N_2889,N_2836);
nor UO_94 (O_94,N_2934,N_2818);
nor UO_95 (O_95,N_2892,N_2939);
or UO_96 (O_96,N_2801,N_2858);
or UO_97 (O_97,N_2830,N_2855);
nand UO_98 (O_98,N_2821,N_2943);
nor UO_99 (O_99,N_2817,N_2885);
and UO_100 (O_100,N_2895,N_2871);
and UO_101 (O_101,N_2861,N_2864);
and UO_102 (O_102,N_2937,N_2839);
and UO_103 (O_103,N_2968,N_2856);
or UO_104 (O_104,N_2885,N_2898);
nand UO_105 (O_105,N_2952,N_2985);
nand UO_106 (O_106,N_2838,N_2855);
nand UO_107 (O_107,N_2932,N_2948);
nor UO_108 (O_108,N_2994,N_2833);
or UO_109 (O_109,N_2995,N_2954);
or UO_110 (O_110,N_2921,N_2944);
nor UO_111 (O_111,N_2818,N_2903);
nor UO_112 (O_112,N_2846,N_2972);
or UO_113 (O_113,N_2818,N_2909);
nand UO_114 (O_114,N_2834,N_2870);
nand UO_115 (O_115,N_2950,N_2996);
nand UO_116 (O_116,N_2874,N_2816);
xor UO_117 (O_117,N_2903,N_2817);
xor UO_118 (O_118,N_2993,N_2805);
xor UO_119 (O_119,N_2944,N_2836);
nor UO_120 (O_120,N_2929,N_2857);
and UO_121 (O_121,N_2840,N_2891);
and UO_122 (O_122,N_2958,N_2897);
nor UO_123 (O_123,N_2922,N_2962);
xor UO_124 (O_124,N_2945,N_2849);
and UO_125 (O_125,N_2978,N_2972);
nand UO_126 (O_126,N_2908,N_2997);
nor UO_127 (O_127,N_2985,N_2801);
nand UO_128 (O_128,N_2875,N_2879);
nor UO_129 (O_129,N_2896,N_2989);
nand UO_130 (O_130,N_2851,N_2995);
nor UO_131 (O_131,N_2913,N_2827);
nor UO_132 (O_132,N_2840,N_2969);
or UO_133 (O_133,N_2831,N_2895);
nand UO_134 (O_134,N_2965,N_2934);
nor UO_135 (O_135,N_2996,N_2874);
nand UO_136 (O_136,N_2932,N_2920);
and UO_137 (O_137,N_2958,N_2973);
and UO_138 (O_138,N_2863,N_2867);
nand UO_139 (O_139,N_2933,N_2967);
and UO_140 (O_140,N_2802,N_2862);
nand UO_141 (O_141,N_2842,N_2890);
nand UO_142 (O_142,N_2884,N_2807);
nand UO_143 (O_143,N_2901,N_2808);
nor UO_144 (O_144,N_2864,N_2856);
or UO_145 (O_145,N_2860,N_2939);
nand UO_146 (O_146,N_2819,N_2938);
nand UO_147 (O_147,N_2840,N_2855);
nor UO_148 (O_148,N_2827,N_2973);
or UO_149 (O_149,N_2919,N_2953);
and UO_150 (O_150,N_2987,N_2937);
nor UO_151 (O_151,N_2883,N_2816);
or UO_152 (O_152,N_2994,N_2888);
nand UO_153 (O_153,N_2924,N_2905);
nor UO_154 (O_154,N_2864,N_2915);
nand UO_155 (O_155,N_2876,N_2959);
and UO_156 (O_156,N_2935,N_2896);
nand UO_157 (O_157,N_2959,N_2909);
and UO_158 (O_158,N_2893,N_2865);
or UO_159 (O_159,N_2845,N_2885);
and UO_160 (O_160,N_2955,N_2912);
nand UO_161 (O_161,N_2858,N_2895);
xnor UO_162 (O_162,N_2998,N_2919);
nor UO_163 (O_163,N_2942,N_2841);
nand UO_164 (O_164,N_2865,N_2978);
and UO_165 (O_165,N_2919,N_2993);
or UO_166 (O_166,N_2812,N_2893);
nor UO_167 (O_167,N_2954,N_2937);
or UO_168 (O_168,N_2812,N_2947);
and UO_169 (O_169,N_2821,N_2946);
nand UO_170 (O_170,N_2940,N_2926);
or UO_171 (O_171,N_2806,N_2978);
nand UO_172 (O_172,N_2985,N_2838);
and UO_173 (O_173,N_2818,N_2949);
or UO_174 (O_174,N_2802,N_2942);
and UO_175 (O_175,N_2962,N_2878);
or UO_176 (O_176,N_2895,N_2884);
nand UO_177 (O_177,N_2900,N_2935);
nor UO_178 (O_178,N_2916,N_2996);
and UO_179 (O_179,N_2824,N_2920);
nand UO_180 (O_180,N_2824,N_2936);
nor UO_181 (O_181,N_2909,N_2802);
and UO_182 (O_182,N_2911,N_2897);
or UO_183 (O_183,N_2802,N_2812);
or UO_184 (O_184,N_2899,N_2832);
and UO_185 (O_185,N_2993,N_2912);
nor UO_186 (O_186,N_2841,N_2957);
or UO_187 (O_187,N_2956,N_2987);
nand UO_188 (O_188,N_2975,N_2861);
nor UO_189 (O_189,N_2981,N_2947);
nand UO_190 (O_190,N_2939,N_2834);
and UO_191 (O_191,N_2933,N_2969);
or UO_192 (O_192,N_2971,N_2924);
nor UO_193 (O_193,N_2915,N_2839);
or UO_194 (O_194,N_2879,N_2983);
or UO_195 (O_195,N_2885,N_2965);
and UO_196 (O_196,N_2872,N_2807);
nand UO_197 (O_197,N_2985,N_2982);
nand UO_198 (O_198,N_2807,N_2811);
nor UO_199 (O_199,N_2837,N_2870);
or UO_200 (O_200,N_2924,N_2931);
nand UO_201 (O_201,N_2853,N_2864);
nand UO_202 (O_202,N_2808,N_2863);
or UO_203 (O_203,N_2822,N_2937);
nor UO_204 (O_204,N_2864,N_2903);
nor UO_205 (O_205,N_2912,N_2825);
nor UO_206 (O_206,N_2899,N_2944);
nand UO_207 (O_207,N_2804,N_2953);
and UO_208 (O_208,N_2852,N_2981);
nand UO_209 (O_209,N_2936,N_2981);
and UO_210 (O_210,N_2801,N_2944);
nor UO_211 (O_211,N_2840,N_2924);
or UO_212 (O_212,N_2886,N_2892);
or UO_213 (O_213,N_2971,N_2925);
or UO_214 (O_214,N_2807,N_2808);
and UO_215 (O_215,N_2906,N_2822);
nand UO_216 (O_216,N_2924,N_2866);
and UO_217 (O_217,N_2969,N_2817);
nand UO_218 (O_218,N_2837,N_2915);
and UO_219 (O_219,N_2977,N_2800);
nor UO_220 (O_220,N_2957,N_2804);
or UO_221 (O_221,N_2850,N_2876);
nand UO_222 (O_222,N_2882,N_2940);
or UO_223 (O_223,N_2960,N_2864);
nor UO_224 (O_224,N_2908,N_2991);
or UO_225 (O_225,N_2947,N_2910);
nor UO_226 (O_226,N_2843,N_2995);
or UO_227 (O_227,N_2892,N_2958);
nor UO_228 (O_228,N_2898,N_2997);
and UO_229 (O_229,N_2896,N_2850);
nor UO_230 (O_230,N_2898,N_2850);
nor UO_231 (O_231,N_2814,N_2954);
or UO_232 (O_232,N_2829,N_2966);
nand UO_233 (O_233,N_2961,N_2962);
or UO_234 (O_234,N_2908,N_2981);
nor UO_235 (O_235,N_2942,N_2909);
nand UO_236 (O_236,N_2811,N_2800);
and UO_237 (O_237,N_2919,N_2915);
nand UO_238 (O_238,N_2800,N_2813);
and UO_239 (O_239,N_2878,N_2944);
nor UO_240 (O_240,N_2870,N_2881);
nand UO_241 (O_241,N_2816,N_2827);
or UO_242 (O_242,N_2833,N_2822);
nand UO_243 (O_243,N_2809,N_2993);
nor UO_244 (O_244,N_2817,N_2861);
and UO_245 (O_245,N_2905,N_2993);
nor UO_246 (O_246,N_2941,N_2984);
nand UO_247 (O_247,N_2901,N_2854);
or UO_248 (O_248,N_2993,N_2885);
and UO_249 (O_249,N_2918,N_2970);
nor UO_250 (O_250,N_2911,N_2830);
nor UO_251 (O_251,N_2857,N_2850);
nand UO_252 (O_252,N_2838,N_2876);
or UO_253 (O_253,N_2986,N_2861);
nand UO_254 (O_254,N_2849,N_2807);
and UO_255 (O_255,N_2822,N_2919);
and UO_256 (O_256,N_2924,N_2955);
and UO_257 (O_257,N_2944,N_2879);
nor UO_258 (O_258,N_2973,N_2862);
or UO_259 (O_259,N_2988,N_2981);
and UO_260 (O_260,N_2890,N_2834);
and UO_261 (O_261,N_2871,N_2805);
nor UO_262 (O_262,N_2830,N_2938);
nand UO_263 (O_263,N_2890,N_2866);
and UO_264 (O_264,N_2948,N_2877);
or UO_265 (O_265,N_2986,N_2964);
or UO_266 (O_266,N_2987,N_2914);
and UO_267 (O_267,N_2915,N_2926);
nor UO_268 (O_268,N_2972,N_2953);
nand UO_269 (O_269,N_2921,N_2822);
or UO_270 (O_270,N_2951,N_2975);
and UO_271 (O_271,N_2895,N_2934);
nand UO_272 (O_272,N_2954,N_2970);
nand UO_273 (O_273,N_2919,N_2965);
or UO_274 (O_274,N_2804,N_2910);
or UO_275 (O_275,N_2887,N_2912);
or UO_276 (O_276,N_2887,N_2899);
nor UO_277 (O_277,N_2849,N_2986);
nand UO_278 (O_278,N_2970,N_2851);
nor UO_279 (O_279,N_2801,N_2826);
nand UO_280 (O_280,N_2822,N_2915);
or UO_281 (O_281,N_2812,N_2999);
nand UO_282 (O_282,N_2874,N_2863);
nor UO_283 (O_283,N_2841,N_2998);
and UO_284 (O_284,N_2809,N_2959);
nor UO_285 (O_285,N_2941,N_2928);
and UO_286 (O_286,N_2886,N_2834);
and UO_287 (O_287,N_2846,N_2911);
and UO_288 (O_288,N_2916,N_2958);
or UO_289 (O_289,N_2954,N_2906);
and UO_290 (O_290,N_2908,N_2961);
nor UO_291 (O_291,N_2879,N_2896);
nor UO_292 (O_292,N_2823,N_2889);
or UO_293 (O_293,N_2915,N_2930);
and UO_294 (O_294,N_2875,N_2839);
nor UO_295 (O_295,N_2970,N_2883);
and UO_296 (O_296,N_2926,N_2876);
nand UO_297 (O_297,N_2880,N_2980);
and UO_298 (O_298,N_2987,N_2959);
nor UO_299 (O_299,N_2986,N_2832);
and UO_300 (O_300,N_2921,N_2978);
nand UO_301 (O_301,N_2885,N_2861);
nor UO_302 (O_302,N_2930,N_2974);
or UO_303 (O_303,N_2862,N_2998);
nand UO_304 (O_304,N_2938,N_2842);
nor UO_305 (O_305,N_2901,N_2956);
nand UO_306 (O_306,N_2909,N_2866);
or UO_307 (O_307,N_2814,N_2803);
or UO_308 (O_308,N_2812,N_2935);
nand UO_309 (O_309,N_2922,N_2899);
nor UO_310 (O_310,N_2809,N_2861);
or UO_311 (O_311,N_2818,N_2854);
nand UO_312 (O_312,N_2970,N_2941);
nor UO_313 (O_313,N_2988,N_2853);
and UO_314 (O_314,N_2930,N_2964);
and UO_315 (O_315,N_2850,N_2853);
nand UO_316 (O_316,N_2865,N_2841);
and UO_317 (O_317,N_2854,N_2842);
or UO_318 (O_318,N_2845,N_2972);
nand UO_319 (O_319,N_2903,N_2895);
nor UO_320 (O_320,N_2919,N_2884);
or UO_321 (O_321,N_2808,N_2868);
nand UO_322 (O_322,N_2997,N_2809);
nor UO_323 (O_323,N_2994,N_2962);
or UO_324 (O_324,N_2843,N_2965);
nand UO_325 (O_325,N_2894,N_2920);
or UO_326 (O_326,N_2870,N_2806);
xnor UO_327 (O_327,N_2977,N_2991);
nor UO_328 (O_328,N_2906,N_2806);
nor UO_329 (O_329,N_2873,N_2846);
nand UO_330 (O_330,N_2926,N_2923);
and UO_331 (O_331,N_2897,N_2940);
nand UO_332 (O_332,N_2949,N_2946);
nor UO_333 (O_333,N_2903,N_2925);
and UO_334 (O_334,N_2834,N_2860);
or UO_335 (O_335,N_2999,N_2818);
or UO_336 (O_336,N_2955,N_2974);
and UO_337 (O_337,N_2873,N_2991);
nand UO_338 (O_338,N_2977,N_2983);
xnor UO_339 (O_339,N_2887,N_2995);
and UO_340 (O_340,N_2812,N_2958);
nand UO_341 (O_341,N_2942,N_2971);
or UO_342 (O_342,N_2940,N_2876);
or UO_343 (O_343,N_2901,N_2836);
or UO_344 (O_344,N_2908,N_2802);
nand UO_345 (O_345,N_2967,N_2821);
nor UO_346 (O_346,N_2801,N_2848);
nor UO_347 (O_347,N_2994,N_2958);
nand UO_348 (O_348,N_2931,N_2842);
nor UO_349 (O_349,N_2958,N_2870);
nor UO_350 (O_350,N_2837,N_2936);
and UO_351 (O_351,N_2996,N_2832);
and UO_352 (O_352,N_2873,N_2996);
and UO_353 (O_353,N_2871,N_2969);
nand UO_354 (O_354,N_2996,N_2904);
xor UO_355 (O_355,N_2835,N_2990);
nor UO_356 (O_356,N_2895,N_2839);
nand UO_357 (O_357,N_2998,N_2963);
and UO_358 (O_358,N_2945,N_2813);
nand UO_359 (O_359,N_2858,N_2985);
or UO_360 (O_360,N_2831,N_2852);
nor UO_361 (O_361,N_2956,N_2954);
and UO_362 (O_362,N_2806,N_2926);
nor UO_363 (O_363,N_2816,N_2835);
or UO_364 (O_364,N_2820,N_2860);
or UO_365 (O_365,N_2840,N_2895);
and UO_366 (O_366,N_2990,N_2800);
nor UO_367 (O_367,N_2844,N_2911);
and UO_368 (O_368,N_2977,N_2949);
or UO_369 (O_369,N_2815,N_2939);
and UO_370 (O_370,N_2931,N_2811);
and UO_371 (O_371,N_2824,N_2848);
nand UO_372 (O_372,N_2989,N_2906);
nand UO_373 (O_373,N_2808,N_2899);
xnor UO_374 (O_374,N_2969,N_2957);
nor UO_375 (O_375,N_2899,N_2942);
nand UO_376 (O_376,N_2971,N_2866);
nand UO_377 (O_377,N_2900,N_2984);
and UO_378 (O_378,N_2884,N_2898);
nand UO_379 (O_379,N_2900,N_2861);
nor UO_380 (O_380,N_2953,N_2868);
nand UO_381 (O_381,N_2902,N_2848);
or UO_382 (O_382,N_2857,N_2930);
or UO_383 (O_383,N_2982,N_2877);
nor UO_384 (O_384,N_2931,N_2823);
and UO_385 (O_385,N_2935,N_2878);
nand UO_386 (O_386,N_2935,N_2872);
and UO_387 (O_387,N_2835,N_2900);
or UO_388 (O_388,N_2959,N_2850);
or UO_389 (O_389,N_2853,N_2887);
and UO_390 (O_390,N_2896,N_2991);
nand UO_391 (O_391,N_2842,N_2889);
xor UO_392 (O_392,N_2963,N_2916);
nand UO_393 (O_393,N_2959,N_2954);
nand UO_394 (O_394,N_2926,N_2828);
or UO_395 (O_395,N_2816,N_2955);
or UO_396 (O_396,N_2875,N_2972);
or UO_397 (O_397,N_2964,N_2948);
and UO_398 (O_398,N_2808,N_2882);
nand UO_399 (O_399,N_2871,N_2811);
nand UO_400 (O_400,N_2838,N_2965);
nand UO_401 (O_401,N_2883,N_2885);
and UO_402 (O_402,N_2939,N_2913);
nand UO_403 (O_403,N_2858,N_2842);
nand UO_404 (O_404,N_2894,N_2927);
nand UO_405 (O_405,N_2843,N_2842);
and UO_406 (O_406,N_2886,N_2857);
nand UO_407 (O_407,N_2810,N_2946);
xnor UO_408 (O_408,N_2848,N_2869);
or UO_409 (O_409,N_2999,N_2871);
or UO_410 (O_410,N_2957,N_2830);
or UO_411 (O_411,N_2945,N_2994);
nand UO_412 (O_412,N_2831,N_2875);
or UO_413 (O_413,N_2863,N_2878);
and UO_414 (O_414,N_2990,N_2991);
or UO_415 (O_415,N_2867,N_2871);
or UO_416 (O_416,N_2974,N_2978);
nand UO_417 (O_417,N_2956,N_2831);
nand UO_418 (O_418,N_2904,N_2886);
nand UO_419 (O_419,N_2951,N_2879);
or UO_420 (O_420,N_2956,N_2883);
and UO_421 (O_421,N_2829,N_2864);
nand UO_422 (O_422,N_2954,N_2922);
and UO_423 (O_423,N_2829,N_2852);
nand UO_424 (O_424,N_2934,N_2821);
nor UO_425 (O_425,N_2915,N_2878);
or UO_426 (O_426,N_2805,N_2925);
or UO_427 (O_427,N_2845,N_2876);
nor UO_428 (O_428,N_2980,N_2864);
xor UO_429 (O_429,N_2988,N_2915);
nor UO_430 (O_430,N_2905,N_2830);
and UO_431 (O_431,N_2810,N_2843);
and UO_432 (O_432,N_2874,N_2802);
or UO_433 (O_433,N_2883,N_2859);
nand UO_434 (O_434,N_2811,N_2806);
nand UO_435 (O_435,N_2880,N_2962);
and UO_436 (O_436,N_2957,N_2839);
or UO_437 (O_437,N_2858,N_2964);
and UO_438 (O_438,N_2951,N_2977);
nor UO_439 (O_439,N_2816,N_2838);
and UO_440 (O_440,N_2976,N_2942);
or UO_441 (O_441,N_2811,N_2865);
nor UO_442 (O_442,N_2844,N_2902);
nand UO_443 (O_443,N_2946,N_2897);
nor UO_444 (O_444,N_2979,N_2937);
nand UO_445 (O_445,N_2977,N_2900);
nand UO_446 (O_446,N_2879,N_2963);
nand UO_447 (O_447,N_2994,N_2826);
and UO_448 (O_448,N_2914,N_2802);
nor UO_449 (O_449,N_2924,N_2952);
nor UO_450 (O_450,N_2992,N_2927);
or UO_451 (O_451,N_2854,N_2815);
and UO_452 (O_452,N_2831,N_2945);
nand UO_453 (O_453,N_2972,N_2876);
nand UO_454 (O_454,N_2855,N_2876);
or UO_455 (O_455,N_2819,N_2934);
and UO_456 (O_456,N_2942,N_2996);
nor UO_457 (O_457,N_2868,N_2943);
and UO_458 (O_458,N_2891,N_2977);
or UO_459 (O_459,N_2979,N_2878);
nor UO_460 (O_460,N_2945,N_2943);
nand UO_461 (O_461,N_2922,N_2996);
or UO_462 (O_462,N_2970,N_2840);
xor UO_463 (O_463,N_2802,N_2863);
or UO_464 (O_464,N_2991,N_2937);
nand UO_465 (O_465,N_2851,N_2824);
nand UO_466 (O_466,N_2880,N_2925);
or UO_467 (O_467,N_2826,N_2930);
nor UO_468 (O_468,N_2840,N_2993);
nor UO_469 (O_469,N_2831,N_2811);
nand UO_470 (O_470,N_2854,N_2988);
xor UO_471 (O_471,N_2939,N_2905);
nor UO_472 (O_472,N_2897,N_2995);
nor UO_473 (O_473,N_2952,N_2886);
xor UO_474 (O_474,N_2845,N_2825);
and UO_475 (O_475,N_2925,N_2800);
nor UO_476 (O_476,N_2929,N_2828);
and UO_477 (O_477,N_2840,N_2896);
or UO_478 (O_478,N_2838,N_2852);
and UO_479 (O_479,N_2964,N_2936);
nand UO_480 (O_480,N_2950,N_2833);
and UO_481 (O_481,N_2885,N_2826);
and UO_482 (O_482,N_2999,N_2994);
nand UO_483 (O_483,N_2868,N_2992);
nand UO_484 (O_484,N_2973,N_2981);
and UO_485 (O_485,N_2937,N_2861);
nor UO_486 (O_486,N_2872,N_2963);
or UO_487 (O_487,N_2894,N_2903);
or UO_488 (O_488,N_2911,N_2975);
nand UO_489 (O_489,N_2904,N_2971);
nand UO_490 (O_490,N_2925,N_2858);
or UO_491 (O_491,N_2976,N_2930);
and UO_492 (O_492,N_2821,N_2887);
or UO_493 (O_493,N_2964,N_2859);
xnor UO_494 (O_494,N_2983,N_2979);
nor UO_495 (O_495,N_2814,N_2994);
nand UO_496 (O_496,N_2935,N_2858);
or UO_497 (O_497,N_2823,N_2809);
nand UO_498 (O_498,N_2916,N_2856);
and UO_499 (O_499,N_2978,N_2990);
endmodule