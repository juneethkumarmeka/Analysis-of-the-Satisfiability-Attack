module basic_500_3000_500_6_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_487,In_170);
and U1 (N_1,In_469,In_267);
xnor U2 (N_2,In_251,In_129);
nor U3 (N_3,In_188,In_50);
nor U4 (N_4,In_136,In_325);
nand U5 (N_5,In_412,In_371);
and U6 (N_6,In_342,In_233);
and U7 (N_7,In_157,In_235);
or U8 (N_8,In_187,In_213);
nor U9 (N_9,In_4,In_231);
or U10 (N_10,In_185,In_149);
nand U11 (N_11,In_112,In_8);
nor U12 (N_12,In_35,In_194);
nand U13 (N_13,In_485,In_102);
nor U14 (N_14,In_491,In_181);
nand U15 (N_15,In_172,In_314);
nor U16 (N_16,In_430,In_227);
and U17 (N_17,In_166,In_139);
nor U18 (N_18,In_254,In_228);
and U19 (N_19,In_328,In_164);
or U20 (N_20,In_162,In_404);
and U21 (N_21,In_106,In_341);
nand U22 (N_22,In_137,In_305);
nand U23 (N_23,In_120,In_224);
nor U24 (N_24,In_17,In_429);
nor U25 (N_25,In_355,In_475);
nor U26 (N_26,In_408,In_62);
nand U27 (N_27,In_0,In_439);
xor U28 (N_28,In_466,In_258);
nand U29 (N_29,In_427,In_163);
nand U30 (N_30,In_452,In_74);
or U31 (N_31,In_222,In_138);
nor U32 (N_32,In_454,In_192);
and U33 (N_33,In_87,In_193);
nand U34 (N_34,In_144,In_257);
nor U35 (N_35,In_195,In_447);
or U36 (N_36,In_101,In_202);
nor U37 (N_37,In_354,In_126);
nand U38 (N_38,In_240,In_303);
nor U39 (N_39,In_19,In_384);
nor U40 (N_40,In_71,In_321);
and U41 (N_41,In_434,In_309);
nor U42 (N_42,In_183,In_155);
and U43 (N_43,In_242,In_255);
nor U44 (N_44,In_85,In_208);
nor U45 (N_45,In_64,In_322);
nor U46 (N_46,In_395,In_245);
and U47 (N_47,In_159,In_400);
nor U48 (N_48,In_189,In_36);
and U49 (N_49,In_394,In_61);
nand U50 (N_50,In_333,In_88);
and U51 (N_51,In_244,In_282);
or U52 (N_52,In_30,In_331);
or U53 (N_53,In_474,In_131);
nand U54 (N_54,In_16,In_368);
nand U55 (N_55,In_463,In_94);
nand U56 (N_56,In_57,In_358);
nor U57 (N_57,In_356,In_277);
nor U58 (N_58,In_75,In_145);
and U59 (N_59,In_81,In_334);
nand U60 (N_60,In_495,In_34);
nor U61 (N_61,In_301,In_169);
nand U62 (N_62,In_241,In_291);
or U63 (N_63,In_117,In_51);
nand U64 (N_64,In_272,In_426);
and U65 (N_65,In_410,In_416);
nor U66 (N_66,In_478,In_488);
or U67 (N_67,In_56,In_46);
or U68 (N_68,In_347,In_498);
nand U69 (N_69,In_393,In_72);
nor U70 (N_70,In_397,In_68);
and U71 (N_71,In_42,In_310);
nor U72 (N_72,In_338,In_23);
nor U73 (N_73,In_362,In_247);
and U74 (N_74,In_148,In_26);
nor U75 (N_75,In_292,In_13);
and U76 (N_76,In_197,In_493);
and U77 (N_77,In_66,In_494);
nor U78 (N_78,In_378,In_216);
nor U79 (N_79,In_108,In_374);
nor U80 (N_80,In_382,In_361);
nand U81 (N_81,In_203,In_421);
nand U82 (N_82,In_38,In_201);
or U83 (N_83,In_73,In_265);
and U84 (N_84,In_154,In_204);
and U85 (N_85,In_48,In_6);
or U86 (N_86,In_340,In_43);
and U87 (N_87,In_103,In_180);
and U88 (N_88,In_389,In_306);
nor U89 (N_89,In_248,In_442);
or U90 (N_90,In_173,In_433);
or U91 (N_91,In_296,In_229);
nor U92 (N_92,In_337,In_21);
or U93 (N_93,In_379,In_302);
nand U94 (N_94,In_445,In_58);
and U95 (N_95,In_67,In_11);
nor U96 (N_96,In_390,In_97);
nand U97 (N_97,In_210,In_191);
nand U98 (N_98,In_111,In_119);
or U99 (N_99,In_349,In_448);
nor U100 (N_100,In_456,In_419);
nand U101 (N_101,In_327,In_330);
nand U102 (N_102,In_152,In_25);
nor U103 (N_103,In_28,In_323);
nand U104 (N_104,In_453,In_190);
and U105 (N_105,In_299,In_158);
xnor U106 (N_106,In_178,In_490);
nor U107 (N_107,In_176,In_405);
and U108 (N_108,In_375,In_264);
and U109 (N_109,In_161,In_403);
or U110 (N_110,In_125,In_196);
and U111 (N_111,In_44,In_122);
nand U112 (N_112,In_449,In_450);
and U113 (N_113,In_268,In_344);
or U114 (N_114,In_319,In_286);
or U115 (N_115,In_263,In_7);
nand U116 (N_116,In_84,In_399);
nor U117 (N_117,In_407,In_440);
xor U118 (N_118,In_116,In_134);
xnor U119 (N_119,In_83,In_33);
or U120 (N_120,In_150,In_486);
nand U121 (N_121,In_441,In_182);
or U122 (N_122,In_114,In_60);
or U123 (N_123,In_65,In_300);
or U124 (N_124,In_460,In_372);
nand U125 (N_125,In_431,In_285);
nor U126 (N_126,In_143,In_91);
nor U127 (N_127,In_212,In_18);
and U128 (N_128,In_262,In_270);
nand U129 (N_129,In_467,In_275);
nor U130 (N_130,In_232,In_100);
nor U131 (N_131,In_381,In_364);
nor U132 (N_132,In_443,In_414);
nand U133 (N_133,In_348,In_96);
nand U134 (N_134,In_9,In_496);
or U135 (N_135,In_470,In_432);
nor U136 (N_136,In_271,In_250);
xor U137 (N_137,In_420,In_468);
and U138 (N_138,In_489,In_332);
nand U139 (N_139,In_477,In_385);
nand U140 (N_140,In_175,In_121);
and U141 (N_141,In_278,In_76);
nand U142 (N_142,In_479,In_200);
nor U143 (N_143,In_160,In_47);
and U144 (N_144,In_401,In_79);
xnor U145 (N_145,In_206,In_53);
or U146 (N_146,In_417,In_77);
nand U147 (N_147,In_353,In_37);
nand U148 (N_148,In_295,In_41);
nand U149 (N_149,In_174,In_132);
nor U150 (N_150,In_3,In_24);
or U151 (N_151,In_165,In_380);
nand U152 (N_152,In_218,In_482);
nor U153 (N_153,In_398,In_20);
and U154 (N_154,In_289,In_446);
xor U155 (N_155,In_459,In_225);
and U156 (N_156,In_437,In_499);
nor U157 (N_157,In_230,In_80);
nand U158 (N_158,In_392,In_223);
or U159 (N_159,In_104,In_352);
or U160 (N_160,In_373,In_465);
xor U161 (N_161,In_326,In_133);
or U162 (N_162,In_12,In_436);
and U163 (N_163,In_177,In_483);
and U164 (N_164,In_52,In_179);
nor U165 (N_165,In_367,In_78);
nand U166 (N_166,In_415,In_238);
or U167 (N_167,In_365,In_127);
nor U168 (N_168,In_461,In_184);
and U169 (N_169,In_281,In_142);
and U170 (N_170,In_313,In_10);
and U171 (N_171,In_307,In_146);
and U172 (N_172,In_135,In_350);
and U173 (N_173,In_249,In_351);
or U174 (N_174,In_59,In_473);
nand U175 (N_175,In_5,In_215);
and U176 (N_176,In_444,In_492);
nand U177 (N_177,In_336,In_92);
and U178 (N_178,In_359,In_1);
and U179 (N_179,In_284,In_205);
nor U180 (N_180,In_413,In_113);
and U181 (N_181,In_424,In_370);
or U182 (N_182,In_409,In_311);
nand U183 (N_183,In_115,In_236);
and U184 (N_184,In_324,In_411);
nor U185 (N_185,In_304,In_217);
nor U186 (N_186,In_207,In_318);
and U187 (N_187,In_105,In_288);
or U188 (N_188,In_383,In_476);
nand U189 (N_189,In_198,In_219);
and U190 (N_190,In_226,In_458);
and U191 (N_191,In_298,In_388);
and U192 (N_192,In_256,In_45);
xnor U193 (N_193,In_260,In_99);
nand U194 (N_194,In_220,In_14);
xor U195 (N_195,In_422,In_329);
and U196 (N_196,In_369,In_156);
nand U197 (N_197,In_15,In_276);
or U198 (N_198,In_147,In_98);
or U199 (N_199,In_472,In_107);
or U200 (N_200,In_199,In_123);
or U201 (N_201,In_435,In_40);
nand U202 (N_202,In_481,In_343);
nand U203 (N_203,In_402,In_54);
or U204 (N_204,In_243,In_308);
and U205 (N_205,In_428,In_280);
or U206 (N_206,In_234,In_49);
and U207 (N_207,In_287,In_391);
nor U208 (N_208,In_438,In_363);
and U209 (N_209,In_386,In_462);
and U210 (N_210,In_118,In_283);
or U211 (N_211,In_451,In_464);
nand U212 (N_212,In_109,In_484);
nand U213 (N_213,In_290,In_32);
nor U214 (N_214,In_130,In_418);
xnor U215 (N_215,In_480,In_22);
or U216 (N_216,In_269,In_246);
nand U217 (N_217,In_312,In_279);
xor U218 (N_218,In_140,In_339);
nand U219 (N_219,In_110,In_345);
or U220 (N_220,In_457,In_316);
nand U221 (N_221,In_261,In_259);
and U222 (N_222,In_186,In_95);
or U223 (N_223,In_335,In_29);
nand U224 (N_224,In_425,In_168);
and U225 (N_225,In_274,In_82);
nor U226 (N_226,In_293,In_315);
or U227 (N_227,In_39,In_317);
or U228 (N_228,In_93,In_273);
or U229 (N_229,In_346,In_471);
nor U230 (N_230,In_237,In_377);
and U231 (N_231,In_153,In_167);
and U232 (N_232,In_376,In_63);
nor U233 (N_233,In_27,In_366);
and U234 (N_234,In_266,In_387);
or U235 (N_235,In_55,In_360);
nor U236 (N_236,In_171,In_151);
and U237 (N_237,In_396,In_214);
or U238 (N_238,In_320,In_209);
or U239 (N_239,In_357,In_294);
and U240 (N_240,In_31,In_239);
and U241 (N_241,In_89,In_86);
nand U242 (N_242,In_124,In_455);
xnor U243 (N_243,In_69,In_211);
or U244 (N_244,In_141,In_297);
nor U245 (N_245,In_423,In_406);
or U246 (N_246,In_252,In_497);
nand U247 (N_247,In_2,In_253);
nor U248 (N_248,In_90,In_128);
nor U249 (N_249,In_70,In_221);
and U250 (N_250,In_108,In_225);
nand U251 (N_251,In_150,In_303);
nand U252 (N_252,In_381,In_32);
nor U253 (N_253,In_285,In_342);
nand U254 (N_254,In_82,In_120);
nand U255 (N_255,In_141,In_64);
nor U256 (N_256,In_243,In_28);
or U257 (N_257,In_462,In_366);
or U258 (N_258,In_106,In_395);
nand U259 (N_259,In_16,In_117);
or U260 (N_260,In_142,In_16);
nor U261 (N_261,In_41,In_491);
or U262 (N_262,In_299,In_312);
and U263 (N_263,In_308,In_116);
and U264 (N_264,In_317,In_208);
nand U265 (N_265,In_268,In_470);
nor U266 (N_266,In_251,In_75);
or U267 (N_267,In_18,In_327);
and U268 (N_268,In_185,In_465);
or U269 (N_269,In_211,In_256);
and U270 (N_270,In_145,In_402);
nor U271 (N_271,In_374,In_405);
nand U272 (N_272,In_447,In_321);
nand U273 (N_273,In_468,In_417);
nand U274 (N_274,In_251,In_33);
xnor U275 (N_275,In_499,In_404);
nor U276 (N_276,In_458,In_219);
or U277 (N_277,In_485,In_339);
and U278 (N_278,In_467,In_191);
and U279 (N_279,In_171,In_85);
and U280 (N_280,In_161,In_287);
nor U281 (N_281,In_418,In_168);
and U282 (N_282,In_172,In_147);
or U283 (N_283,In_7,In_20);
nand U284 (N_284,In_490,In_361);
and U285 (N_285,In_28,In_265);
and U286 (N_286,In_211,In_297);
or U287 (N_287,In_315,In_124);
nand U288 (N_288,In_146,In_280);
nand U289 (N_289,In_198,In_486);
or U290 (N_290,In_354,In_103);
nor U291 (N_291,In_357,In_428);
or U292 (N_292,In_360,In_434);
nor U293 (N_293,In_248,In_480);
nand U294 (N_294,In_428,In_283);
nor U295 (N_295,In_452,In_360);
and U296 (N_296,In_40,In_78);
and U297 (N_297,In_65,In_205);
nor U298 (N_298,In_256,In_138);
nor U299 (N_299,In_361,In_379);
and U300 (N_300,In_371,In_495);
xor U301 (N_301,In_95,In_48);
and U302 (N_302,In_63,In_189);
nor U303 (N_303,In_365,In_165);
xor U304 (N_304,In_99,In_127);
nor U305 (N_305,In_146,In_302);
or U306 (N_306,In_425,In_452);
and U307 (N_307,In_129,In_114);
nand U308 (N_308,In_379,In_486);
nand U309 (N_309,In_356,In_330);
or U310 (N_310,In_368,In_157);
nand U311 (N_311,In_23,In_134);
or U312 (N_312,In_161,In_93);
nor U313 (N_313,In_348,In_273);
or U314 (N_314,In_132,In_423);
nand U315 (N_315,In_376,In_342);
nand U316 (N_316,In_32,In_227);
nand U317 (N_317,In_284,In_455);
or U318 (N_318,In_242,In_287);
nand U319 (N_319,In_171,In_90);
nor U320 (N_320,In_361,In_336);
nor U321 (N_321,In_88,In_109);
nor U322 (N_322,In_127,In_359);
and U323 (N_323,In_360,In_148);
and U324 (N_324,In_166,In_465);
nand U325 (N_325,In_53,In_204);
or U326 (N_326,In_438,In_462);
xor U327 (N_327,In_490,In_306);
nor U328 (N_328,In_279,In_276);
or U329 (N_329,In_14,In_412);
nor U330 (N_330,In_150,In_381);
and U331 (N_331,In_412,In_425);
and U332 (N_332,In_219,In_294);
nor U333 (N_333,In_460,In_459);
nor U334 (N_334,In_70,In_431);
and U335 (N_335,In_390,In_265);
nor U336 (N_336,In_121,In_382);
nand U337 (N_337,In_5,In_493);
nand U338 (N_338,In_398,In_322);
or U339 (N_339,In_330,In_6);
or U340 (N_340,In_474,In_85);
nor U341 (N_341,In_449,In_334);
nor U342 (N_342,In_93,In_7);
or U343 (N_343,In_473,In_269);
xor U344 (N_344,In_324,In_439);
or U345 (N_345,In_305,In_434);
and U346 (N_346,In_149,In_57);
or U347 (N_347,In_22,In_105);
nand U348 (N_348,In_481,In_288);
and U349 (N_349,In_460,In_417);
nor U350 (N_350,In_124,In_216);
and U351 (N_351,In_283,In_55);
and U352 (N_352,In_208,In_274);
and U353 (N_353,In_74,In_245);
and U354 (N_354,In_190,In_153);
and U355 (N_355,In_24,In_448);
or U356 (N_356,In_232,In_123);
nor U357 (N_357,In_36,In_156);
or U358 (N_358,In_22,In_316);
nand U359 (N_359,In_442,In_386);
or U360 (N_360,In_232,In_443);
or U361 (N_361,In_28,In_437);
nor U362 (N_362,In_283,In_142);
and U363 (N_363,In_127,In_312);
nor U364 (N_364,In_150,In_467);
and U365 (N_365,In_29,In_79);
nand U366 (N_366,In_151,In_361);
and U367 (N_367,In_417,In_495);
and U368 (N_368,In_206,In_423);
nor U369 (N_369,In_301,In_99);
and U370 (N_370,In_15,In_246);
nor U371 (N_371,In_68,In_302);
nor U372 (N_372,In_244,In_343);
nor U373 (N_373,In_219,In_320);
xor U374 (N_374,In_486,In_453);
or U375 (N_375,In_467,In_172);
or U376 (N_376,In_294,In_255);
nand U377 (N_377,In_345,In_182);
nand U378 (N_378,In_426,In_227);
or U379 (N_379,In_148,In_468);
nor U380 (N_380,In_48,In_1);
nor U381 (N_381,In_112,In_385);
nor U382 (N_382,In_374,In_411);
and U383 (N_383,In_366,In_482);
nand U384 (N_384,In_362,In_156);
or U385 (N_385,In_51,In_316);
nand U386 (N_386,In_452,In_463);
and U387 (N_387,In_109,In_482);
and U388 (N_388,In_270,In_313);
and U389 (N_389,In_478,In_75);
nand U390 (N_390,In_333,In_412);
or U391 (N_391,In_159,In_242);
or U392 (N_392,In_246,In_240);
and U393 (N_393,In_121,In_235);
or U394 (N_394,In_54,In_130);
nor U395 (N_395,In_273,In_284);
xor U396 (N_396,In_17,In_443);
and U397 (N_397,In_79,In_272);
nand U398 (N_398,In_150,In_326);
or U399 (N_399,In_292,In_140);
or U400 (N_400,In_437,In_450);
and U401 (N_401,In_290,In_81);
nor U402 (N_402,In_282,In_89);
nor U403 (N_403,In_176,In_275);
and U404 (N_404,In_431,In_179);
or U405 (N_405,In_194,In_245);
and U406 (N_406,In_33,In_466);
nand U407 (N_407,In_234,In_218);
nor U408 (N_408,In_314,In_263);
nor U409 (N_409,In_296,In_154);
nand U410 (N_410,In_204,In_370);
nand U411 (N_411,In_146,In_489);
nand U412 (N_412,In_463,In_405);
nand U413 (N_413,In_34,In_485);
or U414 (N_414,In_366,In_421);
nand U415 (N_415,In_270,In_215);
and U416 (N_416,In_407,In_20);
nor U417 (N_417,In_401,In_336);
and U418 (N_418,In_200,In_92);
nor U419 (N_419,In_109,In_67);
or U420 (N_420,In_255,In_177);
or U421 (N_421,In_467,In_410);
nand U422 (N_422,In_451,In_66);
nand U423 (N_423,In_380,In_264);
and U424 (N_424,In_454,In_67);
or U425 (N_425,In_272,In_305);
and U426 (N_426,In_426,In_152);
nor U427 (N_427,In_155,In_213);
nand U428 (N_428,In_303,In_202);
nand U429 (N_429,In_279,In_63);
or U430 (N_430,In_76,In_457);
nor U431 (N_431,In_481,In_154);
nand U432 (N_432,In_101,In_85);
nor U433 (N_433,In_459,In_390);
nand U434 (N_434,In_220,In_17);
and U435 (N_435,In_40,In_284);
nor U436 (N_436,In_186,In_64);
nand U437 (N_437,In_323,In_379);
or U438 (N_438,In_374,In_278);
or U439 (N_439,In_381,In_213);
or U440 (N_440,In_376,In_115);
nand U441 (N_441,In_201,In_365);
or U442 (N_442,In_358,In_402);
or U443 (N_443,In_138,In_240);
nand U444 (N_444,In_444,In_221);
or U445 (N_445,In_321,In_430);
and U446 (N_446,In_171,In_62);
nor U447 (N_447,In_172,In_484);
xnor U448 (N_448,In_23,In_18);
nand U449 (N_449,In_344,In_412);
nor U450 (N_450,In_477,In_438);
xor U451 (N_451,In_299,In_116);
or U452 (N_452,In_116,In_129);
nor U453 (N_453,In_368,In_381);
nand U454 (N_454,In_44,In_222);
nand U455 (N_455,In_9,In_230);
or U456 (N_456,In_159,In_499);
and U457 (N_457,In_441,In_420);
nand U458 (N_458,In_367,In_15);
and U459 (N_459,In_359,In_381);
nor U460 (N_460,In_176,In_241);
or U461 (N_461,In_159,In_150);
and U462 (N_462,In_99,In_424);
nand U463 (N_463,In_79,In_424);
nor U464 (N_464,In_145,In_378);
nand U465 (N_465,In_29,In_36);
nor U466 (N_466,In_391,In_37);
or U467 (N_467,In_311,In_279);
nor U468 (N_468,In_63,In_477);
nand U469 (N_469,In_101,In_373);
nor U470 (N_470,In_134,In_133);
nor U471 (N_471,In_452,In_116);
nand U472 (N_472,In_2,In_335);
and U473 (N_473,In_384,In_412);
and U474 (N_474,In_27,In_344);
and U475 (N_475,In_217,In_128);
and U476 (N_476,In_173,In_87);
nor U477 (N_477,In_132,In_377);
and U478 (N_478,In_498,In_211);
nor U479 (N_479,In_224,In_18);
nor U480 (N_480,In_345,In_389);
or U481 (N_481,In_132,In_491);
nand U482 (N_482,In_363,In_40);
nand U483 (N_483,In_402,In_150);
nor U484 (N_484,In_185,In_453);
nand U485 (N_485,In_154,In_144);
and U486 (N_486,In_182,In_401);
nor U487 (N_487,In_359,In_192);
or U488 (N_488,In_468,In_275);
nor U489 (N_489,In_251,In_226);
nand U490 (N_490,In_419,In_353);
nand U491 (N_491,In_115,In_411);
or U492 (N_492,In_380,In_468);
nor U493 (N_493,In_136,In_236);
nand U494 (N_494,In_131,In_184);
or U495 (N_495,In_321,In_34);
and U496 (N_496,In_4,In_162);
and U497 (N_497,In_256,In_499);
nand U498 (N_498,In_7,In_368);
or U499 (N_499,In_171,In_175);
nand U500 (N_500,N_21,N_218);
or U501 (N_501,N_404,N_269);
and U502 (N_502,N_117,N_321);
or U503 (N_503,N_149,N_489);
and U504 (N_504,N_386,N_130);
nor U505 (N_505,N_338,N_234);
nor U506 (N_506,N_408,N_56);
nand U507 (N_507,N_291,N_146);
or U508 (N_508,N_485,N_206);
xnor U509 (N_509,N_64,N_280);
nand U510 (N_510,N_417,N_313);
and U511 (N_511,N_92,N_351);
or U512 (N_512,N_115,N_203);
or U513 (N_513,N_454,N_184);
or U514 (N_514,N_243,N_466);
nor U515 (N_515,N_390,N_101);
xor U516 (N_516,N_54,N_253);
nand U517 (N_517,N_388,N_139);
or U518 (N_518,N_170,N_204);
and U519 (N_519,N_284,N_488);
nor U520 (N_520,N_202,N_59);
nor U521 (N_521,N_434,N_180);
and U522 (N_522,N_450,N_407);
nor U523 (N_523,N_10,N_228);
nand U524 (N_524,N_199,N_239);
or U525 (N_525,N_493,N_455);
nor U526 (N_526,N_208,N_359);
and U527 (N_527,N_303,N_406);
nand U528 (N_528,N_86,N_481);
nor U529 (N_529,N_175,N_401);
or U530 (N_530,N_99,N_268);
nand U531 (N_531,N_298,N_373);
nand U532 (N_532,N_27,N_110);
nand U533 (N_533,N_151,N_60);
nand U534 (N_534,N_35,N_67);
xor U535 (N_535,N_389,N_377);
and U536 (N_536,N_415,N_128);
nand U537 (N_537,N_132,N_430);
xnor U538 (N_538,N_191,N_307);
nor U539 (N_539,N_25,N_41);
nor U540 (N_540,N_250,N_95);
xor U541 (N_541,N_49,N_440);
nor U542 (N_542,N_111,N_464);
or U543 (N_543,N_379,N_82);
nor U544 (N_544,N_248,N_167);
or U545 (N_545,N_104,N_371);
nor U546 (N_546,N_133,N_397);
or U547 (N_547,N_240,N_182);
and U548 (N_548,N_441,N_78);
and U549 (N_549,N_487,N_26);
and U550 (N_550,N_108,N_442);
nor U551 (N_551,N_312,N_479);
and U552 (N_552,N_426,N_432);
or U553 (N_553,N_84,N_142);
or U554 (N_554,N_452,N_13);
or U555 (N_555,N_224,N_44);
nand U556 (N_556,N_372,N_330);
or U557 (N_557,N_395,N_387);
or U558 (N_558,N_342,N_341);
and U559 (N_559,N_22,N_159);
nand U560 (N_560,N_255,N_403);
and U561 (N_561,N_169,N_309);
or U562 (N_562,N_1,N_102);
nand U563 (N_563,N_369,N_39);
nor U564 (N_564,N_178,N_400);
nand U565 (N_565,N_245,N_305);
nor U566 (N_566,N_433,N_123);
nand U567 (N_567,N_252,N_89);
and U568 (N_568,N_229,N_209);
or U569 (N_569,N_24,N_177);
nor U570 (N_570,N_131,N_244);
nand U571 (N_571,N_290,N_475);
and U572 (N_572,N_308,N_2);
and U573 (N_573,N_439,N_162);
and U574 (N_574,N_30,N_207);
nor U575 (N_575,N_193,N_322);
nor U576 (N_576,N_161,N_381);
or U577 (N_577,N_192,N_411);
or U578 (N_578,N_258,N_339);
nand U579 (N_579,N_136,N_414);
nor U580 (N_580,N_336,N_216);
or U581 (N_581,N_449,N_491);
nor U582 (N_582,N_91,N_398);
and U583 (N_583,N_69,N_460);
and U584 (N_584,N_0,N_468);
and U585 (N_585,N_187,N_219);
or U586 (N_586,N_16,N_85);
nor U587 (N_587,N_221,N_418);
nand U588 (N_588,N_76,N_251);
nand U589 (N_589,N_52,N_137);
nor U590 (N_590,N_57,N_135);
or U591 (N_591,N_384,N_422);
xor U592 (N_592,N_478,N_247);
and U593 (N_593,N_129,N_483);
and U594 (N_594,N_232,N_220);
nor U595 (N_595,N_157,N_141);
or U596 (N_596,N_46,N_265);
and U597 (N_597,N_74,N_292);
and U598 (N_598,N_316,N_348);
or U599 (N_599,N_443,N_168);
and U600 (N_600,N_150,N_448);
nand U601 (N_601,N_471,N_323);
and U602 (N_602,N_246,N_103);
nand U603 (N_603,N_173,N_183);
nand U604 (N_604,N_446,N_147);
nand U605 (N_605,N_282,N_494);
nand U606 (N_606,N_492,N_462);
or U607 (N_607,N_424,N_429);
or U608 (N_608,N_158,N_428);
nand U609 (N_609,N_32,N_278);
nor U610 (N_610,N_267,N_263);
or U611 (N_611,N_90,N_107);
and U612 (N_612,N_394,N_144);
nor U613 (N_613,N_324,N_461);
and U614 (N_614,N_288,N_138);
or U615 (N_615,N_451,N_306);
or U616 (N_616,N_166,N_302);
nand U617 (N_617,N_445,N_3);
or U618 (N_618,N_367,N_419);
nand U619 (N_619,N_45,N_197);
nand U620 (N_620,N_28,N_217);
nand U621 (N_621,N_334,N_71);
nor U622 (N_622,N_38,N_477);
nor U623 (N_623,N_94,N_163);
or U624 (N_624,N_11,N_125);
nand U625 (N_625,N_327,N_29);
or U626 (N_626,N_365,N_285);
nand U627 (N_627,N_4,N_378);
nand U628 (N_628,N_416,N_190);
nor U629 (N_629,N_6,N_9);
nor U630 (N_630,N_374,N_153);
and U631 (N_631,N_259,N_100);
or U632 (N_632,N_380,N_277);
nand U633 (N_633,N_42,N_332);
and U634 (N_634,N_289,N_457);
nand U635 (N_635,N_8,N_370);
and U636 (N_636,N_261,N_116);
or U637 (N_637,N_318,N_435);
and U638 (N_638,N_458,N_33);
or U639 (N_639,N_242,N_5);
and U640 (N_640,N_295,N_212);
and U641 (N_641,N_31,N_200);
nor U642 (N_642,N_65,N_304);
nand U643 (N_643,N_127,N_230);
nand U644 (N_644,N_497,N_17);
or U645 (N_645,N_459,N_156);
and U646 (N_646,N_465,N_171);
nand U647 (N_647,N_366,N_114);
nor U648 (N_648,N_476,N_287);
nor U649 (N_649,N_347,N_335);
xnor U650 (N_650,N_375,N_296);
and U651 (N_651,N_194,N_266);
nand U652 (N_652,N_112,N_317);
nand U653 (N_653,N_499,N_362);
and U654 (N_654,N_353,N_12);
and U655 (N_655,N_205,N_385);
and U656 (N_656,N_176,N_96);
or U657 (N_657,N_421,N_119);
and U658 (N_658,N_281,N_34);
or U659 (N_659,N_354,N_350);
nand U660 (N_660,N_472,N_345);
nand U661 (N_661,N_392,N_473);
nand U662 (N_662,N_198,N_357);
nand U663 (N_663,N_72,N_325);
nor U664 (N_664,N_73,N_37);
nor U665 (N_665,N_469,N_122);
nor U666 (N_666,N_405,N_346);
nor U667 (N_667,N_393,N_196);
or U668 (N_668,N_382,N_299);
nor U669 (N_669,N_225,N_188);
nor U670 (N_670,N_124,N_97);
nand U671 (N_671,N_310,N_14);
or U672 (N_672,N_83,N_257);
nor U673 (N_673,N_231,N_360);
nor U674 (N_674,N_23,N_368);
and U675 (N_675,N_262,N_179);
nand U676 (N_676,N_126,N_344);
nor U677 (N_677,N_154,N_427);
and U678 (N_678,N_376,N_340);
or U679 (N_679,N_185,N_413);
and U680 (N_680,N_227,N_80);
or U681 (N_681,N_396,N_467);
nand U682 (N_682,N_286,N_143);
or U683 (N_683,N_48,N_343);
nand U684 (N_684,N_410,N_140);
nor U685 (N_685,N_36,N_236);
and U686 (N_686,N_301,N_272);
nand U687 (N_687,N_88,N_264);
nand U688 (N_688,N_453,N_256);
and U689 (N_689,N_160,N_201);
or U690 (N_690,N_486,N_186);
nand U691 (N_691,N_189,N_331);
or U692 (N_692,N_444,N_391);
nor U693 (N_693,N_215,N_329);
nand U694 (N_694,N_490,N_355);
nand U695 (N_695,N_436,N_152);
nor U696 (N_696,N_165,N_420);
or U697 (N_697,N_463,N_315);
nand U698 (N_698,N_164,N_121);
nand U699 (N_699,N_79,N_172);
and U700 (N_700,N_63,N_226);
nor U701 (N_701,N_81,N_7);
nand U702 (N_702,N_53,N_474);
nor U703 (N_703,N_274,N_495);
and U704 (N_704,N_349,N_249);
or U705 (N_705,N_43,N_50);
and U706 (N_706,N_326,N_210);
nand U707 (N_707,N_383,N_105);
and U708 (N_708,N_498,N_98);
nor U709 (N_709,N_93,N_337);
and U710 (N_710,N_314,N_356);
and U711 (N_711,N_233,N_235);
or U712 (N_712,N_482,N_412);
nand U713 (N_713,N_40,N_222);
and U714 (N_714,N_275,N_109);
nand U715 (N_715,N_447,N_120);
and U716 (N_716,N_352,N_77);
and U717 (N_717,N_211,N_15);
xor U718 (N_718,N_402,N_70);
and U719 (N_719,N_68,N_113);
nor U720 (N_720,N_87,N_58);
and U721 (N_721,N_20,N_19);
and U722 (N_722,N_480,N_260);
nor U723 (N_723,N_319,N_148);
or U724 (N_724,N_106,N_333);
nor U725 (N_725,N_276,N_311);
nand U726 (N_726,N_47,N_456);
nand U727 (N_727,N_283,N_437);
nand U728 (N_728,N_294,N_237);
nor U729 (N_729,N_75,N_271);
nand U730 (N_730,N_145,N_279);
nand U731 (N_731,N_51,N_320);
or U732 (N_732,N_270,N_399);
nor U733 (N_733,N_425,N_297);
nand U734 (N_734,N_364,N_293);
or U735 (N_735,N_213,N_423);
or U736 (N_736,N_214,N_363);
nor U737 (N_737,N_484,N_181);
xnor U738 (N_738,N_66,N_62);
or U739 (N_739,N_496,N_361);
nor U740 (N_740,N_273,N_300);
and U741 (N_741,N_409,N_18);
nand U742 (N_742,N_223,N_61);
nor U743 (N_743,N_254,N_174);
or U744 (N_744,N_328,N_438);
nand U745 (N_745,N_155,N_358);
and U746 (N_746,N_431,N_195);
nor U747 (N_747,N_238,N_118);
nand U748 (N_748,N_134,N_241);
or U749 (N_749,N_470,N_55);
or U750 (N_750,N_353,N_320);
and U751 (N_751,N_76,N_144);
or U752 (N_752,N_308,N_454);
or U753 (N_753,N_108,N_314);
xor U754 (N_754,N_165,N_150);
and U755 (N_755,N_73,N_88);
nor U756 (N_756,N_113,N_266);
and U757 (N_757,N_24,N_0);
and U758 (N_758,N_50,N_242);
nand U759 (N_759,N_309,N_126);
nand U760 (N_760,N_414,N_14);
and U761 (N_761,N_195,N_59);
or U762 (N_762,N_195,N_210);
and U763 (N_763,N_249,N_389);
xnor U764 (N_764,N_439,N_327);
nand U765 (N_765,N_136,N_413);
nor U766 (N_766,N_384,N_337);
nor U767 (N_767,N_235,N_353);
or U768 (N_768,N_331,N_406);
or U769 (N_769,N_30,N_413);
xor U770 (N_770,N_171,N_351);
and U771 (N_771,N_15,N_229);
or U772 (N_772,N_436,N_89);
xnor U773 (N_773,N_418,N_174);
nand U774 (N_774,N_137,N_65);
nand U775 (N_775,N_233,N_253);
or U776 (N_776,N_419,N_296);
nor U777 (N_777,N_259,N_271);
nand U778 (N_778,N_249,N_176);
nand U779 (N_779,N_341,N_432);
or U780 (N_780,N_0,N_489);
nor U781 (N_781,N_250,N_41);
or U782 (N_782,N_473,N_67);
nand U783 (N_783,N_316,N_148);
or U784 (N_784,N_13,N_150);
or U785 (N_785,N_243,N_445);
xnor U786 (N_786,N_454,N_436);
nor U787 (N_787,N_266,N_419);
or U788 (N_788,N_25,N_419);
or U789 (N_789,N_374,N_308);
and U790 (N_790,N_297,N_14);
nand U791 (N_791,N_67,N_157);
or U792 (N_792,N_215,N_426);
nand U793 (N_793,N_248,N_10);
nand U794 (N_794,N_416,N_212);
and U795 (N_795,N_309,N_311);
and U796 (N_796,N_366,N_227);
nand U797 (N_797,N_89,N_435);
nand U798 (N_798,N_432,N_139);
and U799 (N_799,N_342,N_397);
and U800 (N_800,N_217,N_457);
nor U801 (N_801,N_16,N_248);
and U802 (N_802,N_275,N_448);
nand U803 (N_803,N_218,N_380);
nand U804 (N_804,N_391,N_489);
or U805 (N_805,N_286,N_458);
nand U806 (N_806,N_350,N_211);
and U807 (N_807,N_396,N_472);
nand U808 (N_808,N_186,N_238);
and U809 (N_809,N_488,N_91);
nor U810 (N_810,N_223,N_185);
nor U811 (N_811,N_401,N_15);
nor U812 (N_812,N_285,N_494);
nor U813 (N_813,N_319,N_167);
and U814 (N_814,N_460,N_44);
nor U815 (N_815,N_281,N_423);
nor U816 (N_816,N_363,N_401);
and U817 (N_817,N_108,N_0);
and U818 (N_818,N_260,N_308);
and U819 (N_819,N_62,N_157);
nand U820 (N_820,N_396,N_93);
and U821 (N_821,N_111,N_251);
or U822 (N_822,N_39,N_99);
or U823 (N_823,N_377,N_243);
or U824 (N_824,N_305,N_121);
nand U825 (N_825,N_112,N_23);
or U826 (N_826,N_253,N_301);
or U827 (N_827,N_130,N_413);
nand U828 (N_828,N_354,N_436);
and U829 (N_829,N_409,N_260);
xnor U830 (N_830,N_9,N_363);
nand U831 (N_831,N_444,N_326);
or U832 (N_832,N_478,N_347);
nand U833 (N_833,N_451,N_260);
nor U834 (N_834,N_423,N_83);
and U835 (N_835,N_152,N_19);
xnor U836 (N_836,N_317,N_291);
nand U837 (N_837,N_45,N_294);
nor U838 (N_838,N_39,N_273);
nor U839 (N_839,N_73,N_486);
and U840 (N_840,N_226,N_83);
nor U841 (N_841,N_128,N_413);
nor U842 (N_842,N_494,N_101);
or U843 (N_843,N_299,N_496);
and U844 (N_844,N_140,N_98);
nor U845 (N_845,N_279,N_1);
nor U846 (N_846,N_458,N_176);
and U847 (N_847,N_234,N_499);
nand U848 (N_848,N_366,N_162);
nor U849 (N_849,N_92,N_114);
nand U850 (N_850,N_130,N_197);
and U851 (N_851,N_148,N_149);
and U852 (N_852,N_414,N_116);
nor U853 (N_853,N_471,N_278);
or U854 (N_854,N_300,N_199);
or U855 (N_855,N_41,N_14);
or U856 (N_856,N_376,N_405);
nor U857 (N_857,N_70,N_426);
or U858 (N_858,N_318,N_207);
nand U859 (N_859,N_207,N_439);
and U860 (N_860,N_117,N_101);
nand U861 (N_861,N_168,N_441);
nand U862 (N_862,N_391,N_148);
or U863 (N_863,N_303,N_122);
and U864 (N_864,N_270,N_188);
or U865 (N_865,N_468,N_291);
nor U866 (N_866,N_110,N_399);
and U867 (N_867,N_39,N_488);
or U868 (N_868,N_9,N_38);
xnor U869 (N_869,N_72,N_403);
nand U870 (N_870,N_103,N_426);
nand U871 (N_871,N_308,N_175);
or U872 (N_872,N_86,N_254);
and U873 (N_873,N_335,N_65);
or U874 (N_874,N_442,N_88);
or U875 (N_875,N_390,N_348);
and U876 (N_876,N_162,N_161);
and U877 (N_877,N_465,N_363);
or U878 (N_878,N_425,N_377);
nor U879 (N_879,N_172,N_187);
and U880 (N_880,N_132,N_220);
and U881 (N_881,N_197,N_78);
nor U882 (N_882,N_276,N_305);
nand U883 (N_883,N_222,N_337);
nor U884 (N_884,N_149,N_408);
nand U885 (N_885,N_348,N_485);
or U886 (N_886,N_100,N_362);
and U887 (N_887,N_197,N_303);
or U888 (N_888,N_244,N_307);
nand U889 (N_889,N_268,N_66);
and U890 (N_890,N_441,N_120);
or U891 (N_891,N_353,N_67);
and U892 (N_892,N_232,N_374);
nor U893 (N_893,N_122,N_21);
and U894 (N_894,N_402,N_461);
or U895 (N_895,N_75,N_215);
or U896 (N_896,N_455,N_149);
or U897 (N_897,N_39,N_104);
nand U898 (N_898,N_38,N_133);
nor U899 (N_899,N_100,N_270);
nand U900 (N_900,N_353,N_127);
nor U901 (N_901,N_135,N_5);
or U902 (N_902,N_350,N_54);
and U903 (N_903,N_157,N_332);
nand U904 (N_904,N_262,N_316);
or U905 (N_905,N_274,N_443);
nand U906 (N_906,N_185,N_263);
and U907 (N_907,N_257,N_260);
nand U908 (N_908,N_301,N_137);
or U909 (N_909,N_221,N_411);
nor U910 (N_910,N_477,N_118);
nor U911 (N_911,N_158,N_420);
xor U912 (N_912,N_119,N_112);
nor U913 (N_913,N_10,N_268);
nor U914 (N_914,N_95,N_347);
xor U915 (N_915,N_426,N_451);
and U916 (N_916,N_392,N_22);
and U917 (N_917,N_400,N_453);
nand U918 (N_918,N_359,N_329);
nor U919 (N_919,N_292,N_229);
or U920 (N_920,N_403,N_293);
or U921 (N_921,N_45,N_68);
or U922 (N_922,N_333,N_430);
nand U923 (N_923,N_41,N_163);
or U924 (N_924,N_181,N_77);
or U925 (N_925,N_259,N_93);
and U926 (N_926,N_476,N_19);
nor U927 (N_927,N_48,N_422);
or U928 (N_928,N_393,N_482);
nand U929 (N_929,N_483,N_239);
nand U930 (N_930,N_39,N_212);
and U931 (N_931,N_326,N_457);
and U932 (N_932,N_123,N_96);
nand U933 (N_933,N_453,N_330);
or U934 (N_934,N_275,N_119);
and U935 (N_935,N_13,N_169);
nand U936 (N_936,N_145,N_377);
nand U937 (N_937,N_277,N_75);
nor U938 (N_938,N_391,N_401);
nor U939 (N_939,N_97,N_223);
xor U940 (N_940,N_165,N_183);
and U941 (N_941,N_172,N_152);
or U942 (N_942,N_204,N_333);
and U943 (N_943,N_264,N_207);
or U944 (N_944,N_141,N_252);
and U945 (N_945,N_434,N_404);
or U946 (N_946,N_194,N_352);
and U947 (N_947,N_97,N_220);
and U948 (N_948,N_352,N_183);
and U949 (N_949,N_269,N_52);
or U950 (N_950,N_436,N_14);
or U951 (N_951,N_241,N_192);
nand U952 (N_952,N_254,N_262);
nor U953 (N_953,N_257,N_454);
nor U954 (N_954,N_234,N_344);
nor U955 (N_955,N_31,N_245);
and U956 (N_956,N_349,N_66);
nand U957 (N_957,N_458,N_475);
nor U958 (N_958,N_146,N_449);
nand U959 (N_959,N_50,N_479);
nor U960 (N_960,N_346,N_182);
nor U961 (N_961,N_32,N_84);
and U962 (N_962,N_110,N_41);
nand U963 (N_963,N_311,N_279);
nand U964 (N_964,N_9,N_431);
nor U965 (N_965,N_431,N_384);
or U966 (N_966,N_23,N_229);
and U967 (N_967,N_113,N_279);
or U968 (N_968,N_413,N_60);
nand U969 (N_969,N_406,N_316);
nor U970 (N_970,N_247,N_413);
or U971 (N_971,N_172,N_167);
and U972 (N_972,N_381,N_41);
nand U973 (N_973,N_250,N_234);
nor U974 (N_974,N_2,N_265);
nand U975 (N_975,N_327,N_134);
or U976 (N_976,N_355,N_86);
nor U977 (N_977,N_279,N_415);
and U978 (N_978,N_275,N_406);
xor U979 (N_979,N_394,N_327);
or U980 (N_980,N_421,N_485);
and U981 (N_981,N_239,N_21);
and U982 (N_982,N_412,N_481);
and U983 (N_983,N_101,N_327);
and U984 (N_984,N_14,N_34);
and U985 (N_985,N_449,N_393);
nor U986 (N_986,N_342,N_130);
nor U987 (N_987,N_452,N_347);
nand U988 (N_988,N_214,N_236);
nand U989 (N_989,N_42,N_21);
or U990 (N_990,N_319,N_13);
and U991 (N_991,N_281,N_206);
nor U992 (N_992,N_5,N_456);
and U993 (N_993,N_250,N_98);
nor U994 (N_994,N_355,N_289);
nor U995 (N_995,N_223,N_311);
or U996 (N_996,N_57,N_168);
nand U997 (N_997,N_45,N_447);
nor U998 (N_998,N_205,N_113);
nor U999 (N_999,N_382,N_7);
nand U1000 (N_1000,N_506,N_870);
nand U1001 (N_1001,N_619,N_838);
nand U1002 (N_1002,N_797,N_589);
or U1003 (N_1003,N_894,N_660);
or U1004 (N_1004,N_676,N_526);
nor U1005 (N_1005,N_575,N_509);
nand U1006 (N_1006,N_849,N_898);
or U1007 (N_1007,N_779,N_766);
and U1008 (N_1008,N_523,N_610);
nor U1009 (N_1009,N_918,N_731);
or U1010 (N_1010,N_548,N_588);
nand U1011 (N_1011,N_738,N_728);
and U1012 (N_1012,N_642,N_540);
or U1013 (N_1013,N_763,N_646);
nor U1014 (N_1014,N_744,N_755);
and U1015 (N_1015,N_633,N_969);
nand U1016 (N_1016,N_819,N_916);
or U1017 (N_1017,N_950,N_917);
and U1018 (N_1018,N_514,N_832);
nand U1019 (N_1019,N_530,N_666);
nand U1020 (N_1020,N_972,N_772);
and U1021 (N_1021,N_807,N_611);
and U1022 (N_1022,N_806,N_992);
xnor U1023 (N_1023,N_770,N_576);
nand U1024 (N_1024,N_830,N_892);
and U1025 (N_1025,N_940,N_593);
nand U1026 (N_1026,N_818,N_866);
or U1027 (N_1027,N_764,N_848);
or U1028 (N_1028,N_841,N_835);
xnor U1029 (N_1029,N_953,N_935);
nor U1030 (N_1030,N_618,N_640);
or U1031 (N_1031,N_604,N_775);
or U1032 (N_1032,N_556,N_688);
nor U1033 (N_1033,N_709,N_713);
or U1034 (N_1034,N_761,N_671);
nand U1035 (N_1035,N_789,N_579);
nor U1036 (N_1036,N_977,N_941);
nor U1037 (N_1037,N_773,N_552);
and U1038 (N_1038,N_551,N_510);
and U1039 (N_1039,N_663,N_587);
nor U1040 (N_1040,N_714,N_701);
nor U1041 (N_1041,N_776,N_727);
nor U1042 (N_1042,N_737,N_822);
nor U1043 (N_1043,N_998,N_677);
nand U1044 (N_1044,N_518,N_767);
nor U1045 (N_1045,N_865,N_823);
or U1046 (N_1046,N_853,N_958);
nor U1047 (N_1047,N_783,N_915);
nor U1048 (N_1048,N_811,N_873);
nand U1049 (N_1049,N_921,N_983);
nand U1050 (N_1050,N_905,N_723);
or U1051 (N_1051,N_507,N_607);
nand U1052 (N_1052,N_996,N_769);
nor U1053 (N_1053,N_904,N_956);
nor U1054 (N_1054,N_626,N_900);
nand U1055 (N_1055,N_785,N_988);
and U1056 (N_1056,N_529,N_656);
and U1057 (N_1057,N_524,N_649);
nand U1058 (N_1058,N_750,N_631);
nor U1059 (N_1059,N_585,N_673);
nand U1060 (N_1060,N_707,N_537);
or U1061 (N_1061,N_871,N_515);
nand U1062 (N_1062,N_665,N_754);
or U1063 (N_1063,N_925,N_965);
nor U1064 (N_1064,N_628,N_814);
and U1065 (N_1065,N_934,N_564);
or U1066 (N_1066,N_568,N_795);
xor U1067 (N_1067,N_693,N_605);
and U1068 (N_1068,N_545,N_948);
or U1069 (N_1069,N_602,N_893);
nor U1070 (N_1070,N_828,N_639);
or U1071 (N_1071,N_971,N_520);
nand U1072 (N_1072,N_909,N_923);
xor U1073 (N_1073,N_979,N_682);
nand U1074 (N_1074,N_672,N_573);
nor U1075 (N_1075,N_705,N_842);
nor U1076 (N_1076,N_771,N_730);
nand U1077 (N_1077,N_897,N_538);
nor U1078 (N_1078,N_829,N_534);
nand U1079 (N_1079,N_657,N_597);
nand U1080 (N_1080,N_550,N_800);
and U1081 (N_1081,N_720,N_874);
or U1082 (N_1082,N_875,N_962);
nor U1083 (N_1083,N_691,N_743);
and U1084 (N_1084,N_859,N_946);
and U1085 (N_1085,N_768,N_989);
and U1086 (N_1086,N_792,N_827);
nor U1087 (N_1087,N_651,N_973);
nor U1088 (N_1088,N_532,N_955);
nor U1089 (N_1089,N_986,N_951);
and U1090 (N_1090,N_869,N_836);
or U1091 (N_1091,N_796,N_791);
nand U1092 (N_1092,N_804,N_747);
nor U1093 (N_1093,N_563,N_558);
xnor U1094 (N_1094,N_630,N_997);
nor U1095 (N_1095,N_601,N_999);
nand U1096 (N_1096,N_837,N_906);
or U1097 (N_1097,N_615,N_674);
or U1098 (N_1098,N_994,N_788);
and U1099 (N_1099,N_500,N_777);
or U1100 (N_1100,N_612,N_513);
and U1101 (N_1101,N_799,N_991);
and U1102 (N_1102,N_843,N_781);
nor U1103 (N_1103,N_711,N_694);
and U1104 (N_1104,N_854,N_736);
or U1105 (N_1105,N_503,N_522);
or U1106 (N_1106,N_886,N_793);
and U1107 (N_1107,N_812,N_912);
or U1108 (N_1108,N_528,N_726);
nand U1109 (N_1109,N_759,N_697);
and U1110 (N_1110,N_504,N_722);
nor U1111 (N_1111,N_724,N_982);
nor U1112 (N_1112,N_539,N_745);
or U1113 (N_1113,N_913,N_931);
or U1114 (N_1114,N_749,N_547);
and U1115 (N_1115,N_541,N_732);
nand U1116 (N_1116,N_868,N_845);
nor U1117 (N_1117,N_967,N_881);
or U1118 (N_1118,N_970,N_733);
nor U1119 (N_1119,N_544,N_856);
nor U1120 (N_1120,N_858,N_623);
nor U1121 (N_1121,N_512,N_831);
or U1122 (N_1122,N_809,N_546);
nand U1123 (N_1123,N_942,N_825);
nand U1124 (N_1124,N_715,N_937);
nor U1125 (N_1125,N_938,N_790);
nor U1126 (N_1126,N_926,N_833);
or U1127 (N_1127,N_652,N_696);
nor U1128 (N_1128,N_821,N_895);
and U1129 (N_1129,N_661,N_684);
nor U1130 (N_1130,N_888,N_911);
or U1131 (N_1131,N_620,N_641);
or U1132 (N_1132,N_706,N_553);
or U1133 (N_1133,N_710,N_901);
or U1134 (N_1134,N_824,N_954);
and U1135 (N_1135,N_699,N_778);
nand U1136 (N_1136,N_850,N_527);
nand U1137 (N_1137,N_903,N_648);
or U1138 (N_1138,N_981,N_980);
nand U1139 (N_1139,N_978,N_740);
nand U1140 (N_1140,N_712,N_536);
nand U1141 (N_1141,N_521,N_936);
nor U1142 (N_1142,N_957,N_805);
or U1143 (N_1143,N_653,N_533);
and U1144 (N_1144,N_562,N_774);
nor U1145 (N_1145,N_742,N_861);
or U1146 (N_1146,N_708,N_559);
nand U1147 (N_1147,N_802,N_862);
nand U1148 (N_1148,N_753,N_517);
or U1149 (N_1149,N_879,N_511);
nor U1150 (N_1150,N_683,N_808);
nand U1151 (N_1151,N_698,N_964);
and U1152 (N_1152,N_741,N_643);
or U1153 (N_1153,N_635,N_549);
nand U1154 (N_1154,N_929,N_692);
and U1155 (N_1155,N_867,N_590);
and U1156 (N_1156,N_751,N_690);
or U1157 (N_1157,N_721,N_525);
and U1158 (N_1158,N_974,N_650);
nand U1159 (N_1159,N_907,N_798);
or U1160 (N_1160,N_502,N_687);
nor U1161 (N_1161,N_987,N_542);
and U1162 (N_1162,N_975,N_801);
xor U1163 (N_1163,N_675,N_748);
nand U1164 (N_1164,N_782,N_614);
or U1165 (N_1165,N_944,N_945);
or U1166 (N_1166,N_902,N_908);
nor U1167 (N_1167,N_561,N_784);
nand U1168 (N_1168,N_571,N_885);
nor U1169 (N_1169,N_762,N_896);
nand U1170 (N_1170,N_670,N_968);
xor U1171 (N_1171,N_591,N_924);
nor U1172 (N_1172,N_577,N_780);
or U1173 (N_1173,N_719,N_616);
nand U1174 (N_1174,N_554,N_606);
and U1175 (N_1175,N_876,N_703);
nand U1176 (N_1176,N_949,N_860);
xor U1177 (N_1177,N_622,N_891);
and U1178 (N_1178,N_887,N_592);
nor U1179 (N_1179,N_787,N_932);
and U1180 (N_1180,N_889,N_565);
and U1181 (N_1181,N_716,N_634);
nand U1182 (N_1182,N_725,N_617);
and U1183 (N_1183,N_757,N_846);
nor U1184 (N_1184,N_567,N_679);
nor U1185 (N_1185,N_519,N_746);
nand U1186 (N_1186,N_960,N_560);
or U1187 (N_1187,N_756,N_581);
xor U1188 (N_1188,N_647,N_813);
nor U1189 (N_1189,N_882,N_557);
or U1190 (N_1190,N_717,N_718);
nor U1191 (N_1191,N_735,N_810);
or U1192 (N_1192,N_993,N_939);
and U1193 (N_1193,N_820,N_847);
nor U1194 (N_1194,N_734,N_910);
and U1195 (N_1195,N_943,N_638);
xnor U1196 (N_1196,N_899,N_678);
nand U1197 (N_1197,N_914,N_566);
nor U1198 (N_1198,N_645,N_625);
or U1199 (N_1199,N_855,N_826);
nand U1200 (N_1200,N_995,N_600);
and U1201 (N_1201,N_669,N_985);
nor U1202 (N_1202,N_599,N_840);
and U1203 (N_1203,N_844,N_572);
nor U1204 (N_1204,N_851,N_760);
and U1205 (N_1205,N_516,N_922);
or U1206 (N_1206,N_608,N_621);
nor U1207 (N_1207,N_890,N_505);
nand U1208 (N_1208,N_695,N_668);
nor U1209 (N_1209,N_655,N_919);
or U1210 (N_1210,N_786,N_662);
nand U1211 (N_1211,N_569,N_596);
nand U1212 (N_1212,N_863,N_803);
nand U1213 (N_1213,N_586,N_583);
nor U1214 (N_1214,N_872,N_700);
nor U1215 (N_1215,N_752,N_990);
or U1216 (N_1216,N_880,N_574);
nor U1217 (N_1217,N_883,N_930);
nand U1218 (N_1218,N_667,N_680);
or U1219 (N_1219,N_765,N_839);
nand U1220 (N_1220,N_961,N_702);
nor U1221 (N_1221,N_952,N_578);
and U1222 (N_1222,N_758,N_658);
or U1223 (N_1223,N_976,N_933);
or U1224 (N_1224,N_654,N_535);
nor U1225 (N_1225,N_704,N_927);
xnor U1226 (N_1226,N_595,N_664);
or U1227 (N_1227,N_632,N_816);
nor U1228 (N_1228,N_570,N_584);
and U1229 (N_1229,N_920,N_959);
or U1230 (N_1230,N_963,N_689);
nand U1231 (N_1231,N_884,N_817);
nor U1232 (N_1232,N_685,N_686);
and U1233 (N_1233,N_627,N_864);
nor U1234 (N_1234,N_543,N_877);
or U1235 (N_1235,N_594,N_947);
and U1236 (N_1236,N_794,N_852);
and U1237 (N_1237,N_609,N_624);
and U1238 (N_1238,N_555,N_857);
nand U1239 (N_1239,N_508,N_681);
and U1240 (N_1240,N_580,N_501);
nor U1241 (N_1241,N_815,N_603);
or U1242 (N_1242,N_636,N_729);
nand U1243 (N_1243,N_984,N_613);
nor U1244 (N_1244,N_739,N_637);
nand U1245 (N_1245,N_629,N_834);
and U1246 (N_1246,N_966,N_582);
nor U1247 (N_1247,N_644,N_598);
nand U1248 (N_1248,N_531,N_878);
xor U1249 (N_1249,N_659,N_928);
and U1250 (N_1250,N_664,N_633);
nor U1251 (N_1251,N_626,N_646);
or U1252 (N_1252,N_694,N_886);
nand U1253 (N_1253,N_805,N_663);
and U1254 (N_1254,N_665,N_601);
or U1255 (N_1255,N_621,N_704);
nor U1256 (N_1256,N_938,N_502);
nor U1257 (N_1257,N_887,N_805);
and U1258 (N_1258,N_938,N_844);
nand U1259 (N_1259,N_931,N_599);
nand U1260 (N_1260,N_789,N_766);
xor U1261 (N_1261,N_858,N_627);
nor U1262 (N_1262,N_529,N_799);
or U1263 (N_1263,N_573,N_931);
and U1264 (N_1264,N_700,N_516);
or U1265 (N_1265,N_598,N_658);
nor U1266 (N_1266,N_726,N_971);
nor U1267 (N_1267,N_647,N_518);
nand U1268 (N_1268,N_993,N_640);
or U1269 (N_1269,N_906,N_760);
or U1270 (N_1270,N_751,N_893);
nand U1271 (N_1271,N_697,N_812);
and U1272 (N_1272,N_518,N_696);
nor U1273 (N_1273,N_625,N_705);
nand U1274 (N_1274,N_916,N_930);
nand U1275 (N_1275,N_929,N_555);
or U1276 (N_1276,N_515,N_609);
nand U1277 (N_1277,N_676,N_565);
xnor U1278 (N_1278,N_924,N_579);
or U1279 (N_1279,N_782,N_785);
nor U1280 (N_1280,N_719,N_657);
and U1281 (N_1281,N_617,N_535);
nand U1282 (N_1282,N_625,N_758);
nor U1283 (N_1283,N_534,N_571);
nand U1284 (N_1284,N_769,N_944);
and U1285 (N_1285,N_509,N_591);
nor U1286 (N_1286,N_528,N_561);
xor U1287 (N_1287,N_536,N_774);
nand U1288 (N_1288,N_989,N_727);
or U1289 (N_1289,N_854,N_576);
and U1290 (N_1290,N_904,N_589);
or U1291 (N_1291,N_637,N_607);
and U1292 (N_1292,N_811,N_706);
nand U1293 (N_1293,N_914,N_591);
nand U1294 (N_1294,N_986,N_764);
and U1295 (N_1295,N_947,N_815);
nand U1296 (N_1296,N_935,N_741);
and U1297 (N_1297,N_501,N_551);
and U1298 (N_1298,N_983,N_985);
nor U1299 (N_1299,N_813,N_840);
nand U1300 (N_1300,N_541,N_538);
and U1301 (N_1301,N_790,N_894);
xor U1302 (N_1302,N_940,N_817);
and U1303 (N_1303,N_573,N_767);
or U1304 (N_1304,N_530,N_811);
or U1305 (N_1305,N_852,N_731);
or U1306 (N_1306,N_958,N_724);
nor U1307 (N_1307,N_662,N_614);
or U1308 (N_1308,N_875,N_656);
xor U1309 (N_1309,N_941,N_648);
and U1310 (N_1310,N_725,N_531);
nand U1311 (N_1311,N_635,N_774);
nor U1312 (N_1312,N_984,N_959);
and U1313 (N_1313,N_712,N_734);
nand U1314 (N_1314,N_919,N_750);
or U1315 (N_1315,N_606,N_644);
nor U1316 (N_1316,N_884,N_779);
nand U1317 (N_1317,N_572,N_903);
or U1318 (N_1318,N_535,N_650);
or U1319 (N_1319,N_828,N_693);
and U1320 (N_1320,N_953,N_524);
or U1321 (N_1321,N_555,N_834);
xnor U1322 (N_1322,N_887,N_999);
nand U1323 (N_1323,N_922,N_924);
or U1324 (N_1324,N_547,N_812);
nor U1325 (N_1325,N_652,N_687);
nor U1326 (N_1326,N_520,N_948);
and U1327 (N_1327,N_539,N_678);
or U1328 (N_1328,N_656,N_895);
nand U1329 (N_1329,N_916,N_898);
nor U1330 (N_1330,N_736,N_874);
nand U1331 (N_1331,N_512,N_790);
and U1332 (N_1332,N_643,N_902);
nor U1333 (N_1333,N_562,N_524);
nor U1334 (N_1334,N_510,N_777);
and U1335 (N_1335,N_975,N_777);
nand U1336 (N_1336,N_847,N_845);
and U1337 (N_1337,N_598,N_671);
nor U1338 (N_1338,N_825,N_549);
and U1339 (N_1339,N_831,N_979);
nor U1340 (N_1340,N_970,N_735);
and U1341 (N_1341,N_687,N_683);
or U1342 (N_1342,N_901,N_861);
and U1343 (N_1343,N_535,N_504);
nor U1344 (N_1344,N_609,N_811);
nand U1345 (N_1345,N_850,N_920);
nor U1346 (N_1346,N_893,N_524);
nor U1347 (N_1347,N_698,N_757);
and U1348 (N_1348,N_899,N_941);
nor U1349 (N_1349,N_636,N_820);
or U1350 (N_1350,N_560,N_761);
or U1351 (N_1351,N_692,N_689);
nor U1352 (N_1352,N_618,N_526);
or U1353 (N_1353,N_571,N_684);
nand U1354 (N_1354,N_686,N_808);
or U1355 (N_1355,N_538,N_819);
or U1356 (N_1356,N_535,N_514);
nand U1357 (N_1357,N_547,N_906);
nor U1358 (N_1358,N_540,N_943);
nand U1359 (N_1359,N_904,N_969);
nand U1360 (N_1360,N_592,N_827);
nand U1361 (N_1361,N_500,N_773);
nand U1362 (N_1362,N_689,N_708);
nor U1363 (N_1363,N_874,N_839);
nand U1364 (N_1364,N_788,N_868);
or U1365 (N_1365,N_558,N_709);
or U1366 (N_1366,N_662,N_889);
and U1367 (N_1367,N_812,N_944);
nor U1368 (N_1368,N_879,N_640);
or U1369 (N_1369,N_935,N_552);
nand U1370 (N_1370,N_704,N_972);
and U1371 (N_1371,N_819,N_723);
and U1372 (N_1372,N_989,N_685);
or U1373 (N_1373,N_802,N_794);
nand U1374 (N_1374,N_981,N_699);
and U1375 (N_1375,N_819,N_550);
nand U1376 (N_1376,N_872,N_553);
and U1377 (N_1377,N_951,N_851);
nor U1378 (N_1378,N_699,N_836);
and U1379 (N_1379,N_721,N_852);
nand U1380 (N_1380,N_892,N_742);
nor U1381 (N_1381,N_674,N_638);
nand U1382 (N_1382,N_762,N_508);
nor U1383 (N_1383,N_964,N_921);
nand U1384 (N_1384,N_608,N_837);
or U1385 (N_1385,N_897,N_699);
nand U1386 (N_1386,N_996,N_622);
and U1387 (N_1387,N_870,N_927);
xor U1388 (N_1388,N_522,N_843);
and U1389 (N_1389,N_776,N_823);
or U1390 (N_1390,N_722,N_553);
nor U1391 (N_1391,N_869,N_897);
nor U1392 (N_1392,N_729,N_806);
and U1393 (N_1393,N_916,N_754);
or U1394 (N_1394,N_979,N_573);
xor U1395 (N_1395,N_924,N_605);
and U1396 (N_1396,N_621,N_726);
nor U1397 (N_1397,N_566,N_758);
and U1398 (N_1398,N_844,N_725);
and U1399 (N_1399,N_973,N_637);
or U1400 (N_1400,N_994,N_937);
or U1401 (N_1401,N_994,N_711);
and U1402 (N_1402,N_995,N_677);
and U1403 (N_1403,N_748,N_685);
or U1404 (N_1404,N_641,N_894);
nand U1405 (N_1405,N_937,N_642);
or U1406 (N_1406,N_738,N_512);
or U1407 (N_1407,N_756,N_712);
or U1408 (N_1408,N_809,N_630);
nor U1409 (N_1409,N_912,N_606);
and U1410 (N_1410,N_680,N_885);
nand U1411 (N_1411,N_929,N_761);
or U1412 (N_1412,N_968,N_727);
nor U1413 (N_1413,N_989,N_848);
and U1414 (N_1414,N_802,N_809);
or U1415 (N_1415,N_808,N_525);
nor U1416 (N_1416,N_531,N_950);
or U1417 (N_1417,N_524,N_984);
and U1418 (N_1418,N_526,N_966);
nor U1419 (N_1419,N_923,N_866);
and U1420 (N_1420,N_660,N_753);
nand U1421 (N_1421,N_547,N_723);
nand U1422 (N_1422,N_604,N_623);
nand U1423 (N_1423,N_678,N_851);
nand U1424 (N_1424,N_953,N_518);
and U1425 (N_1425,N_560,N_937);
nor U1426 (N_1426,N_999,N_749);
nand U1427 (N_1427,N_856,N_551);
nor U1428 (N_1428,N_635,N_625);
or U1429 (N_1429,N_615,N_542);
nand U1430 (N_1430,N_915,N_838);
nand U1431 (N_1431,N_652,N_538);
nand U1432 (N_1432,N_908,N_825);
or U1433 (N_1433,N_677,N_742);
nor U1434 (N_1434,N_779,N_515);
nand U1435 (N_1435,N_826,N_608);
xnor U1436 (N_1436,N_721,N_787);
or U1437 (N_1437,N_796,N_943);
nand U1438 (N_1438,N_620,N_976);
nand U1439 (N_1439,N_692,N_975);
nor U1440 (N_1440,N_995,N_802);
nand U1441 (N_1441,N_568,N_553);
nand U1442 (N_1442,N_686,N_768);
nor U1443 (N_1443,N_610,N_531);
or U1444 (N_1444,N_782,N_861);
nand U1445 (N_1445,N_691,N_897);
nand U1446 (N_1446,N_750,N_864);
nor U1447 (N_1447,N_612,N_694);
nand U1448 (N_1448,N_658,N_530);
and U1449 (N_1449,N_899,N_580);
or U1450 (N_1450,N_749,N_793);
nand U1451 (N_1451,N_956,N_991);
or U1452 (N_1452,N_681,N_939);
and U1453 (N_1453,N_590,N_903);
nand U1454 (N_1454,N_782,N_967);
and U1455 (N_1455,N_528,N_992);
nor U1456 (N_1456,N_960,N_609);
nor U1457 (N_1457,N_890,N_739);
nor U1458 (N_1458,N_764,N_675);
nand U1459 (N_1459,N_623,N_637);
xnor U1460 (N_1460,N_531,N_989);
and U1461 (N_1461,N_883,N_648);
or U1462 (N_1462,N_979,N_894);
and U1463 (N_1463,N_714,N_621);
nor U1464 (N_1464,N_931,N_921);
nand U1465 (N_1465,N_766,N_814);
nor U1466 (N_1466,N_546,N_501);
or U1467 (N_1467,N_743,N_579);
nand U1468 (N_1468,N_502,N_580);
nor U1469 (N_1469,N_665,N_875);
and U1470 (N_1470,N_839,N_597);
xnor U1471 (N_1471,N_658,N_963);
nand U1472 (N_1472,N_765,N_794);
nand U1473 (N_1473,N_744,N_758);
or U1474 (N_1474,N_552,N_655);
nand U1475 (N_1475,N_871,N_929);
nor U1476 (N_1476,N_677,N_667);
or U1477 (N_1477,N_593,N_893);
and U1478 (N_1478,N_652,N_827);
nand U1479 (N_1479,N_953,N_775);
or U1480 (N_1480,N_744,N_901);
xor U1481 (N_1481,N_813,N_898);
nand U1482 (N_1482,N_772,N_782);
or U1483 (N_1483,N_687,N_719);
or U1484 (N_1484,N_867,N_702);
and U1485 (N_1485,N_527,N_871);
nor U1486 (N_1486,N_677,N_993);
or U1487 (N_1487,N_867,N_523);
nand U1488 (N_1488,N_967,N_508);
xor U1489 (N_1489,N_964,N_954);
or U1490 (N_1490,N_776,N_580);
and U1491 (N_1491,N_797,N_910);
nand U1492 (N_1492,N_987,N_967);
or U1493 (N_1493,N_934,N_687);
nor U1494 (N_1494,N_893,N_613);
or U1495 (N_1495,N_788,N_809);
nor U1496 (N_1496,N_999,N_612);
and U1497 (N_1497,N_791,N_831);
or U1498 (N_1498,N_882,N_501);
and U1499 (N_1499,N_679,N_850);
and U1500 (N_1500,N_1274,N_1088);
or U1501 (N_1501,N_1367,N_1357);
nand U1502 (N_1502,N_1152,N_1416);
nor U1503 (N_1503,N_1175,N_1209);
or U1504 (N_1504,N_1070,N_1306);
nor U1505 (N_1505,N_1056,N_1471);
nor U1506 (N_1506,N_1151,N_1444);
or U1507 (N_1507,N_1316,N_1079);
nand U1508 (N_1508,N_1154,N_1137);
nor U1509 (N_1509,N_1053,N_1338);
or U1510 (N_1510,N_1374,N_1269);
nor U1511 (N_1511,N_1321,N_1470);
nand U1512 (N_1512,N_1363,N_1352);
and U1513 (N_1513,N_1021,N_1093);
or U1514 (N_1514,N_1473,N_1383);
or U1515 (N_1515,N_1436,N_1465);
and U1516 (N_1516,N_1227,N_1409);
or U1517 (N_1517,N_1287,N_1210);
and U1518 (N_1518,N_1136,N_1384);
nor U1519 (N_1519,N_1236,N_1207);
and U1520 (N_1520,N_1013,N_1442);
nand U1521 (N_1521,N_1340,N_1081);
nand U1522 (N_1522,N_1171,N_1028);
nand U1523 (N_1523,N_1371,N_1423);
nand U1524 (N_1524,N_1127,N_1094);
and U1525 (N_1525,N_1435,N_1372);
or U1526 (N_1526,N_1391,N_1303);
and U1527 (N_1527,N_1092,N_1205);
nor U1528 (N_1528,N_1069,N_1189);
nor U1529 (N_1529,N_1424,N_1407);
or U1530 (N_1530,N_1030,N_1385);
and U1531 (N_1531,N_1048,N_1454);
xor U1532 (N_1532,N_1188,N_1035);
and U1533 (N_1533,N_1421,N_1472);
and U1534 (N_1534,N_1323,N_1285);
or U1535 (N_1535,N_1190,N_1174);
nor U1536 (N_1536,N_1410,N_1301);
nor U1537 (N_1537,N_1312,N_1004);
or U1538 (N_1538,N_1144,N_1119);
or U1539 (N_1539,N_1022,N_1243);
and U1540 (N_1540,N_1336,N_1467);
nor U1541 (N_1541,N_1333,N_1109);
nor U1542 (N_1542,N_1215,N_1031);
nor U1543 (N_1543,N_1469,N_1002);
nand U1544 (N_1544,N_1441,N_1033);
xor U1545 (N_1545,N_1139,N_1293);
or U1546 (N_1546,N_1439,N_1335);
nor U1547 (N_1547,N_1368,N_1281);
or U1548 (N_1548,N_1296,N_1403);
nand U1549 (N_1549,N_1085,N_1365);
and U1550 (N_1550,N_1198,N_1123);
and U1551 (N_1551,N_1286,N_1430);
nor U1552 (N_1552,N_1149,N_1478);
or U1553 (N_1553,N_1034,N_1150);
or U1554 (N_1554,N_1219,N_1107);
nor U1555 (N_1555,N_1102,N_1422);
nand U1556 (N_1556,N_1218,N_1288);
nor U1557 (N_1557,N_1006,N_1178);
and U1558 (N_1558,N_1214,N_1073);
or U1559 (N_1559,N_1495,N_1075);
nand U1560 (N_1560,N_1114,N_1350);
nand U1561 (N_1561,N_1404,N_1246);
or U1562 (N_1562,N_1084,N_1086);
nor U1563 (N_1563,N_1164,N_1052);
nand U1564 (N_1564,N_1179,N_1455);
nand U1565 (N_1565,N_1019,N_1361);
nor U1566 (N_1566,N_1419,N_1279);
or U1567 (N_1567,N_1427,N_1394);
nand U1568 (N_1568,N_1128,N_1401);
nor U1569 (N_1569,N_1124,N_1309);
or U1570 (N_1570,N_1145,N_1155);
or U1571 (N_1571,N_1320,N_1029);
nor U1572 (N_1572,N_1011,N_1110);
and U1573 (N_1573,N_1396,N_1345);
nor U1574 (N_1574,N_1337,N_1297);
and U1575 (N_1575,N_1451,N_1222);
nand U1576 (N_1576,N_1282,N_1483);
nand U1577 (N_1577,N_1169,N_1104);
nand U1578 (N_1578,N_1496,N_1118);
nor U1579 (N_1579,N_1378,N_1327);
or U1580 (N_1580,N_1057,N_1453);
or U1581 (N_1581,N_1488,N_1298);
and U1582 (N_1582,N_1490,N_1121);
xor U1583 (N_1583,N_1461,N_1484);
or U1584 (N_1584,N_1186,N_1330);
nand U1585 (N_1585,N_1414,N_1097);
nor U1586 (N_1586,N_1356,N_1200);
nand U1587 (N_1587,N_1162,N_1283);
or U1588 (N_1588,N_1456,N_1364);
nor U1589 (N_1589,N_1314,N_1193);
and U1590 (N_1590,N_1066,N_1308);
nand U1591 (N_1591,N_1299,N_1494);
nand U1592 (N_1592,N_1252,N_1106);
and U1593 (N_1593,N_1014,N_1305);
or U1594 (N_1594,N_1060,N_1242);
nor U1595 (N_1595,N_1055,N_1077);
or U1596 (N_1596,N_1418,N_1051);
or U1597 (N_1597,N_1458,N_1452);
or U1598 (N_1598,N_1485,N_1182);
and U1599 (N_1599,N_1428,N_1295);
and U1600 (N_1600,N_1486,N_1217);
nand U1601 (N_1601,N_1388,N_1225);
or U1602 (N_1602,N_1201,N_1208);
nor U1603 (N_1603,N_1163,N_1477);
nor U1604 (N_1604,N_1067,N_1277);
nand U1605 (N_1605,N_1250,N_1291);
and U1606 (N_1606,N_1042,N_1377);
nand U1607 (N_1607,N_1161,N_1278);
nand U1608 (N_1608,N_1074,N_1290);
and U1609 (N_1609,N_1313,N_1474);
nand U1610 (N_1610,N_1445,N_1234);
or U1611 (N_1611,N_1349,N_1310);
and U1612 (N_1612,N_1417,N_1261);
and U1613 (N_1613,N_1353,N_1420);
xor U1614 (N_1614,N_1468,N_1392);
and U1615 (N_1615,N_1146,N_1112);
nor U1616 (N_1616,N_1156,N_1159);
xor U1617 (N_1617,N_1206,N_1322);
and U1618 (N_1618,N_1181,N_1224);
or U1619 (N_1619,N_1005,N_1180);
or U1620 (N_1620,N_1008,N_1023);
and U1621 (N_1621,N_1091,N_1235);
xor U1622 (N_1622,N_1275,N_1213);
nand U1623 (N_1623,N_1173,N_1499);
and U1624 (N_1624,N_1177,N_1223);
or U1625 (N_1625,N_1111,N_1389);
nor U1626 (N_1626,N_1487,N_1462);
or U1627 (N_1627,N_1264,N_1370);
nand U1628 (N_1628,N_1348,N_1203);
nor U1629 (N_1629,N_1165,N_1440);
nand U1630 (N_1630,N_1492,N_1226);
nor U1631 (N_1631,N_1204,N_1239);
and U1632 (N_1632,N_1071,N_1280);
and U1633 (N_1633,N_1344,N_1354);
nor U1634 (N_1634,N_1411,N_1433);
nand U1635 (N_1635,N_1415,N_1263);
and U1636 (N_1636,N_1284,N_1294);
and U1637 (N_1637,N_1481,N_1302);
and U1638 (N_1638,N_1038,N_1270);
or U1639 (N_1639,N_1183,N_1100);
nand U1640 (N_1640,N_1429,N_1115);
and U1641 (N_1641,N_1395,N_1015);
nor U1642 (N_1642,N_1362,N_1170);
nand U1643 (N_1643,N_1341,N_1397);
nand U1644 (N_1644,N_1037,N_1120);
or U1645 (N_1645,N_1130,N_1408);
nand U1646 (N_1646,N_1447,N_1311);
xnor U1647 (N_1647,N_1065,N_1001);
nor U1648 (N_1648,N_1230,N_1491);
nor U1649 (N_1649,N_1431,N_1425);
nor U1650 (N_1650,N_1343,N_1498);
and U1651 (N_1651,N_1116,N_1047);
nand U1652 (N_1652,N_1272,N_1449);
nor U1653 (N_1653,N_1167,N_1406);
nor U1654 (N_1654,N_1135,N_1003);
nand U1655 (N_1655,N_1158,N_1479);
or U1656 (N_1656,N_1221,N_1450);
nor U1657 (N_1657,N_1108,N_1342);
nor U1658 (N_1658,N_1398,N_1131);
nand U1659 (N_1659,N_1258,N_1260);
nor U1660 (N_1660,N_1434,N_1262);
or U1661 (N_1661,N_1393,N_1054);
nand U1662 (N_1662,N_1319,N_1228);
or U1663 (N_1663,N_1039,N_1466);
or U1664 (N_1664,N_1399,N_1475);
nand U1665 (N_1665,N_1266,N_1078);
nand U1666 (N_1666,N_1493,N_1099);
nand U1667 (N_1667,N_1233,N_1460);
nor U1668 (N_1668,N_1103,N_1132);
nand U1669 (N_1669,N_1082,N_1315);
nand U1670 (N_1670,N_1489,N_1045);
nand U1671 (N_1671,N_1328,N_1253);
nand U1672 (N_1672,N_1089,N_1096);
nor U1673 (N_1673,N_1018,N_1194);
nor U1674 (N_1674,N_1050,N_1192);
nor U1675 (N_1675,N_1355,N_1049);
nor U1676 (N_1676,N_1366,N_1185);
nand U1677 (N_1677,N_1304,N_1009);
nor U1678 (N_1678,N_1231,N_1068);
nor U1679 (N_1679,N_1199,N_1497);
nor U1680 (N_1680,N_1373,N_1212);
nor U1681 (N_1681,N_1027,N_1020);
nor U1682 (N_1682,N_1405,N_1160);
nand U1683 (N_1683,N_1245,N_1375);
nor U1684 (N_1684,N_1172,N_1044);
or U1685 (N_1685,N_1147,N_1237);
nor U1686 (N_1686,N_1032,N_1090);
nor U1687 (N_1687,N_1025,N_1346);
nor U1688 (N_1688,N_1351,N_1238);
nand U1689 (N_1689,N_1457,N_1437);
or U1690 (N_1690,N_1197,N_1211);
nand U1691 (N_1691,N_1248,N_1380);
and U1692 (N_1692,N_1413,N_1292);
and U1693 (N_1693,N_1476,N_1360);
nand U1694 (N_1694,N_1000,N_1016);
or U1695 (N_1695,N_1064,N_1369);
nor U1696 (N_1696,N_1438,N_1443);
nor U1697 (N_1697,N_1463,N_1184);
nor U1698 (N_1698,N_1010,N_1347);
nand U1699 (N_1699,N_1300,N_1191);
nor U1700 (N_1700,N_1202,N_1251);
and U1701 (N_1701,N_1339,N_1072);
and U1702 (N_1702,N_1166,N_1256);
or U1703 (N_1703,N_1229,N_1113);
nand U1704 (N_1704,N_1059,N_1024);
nor U1705 (N_1705,N_1259,N_1058);
or U1706 (N_1706,N_1387,N_1358);
nand U1707 (N_1707,N_1267,N_1040);
nand U1708 (N_1708,N_1105,N_1482);
and U1709 (N_1709,N_1400,N_1083);
and U1710 (N_1710,N_1026,N_1244);
nand U1711 (N_1711,N_1036,N_1432);
or U1712 (N_1712,N_1138,N_1326);
and U1713 (N_1713,N_1125,N_1232);
or U1714 (N_1714,N_1168,N_1334);
xor U1715 (N_1715,N_1257,N_1157);
or U1716 (N_1716,N_1041,N_1087);
nor U1717 (N_1717,N_1426,N_1076);
or U1718 (N_1718,N_1061,N_1216);
nand U1719 (N_1719,N_1402,N_1122);
nand U1720 (N_1720,N_1480,N_1332);
and U1721 (N_1721,N_1381,N_1012);
or U1722 (N_1722,N_1148,N_1459);
nor U1723 (N_1723,N_1153,N_1133);
nor U1724 (N_1724,N_1062,N_1134);
or U1725 (N_1725,N_1095,N_1129);
or U1726 (N_1726,N_1098,N_1142);
or U1727 (N_1727,N_1126,N_1195);
or U1728 (N_1728,N_1017,N_1063);
or U1729 (N_1729,N_1412,N_1080);
nor U1730 (N_1730,N_1143,N_1046);
nand U1731 (N_1731,N_1464,N_1043);
and U1732 (N_1732,N_1390,N_1220);
or U1733 (N_1733,N_1382,N_1241);
nand U1734 (N_1734,N_1176,N_1117);
nor U1735 (N_1735,N_1329,N_1289);
nor U1736 (N_1736,N_1446,N_1101);
nor U1737 (N_1737,N_1254,N_1265);
or U1738 (N_1738,N_1379,N_1386);
nand U1739 (N_1739,N_1325,N_1307);
nor U1740 (N_1740,N_1249,N_1376);
nand U1741 (N_1741,N_1324,N_1196);
or U1742 (N_1742,N_1141,N_1448);
or U1743 (N_1743,N_1331,N_1273);
or U1744 (N_1744,N_1318,N_1268);
nor U1745 (N_1745,N_1271,N_1007);
nor U1746 (N_1746,N_1359,N_1240);
xor U1747 (N_1747,N_1276,N_1247);
and U1748 (N_1748,N_1140,N_1255);
nand U1749 (N_1749,N_1187,N_1317);
and U1750 (N_1750,N_1233,N_1401);
nor U1751 (N_1751,N_1371,N_1189);
or U1752 (N_1752,N_1154,N_1138);
and U1753 (N_1753,N_1085,N_1025);
xnor U1754 (N_1754,N_1436,N_1136);
or U1755 (N_1755,N_1011,N_1075);
nand U1756 (N_1756,N_1097,N_1478);
nand U1757 (N_1757,N_1330,N_1134);
nor U1758 (N_1758,N_1295,N_1483);
and U1759 (N_1759,N_1288,N_1124);
nor U1760 (N_1760,N_1213,N_1443);
xnor U1761 (N_1761,N_1310,N_1286);
nand U1762 (N_1762,N_1125,N_1258);
nand U1763 (N_1763,N_1325,N_1324);
or U1764 (N_1764,N_1140,N_1364);
and U1765 (N_1765,N_1499,N_1020);
nand U1766 (N_1766,N_1192,N_1172);
nand U1767 (N_1767,N_1362,N_1056);
and U1768 (N_1768,N_1116,N_1472);
or U1769 (N_1769,N_1287,N_1497);
nor U1770 (N_1770,N_1225,N_1013);
nand U1771 (N_1771,N_1057,N_1016);
nor U1772 (N_1772,N_1003,N_1152);
nor U1773 (N_1773,N_1310,N_1000);
and U1774 (N_1774,N_1219,N_1354);
or U1775 (N_1775,N_1245,N_1074);
and U1776 (N_1776,N_1015,N_1270);
nor U1777 (N_1777,N_1388,N_1458);
nand U1778 (N_1778,N_1228,N_1103);
nand U1779 (N_1779,N_1469,N_1234);
nand U1780 (N_1780,N_1327,N_1462);
or U1781 (N_1781,N_1270,N_1373);
or U1782 (N_1782,N_1276,N_1013);
nand U1783 (N_1783,N_1298,N_1325);
nor U1784 (N_1784,N_1133,N_1225);
nand U1785 (N_1785,N_1026,N_1066);
and U1786 (N_1786,N_1177,N_1450);
nor U1787 (N_1787,N_1308,N_1098);
nand U1788 (N_1788,N_1045,N_1416);
or U1789 (N_1789,N_1373,N_1273);
or U1790 (N_1790,N_1263,N_1444);
or U1791 (N_1791,N_1103,N_1375);
nand U1792 (N_1792,N_1054,N_1025);
or U1793 (N_1793,N_1034,N_1003);
and U1794 (N_1794,N_1413,N_1015);
nand U1795 (N_1795,N_1076,N_1151);
nand U1796 (N_1796,N_1235,N_1411);
and U1797 (N_1797,N_1195,N_1059);
and U1798 (N_1798,N_1348,N_1301);
and U1799 (N_1799,N_1336,N_1340);
nor U1800 (N_1800,N_1340,N_1310);
or U1801 (N_1801,N_1037,N_1215);
nor U1802 (N_1802,N_1314,N_1408);
and U1803 (N_1803,N_1053,N_1231);
and U1804 (N_1804,N_1255,N_1227);
and U1805 (N_1805,N_1174,N_1129);
and U1806 (N_1806,N_1081,N_1379);
nand U1807 (N_1807,N_1036,N_1311);
and U1808 (N_1808,N_1463,N_1059);
and U1809 (N_1809,N_1441,N_1008);
nand U1810 (N_1810,N_1274,N_1453);
nand U1811 (N_1811,N_1417,N_1467);
nand U1812 (N_1812,N_1315,N_1489);
nand U1813 (N_1813,N_1494,N_1047);
and U1814 (N_1814,N_1051,N_1058);
nand U1815 (N_1815,N_1046,N_1121);
nor U1816 (N_1816,N_1191,N_1295);
and U1817 (N_1817,N_1161,N_1213);
and U1818 (N_1818,N_1457,N_1224);
or U1819 (N_1819,N_1359,N_1233);
and U1820 (N_1820,N_1425,N_1450);
nor U1821 (N_1821,N_1038,N_1286);
and U1822 (N_1822,N_1237,N_1339);
nand U1823 (N_1823,N_1353,N_1093);
nor U1824 (N_1824,N_1252,N_1047);
nand U1825 (N_1825,N_1366,N_1418);
xnor U1826 (N_1826,N_1061,N_1450);
nor U1827 (N_1827,N_1158,N_1462);
nand U1828 (N_1828,N_1468,N_1081);
nor U1829 (N_1829,N_1355,N_1475);
or U1830 (N_1830,N_1291,N_1126);
and U1831 (N_1831,N_1156,N_1458);
and U1832 (N_1832,N_1248,N_1403);
nor U1833 (N_1833,N_1383,N_1386);
nand U1834 (N_1834,N_1056,N_1258);
or U1835 (N_1835,N_1294,N_1434);
and U1836 (N_1836,N_1212,N_1438);
or U1837 (N_1837,N_1477,N_1236);
or U1838 (N_1838,N_1040,N_1175);
nor U1839 (N_1839,N_1204,N_1124);
or U1840 (N_1840,N_1425,N_1096);
nand U1841 (N_1841,N_1055,N_1054);
and U1842 (N_1842,N_1352,N_1204);
and U1843 (N_1843,N_1175,N_1310);
nand U1844 (N_1844,N_1256,N_1361);
or U1845 (N_1845,N_1151,N_1222);
nand U1846 (N_1846,N_1474,N_1247);
and U1847 (N_1847,N_1341,N_1491);
nand U1848 (N_1848,N_1476,N_1377);
and U1849 (N_1849,N_1425,N_1242);
or U1850 (N_1850,N_1232,N_1430);
nand U1851 (N_1851,N_1431,N_1324);
nand U1852 (N_1852,N_1203,N_1327);
or U1853 (N_1853,N_1025,N_1249);
and U1854 (N_1854,N_1110,N_1386);
or U1855 (N_1855,N_1448,N_1261);
or U1856 (N_1856,N_1131,N_1368);
or U1857 (N_1857,N_1024,N_1223);
and U1858 (N_1858,N_1133,N_1217);
nand U1859 (N_1859,N_1181,N_1139);
and U1860 (N_1860,N_1439,N_1240);
nand U1861 (N_1861,N_1304,N_1014);
nand U1862 (N_1862,N_1482,N_1333);
and U1863 (N_1863,N_1121,N_1126);
and U1864 (N_1864,N_1498,N_1271);
and U1865 (N_1865,N_1369,N_1452);
nor U1866 (N_1866,N_1468,N_1035);
and U1867 (N_1867,N_1247,N_1080);
nor U1868 (N_1868,N_1415,N_1216);
nor U1869 (N_1869,N_1042,N_1167);
and U1870 (N_1870,N_1283,N_1327);
or U1871 (N_1871,N_1007,N_1075);
nand U1872 (N_1872,N_1191,N_1482);
and U1873 (N_1873,N_1321,N_1480);
nor U1874 (N_1874,N_1113,N_1191);
or U1875 (N_1875,N_1480,N_1323);
or U1876 (N_1876,N_1196,N_1280);
nor U1877 (N_1877,N_1349,N_1482);
or U1878 (N_1878,N_1022,N_1431);
or U1879 (N_1879,N_1435,N_1163);
nor U1880 (N_1880,N_1352,N_1323);
nand U1881 (N_1881,N_1155,N_1412);
nand U1882 (N_1882,N_1214,N_1131);
and U1883 (N_1883,N_1309,N_1473);
and U1884 (N_1884,N_1180,N_1109);
nor U1885 (N_1885,N_1432,N_1382);
nor U1886 (N_1886,N_1453,N_1286);
nand U1887 (N_1887,N_1275,N_1150);
nand U1888 (N_1888,N_1382,N_1415);
or U1889 (N_1889,N_1010,N_1172);
or U1890 (N_1890,N_1277,N_1135);
or U1891 (N_1891,N_1046,N_1147);
or U1892 (N_1892,N_1236,N_1424);
nand U1893 (N_1893,N_1097,N_1376);
and U1894 (N_1894,N_1417,N_1382);
or U1895 (N_1895,N_1040,N_1274);
nand U1896 (N_1896,N_1365,N_1370);
or U1897 (N_1897,N_1343,N_1106);
or U1898 (N_1898,N_1311,N_1259);
xor U1899 (N_1899,N_1288,N_1130);
nor U1900 (N_1900,N_1380,N_1224);
or U1901 (N_1901,N_1280,N_1445);
nor U1902 (N_1902,N_1157,N_1208);
and U1903 (N_1903,N_1104,N_1166);
and U1904 (N_1904,N_1479,N_1206);
nor U1905 (N_1905,N_1359,N_1147);
or U1906 (N_1906,N_1420,N_1033);
nor U1907 (N_1907,N_1482,N_1236);
nand U1908 (N_1908,N_1002,N_1452);
or U1909 (N_1909,N_1418,N_1332);
and U1910 (N_1910,N_1229,N_1266);
nor U1911 (N_1911,N_1411,N_1213);
nor U1912 (N_1912,N_1493,N_1457);
nor U1913 (N_1913,N_1180,N_1499);
and U1914 (N_1914,N_1128,N_1156);
and U1915 (N_1915,N_1328,N_1455);
or U1916 (N_1916,N_1156,N_1300);
nand U1917 (N_1917,N_1399,N_1392);
and U1918 (N_1918,N_1389,N_1400);
or U1919 (N_1919,N_1458,N_1238);
nand U1920 (N_1920,N_1383,N_1173);
and U1921 (N_1921,N_1210,N_1174);
nand U1922 (N_1922,N_1057,N_1206);
or U1923 (N_1923,N_1015,N_1096);
and U1924 (N_1924,N_1151,N_1376);
nand U1925 (N_1925,N_1178,N_1053);
or U1926 (N_1926,N_1152,N_1014);
and U1927 (N_1927,N_1019,N_1023);
or U1928 (N_1928,N_1375,N_1457);
or U1929 (N_1929,N_1465,N_1114);
or U1930 (N_1930,N_1087,N_1486);
nor U1931 (N_1931,N_1161,N_1374);
nor U1932 (N_1932,N_1076,N_1291);
nand U1933 (N_1933,N_1413,N_1391);
and U1934 (N_1934,N_1216,N_1157);
nor U1935 (N_1935,N_1058,N_1177);
nand U1936 (N_1936,N_1041,N_1411);
nand U1937 (N_1937,N_1487,N_1157);
and U1938 (N_1938,N_1362,N_1319);
nand U1939 (N_1939,N_1169,N_1176);
and U1940 (N_1940,N_1439,N_1279);
nor U1941 (N_1941,N_1067,N_1041);
nand U1942 (N_1942,N_1266,N_1298);
and U1943 (N_1943,N_1353,N_1004);
nor U1944 (N_1944,N_1206,N_1200);
and U1945 (N_1945,N_1390,N_1011);
nand U1946 (N_1946,N_1318,N_1248);
nand U1947 (N_1947,N_1295,N_1317);
nand U1948 (N_1948,N_1460,N_1186);
and U1949 (N_1949,N_1244,N_1359);
and U1950 (N_1950,N_1011,N_1217);
or U1951 (N_1951,N_1444,N_1420);
nand U1952 (N_1952,N_1226,N_1003);
nor U1953 (N_1953,N_1032,N_1333);
nand U1954 (N_1954,N_1337,N_1230);
or U1955 (N_1955,N_1017,N_1328);
and U1956 (N_1956,N_1430,N_1448);
and U1957 (N_1957,N_1191,N_1396);
nand U1958 (N_1958,N_1170,N_1339);
or U1959 (N_1959,N_1234,N_1431);
and U1960 (N_1960,N_1260,N_1060);
nor U1961 (N_1961,N_1085,N_1036);
or U1962 (N_1962,N_1278,N_1149);
or U1963 (N_1963,N_1498,N_1188);
and U1964 (N_1964,N_1487,N_1083);
nand U1965 (N_1965,N_1402,N_1256);
or U1966 (N_1966,N_1301,N_1388);
and U1967 (N_1967,N_1178,N_1148);
or U1968 (N_1968,N_1280,N_1278);
nor U1969 (N_1969,N_1473,N_1085);
and U1970 (N_1970,N_1159,N_1022);
or U1971 (N_1971,N_1483,N_1211);
and U1972 (N_1972,N_1498,N_1013);
nor U1973 (N_1973,N_1270,N_1446);
and U1974 (N_1974,N_1167,N_1335);
nand U1975 (N_1975,N_1490,N_1493);
nor U1976 (N_1976,N_1005,N_1450);
or U1977 (N_1977,N_1011,N_1226);
nor U1978 (N_1978,N_1281,N_1024);
or U1979 (N_1979,N_1308,N_1409);
and U1980 (N_1980,N_1417,N_1409);
or U1981 (N_1981,N_1295,N_1267);
nand U1982 (N_1982,N_1223,N_1445);
nand U1983 (N_1983,N_1012,N_1247);
nor U1984 (N_1984,N_1412,N_1346);
nor U1985 (N_1985,N_1237,N_1284);
and U1986 (N_1986,N_1284,N_1278);
and U1987 (N_1987,N_1493,N_1069);
nand U1988 (N_1988,N_1012,N_1000);
nand U1989 (N_1989,N_1136,N_1421);
or U1990 (N_1990,N_1047,N_1414);
nor U1991 (N_1991,N_1437,N_1359);
or U1992 (N_1992,N_1415,N_1345);
nand U1993 (N_1993,N_1160,N_1259);
nor U1994 (N_1994,N_1309,N_1076);
nand U1995 (N_1995,N_1250,N_1088);
nand U1996 (N_1996,N_1248,N_1070);
and U1997 (N_1997,N_1201,N_1311);
nand U1998 (N_1998,N_1422,N_1449);
nor U1999 (N_1999,N_1171,N_1258);
and U2000 (N_2000,N_1596,N_1858);
nand U2001 (N_2001,N_1820,N_1545);
and U2002 (N_2002,N_1878,N_1649);
or U2003 (N_2003,N_1584,N_1635);
nor U2004 (N_2004,N_1941,N_1560);
nor U2005 (N_2005,N_1842,N_1885);
nor U2006 (N_2006,N_1846,N_1918);
nor U2007 (N_2007,N_1511,N_1769);
and U2008 (N_2008,N_1826,N_1685);
or U2009 (N_2009,N_1542,N_1625);
nand U2010 (N_2010,N_1653,N_1686);
nand U2011 (N_2011,N_1541,N_1627);
nand U2012 (N_2012,N_1548,N_1671);
or U2013 (N_2013,N_1574,N_1978);
and U2014 (N_2014,N_1946,N_1646);
nor U2015 (N_2015,N_1644,N_1888);
nor U2016 (N_2016,N_1818,N_1933);
nor U2017 (N_2017,N_1891,N_1944);
and U2018 (N_2018,N_1934,N_1904);
nand U2019 (N_2019,N_1534,N_1506);
and U2020 (N_2020,N_1722,N_1865);
and U2021 (N_2021,N_1650,N_1823);
and U2022 (N_2022,N_1739,N_1923);
or U2023 (N_2023,N_1977,N_1965);
nor U2024 (N_2024,N_1777,N_1830);
nand U2025 (N_2025,N_1929,N_1629);
and U2026 (N_2026,N_1753,N_1822);
or U2027 (N_2027,N_1603,N_1790);
or U2028 (N_2028,N_1768,N_1515);
nor U2029 (N_2029,N_1659,N_1870);
and U2030 (N_2030,N_1866,N_1984);
nor U2031 (N_2031,N_1905,N_1553);
nand U2032 (N_2032,N_1704,N_1743);
nand U2033 (N_2033,N_1791,N_1660);
nand U2034 (N_2034,N_1589,N_1680);
nand U2035 (N_2035,N_1639,N_1779);
nor U2036 (N_2036,N_1926,N_1950);
nor U2037 (N_2037,N_1949,N_1549);
nand U2038 (N_2038,N_1519,N_1664);
nand U2039 (N_2039,N_1618,N_1691);
nor U2040 (N_2040,N_1834,N_1938);
and U2041 (N_2041,N_1624,N_1705);
nand U2042 (N_2042,N_1725,N_1766);
and U2043 (N_2043,N_1893,N_1601);
and U2044 (N_2044,N_1890,N_1637);
or U2045 (N_2045,N_1586,N_1504);
and U2046 (N_2046,N_1873,N_1764);
nor U2047 (N_2047,N_1523,N_1814);
nand U2048 (N_2048,N_1699,N_1505);
or U2049 (N_2049,N_1718,N_1735);
nor U2050 (N_2050,N_1916,N_1892);
nand U2051 (N_2051,N_1695,N_1656);
or U2052 (N_2052,N_1552,N_1837);
nand U2053 (N_2053,N_1808,N_1781);
nor U2054 (N_2054,N_1991,N_1620);
nand U2055 (N_2055,N_1719,N_1501);
nand U2056 (N_2056,N_1975,N_1784);
nor U2057 (N_2057,N_1831,N_1547);
nand U2058 (N_2058,N_1930,N_1585);
nand U2059 (N_2059,N_1692,N_1652);
nor U2060 (N_2060,N_1785,N_1630);
and U2061 (N_2061,N_1937,N_1703);
nor U2062 (N_2062,N_1587,N_1971);
or U2063 (N_2063,N_1513,N_1920);
nor U2064 (N_2064,N_1828,N_1696);
nor U2065 (N_2065,N_1988,N_1898);
nor U2066 (N_2066,N_1868,N_1895);
nand U2067 (N_2067,N_1881,N_1853);
nand U2068 (N_2068,N_1765,N_1875);
and U2069 (N_2069,N_1894,N_1788);
nand U2070 (N_2070,N_1593,N_1883);
nand U2071 (N_2071,N_1919,N_1578);
and U2072 (N_2072,N_1774,N_1507);
and U2073 (N_2073,N_1538,N_1848);
or U2074 (N_2074,N_1861,N_1573);
nand U2075 (N_2075,N_1961,N_1631);
nor U2076 (N_2076,N_1537,N_1567);
and U2077 (N_2077,N_1835,N_1517);
and U2078 (N_2078,N_1800,N_1986);
xnor U2079 (N_2079,N_1947,N_1819);
nor U2080 (N_2080,N_1924,N_1754);
nand U2081 (N_2081,N_1687,N_1674);
nor U2082 (N_2082,N_1841,N_1909);
nand U2083 (N_2083,N_1702,N_1803);
and U2084 (N_2084,N_1717,N_1518);
and U2085 (N_2085,N_1747,N_1780);
xor U2086 (N_2086,N_1748,N_1693);
nand U2087 (N_2087,N_1707,N_1556);
xor U2088 (N_2088,N_1760,N_1694);
and U2089 (N_2089,N_1623,N_1546);
nor U2090 (N_2090,N_1806,N_1733);
nor U2091 (N_2091,N_1599,N_1771);
and U2092 (N_2092,N_1973,N_1773);
and U2093 (N_2093,N_1964,N_1901);
and U2094 (N_2094,N_1613,N_1897);
and U2095 (N_2095,N_1647,N_1642);
nor U2096 (N_2096,N_1921,N_1762);
or U2097 (N_2097,N_1638,N_1665);
nor U2098 (N_2098,N_1911,N_1690);
nor U2099 (N_2099,N_1662,N_1927);
nor U2100 (N_2100,N_1999,N_1772);
nand U2101 (N_2101,N_1740,N_1915);
or U2102 (N_2102,N_1500,N_1914);
and U2103 (N_2103,N_1676,N_1634);
and U2104 (N_2104,N_1713,N_1510);
nand U2105 (N_2105,N_1522,N_1816);
or U2106 (N_2106,N_1607,N_1956);
nand U2107 (N_2107,N_1524,N_1948);
or U2108 (N_2108,N_1540,N_1606);
and U2109 (N_2109,N_1698,N_1708);
nand U2110 (N_2110,N_1532,N_1903);
nand U2111 (N_2111,N_1854,N_1786);
or U2112 (N_2112,N_1626,N_1939);
nor U2113 (N_2113,N_1966,N_1763);
nand U2114 (N_2114,N_1670,N_1809);
nor U2115 (N_2115,N_1855,N_1727);
or U2116 (N_2116,N_1571,N_1610);
nand U2117 (N_2117,N_1990,N_1579);
nor U2118 (N_2118,N_1526,N_1654);
nor U2119 (N_2119,N_1677,N_1730);
or U2120 (N_2120,N_1940,N_1935);
nor U2121 (N_2121,N_1840,N_1576);
nand U2122 (N_2122,N_1955,N_1856);
nand U2123 (N_2123,N_1968,N_1648);
nor U2124 (N_2124,N_1932,N_1509);
nand U2125 (N_2125,N_1736,N_1661);
nor U2126 (N_2126,N_1528,N_1793);
nor U2127 (N_2127,N_1770,N_1817);
and U2128 (N_2128,N_1759,N_1732);
and U2129 (N_2129,N_1863,N_1738);
or U2130 (N_2130,N_1952,N_1628);
nand U2131 (N_2131,N_1776,N_1796);
nor U2132 (N_2132,N_1907,N_1666);
and U2133 (N_2133,N_1844,N_1925);
nand U2134 (N_2134,N_1829,N_1997);
and U2135 (N_2135,N_1512,N_1896);
nor U2136 (N_2136,N_1550,N_1521);
nor U2137 (N_2137,N_1825,N_1751);
nor U2138 (N_2138,N_1859,N_1602);
nor U2139 (N_2139,N_1900,N_1590);
xor U2140 (N_2140,N_1804,N_1516);
or U2141 (N_2141,N_1689,N_1668);
and U2142 (N_2142,N_1712,N_1663);
and U2143 (N_2143,N_1864,N_1636);
nand U2144 (N_2144,N_1969,N_1643);
nand U2145 (N_2145,N_1787,N_1622);
xor U2146 (N_2146,N_1993,N_1962);
nand U2147 (N_2147,N_1852,N_1569);
nand U2148 (N_2148,N_1728,N_1797);
nor U2149 (N_2149,N_1675,N_1899);
nand U2150 (N_2150,N_1839,N_1614);
nand U2151 (N_2151,N_1598,N_1581);
or U2152 (N_2152,N_1734,N_1872);
and U2153 (N_2153,N_1688,N_1979);
or U2154 (N_2154,N_1641,N_1913);
nor U2155 (N_2155,N_1715,N_1994);
nor U2156 (N_2156,N_1700,N_1562);
or U2157 (N_2157,N_1742,N_1720);
and U2158 (N_2158,N_1681,N_1721);
nor U2159 (N_2159,N_1611,N_1758);
nand U2160 (N_2160,N_1615,N_1824);
nand U2161 (N_2161,N_1802,N_1783);
or U2162 (N_2162,N_1529,N_1530);
nand U2163 (N_2163,N_1651,N_1608);
or U2164 (N_2164,N_1959,N_1957);
nand U2165 (N_2165,N_1503,N_1943);
and U2166 (N_2166,N_1805,N_1967);
and U2167 (N_2167,N_1869,N_1794);
or U2168 (N_2168,N_1810,N_1731);
nand U2169 (N_2169,N_1591,N_1879);
or U2170 (N_2170,N_1821,N_1902);
or U2171 (N_2171,N_1672,N_1554);
nor U2172 (N_2172,N_1767,N_1750);
and U2173 (N_2173,N_1600,N_1527);
nand U2174 (N_2174,N_1544,N_1867);
nand U2175 (N_2175,N_1678,N_1827);
and U2176 (N_2176,N_1551,N_1577);
nand U2177 (N_2177,N_1884,N_1525);
nand U2178 (N_2178,N_1682,N_1726);
nor U2179 (N_2179,N_1756,N_1535);
or U2180 (N_2180,N_1813,N_1951);
nor U2181 (N_2181,N_1561,N_1565);
or U2182 (N_2182,N_1857,N_1807);
nand U2183 (N_2183,N_1958,N_1605);
or U2184 (N_2184,N_1609,N_1755);
nand U2185 (N_2185,N_1782,N_1953);
nor U2186 (N_2186,N_1928,N_1850);
or U2187 (N_2187,N_1876,N_1683);
and U2188 (N_2188,N_1849,N_1972);
nor U2189 (N_2189,N_1640,N_1558);
nor U2190 (N_2190,N_1983,N_1812);
nand U2191 (N_2191,N_1931,N_1566);
nand U2192 (N_2192,N_1621,N_1917);
or U2193 (N_2193,N_1531,N_1594);
or U2194 (N_2194,N_1655,N_1886);
and U2195 (N_2195,N_1679,N_1536);
or U2196 (N_2196,N_1746,N_1619);
and U2197 (N_2197,N_1757,N_1843);
nand U2198 (N_2198,N_1880,N_1714);
nor U2199 (N_2199,N_1709,N_1737);
and U2200 (N_2200,N_1980,N_1998);
nand U2201 (N_2201,N_1710,N_1974);
xor U2202 (N_2202,N_1862,N_1989);
nand U2203 (N_2203,N_1741,N_1580);
nor U2204 (N_2204,N_1912,N_1570);
or U2205 (N_2205,N_1723,N_1954);
or U2206 (N_2206,N_1711,N_1658);
nand U2207 (N_2207,N_1555,N_1533);
and U2208 (N_2208,N_1724,N_1789);
nand U2209 (N_2209,N_1799,N_1706);
nor U2210 (N_2210,N_1992,N_1910);
nor U2211 (N_2211,N_1612,N_1568);
nand U2212 (N_2212,N_1595,N_1798);
or U2213 (N_2213,N_1563,N_1539);
nand U2214 (N_2214,N_1701,N_1833);
or U2215 (N_2215,N_1889,N_1744);
and U2216 (N_2216,N_1582,N_1572);
or U2217 (N_2217,N_1684,N_1752);
and U2218 (N_2218,N_1557,N_1922);
or U2219 (N_2219,N_1514,N_1845);
nand U2220 (N_2220,N_1795,N_1508);
nand U2221 (N_2221,N_1970,N_1887);
and U2222 (N_2222,N_1616,N_1583);
and U2223 (N_2223,N_1564,N_1645);
nor U2224 (N_2224,N_1987,N_1906);
or U2225 (N_2225,N_1775,N_1667);
xnor U2226 (N_2226,N_1982,N_1942);
nand U2227 (N_2227,N_1543,N_1588);
and U2228 (N_2228,N_1657,N_1559);
nor U2229 (N_2229,N_1877,N_1575);
and U2230 (N_2230,N_1801,N_1745);
and U2231 (N_2231,N_1995,N_1632);
and U2232 (N_2232,N_1996,N_1832);
nand U2233 (N_2233,N_1729,N_1597);
or U2234 (N_2234,N_1633,N_1592);
nand U2235 (N_2235,N_1847,N_1981);
or U2236 (N_2236,N_1669,N_1811);
and U2237 (N_2237,N_1716,N_1815);
nand U2238 (N_2238,N_1836,N_1617);
or U2239 (N_2239,N_1976,N_1960);
nor U2240 (N_2240,N_1520,N_1673);
nor U2241 (N_2241,N_1945,N_1874);
nor U2242 (N_2242,N_1860,N_1882);
and U2243 (N_2243,N_1838,N_1985);
nor U2244 (N_2244,N_1851,N_1604);
nor U2245 (N_2245,N_1871,N_1963);
nand U2246 (N_2246,N_1778,N_1697);
nand U2247 (N_2247,N_1761,N_1908);
nand U2248 (N_2248,N_1502,N_1749);
or U2249 (N_2249,N_1792,N_1936);
nor U2250 (N_2250,N_1854,N_1510);
nand U2251 (N_2251,N_1624,N_1569);
nand U2252 (N_2252,N_1560,N_1917);
nor U2253 (N_2253,N_1592,N_1875);
nand U2254 (N_2254,N_1588,N_1605);
nand U2255 (N_2255,N_1725,N_1795);
or U2256 (N_2256,N_1678,N_1953);
and U2257 (N_2257,N_1942,N_1736);
and U2258 (N_2258,N_1993,N_1595);
or U2259 (N_2259,N_1751,N_1962);
nor U2260 (N_2260,N_1612,N_1610);
and U2261 (N_2261,N_1737,N_1946);
or U2262 (N_2262,N_1539,N_1819);
nor U2263 (N_2263,N_1808,N_1531);
and U2264 (N_2264,N_1752,N_1964);
nand U2265 (N_2265,N_1514,N_1752);
nor U2266 (N_2266,N_1504,N_1682);
and U2267 (N_2267,N_1580,N_1855);
and U2268 (N_2268,N_1988,N_1721);
xnor U2269 (N_2269,N_1802,N_1776);
nor U2270 (N_2270,N_1666,N_1910);
and U2271 (N_2271,N_1697,N_1731);
or U2272 (N_2272,N_1779,N_1921);
or U2273 (N_2273,N_1926,N_1522);
nand U2274 (N_2274,N_1673,N_1777);
nand U2275 (N_2275,N_1552,N_1683);
nand U2276 (N_2276,N_1915,N_1937);
xnor U2277 (N_2277,N_1588,N_1909);
and U2278 (N_2278,N_1996,N_1580);
nor U2279 (N_2279,N_1587,N_1745);
xnor U2280 (N_2280,N_1865,N_1771);
nand U2281 (N_2281,N_1549,N_1546);
nand U2282 (N_2282,N_1961,N_1842);
nand U2283 (N_2283,N_1539,N_1760);
nand U2284 (N_2284,N_1757,N_1845);
xor U2285 (N_2285,N_1777,N_1892);
nor U2286 (N_2286,N_1523,N_1795);
and U2287 (N_2287,N_1718,N_1803);
nor U2288 (N_2288,N_1796,N_1665);
nand U2289 (N_2289,N_1566,N_1647);
and U2290 (N_2290,N_1771,N_1674);
and U2291 (N_2291,N_1707,N_1735);
xnor U2292 (N_2292,N_1901,N_1708);
and U2293 (N_2293,N_1537,N_1601);
nor U2294 (N_2294,N_1771,N_1737);
and U2295 (N_2295,N_1917,N_1763);
nand U2296 (N_2296,N_1525,N_1914);
or U2297 (N_2297,N_1874,N_1964);
nor U2298 (N_2298,N_1984,N_1539);
or U2299 (N_2299,N_1961,N_1784);
and U2300 (N_2300,N_1814,N_1862);
or U2301 (N_2301,N_1896,N_1852);
nor U2302 (N_2302,N_1815,N_1603);
or U2303 (N_2303,N_1611,N_1697);
or U2304 (N_2304,N_1504,N_1879);
or U2305 (N_2305,N_1754,N_1795);
nor U2306 (N_2306,N_1613,N_1964);
or U2307 (N_2307,N_1612,N_1931);
or U2308 (N_2308,N_1953,N_1512);
or U2309 (N_2309,N_1877,N_1597);
nand U2310 (N_2310,N_1980,N_1957);
or U2311 (N_2311,N_1610,N_1765);
nand U2312 (N_2312,N_1784,N_1860);
nor U2313 (N_2313,N_1861,N_1648);
or U2314 (N_2314,N_1544,N_1747);
or U2315 (N_2315,N_1857,N_1819);
nand U2316 (N_2316,N_1783,N_1867);
or U2317 (N_2317,N_1855,N_1572);
nand U2318 (N_2318,N_1527,N_1766);
or U2319 (N_2319,N_1794,N_1528);
nor U2320 (N_2320,N_1988,N_1863);
and U2321 (N_2321,N_1804,N_1520);
xor U2322 (N_2322,N_1894,N_1575);
and U2323 (N_2323,N_1965,N_1625);
or U2324 (N_2324,N_1994,N_1691);
or U2325 (N_2325,N_1765,N_1987);
and U2326 (N_2326,N_1609,N_1857);
nand U2327 (N_2327,N_1614,N_1732);
xor U2328 (N_2328,N_1944,N_1809);
nor U2329 (N_2329,N_1992,N_1899);
or U2330 (N_2330,N_1988,N_1568);
nor U2331 (N_2331,N_1926,N_1794);
and U2332 (N_2332,N_1841,N_1635);
nor U2333 (N_2333,N_1594,N_1540);
nand U2334 (N_2334,N_1758,N_1576);
and U2335 (N_2335,N_1829,N_1981);
or U2336 (N_2336,N_1639,N_1868);
or U2337 (N_2337,N_1613,N_1668);
or U2338 (N_2338,N_1770,N_1997);
nand U2339 (N_2339,N_1846,N_1541);
and U2340 (N_2340,N_1648,N_1790);
nor U2341 (N_2341,N_1805,N_1503);
and U2342 (N_2342,N_1853,N_1855);
and U2343 (N_2343,N_1628,N_1715);
and U2344 (N_2344,N_1805,N_1770);
and U2345 (N_2345,N_1569,N_1700);
nand U2346 (N_2346,N_1972,N_1521);
and U2347 (N_2347,N_1937,N_1863);
or U2348 (N_2348,N_1708,N_1867);
and U2349 (N_2349,N_1791,N_1654);
nor U2350 (N_2350,N_1632,N_1607);
and U2351 (N_2351,N_1902,N_1996);
nor U2352 (N_2352,N_1892,N_1690);
or U2353 (N_2353,N_1776,N_1995);
nor U2354 (N_2354,N_1673,N_1954);
and U2355 (N_2355,N_1525,N_1909);
or U2356 (N_2356,N_1923,N_1706);
and U2357 (N_2357,N_1658,N_1742);
nor U2358 (N_2358,N_1673,N_1994);
or U2359 (N_2359,N_1941,N_1612);
or U2360 (N_2360,N_1602,N_1643);
or U2361 (N_2361,N_1590,N_1715);
or U2362 (N_2362,N_1522,N_1501);
and U2363 (N_2363,N_1658,N_1970);
nand U2364 (N_2364,N_1905,N_1919);
and U2365 (N_2365,N_1529,N_1557);
nand U2366 (N_2366,N_1523,N_1717);
or U2367 (N_2367,N_1614,N_1951);
nand U2368 (N_2368,N_1785,N_1537);
nand U2369 (N_2369,N_1807,N_1522);
nand U2370 (N_2370,N_1808,N_1673);
nor U2371 (N_2371,N_1669,N_1756);
and U2372 (N_2372,N_1566,N_1576);
nor U2373 (N_2373,N_1761,N_1503);
nand U2374 (N_2374,N_1724,N_1622);
or U2375 (N_2375,N_1513,N_1608);
nand U2376 (N_2376,N_1919,N_1684);
nand U2377 (N_2377,N_1599,N_1661);
and U2378 (N_2378,N_1968,N_1953);
xnor U2379 (N_2379,N_1715,N_1892);
nand U2380 (N_2380,N_1911,N_1973);
nor U2381 (N_2381,N_1970,N_1911);
nor U2382 (N_2382,N_1717,N_1535);
nand U2383 (N_2383,N_1651,N_1919);
nand U2384 (N_2384,N_1825,N_1837);
nor U2385 (N_2385,N_1531,N_1813);
and U2386 (N_2386,N_1797,N_1618);
and U2387 (N_2387,N_1535,N_1773);
xor U2388 (N_2388,N_1687,N_1599);
xor U2389 (N_2389,N_1732,N_1919);
or U2390 (N_2390,N_1941,N_1917);
nor U2391 (N_2391,N_1838,N_1809);
or U2392 (N_2392,N_1939,N_1604);
and U2393 (N_2393,N_1864,N_1778);
nor U2394 (N_2394,N_1968,N_1881);
and U2395 (N_2395,N_1983,N_1878);
or U2396 (N_2396,N_1667,N_1821);
nor U2397 (N_2397,N_1656,N_1991);
nor U2398 (N_2398,N_1552,N_1616);
and U2399 (N_2399,N_1505,N_1502);
nand U2400 (N_2400,N_1588,N_1871);
or U2401 (N_2401,N_1891,N_1614);
nand U2402 (N_2402,N_1835,N_1960);
and U2403 (N_2403,N_1714,N_1624);
or U2404 (N_2404,N_1983,N_1741);
or U2405 (N_2405,N_1544,N_1711);
and U2406 (N_2406,N_1742,N_1786);
nor U2407 (N_2407,N_1593,N_1814);
nand U2408 (N_2408,N_1634,N_1859);
nor U2409 (N_2409,N_1842,N_1700);
or U2410 (N_2410,N_1648,N_1594);
nor U2411 (N_2411,N_1627,N_1992);
xor U2412 (N_2412,N_1731,N_1909);
or U2413 (N_2413,N_1550,N_1733);
xor U2414 (N_2414,N_1627,N_1830);
and U2415 (N_2415,N_1745,N_1888);
nand U2416 (N_2416,N_1643,N_1876);
and U2417 (N_2417,N_1618,N_1678);
or U2418 (N_2418,N_1869,N_1753);
nor U2419 (N_2419,N_1612,N_1697);
and U2420 (N_2420,N_1554,N_1680);
nand U2421 (N_2421,N_1793,N_1600);
nand U2422 (N_2422,N_1730,N_1836);
nor U2423 (N_2423,N_1664,N_1915);
nor U2424 (N_2424,N_1663,N_1935);
or U2425 (N_2425,N_1976,N_1503);
nand U2426 (N_2426,N_1958,N_1528);
nand U2427 (N_2427,N_1730,N_1913);
nand U2428 (N_2428,N_1729,N_1697);
and U2429 (N_2429,N_1903,N_1582);
xnor U2430 (N_2430,N_1909,N_1631);
nand U2431 (N_2431,N_1769,N_1575);
and U2432 (N_2432,N_1761,N_1817);
nor U2433 (N_2433,N_1942,N_1525);
nand U2434 (N_2434,N_1845,N_1611);
or U2435 (N_2435,N_1844,N_1886);
nor U2436 (N_2436,N_1968,N_1925);
and U2437 (N_2437,N_1679,N_1964);
nand U2438 (N_2438,N_1950,N_1923);
nand U2439 (N_2439,N_1749,N_1631);
and U2440 (N_2440,N_1856,N_1731);
nor U2441 (N_2441,N_1885,N_1880);
nor U2442 (N_2442,N_1716,N_1794);
nand U2443 (N_2443,N_1833,N_1627);
or U2444 (N_2444,N_1963,N_1551);
nor U2445 (N_2445,N_1777,N_1604);
or U2446 (N_2446,N_1893,N_1828);
and U2447 (N_2447,N_1724,N_1624);
nand U2448 (N_2448,N_1527,N_1684);
or U2449 (N_2449,N_1502,N_1903);
and U2450 (N_2450,N_1709,N_1835);
xor U2451 (N_2451,N_1694,N_1794);
or U2452 (N_2452,N_1967,N_1695);
nor U2453 (N_2453,N_1699,N_1600);
nand U2454 (N_2454,N_1925,N_1634);
or U2455 (N_2455,N_1638,N_1910);
and U2456 (N_2456,N_1975,N_1866);
or U2457 (N_2457,N_1609,N_1997);
and U2458 (N_2458,N_1810,N_1546);
xnor U2459 (N_2459,N_1872,N_1892);
nand U2460 (N_2460,N_1852,N_1699);
nor U2461 (N_2461,N_1517,N_1883);
nor U2462 (N_2462,N_1786,N_1604);
nor U2463 (N_2463,N_1997,N_1605);
and U2464 (N_2464,N_1971,N_1716);
and U2465 (N_2465,N_1588,N_1918);
nand U2466 (N_2466,N_1880,N_1767);
and U2467 (N_2467,N_1731,N_1591);
nor U2468 (N_2468,N_1601,N_1608);
and U2469 (N_2469,N_1877,N_1991);
nand U2470 (N_2470,N_1635,N_1798);
and U2471 (N_2471,N_1748,N_1940);
or U2472 (N_2472,N_1540,N_1728);
nand U2473 (N_2473,N_1822,N_1956);
and U2474 (N_2474,N_1791,N_1695);
nand U2475 (N_2475,N_1830,N_1814);
nor U2476 (N_2476,N_1578,N_1983);
and U2477 (N_2477,N_1599,N_1839);
nor U2478 (N_2478,N_1852,N_1894);
or U2479 (N_2479,N_1727,N_1535);
nor U2480 (N_2480,N_1653,N_1642);
and U2481 (N_2481,N_1874,N_1816);
and U2482 (N_2482,N_1960,N_1551);
or U2483 (N_2483,N_1521,N_1863);
and U2484 (N_2484,N_1823,N_1907);
and U2485 (N_2485,N_1505,N_1870);
or U2486 (N_2486,N_1608,N_1836);
xnor U2487 (N_2487,N_1826,N_1871);
or U2488 (N_2488,N_1919,N_1737);
nor U2489 (N_2489,N_1846,N_1543);
nor U2490 (N_2490,N_1571,N_1942);
nor U2491 (N_2491,N_1745,N_1944);
nor U2492 (N_2492,N_1886,N_1538);
nor U2493 (N_2493,N_1826,N_1916);
or U2494 (N_2494,N_1932,N_1633);
and U2495 (N_2495,N_1935,N_1503);
or U2496 (N_2496,N_1687,N_1987);
nor U2497 (N_2497,N_1778,N_1594);
and U2498 (N_2498,N_1536,N_1987);
and U2499 (N_2499,N_1782,N_1664);
nand U2500 (N_2500,N_2054,N_2464);
nand U2501 (N_2501,N_2307,N_2404);
or U2502 (N_2502,N_2119,N_2298);
nor U2503 (N_2503,N_2351,N_2034);
or U2504 (N_2504,N_2094,N_2201);
nand U2505 (N_2505,N_2337,N_2282);
nor U2506 (N_2506,N_2217,N_2277);
or U2507 (N_2507,N_2406,N_2388);
nor U2508 (N_2508,N_2036,N_2010);
nor U2509 (N_2509,N_2371,N_2232);
nor U2510 (N_2510,N_2432,N_2085);
or U2511 (N_2511,N_2127,N_2383);
and U2512 (N_2512,N_2113,N_2385);
or U2513 (N_2513,N_2465,N_2005);
or U2514 (N_2514,N_2462,N_2120);
nor U2515 (N_2515,N_2394,N_2180);
nand U2516 (N_2516,N_2349,N_2227);
nor U2517 (N_2517,N_2409,N_2083);
nor U2518 (N_2518,N_2086,N_2314);
or U2519 (N_2519,N_2389,N_2016);
nor U2520 (N_2520,N_2318,N_2338);
or U2521 (N_2521,N_2025,N_2096);
or U2522 (N_2522,N_2274,N_2087);
nand U2523 (N_2523,N_2348,N_2487);
xnor U2524 (N_2524,N_2002,N_2491);
or U2525 (N_2525,N_2151,N_2142);
and U2526 (N_2526,N_2177,N_2440);
or U2527 (N_2527,N_2329,N_2181);
and U2528 (N_2528,N_2251,N_2417);
or U2529 (N_2529,N_2157,N_2077);
or U2530 (N_2530,N_2035,N_2423);
nor U2531 (N_2531,N_2270,N_2345);
or U2532 (N_2532,N_2310,N_2078);
nand U2533 (N_2533,N_2066,N_2281);
or U2534 (N_2534,N_2308,N_2279);
and U2535 (N_2535,N_2458,N_2263);
nor U2536 (N_2536,N_2296,N_2214);
nand U2537 (N_2537,N_2246,N_2355);
nand U2538 (N_2538,N_2390,N_2164);
nor U2539 (N_2539,N_2340,N_2288);
and U2540 (N_2540,N_2323,N_2006);
or U2541 (N_2541,N_2075,N_2468);
nand U2542 (N_2542,N_2369,N_2115);
or U2543 (N_2543,N_2199,N_2461);
nand U2544 (N_2544,N_2488,N_2029);
nor U2545 (N_2545,N_2499,N_2101);
and U2546 (N_2546,N_2073,N_2255);
and U2547 (N_2547,N_2140,N_2291);
or U2548 (N_2548,N_2289,N_2426);
nand U2549 (N_2549,N_2474,N_2249);
or U2550 (N_2550,N_2354,N_2108);
xnor U2551 (N_2551,N_2293,N_2490);
or U2552 (N_2552,N_2254,N_2100);
and U2553 (N_2553,N_2334,N_2187);
and U2554 (N_2554,N_2141,N_2067);
nor U2555 (N_2555,N_2366,N_2200);
and U2556 (N_2556,N_2379,N_2081);
nand U2557 (N_2557,N_2273,N_2301);
and U2558 (N_2558,N_2074,N_2215);
or U2559 (N_2559,N_2186,N_2204);
nand U2560 (N_2560,N_2213,N_2221);
nor U2561 (N_2561,N_2429,N_2012);
or U2562 (N_2562,N_2033,N_2359);
nand U2563 (N_2563,N_2168,N_2292);
and U2564 (N_2564,N_2072,N_2216);
and U2565 (N_2565,N_2211,N_2138);
nand U2566 (N_2566,N_2320,N_2102);
xnor U2567 (N_2567,N_2150,N_2370);
nor U2568 (N_2568,N_2088,N_2469);
and U2569 (N_2569,N_2003,N_2226);
nor U2570 (N_2570,N_2401,N_2433);
and U2571 (N_2571,N_2365,N_2079);
nor U2572 (N_2572,N_2363,N_2117);
and U2573 (N_2573,N_2357,N_2449);
nor U2574 (N_2574,N_2387,N_2299);
or U2575 (N_2575,N_2418,N_2239);
or U2576 (N_2576,N_2341,N_2410);
and U2577 (N_2577,N_2009,N_2228);
nand U2578 (N_2578,N_2466,N_2436);
or U2579 (N_2579,N_2172,N_2328);
nand U2580 (N_2580,N_2122,N_2146);
nand U2581 (N_2581,N_2070,N_2060);
and U2582 (N_2582,N_2159,N_2287);
xor U2583 (N_2583,N_2059,N_2495);
or U2584 (N_2584,N_2421,N_2037);
or U2585 (N_2585,N_2017,N_2062);
nand U2586 (N_2586,N_2111,N_2104);
or U2587 (N_2587,N_2399,N_2128);
nand U2588 (N_2588,N_2040,N_2424);
and U2589 (N_2589,N_2250,N_2256);
nand U2590 (N_2590,N_2326,N_2405);
or U2591 (N_2591,N_2472,N_2173);
and U2592 (N_2592,N_2121,N_2098);
and U2593 (N_2593,N_2032,N_2391);
or U2594 (N_2594,N_2346,N_2286);
and U2595 (N_2595,N_2428,N_2445);
xor U2596 (N_2596,N_2455,N_2191);
or U2597 (N_2597,N_2198,N_2144);
nand U2598 (N_2598,N_2044,N_2243);
or U2599 (N_2599,N_2482,N_2265);
and U2600 (N_2600,N_2361,N_2219);
and U2601 (N_2601,N_2295,N_2375);
nand U2602 (N_2602,N_2107,N_2386);
and U2603 (N_2603,N_2306,N_2209);
or U2604 (N_2604,N_2343,N_2166);
nand U2605 (N_2605,N_2378,N_2097);
nor U2606 (N_2606,N_2007,N_2076);
or U2607 (N_2607,N_2133,N_2064);
nor U2608 (N_2608,N_2099,N_2347);
and U2609 (N_2609,N_2413,N_2480);
xor U2610 (N_2610,N_2224,N_2161);
or U2611 (N_2611,N_2210,N_2152);
and U2612 (N_2612,N_2312,N_2145);
nor U2613 (N_2613,N_2027,N_2171);
nand U2614 (N_2614,N_2169,N_2350);
nand U2615 (N_2615,N_2470,N_2234);
nand U2616 (N_2616,N_2089,N_2008);
or U2617 (N_2617,N_2330,N_2207);
nand U2618 (N_2618,N_2014,N_2158);
nand U2619 (N_2619,N_2130,N_2407);
nand U2620 (N_2620,N_2167,N_2065);
and U2621 (N_2621,N_2460,N_2202);
or U2622 (N_2622,N_2283,N_2155);
nand U2623 (N_2623,N_2176,N_2114);
or U2624 (N_2624,N_2162,N_2353);
nand U2625 (N_2625,N_2484,N_2303);
nor U2626 (N_2626,N_2045,N_2396);
nor U2627 (N_2627,N_2425,N_2205);
nor U2628 (N_2628,N_2206,N_2230);
or U2629 (N_2629,N_2367,N_2236);
and U2630 (N_2630,N_2103,N_2061);
nand U2631 (N_2631,N_2023,N_2368);
xnor U2632 (N_2632,N_2362,N_2473);
nor U2633 (N_2633,N_2190,N_2153);
xnor U2634 (N_2634,N_2165,N_2233);
nand U2635 (N_2635,N_2011,N_2313);
or U2636 (N_2636,N_2364,N_2196);
or U2637 (N_2637,N_2414,N_2446);
and U2638 (N_2638,N_2327,N_2319);
nor U2639 (N_2639,N_2380,N_2360);
or U2640 (N_2640,N_2056,N_2193);
and U2641 (N_2641,N_2498,N_2280);
or U2642 (N_2642,N_2080,N_2124);
nand U2643 (N_2643,N_2112,N_2197);
nand U2644 (N_2644,N_2048,N_2271);
and U2645 (N_2645,N_2245,N_2231);
nand U2646 (N_2646,N_2203,N_2454);
or U2647 (N_2647,N_2188,N_2477);
nor U2648 (N_2648,N_2252,N_2212);
or U2649 (N_2649,N_2049,N_2438);
nor U2650 (N_2650,N_2038,N_2185);
or U2651 (N_2651,N_2090,N_2106);
nor U2652 (N_2652,N_2134,N_2058);
or U2653 (N_2653,N_2195,N_2358);
and U2654 (N_2654,N_2235,N_2093);
nand U2655 (N_2655,N_2039,N_2430);
nand U2656 (N_2656,N_2109,N_2492);
and U2657 (N_2657,N_2194,N_2384);
nor U2658 (N_2658,N_2435,N_2021);
nor U2659 (N_2659,N_2459,N_2092);
and U2660 (N_2660,N_2131,N_2451);
or U2661 (N_2661,N_2031,N_2486);
nor U2662 (N_2662,N_2456,N_2163);
or U2663 (N_2663,N_2137,N_2020);
or U2664 (N_2664,N_2400,N_2237);
nand U2665 (N_2665,N_2170,N_2290);
or U2666 (N_2666,N_2053,N_2463);
and U2667 (N_2667,N_2448,N_2397);
or U2668 (N_2668,N_2052,N_2339);
nand U2669 (N_2669,N_2024,N_2336);
or U2670 (N_2670,N_2091,N_2116);
nor U2671 (N_2671,N_2489,N_2223);
or U2672 (N_2672,N_2278,N_2218);
nor U2673 (N_2673,N_2257,N_2377);
or U2674 (N_2674,N_2304,N_2485);
nor U2675 (N_2675,N_2125,N_2483);
nand U2676 (N_2676,N_2497,N_2325);
and U2677 (N_2677,N_2356,N_2395);
or U2678 (N_2678,N_2147,N_2324);
nand U2679 (N_2679,N_2174,N_2297);
or U2680 (N_2680,N_2043,N_2179);
or U2681 (N_2681,N_2476,N_2261);
or U2682 (N_2682,N_2285,N_2276);
nor U2683 (N_2683,N_2392,N_2478);
or U2684 (N_2684,N_2220,N_2335);
nand U2685 (N_2685,N_2266,N_2332);
or U2686 (N_2686,N_2015,N_2132);
nand U2687 (N_2687,N_2178,N_2022);
xnor U2688 (N_2688,N_2105,N_2305);
or U2689 (N_2689,N_2260,N_2019);
nor U2690 (N_2690,N_2434,N_2057);
nand U2691 (N_2691,N_2442,N_2042);
nor U2692 (N_2692,N_2018,N_2148);
nand U2693 (N_2693,N_2479,N_2262);
nand U2694 (N_2694,N_2457,N_2129);
and U2695 (N_2695,N_2309,N_2183);
or U2696 (N_2696,N_2055,N_2415);
and U2697 (N_2697,N_2192,N_2381);
xor U2698 (N_2698,N_2275,N_2082);
nor U2699 (N_2699,N_2135,N_2452);
nor U2700 (N_2700,N_2222,N_2139);
or U2701 (N_2701,N_2344,N_2450);
nand U2702 (N_2702,N_2030,N_2481);
nor U2703 (N_2703,N_2416,N_2041);
or U2704 (N_2704,N_2373,N_2259);
nor U2705 (N_2705,N_2241,N_2422);
or U2706 (N_2706,N_2013,N_2149);
and U2707 (N_2707,N_2268,N_2331);
nand U2708 (N_2708,N_2431,N_2123);
nand U2709 (N_2709,N_2154,N_2284);
and U2710 (N_2710,N_2126,N_2240);
or U2711 (N_2711,N_2447,N_2496);
nor U2712 (N_2712,N_2136,N_2372);
and U2713 (N_2713,N_2412,N_2467);
or U2714 (N_2714,N_2028,N_2051);
nand U2715 (N_2715,N_2068,N_2316);
or U2716 (N_2716,N_2493,N_2352);
or U2717 (N_2717,N_2403,N_2267);
and U2718 (N_2718,N_2175,N_2302);
and U2719 (N_2719,N_2411,N_2071);
and U2720 (N_2720,N_2000,N_2311);
and U2721 (N_2721,N_2471,N_2253);
nor U2722 (N_2722,N_2182,N_2315);
and U2723 (N_2723,N_2248,N_2160);
nand U2724 (N_2724,N_2374,N_2342);
nand U2725 (N_2725,N_2376,N_2238);
nor U2726 (N_2726,N_2382,N_2244);
nor U2727 (N_2727,N_2063,N_2264);
nor U2728 (N_2728,N_2427,N_2322);
or U2729 (N_2729,N_2095,N_2156);
nor U2730 (N_2730,N_2333,N_2439);
xnor U2731 (N_2731,N_2272,N_2393);
nor U2732 (N_2732,N_2437,N_2419);
or U2733 (N_2733,N_2069,N_2046);
or U2734 (N_2734,N_2184,N_2050);
or U2735 (N_2735,N_2118,N_2321);
nand U2736 (N_2736,N_2420,N_2047);
nand U2737 (N_2737,N_2294,N_2225);
nand U2738 (N_2738,N_2229,N_2026);
or U2739 (N_2739,N_2247,N_2300);
and U2740 (N_2740,N_2453,N_2084);
or U2741 (N_2741,N_2398,N_2408);
nand U2742 (N_2742,N_2143,N_2402);
nand U2743 (N_2743,N_2475,N_2494);
xnor U2744 (N_2744,N_2317,N_2189);
nand U2745 (N_2745,N_2110,N_2242);
and U2746 (N_2746,N_2001,N_2004);
and U2747 (N_2747,N_2443,N_2208);
or U2748 (N_2748,N_2258,N_2441);
nand U2749 (N_2749,N_2269,N_2444);
and U2750 (N_2750,N_2406,N_2007);
nand U2751 (N_2751,N_2056,N_2027);
or U2752 (N_2752,N_2401,N_2007);
nor U2753 (N_2753,N_2264,N_2444);
nor U2754 (N_2754,N_2409,N_2233);
and U2755 (N_2755,N_2044,N_2126);
nor U2756 (N_2756,N_2223,N_2476);
or U2757 (N_2757,N_2462,N_2211);
and U2758 (N_2758,N_2136,N_2204);
nor U2759 (N_2759,N_2118,N_2222);
and U2760 (N_2760,N_2116,N_2233);
nor U2761 (N_2761,N_2290,N_2187);
nand U2762 (N_2762,N_2338,N_2294);
nor U2763 (N_2763,N_2077,N_2462);
nand U2764 (N_2764,N_2152,N_2433);
nand U2765 (N_2765,N_2131,N_2118);
and U2766 (N_2766,N_2284,N_2085);
and U2767 (N_2767,N_2422,N_2009);
and U2768 (N_2768,N_2374,N_2404);
or U2769 (N_2769,N_2441,N_2094);
or U2770 (N_2770,N_2421,N_2265);
nor U2771 (N_2771,N_2106,N_2473);
and U2772 (N_2772,N_2075,N_2198);
nand U2773 (N_2773,N_2002,N_2293);
xor U2774 (N_2774,N_2082,N_2420);
nor U2775 (N_2775,N_2274,N_2354);
or U2776 (N_2776,N_2311,N_2483);
xor U2777 (N_2777,N_2299,N_2482);
and U2778 (N_2778,N_2450,N_2136);
nand U2779 (N_2779,N_2227,N_2337);
nand U2780 (N_2780,N_2417,N_2205);
or U2781 (N_2781,N_2329,N_2251);
or U2782 (N_2782,N_2426,N_2338);
and U2783 (N_2783,N_2160,N_2183);
or U2784 (N_2784,N_2343,N_2155);
or U2785 (N_2785,N_2075,N_2052);
and U2786 (N_2786,N_2302,N_2095);
or U2787 (N_2787,N_2283,N_2182);
or U2788 (N_2788,N_2110,N_2178);
and U2789 (N_2789,N_2077,N_2426);
or U2790 (N_2790,N_2109,N_2067);
nand U2791 (N_2791,N_2189,N_2492);
nand U2792 (N_2792,N_2415,N_2491);
and U2793 (N_2793,N_2280,N_2004);
nor U2794 (N_2794,N_2412,N_2334);
nand U2795 (N_2795,N_2444,N_2343);
and U2796 (N_2796,N_2164,N_2418);
nand U2797 (N_2797,N_2056,N_2429);
nor U2798 (N_2798,N_2100,N_2451);
or U2799 (N_2799,N_2263,N_2252);
and U2800 (N_2800,N_2265,N_2203);
nor U2801 (N_2801,N_2051,N_2433);
nand U2802 (N_2802,N_2266,N_2030);
or U2803 (N_2803,N_2058,N_2281);
nand U2804 (N_2804,N_2359,N_2482);
nor U2805 (N_2805,N_2225,N_2319);
or U2806 (N_2806,N_2358,N_2296);
or U2807 (N_2807,N_2055,N_2490);
nand U2808 (N_2808,N_2120,N_2223);
and U2809 (N_2809,N_2304,N_2045);
or U2810 (N_2810,N_2467,N_2247);
and U2811 (N_2811,N_2210,N_2128);
nand U2812 (N_2812,N_2192,N_2257);
or U2813 (N_2813,N_2119,N_2078);
nor U2814 (N_2814,N_2155,N_2121);
nor U2815 (N_2815,N_2213,N_2047);
xor U2816 (N_2816,N_2315,N_2426);
nand U2817 (N_2817,N_2394,N_2127);
nand U2818 (N_2818,N_2431,N_2269);
nand U2819 (N_2819,N_2205,N_2107);
and U2820 (N_2820,N_2262,N_2270);
nand U2821 (N_2821,N_2013,N_2294);
or U2822 (N_2822,N_2475,N_2341);
and U2823 (N_2823,N_2253,N_2364);
nand U2824 (N_2824,N_2096,N_2407);
or U2825 (N_2825,N_2073,N_2061);
nor U2826 (N_2826,N_2221,N_2406);
and U2827 (N_2827,N_2413,N_2099);
nand U2828 (N_2828,N_2197,N_2037);
nor U2829 (N_2829,N_2442,N_2150);
or U2830 (N_2830,N_2449,N_2013);
nand U2831 (N_2831,N_2002,N_2246);
or U2832 (N_2832,N_2373,N_2380);
nand U2833 (N_2833,N_2289,N_2305);
nand U2834 (N_2834,N_2097,N_2043);
and U2835 (N_2835,N_2084,N_2145);
or U2836 (N_2836,N_2133,N_2198);
nor U2837 (N_2837,N_2019,N_2472);
nand U2838 (N_2838,N_2498,N_2128);
or U2839 (N_2839,N_2039,N_2198);
nor U2840 (N_2840,N_2344,N_2485);
nor U2841 (N_2841,N_2208,N_2026);
nor U2842 (N_2842,N_2442,N_2334);
or U2843 (N_2843,N_2383,N_2296);
and U2844 (N_2844,N_2075,N_2081);
and U2845 (N_2845,N_2397,N_2394);
or U2846 (N_2846,N_2280,N_2006);
nor U2847 (N_2847,N_2156,N_2330);
nor U2848 (N_2848,N_2044,N_2270);
or U2849 (N_2849,N_2390,N_2234);
or U2850 (N_2850,N_2079,N_2002);
or U2851 (N_2851,N_2417,N_2465);
and U2852 (N_2852,N_2107,N_2436);
or U2853 (N_2853,N_2280,N_2126);
nor U2854 (N_2854,N_2149,N_2421);
or U2855 (N_2855,N_2265,N_2243);
nand U2856 (N_2856,N_2219,N_2372);
nand U2857 (N_2857,N_2325,N_2253);
xor U2858 (N_2858,N_2017,N_2116);
nor U2859 (N_2859,N_2461,N_2279);
nand U2860 (N_2860,N_2165,N_2020);
nor U2861 (N_2861,N_2233,N_2294);
or U2862 (N_2862,N_2158,N_2402);
or U2863 (N_2863,N_2110,N_2193);
nand U2864 (N_2864,N_2215,N_2329);
or U2865 (N_2865,N_2004,N_2476);
or U2866 (N_2866,N_2158,N_2466);
and U2867 (N_2867,N_2339,N_2303);
nor U2868 (N_2868,N_2016,N_2321);
or U2869 (N_2869,N_2448,N_2238);
nor U2870 (N_2870,N_2209,N_2377);
or U2871 (N_2871,N_2038,N_2371);
nand U2872 (N_2872,N_2036,N_2292);
nor U2873 (N_2873,N_2375,N_2180);
or U2874 (N_2874,N_2348,N_2216);
and U2875 (N_2875,N_2181,N_2492);
and U2876 (N_2876,N_2065,N_2216);
nor U2877 (N_2877,N_2114,N_2095);
nand U2878 (N_2878,N_2088,N_2336);
or U2879 (N_2879,N_2382,N_2281);
or U2880 (N_2880,N_2119,N_2485);
or U2881 (N_2881,N_2453,N_2463);
and U2882 (N_2882,N_2225,N_2157);
nand U2883 (N_2883,N_2149,N_2470);
nand U2884 (N_2884,N_2427,N_2099);
and U2885 (N_2885,N_2435,N_2142);
and U2886 (N_2886,N_2195,N_2469);
and U2887 (N_2887,N_2166,N_2012);
and U2888 (N_2888,N_2005,N_2179);
nand U2889 (N_2889,N_2155,N_2246);
or U2890 (N_2890,N_2457,N_2316);
nor U2891 (N_2891,N_2067,N_2343);
or U2892 (N_2892,N_2364,N_2125);
nand U2893 (N_2893,N_2454,N_2367);
and U2894 (N_2894,N_2329,N_2162);
nand U2895 (N_2895,N_2134,N_2403);
and U2896 (N_2896,N_2263,N_2173);
and U2897 (N_2897,N_2490,N_2314);
or U2898 (N_2898,N_2454,N_2291);
and U2899 (N_2899,N_2027,N_2291);
nor U2900 (N_2900,N_2222,N_2221);
nand U2901 (N_2901,N_2317,N_2060);
nor U2902 (N_2902,N_2498,N_2260);
and U2903 (N_2903,N_2414,N_2231);
or U2904 (N_2904,N_2226,N_2326);
nor U2905 (N_2905,N_2318,N_2347);
or U2906 (N_2906,N_2136,N_2210);
or U2907 (N_2907,N_2003,N_2063);
nor U2908 (N_2908,N_2128,N_2357);
nand U2909 (N_2909,N_2095,N_2267);
nor U2910 (N_2910,N_2098,N_2438);
and U2911 (N_2911,N_2440,N_2315);
nor U2912 (N_2912,N_2478,N_2056);
nand U2913 (N_2913,N_2403,N_2020);
nor U2914 (N_2914,N_2069,N_2148);
or U2915 (N_2915,N_2160,N_2424);
nor U2916 (N_2916,N_2289,N_2242);
and U2917 (N_2917,N_2016,N_2441);
nor U2918 (N_2918,N_2105,N_2397);
nor U2919 (N_2919,N_2007,N_2378);
nor U2920 (N_2920,N_2229,N_2386);
and U2921 (N_2921,N_2215,N_2085);
nor U2922 (N_2922,N_2000,N_2122);
nor U2923 (N_2923,N_2278,N_2258);
nand U2924 (N_2924,N_2398,N_2182);
nand U2925 (N_2925,N_2313,N_2074);
xor U2926 (N_2926,N_2199,N_2052);
or U2927 (N_2927,N_2252,N_2467);
and U2928 (N_2928,N_2023,N_2059);
nor U2929 (N_2929,N_2033,N_2228);
nor U2930 (N_2930,N_2063,N_2175);
or U2931 (N_2931,N_2174,N_2224);
and U2932 (N_2932,N_2159,N_2343);
nor U2933 (N_2933,N_2418,N_2342);
nand U2934 (N_2934,N_2079,N_2284);
or U2935 (N_2935,N_2167,N_2168);
nand U2936 (N_2936,N_2485,N_2336);
and U2937 (N_2937,N_2223,N_2149);
and U2938 (N_2938,N_2364,N_2109);
and U2939 (N_2939,N_2204,N_2252);
nand U2940 (N_2940,N_2427,N_2129);
xnor U2941 (N_2941,N_2060,N_2097);
xnor U2942 (N_2942,N_2333,N_2242);
nand U2943 (N_2943,N_2024,N_2131);
nor U2944 (N_2944,N_2181,N_2434);
or U2945 (N_2945,N_2127,N_2180);
and U2946 (N_2946,N_2059,N_2302);
nand U2947 (N_2947,N_2354,N_2034);
nand U2948 (N_2948,N_2020,N_2374);
and U2949 (N_2949,N_2265,N_2349);
or U2950 (N_2950,N_2370,N_2337);
or U2951 (N_2951,N_2370,N_2218);
nor U2952 (N_2952,N_2225,N_2334);
nor U2953 (N_2953,N_2187,N_2497);
and U2954 (N_2954,N_2316,N_2012);
nand U2955 (N_2955,N_2311,N_2460);
nor U2956 (N_2956,N_2175,N_2199);
or U2957 (N_2957,N_2221,N_2447);
nor U2958 (N_2958,N_2312,N_2112);
and U2959 (N_2959,N_2078,N_2053);
nand U2960 (N_2960,N_2314,N_2072);
nor U2961 (N_2961,N_2172,N_2189);
nand U2962 (N_2962,N_2280,N_2037);
or U2963 (N_2963,N_2358,N_2449);
nand U2964 (N_2964,N_2236,N_2488);
nor U2965 (N_2965,N_2081,N_2413);
or U2966 (N_2966,N_2111,N_2408);
nand U2967 (N_2967,N_2357,N_2293);
or U2968 (N_2968,N_2148,N_2143);
nand U2969 (N_2969,N_2459,N_2360);
nand U2970 (N_2970,N_2363,N_2340);
or U2971 (N_2971,N_2135,N_2425);
or U2972 (N_2972,N_2087,N_2366);
nand U2973 (N_2973,N_2189,N_2446);
nor U2974 (N_2974,N_2092,N_2318);
or U2975 (N_2975,N_2197,N_2006);
nor U2976 (N_2976,N_2231,N_2022);
and U2977 (N_2977,N_2176,N_2123);
nor U2978 (N_2978,N_2184,N_2260);
nand U2979 (N_2979,N_2122,N_2349);
or U2980 (N_2980,N_2059,N_2156);
nor U2981 (N_2981,N_2499,N_2364);
nand U2982 (N_2982,N_2381,N_2473);
or U2983 (N_2983,N_2314,N_2309);
nand U2984 (N_2984,N_2097,N_2085);
nand U2985 (N_2985,N_2218,N_2146);
or U2986 (N_2986,N_2378,N_2046);
nand U2987 (N_2987,N_2043,N_2198);
nand U2988 (N_2988,N_2321,N_2452);
or U2989 (N_2989,N_2222,N_2436);
nor U2990 (N_2990,N_2026,N_2446);
nor U2991 (N_2991,N_2341,N_2128);
or U2992 (N_2992,N_2209,N_2460);
nor U2993 (N_2993,N_2049,N_2458);
nor U2994 (N_2994,N_2224,N_2471);
nand U2995 (N_2995,N_2224,N_2373);
nand U2996 (N_2996,N_2103,N_2003);
or U2997 (N_2997,N_2267,N_2017);
or U2998 (N_2998,N_2081,N_2003);
nor U2999 (N_2999,N_2282,N_2334);
nand UO_0 (O_0,N_2992,N_2609);
nor UO_1 (O_1,N_2963,N_2721);
nand UO_2 (O_2,N_2686,N_2675);
and UO_3 (O_3,N_2937,N_2596);
xor UO_4 (O_4,N_2723,N_2667);
or UO_5 (O_5,N_2767,N_2505);
nor UO_6 (O_6,N_2644,N_2769);
and UO_7 (O_7,N_2926,N_2735);
nand UO_8 (O_8,N_2687,N_2717);
and UO_9 (O_9,N_2745,N_2821);
or UO_10 (O_10,N_2594,N_2840);
nor UO_11 (O_11,N_2814,N_2957);
and UO_12 (O_12,N_2872,N_2984);
and UO_13 (O_13,N_2693,N_2981);
nand UO_14 (O_14,N_2697,N_2583);
and UO_15 (O_15,N_2616,N_2944);
or UO_16 (O_16,N_2884,N_2706);
and UO_17 (O_17,N_2638,N_2980);
nor UO_18 (O_18,N_2584,N_2779);
nor UO_19 (O_19,N_2664,N_2913);
nand UO_20 (O_20,N_2783,N_2865);
nand UO_21 (O_21,N_2927,N_2986);
and UO_22 (O_22,N_2990,N_2808);
nor UO_23 (O_23,N_2979,N_2756);
nor UO_24 (O_24,N_2677,N_2772);
or UO_25 (O_25,N_2539,N_2683);
nand UO_26 (O_26,N_2995,N_2829);
nor UO_27 (O_27,N_2806,N_2509);
xnor UO_28 (O_28,N_2588,N_2738);
nand UO_29 (O_29,N_2757,N_2670);
nor UO_30 (O_30,N_2946,N_2819);
nor UO_31 (O_31,N_2850,N_2862);
or UO_32 (O_32,N_2982,N_2917);
nor UO_33 (O_33,N_2999,N_2689);
nand UO_34 (O_34,N_2930,N_2654);
nand UO_35 (O_35,N_2537,N_2655);
nor UO_36 (O_36,N_2665,N_2878);
nand UO_37 (O_37,N_2776,N_2582);
and UO_38 (O_38,N_2501,N_2731);
nor UO_39 (O_39,N_2621,N_2998);
and UO_40 (O_40,N_2650,N_2587);
nand UO_41 (O_41,N_2719,N_2612);
or UO_42 (O_42,N_2837,N_2524);
nor UO_43 (O_43,N_2971,N_2941);
or UO_44 (O_44,N_2606,N_2647);
and UO_45 (O_45,N_2567,N_2754);
or UO_46 (O_46,N_2773,N_2935);
or UO_47 (O_47,N_2768,N_2860);
or UO_48 (O_48,N_2880,N_2764);
or UO_49 (O_49,N_2591,N_2945);
xor UO_50 (O_50,N_2698,N_2578);
or UO_51 (O_51,N_2744,N_2958);
and UO_52 (O_52,N_2901,N_2885);
or UO_53 (O_53,N_2888,N_2737);
or UO_54 (O_54,N_2960,N_2909);
nand UO_55 (O_55,N_2815,N_2568);
or UO_56 (O_56,N_2516,N_2900);
nand UO_57 (O_57,N_2694,N_2752);
nand UO_58 (O_58,N_2922,N_2747);
nor UO_59 (O_59,N_2997,N_2955);
nor UO_60 (O_60,N_2956,N_2845);
and UO_61 (O_61,N_2891,N_2780);
nand UO_62 (O_62,N_2666,N_2912);
nor UO_63 (O_63,N_2874,N_2548);
nand UO_64 (O_64,N_2577,N_2809);
or UO_65 (O_65,N_2939,N_2630);
or UO_66 (O_66,N_2503,N_2640);
nand UO_67 (O_67,N_2691,N_2550);
xnor UO_68 (O_68,N_2519,N_2574);
and UO_69 (O_69,N_2546,N_2728);
nand UO_70 (O_70,N_2763,N_2771);
and UO_71 (O_71,N_2961,N_2620);
or UO_72 (O_72,N_2749,N_2551);
or UO_73 (O_73,N_2634,N_2856);
and UO_74 (O_74,N_2718,N_2972);
or UO_75 (O_75,N_2557,N_2590);
and UO_76 (O_76,N_2828,N_2572);
or UO_77 (O_77,N_2753,N_2879);
nor UO_78 (O_78,N_2528,N_2841);
xnor UO_79 (O_79,N_2940,N_2619);
nand UO_80 (O_80,N_2506,N_2942);
or UO_81 (O_81,N_2983,N_2576);
nand UO_82 (O_82,N_2645,N_2510);
or UO_83 (O_83,N_2766,N_2886);
nand UO_84 (O_84,N_2720,N_2710);
and UO_85 (O_85,N_2925,N_2993);
or UO_86 (O_86,N_2549,N_2529);
nand UO_87 (O_87,N_2920,N_2652);
nor UO_88 (O_88,N_2736,N_2923);
nand UO_89 (O_89,N_2540,N_2857);
or UO_90 (O_90,N_2522,N_2974);
and UO_91 (O_91,N_2797,N_2561);
nand UO_92 (O_92,N_2949,N_2866);
nor UO_93 (O_93,N_2905,N_2989);
or UO_94 (O_94,N_2623,N_2858);
or UO_95 (O_95,N_2595,N_2629);
or UO_96 (O_96,N_2834,N_2605);
nand UO_97 (O_97,N_2727,N_2663);
or UO_98 (O_98,N_2904,N_2504);
and UO_99 (O_99,N_2725,N_2592);
nor UO_100 (O_100,N_2831,N_2690);
or UO_101 (O_101,N_2967,N_2802);
nor UO_102 (O_102,N_2661,N_2870);
nor UO_103 (O_103,N_2931,N_2660);
or UO_104 (O_104,N_2805,N_2914);
nand UO_105 (O_105,N_2867,N_2580);
nor UO_106 (O_106,N_2688,N_2788);
nand UO_107 (O_107,N_2796,N_2807);
or UO_108 (O_108,N_2948,N_2893);
nand UO_109 (O_109,N_2896,N_2599);
nand UO_110 (O_110,N_2545,N_2542);
or UO_111 (O_111,N_2818,N_2607);
nand UO_112 (O_112,N_2649,N_2765);
nand UO_113 (O_113,N_2804,N_2936);
nor UO_114 (O_114,N_2799,N_2921);
nor UO_115 (O_115,N_2603,N_2864);
nor UO_116 (O_116,N_2659,N_2748);
nand UO_117 (O_117,N_2742,N_2916);
and UO_118 (O_118,N_2733,N_2672);
or UO_119 (O_119,N_2934,N_2679);
and UO_120 (O_120,N_2525,N_2556);
nor UO_121 (O_121,N_2810,N_2969);
nand UO_122 (O_122,N_2657,N_2684);
or UO_123 (O_123,N_2502,N_2611);
and UO_124 (O_124,N_2575,N_2873);
nand UO_125 (O_125,N_2787,N_2637);
and UO_126 (O_126,N_2825,N_2844);
nor UO_127 (O_127,N_2598,N_2785);
or UO_128 (O_128,N_2669,N_2615);
and UO_129 (O_129,N_2523,N_2911);
or UO_130 (O_130,N_2680,N_2890);
nor UO_131 (O_131,N_2863,N_2758);
nor UO_132 (O_132,N_2964,N_2579);
or UO_133 (O_133,N_2970,N_2869);
nor UO_134 (O_134,N_2826,N_2947);
nand UO_135 (O_135,N_2518,N_2755);
nor UO_136 (O_136,N_2854,N_2932);
or UO_137 (O_137,N_2976,N_2602);
and UO_138 (O_138,N_2813,N_2521);
nand UO_139 (O_139,N_2653,N_2526);
or UO_140 (O_140,N_2835,N_2762);
and UO_141 (O_141,N_2994,N_2908);
nor UO_142 (O_142,N_2790,N_2950);
nor UO_143 (O_143,N_2954,N_2830);
nand UO_144 (O_144,N_2722,N_2784);
or UO_145 (O_145,N_2585,N_2789);
nor UO_146 (O_146,N_2875,N_2559);
or UO_147 (O_147,N_2538,N_2848);
or UO_148 (O_148,N_2534,N_2739);
nand UO_149 (O_149,N_2743,N_2833);
and UO_150 (O_150,N_2681,N_2730);
nor UO_151 (O_151,N_2631,N_2881);
or UO_152 (O_152,N_2646,N_2651);
nand UO_153 (O_153,N_2715,N_2533);
and UO_154 (O_154,N_2581,N_2760);
and UO_155 (O_155,N_2962,N_2793);
nand UO_156 (O_156,N_2877,N_2702);
nand UO_157 (O_157,N_2641,N_2953);
nand UO_158 (O_158,N_2778,N_2692);
nand UO_159 (O_159,N_2859,N_2622);
nand UO_160 (O_160,N_2968,N_2662);
or UO_161 (O_161,N_2894,N_2625);
nor UO_162 (O_162,N_2987,N_2973);
or UO_163 (O_163,N_2714,N_2648);
and UO_164 (O_164,N_2500,N_2846);
and UO_165 (O_165,N_2696,N_2824);
nor UO_166 (O_166,N_2811,N_2724);
and UO_167 (O_167,N_2823,N_2674);
or UO_168 (O_168,N_2565,N_2713);
or UO_169 (O_169,N_2907,N_2853);
and UO_170 (O_170,N_2673,N_2889);
and UO_171 (O_171,N_2952,N_2560);
nand UO_172 (O_172,N_2531,N_2978);
and UO_173 (O_173,N_2658,N_2635);
and UO_174 (O_174,N_2562,N_2847);
or UO_175 (O_175,N_2801,N_2708);
xnor UO_176 (O_176,N_2803,N_2544);
and UO_177 (O_177,N_2513,N_2820);
nand UO_178 (O_178,N_2601,N_2938);
nor UO_179 (O_179,N_2527,N_2676);
or UO_180 (O_180,N_2751,N_2951);
nor UO_181 (O_181,N_2924,N_2816);
nand UO_182 (O_182,N_2919,N_2943);
nand UO_183 (O_183,N_2558,N_2685);
nor UO_184 (O_184,N_2508,N_2918);
or UO_185 (O_185,N_2903,N_2827);
nor UO_186 (O_186,N_2515,N_2627);
and UO_187 (O_187,N_2897,N_2852);
or UO_188 (O_188,N_2800,N_2741);
and UO_189 (O_189,N_2514,N_2832);
or UO_190 (O_190,N_2928,N_2794);
nor UO_191 (O_191,N_2552,N_2839);
or UO_192 (O_192,N_2732,N_2547);
nand UO_193 (O_193,N_2617,N_2700);
or UO_194 (O_194,N_2775,N_2883);
and UO_195 (O_195,N_2610,N_2705);
xor UO_196 (O_196,N_2608,N_2899);
or UO_197 (O_197,N_2770,N_2991);
or UO_198 (O_198,N_2792,N_2569);
and UO_199 (O_199,N_2618,N_2761);
nand UO_200 (O_200,N_2786,N_2977);
nor UO_201 (O_201,N_2855,N_2633);
nor UO_202 (O_202,N_2929,N_2678);
and UO_203 (O_203,N_2536,N_2517);
or UO_204 (O_204,N_2704,N_2520);
or UO_205 (O_205,N_2632,N_2566);
or UO_206 (O_206,N_2511,N_2750);
nand UO_207 (O_207,N_2682,N_2734);
nor UO_208 (O_208,N_2965,N_2701);
and UO_209 (O_209,N_2712,N_2711);
or UO_210 (O_210,N_2795,N_2791);
and UO_211 (O_211,N_2586,N_2555);
or UO_212 (O_212,N_2975,N_2570);
nand UO_213 (O_213,N_2985,N_2563);
xor UO_214 (O_214,N_2553,N_2861);
nor UO_215 (O_215,N_2571,N_2851);
nand UO_216 (O_216,N_2892,N_2628);
and UO_217 (O_217,N_2774,N_2726);
and UO_218 (O_218,N_2849,N_2671);
or UO_219 (O_219,N_2699,N_2600);
and UO_220 (O_220,N_2996,N_2871);
xor UO_221 (O_221,N_2740,N_2703);
and UO_222 (O_222,N_2882,N_2613);
and UO_223 (O_223,N_2573,N_2642);
nor UO_224 (O_224,N_2593,N_2822);
nand UO_225 (O_225,N_2746,N_2639);
xor UO_226 (O_226,N_2656,N_2507);
and UO_227 (O_227,N_2988,N_2898);
nand UO_228 (O_228,N_2624,N_2695);
or UO_229 (O_229,N_2626,N_2959);
nand UO_230 (O_230,N_2535,N_2716);
and UO_231 (O_231,N_2812,N_2817);
or UO_232 (O_232,N_2543,N_2843);
or UO_233 (O_233,N_2966,N_2777);
nand UO_234 (O_234,N_2643,N_2614);
nor UO_235 (O_235,N_2759,N_2512);
nor UO_236 (O_236,N_2868,N_2707);
and UO_237 (O_237,N_2709,N_2915);
nor UO_238 (O_238,N_2729,N_2541);
nor UO_239 (O_239,N_2589,N_2876);
or UO_240 (O_240,N_2838,N_2902);
and UO_241 (O_241,N_2604,N_2887);
xor UO_242 (O_242,N_2836,N_2906);
nand UO_243 (O_243,N_2564,N_2668);
nand UO_244 (O_244,N_2530,N_2895);
nor UO_245 (O_245,N_2910,N_2842);
nand UO_246 (O_246,N_2532,N_2933);
and UO_247 (O_247,N_2798,N_2554);
or UO_248 (O_248,N_2597,N_2781);
nand UO_249 (O_249,N_2782,N_2636);
or UO_250 (O_250,N_2711,N_2615);
nand UO_251 (O_251,N_2882,N_2818);
nand UO_252 (O_252,N_2954,N_2530);
or UO_253 (O_253,N_2891,N_2786);
and UO_254 (O_254,N_2646,N_2764);
nand UO_255 (O_255,N_2736,N_2714);
nor UO_256 (O_256,N_2754,N_2909);
nand UO_257 (O_257,N_2873,N_2631);
nand UO_258 (O_258,N_2938,N_2553);
nor UO_259 (O_259,N_2922,N_2667);
nor UO_260 (O_260,N_2951,N_2683);
or UO_261 (O_261,N_2903,N_2882);
or UO_262 (O_262,N_2910,N_2771);
or UO_263 (O_263,N_2617,N_2844);
xnor UO_264 (O_264,N_2605,N_2973);
xor UO_265 (O_265,N_2670,N_2639);
nand UO_266 (O_266,N_2996,N_2758);
or UO_267 (O_267,N_2850,N_2643);
and UO_268 (O_268,N_2731,N_2883);
and UO_269 (O_269,N_2974,N_2886);
nand UO_270 (O_270,N_2536,N_2864);
nor UO_271 (O_271,N_2868,N_2983);
nand UO_272 (O_272,N_2617,N_2562);
or UO_273 (O_273,N_2719,N_2645);
nand UO_274 (O_274,N_2763,N_2651);
or UO_275 (O_275,N_2661,N_2784);
nand UO_276 (O_276,N_2608,N_2803);
nor UO_277 (O_277,N_2987,N_2897);
xor UO_278 (O_278,N_2503,N_2952);
nor UO_279 (O_279,N_2532,N_2529);
and UO_280 (O_280,N_2603,N_2744);
xnor UO_281 (O_281,N_2854,N_2642);
nor UO_282 (O_282,N_2926,N_2767);
nor UO_283 (O_283,N_2697,N_2524);
nand UO_284 (O_284,N_2818,N_2511);
and UO_285 (O_285,N_2863,N_2791);
nand UO_286 (O_286,N_2678,N_2826);
and UO_287 (O_287,N_2790,N_2686);
nor UO_288 (O_288,N_2845,N_2564);
nand UO_289 (O_289,N_2581,N_2844);
or UO_290 (O_290,N_2750,N_2974);
or UO_291 (O_291,N_2783,N_2961);
xor UO_292 (O_292,N_2542,N_2661);
nand UO_293 (O_293,N_2849,N_2528);
or UO_294 (O_294,N_2960,N_2875);
or UO_295 (O_295,N_2991,N_2929);
and UO_296 (O_296,N_2590,N_2699);
and UO_297 (O_297,N_2698,N_2838);
nor UO_298 (O_298,N_2832,N_2717);
nor UO_299 (O_299,N_2788,N_2724);
nor UO_300 (O_300,N_2733,N_2847);
and UO_301 (O_301,N_2889,N_2879);
xor UO_302 (O_302,N_2627,N_2544);
or UO_303 (O_303,N_2932,N_2943);
or UO_304 (O_304,N_2941,N_2873);
and UO_305 (O_305,N_2500,N_2711);
and UO_306 (O_306,N_2679,N_2662);
or UO_307 (O_307,N_2979,N_2680);
nand UO_308 (O_308,N_2954,N_2620);
nor UO_309 (O_309,N_2746,N_2742);
nor UO_310 (O_310,N_2912,N_2572);
nor UO_311 (O_311,N_2811,N_2966);
or UO_312 (O_312,N_2803,N_2751);
nand UO_313 (O_313,N_2750,N_2753);
or UO_314 (O_314,N_2710,N_2811);
and UO_315 (O_315,N_2678,N_2607);
or UO_316 (O_316,N_2826,N_2569);
or UO_317 (O_317,N_2576,N_2848);
nand UO_318 (O_318,N_2999,N_2827);
or UO_319 (O_319,N_2750,N_2840);
or UO_320 (O_320,N_2549,N_2612);
or UO_321 (O_321,N_2835,N_2861);
or UO_322 (O_322,N_2949,N_2573);
or UO_323 (O_323,N_2526,N_2765);
nor UO_324 (O_324,N_2624,N_2801);
nor UO_325 (O_325,N_2607,N_2562);
or UO_326 (O_326,N_2672,N_2705);
nand UO_327 (O_327,N_2631,N_2987);
or UO_328 (O_328,N_2765,N_2838);
or UO_329 (O_329,N_2775,N_2990);
or UO_330 (O_330,N_2656,N_2514);
and UO_331 (O_331,N_2920,N_2794);
nand UO_332 (O_332,N_2520,N_2733);
nor UO_333 (O_333,N_2952,N_2937);
or UO_334 (O_334,N_2666,N_2662);
nand UO_335 (O_335,N_2715,N_2950);
and UO_336 (O_336,N_2876,N_2529);
nand UO_337 (O_337,N_2554,N_2804);
nor UO_338 (O_338,N_2675,N_2826);
nor UO_339 (O_339,N_2858,N_2983);
nor UO_340 (O_340,N_2552,N_2863);
nor UO_341 (O_341,N_2591,N_2745);
nand UO_342 (O_342,N_2875,N_2714);
and UO_343 (O_343,N_2741,N_2867);
or UO_344 (O_344,N_2592,N_2515);
or UO_345 (O_345,N_2896,N_2768);
and UO_346 (O_346,N_2848,N_2710);
nor UO_347 (O_347,N_2945,N_2896);
nor UO_348 (O_348,N_2637,N_2525);
nor UO_349 (O_349,N_2579,N_2896);
or UO_350 (O_350,N_2974,N_2852);
nor UO_351 (O_351,N_2990,N_2954);
nand UO_352 (O_352,N_2981,N_2637);
or UO_353 (O_353,N_2845,N_2735);
nor UO_354 (O_354,N_2898,N_2840);
nor UO_355 (O_355,N_2793,N_2771);
and UO_356 (O_356,N_2597,N_2611);
and UO_357 (O_357,N_2810,N_2567);
and UO_358 (O_358,N_2896,N_2862);
and UO_359 (O_359,N_2835,N_2824);
nor UO_360 (O_360,N_2568,N_2644);
nor UO_361 (O_361,N_2562,N_2891);
or UO_362 (O_362,N_2547,N_2726);
nand UO_363 (O_363,N_2502,N_2882);
or UO_364 (O_364,N_2692,N_2649);
or UO_365 (O_365,N_2782,N_2656);
nor UO_366 (O_366,N_2898,N_2958);
and UO_367 (O_367,N_2699,N_2776);
or UO_368 (O_368,N_2659,N_2539);
nand UO_369 (O_369,N_2925,N_2781);
or UO_370 (O_370,N_2755,N_2788);
nand UO_371 (O_371,N_2902,N_2803);
or UO_372 (O_372,N_2899,N_2834);
nor UO_373 (O_373,N_2635,N_2694);
nor UO_374 (O_374,N_2510,N_2876);
nor UO_375 (O_375,N_2729,N_2537);
and UO_376 (O_376,N_2628,N_2651);
and UO_377 (O_377,N_2915,N_2578);
or UO_378 (O_378,N_2749,N_2589);
nor UO_379 (O_379,N_2571,N_2977);
nand UO_380 (O_380,N_2853,N_2517);
nor UO_381 (O_381,N_2501,N_2646);
or UO_382 (O_382,N_2826,N_2610);
and UO_383 (O_383,N_2825,N_2801);
and UO_384 (O_384,N_2917,N_2619);
and UO_385 (O_385,N_2977,N_2998);
and UO_386 (O_386,N_2828,N_2954);
or UO_387 (O_387,N_2562,N_2917);
nand UO_388 (O_388,N_2897,N_2730);
and UO_389 (O_389,N_2600,N_2717);
and UO_390 (O_390,N_2699,N_2815);
nor UO_391 (O_391,N_2897,N_2924);
nor UO_392 (O_392,N_2772,N_2675);
nand UO_393 (O_393,N_2828,N_2610);
and UO_394 (O_394,N_2737,N_2724);
and UO_395 (O_395,N_2591,N_2971);
nor UO_396 (O_396,N_2851,N_2840);
and UO_397 (O_397,N_2701,N_2754);
nand UO_398 (O_398,N_2765,N_2850);
or UO_399 (O_399,N_2987,N_2790);
and UO_400 (O_400,N_2807,N_2536);
nand UO_401 (O_401,N_2661,N_2928);
nand UO_402 (O_402,N_2975,N_2680);
and UO_403 (O_403,N_2675,N_2562);
nand UO_404 (O_404,N_2764,N_2672);
or UO_405 (O_405,N_2753,N_2788);
or UO_406 (O_406,N_2772,N_2999);
nand UO_407 (O_407,N_2534,N_2553);
nand UO_408 (O_408,N_2623,N_2544);
or UO_409 (O_409,N_2972,N_2768);
nand UO_410 (O_410,N_2779,N_2762);
or UO_411 (O_411,N_2684,N_2870);
nand UO_412 (O_412,N_2954,N_2952);
nand UO_413 (O_413,N_2849,N_2737);
and UO_414 (O_414,N_2508,N_2542);
and UO_415 (O_415,N_2616,N_2852);
nor UO_416 (O_416,N_2837,N_2521);
and UO_417 (O_417,N_2779,N_2980);
nor UO_418 (O_418,N_2697,N_2981);
nand UO_419 (O_419,N_2954,N_2801);
and UO_420 (O_420,N_2577,N_2673);
and UO_421 (O_421,N_2538,N_2944);
or UO_422 (O_422,N_2745,N_2768);
nor UO_423 (O_423,N_2869,N_2851);
xor UO_424 (O_424,N_2907,N_2905);
nand UO_425 (O_425,N_2522,N_2566);
and UO_426 (O_426,N_2974,N_2726);
nand UO_427 (O_427,N_2828,N_2767);
or UO_428 (O_428,N_2814,N_2714);
nand UO_429 (O_429,N_2984,N_2996);
and UO_430 (O_430,N_2693,N_2970);
and UO_431 (O_431,N_2978,N_2770);
and UO_432 (O_432,N_2542,N_2907);
nor UO_433 (O_433,N_2940,N_2988);
nor UO_434 (O_434,N_2943,N_2951);
nor UO_435 (O_435,N_2586,N_2972);
or UO_436 (O_436,N_2687,N_2813);
and UO_437 (O_437,N_2748,N_2902);
nor UO_438 (O_438,N_2806,N_2670);
or UO_439 (O_439,N_2553,N_2822);
or UO_440 (O_440,N_2680,N_2796);
nor UO_441 (O_441,N_2640,N_2993);
and UO_442 (O_442,N_2756,N_2723);
nand UO_443 (O_443,N_2669,N_2591);
nand UO_444 (O_444,N_2843,N_2842);
nor UO_445 (O_445,N_2545,N_2649);
or UO_446 (O_446,N_2730,N_2555);
nor UO_447 (O_447,N_2558,N_2659);
or UO_448 (O_448,N_2587,N_2847);
or UO_449 (O_449,N_2528,N_2754);
or UO_450 (O_450,N_2942,N_2800);
nand UO_451 (O_451,N_2571,N_2593);
or UO_452 (O_452,N_2509,N_2894);
xnor UO_453 (O_453,N_2987,N_2554);
nor UO_454 (O_454,N_2738,N_2948);
or UO_455 (O_455,N_2810,N_2839);
xnor UO_456 (O_456,N_2692,N_2887);
nand UO_457 (O_457,N_2787,N_2811);
nor UO_458 (O_458,N_2533,N_2831);
or UO_459 (O_459,N_2865,N_2565);
nand UO_460 (O_460,N_2990,N_2714);
nand UO_461 (O_461,N_2789,N_2862);
and UO_462 (O_462,N_2581,N_2947);
nor UO_463 (O_463,N_2664,N_2955);
nor UO_464 (O_464,N_2707,N_2642);
or UO_465 (O_465,N_2646,N_2589);
nor UO_466 (O_466,N_2862,N_2561);
or UO_467 (O_467,N_2655,N_2913);
or UO_468 (O_468,N_2697,N_2933);
or UO_469 (O_469,N_2764,N_2884);
or UO_470 (O_470,N_2699,N_2936);
and UO_471 (O_471,N_2733,N_2820);
or UO_472 (O_472,N_2741,N_2913);
nor UO_473 (O_473,N_2938,N_2587);
or UO_474 (O_474,N_2967,N_2637);
and UO_475 (O_475,N_2579,N_2689);
nor UO_476 (O_476,N_2973,N_2594);
xnor UO_477 (O_477,N_2769,N_2909);
and UO_478 (O_478,N_2687,N_2973);
and UO_479 (O_479,N_2832,N_2566);
nand UO_480 (O_480,N_2605,N_2756);
or UO_481 (O_481,N_2714,N_2909);
and UO_482 (O_482,N_2712,N_2607);
nor UO_483 (O_483,N_2645,N_2671);
and UO_484 (O_484,N_2850,N_2726);
nor UO_485 (O_485,N_2998,N_2893);
nor UO_486 (O_486,N_2585,N_2782);
nand UO_487 (O_487,N_2913,N_2687);
or UO_488 (O_488,N_2659,N_2968);
and UO_489 (O_489,N_2671,N_2825);
nor UO_490 (O_490,N_2598,N_2740);
or UO_491 (O_491,N_2691,N_2653);
or UO_492 (O_492,N_2619,N_2508);
or UO_493 (O_493,N_2952,N_2639);
nor UO_494 (O_494,N_2908,N_2903);
nor UO_495 (O_495,N_2872,N_2768);
nand UO_496 (O_496,N_2979,N_2671);
nand UO_497 (O_497,N_2773,N_2836);
nand UO_498 (O_498,N_2743,N_2529);
and UO_499 (O_499,N_2513,N_2677);
endmodule