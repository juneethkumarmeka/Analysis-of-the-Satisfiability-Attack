module basic_5000_50000_5000_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_4007,In_865);
nor U1 (N_1,In_36,In_2315);
or U2 (N_2,In_4507,In_2616);
xnor U3 (N_3,In_706,In_4177);
nand U4 (N_4,In_2849,In_2542);
nand U5 (N_5,In_1407,In_2322);
nor U6 (N_6,In_2247,In_3422);
xnor U7 (N_7,In_4046,In_4040);
nand U8 (N_8,In_2957,In_4472);
nor U9 (N_9,In_3513,In_4923);
and U10 (N_10,In_392,In_768);
or U11 (N_11,In_3267,In_3723);
or U12 (N_12,In_4903,In_3197);
or U13 (N_13,In_181,In_2496);
or U14 (N_14,In_973,In_149);
or U15 (N_15,In_1577,In_778);
nor U16 (N_16,In_2044,In_2975);
nor U17 (N_17,In_1143,In_1463);
nand U18 (N_18,In_296,In_3432);
or U19 (N_19,In_2767,In_665);
nand U20 (N_20,In_2652,In_2833);
and U21 (N_21,In_2532,In_4250);
nand U22 (N_22,In_2318,In_4152);
nor U23 (N_23,In_4257,In_4092);
xor U24 (N_24,In_2225,In_3932);
xnor U25 (N_25,In_1371,In_1097);
or U26 (N_26,In_4188,In_4605);
nand U27 (N_27,In_1446,In_1759);
nand U28 (N_28,In_984,In_2875);
nand U29 (N_29,In_1746,In_2677);
or U30 (N_30,In_2450,In_1808);
and U31 (N_31,In_1422,In_1164);
or U32 (N_32,In_2148,In_2891);
xor U33 (N_33,In_1559,In_560);
or U34 (N_34,In_2104,In_2385);
or U35 (N_35,In_1743,In_1615);
nand U36 (N_36,In_4198,In_3185);
nand U37 (N_37,In_1256,In_3878);
and U38 (N_38,In_3320,In_564);
and U39 (N_39,In_1061,In_1079);
nand U40 (N_40,In_2224,In_1169);
and U41 (N_41,In_607,In_2343);
or U42 (N_42,In_4506,In_4193);
nand U43 (N_43,In_525,In_4110);
nand U44 (N_44,In_4947,In_1089);
nand U45 (N_45,In_4070,In_4163);
and U46 (N_46,In_4900,In_4212);
and U47 (N_47,In_3011,In_3374);
nand U48 (N_48,In_1728,In_3092);
xor U49 (N_49,In_644,In_4864);
or U50 (N_50,In_801,In_2910);
and U51 (N_51,In_3879,In_2111);
nand U52 (N_52,In_3576,In_1328);
nand U53 (N_53,In_4622,In_2527);
and U54 (N_54,In_2878,In_4379);
or U55 (N_55,In_692,In_3844);
nand U56 (N_56,In_545,In_1600);
xor U57 (N_57,In_2831,In_3045);
nor U58 (N_58,In_4448,In_68);
and U59 (N_59,In_566,In_854);
nor U60 (N_60,In_1483,In_1421);
and U61 (N_61,In_1306,In_4464);
and U62 (N_62,In_1846,In_1500);
and U63 (N_63,In_4280,In_2331);
xor U64 (N_64,In_4461,In_3999);
or U65 (N_65,In_3025,In_1788);
nor U66 (N_66,In_3854,In_2627);
or U67 (N_67,In_4319,In_2893);
and U68 (N_68,In_1354,In_914);
and U69 (N_69,In_4227,In_111);
and U70 (N_70,In_659,In_1823);
and U71 (N_71,In_4905,In_1845);
or U72 (N_72,In_1327,In_2010);
nand U73 (N_73,In_4490,In_2839);
or U74 (N_74,In_1382,In_1054);
or U75 (N_75,In_2869,In_1213);
and U76 (N_76,In_871,In_572);
and U77 (N_77,In_3221,In_1758);
and U78 (N_78,In_457,In_1198);
and U79 (N_79,In_4732,In_1637);
or U80 (N_80,In_2801,In_3481);
xnor U81 (N_81,In_4997,In_4946);
nand U82 (N_82,In_959,In_3289);
nand U83 (N_83,In_4413,In_2358);
and U84 (N_84,In_342,In_329);
nand U85 (N_85,In_4189,In_1031);
xnor U86 (N_86,In_265,In_2584);
xor U87 (N_87,In_1283,In_4321);
nor U88 (N_88,In_4024,In_215);
xnor U89 (N_89,In_2077,In_3590);
and U90 (N_90,In_2959,In_1598);
nand U91 (N_91,In_2942,In_1580);
nand U92 (N_92,In_3687,In_4801);
xnor U93 (N_93,In_2775,In_1452);
nor U94 (N_94,In_2666,In_4361);
xnor U95 (N_95,In_2887,In_2582);
xnor U96 (N_96,In_2492,In_4534);
or U97 (N_97,In_2459,In_1990);
xor U98 (N_98,In_1352,In_3913);
or U99 (N_99,In_202,In_1609);
nand U100 (N_100,In_4840,In_1958);
nor U101 (N_101,In_77,In_509);
nand U102 (N_102,In_2033,In_637);
nand U103 (N_103,In_2489,In_4333);
or U104 (N_104,In_1875,In_3961);
nor U105 (N_105,In_172,In_2463);
xnor U106 (N_106,In_1032,In_4150);
nand U107 (N_107,In_1247,In_4038);
nand U108 (N_108,In_1429,In_398);
xor U109 (N_109,In_4744,In_4045);
nor U110 (N_110,In_755,In_3997);
nor U111 (N_111,In_3690,In_2451);
nor U112 (N_112,In_482,In_4465);
nand U113 (N_113,In_1066,In_4255);
nand U114 (N_114,In_4484,In_4010);
or U115 (N_115,In_1204,In_3281);
or U116 (N_116,In_1961,In_1632);
nor U117 (N_117,In_4775,In_3433);
and U118 (N_118,In_2600,In_1687);
nor U119 (N_119,In_146,In_1779);
and U120 (N_120,In_3872,In_3528);
nor U121 (N_121,In_4301,In_4228);
or U122 (N_122,In_4182,In_4850);
nand U123 (N_123,In_688,In_4416);
and U124 (N_124,In_936,In_1850);
xnor U125 (N_125,In_294,In_1832);
nor U126 (N_126,In_1474,In_5);
nor U127 (N_127,In_3215,In_3988);
nor U128 (N_128,In_3660,In_4354);
nor U129 (N_129,In_1602,In_2609);
and U130 (N_130,In_428,In_4305);
nor U131 (N_131,In_2798,In_1172);
or U132 (N_132,In_2954,In_738);
or U133 (N_133,In_910,In_3656);
and U134 (N_134,In_4501,In_3860);
and U135 (N_135,In_127,In_3019);
nor U136 (N_136,In_4517,In_95);
nor U137 (N_137,In_3897,In_3337);
nand U138 (N_138,In_3689,In_2591);
or U139 (N_139,In_2231,In_4794);
and U140 (N_140,In_3369,In_1005);
or U141 (N_141,In_2311,In_460);
nor U142 (N_142,In_3884,In_1585);
nand U143 (N_143,In_930,In_255);
xnor U144 (N_144,In_1806,In_2997);
nand U145 (N_145,In_810,In_2294);
or U146 (N_146,In_776,In_3220);
or U147 (N_147,In_3,In_3001);
nand U148 (N_148,In_1425,In_1925);
nor U149 (N_149,In_1595,In_427);
and U150 (N_150,In_3269,In_2137);
nor U151 (N_151,In_4600,In_4433);
or U152 (N_152,In_2120,In_2785);
or U153 (N_153,In_130,In_2818);
nor U154 (N_154,In_4486,In_3066);
nor U155 (N_155,In_282,In_2503);
and U156 (N_156,In_4899,In_3174);
nor U157 (N_157,In_947,In_2668);
or U158 (N_158,In_3040,In_839);
nor U159 (N_159,In_4398,In_2288);
xnor U160 (N_160,In_1071,In_4446);
nor U161 (N_161,In_1836,In_4214);
nand U162 (N_162,In_2632,In_2301);
nor U163 (N_163,In_4488,In_4951);
nor U164 (N_164,In_3128,In_3798);
or U165 (N_165,In_3126,In_132);
nor U166 (N_166,In_4555,In_4356);
nor U167 (N_167,In_4706,In_2351);
nor U168 (N_168,In_2170,In_3136);
nand U169 (N_169,In_4930,In_4295);
nand U170 (N_170,In_2447,In_4241);
and U171 (N_171,In_4693,In_2919);
xnor U172 (N_172,In_3072,In_2825);
nand U173 (N_173,In_1130,In_2475);
xor U174 (N_174,In_220,In_3495);
and U175 (N_175,In_4877,In_2992);
nand U176 (N_176,In_4013,In_3627);
xnor U177 (N_177,In_4273,In_1922);
and U178 (N_178,In_2226,In_1184);
or U179 (N_179,In_1424,In_927);
and U180 (N_180,In_860,In_842);
and U181 (N_181,In_3606,In_4828);
or U182 (N_182,In_2158,In_1509);
and U183 (N_183,In_1868,In_2750);
and U184 (N_184,In_987,In_901);
nand U185 (N_185,In_2398,In_1178);
xnor U186 (N_186,In_1106,In_1085);
nand U187 (N_187,In_1488,In_3377);
or U188 (N_188,In_1335,In_3679);
and U189 (N_189,In_832,In_3052);
nand U190 (N_190,In_1332,In_2961);
or U191 (N_191,In_4317,In_1299);
xnor U192 (N_192,In_2483,In_195);
xor U193 (N_193,In_4130,In_2530);
xnor U194 (N_194,In_4759,In_3848);
or U195 (N_195,In_4875,In_2159);
nor U196 (N_196,In_430,In_3863);
nor U197 (N_197,In_1197,In_2424);
nor U198 (N_198,In_4406,In_4719);
nand U199 (N_199,In_1456,In_3112);
or U200 (N_200,In_2222,In_2643);
xor U201 (N_201,In_1158,In_1271);
nand U202 (N_202,In_4672,In_4051);
xor U203 (N_203,In_1928,In_1040);
nand U204 (N_204,In_4965,In_1828);
or U205 (N_205,In_4290,In_4624);
nor U206 (N_206,In_231,In_2131);
and U207 (N_207,In_3584,In_948);
or U208 (N_208,In_1926,In_245);
nand U209 (N_209,In_2661,In_1529);
and U210 (N_210,In_3789,In_3657);
nor U211 (N_211,In_384,In_2876);
or U212 (N_212,In_1028,In_870);
nor U213 (N_213,In_1343,In_1813);
or U214 (N_214,In_4680,In_2040);
nor U215 (N_215,In_438,In_4683);
xor U216 (N_216,In_4279,In_102);
or U217 (N_217,In_3504,In_4608);
nor U218 (N_218,In_2977,In_3399);
or U219 (N_219,In_451,In_287);
xnor U220 (N_220,In_1947,In_4405);
nor U221 (N_221,In_615,In_3993);
or U222 (N_222,In_1975,In_4854);
nand U223 (N_223,In_3198,In_884);
or U224 (N_224,In_4566,In_1716);
nor U225 (N_225,In_1692,In_2710);
nand U226 (N_226,In_3016,In_1113);
and U227 (N_227,In_4039,In_4169);
nor U228 (N_228,In_1882,In_3697);
nand U229 (N_229,In_4986,In_1860);
nor U230 (N_230,In_2923,In_40);
nand U231 (N_231,In_2518,In_3230);
and U232 (N_232,In_426,In_455);
nand U233 (N_233,In_1165,In_266);
and U234 (N_234,In_903,In_1901);
xnor U235 (N_235,In_3845,In_1511);
and U236 (N_236,In_2096,In_2468);
and U237 (N_237,In_3043,In_4787);
xnor U238 (N_238,In_3039,In_1963);
and U239 (N_239,In_3796,In_4991);
and U240 (N_240,In_4300,In_2127);
nor U241 (N_241,In_2610,In_4573);
and U242 (N_242,In_1399,In_4190);
and U243 (N_243,In_198,In_4422);
nand U244 (N_244,In_1155,In_4473);
and U245 (N_245,In_4862,In_4889);
and U246 (N_246,In_791,In_3573);
xnor U247 (N_247,In_4952,In_4498);
nand U248 (N_248,In_813,In_1401);
nor U249 (N_249,In_544,In_4171);
or U250 (N_250,In_3818,In_4286);
or U251 (N_251,In_4563,In_2336);
xnor U252 (N_252,In_1516,In_210);
xor U253 (N_253,In_517,In_1237);
xnor U254 (N_254,In_3775,In_4391);
and U255 (N_255,In_749,In_370);
or U256 (N_256,In_2707,In_4147);
nor U257 (N_257,In_3014,In_823);
nand U258 (N_258,In_1621,In_4876);
xor U259 (N_259,In_3836,In_4987);
nor U260 (N_260,In_4209,In_513);
and U261 (N_261,In_2725,In_2570);
or U262 (N_262,In_489,In_3060);
and U263 (N_263,In_1867,In_3133);
nor U264 (N_264,In_3375,In_642);
xor U265 (N_265,In_916,In_2602);
xor U266 (N_266,In_4599,In_1611);
nor U267 (N_267,In_1026,In_3499);
nand U268 (N_268,In_4996,In_4256);
or U269 (N_269,In_4972,In_3241);
nor U270 (N_270,In_1334,In_840);
nor U271 (N_271,In_4251,In_1274);
or U272 (N_272,In_4106,In_2441);
or U273 (N_273,In_4418,In_4577);
nand U274 (N_274,In_3274,In_1392);
xnor U275 (N_275,In_1517,In_2233);
or U276 (N_276,In_2917,In_2230);
and U277 (N_277,In_2114,In_3955);
nand U278 (N_278,In_2426,In_3936);
and U279 (N_279,In_596,In_1586);
nand U280 (N_280,In_777,In_1000);
and U281 (N_281,In_3239,In_3098);
or U282 (N_282,In_1210,In_1396);
nor U283 (N_283,In_1034,In_4127);
or U284 (N_284,In_2282,In_4205);
xnor U285 (N_285,In_598,In_1329);
or U286 (N_286,In_4841,In_3880);
nand U287 (N_287,In_2238,In_3079);
xnor U288 (N_288,In_2009,In_1489);
xnor U289 (N_289,In_4340,In_9);
and U290 (N_290,In_4885,In_4457);
or U291 (N_291,In_4469,In_3090);
xnor U292 (N_292,In_15,In_2372);
or U293 (N_293,In_4648,In_4913);
or U294 (N_294,In_1398,In_3950);
nor U295 (N_295,In_2299,In_2332);
nand U296 (N_296,In_1643,In_710);
or U297 (N_297,In_1709,In_4908);
or U298 (N_298,In_879,In_4896);
nor U299 (N_299,In_2458,In_1555);
and U300 (N_300,In_1154,In_1839);
nand U301 (N_301,In_3329,In_2605);
nor U302 (N_302,In_238,In_1578);
and U303 (N_303,In_3982,In_2759);
nor U304 (N_304,In_2354,In_4204);
nor U305 (N_305,In_2041,In_2547);
nor U306 (N_306,In_782,In_485);
and U307 (N_307,In_444,In_635);
nor U308 (N_308,In_2442,In_2142);
nor U309 (N_309,In_1261,In_2173);
and U310 (N_310,In_1704,In_2440);
and U311 (N_311,In_145,In_2933);
nor U312 (N_312,In_4065,In_3813);
and U313 (N_313,In_170,In_4613);
or U314 (N_314,In_2268,In_1182);
nor U315 (N_315,In_2918,In_4494);
and U316 (N_316,In_887,In_22);
xnor U317 (N_317,In_2550,In_2007);
nor U318 (N_318,In_1152,In_3986);
nor U319 (N_319,In_14,In_4940);
xnor U320 (N_320,In_1804,In_4967);
nand U321 (N_321,In_522,In_3334);
or U322 (N_322,In_974,In_403);
xor U323 (N_323,In_1757,In_1902);
or U324 (N_324,In_54,In_2378);
and U325 (N_325,In_3028,In_2204);
and U326 (N_326,In_1739,In_4958);
or U327 (N_327,In_322,In_4466);
and U328 (N_328,In_4233,In_1742);
and U329 (N_329,In_2514,In_4649);
xnor U330 (N_330,In_1008,In_3492);
and U331 (N_331,In_4492,In_174);
or U332 (N_332,In_1263,In_3317);
xnor U333 (N_333,In_1098,In_3871);
xor U334 (N_334,In_4692,In_4890);
or U335 (N_335,In_1272,In_1486);
nor U336 (N_336,In_4268,In_3827);
and U337 (N_337,In_703,In_4096);
nand U338 (N_338,In_4332,In_4539);
xor U339 (N_339,In_3242,In_1729);
or U340 (N_340,In_1367,In_3084);
nor U341 (N_341,In_2344,In_1118);
xnor U342 (N_342,In_1862,In_1219);
xnor U343 (N_343,In_781,In_3340);
nand U344 (N_344,In_2912,In_1645);
xor U345 (N_345,In_4660,In_254);
or U346 (N_346,In_3757,In_2218);
and U347 (N_347,In_961,In_2296);
nor U348 (N_348,In_2903,In_331);
nand U349 (N_349,In_3109,In_3059);
nand U350 (N_350,In_2774,In_2108);
nor U351 (N_351,In_3471,In_4653);
nand U352 (N_352,In_233,In_3416);
xor U353 (N_353,In_4170,In_2967);
nor U354 (N_354,In_783,In_1858);
nand U355 (N_355,In_2200,In_2117);
nand U356 (N_356,In_3453,In_1464);
or U357 (N_357,In_2254,In_4859);
xor U358 (N_358,In_2464,In_1968);
xor U359 (N_359,In_1468,In_695);
xnor U360 (N_360,In_3135,In_4387);
and U361 (N_361,In_4695,In_4629);
xor U362 (N_362,In_3105,In_135);
xnor U363 (N_363,In_388,In_625);
nand U364 (N_364,In_2884,In_277);
or U365 (N_365,In_4310,In_3386);
nor U366 (N_366,In_516,In_1535);
and U367 (N_367,In_704,In_3167);
and U368 (N_368,In_98,In_2481);
or U369 (N_369,In_2068,In_2312);
or U370 (N_370,In_3296,In_4725);
or U371 (N_371,In_1833,In_970);
and U372 (N_372,In_4620,In_846);
and U373 (N_373,In_2211,In_1548);
xnor U374 (N_374,In_1871,In_2913);
nor U375 (N_375,In_4554,In_1979);
xor U376 (N_376,In_4617,In_3976);
nand U377 (N_377,In_3265,In_3791);
or U378 (N_378,In_2676,In_3862);
xnor U379 (N_379,In_2597,In_476);
nand U380 (N_380,In_733,In_3930);
or U381 (N_381,In_66,In_2045);
or U382 (N_382,In_675,In_4338);
or U383 (N_383,In_1762,In_1104);
nand U384 (N_384,In_1503,In_4012);
or U385 (N_385,In_709,In_1207);
and U386 (N_386,In_4119,In_4852);
nor U387 (N_387,In_662,In_3632);
or U388 (N_388,In_942,In_37);
nor U389 (N_389,In_4666,In_4078);
and U390 (N_390,In_956,In_2726);
and U391 (N_391,In_4380,In_1647);
nand U392 (N_392,In_655,In_2216);
or U393 (N_393,In_492,In_1674);
and U394 (N_394,In_2032,In_4861);
and U395 (N_395,In_2874,In_50);
xor U396 (N_396,In_3543,In_4528);
and U397 (N_397,In_1810,In_3217);
nand U398 (N_398,In_4746,In_4519);
nand U399 (N_399,In_3933,In_2566);
or U400 (N_400,In_3285,In_1437);
nand U401 (N_401,In_2840,In_1007);
nor U402 (N_402,In_99,In_1983);
and U403 (N_403,In_4602,In_3083);
xor U404 (N_404,In_4008,In_1619);
nor U405 (N_405,In_1605,In_3366);
xnor U406 (N_406,In_327,In_3168);
nand U407 (N_407,In_2403,In_2501);
nor U408 (N_408,In_4830,In_311);
nor U409 (N_409,In_1091,In_1235);
and U410 (N_410,In_4242,In_2136);
nor U411 (N_411,In_977,In_124);
and U412 (N_412,In_3462,In_4067);
nand U413 (N_413,In_2916,In_1);
or U414 (N_414,In_3892,In_4057);
and U415 (N_415,In_1218,In_2485);
or U416 (N_416,In_1147,In_3355);
and U417 (N_417,In_3315,In_3900);
or U418 (N_418,In_4284,In_589);
nand U419 (N_419,In_4638,In_2210);
nand U420 (N_420,In_339,In_3390);
and U421 (N_421,In_1812,In_3521);
nor U422 (N_422,In_4703,In_279);
or U423 (N_423,In_1403,In_1183);
xnor U424 (N_424,In_4056,In_3391);
xnor U425 (N_425,In_2388,In_1059);
xnor U426 (N_426,In_767,In_3373);
xnor U427 (N_427,In_4195,In_163);
and U428 (N_428,In_2494,In_3461);
and U429 (N_429,In_1814,In_4542);
nand U430 (N_430,In_2162,In_886);
xnor U431 (N_431,In_1162,In_4640);
xnor U432 (N_432,In_850,In_4705);
nor U433 (N_433,In_4834,In_1607);
xnor U434 (N_434,In_4781,In_536);
or U435 (N_435,In_1805,In_4961);
nor U436 (N_436,In_3938,In_104);
nor U437 (N_437,In_3186,In_4825);
xor U438 (N_438,In_2411,In_483);
xor U439 (N_439,In_2928,In_4087);
and U440 (N_440,In_4770,In_2686);
nor U441 (N_441,In_1221,In_2734);
nor U442 (N_442,In_4676,In_657);
or U443 (N_443,In_1043,In_4687);
xnor U444 (N_444,In_212,In_2327);
nor U445 (N_445,In_2963,In_2964);
or U446 (N_446,In_4589,In_2988);
nor U447 (N_447,In_4607,In_17);
xnor U448 (N_448,In_4259,In_1683);
nand U449 (N_449,In_118,In_1231);
nand U450 (N_450,In_2085,In_2456);
nor U451 (N_451,In_3866,In_1859);
and U452 (N_452,In_2663,In_570);
nor U453 (N_453,In_844,In_4202);
nor U454 (N_454,In_373,In_2662);
or U455 (N_455,In_3536,In_439);
or U456 (N_456,In_2735,In_2938);
nand U457 (N_457,In_4580,In_115);
nor U458 (N_458,In_3063,In_629);
and U459 (N_459,In_1259,In_1712);
or U460 (N_460,In_2578,In_1795);
nand U461 (N_461,In_1127,In_2821);
xnor U462 (N_462,In_87,In_414);
and U463 (N_463,In_769,In_1853);
xor U464 (N_464,In_1929,In_3099);
nand U465 (N_465,In_18,In_4757);
nor U466 (N_466,In_1870,In_3987);
nor U467 (N_467,In_2573,In_1505);
xnor U468 (N_468,In_3520,In_3407);
and U469 (N_469,In_2708,In_4026);
nand U470 (N_470,In_784,In_3605);
nor U471 (N_471,In_3840,In_3563);
and U472 (N_472,In_2274,In_4655);
nand U473 (N_473,In_200,In_2395);
xnor U474 (N_474,In_4503,In_2554);
nand U475 (N_475,In_4281,In_1439);
nor U476 (N_476,In_3677,In_1051);
nand U477 (N_477,In_196,In_1393);
and U478 (N_478,In_2581,In_2647);
or U479 (N_479,In_3895,In_2792);
and U480 (N_480,In_383,In_2860);
xnor U481 (N_481,In_1270,In_4218);
nand U482 (N_482,In_3140,In_1648);
or U483 (N_483,In_3851,In_173);
nand U484 (N_484,In_2352,In_3608);
nor U485 (N_485,In_4557,In_3952);
or U486 (N_486,In_1078,In_134);
or U487 (N_487,In_3142,In_240);
nand U488 (N_488,In_4254,In_4055);
nor U489 (N_489,In_1669,In_2989);
or U490 (N_490,In_3405,In_933);
and U491 (N_491,In_4715,In_2285);
xnor U492 (N_492,In_2665,In_4033);
xor U493 (N_493,In_4062,In_4107);
or U494 (N_494,In_330,In_3778);
or U495 (N_495,In_2653,In_4451);
and U496 (N_496,In_1727,In_774);
nand U497 (N_497,In_3323,In_4061);
nor U498 (N_498,In_3947,In_4347);
and U499 (N_499,In_2264,In_1948);
or U500 (N_500,In_458,In_3360);
xor U501 (N_501,In_1864,In_1443);
or U502 (N_502,In_1388,In_3282);
nand U503 (N_503,In_4000,In_318);
and U504 (N_504,In_1524,In_3061);
nand U505 (N_505,In_4266,In_2405);
nor U506 (N_506,In_1995,In_401);
or U507 (N_507,In_3876,In_4704);
xor U508 (N_508,In_1056,In_1462);
or U509 (N_509,In_1432,In_4924);
nor U510 (N_510,In_790,In_3469);
nor U511 (N_511,In_2425,In_154);
nand U512 (N_512,In_3152,In_3246);
and U513 (N_513,In_909,In_2232);
or U514 (N_514,In_3946,In_1735);
or U515 (N_515,In_872,In_3021);
and U516 (N_516,In_168,In_4582);
nand U517 (N_517,In_1175,In_3922);
xnor U518 (N_518,In_236,In_912);
and U519 (N_519,In_736,In_3137);
nand U520 (N_520,In_845,In_1916);
or U521 (N_521,In_4808,In_94);
nand U522 (N_522,In_2531,In_2816);
and U523 (N_523,In_290,In_4977);
nand U524 (N_524,In_286,In_2644);
and U525 (N_525,In_216,In_4271);
nand U526 (N_526,In_503,In_4785);
and U527 (N_527,In_4341,In_3078);
xnor U528 (N_528,In_1955,In_1374);
and U529 (N_529,In_2754,In_4264);
xor U530 (N_530,In_4025,In_1826);
xnor U531 (N_531,In_1939,In_4741);
and U532 (N_532,In_1016,In_4523);
xnor U533 (N_533,In_1453,In_2687);
nor U534 (N_534,In_257,In_1738);
nor U535 (N_535,In_291,In_3149);
nand U536 (N_536,In_1601,In_4291);
and U537 (N_537,In_2400,In_2850);
nor U538 (N_538,In_4041,In_3344);
and U539 (N_539,In_3760,In_2191);
nand U540 (N_540,In_3224,In_2585);
nand U541 (N_541,In_1417,In_1921);
nand U542 (N_542,In_4088,In_3120);
nor U543 (N_543,In_4407,In_1288);
and U544 (N_544,In_159,In_2900);
nand U545 (N_545,In_199,In_3834);
nand U546 (N_546,In_3297,In_1081);
or U547 (N_547,In_4588,In_1659);
and U548 (N_548,In_1321,In_4176);
nor U549 (N_549,In_369,In_4532);
nand U550 (N_550,In_1167,In_1360);
and U551 (N_551,In_371,In_2076);
nor U552 (N_552,In_234,In_1369);
xnor U553 (N_553,In_3254,In_4186);
nand U554 (N_554,In_4630,In_2383);
and U555 (N_555,In_2046,In_2269);
xnor U556 (N_556,In_1530,In_93);
or U557 (N_557,In_4316,In_1946);
nand U558 (N_558,In_2556,In_530);
nand U559 (N_559,In_3474,In_1513);
xor U560 (N_560,In_3284,In_1465);
or U561 (N_561,In_417,In_3972);
or U562 (N_562,In_1531,In_1625);
or U563 (N_563,In_3227,In_1294);
or U564 (N_564,In_4358,In_979);
xnor U565 (N_565,In_698,In_1905);
nand U566 (N_566,In_1831,In_1494);
nand U567 (N_567,In_2365,In_2145);
and U568 (N_568,In_1656,In_568);
nor U569 (N_569,In_3219,In_3935);
or U570 (N_570,In_4904,In_529);
xnor U571 (N_571,In_1298,In_2439);
and U572 (N_572,In_1697,In_3645);
nor U573 (N_573,In_506,In_1628);
nand U574 (N_574,In_2854,In_1404);
xnor U575 (N_575,In_469,In_1707);
xor U576 (N_576,In_1668,In_4627);
xnor U577 (N_577,In_4783,In_2024);
nand U578 (N_578,In_794,In_4917);
nand U579 (N_579,In_2128,In_907);
nor U580 (N_580,In_2746,In_2345);
or U581 (N_581,In_1942,In_3569);
xnor U582 (N_582,In_1286,In_3953);
nor U583 (N_583,In_1088,In_3073);
xnor U584 (N_584,In_2067,In_4443);
nand U585 (N_585,In_1222,In_4482);
nor U586 (N_586,In_3214,In_3434);
nand U587 (N_587,In_3853,In_4945);
nor U588 (N_588,In_2449,In_4644);
and U589 (N_589,In_3904,In_2683);
nand U590 (N_590,In_142,In_3510);
xnor U591 (N_591,In_4248,In_2946);
nor U592 (N_592,In_184,In_207);
xnor U593 (N_593,In_4837,In_4593);
nor U594 (N_594,In_344,In_4094);
xnor U595 (N_595,In_1326,In_4718);
and U596 (N_596,In_3561,In_3050);
xnor U597 (N_597,In_1851,In_4276);
nor U598 (N_598,In_53,In_955);
nor U599 (N_599,In_668,In_1394);
and U600 (N_600,In_326,In_164);
or U601 (N_601,In_672,In_1243);
nand U602 (N_602,In_3957,In_280);
xor U603 (N_603,In_2969,In_4386);
xor U604 (N_604,In_1514,In_2023);
nand U605 (N_605,In_4385,In_3577);
xor U606 (N_606,In_2940,In_3156);
nor U607 (N_607,In_3829,In_1967);
xnor U608 (N_608,In_993,In_100);
and U609 (N_609,In_524,In_3038);
xnor U610 (N_610,In_2921,In_363);
xor U611 (N_611,In_1414,In_1236);
nand U612 (N_612,In_2499,In_162);
nand U613 (N_613,In_59,In_3415);
and U614 (N_614,In_1708,In_1391);
xor U615 (N_615,In_463,In_1676);
or U616 (N_616,In_4217,In_3814);
nor U617 (N_617,In_474,In_3324);
nand U618 (N_618,In_4688,In_2589);
nand U619 (N_619,In_3313,In_4720);
xor U620 (N_620,In_4395,In_1993);
xnor U621 (N_621,In_3303,In_67);
or U622 (N_622,In_4681,In_3264);
nand U623 (N_623,In_3222,In_4304);
xor U624 (N_624,In_3692,In_3054);
nor U625 (N_625,In_4174,In_1212);
or U626 (N_626,In_1310,In_1311);
and U627 (N_627,In_937,In_3793);
nand U628 (N_628,In_3439,In_3546);
nand U629 (N_629,In_3328,In_4510);
xor U630 (N_630,In_3258,In_2263);
nor U631 (N_631,In_1339,In_986);
and U632 (N_632,In_3704,In_1815);
nor U633 (N_633,In_1966,In_1470);
nand U634 (N_634,In_4805,In_1888);
xor U635 (N_635,In_1653,In_1614);
and U636 (N_636,In_2014,In_4444);
nand U637 (N_637,In_2980,In_3456);
or U638 (N_638,In_3455,In_531);
or U639 (N_639,In_1636,In_3738);
nand U640 (N_640,In_2953,In_4954);
nor U641 (N_641,In_3480,In_1315);
or U642 (N_642,In_2693,In_3786);
xor U643 (N_643,In_1748,In_1023);
nand U644 (N_644,In_4754,In_4818);
nand U645 (N_645,In_4192,In_1652);
nand U646 (N_646,In_3550,In_3625);
and U647 (N_647,In_900,In_3209);
xor U648 (N_648,In_3822,In_1080);
nand U649 (N_649,In_3143,In_1269);
or U650 (N_650,In_2976,In_4700);
nor U651 (N_651,In_3086,In_4458);
nor U652 (N_652,In_3909,In_4819);
nand U653 (N_653,In_2659,In_2502);
nand U654 (N_654,In_3428,In_614);
xnor U655 (N_655,In_3223,In_1381);
nand U656 (N_656,In_2670,In_3631);
nor U657 (N_657,In_3585,In_1571);
xnor U658 (N_658,In_3729,In_2337);
xor U659 (N_659,In_2786,In_2083);
and U660 (N_660,In_4359,In_1240);
xor U661 (N_661,In_1139,In_4099);
and U662 (N_662,In_2806,In_367);
xor U663 (N_663,In_3555,In_466);
xor U664 (N_664,In_26,In_3408);
and U665 (N_665,In_2638,In_496);
xnor U666 (N_666,In_1883,In_2956);
and U667 (N_667,In_3410,In_719);
nor U668 (N_668,In_4404,In_2592);
or U669 (N_669,In_3356,In_3650);
nor U670 (N_670,In_261,In_1924);
nand U671 (N_671,In_1694,In_4128);
xnor U672 (N_672,In_4173,In_4097);
xor U673 (N_673,In_4042,In_3488);
xor U674 (N_674,In_197,In_2970);
xor U675 (N_675,In_2523,In_4726);
and U676 (N_676,In_3623,In_1761);
xor U677 (N_677,In_3838,In_1969);
nor U678 (N_678,In_2699,In_1807);
and U679 (N_679,In_559,In_4793);
or U680 (N_680,In_193,In_1914);
nor U681 (N_681,In_2624,In_1733);
nand U682 (N_682,In_1171,In_2164);
nand U683 (N_683,In_2812,In_3659);
nor U684 (N_684,In_3752,In_2811);
nor U685 (N_685,In_4277,In_2397);
xor U686 (N_686,In_1732,In_2025);
or U687 (N_687,In_3106,In_1273);
nand U688 (N_688,In_2133,In_4146);
nor U689 (N_689,In_3534,In_408);
nand U690 (N_690,In_3358,In_3559);
nor U691 (N_691,In_3842,In_2819);
nor U692 (N_692,In_571,In_29);
nand U693 (N_693,In_4916,In_1791);
and U694 (N_694,In_4860,In_838);
or U695 (N_695,In_4285,In_3062);
or U696 (N_696,In_4778,In_3256);
xor U697 (N_697,In_1282,In_1469);
or U698 (N_698,In_360,In_2061);
nor U699 (N_699,In_2177,In_638);
nand U700 (N_700,In_1409,In_2252);
or U701 (N_701,In_2680,In_3074);
nor U702 (N_702,In_253,In_2607);
nor U703 (N_703,In_3991,In_3351);
or U704 (N_704,In_565,In_1873);
nor U705 (N_705,In_1083,In_4774);
xnor U706 (N_706,In_1837,In_4739);
and U707 (N_707,In_1402,In_3661);
or U708 (N_708,In_4125,In_2064);
nand U709 (N_709,In_2999,In_2297);
or U710 (N_710,In_3591,In_3739);
xor U711 (N_711,In_1506,In_4392);
and U712 (N_712,In_3787,In_4104);
nor U713 (N_713,In_437,In_180);
xor U714 (N_714,In_2658,In_1649);
nand U715 (N_715,In_4004,In_3199);
nor U716 (N_716,In_2993,In_2123);
nand U717 (N_717,In_89,In_3447);
and U718 (N_718,In_4839,In_4123);
nor U719 (N_719,In_450,In_4496);
nand U720 (N_720,In_3803,In_3160);
nor U721 (N_721,In_4995,In_4371);
and U722 (N_722,In_144,In_2151);
and U723 (N_723,In_4129,In_889);
xor U724 (N_724,In_4929,In_4901);
nand U725 (N_725,In_2081,In_3484);
nand U726 (N_726,In_2052,In_301);
or U727 (N_727,In_56,In_2901);
nor U728 (N_728,In_550,In_966);
or U729 (N_729,In_1323,In_4550);
nand U730 (N_730,In_922,In_3506);
nand U731 (N_731,In_1099,In_468);
or U732 (N_732,In_1776,In_1734);
or U733 (N_733,In_2905,In_2565);
or U734 (N_734,In_4475,In_2129);
nor U735 (N_735,In_3187,In_4114);
or U736 (N_736,In_3629,In_3406);
or U737 (N_737,In_3497,In_4102);
nand U738 (N_738,In_1123,In_1629);
xnor U739 (N_739,In_2829,In_3685);
and U740 (N_740,In_2823,In_4618);
or U741 (N_741,In_2561,In_4982);
xnor U742 (N_742,In_4275,In_558);
nand U743 (N_743,In_2392,In_4439);
and U744 (N_744,In_4980,In_878);
nand U745 (N_745,In_1811,In_1566);
xor U746 (N_746,In_4804,In_3776);
nor U747 (N_747,In_4826,In_647);
and U748 (N_748,In_2889,In_1992);
xnor U749 (N_749,In_1094,In_4336);
xor U750 (N_750,In_2651,In_185);
or U751 (N_751,In_1908,In_646);
and U752 (N_752,In_2460,In_1304);
nor U753 (N_753,In_119,In_2369);
nor U754 (N_754,In_2780,In_3365);
or U755 (N_755,In_143,In_2124);
or U756 (N_756,In_2251,In_1638);
and U757 (N_757,In_3467,In_3523);
nand U758 (N_758,In_4441,In_3846);
xor U759 (N_759,In_1703,In_1677);
and U760 (N_760,In_2237,In_2241);
or U761 (N_761,In_3908,In_1361);
or U762 (N_762,In_3165,In_4716);
or U763 (N_763,In_2788,In_972);
nand U764 (N_764,In_2229,In_49);
and U765 (N_765,In_2165,In_3524);
or U766 (N_766,In_4428,In_1896);
and U767 (N_767,In_687,In_1415);
nand U768 (N_768,In_775,In_2642);
nand U769 (N_769,In_3418,In_2800);
xor U770 (N_770,In_4415,In_1126);
and U771 (N_771,In_2350,In_1502);
nand U772 (N_772,In_2855,In_3886);
nand U773 (N_773,In_3795,In_633);
or U774 (N_774,In_4334,In_3587);
or U775 (N_775,In_734,In_2747);
and U776 (N_776,In_247,In_645);
nand U777 (N_777,In_1140,In_4373);
nand U778 (N_778,In_2730,In_4820);
and U779 (N_779,In_1342,In_2859);
xnor U780 (N_780,In_4136,In_1317);
and U781 (N_781,In_2206,In_1313);
xnor U782 (N_782,In_2433,In_1682);
nand U783 (N_783,In_186,In_1426);
or U784 (N_784,In_4297,In_519);
or U785 (N_785,In_1655,In_2368);
xnor U786 (N_786,In_45,In_214);
or U787 (N_787,In_2212,In_691);
nand U788 (N_788,In_84,In_3994);
and U789 (N_789,In_3277,In_1817);
or U790 (N_790,In_385,In_4772);
and U791 (N_791,In_347,In_2065);
and U792 (N_792,In_3007,In_3244);
nand U793 (N_793,In_1238,In_1886);
xor U794 (N_794,In_3412,In_1802);
or U795 (N_795,In_581,In_1977);
xnor U796 (N_796,In_1436,In_2291);
and U797 (N_797,In_4253,In_2484);
nor U798 (N_798,In_3861,In_3525);
xnor U799 (N_799,In_2622,In_1442);
xor U800 (N_800,In_305,In_3364);
or U801 (N_801,In_820,In_648);
nor U802 (N_802,In_467,In_2037);
xor U803 (N_803,In_2899,In_4463);
and U804 (N_804,In_1202,In_1552);
or U805 (N_805,In_811,In_12);
xnor U806 (N_806,In_4651,In_178);
and U807 (N_807,In_1857,In_2195);
nand U808 (N_808,In_334,In_3110);
or U809 (N_809,In_4886,In_521);
nor U810 (N_810,In_3712,In_3821);
xor U811 (N_811,In_4615,In_112);
xnor U812 (N_812,In_3582,In_1019);
xor U813 (N_813,In_2843,In_3298);
or U814 (N_814,In_4760,In_1635);
xnor U815 (N_815,In_4844,In_2348);
nor U816 (N_816,In_1413,In_4274);
xnor U817 (N_817,In_480,In_3945);
nand U818 (N_818,In_1563,In_4206);
and U819 (N_819,In_3273,In_188);
or U820 (N_820,In_1540,In_3671);
or U821 (N_821,In_2027,In_1217);
or U822 (N_822,In_4153,In_4179);
xnor U823 (N_823,In_1117,In_4753);
or U824 (N_824,In_2679,In_2134);
and U825 (N_825,In_619,In_2141);
nand U826 (N_826,In_1395,In_895);
nand U827 (N_827,In_1194,In_918);
and U828 (N_828,In_2380,In_2054);
nor U829 (N_829,In_4191,In_1984);
and U830 (N_830,In_1553,In_4802);
or U831 (N_831,In_507,In_4364);
nor U832 (N_832,In_2386,In_3423);
xor U833 (N_833,In_4003,In_949);
or U834 (N_834,In_359,In_636);
nor U835 (N_835,In_3713,In_3517);
and U836 (N_836,In_3225,In_3114);
nor U837 (N_837,In_3250,In_1092);
or U838 (N_838,In_1970,In_2576);
xor U839 (N_839,In_3726,In_1863);
xnor U840 (N_840,In_3551,In_951);
nor U841 (N_841,In_3676,In_4060);
and U842 (N_842,In_30,In_1534);
xnor U843 (N_843,In_1550,In_3169);
and U844 (N_844,In_3087,In_4440);
or U845 (N_845,In_3158,In_3843);
and U846 (N_846,In_4390,In_4436);
and U847 (N_847,In_2138,In_2409);
nor U848 (N_848,In_1688,In_4044);
or U849 (N_849,In_535,In_608);
and U850 (N_850,In_779,In_1132);
xnor U851 (N_851,In_577,In_1889);
xnor U852 (N_852,In_552,In_868);
nand U853 (N_853,In_4384,In_676);
nor U854 (N_854,In_3751,In_4118);
nand U855 (N_855,In_4158,In_3593);
and U856 (N_856,In_106,In_945);
xor U857 (N_857,In_4483,In_3898);
xnor U858 (N_858,In_555,In_4283);
or U859 (N_859,In_2379,In_3420);
nor U860 (N_860,In_4611,In_3995);
or U861 (N_861,In_3647,In_1036);
xor U862 (N_862,In_2844,In_4424);
or U863 (N_863,In_1696,In_2911);
nand U864 (N_864,In_232,In_1009);
xor U865 (N_865,In_2712,In_3445);
nor U866 (N_866,In_1723,In_2983);
or U867 (N_867,In_2394,In_1296);
or U868 (N_868,In_722,In_2339);
nand U869 (N_869,In_1633,In_4675);
nand U870 (N_870,In_2228,In_4072);
nand U871 (N_871,In_1262,In_4764);
and U872 (N_872,In_153,In_2646);
nor U873 (N_873,In_753,In_902);
nand U874 (N_874,In_1981,In_3262);
or U875 (N_875,In_4215,In_861);
xor U876 (N_876,In_3253,In_1074);
or U877 (N_877,In_4412,In_4558);
or U878 (N_878,In_3145,In_4601);
nor U879 (N_879,In_4891,In_1438);
or U880 (N_880,In_4023,In_2721);
nand U881 (N_881,In_3003,In_1606);
xor U882 (N_882,In_3554,In_2794);
nor U883 (N_883,In_3833,In_2213);
and U884 (N_884,In_1378,In_1033);
nor U885 (N_885,In_2985,In_876);
nand U886 (N_886,In_4162,In_406);
or U887 (N_887,In_3779,In_1498);
xnor U888 (N_888,In_2931,In_2998);
xnor U889 (N_889,In_73,In_3157);
nor U890 (N_890,In_2172,In_1821);
nand U891 (N_891,In_1062,In_3451);
xor U892 (N_892,In_1865,In_1181);
and U893 (N_893,In_241,In_4421);
nor U894 (N_894,In_4235,In_1872);
or U895 (N_895,In_2220,In_3716);
or U896 (N_896,In_1330,In_2965);
xnor U897 (N_897,In_892,In_2894);
and U898 (N_898,In_4707,In_4710);
nor U899 (N_899,In_4647,In_4372);
and U900 (N_900,In_3179,In_4337);
xnor U901 (N_901,In_1122,In_2320);
and U902 (N_902,In_2001,In_2452);
nor U903 (N_903,In_3388,In_7);
or U904 (N_904,In_1187,In_2500);
or U905 (N_905,In_3526,In_2080);
nand U906 (N_906,In_3825,In_4141);
nand U907 (N_907,In_1698,In_623);
xnor U908 (N_908,In_1740,In_1101);
and U909 (N_909,In_2335,In_3309);
nand U910 (N_910,In_2071,In_1866);
or U911 (N_911,In_4445,In_3941);
or U912 (N_912,In_2246,In_606);
or U913 (N_913,In_721,In_3977);
and U914 (N_914,In_4408,In_4752);
nor U915 (N_915,In_323,In_3437);
or U916 (N_916,In_1082,In_1906);
nand U917 (N_917,In_4388,In_1900);
nand U918 (N_918,In_3192,In_1999);
xor U919 (N_919,In_4921,In_2035);
and U920 (N_920,In_4468,In_4197);
and U921 (N_921,In_4974,In_2063);
xnor U922 (N_922,In_3556,In_2630);
and U923 (N_923,In_315,In_3758);
or U924 (N_924,In_1266,In_3130);
nor U925 (N_925,In_4581,In_3435);
and U926 (N_926,In_3925,In_3260);
or U927 (N_927,In_4909,In_523);
or U928 (N_928,In_1063,In_263);
nor U929 (N_929,In_3812,In_2696);
nand U930 (N_930,In_1496,In_3427);
nor U931 (N_931,In_391,In_411);
xor U932 (N_932,In_3985,In_1372);
or U933 (N_933,In_4294,In_3567);
nor U934 (N_934,In_494,In_2406);
or U935 (N_935,In_4016,In_855);
xnor U936 (N_936,In_4926,In_2594);
and U937 (N_937,In_1852,In_1624);
nor U938 (N_938,In_2367,In_3017);
xor U939 (N_939,In_1254,In_3032);
and U940 (N_940,In_3500,In_1903);
xor U941 (N_941,In_2948,In_4121);
xor U942 (N_942,In_4988,In_2089);
or U943 (N_943,In_4512,In_2902);
nor U944 (N_944,In_76,In_4077);
nand U945 (N_945,In_915,In_1528);
xnor U946 (N_946,In_3426,In_4799);
nor U947 (N_947,In_4727,In_3518);
and U948 (N_948,In_1749,In_771);
nand U949 (N_949,In_1255,In_3013);
xnor U950 (N_950,In_563,In_4748);
xor U951 (N_951,In_79,In_2870);
xor U952 (N_952,In_416,In_3000);
nor U953 (N_953,In_2039,In_1681);
nor U954 (N_954,In_1058,In_3363);
and U955 (N_955,In_3419,In_486);
or U956 (N_956,In_4847,In_2360);
nor U957 (N_957,In_4142,In_3665);
or U958 (N_958,In_150,In_3034);
nand U959 (N_959,In_1351,In_3902);
and U960 (N_960,In_4156,In_4777);
nor U961 (N_961,In_4282,In_556);
nand U962 (N_962,In_4116,In_2219);
or U963 (N_963,In_189,In_3589);
xnor U964 (N_964,In_3750,In_2214);
xnor U965 (N_965,In_2515,In_2601);
nor U966 (N_966,In_2022,In_3560);
nor U967 (N_967,In_1234,In_1277);
or U968 (N_968,In_2817,In_4246);
xnor U969 (N_969,In_3460,In_605);
xnor U970 (N_970,In_4873,In_4144);
and U971 (N_971,In_3618,In_3163);
xnor U972 (N_972,In_1987,In_1803);
or U973 (N_973,In_1045,In_2149);
or U974 (N_974,In_355,In_498);
or U975 (N_975,In_4667,In_4154);
xor U976 (N_976,In_1109,In_2966);
and U977 (N_977,In_857,In_740);
xor U978 (N_978,In_2422,In_4243);
nand U979 (N_979,In_2259,In_3754);
nor U980 (N_980,In_1108,In_3545);
and U981 (N_981,In_349,In_1623);
and U982 (N_982,In_2376,In_2703);
or U983 (N_983,In_4822,In_1472);
nor U984 (N_984,In_3586,In_4792);
xor U985 (N_985,In_4636,In_4309);
nor U986 (N_986,In_2307,In_1907);
or U987 (N_987,In_621,In_4500);
nor U988 (N_988,In_3724,In_4941);
xnor U989 (N_989,In_3378,In_4766);
nor U990 (N_990,In_3448,In_4603);
or U991 (N_991,In_2053,In_4157);
or U992 (N_992,In_1191,In_2895);
and U993 (N_993,In_4970,In_2006);
nor U994 (N_994,In_3973,In_4567);
xor U995 (N_995,In_1919,In_4894);
or U996 (N_996,In_4842,In_2771);
or U997 (N_997,In_4664,In_138);
and U998 (N_998,In_762,In_3785);
nand U999 (N_999,In_3228,In_1767);
nand U1000 (N_1000,In_2135,In_3960);
xnor U1001 (N_1001,In_440,In_3233);
and U1002 (N_1002,In_1133,In_4898);
nand U1003 (N_1003,In_462,In_3788);
nor U1004 (N_1004,In_1780,In_3519);
nand U1005 (N_1005,In_4696,In_1838);
nand U1006 (N_1006,In_2116,In_4505);
or U1007 (N_1007,In_3342,In_3401);
or U1008 (N_1008,In_815,In_3652);
or U1009 (N_1009,In_1389,In_705);
nand U1010 (N_1010,In_3501,In_924);
and U1011 (N_1011,In_4376,In_1318);
nor U1012 (N_1012,In_129,In_3020);
nand U1013 (N_1013,In_442,In_3316);
or U1014 (N_1014,In_4920,In_1544);
and U1015 (N_1015,In_1166,In_103);
or U1016 (N_1016,In_3398,In_4299);
xor U1017 (N_1017,In_1897,In_4148);
or U1018 (N_1018,In_2672,In_2711);
xor U1019 (N_1019,In_858,In_3493);
nand U1020 (N_1020,In_3527,In_3367);
nor U1021 (N_1021,In_4513,In_785);
and U1022 (N_1022,In_2804,In_307);
and U1023 (N_1023,In_2834,In_1691);
and U1024 (N_1024,In_3837,In_262);
xnor U1025 (N_1025,In_1769,In_402);
nor U1026 (N_1026,In_2562,In_2420);
and U1027 (N_1027,In_1665,In_3646);
nand U1028 (N_1028,In_2749,In_2718);
nor U1029 (N_1029,In_723,In_2766);
and U1030 (N_1030,In_2863,In_4747);
xor U1031 (N_1031,In_3081,In_4562);
or U1032 (N_1032,In_3974,In_1885);
and U1033 (N_1033,In_2466,In_3709);
or U1034 (N_1034,In_3740,In_3308);
nand U1035 (N_1035,In_732,In_2904);
nor U1036 (N_1036,In_4208,In_409);
nand U1037 (N_1037,In_65,In_1170);
nor U1038 (N_1038,In_908,In_3965);
or U1039 (N_1039,In_2474,In_3730);
xor U1040 (N_1040,In_1333,In_1843);
nor U1041 (N_1041,In_3603,In_1626);
nor U1042 (N_1042,In_3044,In_3686);
xor U1043 (N_1043,In_639,In_1145);
nor U1044 (N_1044,In_620,In_2097);
or U1045 (N_1045,In_952,In_3990);
xor U1046 (N_1046,In_534,In_1945);
nand U1047 (N_1047,In_874,In_4470);
or U1048 (N_1048,In_4597,In_3915);
or U1049 (N_1049,In_2896,In_423);
or U1050 (N_1050,In_447,In_2545);
xor U1051 (N_1051,In_885,In_4949);
xor U1052 (N_1052,In_3981,In_2402);
and U1053 (N_1053,In_4219,In_1180);
or U1054 (N_1054,In_1131,In_1119);
xor U1055 (N_1055,In_2784,In_219);
or U1056 (N_1056,In_4928,In_1634);
and U1057 (N_1057,In_2762,In_1923);
and U1058 (N_1058,In_1721,In_3578);
nand U1059 (N_1059,In_773,In_882);
or U1060 (N_1060,In_1347,In_4823);
nor U1061 (N_1061,In_2742,In_396);
and U1062 (N_1062,In_354,In_1877);
xnor U1063 (N_1063,In_4994,In_3756);
or U1064 (N_1064,In_2611,In_3266);
nor U1065 (N_1065,In_4432,In_192);
nand U1066 (N_1066,In_793,In_1592);
and U1067 (N_1067,In_1253,In_3594);
nand U1068 (N_1068,In_1345,In_2098);
nand U1069 (N_1069,In_2548,In_3728);
xnor U1070 (N_1070,In_4831,In_2720);
or U1071 (N_1071,In_3639,In_448);
xnor U1072 (N_1072,In_3279,In_2239);
nor U1073 (N_1073,In_1383,In_3771);
nor U1074 (N_1074,In_939,In_4978);
xor U1075 (N_1075,In_3931,In_803);
and U1076 (N_1076,In_3873,In_2559);
or U1077 (N_1077,In_2377,In_1337);
nor U1078 (N_1078,In_630,In_2234);
xor U1079 (N_1079,In_2675,In_288);
or U1080 (N_1080,In_2598,In_1225);
and U1081 (N_1081,In_4247,In_4882);
nand U1082 (N_1082,In_3395,In_1473);
and U1083 (N_1083,In_685,In_2021);
xnor U1084 (N_1084,In_2538,In_789);
or U1085 (N_1085,In_1565,In_3613);
or U1086 (N_1086,In_4975,In_2166);
nand U1087 (N_1087,In_1988,In_1792);
nand U1088 (N_1088,In_1532,In_1416);
or U1089 (N_1089,In_2569,In_4973);
and U1090 (N_1090,In_866,In_4750);
nor U1091 (N_1091,In_2030,In_1574);
or U1092 (N_1092,In_4932,In_696);
nor U1093 (N_1093,In_4574,In_3722);
nor U1094 (N_1094,In_2664,In_1027);
xnor U1095 (N_1095,In_4222,In_3907);
nor U1096 (N_1096,In_4504,In_2773);
nand U1097 (N_1097,In_3718,In_4383);
nand U1098 (N_1098,In_2649,In_4499);
nor U1099 (N_1099,In_4199,In_2727);
and U1100 (N_1100,In_3218,In_584);
xnor U1101 (N_1101,In_2736,In_4351);
nand U1102 (N_1102,In_4133,In_4811);
nor U1103 (N_1103,In_683,In_3549);
and U1104 (N_1104,In_137,In_281);
nand U1105 (N_1105,In_4330,In_990);
nor U1106 (N_1106,In_2864,In_944);
or U1107 (N_1107,In_2763,In_3183);
xor U1108 (N_1108,In_4796,In_3581);
xor U1109 (N_1109,In_1230,In_1057);
and U1110 (N_1110,In_4552,In_3514);
nor U1111 (N_1111,In_3865,In_109);
nor U1112 (N_1112,In_3830,In_292);
nand U1113 (N_1113,In_4669,In_4050);
and U1114 (N_1114,In_760,In_1035);
nor U1115 (N_1115,In_551,In_1450);
or U1116 (N_1116,In_3969,In_491);
xor U1117 (N_1117,In_258,In_1454);
or U1118 (N_1118,In_390,In_2603);
xor U1119 (N_1119,In_4670,In_888);
xnor U1120 (N_1120,In_1012,In_3828);
or U1121 (N_1121,In_693,In_3475);
or U1122 (N_1122,In_928,In_4323);
and U1123 (N_1123,In_831,In_931);
xnor U1124 (N_1124,In_3856,In_3470);
or U1125 (N_1125,In_3175,In_1965);
or U1126 (N_1126,In_2334,In_4902);
nor U1127 (N_1127,In_4329,In_3894);
nor U1128 (N_1128,In_4030,In_2357);
xnor U1129 (N_1129,In_80,In_4074);
xor U1130 (N_1130,In_2155,In_798);
nand U1131 (N_1131,In_4654,In_3268);
xnor U1132 (N_1132,In_2384,In_1912);
nor U1133 (N_1133,In_4773,In_3850);
or U1134 (N_1134,In_4027,In_35);
nand U1135 (N_1135,In_4037,In_971);
or U1136 (N_1136,In_528,In_2748);
nor U1137 (N_1137,In_1477,In_4816);
or U1138 (N_1138,In_3343,In_756);
nand U1139 (N_1139,In_4610,In_395);
and U1140 (N_1140,In_2564,In_2043);
nor U1141 (N_1141,In_541,In_3338);
nor U1142 (N_1142,In_1116,In_302);
nor U1143 (N_1143,In_880,In_1731);
and U1144 (N_1144,In_742,In_3202);
and U1145 (N_1145,In_3648,In_1444);
nor U1146 (N_1146,In_177,In_4265);
xnor U1147 (N_1147,In_2982,In_3051);
nor U1148 (N_1148,In_4103,In_2719);
and U1149 (N_1149,In_1994,In_1512);
xor U1150 (N_1150,In_1206,In_2733);
or U1151 (N_1151,In_3864,In_4578);
or U1152 (N_1152,In_3104,In_2183);
nand U1153 (N_1153,In_3727,In_338);
and U1154 (N_1154,In_4352,In_609);
nand U1155 (N_1155,In_4570,In_1890);
and U1156 (N_1156,In_4855,In_1997);
nand U1157 (N_1157,In_3065,In_4480);
nand U1158 (N_1158,In_425,In_4767);
xnor U1159 (N_1159,In_2636,In_2596);
nor U1160 (N_1160,In_1554,In_3094);
nor U1161 (N_1161,In_3983,In_2473);
nor U1162 (N_1162,In_3147,In_4335);
xor U1163 (N_1163,In_2244,In_120);
nand U1164 (N_1164,In_697,In_1338);
and U1165 (N_1165,In_4966,In_4521);
nor U1166 (N_1166,In_1137,In_4140);
or U1167 (N_1167,In_2286,In_376);
nand U1168 (N_1168,In_3503,In_2390);
or U1169 (N_1169,In_1747,In_2236);
or U1170 (N_1170,In_4596,In_3107);
and U1171 (N_1171,In_3022,In_2248);
nor U1172 (N_1172,In_2181,In_4328);
or U1173 (N_1173,In_1013,In_4021);
xnor U1174 (N_1174,In_4237,In_2639);
nand U1175 (N_1175,In_116,In_795);
xor U1176 (N_1176,In_4478,In_500);
and U1177 (N_1177,In_3409,In_2261);
xor U1178 (N_1178,In_82,In_3512);
nor U1179 (N_1179,In_3177,In_8);
xnor U1180 (N_1180,In_3276,In_808);
xnor U1181 (N_1181,In_1725,In_4671);
nand U1182 (N_1182,In_913,In_4733);
nor U1183 (N_1183,In_1702,In_932);
xnor U1184 (N_1184,In_4261,In_3023);
nand U1185 (N_1185,In_573,In_4134);
xor U1186 (N_1186,In_434,In_3288);
nand U1187 (N_1187,In_225,In_4502);
nor U1188 (N_1188,In_2416,In_2528);
nand U1189 (N_1189,In_2382,In_4661);
nor U1190 (N_1190,In_1711,In_3048);
nor U1191 (N_1191,In_4349,In_4836);
nor U1192 (N_1192,In_4518,In_2832);
and U1193 (N_1193,In_1667,In_2635);
nand U1194 (N_1194,In_960,In_2163);
and U1195 (N_1195,In_3301,In_4403);
nor U1196 (N_1196,In_3468,In_2776);
and U1197 (N_1197,In_1151,In_4117);
and U1198 (N_1198,In_1583,In_264);
xnor U1199 (N_1199,In_81,In_2520);
xnor U1200 (N_1200,In_3819,In_3694);
nor U1201 (N_1201,In_4779,In_1185);
and U1202 (N_1202,In_975,In_1455);
nor U1203 (N_1203,In_1657,In_2932);
xnor U1204 (N_1204,In_3380,In_4211);
nand U1205 (N_1205,In_3131,In_3673);
or U1206 (N_1206,In_4869,In_821);
nand U1207 (N_1207,In_4236,In_204);
xnor U1208 (N_1208,In_2366,In_822);
xor U1209 (N_1209,In_4937,In_1475);
or U1210 (N_1210,In_1705,In_495);
nor U1211 (N_1211,In_4708,In_2709);
and U1212 (N_1212,In_2613,In_1641);
nor U1213 (N_1213,In_3636,In_3006);
and U1214 (N_1214,In_4262,In_2753);
xor U1215 (N_1215,In_2272,In_4922);
and U1216 (N_1216,In_3443,In_1936);
nor U1217 (N_1217,In_3695,In_2628);
nand U1218 (N_1218,In_2305,In_1305);
nand U1219 (N_1219,In_2362,In_3188);
and U1220 (N_1220,In_2434,In_4536);
or U1221 (N_1221,In_394,In_1699);
nor U1222 (N_1222,In_765,In_4438);
or U1223 (N_1223,In_1480,In_562);
nand U1224 (N_1224,In_817,In_289);
nand U1225 (N_1225,In_4258,In_3734);
nand U1226 (N_1226,In_4829,In_47);
xnor U1227 (N_1227,In_2790,In_160);
nand U1228 (N_1228,In_361,In_2431);
and U1229 (N_1229,In_400,In_4678);
xnor U1230 (N_1230,In_4381,In_2193);
nand U1231 (N_1231,In_4288,In_4160);
nand U1232 (N_1232,In_3206,In_758);
xor U1233 (N_1233,In_2575,In_652);
nor U1234 (N_1234,In_4249,In_3012);
nor U1235 (N_1235,In_227,In_2346);
and U1236 (N_1236,In_19,In_3080);
nor U1237 (N_1237,In_4749,In_2192);
nand U1238 (N_1238,In_3154,In_591);
nand U1239 (N_1239,In_4452,In_4348);
nor U1240 (N_1240,In_1996,In_3966);
and U1241 (N_1241,In_1590,In_1938);
nand U1242 (N_1242,In_3790,In_4571);
nor U1243 (N_1243,In_2714,In_78);
or U1244 (N_1244,In_3383,In_4172);
and U1245 (N_1245,In_3030,In_24);
or U1246 (N_1246,In_805,In_4287);
nand U1247 (N_1247,In_2355,In_2399);
xnor U1248 (N_1248,In_389,In_2073);
xnor U1249 (N_1249,In_2042,In_2713);
and U1250 (N_1250,In_1785,In_569);
or U1251 (N_1251,In_2430,In_4101);
or U1252 (N_1252,In_595,In_1275);
and U1253 (N_1253,In_2637,In_537);
nand U1254 (N_1254,In_4396,In_1719);
and U1255 (N_1255,In_4565,In_4737);
or U1256 (N_1256,In_2000,In_4650);
xnor U1257 (N_1257,In_3693,In_2476);
nand U1258 (N_1258,In_1750,In_3668);
xor U1259 (N_1259,In_4292,In_4540);
and U1260 (N_1260,In_1192,In_4537);
xor U1261 (N_1261,In_1830,In_2822);
xor U1262 (N_1262,In_1887,In_101);
nor U1263 (N_1263,In_2168,In_293);
nor U1264 (N_1264,In_4551,In_4223);
and U1265 (N_1265,In_2099,In_477);
xor U1266 (N_1266,In_3820,In_4430);
and U1267 (N_1267,In_2968,In_4742);
xnor U1268 (N_1268,In_3211,In_436);
nand U1269 (N_1269,In_650,In_1855);
xor U1270 (N_1270,In_1542,In_3018);
nand U1271 (N_1271,In_2469,In_1539);
and U1272 (N_1272,In_1276,In_3354);
xor U1273 (N_1273,In_3307,In_4765);
or U1274 (N_1274,In_1701,In_432);
or U1275 (N_1275,In_1686,In_2436);
or U1276 (N_1276,In_1910,In_4053);
nor U1277 (N_1277,In_4702,In_3055);
and U1278 (N_1278,In_2119,In_2927);
and U1279 (N_1279,In_4090,In_4957);
and U1280 (N_1280,In_953,In_751);
and U1281 (N_1281,In_3182,In_4530);
or U1282 (N_1282,In_1331,In_2408);
or U1283 (N_1283,In_3792,In_1115);
and U1284 (N_1284,In_1227,In_4606);
xor U1285 (N_1285,In_3057,In_4635);
nor U1286 (N_1286,In_1654,In_2793);
nand U1287 (N_1287,In_1248,In_3121);
and U1288 (N_1288,In_2949,In_2978);
and U1289 (N_1289,In_1893,In_4959);
nor U1290 (N_1290,In_499,In_2471);
and U1291 (N_1291,In_1112,In_610);
or U1292 (N_1292,In_4584,In_2329);
nand U1293 (N_1293,In_2862,In_3910);
nor U1294 (N_1294,In_1519,In_4788);
xnor U1295 (N_1295,In_538,In_3085);
or U1296 (N_1296,In_4944,In_343);
xor U1297 (N_1297,In_725,In_4120);
or U1298 (N_1298,In_1662,In_1879);
nand U1299 (N_1299,In_2110,In_681);
or U1300 (N_1300,In_1751,In_1223);
and U1301 (N_1301,In_3869,In_1790);
nand U1302 (N_1302,In_4165,In_3385);
and U1303 (N_1303,In_3958,In_4763);
and U1304 (N_1304,In_2429,In_3507);
or U1305 (N_1305,In_4063,In_3509);
or U1306 (N_1306,In_1775,In_152);
nor U1307 (N_1307,In_3684,In_3816);
xnor U1308 (N_1308,In_1546,In_1551);
and U1309 (N_1309,In_4485,In_4231);
and U1310 (N_1310,In_1770,In_3731);
xor U1311 (N_1311,In_582,In_4884);
and U1312 (N_1312,In_303,In_2412);
and U1313 (N_1313,In_2287,In_4131);
nand U1314 (N_1314,In_1971,In_217);
nor U1315 (N_1315,In_4194,In_700);
and U1316 (N_1316,In_4663,In_3494);
nor U1317 (N_1317,In_1046,In_3123);
and U1318 (N_1318,In_4809,In_3912);
nor U1319 (N_1319,In_88,In_2583);
nand U1320 (N_1320,In_4856,In_2090);
or U1321 (N_1321,In_61,In_415);
and U1322 (N_1322,In_4476,In_3332);
xnor U1323 (N_1323,In_2488,In_2353);
xor U1324 (N_1324,In_206,In_2454);
nand U1325 (N_1325,In_4849,In_3058);
and U1326 (N_1326,In_2308,In_1458);
nand U1327 (N_1327,In_2031,In_2922);
and U1328 (N_1328,In_4933,In_1075);
nand U1329 (N_1329,In_4709,In_141);
or U1330 (N_1330,In_25,In_4897);
and U1331 (N_1331,In_3305,In_2586);
nand U1332 (N_1332,In_4858,In_4307);
and U1333 (N_1333,In_2480,In_2505);
and U1334 (N_1334,In_1177,In_1200);
or U1335 (N_1335,In_2882,In_1639);
and U1336 (N_1336,In_1358,In_4036);
xor U1337 (N_1337,In_3394,In_4592);
xnor U1338 (N_1338,In_2587,In_1176);
nand U1339 (N_1339,In_2341,In_1493);
xnor U1340 (N_1340,In_1406,In_574);
and U1341 (N_1341,In_4938,In_1847);
xnor U1342 (N_1342,In_2342,In_575);
nand U1343 (N_1343,In_926,In_350);
nor U1344 (N_1344,In_4813,In_38);
and U1345 (N_1345,In_4509,In_2608);
nor U1346 (N_1346,In_2103,In_2401);
nor U1347 (N_1347,In_3643,In_3959);
and U1348 (N_1348,In_306,In_2157);
and U1349 (N_1349,In_4758,In_4143);
and U1350 (N_1350,In_4879,In_923);
nor U1351 (N_1351,In_3633,In_2250);
or U1352 (N_1352,In_3638,In_1232);
nand U1353 (N_1353,In_1492,In_1658);
nor U1354 (N_1354,In_3111,In_2612);
xnor U1355 (N_1355,In_2018,In_2249);
or U1356 (N_1356,In_2479,In_3670);
or U1357 (N_1357,In_284,In_4694);
xnor U1358 (N_1358,In_1744,In_3243);
or U1359 (N_1359,In_260,In_3392);
and U1360 (N_1360,In_4868,In_3015);
xor U1361 (N_1361,In_1951,In_1020);
nor U1362 (N_1362,In_1726,In_2359);
and U1363 (N_1363,In_4548,In_3674);
and U1364 (N_1364,In_251,In_786);
nor U1365 (N_1365,In_1068,In_3721);
xor U1366 (N_1366,In_628,In_3361);
xor U1367 (N_1367,In_4835,In_4069);
or U1368 (N_1368,In_2657,In_2805);
and U1369 (N_1369,In_1881,In_379);
or U1370 (N_1370,In_3630,In_863);
nand U1371 (N_1371,In_894,In_375);
and U1372 (N_1372,In_3482,In_3759);
or U1373 (N_1373,In_2705,In_3558);
nand U1374 (N_1374,In_2994,In_2415);
or U1375 (N_1375,In_4071,In_3496);
or U1376 (N_1376,In_1086,In_3370);
nor U1377 (N_1377,In_2689,In_1447);
nor U1378 (N_1378,In_3379,In_4587);
nand U1379 (N_1379,In_3835,In_3138);
nand U1380 (N_1380,In_4984,In_3720);
nand U1381 (N_1381,In_1195,In_3291);
xor U1382 (N_1382,In_3891,In_3920);
or U1383 (N_1383,In_4919,In_3553);
and U1384 (N_1384,In_4789,In_2926);
nor U1385 (N_1385,In_2223,In_3620);
nand U1386 (N_1386,In_3855,In_3905);
or U1387 (N_1387,In_4880,In_441);
nand U1388 (N_1388,In_669,In_3548);
nor U1389 (N_1389,In_3314,In_510);
nand U1390 (N_1390,In_3634,In_1252);
nor U1391 (N_1391,In_1976,In_2857);
nand U1392 (N_1392,In_578,In_4721);
and U1393 (N_1393,In_63,In_3438);
or U1394 (N_1394,In_1320,In_3663);
and U1395 (N_1395,In_4311,In_3951);
nand U1396 (N_1396,In_1956,In_1950);
or U1397 (N_1397,In_1884,In_3826);
and U1398 (N_1398,In_1038,In_4252);
and U1399 (N_1399,In_4229,In_3683);
xor U1400 (N_1400,In_1679,In_3893);
xnor U1401 (N_1401,In_1385,In_1479);
nand U1402 (N_1402,In_3148,In_348);
nor U1403 (N_1403,In_1188,In_4761);
nor U1404 (N_1404,In_3911,In_1348);
nor U1405 (N_1405,In_4892,In_3261);
or U1406 (N_1406,In_3688,In_2764);
nand U1407 (N_1407,In_4427,In_205);
or U1408 (N_1408,In_4083,In_3654);
or U1409 (N_1409,In_3009,In_1284);
and U1410 (N_1410,In_1368,In_3797);
or U1411 (N_1411,In_905,In_2443);
nand U1412 (N_1412,In_2694,In_3161);
xnor U1413 (N_1413,In_2778,In_3024);
nor U1414 (N_1414,In_1547,In_2716);
and U1415 (N_1415,In_841,In_3005);
and U1416 (N_1416,In_1067,In_1220);
nor U1417 (N_1417,In_2674,In_4151);
or U1418 (N_1418,In_1478,In_459);
xor U1419 (N_1419,In_3194,In_3259);
nand U1420 (N_1420,In_3068,In_1834);
and U1421 (N_1421,In_3184,In_1765);
nand U1422 (N_1422,In_2761,In_4029);
and U1423 (N_1423,In_983,In_2275);
and U1424 (N_1424,In_4181,In_1579);
and U1425 (N_1425,In_711,In_3944);
nor U1426 (N_1426,In_664,In_187);
nor U1427 (N_1427,In_1986,In_505);
nor U1428 (N_1428,In_3478,In_3571);
or U1429 (N_1429,In_824,In_4586);
or U1430 (N_1430,In_1141,In_920);
nand U1431 (N_1431,In_4729,In_2302);
nor U1432 (N_1432,In_1095,In_3600);
nand U1433 (N_1433,In_3903,In_4520);
nand U1434 (N_1434,In_333,In_3076);
nor U1435 (N_1435,In_897,In_2745);
and U1436 (N_1436,In_3286,In_4832);
nor U1437 (N_1437,In_3680,In_3877);
and U1438 (N_1438,In_4846,In_852);
or U1439 (N_1439,In_316,In_2482);
and U1440 (N_1440,In_766,In_2281);
and U1441 (N_1441,In_3541,In_1515);
nand U1442 (N_1442,In_3339,In_1281);
nor U1443 (N_1443,In_1829,In_1593);
or U1444 (N_1444,In_622,In_2490);
nand U1445 (N_1445,In_1543,In_4514);
xnor U1446 (N_1446,In_404,In_2146);
xor U1447 (N_1447,In_4081,In_2604);
xnor U1448 (N_1448,In_2537,In_2553);
and U1449 (N_1449,In_3899,In_3714);
nor U1450 (N_1450,In_1397,In_2943);
xnor U1451 (N_1451,In_3381,In_433);
or U1452 (N_1452,In_3477,In_4728);
or U1453 (N_1453,In_3737,In_2555);
xor U1454 (N_1454,In_3190,In_4682);
nand U1455 (N_1455,In_4098,In_588);
and U1456 (N_1456,In_2109,In_275);
xor U1457 (N_1457,In_136,In_365);
nand U1458 (N_1458,In_4658,In_1102);
or U1459 (N_1459,In_3575,In_580);
and U1460 (N_1460,In_730,In_4343);
and U1461 (N_1461,In_3896,In_4762);
xnor U1462 (N_1462,In_3056,In_670);
nand U1463 (N_1463,In_1599,In_2087);
nor U1464 (N_1464,In_804,In_3203);
nor U1465 (N_1465,In_2207,In_4583);
nor U1466 (N_1466,In_4018,In_1476);
xnor U1467 (N_1467,In_2688,In_3773);
or U1468 (N_1468,In_2049,In_4481);
nor U1469 (N_1469,In_2827,In_2660);
nor U1470 (N_1470,In_579,In_2066);
nor U1471 (N_1471,In_3942,In_752);
nand U1472 (N_1472,In_2549,In_4590);
nand U1473 (N_1473,In_4303,In_4950);
xnor U1474 (N_1474,In_4526,In_4115);
or U1475 (N_1475,In_1257,In_2437);
and U1476 (N_1476,In_3580,In_4313);
xor U1477 (N_1477,In_847,In_1507);
xnor U1478 (N_1478,In_85,In_583);
xnor U1479 (N_1479,In_3459,In_2036);
or U1480 (N_1480,In_1295,In_978);
nand U1481 (N_1481,In_3053,In_788);
or U1482 (N_1482,In_2886,In_4429);
nand U1483 (N_1483,In_4497,In_4963);
nor U1484 (N_1484,In_3998,In_4474);
or U1485 (N_1485,In_2019,In_3033);
and U1486 (N_1486,In_3658,In_2493);
nand U1487 (N_1487,In_508,In_3402);
xnor U1488 (N_1488,In_2310,In_2738);
nand U1489 (N_1489,In_2374,In_4848);
nand U1490 (N_1490,In_1114,In_587);
or U1491 (N_1491,In_1533,In_3596);
or U1492 (N_1492,In_2062,In_4511);
nor U1493 (N_1493,In_2552,In_1111);
xor U1494 (N_1494,In_1789,In_934);
xnor U1495 (N_1495,In_4342,In_2990);
xnor U1496 (N_1496,In_3928,In_4723);
or U1497 (N_1497,In_52,In_4034);
or U1498 (N_1498,In_1050,In_353);
nand U1499 (N_1499,In_2593,In_3321);
nand U1500 (N_1500,In_1229,In_3881);
nor U1501 (N_1501,In_3251,In_3166);
and U1502 (N_1502,In_4368,In_989);
and U1503 (N_1503,In_182,In_276);
nor U1504 (N_1504,In_1538,In_1090);
and U1505 (N_1505,In_1700,In_4178);
nor U1506 (N_1506,In_4838,In_4005);
or U1507 (N_1507,In_548,In_407);
or U1508 (N_1508,In_518,In_4318);
and U1509 (N_1509,In_812,In_2853);
xnor U1510 (N_1510,In_1134,In_2495);
nor U1511 (N_1511,In_2034,In_1344);
nand U1512 (N_1512,In_1874,In_2606);
nand U1513 (N_1513,In_3653,In_3882);
and U1514 (N_1514,In_3564,In_2446);
or U1515 (N_1515,In_328,In_3824);
nand U1516 (N_1516,In_3196,In_176);
xnor U1517 (N_1517,In_2107,In_3027);
and U1518 (N_1518,In_1457,In_4734);
nand U1519 (N_1519,In_3441,In_64);
nor U1520 (N_1520,In_3921,In_2088);
xor U1521 (N_1521,In_2477,In_4910);
xor U1522 (N_1522,In_4014,In_1597);
nand U1523 (N_1523,In_4260,In_1989);
nand U1524 (N_1524,In_3146,In_3815);
or U1525 (N_1525,In_3486,In_4934);
nor U1526 (N_1526,In_4999,In_2060);
and U1527 (N_1527,In_4979,In_853);
xnor U1528 (N_1528,In_1835,In_3124);
and U1529 (N_1529,In_3485,In_256);
or U1530 (N_1530,In_3449,In_4302);
xor U1531 (N_1531,In_4213,In_2055);
and U1532 (N_1532,In_3442,In_3141);
xnor U1533 (N_1533,In_3772,In_632);
or U1534 (N_1534,In_2279,In_1772);
nand U1535 (N_1535,In_449,In_1308);
nand U1536 (N_1536,In_549,In_1953);
nor U1537 (N_1537,In_746,In_3667);
nand U1538 (N_1538,In_1717,In_4782);
and U1539 (N_1539,In_2082,In_772);
xnor U1540 (N_1540,In_543,In_4491);
xnor U1541 (N_1541,In_3805,In_1763);
nor U1542 (N_1542,In_4224,In_3353);
nor U1543 (N_1543,In_4272,In_3615);
nor U1544 (N_1544,In_3583,In_3566);
nand U1545 (N_1545,In_3089,In_2791);
and U1546 (N_1546,In_2,In_2262);
nand U1547 (N_1547,In_2701,In_1100);
xor U1548 (N_1548,In_4079,In_2626);
or U1549 (N_1549,In_1622,In_1341);
or U1550 (N_1550,In_2347,In_3247);
nor U1551 (N_1551,In_1801,In_1149);
nand U1552 (N_1552,In_2525,In_2572);
nand U1553 (N_1553,In_2868,In_1861);
nor U1554 (N_1554,In_4740,In_2154);
or U1555 (N_1555,In_4105,In_1150);
nand U1556 (N_1556,In_770,In_3150);
nor U1557 (N_1557,In_3889,In_3129);
nor U1558 (N_1558,In_848,In_2290);
xnor U1559 (N_1559,In_3637,In_1822);
nand U1560 (N_1560,In_2846,In_4939);
nand U1561 (N_1561,In_2509,In_1041);
and U1562 (N_1562,In_2101,In_3735);
nor U1563 (N_1563,In_1620,In_2813);
xnor U1564 (N_1564,In_156,In_2011);
or U1565 (N_1565,In_2879,In_1267);
nor U1566 (N_1566,In_166,In_2242);
xor U1567 (N_1567,In_3616,In_2536);
and U1568 (N_1568,In_28,In_2986);
xor U1569 (N_1569,In_4993,In_70);
nor U1570 (N_1570,In_3207,In_567);
nor U1571 (N_1571,In_3516,In_3035);
and U1572 (N_1572,In_3767,In_4736);
or U1573 (N_1573,In_169,In_4419);
xor U1574 (N_1574,In_1782,In_3077);
xor U1575 (N_1575,In_764,In_2208);
nand U1576 (N_1576,In_3159,In_4437);
xnor U1577 (N_1577,In_3774,In_3706);
nor U1578 (N_1578,In_2391,In_4032);
nand U1579 (N_1579,In_1186,In_3465);
nor U1580 (N_1580,In_223,In_702);
and U1581 (N_1581,In_2962,In_1737);
nor U1582 (N_1582,In_2319,In_285);
xnor U1583 (N_1583,In_1433,In_4575);
nand U1584 (N_1584,In_3299,In_2478);
or U1585 (N_1585,In_1461,In_3602);
nand U1586 (N_1586,In_191,In_309);
nand U1587 (N_1587,In_996,In_1070);
nor U1588 (N_1588,In_4833,In_1722);
nor U1589 (N_1589,In_4315,In_3417);
and U1590 (N_1590,In_3236,In_1661);
or U1591 (N_1591,In_4091,In_4691);
xor U1592 (N_1592,In_1960,In_244);
xor U1593 (N_1593,In_3808,In_4579);
nor U1594 (N_1594,In_295,In_62);
and U1595 (N_1595,In_3939,In_4225);
nand U1596 (N_1596,In_1430,In_3919);
and U1597 (N_1597,In_2782,In_1160);
nand U1598 (N_1598,In_3322,In_1943);
nor U1599 (N_1599,In_4244,In_4989);
or U1600 (N_1600,In_893,In_4731);
or U1601 (N_1601,In_454,In_3037);
nor U1602 (N_1602,In_2227,In_3612);
nor U1603 (N_1603,In_3614,In_533);
nand U1604 (N_1604,In_3362,In_3948);
xor U1605 (N_1605,In_3574,In_1490);
and U1606 (N_1606,In_2737,In_1427);
xnor U1607 (N_1607,In_859,In_1588);
nand U1608 (N_1608,In_2300,In_3153);
xnor U1609 (N_1609,In_2769,In_1300);
or U1610 (N_1610,In_4442,In_661);
or U1611 (N_1611,In_123,In_4717);
nor U1612 (N_1612,In_678,In_122);
nand U1613 (N_1613,In_4411,In_3984);
or U1614 (N_1614,In_1773,In_4414);
or U1615 (N_1615,In_4843,In_1014);
nor U1616 (N_1616,In_2739,In_1518);
or U1617 (N_1617,In_4543,In_2952);
xnor U1618 (N_1618,In_147,In_4410);
and U1619 (N_1619,In_1285,In_3300);
or U1620 (N_1620,In_1103,In_3290);
nor U1621 (N_1621,In_4971,In_690);
and U1622 (N_1622,In_3164,In_1076);
nor U1623 (N_1623,In_3890,In_3108);
and U1624 (N_1624,In_4942,In_4450);
xor U1625 (N_1625,In_1680,In_3347);
or U1626 (N_1626,In_1998,In_4771);
nand U1627 (N_1627,In_3699,In_2906);
nor U1628 (N_1628,In_1073,In_1064);
or U1629 (N_1629,In_336,In_1138);
and U1630 (N_1630,In_2095,In_3144);
nor U1631 (N_1631,In_714,In_1435);
and U1632 (N_1632,In_627,In_720);
nand U1633 (N_1633,In_849,In_2820);
or U1634 (N_1634,In_3868,In_2706);
or U1635 (N_1635,In_2267,In_3336);
xnor U1636 (N_1636,In_827,In_4769);
or U1637 (N_1637,In_259,In_57);
xor U1638 (N_1638,In_2654,In_3134);
xnor U1639 (N_1639,In_1650,In_4076);
nand U1640 (N_1640,In_2140,In_954);
and U1641 (N_1641,In_267,In_114);
or U1642 (N_1642,In_3436,In_420);
or U1643 (N_1643,In_3002,In_4878);
or U1644 (N_1644,In_1673,In_649);
and U1645 (N_1645,In_4724,In_660);
and U1646 (N_1646,In_242,In_3042);
nand U1647 (N_1647,In_3852,In_2086);
or U1648 (N_1648,In_1069,In_2858);
xor U1649 (N_1649,In_3901,In_3189);
xor U1650 (N_1650,In_4035,In_4800);
nand U1651 (N_1651,In_666,In_3736);
nor U1652 (N_1652,In_4382,In_1660);
and U1653 (N_1653,In_2462,In_4953);
nor U1654 (N_1654,In_1581,In_1596);
xnor U1655 (N_1655,In_2768,In_1799);
and U1656 (N_1656,In_456,In_1024);
nor U1657 (N_1657,In_4756,In_1841);
or U1658 (N_1658,In_243,In_4803);
xor U1659 (N_1659,In_2102,In_677);
xnor U1660 (N_1660,In_3352,In_1755);
or U1661 (N_1661,In_4489,In_4363);
xnor U1662 (N_1662,In_1689,In_3031);
or U1663 (N_1663,In_1844,In_814);
nor U1664 (N_1664,In_209,In_1561);
nand U1665 (N_1665,In_1302,In_3711);
or U1666 (N_1666,In_2273,In_2907);
xnor U1667 (N_1667,In_1985,In_4184);
or U1668 (N_1668,In_4956,In_3628);
nand U1669 (N_1669,In_4298,In_1849);
nor U1670 (N_1670,In_1909,In_4791);
xnor U1671 (N_1671,In_237,In_2498);
nand U1672 (N_1672,In_1077,In_925);
nand U1673 (N_1673,In_3404,In_1937);
nand U1674 (N_1674,In_4866,In_4559);
xor U1675 (N_1675,In_2240,In_4544);
nand U1676 (N_1676,In_969,In_3454);
nand U1677 (N_1677,In_1044,In_2186);
or U1678 (N_1678,In_4545,In_3464);
nor U1679 (N_1679,In_3753,In_728);
nor U1680 (N_1680,In_2623,In_2698);
or U1681 (N_1681,In_4002,In_3400);
nor U1682 (N_1682,In_2650,In_2276);
nand U1683 (N_1683,In_3800,In_3387);
nand U1684 (N_1684,In_1787,In_90);
xor U1685 (N_1685,In_2648,In_1386);
and U1686 (N_1686,In_3389,In_2941);
nor U1687 (N_1687,In_2038,In_4535);
nand U1688 (N_1688,In_3743,In_4525);
nor U1689 (N_1689,In_2079,In_4011);
nor U1690 (N_1690,In_1557,In_4327);
nor U1691 (N_1691,In_4522,In_4400);
and U1692 (N_1692,In_270,In_2671);
xnor U1693 (N_1693,In_3371,In_3547);
or U1694 (N_1694,In_3151,In_3170);
nand U1695 (N_1695,In_1279,In_2824);
nor U1696 (N_1696,In_689,In_3212);
xnor U1697 (N_1697,In_2704,In_1359);
nor U1698 (N_1698,In_1964,In_1491);
or U1699 (N_1699,In_2470,In_2512);
nor U1700 (N_1700,In_3832,In_4547);
nand U1701 (N_1701,In_397,In_1526);
nand U1702 (N_1702,In_4990,In_1664);
xnor U1703 (N_1703,In_74,In_4357);
and U1704 (N_1704,In_2830,In_729);
nor U1705 (N_1705,In_2936,In_443);
nor U1706 (N_1706,In_3200,In_1545);
xor U1707 (N_1707,In_2258,In_4735);
or U1708 (N_1708,In_1927,In_2457);
and U1709 (N_1709,In_1203,In_3064);
xnor U1710 (N_1710,In_3041,In_1589);
nor U1711 (N_1711,In_2050,In_3867);
nor U1712 (N_1712,In_4493,In_1324);
and U1713 (N_1713,In_3943,In_2058);
or U1714 (N_1714,In_667,In_337);
or U1715 (N_1715,In_1651,In_3331);
or U1716 (N_1716,In_312,In_4948);
xnor U1717 (N_1717,In_2143,In_3610);
or U1718 (N_1718,In_3635,In_2557);
or U1719 (N_1719,In_91,In_1370);
nor U1720 (N_1720,In_875,In_4722);
xnor U1721 (N_1721,In_4943,In_4743);
nor U1722 (N_1722,In_3809,In_2144);
nand U1723 (N_1723,In_3956,In_3403);
and U1724 (N_1724,In_2621,In_929);
and U1725 (N_1725,In_4798,In_2338);
and U1726 (N_1726,In_4533,In_4556);
nor U1727 (N_1727,In_3762,In_4810);
or U1728 (N_1728,In_4918,In_2180);
and U1729 (N_1729,In_1666,In_34);
and U1730 (N_1730,In_613,In_946);
xor U1731 (N_1731,In_3847,In_1246);
xnor U1732 (N_1732,In_3489,In_110);
and U1733 (N_1733,In_2558,In_3611);
nor U1734 (N_1734,In_2972,In_158);
nor U1735 (N_1735,In_2472,In_179);
nand U1736 (N_1736,In_1510,In_4306);
or U1737 (N_1737,In_3607,In_2414);
or U1738 (N_1738,In_2317,In_626);
and U1739 (N_1739,In_601,In_412);
and U1740 (N_1740,In_2194,In_2069);
nand U1741 (N_1741,In_3287,In_1226);
nor U1742 (N_1742,In_4175,In_2543);
or U1743 (N_1743,In_1675,In_512);
or U1744 (N_1744,In_985,In_965);
and U1745 (N_1745,In_372,In_2325);
nor U1746 (N_1746,In_4320,In_2722);
and U1747 (N_1747,In_2253,In_4234);
or U1748 (N_1748,In_943,In_3472);
and U1749 (N_1749,In_3601,In_1777);
nor U1750 (N_1750,In_3857,In_3641);
nand U1751 (N_1751,In_358,In_2728);
or U1752 (N_1752,In_4,In_1319);
and U1753 (N_1753,In_4374,In_1365);
and U1754 (N_1754,In_686,In_1208);
xor U1755 (N_1755,In_3746,In_3539);
nor U1756 (N_1756,In_542,In_4180);
and U1757 (N_1757,In_836,In_55);
nand U1758 (N_1758,In_3572,In_3231);
and U1759 (N_1759,In_3599,In_2743);
and U1760 (N_1760,In_2810,In_4389);
xor U1761 (N_1761,In_157,In_586);
or U1762 (N_1762,In_3491,In_171);
and U1763 (N_1763,In_1484,In_3923);
nand U1764 (N_1764,In_2243,In_1824);
xnor U1765 (N_1765,In_2925,In_3450);
nor U1766 (N_1766,In_3557,In_3103);
nor U1767 (N_1767,In_125,In_3579);
and U1768 (N_1768,In_679,In_2201);
or U1769 (N_1769,In_4776,In_1745);
nor U1770 (N_1770,In_435,In_2217);
and U1771 (N_1771,In_317,In_3191);
xnor U1772 (N_1772,In_1168,In_2432);
nor U1773 (N_1773,In_1244,In_968);
nand U1774 (N_1774,In_1015,In_3213);
nor U1775 (N_1775,In_1129,In_4915);
or U1776 (N_1776,In_1497,In_133);
nor U1777 (N_1777,In_1718,In_2534);
nand U1778 (N_1778,In_1144,In_27);
xnor U1779 (N_1779,In_1568,In_4699);
nor U1780 (N_1780,In_464,In_3127);
or U1781 (N_1781,In_826,In_2002);
and U1782 (N_1782,In_3597,In_2590);
or U1783 (N_1783,In_3747,In_1714);
nor U1784 (N_1784,In_2909,In_3916);
nand U1785 (N_1785,In_4795,In_310);
xnor U1786 (N_1786,In_3996,In_2629);
nor U1787 (N_1787,In_1052,In_2328);
and U1788 (N_1788,In_2417,In_3624);
and U1789 (N_1789,In_967,In_3411);
nor U1790 (N_1790,In_140,In_2028);
nand U1791 (N_1791,In_4100,In_1576);
and U1792 (N_1792,In_3235,In_2772);
or U1793 (N_1793,In_2571,In_3319);
and U1794 (N_1794,In_4911,In_1794);
xor U1795 (N_1795,In_1142,In_1818);
nor U1796 (N_1796,In_4698,In_3293);
and U1797 (N_1797,In_2984,In_2533);
nand U1798 (N_1798,In_4888,In_4009);
and U1799 (N_1799,In_3565,In_0);
xor U1800 (N_1800,In_2280,In_2418);
xor U1801 (N_1801,In_3075,In_2944);
and U1802 (N_1802,In_4278,In_3964);
nor U1803 (N_1803,In_3234,In_1710);
or U1804 (N_1804,In_2118,In_4927);
or U1805 (N_1805,In_3655,In_4495);
xnor U1806 (N_1806,In_3204,In_4397);
and U1807 (N_1807,In_3708,In_3807);
nor U1808 (N_1808,In_2645,In_3678);
nand U1809 (N_1809,In_2091,In_2551);
xnor U1810 (N_1810,In_3949,In_1591);
and U1811 (N_1811,In_3542,In_1783);
or U1812 (N_1812,In_239,In_818);
or U1813 (N_1813,In_2690,In_224);
nand U1814 (N_1814,In_3810,In_4126);
and U1815 (N_1815,In_4435,In_335);
or U1816 (N_1816,In_1387,In_4449);
nor U1817 (N_1817,In_313,In_377);
or U1818 (N_1818,In_3294,In_4462);
nor U1819 (N_1819,In_2809,In_4609);
and U1820 (N_1820,In_4598,In_4751);
or U1821 (N_1821,In_4187,In_2885);
nor U1822 (N_1822,In_2700,In_4200);
nand U1823 (N_1823,In_4420,In_4293);
nor U1824 (N_1824,In_3979,In_1017);
and U1825 (N_1825,In_3717,In_2504);
or U1826 (N_1826,In_324,In_1441);
and U1827 (N_1827,In_3216,In_2920);
nor U1828 (N_1828,In_3621,In_2051);
or U1829 (N_1829,In_1022,In_594);
and U1830 (N_1830,In_2544,In_4080);
nand U1831 (N_1831,In_1784,In_1030);
nor U1832 (N_1832,In_211,In_2215);
nand U1833 (N_1833,In_2130,In_1671);
xnor U1834 (N_1834,In_1959,In_3992);
or U1835 (N_1835,In_4538,In_3396);
nor U1836 (N_1836,In_1121,In_2445);
xnor U1837 (N_1837,In_717,In_963);
or U1838 (N_1838,In_3070,In_2176);
or U1839 (N_1839,In_2950,In_2375);
xor U1840 (N_1840,In_4049,In_713);
and U1841 (N_1841,In_2012,In_3429);
or U1842 (N_1842,In_4245,In_4549);
xnor U1843 (N_1843,In_3696,In_2370);
nand U1844 (N_1844,In_1357,In_2702);
and U1845 (N_1845,In_151,In_708);
nor U1846 (N_1846,In_3609,In_2277);
nand U1847 (N_1847,In_616,In_2673);
or U1848 (N_1848,In_75,In_4048);
xor U1849 (N_1849,In_501,In_2371);
xor U1850 (N_1850,In_3326,In_4863);
nand U1851 (N_1851,In_3272,In_2306);
and U1852 (N_1852,In_2872,In_235);
nand U1853 (N_1853,In_1646,In_4964);
or U1854 (N_1854,In_1366,In_3741);
nand U1855 (N_1855,In_1809,In_4591);
xnor U1856 (N_1856,In_2897,In_3732);
or U1857 (N_1857,In_4814,In_3568);
nor U1858 (N_1858,In_1556,In_3173);
xnor U1859 (N_1859,In_11,In_2521);
xnor U1860 (N_1860,In_2156,In_1419);
nand U1861 (N_1861,In_2929,In_1289);
nor U1862 (N_1862,In_1011,In_3662);
nor U1863 (N_1863,In_4043,In_2005);
or U1864 (N_1864,In_739,In_2802);
xor U1865 (N_1865,In_3934,In_2057);
and U1866 (N_1866,In_3742,In_4216);
and U1867 (N_1867,In_592,In_1350);
nor U1868 (N_1868,In_2574,In_2075);
nand U1869 (N_1869,In_3769,In_490);
or U1870 (N_1870,In_2381,In_3963);
nor U1871 (N_1871,In_2070,In_2815);
and U1872 (N_1872,In_641,In_1481);
nand U1873 (N_1873,In_2175,In_1678);
nor U1874 (N_1874,In_2059,In_1251);
xnor U1875 (N_1875,In_2497,In_671);
xnor U1876 (N_1876,In_2995,In_1072);
nor U1877 (N_1877,In_3487,In_1434);
nor U1878 (N_1878,In_1420,In_547);
nor U1879 (N_1879,In_1525,In_461);
nor U1880 (N_1880,In_229,In_3458);
nor U1881 (N_1881,In_3691,In_2838);
or U1882 (N_1882,In_2619,In_387);
or U1883 (N_1883,In_3672,In_2526);
nor U1884 (N_1884,In_1610,In_891);
or U1885 (N_1885,In_3205,In_2974);
nor U1886 (N_1886,In_4643,In_1991);
xor U1887 (N_1887,In_41,In_553);
and U1888 (N_1888,In_4210,In_511);
nand U1889 (N_1889,In_3345,In_1932);
xnor U1890 (N_1890,In_1205,In_4712);
xnor U1891 (N_1891,In_3763,In_819);
nand U1892 (N_1892,In_51,In_3817);
nand U1893 (N_1893,In_1869,In_835);
and U1894 (N_1894,In_899,In_754);
xnor U1895 (N_1895,In_1190,In_1891);
nand U1896 (N_1896,In_2389,In_3049);
nand U1897 (N_1897,In_991,In_230);
nor U1898 (N_1898,In_3962,In_3535);
xnor U1899 (N_1899,In_833,In_1048);
or U1900 (N_1900,In_834,In_3508);
nor U1901 (N_1901,In_1264,In_299);
xor U1902 (N_1902,In_4149,In_2303);
and U1903 (N_1903,In_2020,In_2755);
or U1904 (N_1904,In_4015,In_3702);
xnor U1905 (N_1905,In_1146,In_3883);
and U1906 (N_1906,In_380,In_413);
xnor U1907 (N_1907,In_1670,In_1693);
or U1908 (N_1908,In_727,In_3029);
nor U1909 (N_1909,In_4936,In_4619);
nor U1910 (N_1910,In_2845,In_1973);
nor U1911 (N_1911,In_4976,In_3359);
nand U1912 (N_1912,In_4604,In_3978);
nor U1913 (N_1913,In_3171,In_3263);
and U1914 (N_1914,In_3926,In_640);
xor U1915 (N_1915,In_201,In_484);
xor U1916 (N_1916,In_3368,In_2667);
and U1917 (N_1917,In_603,In_3707);
nand U1918 (N_1918,In_4628,In_3397);
nor U1919 (N_1919,In_1582,In_3801);
or U1920 (N_1920,In_128,In_4360);
nor U1921 (N_1921,In_3700,In_1314);
nor U1922 (N_1922,In_3115,In_3348);
nand U1923 (N_1923,In_2852,In_2393);
nand U1924 (N_1924,In_1915,In_1562);
xor U1925 (N_1925,In_663,In_631);
nor U1926 (N_1926,In_4962,In_2958);
or U1927 (N_1927,In_222,In_421);
or U1928 (N_1928,In_2209,In_2535);
or U1929 (N_1929,In_2826,In_3238);
nor U1930 (N_1930,In_2292,In_3452);
nor U1931 (N_1931,In_249,In_3181);
nand U1932 (N_1932,In_71,In_2487);
nor U1933 (N_1933,In_809,In_2326);
nor U1934 (N_1934,In_1754,In_674);
xnor U1935 (N_1935,In_4646,In_399);
or U1936 (N_1936,In_1001,In_718);
nand U1937 (N_1937,In_2304,In_1379);
and U1938 (N_1938,In_3622,In_3483);
and U1939 (N_1939,In_2174,In_4568);
xor U1940 (N_1940,In_1373,In_3100);
and U1941 (N_1941,In_1163,In_3155);
nor U1942 (N_1942,In_1301,In_3755);
xor U1943 (N_1943,In_97,In_2947);
nor U1944 (N_1944,In_1303,In_1380);
nand U1945 (N_1945,In_3310,In_1384);
nand U1946 (N_1946,In_3132,In_3082);
or U1947 (N_1947,In_4981,In_2321);
or U1948 (N_1948,In_1060,In_351);
nor U1949 (N_1949,In_957,In_2924);
nand U1950 (N_1950,In_1724,In_2508);
and U1951 (N_1951,In_3544,In_3675);
xnor U1952 (N_1952,In_2783,In_92);
and U1953 (N_1953,In_3744,In_1148);
or U1954 (N_1954,In_2620,In_4138);
nand U1955 (N_1955,In_1768,In_2519);
nand U1956 (N_1956,In_4612,In_744);
or U1957 (N_1957,In_4322,In_2017);
and U1958 (N_1958,In_921,In_3980);
or U1959 (N_1959,In_4426,In_4477);
nand U1960 (N_1960,In_148,In_2837);
xor U1961 (N_1961,In_1521,In_825);
nor U1962 (N_1962,In_2934,In_2881);
and U1963 (N_1963,In_1418,In_4122);
or U1964 (N_1964,In_3502,In_3505);
nor U1965 (N_1965,In_4132,In_1174);
nand U1966 (N_1966,In_4086,In_4807);
nor U1967 (N_1967,In_1290,In_3446);
or U1968 (N_1968,In_4529,In_2349);
xnor U1969 (N_1969,In_806,In_1941);
and U1970 (N_1970,In_3765,In_2951);
xnor U1971 (N_1971,In_4992,In_3357);
or U1972 (N_1972,In_1087,In_4455);
and U1973 (N_1973,In_300,In_10);
nor U1974 (N_1974,In_3327,In_2455);
nand U1975 (N_1975,In_682,In_2094);
nand U1976 (N_1976,In_982,In_590);
nand U1977 (N_1977,In_1107,In_1096);
nor U1978 (N_1978,In_2047,In_356);
nor U1979 (N_1979,In_3532,In_4887);
nor U1980 (N_1980,In_1608,In_3725);
or U1981 (N_1981,In_1377,In_4569);
nor U1982 (N_1982,In_1944,In_21);
or U1983 (N_1983,In_481,In_2541);
nand U1984 (N_1984,In_346,In_4870);
and U1985 (N_1985,In_1157,In_3490);
nor U1986 (N_1986,In_3642,In_1364);
nand U1987 (N_1987,In_4689,In_2866);
nand U1988 (N_1988,In_2678,In_3954);
nor U1989 (N_1989,In_4871,In_297);
nand U1990 (N_1990,In_4093,In_3831);
or U1991 (N_1991,In_314,In_3522);
nor U1992 (N_1992,In_873,In_3306);
nor U1993 (N_1993,In_378,In_2847);
xor U1994 (N_1994,In_4786,In_1448);
and U1995 (N_1995,In_4377,In_2588);
nand U1996 (N_1996,In_1065,In_1431);
or U1997 (N_1997,In_4487,In_3651);
nand U1998 (N_1998,In_796,In_4085);
and U1999 (N_1999,In_3644,In_1594);
xor U2000 (N_2000,In_3538,In_4353);
and U2001 (N_2001,In_1199,In_599);
nor U2002 (N_2002,In_3770,In_272);
nor U2003 (N_2003,In_4084,In_881);
nor U2004 (N_2004,In_69,In_1242);
nor U2005 (N_2005,In_1084,In_3511);
xnor U2006 (N_2006,In_381,In_2741);
xor U2007 (N_2007,In_1713,In_1173);
nor U2008 (N_2008,In_3325,In_2314);
or U2009 (N_2009,In_2877,In_2848);
nand U2010 (N_2010,In_320,In_2324);
nor U2011 (N_2011,In_3870,In_3046);
nor U2012 (N_2012,In_816,In_3424);
or U2013 (N_2013,In_2004,In_3466);
or U2014 (N_2014,In_2615,In_3705);
nor U2015 (N_2015,In_2056,In_4935);
nand U2016 (N_2016,In_2356,In_1876);
and U2017 (N_2017,In_3444,In_2161);
xnor U2018 (N_2018,In_3393,In_364);
or U2019 (N_2019,In_4423,In_250);
or U2020 (N_2020,In_4350,In_3875);
nor U2021 (N_2021,In_1400,In_4155);
nand U2022 (N_2022,In_828,In_246);
and U2023 (N_2023,In_1445,In_3766);
or U2024 (N_2024,In_58,In_4585);
nand U2025 (N_2025,In_1423,In_4111);
or U2026 (N_2026,In_4221,In_1978);
and U2027 (N_2027,In_3749,In_3176);
nand U2028 (N_2028,In_452,In_1278);
nor U2029 (N_2029,In_4745,In_540);
nand U2030 (N_2030,In_1642,In_2265);
and U2031 (N_2031,In_2795,In_352);
xor U2032 (N_2032,In_2404,In_2364);
nor U2033 (N_2033,In_2797,In_273);
nand U2034 (N_2034,In_4711,In_4066);
or U2035 (N_2035,In_1362,In_917);
or U2036 (N_2036,In_4576,In_4196);
xor U2037 (N_2037,In_3914,In_4479);
xor U2038 (N_2038,In_1980,In_1706);
or U2039 (N_2039,In_1196,In_3180);
or U2040 (N_2040,In_2184,In_3304);
nor U2041 (N_2041,In_3302,In_2293);
nor U2042 (N_2042,In_3091,In_1110);
or U2043 (N_2043,In_4325,In_2333);
or U2044 (N_2044,In_2410,In_4969);
nand U2045 (N_2045,In_493,In_1280);
xor U2046 (N_2046,In_654,In_271);
or U2047 (N_2047,In_1972,In_4697);
nor U2048 (N_2048,In_155,In_504);
nand U2049 (N_2049,In_1316,In_1894);
nor U2050 (N_2050,In_1006,In_4912);
xor U2051 (N_2051,In_994,In_4312);
xnor U2052 (N_2052,In_1216,In_4425);
and U2053 (N_2053,In_2160,In_883);
xor U2054 (N_2054,In_2428,In_431);
xnor U2055 (N_2055,In_4137,In_4797);
xor U2056 (N_2056,In_1460,In_624);
xor U2057 (N_2057,In_2153,In_1584);
or U2058 (N_2058,In_3479,In_410);
nand U2059 (N_2059,In_16,In_2188);
nand U2060 (N_2060,In_1575,In_2799);
or U2061 (N_2061,In_2511,In_1522);
nand U2062 (N_2062,In_4827,In_1120);
xnor U2063 (N_2063,In_735,In_759);
nor U2064 (N_2064,In_2803,In_1161);
xor U2065 (N_2065,In_23,In_4755);
nor U2066 (N_2066,In_4238,In_3116);
nor U2067 (N_2067,In_3733,In_3232);
nand U2068 (N_2068,In_2991,In_3384);
and U2069 (N_2069,In_1029,In_108);
nor U2070 (N_2070,In_479,In_3681);
or U2071 (N_2071,In_3210,In_4968);
nand U2072 (N_2072,In_1105,In_3275);
nor U2073 (N_2073,In_4685,In_4634);
xor U2074 (N_2074,In_4790,In_1760);
nand U2075 (N_2075,In_4456,In_2015);
or U2076 (N_2076,In_2278,In_1644);
or U2077 (N_2077,In_2669,In_386);
or U2078 (N_2078,In_699,In_1291);
or U2079 (N_2079,In_2295,In_877);
or U2080 (N_2080,In_4594,In_2413);
xnor U2081 (N_2081,In_2132,In_3761);
nor U2082 (N_2082,In_4690,In_3592);
or U2083 (N_2083,In_3208,In_1215);
and U2084 (N_2084,In_1495,In_3425);
nor U2085 (N_2085,In_472,In_1128);
or U2086 (N_2086,In_2981,In_3669);
xor U2087 (N_2087,In_3849,In_1935);
nand U2088 (N_2088,In_1613,In_4161);
and U2089 (N_2089,In_4167,In_2939);
xor U2090 (N_2090,In_4453,In_2516);
nor U2091 (N_2091,In_940,In_2461);
or U2092 (N_2092,In_3515,In_3097);
nand U2093 (N_2093,In_898,In_2182);
or U2094 (N_2094,In_3617,In_3906);
or U2095 (N_2095,In_2256,In_716);
or U2096 (N_2096,In_4561,In_680);
xnor U2097 (N_2097,In_3125,In_4713);
or U2098 (N_2098,In_3682,In_2751);
nand U2099 (N_2099,In_3927,In_4064);
nor U2100 (N_2100,In_3476,In_2106);
nor U2101 (N_2101,In_1159,In_2888);
and U2102 (N_2102,In_1736,In_3598);
nand U2103 (N_2103,In_745,In_2197);
nor U2104 (N_2104,In_1527,In_741);
xor U2105 (N_2105,In_1136,In_950);
nor U2106 (N_2106,In_4159,In_3540);
xor U2107 (N_2107,In_1428,In_3531);
nor U2108 (N_2108,In_3989,In_3113);
or U2109 (N_2109,In_1816,In_1603);
or U2110 (N_2110,In_4139,In_32);
xor U2111 (N_2111,In_2205,In_1752);
xnor U2112 (N_2112,In_515,In_4983);
nor U2113 (N_2113,In_1880,In_546);
nor U2114 (N_2114,In_787,In_585);
or U2115 (N_2115,In_1520,In_4621);
nor U2116 (N_2116,In_2316,In_980);
nand U2117 (N_2117,In_514,In_4006);
nor U2118 (N_2118,In_2729,In_2796);
nand U2119 (N_2119,In_1307,In_1055);
and U2120 (N_2120,In_634,In_763);
and U2121 (N_2121,In_4052,In_561);
xnor U2122 (N_2122,In_4780,In_2633);
nand U2123 (N_2123,In_3245,In_4872);
nand U2124 (N_2124,In_3119,In_2861);
or U2125 (N_2125,In_4955,In_2363);
or U2126 (N_2126,In_429,In_1340);
and U2127 (N_2127,In_4028,In_2257);
xor U2128 (N_2128,In_3430,In_1957);
nand U2129 (N_2129,In_3799,In_1297);
or U2130 (N_2130,In_1854,In_3311);
and U2131 (N_2131,In_3968,In_4355);
nand U2132 (N_2132,In_4665,In_2655);
nand U2133 (N_2133,In_2444,In_4998);
or U2134 (N_2134,In_3784,In_4113);
nor U2135 (N_2135,In_4893,In_497);
xor U2136 (N_2136,In_2423,In_4616);
nand U2137 (N_2137,In_653,In_4239);
or U2138 (N_2138,In_126,In_2724);
nand U2139 (N_2139,In_2465,In_2987);
nor U2140 (N_2140,In_1917,In_1504);
and U2141 (N_2141,In_2539,In_830);
nor U2142 (N_2142,In_3341,In_2681);
xnor U2143 (N_2143,In_2271,In_1933);
xnor U2144 (N_2144,In_2577,In_1764);
or U2145 (N_2145,In_4657,In_4431);
nor U2146 (N_2146,In_1002,In_4652);
nand U2147 (N_2147,In_4022,In_1018);
nand U2148 (N_2148,In_1047,In_864);
or U2149 (N_2149,In_2078,In_3537);
xor U2150 (N_2150,In_4738,In_526);
nand U2151 (N_2151,In_2851,In_2915);
and U2152 (N_2152,In_2524,In_3139);
nand U2153 (N_2153,In_1934,In_4164);
xnor U2154 (N_2154,In_3271,In_1895);
nor U2155 (N_2155,In_1353,In_1499);
nor U2156 (N_2156,In_4553,In_1508);
nor U2157 (N_2157,In_1408,In_792);
or U2158 (N_2158,In_715,In_3562);
xnor U2159 (N_2159,In_3295,In_694);
and U2160 (N_2160,In_86,In_3806);
and U2161 (N_2161,In_4001,In_4031);
nor U2162 (N_2162,In_2828,In_1753);
and U2163 (N_2163,In_190,In_4296);
and U2164 (N_2164,In_2139,In_576);
nor U2165 (N_2165,In_453,In_4960);
nor U2166 (N_2166,In_4668,In_2890);
and U2167 (N_2167,In_2178,In_684);
nand U2168 (N_2168,In_3764,In_2387);
xor U2169 (N_2169,In_3292,In_976);
xor U2170 (N_2170,In_2084,In_321);
nor U2171 (N_2171,In_3498,In_3350);
nor U2172 (N_2172,In_1899,In_3839);
and U2173 (N_2173,In_3270,In_2695);
nor U2174 (N_2174,In_4059,In_1567);
nand U2175 (N_2175,In_658,In_4270);
xor U2176 (N_2176,In_4447,In_4095);
nor U2177 (N_2177,In_1376,In_3666);
and U2178 (N_2178,In_2740,In_4308);
or U2179 (N_2179,In_1053,In_4853);
nor U2180 (N_2180,In_2510,In_2634);
nor U2181 (N_2181,In_557,In_4633);
and U2182 (N_2182,In_2656,In_4289);
nand U2183 (N_2183,In_470,In_4073);
xor U2184 (N_2184,In_2147,In_2789);
xor U2185 (N_2185,In_2955,In_2323);
nor U2186 (N_2186,In_1459,In_829);
or U2187 (N_2187,In_4907,In_4054);
nand U2188 (N_2188,In_4401,In_1730);
nand U2189 (N_2189,In_4784,In_1287);
and U2190 (N_2190,In_107,In_3918);
and U2191 (N_2191,In_3887,In_1037);
nand U2192 (N_2192,In_4632,In_995);
and U2193 (N_2193,In_4817,In_2758);
or U2194 (N_2194,In_1570,In_3318);
nand U2195 (N_2195,In_3619,In_4812);
xnor U2196 (N_2196,In_707,In_4089);
nor U2197 (N_2197,In_748,In_2723);
xor U2198 (N_2198,In_2074,In_4331);
nor U2199 (N_2199,In_750,In_4417);
and U2200 (N_2200,In_1690,In_228);
or U2201 (N_2201,In_4637,In_4367);
and U2202 (N_2202,In_4375,In_2641);
xor U2203 (N_2203,In_2486,In_2756);
nand U2204 (N_2204,In_161,In_221);
xor U2205 (N_2205,In_445,In_800);
and U2206 (N_2206,In_712,In_4595);
and U2207 (N_2207,In_656,In_3333);
and U2208 (N_2208,In_3248,In_226);
or U2209 (N_2209,In_3440,In_3698);
nand U2210 (N_2210,In_4701,In_1842);
nor U2211 (N_2211,In_701,In_1309);
and U2212 (N_2212,In_4369,In_611);
xnor U2213 (N_2213,In_2092,In_1878);
nand U2214 (N_2214,In_4344,In_2507);
xnor U2215 (N_2215,In_4365,In_1549);
xnor U2216 (N_2216,In_4895,In_502);
xnor U2217 (N_2217,In_3457,In_2914);
or U2218 (N_2218,In_904,In_393);
or U2219 (N_2219,In_96,In_1793);
xor U2220 (N_2220,In_121,In_3748);
or U2221 (N_2221,In_3929,In_278);
or U2222 (N_2222,In_2396,In_2697);
nand U2223 (N_2223,In_4623,In_1982);
xnor U2224 (N_2224,In_4679,In_938);
and U2225 (N_2225,In_600,In_2841);
or U2226 (N_2226,In_743,In_117);
xor U2227 (N_2227,In_2245,In_2171);
nor U2228 (N_2228,In_3530,In_3346);
nor U2229 (N_2229,In_1825,In_651);
and U2230 (N_2230,In_374,In_4109);
and U2231 (N_2231,In_2595,In_1974);
or U2232 (N_2232,In_4112,In_2770);
xor U2233 (N_2233,In_3529,In_4867);
xnor U2234 (N_2234,In_20,In_602);
nand U2235 (N_2235,In_604,In_3067);
or U2236 (N_2236,In_1962,In_997);
and U2237 (N_2237,In_3117,In_3240);
xor U2238 (N_2238,In_1245,In_471);
nor U2239 (N_2239,In_4378,In_345);
xnor U2240 (N_2240,In_3781,In_382);
xor U2241 (N_2241,In_3172,In_2283);
nor U2242 (N_2242,In_4684,In_1797);
nor U2243 (N_2243,In_422,In_4631);
and U2244 (N_2244,In_1025,In_757);
or U2245 (N_2245,In_2777,In_2330);
nor U2246 (N_2246,In_4124,In_2691);
nor U2247 (N_2247,In_2255,In_3715);
or U2248 (N_2248,In_2599,In_2126);
and U2249 (N_2249,In_3069,In_4931);
nand U2250 (N_2250,In_3118,In_2266);
nand U2251 (N_2251,In_1573,In_1778);
nor U2252 (N_2252,In_3312,In_2617);
and U2253 (N_2253,In_3431,In_2029);
nand U2254 (N_2254,In_999,In_3102);
nand U2255 (N_2255,In_325,In_248);
nor U2256 (N_2256,In_1322,In_1892);
nand U2257 (N_2257,In_1796,In_3349);
nor U2258 (N_2258,In_1952,In_1201);
xor U2259 (N_2259,In_2361,In_981);
nand U2260 (N_2260,In_1564,In_2105);
or U2261 (N_2261,In_1189,In_4135);
nor U2262 (N_2262,In_3604,In_4207);
and U2263 (N_2263,In_1756,In_3874);
and U2264 (N_2264,In_2971,In_2196);
nor U2265 (N_2265,In_2529,In_2937);
xnor U2266 (N_2266,In_2732,In_252);
nand U2267 (N_2267,In_46,In_1214);
and U2268 (N_2268,In_1260,In_1537);
nor U2269 (N_2269,In_2836,In_4730);
or U2270 (N_2270,In_2185,In_2407);
and U2271 (N_2271,In_1249,In_3971);
xnor U2272 (N_2272,In_3811,In_1268);
nand U2273 (N_2273,In_1898,In_4874);
and U2274 (N_2274,In_3278,In_194);
nand U2275 (N_2275,In_802,In_1153);
and U2276 (N_2276,In_2427,In_4402);
nor U2277 (N_2277,In_1467,In_1093);
xnor U2278 (N_2278,In_2930,In_1640);
xor U2279 (N_2279,In_737,In_998);
xnor U2280 (N_2280,In_31,In_4460);
or U2281 (N_2281,In_4108,In_1241);
or U2282 (N_2282,In_1042,In_1572);
and U2283 (N_2283,In_2013,In_1451);
xnor U2284 (N_2284,In_2121,In_2115);
nand U2285 (N_2285,In_1501,In_1819);
or U2286 (N_2286,In_1292,In_2898);
xor U2287 (N_2287,In_2787,In_1954);
nor U2288 (N_2288,In_2880,In_175);
nor U2289 (N_2289,In_368,In_2016);
nor U2290 (N_2290,In_2807,In_1715);
nand U2291 (N_2291,In_4269,In_3780);
nand U2292 (N_2292,In_1440,In_1293);
and U2293 (N_2293,In_4201,In_1536);
nand U2294 (N_2294,In_1920,In_4267);
and U2295 (N_2295,In_4674,In_1904);
nor U2296 (N_2296,In_3010,In_3071);
or U2297 (N_2297,In_1363,In_2221);
nand U2298 (N_2298,In_13,In_2560);
and U2299 (N_2299,In_2112,In_906);
nor U2300 (N_2300,In_3858,In_1741);
or U2301 (N_2301,In_2856,In_4560);
and U2302 (N_2302,In_4626,In_3967);
xor U2303 (N_2303,In_4531,In_2513);
or U2304 (N_2304,In_3026,In_1485);
or U2305 (N_2305,In_183,In_3372);
or U2306 (N_2306,In_1931,In_3649);
xor U2307 (N_2307,In_4454,In_4168);
or U2308 (N_2308,In_2996,In_4075);
and U2309 (N_2309,In_4399,In_1617);
nor U2310 (N_2310,In_2008,In_42);
and U2311 (N_2311,In_3226,In_131);
xor U2312 (N_2312,In_1482,In_2202);
nor U2313 (N_2313,In_33,In_2373);
xnor U2314 (N_2314,In_2198,In_597);
nand U2315 (N_2315,In_3257,In_612);
nand U2316 (N_2316,In_3924,In_2048);
or U2317 (N_2317,In_3719,In_4394);
or U2318 (N_2318,In_4686,In_4082);
nor U2319 (N_2319,In_2235,In_935);
xor U2320 (N_2320,In_2625,In_3885);
xor U2321 (N_2321,In_3376,In_4914);
xnor U2322 (N_2322,In_4020,In_139);
nand U2323 (N_2323,In_747,In_962);
or U2324 (N_2324,In_298,In_213);
and U2325 (N_2325,In_4467,In_911);
nor U2326 (N_2326,In_2190,In_1820);
nand U2327 (N_2327,In_4362,In_2715);
and U2328 (N_2328,In_3552,In_1612);
and U2329 (N_2329,In_2618,In_4714);
nand U2330 (N_2330,In_862,In_4459);
and U2331 (N_2331,In_3178,In_475);
nor U2332 (N_2332,In_60,In_405);
or U2333 (N_2333,In_6,In_1560);
and U2334 (N_2334,In_4625,In_958);
or U2335 (N_2335,In_2453,In_724);
nand U2336 (N_2336,In_2100,In_2757);
xnor U2337 (N_2337,In_2448,In_2765);
nor U2338 (N_2338,In_2122,In_3162);
or U2339 (N_2339,In_3745,In_2892);
nor U2340 (N_2340,In_3413,In_4845);
nand U2341 (N_2341,In_780,In_3975);
xnor U2342 (N_2342,In_539,In_3237);
xnor U2343 (N_2343,In_2438,In_3280);
xor U2344 (N_2344,In_3703,In_643);
nor U2345 (N_2345,In_4434,In_3664);
and U2346 (N_2346,In_3888,In_4240);
or U2347 (N_2347,In_4326,In_2125);
xnor U2348 (N_2348,In_4985,In_4639);
and U2349 (N_2349,In_1265,In_4183);
xor U2350 (N_2350,In_2093,In_2835);
xnor U2351 (N_2351,In_165,In_1349);
and U2352 (N_2352,In_1618,In_4865);
nand U2353 (N_2353,In_3095,In_520);
nor U2354 (N_2354,In_1523,In_1630);
nand U2355 (N_2355,In_39,In_2203);
xnor U2356 (N_2356,In_2187,In_4541);
nand U2357 (N_2357,In_4677,In_366);
nand U2358 (N_2358,In_3463,In_2152);
and U2359 (N_2359,In_4572,In_761);
or U2360 (N_2360,In_2960,In_2717);
xor U2361 (N_2361,In_268,In_2979);
nor U2362 (N_2362,In_2973,In_2467);
nor U2363 (N_2363,In_2568,In_1405);
nor U2364 (N_2364,In_3859,In_4564);
xnor U2365 (N_2365,In_1049,In_2189);
nand U2366 (N_2366,In_3047,In_4515);
and U2367 (N_2367,In_2873,In_3823);
xor U2368 (N_2368,In_617,In_807);
nor U2369 (N_2369,In_1010,In_1125);
xnor U2370 (N_2370,In_424,In_1003);
nor U2371 (N_2371,In_992,In_1949);
xor U2372 (N_2372,In_2744,In_3096);
and U2373 (N_2373,In_1627,In_4366);
xor U2374 (N_2374,In_3533,In_1411);
nand U2375 (N_2375,In_43,In_3382);
nor U2376 (N_2376,In_1913,In_3036);
xor U2377 (N_2377,In_2072,In_218);
xnor U2378 (N_2378,In_1312,In_3710);
nand U2379 (N_2379,In_3595,In_1672);
nor U2380 (N_2380,In_1193,In_2640);
nor U2381 (N_2381,In_4145,In_1786);
or U2382 (N_2382,In_1840,In_1911);
nor U2383 (N_2383,In_4546,In_3626);
or U2384 (N_2384,In_2865,In_3201);
nor U2385 (N_2385,In_2421,In_3088);
and U2386 (N_2386,In_3008,In_3970);
nor U2387 (N_2387,In_1356,In_4226);
nand U2388 (N_2388,In_2935,In_869);
and U2389 (N_2389,In_3777,In_1720);
xor U2390 (N_2390,In_3802,In_2631);
nand U2391 (N_2391,In_3794,In_2814);
and U2392 (N_2392,In_2808,In_2540);
nand U2393 (N_2393,In_4824,In_308);
nor U2394 (N_2394,In_340,In_4815);
or U2395 (N_2395,In_1325,In_487);
nand U2396 (N_2396,In_1250,In_2199);
nor U2397 (N_2397,In_3004,In_465);
nor U2398 (N_2398,In_2908,In_618);
and U2399 (N_2399,In_4230,In_208);
xnor U2400 (N_2400,In_4673,In_2284);
nor U2401 (N_2401,In_3093,In_3768);
nand U2402 (N_2402,In_3841,In_3917);
or U2403 (N_2403,In_1124,In_4857);
or U2404 (N_2404,In_167,In_2546);
nand U2405 (N_2405,In_1021,In_2760);
nand U2406 (N_2406,In_4851,In_2883);
nor U2407 (N_2407,In_3330,In_4471);
xnor U2408 (N_2408,In_2522,In_890);
and U2409 (N_2409,In_2579,In_1781);
nand U2410 (N_2410,In_1930,In_2682);
nor U2411 (N_2411,In_1004,In_3783);
nor U2412 (N_2412,In_941,In_4768);
nor U2413 (N_2413,In_357,In_4614);
xor U2414 (N_2414,In_1471,In_4017);
nor U2415 (N_2415,In_3255,In_4220);
nor U2416 (N_2416,In_4508,In_304);
and U2417 (N_2417,In_3937,In_1239);
xor U2418 (N_2418,In_4232,In_4821);
and U2419 (N_2419,In_2692,In_1918);
and U2420 (N_2420,In_105,In_2563);
nor U2421 (N_2421,In_1390,In_2169);
or U2422 (N_2422,In_726,In_843);
or U2423 (N_2423,In_4516,In_1848);
nand U2424 (N_2424,In_1558,In_488);
nand U2425 (N_2425,In_1587,In_1209);
and U2426 (N_2426,In_4058,In_4925);
or U2427 (N_2427,In_4656,In_1466);
or U2428 (N_2428,In_4166,In_2871);
nor U2429 (N_2429,In_3335,In_269);
xnor U2430 (N_2430,In_4641,In_2781);
or U2431 (N_2431,In_2289,In_2113);
xor U2432 (N_2432,In_4346,In_2731);
and U2433 (N_2433,In_1355,In_1487);
nand U2434 (N_2434,In_896,In_2309);
nor U2435 (N_2435,In_3249,In_3804);
xor U2436 (N_2436,In_4881,In_4068);
xnor U2437 (N_2437,In_1410,In_2580);
or U2438 (N_2438,In_341,In_4263);
and U2439 (N_2439,In_2150,In_1156);
nor U2440 (N_2440,In_1771,In_362);
nor U2441 (N_2441,In_1798,In_3782);
xnor U2442 (N_2442,In_1228,In_274);
xnor U2443 (N_2443,In_1211,In_113);
nor U2444 (N_2444,In_3122,In_4806);
or U2445 (N_2445,In_1766,In_2614);
xnor U2446 (N_2446,In_3640,In_2685);
xor U2447 (N_2447,In_1827,In_4370);
or U2448 (N_2448,In_1569,In_3101);
nand U2449 (N_2449,In_1039,In_1800);
xnor U2450 (N_2450,In_3588,In_593);
nor U2451 (N_2451,In_2842,In_2298);
and U2452 (N_2452,In_4659,In_2567);
and U2453 (N_2453,In_4409,In_1616);
nand U2454 (N_2454,In_1449,In_3195);
xnor U2455 (N_2455,In_2506,In_1233);
xor U2456 (N_2456,In_797,In_473);
xor U2457 (N_2457,In_2167,In_4203);
nand U2458 (N_2458,In_83,In_1856);
xnor U2459 (N_2459,In_332,In_867);
xnor U2460 (N_2460,In_1774,In_319);
or U2461 (N_2461,In_2419,In_44);
and U2462 (N_2462,In_3421,In_4185);
and U2463 (N_2463,In_3570,In_4883);
and U2464 (N_2464,In_988,In_2260);
nor U2465 (N_2465,In_446,In_4393);
nand U2466 (N_2466,In_418,In_2313);
and U2467 (N_2467,In_2779,In_4645);
and U2468 (N_2468,In_2752,In_283);
xor U2469 (N_2469,In_2340,In_3229);
or U2470 (N_2470,In_72,In_3473);
nor U2471 (N_2471,In_1685,In_2270);
nor U2472 (N_2472,In_2491,In_3193);
nor U2473 (N_2473,In_203,In_1541);
nor U2474 (N_2474,In_4019,In_2026);
nand U2475 (N_2475,In_1375,In_851);
nor U2476 (N_2476,In_1604,In_532);
xnor U2477 (N_2477,In_2003,In_4527);
xor U2478 (N_2478,In_3414,In_4314);
nor U2479 (N_2479,In_837,In_1135);
nor U2480 (N_2480,In_1346,In_3701);
nand U2481 (N_2481,In_964,In_4345);
nand U2482 (N_2482,In_4324,In_48);
xnor U2483 (N_2483,In_919,In_2867);
nand U2484 (N_2484,In_1940,In_731);
nand U2485 (N_2485,In_1695,In_4339);
nand U2486 (N_2486,In_856,In_2517);
nor U2487 (N_2487,In_2945,In_554);
nand U2488 (N_2488,In_419,In_4662);
and U2489 (N_2489,In_2435,In_799);
nor U2490 (N_2490,In_3252,In_1684);
and U2491 (N_2491,In_1412,In_673);
nand U2492 (N_2492,In_2179,In_2684);
and U2493 (N_2493,In_3940,In_1224);
nor U2494 (N_2494,In_1663,In_1631);
nor U2495 (N_2495,In_478,In_1179);
nand U2496 (N_2496,In_4047,In_4524);
nor U2497 (N_2497,In_1336,In_4906);
or U2498 (N_2498,In_3283,In_1258);
or U2499 (N_2499,In_4642,In_527);
nand U2500 (N_2500,In_3927,In_2074);
and U2501 (N_2501,In_4631,In_3894);
and U2502 (N_2502,In_2874,In_4671);
nand U2503 (N_2503,In_639,In_612);
xnor U2504 (N_2504,In_2871,In_2000);
or U2505 (N_2505,In_4772,In_3958);
xnor U2506 (N_2506,In_4603,In_50);
or U2507 (N_2507,In_1702,In_1428);
or U2508 (N_2508,In_548,In_4942);
or U2509 (N_2509,In_3234,In_2382);
xnor U2510 (N_2510,In_2829,In_643);
nor U2511 (N_2511,In_2145,In_4129);
and U2512 (N_2512,In_4260,In_1635);
nand U2513 (N_2513,In_2569,In_3028);
xor U2514 (N_2514,In_4610,In_983);
nand U2515 (N_2515,In_1556,In_1248);
or U2516 (N_2516,In_2556,In_2397);
or U2517 (N_2517,In_2864,In_4850);
nand U2518 (N_2518,In_2372,In_965);
xnor U2519 (N_2519,In_2225,In_127);
xor U2520 (N_2520,In_2590,In_1719);
xnor U2521 (N_2521,In_4314,In_4003);
nand U2522 (N_2522,In_1970,In_660);
xor U2523 (N_2523,In_481,In_1908);
nand U2524 (N_2524,In_3478,In_1575);
nor U2525 (N_2525,In_907,In_2552);
nand U2526 (N_2526,In_3758,In_3786);
nor U2527 (N_2527,In_1615,In_2599);
and U2528 (N_2528,In_1818,In_1754);
xor U2529 (N_2529,In_3112,In_1594);
nand U2530 (N_2530,In_3799,In_4001);
and U2531 (N_2531,In_1796,In_1265);
nor U2532 (N_2532,In_690,In_747);
xor U2533 (N_2533,In_4470,In_303);
nand U2534 (N_2534,In_2842,In_3127);
nor U2535 (N_2535,In_1169,In_3560);
and U2536 (N_2536,In_4185,In_4866);
nor U2537 (N_2537,In_2181,In_2542);
nor U2538 (N_2538,In_2963,In_982);
nand U2539 (N_2539,In_1262,In_2154);
xnor U2540 (N_2540,In_605,In_4594);
or U2541 (N_2541,In_537,In_4589);
nor U2542 (N_2542,In_4347,In_3760);
and U2543 (N_2543,In_1409,In_3498);
nand U2544 (N_2544,In_3075,In_2060);
xnor U2545 (N_2545,In_4544,In_783);
and U2546 (N_2546,In_4602,In_4615);
xor U2547 (N_2547,In_3998,In_397);
or U2548 (N_2548,In_372,In_145);
xnor U2549 (N_2549,In_3238,In_390);
xor U2550 (N_2550,In_3792,In_494);
nor U2551 (N_2551,In_2243,In_411);
xor U2552 (N_2552,In_3351,In_4679);
and U2553 (N_2553,In_2332,In_215);
and U2554 (N_2554,In_4064,In_3597);
and U2555 (N_2555,In_4269,In_4723);
nand U2556 (N_2556,In_4271,In_4186);
xnor U2557 (N_2557,In_4052,In_1270);
nand U2558 (N_2558,In_2982,In_4811);
or U2559 (N_2559,In_3718,In_637);
and U2560 (N_2560,In_1500,In_925);
or U2561 (N_2561,In_104,In_4328);
xor U2562 (N_2562,In_4846,In_2062);
and U2563 (N_2563,In_2756,In_1126);
xor U2564 (N_2564,In_1222,In_4406);
or U2565 (N_2565,In_4490,In_514);
or U2566 (N_2566,In_4103,In_3368);
or U2567 (N_2567,In_2558,In_1210);
or U2568 (N_2568,In_3836,In_384);
nor U2569 (N_2569,In_340,In_3419);
or U2570 (N_2570,In_3168,In_2907);
or U2571 (N_2571,In_3553,In_3819);
and U2572 (N_2572,In_4806,In_3200);
nor U2573 (N_2573,In_1682,In_1852);
nand U2574 (N_2574,In_4054,In_820);
xnor U2575 (N_2575,In_1594,In_4963);
and U2576 (N_2576,In_628,In_4116);
xnor U2577 (N_2577,In_2703,In_4116);
xnor U2578 (N_2578,In_2906,In_4850);
xnor U2579 (N_2579,In_2670,In_4497);
or U2580 (N_2580,In_4648,In_1373);
and U2581 (N_2581,In_662,In_1465);
and U2582 (N_2582,In_1919,In_2847);
or U2583 (N_2583,In_1432,In_4748);
nand U2584 (N_2584,In_3278,In_830);
nand U2585 (N_2585,In_3895,In_1257);
nand U2586 (N_2586,In_2112,In_2127);
and U2587 (N_2587,In_132,In_4452);
nor U2588 (N_2588,In_48,In_165);
or U2589 (N_2589,In_946,In_473);
nand U2590 (N_2590,In_3199,In_3866);
nand U2591 (N_2591,In_2943,In_1552);
nand U2592 (N_2592,In_443,In_2026);
or U2593 (N_2593,In_833,In_562);
xnor U2594 (N_2594,In_2252,In_662);
nand U2595 (N_2595,In_2873,In_4354);
nand U2596 (N_2596,In_3535,In_2769);
and U2597 (N_2597,In_4541,In_863);
or U2598 (N_2598,In_642,In_384);
or U2599 (N_2599,In_4307,In_4624);
and U2600 (N_2600,In_3838,In_2034);
xnor U2601 (N_2601,In_1861,In_78);
or U2602 (N_2602,In_3729,In_4230);
and U2603 (N_2603,In_388,In_2634);
xnor U2604 (N_2604,In_1561,In_1872);
or U2605 (N_2605,In_3798,In_4166);
xnor U2606 (N_2606,In_2413,In_2647);
nor U2607 (N_2607,In_37,In_2650);
and U2608 (N_2608,In_4429,In_212);
nor U2609 (N_2609,In_489,In_2724);
xor U2610 (N_2610,In_295,In_2376);
nand U2611 (N_2611,In_2191,In_4429);
nor U2612 (N_2612,In_2778,In_64);
or U2613 (N_2613,In_1158,In_3799);
or U2614 (N_2614,In_1172,In_705);
xnor U2615 (N_2615,In_747,In_710);
or U2616 (N_2616,In_2984,In_1317);
and U2617 (N_2617,In_3724,In_1579);
nor U2618 (N_2618,In_4974,In_2485);
nor U2619 (N_2619,In_4049,In_1445);
nor U2620 (N_2620,In_4081,In_3881);
nand U2621 (N_2621,In_2111,In_4081);
nor U2622 (N_2622,In_1247,In_1954);
xor U2623 (N_2623,In_1709,In_1565);
and U2624 (N_2624,In_1217,In_4093);
nand U2625 (N_2625,In_1840,In_3401);
nand U2626 (N_2626,In_1258,In_738);
and U2627 (N_2627,In_690,In_3880);
or U2628 (N_2628,In_1780,In_1272);
nor U2629 (N_2629,In_2384,In_4536);
nand U2630 (N_2630,In_1945,In_4340);
xnor U2631 (N_2631,In_1672,In_1921);
nor U2632 (N_2632,In_4846,In_2159);
xor U2633 (N_2633,In_2303,In_911);
or U2634 (N_2634,In_2730,In_3359);
nand U2635 (N_2635,In_3270,In_1724);
xor U2636 (N_2636,In_381,In_1035);
nand U2637 (N_2637,In_2930,In_4817);
nand U2638 (N_2638,In_2639,In_1614);
and U2639 (N_2639,In_4797,In_674);
and U2640 (N_2640,In_700,In_2320);
xor U2641 (N_2641,In_980,In_683);
nor U2642 (N_2642,In_1781,In_3249);
nand U2643 (N_2643,In_4209,In_1395);
or U2644 (N_2644,In_4159,In_238);
nor U2645 (N_2645,In_2689,In_1678);
xnor U2646 (N_2646,In_1765,In_3714);
nand U2647 (N_2647,In_57,In_2354);
nor U2648 (N_2648,In_4075,In_4066);
nor U2649 (N_2649,In_1516,In_874);
or U2650 (N_2650,In_3143,In_3396);
xor U2651 (N_2651,In_585,In_998);
or U2652 (N_2652,In_4656,In_3692);
nand U2653 (N_2653,In_4635,In_4961);
xnor U2654 (N_2654,In_4887,In_4713);
nand U2655 (N_2655,In_1564,In_1234);
nor U2656 (N_2656,In_1913,In_2410);
or U2657 (N_2657,In_4096,In_1995);
or U2658 (N_2658,In_1292,In_1529);
nand U2659 (N_2659,In_4831,In_987);
xor U2660 (N_2660,In_3463,In_1783);
nor U2661 (N_2661,In_2518,In_3184);
and U2662 (N_2662,In_3119,In_394);
and U2663 (N_2663,In_3276,In_1491);
xnor U2664 (N_2664,In_1489,In_1872);
nand U2665 (N_2665,In_2109,In_1245);
nor U2666 (N_2666,In_1304,In_2421);
or U2667 (N_2667,In_4260,In_2430);
and U2668 (N_2668,In_2861,In_1759);
nor U2669 (N_2669,In_424,In_3922);
and U2670 (N_2670,In_588,In_4973);
nand U2671 (N_2671,In_3614,In_4427);
and U2672 (N_2672,In_297,In_1794);
and U2673 (N_2673,In_3791,In_2979);
or U2674 (N_2674,In_720,In_3058);
or U2675 (N_2675,In_4122,In_4879);
nand U2676 (N_2676,In_1380,In_3746);
and U2677 (N_2677,In_3597,In_499);
or U2678 (N_2678,In_4121,In_2150);
xor U2679 (N_2679,In_1765,In_4197);
and U2680 (N_2680,In_3381,In_1113);
or U2681 (N_2681,In_1621,In_3205);
and U2682 (N_2682,In_458,In_2844);
or U2683 (N_2683,In_256,In_3002);
nand U2684 (N_2684,In_2769,In_2383);
or U2685 (N_2685,In_2966,In_4204);
nor U2686 (N_2686,In_4488,In_4173);
nand U2687 (N_2687,In_133,In_450);
nor U2688 (N_2688,In_220,In_3991);
or U2689 (N_2689,In_424,In_4865);
or U2690 (N_2690,In_2316,In_3996);
nand U2691 (N_2691,In_4572,In_646);
xor U2692 (N_2692,In_4711,In_1917);
nor U2693 (N_2693,In_3687,In_2331);
and U2694 (N_2694,In_3507,In_2333);
xnor U2695 (N_2695,In_4659,In_949);
nand U2696 (N_2696,In_4335,In_396);
nor U2697 (N_2697,In_3418,In_918);
or U2698 (N_2698,In_1166,In_2127);
xnor U2699 (N_2699,In_4581,In_1695);
and U2700 (N_2700,In_1486,In_2148);
nand U2701 (N_2701,In_476,In_2332);
and U2702 (N_2702,In_4792,In_4584);
nor U2703 (N_2703,In_4716,In_2498);
or U2704 (N_2704,In_4175,In_1516);
nand U2705 (N_2705,In_652,In_4137);
or U2706 (N_2706,In_897,In_4665);
xor U2707 (N_2707,In_3483,In_2201);
nor U2708 (N_2708,In_4940,In_1904);
nand U2709 (N_2709,In_702,In_184);
xnor U2710 (N_2710,In_2249,In_2988);
nor U2711 (N_2711,In_4893,In_654);
nor U2712 (N_2712,In_4467,In_599);
or U2713 (N_2713,In_1649,In_1363);
nand U2714 (N_2714,In_2220,In_1728);
xnor U2715 (N_2715,In_2543,In_2768);
nand U2716 (N_2716,In_4886,In_1865);
xnor U2717 (N_2717,In_1229,In_3762);
or U2718 (N_2718,In_4444,In_3661);
nand U2719 (N_2719,In_3123,In_4944);
nor U2720 (N_2720,In_4071,In_4061);
xor U2721 (N_2721,In_4147,In_2757);
or U2722 (N_2722,In_4731,In_696);
nor U2723 (N_2723,In_2425,In_4443);
and U2724 (N_2724,In_4391,In_1601);
and U2725 (N_2725,In_3355,In_466);
nor U2726 (N_2726,In_1346,In_185);
nand U2727 (N_2727,In_3390,In_65);
or U2728 (N_2728,In_1721,In_4648);
and U2729 (N_2729,In_4889,In_4407);
and U2730 (N_2730,In_4592,In_773);
nor U2731 (N_2731,In_325,In_4379);
nor U2732 (N_2732,In_960,In_3931);
and U2733 (N_2733,In_2677,In_4989);
and U2734 (N_2734,In_4411,In_1782);
nand U2735 (N_2735,In_2519,In_1837);
xor U2736 (N_2736,In_2547,In_1884);
xor U2737 (N_2737,In_4297,In_2976);
nor U2738 (N_2738,In_3479,In_2366);
xnor U2739 (N_2739,In_1327,In_4136);
and U2740 (N_2740,In_2931,In_2533);
or U2741 (N_2741,In_3216,In_2499);
xor U2742 (N_2742,In_3848,In_2734);
xnor U2743 (N_2743,In_2291,In_853);
or U2744 (N_2744,In_4783,In_836);
nand U2745 (N_2745,In_4169,In_4489);
nor U2746 (N_2746,In_3925,In_3906);
and U2747 (N_2747,In_2265,In_4212);
or U2748 (N_2748,In_2448,In_199);
and U2749 (N_2749,In_2709,In_2033);
nor U2750 (N_2750,In_2262,In_4945);
and U2751 (N_2751,In_1200,In_4209);
nand U2752 (N_2752,In_3861,In_3371);
and U2753 (N_2753,In_169,In_3822);
nor U2754 (N_2754,In_3724,In_2451);
or U2755 (N_2755,In_3052,In_2182);
and U2756 (N_2756,In_2270,In_295);
nor U2757 (N_2757,In_2918,In_1612);
xor U2758 (N_2758,In_3786,In_4570);
and U2759 (N_2759,In_4526,In_295);
xnor U2760 (N_2760,In_4529,In_100);
xor U2761 (N_2761,In_2946,In_2939);
xnor U2762 (N_2762,In_4003,In_2707);
or U2763 (N_2763,In_4156,In_3085);
nand U2764 (N_2764,In_1013,In_2943);
nand U2765 (N_2765,In_3960,In_3384);
or U2766 (N_2766,In_51,In_183);
xnor U2767 (N_2767,In_2793,In_4244);
nor U2768 (N_2768,In_4635,In_76);
or U2769 (N_2769,In_1387,In_1268);
or U2770 (N_2770,In_3942,In_563);
nor U2771 (N_2771,In_4657,In_4967);
nor U2772 (N_2772,In_2913,In_418);
nand U2773 (N_2773,In_397,In_3573);
nand U2774 (N_2774,In_714,In_3072);
nor U2775 (N_2775,In_2531,In_2625);
and U2776 (N_2776,In_1434,In_3753);
or U2777 (N_2777,In_2443,In_1903);
or U2778 (N_2778,In_2118,In_301);
nand U2779 (N_2779,In_355,In_3841);
or U2780 (N_2780,In_4712,In_1307);
nor U2781 (N_2781,In_115,In_1217);
xor U2782 (N_2782,In_2160,In_2888);
nor U2783 (N_2783,In_3380,In_4338);
or U2784 (N_2784,In_2135,In_964);
and U2785 (N_2785,In_4291,In_1088);
nand U2786 (N_2786,In_2105,In_3727);
nor U2787 (N_2787,In_3899,In_1352);
or U2788 (N_2788,In_947,In_3911);
nor U2789 (N_2789,In_4753,In_3901);
nor U2790 (N_2790,In_4154,In_4500);
or U2791 (N_2791,In_4350,In_2282);
nor U2792 (N_2792,In_456,In_4935);
or U2793 (N_2793,In_545,In_920);
and U2794 (N_2794,In_3209,In_1601);
and U2795 (N_2795,In_1531,In_1942);
xnor U2796 (N_2796,In_1054,In_1111);
nand U2797 (N_2797,In_3790,In_419);
or U2798 (N_2798,In_4500,In_2349);
nor U2799 (N_2799,In_2956,In_11);
nand U2800 (N_2800,In_3020,In_4593);
nand U2801 (N_2801,In_2853,In_779);
or U2802 (N_2802,In_12,In_1424);
and U2803 (N_2803,In_1920,In_4180);
xnor U2804 (N_2804,In_705,In_2322);
or U2805 (N_2805,In_2140,In_2752);
and U2806 (N_2806,In_2265,In_4159);
xor U2807 (N_2807,In_3465,In_4597);
xnor U2808 (N_2808,In_4306,In_4296);
nand U2809 (N_2809,In_2594,In_2850);
nand U2810 (N_2810,In_2175,In_1068);
xor U2811 (N_2811,In_4241,In_2524);
nor U2812 (N_2812,In_3750,In_4435);
xor U2813 (N_2813,In_4603,In_2728);
and U2814 (N_2814,In_3789,In_4426);
nor U2815 (N_2815,In_2441,In_2587);
nand U2816 (N_2816,In_2323,In_4055);
nor U2817 (N_2817,In_3936,In_3802);
and U2818 (N_2818,In_4317,In_236);
or U2819 (N_2819,In_99,In_3321);
and U2820 (N_2820,In_303,In_2533);
nor U2821 (N_2821,In_1495,In_455);
nand U2822 (N_2822,In_3932,In_499);
xor U2823 (N_2823,In_4894,In_2947);
and U2824 (N_2824,In_1201,In_2858);
xnor U2825 (N_2825,In_2162,In_160);
nor U2826 (N_2826,In_970,In_2990);
or U2827 (N_2827,In_1251,In_2482);
and U2828 (N_2828,In_1449,In_4947);
xor U2829 (N_2829,In_4224,In_1953);
or U2830 (N_2830,In_4704,In_2626);
or U2831 (N_2831,In_2217,In_4678);
or U2832 (N_2832,In_2654,In_4147);
nand U2833 (N_2833,In_3916,In_1560);
and U2834 (N_2834,In_123,In_3854);
nor U2835 (N_2835,In_1963,In_638);
nor U2836 (N_2836,In_2682,In_1411);
xor U2837 (N_2837,In_3121,In_3970);
nand U2838 (N_2838,In_2880,In_3744);
and U2839 (N_2839,In_4032,In_1243);
and U2840 (N_2840,In_1134,In_4380);
nand U2841 (N_2841,In_3844,In_2979);
nor U2842 (N_2842,In_3334,In_1085);
xor U2843 (N_2843,In_4099,In_3930);
xor U2844 (N_2844,In_3966,In_4816);
nand U2845 (N_2845,In_3730,In_1686);
and U2846 (N_2846,In_1178,In_130);
and U2847 (N_2847,In_431,In_3685);
or U2848 (N_2848,In_1264,In_1621);
xnor U2849 (N_2849,In_3661,In_965);
nor U2850 (N_2850,In_3015,In_2570);
nand U2851 (N_2851,In_3462,In_3809);
xor U2852 (N_2852,In_1987,In_1060);
nand U2853 (N_2853,In_4307,In_2604);
nand U2854 (N_2854,In_375,In_1018);
nor U2855 (N_2855,In_482,In_2190);
or U2856 (N_2856,In_2175,In_4422);
or U2857 (N_2857,In_267,In_2269);
xor U2858 (N_2858,In_281,In_209);
nor U2859 (N_2859,In_1622,In_3322);
nand U2860 (N_2860,In_1674,In_1284);
nand U2861 (N_2861,In_3269,In_3206);
xor U2862 (N_2862,In_394,In_321);
nor U2863 (N_2863,In_4555,In_1812);
nor U2864 (N_2864,In_4461,In_1548);
and U2865 (N_2865,In_2045,In_1358);
and U2866 (N_2866,In_4770,In_3712);
nor U2867 (N_2867,In_3629,In_3635);
or U2868 (N_2868,In_278,In_4260);
or U2869 (N_2869,In_3906,In_3998);
and U2870 (N_2870,In_1534,In_1126);
nand U2871 (N_2871,In_3004,In_4619);
nand U2872 (N_2872,In_3099,In_2215);
nor U2873 (N_2873,In_1109,In_3091);
nor U2874 (N_2874,In_65,In_2469);
or U2875 (N_2875,In_2054,In_697);
xnor U2876 (N_2876,In_4608,In_3259);
nand U2877 (N_2877,In_297,In_1816);
or U2878 (N_2878,In_257,In_1589);
xnor U2879 (N_2879,In_4067,In_1582);
nor U2880 (N_2880,In_2010,In_1574);
and U2881 (N_2881,In_3284,In_4976);
xor U2882 (N_2882,In_1037,In_2425);
nand U2883 (N_2883,In_3363,In_806);
nand U2884 (N_2884,In_521,In_4800);
nor U2885 (N_2885,In_1704,In_3755);
xor U2886 (N_2886,In_362,In_3180);
nor U2887 (N_2887,In_2116,In_1602);
and U2888 (N_2888,In_4078,In_3029);
nand U2889 (N_2889,In_2420,In_3939);
xnor U2890 (N_2890,In_4971,In_2734);
xnor U2891 (N_2891,In_4269,In_1920);
nand U2892 (N_2892,In_306,In_737);
nor U2893 (N_2893,In_1398,In_1421);
or U2894 (N_2894,In_3970,In_2605);
nor U2895 (N_2895,In_2786,In_1470);
or U2896 (N_2896,In_1785,In_2334);
xor U2897 (N_2897,In_3105,In_2459);
nor U2898 (N_2898,In_1581,In_3114);
nor U2899 (N_2899,In_2077,In_3793);
nor U2900 (N_2900,In_817,In_1956);
nand U2901 (N_2901,In_689,In_1834);
xnor U2902 (N_2902,In_303,In_2341);
and U2903 (N_2903,In_4989,In_3569);
and U2904 (N_2904,In_2518,In_3477);
xnor U2905 (N_2905,In_3498,In_1927);
nor U2906 (N_2906,In_4967,In_2332);
or U2907 (N_2907,In_4775,In_2329);
xnor U2908 (N_2908,In_1214,In_4118);
xor U2909 (N_2909,In_3688,In_1231);
and U2910 (N_2910,In_1526,In_513);
xor U2911 (N_2911,In_2140,In_489);
xnor U2912 (N_2912,In_706,In_1149);
nand U2913 (N_2913,In_4873,In_4299);
nor U2914 (N_2914,In_1351,In_3273);
xor U2915 (N_2915,In_3290,In_3297);
and U2916 (N_2916,In_4831,In_1625);
and U2917 (N_2917,In_2482,In_4520);
or U2918 (N_2918,In_1970,In_3770);
or U2919 (N_2919,In_4106,In_4516);
nand U2920 (N_2920,In_3335,In_1446);
nand U2921 (N_2921,In_4842,In_3080);
or U2922 (N_2922,In_4627,In_3393);
nand U2923 (N_2923,In_1312,In_4049);
xor U2924 (N_2924,In_566,In_322);
and U2925 (N_2925,In_4011,In_350);
nand U2926 (N_2926,In_2874,In_587);
xnor U2927 (N_2927,In_3548,In_1862);
nor U2928 (N_2928,In_4567,In_1228);
nor U2929 (N_2929,In_2107,In_4262);
and U2930 (N_2930,In_999,In_1504);
nand U2931 (N_2931,In_3254,In_4462);
xnor U2932 (N_2932,In_3433,In_44);
xnor U2933 (N_2933,In_3287,In_1895);
xor U2934 (N_2934,In_1219,In_235);
xnor U2935 (N_2935,In_4233,In_2998);
and U2936 (N_2936,In_1379,In_3348);
or U2937 (N_2937,In_3529,In_436);
nor U2938 (N_2938,In_718,In_1994);
or U2939 (N_2939,In_4034,In_791);
xor U2940 (N_2940,In_1766,In_1761);
nand U2941 (N_2941,In_3458,In_1950);
or U2942 (N_2942,In_816,In_2296);
or U2943 (N_2943,In_1423,In_3822);
nor U2944 (N_2944,In_1520,In_1303);
or U2945 (N_2945,In_4855,In_3479);
or U2946 (N_2946,In_2348,In_2687);
xor U2947 (N_2947,In_2239,In_4892);
nand U2948 (N_2948,In_1990,In_2477);
and U2949 (N_2949,In_4352,In_4134);
or U2950 (N_2950,In_2081,In_4086);
nand U2951 (N_2951,In_4294,In_3518);
or U2952 (N_2952,In_2263,In_3781);
xnor U2953 (N_2953,In_1302,In_3448);
or U2954 (N_2954,In_3592,In_65);
and U2955 (N_2955,In_2986,In_1367);
nand U2956 (N_2956,In_226,In_4044);
nor U2957 (N_2957,In_1134,In_1728);
nand U2958 (N_2958,In_1692,In_4132);
xor U2959 (N_2959,In_1489,In_2696);
nor U2960 (N_2960,In_2478,In_24);
and U2961 (N_2961,In_2242,In_1008);
or U2962 (N_2962,In_3507,In_275);
nand U2963 (N_2963,In_1877,In_3453);
or U2964 (N_2964,In_413,In_1148);
nor U2965 (N_2965,In_2599,In_1790);
nor U2966 (N_2966,In_1239,In_3814);
xnor U2967 (N_2967,In_4567,In_2903);
xor U2968 (N_2968,In_3122,In_1080);
and U2969 (N_2969,In_825,In_1176);
and U2970 (N_2970,In_3469,In_3233);
and U2971 (N_2971,In_1257,In_3317);
nand U2972 (N_2972,In_1365,In_2119);
nor U2973 (N_2973,In_460,In_1492);
nor U2974 (N_2974,In_1126,In_1332);
xor U2975 (N_2975,In_3853,In_62);
or U2976 (N_2976,In_3447,In_1021);
nand U2977 (N_2977,In_919,In_438);
or U2978 (N_2978,In_1554,In_1781);
or U2979 (N_2979,In_4519,In_3037);
or U2980 (N_2980,In_1097,In_833);
nand U2981 (N_2981,In_3561,In_3011);
and U2982 (N_2982,In_3082,In_3403);
nand U2983 (N_2983,In_2609,In_3801);
nor U2984 (N_2984,In_702,In_2338);
xnor U2985 (N_2985,In_324,In_3141);
nand U2986 (N_2986,In_849,In_1011);
nor U2987 (N_2987,In_4703,In_51);
or U2988 (N_2988,In_1669,In_3464);
or U2989 (N_2989,In_634,In_4933);
nor U2990 (N_2990,In_1157,In_418);
and U2991 (N_2991,In_4154,In_4513);
xnor U2992 (N_2992,In_2002,In_2917);
and U2993 (N_2993,In_3161,In_834);
and U2994 (N_2994,In_1608,In_869);
nor U2995 (N_2995,In_4276,In_1508);
nor U2996 (N_2996,In_856,In_674);
xnor U2997 (N_2997,In_2512,In_3729);
nand U2998 (N_2998,In_115,In_1720);
or U2999 (N_2999,In_4446,In_4205);
and U3000 (N_3000,In_1741,In_3760);
or U3001 (N_3001,In_3204,In_2479);
nand U3002 (N_3002,In_2600,In_1582);
xor U3003 (N_3003,In_3817,In_1638);
nand U3004 (N_3004,In_1789,In_2698);
xnor U3005 (N_3005,In_2014,In_2160);
nand U3006 (N_3006,In_4169,In_4249);
and U3007 (N_3007,In_4910,In_377);
and U3008 (N_3008,In_334,In_1933);
nor U3009 (N_3009,In_3540,In_3454);
xor U3010 (N_3010,In_1761,In_1042);
or U3011 (N_3011,In_3931,In_4275);
nor U3012 (N_3012,In_1984,In_2365);
nand U3013 (N_3013,In_280,In_3343);
and U3014 (N_3014,In_765,In_1266);
or U3015 (N_3015,In_1691,In_503);
xnor U3016 (N_3016,In_1885,In_31);
xor U3017 (N_3017,In_2371,In_2783);
or U3018 (N_3018,In_3837,In_2724);
nand U3019 (N_3019,In_3073,In_4445);
nor U3020 (N_3020,In_1075,In_1218);
nor U3021 (N_3021,In_2717,In_1651);
nor U3022 (N_3022,In_582,In_3449);
and U3023 (N_3023,In_888,In_3813);
nor U3024 (N_3024,In_57,In_2118);
or U3025 (N_3025,In_1962,In_2626);
and U3026 (N_3026,In_4012,In_3367);
xnor U3027 (N_3027,In_4878,In_2008);
xnor U3028 (N_3028,In_1841,In_2020);
or U3029 (N_3029,In_2957,In_1465);
xnor U3030 (N_3030,In_704,In_4970);
and U3031 (N_3031,In_2864,In_1277);
and U3032 (N_3032,In_2007,In_341);
and U3033 (N_3033,In_968,In_268);
and U3034 (N_3034,In_2038,In_4328);
nor U3035 (N_3035,In_1036,In_2940);
nand U3036 (N_3036,In_2641,In_4986);
xor U3037 (N_3037,In_2913,In_3327);
nor U3038 (N_3038,In_2980,In_3028);
nor U3039 (N_3039,In_2485,In_1389);
xor U3040 (N_3040,In_683,In_382);
xnor U3041 (N_3041,In_4152,In_1499);
nand U3042 (N_3042,In_1616,In_3735);
xnor U3043 (N_3043,In_1031,In_3423);
and U3044 (N_3044,In_2803,In_2568);
nor U3045 (N_3045,In_715,In_3306);
and U3046 (N_3046,In_2660,In_4080);
nor U3047 (N_3047,In_1510,In_3676);
and U3048 (N_3048,In_1036,In_4525);
and U3049 (N_3049,In_2039,In_4929);
nor U3050 (N_3050,In_4356,In_3369);
nor U3051 (N_3051,In_645,In_4605);
or U3052 (N_3052,In_520,In_775);
and U3053 (N_3053,In_432,In_4714);
xor U3054 (N_3054,In_4848,In_1386);
or U3055 (N_3055,In_4921,In_3164);
xnor U3056 (N_3056,In_2812,In_1024);
nor U3057 (N_3057,In_1156,In_4692);
and U3058 (N_3058,In_4282,In_4028);
nor U3059 (N_3059,In_1260,In_2850);
nand U3060 (N_3060,In_309,In_381);
and U3061 (N_3061,In_4202,In_3743);
and U3062 (N_3062,In_4319,In_629);
nor U3063 (N_3063,In_4522,In_776);
or U3064 (N_3064,In_4814,In_4705);
xor U3065 (N_3065,In_1065,In_1255);
and U3066 (N_3066,In_3791,In_4211);
nor U3067 (N_3067,In_4704,In_327);
nand U3068 (N_3068,In_2917,In_52);
or U3069 (N_3069,In_4485,In_815);
and U3070 (N_3070,In_3318,In_3144);
nor U3071 (N_3071,In_4185,In_4656);
or U3072 (N_3072,In_3325,In_2016);
or U3073 (N_3073,In_1788,In_147);
nand U3074 (N_3074,In_965,In_4439);
xnor U3075 (N_3075,In_140,In_1064);
or U3076 (N_3076,In_3127,In_4346);
xor U3077 (N_3077,In_793,In_2622);
xnor U3078 (N_3078,In_2478,In_269);
nor U3079 (N_3079,In_3229,In_1185);
and U3080 (N_3080,In_2519,In_46);
xnor U3081 (N_3081,In_1937,In_908);
or U3082 (N_3082,In_298,In_3872);
nor U3083 (N_3083,In_184,In_3290);
or U3084 (N_3084,In_1714,In_582);
and U3085 (N_3085,In_1458,In_3096);
nor U3086 (N_3086,In_293,In_4617);
xor U3087 (N_3087,In_3298,In_1424);
nor U3088 (N_3088,In_988,In_1848);
or U3089 (N_3089,In_1593,In_270);
and U3090 (N_3090,In_353,In_478);
nor U3091 (N_3091,In_4506,In_3448);
and U3092 (N_3092,In_2805,In_573);
or U3093 (N_3093,In_80,In_3498);
nand U3094 (N_3094,In_3777,In_3087);
and U3095 (N_3095,In_2520,In_946);
or U3096 (N_3096,In_3444,In_4619);
nand U3097 (N_3097,In_1860,In_4340);
and U3098 (N_3098,In_4495,In_2097);
xor U3099 (N_3099,In_3249,In_4343);
xnor U3100 (N_3100,In_265,In_1385);
xnor U3101 (N_3101,In_4426,In_2777);
and U3102 (N_3102,In_2351,In_4799);
and U3103 (N_3103,In_406,In_909);
nand U3104 (N_3104,In_559,In_4461);
and U3105 (N_3105,In_1257,In_4821);
xor U3106 (N_3106,In_32,In_3439);
and U3107 (N_3107,In_1461,In_815);
nor U3108 (N_3108,In_2069,In_3728);
or U3109 (N_3109,In_2375,In_2000);
or U3110 (N_3110,In_3027,In_2739);
nand U3111 (N_3111,In_3402,In_4240);
xor U3112 (N_3112,In_2215,In_2075);
xnor U3113 (N_3113,In_1423,In_4149);
and U3114 (N_3114,In_4325,In_2752);
nand U3115 (N_3115,In_47,In_1786);
nor U3116 (N_3116,In_365,In_159);
or U3117 (N_3117,In_4763,In_3119);
nand U3118 (N_3118,In_1822,In_3371);
nand U3119 (N_3119,In_3957,In_4503);
nor U3120 (N_3120,In_2829,In_647);
and U3121 (N_3121,In_2788,In_163);
or U3122 (N_3122,In_648,In_330);
or U3123 (N_3123,In_4195,In_2220);
nor U3124 (N_3124,In_1297,In_826);
nand U3125 (N_3125,In_800,In_4216);
nand U3126 (N_3126,In_1673,In_1073);
and U3127 (N_3127,In_4873,In_1080);
nor U3128 (N_3128,In_2899,In_3534);
nor U3129 (N_3129,In_3614,In_2137);
and U3130 (N_3130,In_4520,In_2337);
nand U3131 (N_3131,In_3315,In_3964);
or U3132 (N_3132,In_1613,In_1599);
nor U3133 (N_3133,In_3224,In_3000);
xor U3134 (N_3134,In_840,In_491);
nand U3135 (N_3135,In_2469,In_2717);
or U3136 (N_3136,In_1066,In_1011);
nor U3137 (N_3137,In_1043,In_2507);
and U3138 (N_3138,In_2517,In_3465);
xnor U3139 (N_3139,In_2787,In_1941);
or U3140 (N_3140,In_4409,In_43);
xor U3141 (N_3141,In_3070,In_2836);
xor U3142 (N_3142,In_4924,In_2034);
and U3143 (N_3143,In_3536,In_3132);
nor U3144 (N_3144,In_915,In_403);
nand U3145 (N_3145,In_2971,In_4876);
and U3146 (N_3146,In_4945,In_3073);
or U3147 (N_3147,In_46,In_4157);
nand U3148 (N_3148,In_4344,In_1433);
nand U3149 (N_3149,In_2672,In_284);
nand U3150 (N_3150,In_430,In_2525);
nand U3151 (N_3151,In_1467,In_2085);
xnor U3152 (N_3152,In_482,In_2408);
or U3153 (N_3153,In_4771,In_2874);
nand U3154 (N_3154,In_2878,In_3697);
nand U3155 (N_3155,In_781,In_177);
nor U3156 (N_3156,In_2138,In_1433);
or U3157 (N_3157,In_670,In_2932);
nor U3158 (N_3158,In_1083,In_3560);
xnor U3159 (N_3159,In_1316,In_2684);
and U3160 (N_3160,In_3223,In_1022);
or U3161 (N_3161,In_4816,In_191);
and U3162 (N_3162,In_3501,In_115);
or U3163 (N_3163,In_2910,In_1655);
or U3164 (N_3164,In_1137,In_1976);
or U3165 (N_3165,In_2339,In_4663);
xnor U3166 (N_3166,In_1672,In_1604);
nand U3167 (N_3167,In_2093,In_130);
xor U3168 (N_3168,In_1416,In_1820);
or U3169 (N_3169,In_170,In_110);
nand U3170 (N_3170,In_4218,In_2159);
nand U3171 (N_3171,In_1133,In_218);
and U3172 (N_3172,In_2415,In_167);
or U3173 (N_3173,In_1028,In_3796);
and U3174 (N_3174,In_466,In_4233);
nor U3175 (N_3175,In_4405,In_2042);
and U3176 (N_3176,In_4341,In_4682);
and U3177 (N_3177,In_506,In_1838);
xor U3178 (N_3178,In_1984,In_2232);
nor U3179 (N_3179,In_3953,In_1267);
nand U3180 (N_3180,In_2903,In_1409);
and U3181 (N_3181,In_1675,In_2385);
or U3182 (N_3182,In_2930,In_3608);
xor U3183 (N_3183,In_1817,In_397);
and U3184 (N_3184,In_4277,In_310);
or U3185 (N_3185,In_4777,In_2633);
nand U3186 (N_3186,In_4680,In_121);
nand U3187 (N_3187,In_2165,In_2329);
nand U3188 (N_3188,In_3011,In_1198);
xor U3189 (N_3189,In_1394,In_35);
nor U3190 (N_3190,In_24,In_1250);
nor U3191 (N_3191,In_3666,In_4328);
nand U3192 (N_3192,In_1986,In_903);
or U3193 (N_3193,In_4422,In_3776);
nand U3194 (N_3194,In_3202,In_23);
and U3195 (N_3195,In_4245,In_3596);
xor U3196 (N_3196,In_3691,In_3753);
xnor U3197 (N_3197,In_2716,In_1415);
and U3198 (N_3198,In_1440,In_233);
and U3199 (N_3199,In_2301,In_4954);
xnor U3200 (N_3200,In_345,In_2232);
nor U3201 (N_3201,In_4441,In_2393);
nor U3202 (N_3202,In_2759,In_2953);
or U3203 (N_3203,In_4828,In_4368);
nor U3204 (N_3204,In_129,In_1409);
xnor U3205 (N_3205,In_2453,In_3902);
and U3206 (N_3206,In_2443,In_1496);
or U3207 (N_3207,In_3214,In_1021);
nor U3208 (N_3208,In_3689,In_2550);
xnor U3209 (N_3209,In_4192,In_4215);
or U3210 (N_3210,In_3136,In_779);
nor U3211 (N_3211,In_4524,In_1560);
xnor U3212 (N_3212,In_4131,In_4679);
xnor U3213 (N_3213,In_2713,In_2818);
and U3214 (N_3214,In_3874,In_2547);
nand U3215 (N_3215,In_1794,In_1163);
nand U3216 (N_3216,In_2435,In_1513);
nand U3217 (N_3217,In_4364,In_2723);
nand U3218 (N_3218,In_4998,In_3113);
xnor U3219 (N_3219,In_2195,In_4835);
or U3220 (N_3220,In_1305,In_2533);
nor U3221 (N_3221,In_259,In_1506);
nor U3222 (N_3222,In_313,In_1182);
nor U3223 (N_3223,In_2267,In_158);
and U3224 (N_3224,In_4492,In_276);
nand U3225 (N_3225,In_2773,In_951);
or U3226 (N_3226,In_1248,In_3655);
nor U3227 (N_3227,In_4997,In_3396);
nor U3228 (N_3228,In_3661,In_2148);
or U3229 (N_3229,In_3571,In_150);
nand U3230 (N_3230,In_2475,In_931);
and U3231 (N_3231,In_2119,In_1389);
nor U3232 (N_3232,In_4403,In_3460);
nand U3233 (N_3233,In_4055,In_1713);
nor U3234 (N_3234,In_3185,In_1620);
or U3235 (N_3235,In_1083,In_3361);
nand U3236 (N_3236,In_1430,In_3625);
or U3237 (N_3237,In_3188,In_1065);
and U3238 (N_3238,In_1164,In_8);
nand U3239 (N_3239,In_90,In_2862);
nor U3240 (N_3240,In_3975,In_1323);
or U3241 (N_3241,In_4575,In_3734);
xnor U3242 (N_3242,In_1499,In_4046);
and U3243 (N_3243,In_181,In_2150);
nand U3244 (N_3244,In_834,In_1180);
or U3245 (N_3245,In_1628,In_532);
nand U3246 (N_3246,In_2883,In_2850);
or U3247 (N_3247,In_3062,In_4713);
or U3248 (N_3248,In_1724,In_4271);
or U3249 (N_3249,In_3657,In_3705);
or U3250 (N_3250,In_540,In_4625);
or U3251 (N_3251,In_3074,In_2789);
xnor U3252 (N_3252,In_690,In_678);
xnor U3253 (N_3253,In_2083,In_1036);
or U3254 (N_3254,In_4232,In_592);
and U3255 (N_3255,In_1508,In_4515);
or U3256 (N_3256,In_185,In_721);
or U3257 (N_3257,In_421,In_3049);
and U3258 (N_3258,In_1257,In_4324);
nand U3259 (N_3259,In_500,In_711);
nand U3260 (N_3260,In_2267,In_680);
nor U3261 (N_3261,In_3217,In_704);
or U3262 (N_3262,In_4188,In_4901);
or U3263 (N_3263,In_4186,In_2114);
and U3264 (N_3264,In_669,In_189);
and U3265 (N_3265,In_4589,In_665);
and U3266 (N_3266,In_3931,In_4987);
or U3267 (N_3267,In_883,In_4374);
or U3268 (N_3268,In_591,In_2743);
xor U3269 (N_3269,In_1754,In_1253);
or U3270 (N_3270,In_2380,In_443);
nand U3271 (N_3271,In_2086,In_27);
and U3272 (N_3272,In_153,In_458);
nor U3273 (N_3273,In_1538,In_3163);
and U3274 (N_3274,In_4942,In_2881);
nor U3275 (N_3275,In_3321,In_4338);
or U3276 (N_3276,In_780,In_219);
nor U3277 (N_3277,In_4695,In_4646);
nor U3278 (N_3278,In_3604,In_2398);
and U3279 (N_3279,In_1915,In_3580);
nand U3280 (N_3280,In_4995,In_3899);
and U3281 (N_3281,In_952,In_1729);
nand U3282 (N_3282,In_2395,In_2666);
nor U3283 (N_3283,In_4703,In_77);
and U3284 (N_3284,In_346,In_2124);
nor U3285 (N_3285,In_1851,In_3068);
nor U3286 (N_3286,In_3675,In_1833);
nor U3287 (N_3287,In_4829,In_1390);
and U3288 (N_3288,In_3737,In_1692);
or U3289 (N_3289,In_4729,In_2727);
or U3290 (N_3290,In_2761,In_4569);
or U3291 (N_3291,In_1460,In_3150);
xnor U3292 (N_3292,In_890,In_139);
and U3293 (N_3293,In_1505,In_3244);
and U3294 (N_3294,In_302,In_3295);
xnor U3295 (N_3295,In_3575,In_4026);
and U3296 (N_3296,In_3943,In_3332);
or U3297 (N_3297,In_320,In_2974);
nor U3298 (N_3298,In_1285,In_3467);
nand U3299 (N_3299,In_924,In_3588);
and U3300 (N_3300,In_1200,In_1099);
nor U3301 (N_3301,In_264,In_619);
nor U3302 (N_3302,In_2187,In_3732);
and U3303 (N_3303,In_1571,In_924);
and U3304 (N_3304,In_1230,In_4248);
or U3305 (N_3305,In_468,In_797);
xor U3306 (N_3306,In_4095,In_1575);
nor U3307 (N_3307,In_1757,In_4106);
or U3308 (N_3308,In_2221,In_947);
nor U3309 (N_3309,In_2237,In_596);
nand U3310 (N_3310,In_1522,In_3864);
nand U3311 (N_3311,In_3205,In_3945);
nand U3312 (N_3312,In_886,In_3688);
nor U3313 (N_3313,In_2325,In_1359);
or U3314 (N_3314,In_544,In_415);
or U3315 (N_3315,In_932,In_3972);
xor U3316 (N_3316,In_985,In_177);
nor U3317 (N_3317,In_2932,In_4657);
nor U3318 (N_3318,In_4876,In_929);
nor U3319 (N_3319,In_3080,In_4862);
or U3320 (N_3320,In_3193,In_1028);
nand U3321 (N_3321,In_1870,In_2863);
or U3322 (N_3322,In_2167,In_1434);
xnor U3323 (N_3323,In_4437,In_3271);
nor U3324 (N_3324,In_2422,In_1287);
xnor U3325 (N_3325,In_2712,In_3275);
nor U3326 (N_3326,In_897,In_3216);
nor U3327 (N_3327,In_1933,In_3992);
nand U3328 (N_3328,In_3087,In_2653);
or U3329 (N_3329,In_2169,In_2460);
or U3330 (N_3330,In_2636,In_3071);
xnor U3331 (N_3331,In_3340,In_3097);
nor U3332 (N_3332,In_563,In_2709);
nand U3333 (N_3333,In_911,In_1345);
nor U3334 (N_3334,In_2137,In_366);
nand U3335 (N_3335,In_3363,In_2373);
nand U3336 (N_3336,In_2865,In_2052);
nand U3337 (N_3337,In_428,In_3002);
xnor U3338 (N_3338,In_2895,In_4837);
and U3339 (N_3339,In_2601,In_537);
xnor U3340 (N_3340,In_2429,In_2194);
nand U3341 (N_3341,In_1152,In_4578);
and U3342 (N_3342,In_3993,In_2299);
nor U3343 (N_3343,In_735,In_1608);
xnor U3344 (N_3344,In_4230,In_2069);
nor U3345 (N_3345,In_3215,In_238);
or U3346 (N_3346,In_3016,In_2935);
xor U3347 (N_3347,In_1949,In_60);
and U3348 (N_3348,In_4679,In_1999);
or U3349 (N_3349,In_2305,In_2234);
and U3350 (N_3350,In_1587,In_2950);
or U3351 (N_3351,In_1317,In_3362);
nand U3352 (N_3352,In_3198,In_4892);
xor U3353 (N_3353,In_123,In_163);
xnor U3354 (N_3354,In_3832,In_2869);
nand U3355 (N_3355,In_2117,In_2535);
nor U3356 (N_3356,In_1463,In_1166);
nand U3357 (N_3357,In_1059,In_3311);
nand U3358 (N_3358,In_1774,In_4764);
nor U3359 (N_3359,In_3605,In_864);
nor U3360 (N_3360,In_1057,In_2195);
or U3361 (N_3361,In_4126,In_1343);
nor U3362 (N_3362,In_1298,In_647);
and U3363 (N_3363,In_997,In_4694);
nand U3364 (N_3364,In_4405,In_972);
xor U3365 (N_3365,In_2385,In_3644);
xnor U3366 (N_3366,In_1794,In_2704);
nor U3367 (N_3367,In_4109,In_4720);
or U3368 (N_3368,In_1407,In_3800);
or U3369 (N_3369,In_4695,In_87);
xnor U3370 (N_3370,In_2436,In_1344);
and U3371 (N_3371,In_2316,In_4070);
or U3372 (N_3372,In_778,In_2393);
nand U3373 (N_3373,In_4600,In_1194);
nand U3374 (N_3374,In_1906,In_4519);
and U3375 (N_3375,In_3442,In_2758);
xnor U3376 (N_3376,In_760,In_3615);
or U3377 (N_3377,In_4747,In_4047);
nor U3378 (N_3378,In_994,In_227);
nand U3379 (N_3379,In_4903,In_264);
xor U3380 (N_3380,In_1459,In_4111);
nand U3381 (N_3381,In_2077,In_1744);
and U3382 (N_3382,In_3783,In_3304);
nor U3383 (N_3383,In_1729,In_3583);
or U3384 (N_3384,In_2130,In_4623);
and U3385 (N_3385,In_1067,In_4260);
nand U3386 (N_3386,In_3109,In_4254);
nand U3387 (N_3387,In_4182,In_2627);
xnor U3388 (N_3388,In_3411,In_4256);
xnor U3389 (N_3389,In_4104,In_4975);
nor U3390 (N_3390,In_4465,In_2757);
nor U3391 (N_3391,In_2019,In_3205);
or U3392 (N_3392,In_4533,In_3472);
nor U3393 (N_3393,In_2432,In_571);
nand U3394 (N_3394,In_1201,In_4497);
xnor U3395 (N_3395,In_1564,In_1179);
nor U3396 (N_3396,In_581,In_1102);
xnor U3397 (N_3397,In_3473,In_727);
xor U3398 (N_3398,In_3634,In_4382);
xnor U3399 (N_3399,In_1363,In_3186);
and U3400 (N_3400,In_996,In_1704);
nand U3401 (N_3401,In_3664,In_2758);
nand U3402 (N_3402,In_573,In_4066);
and U3403 (N_3403,In_397,In_3866);
xor U3404 (N_3404,In_3579,In_4396);
or U3405 (N_3405,In_1586,In_2630);
and U3406 (N_3406,In_4996,In_357);
and U3407 (N_3407,In_3008,In_2633);
and U3408 (N_3408,In_3951,In_161);
and U3409 (N_3409,In_2875,In_3135);
nor U3410 (N_3410,In_2765,In_471);
nor U3411 (N_3411,In_4253,In_890);
nand U3412 (N_3412,In_983,In_1018);
xor U3413 (N_3413,In_4322,In_4469);
or U3414 (N_3414,In_2016,In_4981);
or U3415 (N_3415,In_3594,In_2133);
nand U3416 (N_3416,In_3645,In_3837);
or U3417 (N_3417,In_286,In_1127);
nor U3418 (N_3418,In_3181,In_1512);
nand U3419 (N_3419,In_35,In_868);
and U3420 (N_3420,In_2907,In_365);
nand U3421 (N_3421,In_4506,In_3035);
and U3422 (N_3422,In_912,In_2691);
nand U3423 (N_3423,In_2240,In_3224);
or U3424 (N_3424,In_1629,In_1095);
nor U3425 (N_3425,In_2144,In_183);
nor U3426 (N_3426,In_4517,In_3658);
or U3427 (N_3427,In_4094,In_3538);
xor U3428 (N_3428,In_4688,In_3000);
and U3429 (N_3429,In_3822,In_1727);
nand U3430 (N_3430,In_4576,In_3036);
nand U3431 (N_3431,In_4959,In_232);
xor U3432 (N_3432,In_3217,In_657);
xnor U3433 (N_3433,In_4321,In_838);
nand U3434 (N_3434,In_4549,In_973);
nor U3435 (N_3435,In_4485,In_17);
xor U3436 (N_3436,In_889,In_3887);
or U3437 (N_3437,In_2186,In_4934);
xor U3438 (N_3438,In_2663,In_217);
and U3439 (N_3439,In_3250,In_2845);
nand U3440 (N_3440,In_1317,In_2429);
xnor U3441 (N_3441,In_4156,In_313);
and U3442 (N_3442,In_4953,In_1195);
xnor U3443 (N_3443,In_4744,In_3753);
nand U3444 (N_3444,In_4515,In_1326);
or U3445 (N_3445,In_405,In_3834);
xnor U3446 (N_3446,In_4106,In_2209);
nor U3447 (N_3447,In_3504,In_2146);
nand U3448 (N_3448,In_244,In_106);
nor U3449 (N_3449,In_2956,In_2439);
and U3450 (N_3450,In_3318,In_284);
and U3451 (N_3451,In_58,In_2383);
or U3452 (N_3452,In_2567,In_83);
xnor U3453 (N_3453,In_1669,In_3706);
and U3454 (N_3454,In_1533,In_3181);
or U3455 (N_3455,In_1313,In_4890);
or U3456 (N_3456,In_4897,In_1663);
nand U3457 (N_3457,In_4674,In_2119);
xnor U3458 (N_3458,In_3354,In_3329);
and U3459 (N_3459,In_1244,In_3);
xnor U3460 (N_3460,In_4955,In_4681);
or U3461 (N_3461,In_4091,In_3654);
xor U3462 (N_3462,In_2328,In_4468);
and U3463 (N_3463,In_675,In_3171);
nand U3464 (N_3464,In_2180,In_593);
or U3465 (N_3465,In_4666,In_4662);
and U3466 (N_3466,In_1222,In_4676);
nand U3467 (N_3467,In_1180,In_3712);
and U3468 (N_3468,In_3450,In_4250);
and U3469 (N_3469,In_4787,In_3214);
nor U3470 (N_3470,In_2204,In_2323);
nor U3471 (N_3471,In_4241,In_4083);
nand U3472 (N_3472,In_425,In_1458);
xnor U3473 (N_3473,In_894,In_3379);
nand U3474 (N_3474,In_8,In_3481);
xnor U3475 (N_3475,In_3235,In_3357);
nand U3476 (N_3476,In_4508,In_1689);
and U3477 (N_3477,In_2983,In_4551);
xor U3478 (N_3478,In_4857,In_4552);
xor U3479 (N_3479,In_2670,In_4341);
or U3480 (N_3480,In_4891,In_24);
and U3481 (N_3481,In_2345,In_1075);
nor U3482 (N_3482,In_4606,In_4656);
nor U3483 (N_3483,In_973,In_2864);
and U3484 (N_3484,In_1185,In_1806);
or U3485 (N_3485,In_2467,In_1882);
nand U3486 (N_3486,In_833,In_3947);
nor U3487 (N_3487,In_1415,In_2537);
xor U3488 (N_3488,In_985,In_4734);
and U3489 (N_3489,In_3051,In_762);
or U3490 (N_3490,In_3719,In_1643);
nor U3491 (N_3491,In_4451,In_2658);
nor U3492 (N_3492,In_3571,In_1133);
nand U3493 (N_3493,In_3066,In_3526);
xor U3494 (N_3494,In_3777,In_1009);
xor U3495 (N_3495,In_4638,In_468);
xnor U3496 (N_3496,In_4232,In_3998);
and U3497 (N_3497,In_4711,In_186);
xnor U3498 (N_3498,In_4089,In_1056);
nand U3499 (N_3499,In_1132,In_1678);
nor U3500 (N_3500,In_1284,In_1404);
nor U3501 (N_3501,In_433,In_1880);
and U3502 (N_3502,In_8,In_4978);
and U3503 (N_3503,In_233,In_2098);
or U3504 (N_3504,In_1636,In_1000);
nor U3505 (N_3505,In_591,In_2195);
nor U3506 (N_3506,In_4618,In_46);
or U3507 (N_3507,In_2193,In_1735);
or U3508 (N_3508,In_2825,In_4127);
and U3509 (N_3509,In_4415,In_4411);
or U3510 (N_3510,In_419,In_2281);
nand U3511 (N_3511,In_937,In_4385);
nand U3512 (N_3512,In_2299,In_3982);
and U3513 (N_3513,In_1886,In_4431);
and U3514 (N_3514,In_4820,In_100);
and U3515 (N_3515,In_2625,In_905);
nor U3516 (N_3516,In_1586,In_1974);
and U3517 (N_3517,In_3330,In_3790);
nand U3518 (N_3518,In_705,In_3329);
nor U3519 (N_3519,In_1991,In_3549);
xor U3520 (N_3520,In_1874,In_2790);
nor U3521 (N_3521,In_3563,In_642);
or U3522 (N_3522,In_4001,In_1035);
nor U3523 (N_3523,In_1006,In_2088);
nor U3524 (N_3524,In_2116,In_2635);
or U3525 (N_3525,In_980,In_1281);
or U3526 (N_3526,In_2632,In_3707);
nand U3527 (N_3527,In_977,In_3308);
nor U3528 (N_3528,In_3526,In_3623);
or U3529 (N_3529,In_2157,In_3700);
xor U3530 (N_3530,In_4356,In_740);
xnor U3531 (N_3531,In_2058,In_3985);
nand U3532 (N_3532,In_4683,In_122);
nor U3533 (N_3533,In_408,In_2868);
xnor U3534 (N_3534,In_3582,In_3007);
xor U3535 (N_3535,In_440,In_4236);
nand U3536 (N_3536,In_1409,In_1856);
nor U3537 (N_3537,In_1125,In_1972);
nor U3538 (N_3538,In_2572,In_4566);
nor U3539 (N_3539,In_2008,In_1893);
nor U3540 (N_3540,In_242,In_457);
nand U3541 (N_3541,In_1389,In_621);
and U3542 (N_3542,In_413,In_556);
or U3543 (N_3543,In_1893,In_1473);
nor U3544 (N_3544,In_118,In_1383);
nor U3545 (N_3545,In_2269,In_4049);
xnor U3546 (N_3546,In_3454,In_3660);
nor U3547 (N_3547,In_1426,In_1734);
nand U3548 (N_3548,In_2767,In_1453);
nor U3549 (N_3549,In_3743,In_354);
nor U3550 (N_3550,In_3295,In_4628);
nor U3551 (N_3551,In_588,In_89);
and U3552 (N_3552,In_145,In_494);
or U3553 (N_3553,In_416,In_2334);
nand U3554 (N_3554,In_2324,In_3627);
or U3555 (N_3555,In_4372,In_1483);
and U3556 (N_3556,In_16,In_2103);
xor U3557 (N_3557,In_1882,In_3853);
nor U3558 (N_3558,In_4824,In_381);
and U3559 (N_3559,In_433,In_4094);
xnor U3560 (N_3560,In_3574,In_325);
and U3561 (N_3561,In_754,In_2338);
nand U3562 (N_3562,In_1480,In_4823);
xnor U3563 (N_3563,In_1918,In_2644);
and U3564 (N_3564,In_4498,In_3027);
and U3565 (N_3565,In_374,In_4900);
and U3566 (N_3566,In_3380,In_472);
or U3567 (N_3567,In_4439,In_99);
nand U3568 (N_3568,In_3812,In_3248);
nor U3569 (N_3569,In_2767,In_3032);
xnor U3570 (N_3570,In_2913,In_1001);
or U3571 (N_3571,In_3142,In_986);
nand U3572 (N_3572,In_901,In_1494);
and U3573 (N_3573,In_4093,In_3054);
xnor U3574 (N_3574,In_3656,In_2158);
nand U3575 (N_3575,In_433,In_3897);
nor U3576 (N_3576,In_2120,In_1284);
or U3577 (N_3577,In_48,In_2978);
xnor U3578 (N_3578,In_3703,In_3986);
xnor U3579 (N_3579,In_1556,In_70);
nand U3580 (N_3580,In_2390,In_2741);
or U3581 (N_3581,In_981,In_1163);
and U3582 (N_3582,In_1422,In_4197);
nor U3583 (N_3583,In_1368,In_387);
and U3584 (N_3584,In_2308,In_3178);
nand U3585 (N_3585,In_4968,In_1787);
nor U3586 (N_3586,In_4692,In_2779);
nor U3587 (N_3587,In_2170,In_4142);
xor U3588 (N_3588,In_1112,In_2182);
nand U3589 (N_3589,In_2066,In_2437);
or U3590 (N_3590,In_439,In_2110);
and U3591 (N_3591,In_3637,In_4247);
or U3592 (N_3592,In_3652,In_2313);
nor U3593 (N_3593,In_4925,In_2336);
or U3594 (N_3594,In_2522,In_3436);
and U3595 (N_3595,In_1851,In_996);
nand U3596 (N_3596,In_255,In_1993);
nand U3597 (N_3597,In_4790,In_3622);
nor U3598 (N_3598,In_1394,In_3336);
and U3599 (N_3599,In_1012,In_258);
or U3600 (N_3600,In_2345,In_2608);
nand U3601 (N_3601,In_311,In_1647);
nor U3602 (N_3602,In_521,In_3157);
or U3603 (N_3603,In_620,In_668);
and U3604 (N_3604,In_215,In_3857);
nand U3605 (N_3605,In_1889,In_3549);
nand U3606 (N_3606,In_4304,In_457);
xor U3607 (N_3607,In_2425,In_189);
xnor U3608 (N_3608,In_4712,In_4008);
or U3609 (N_3609,In_3254,In_4129);
nor U3610 (N_3610,In_2978,In_3741);
nand U3611 (N_3611,In_3949,In_4361);
xnor U3612 (N_3612,In_3587,In_4256);
or U3613 (N_3613,In_3504,In_3394);
or U3614 (N_3614,In_2171,In_46);
and U3615 (N_3615,In_1428,In_1289);
and U3616 (N_3616,In_893,In_3460);
and U3617 (N_3617,In_775,In_3385);
nand U3618 (N_3618,In_1979,In_235);
nand U3619 (N_3619,In_1732,In_3808);
nor U3620 (N_3620,In_3828,In_2969);
and U3621 (N_3621,In_3364,In_2128);
nand U3622 (N_3622,In_1866,In_1309);
and U3623 (N_3623,In_3827,In_1311);
nor U3624 (N_3624,In_38,In_1372);
and U3625 (N_3625,In_3102,In_4573);
or U3626 (N_3626,In_1051,In_4022);
nand U3627 (N_3627,In_1949,In_1119);
and U3628 (N_3628,In_3700,In_3717);
and U3629 (N_3629,In_2073,In_2472);
and U3630 (N_3630,In_405,In_1233);
nand U3631 (N_3631,In_4650,In_2165);
xor U3632 (N_3632,In_3965,In_4036);
nor U3633 (N_3633,In_800,In_402);
xnor U3634 (N_3634,In_1332,In_2964);
or U3635 (N_3635,In_36,In_2080);
and U3636 (N_3636,In_662,In_4778);
nand U3637 (N_3637,In_2132,In_2125);
and U3638 (N_3638,In_1764,In_2129);
nor U3639 (N_3639,In_1399,In_459);
xnor U3640 (N_3640,In_2154,In_4654);
nor U3641 (N_3641,In_2037,In_918);
and U3642 (N_3642,In_4107,In_3069);
nor U3643 (N_3643,In_4374,In_2315);
or U3644 (N_3644,In_4512,In_1102);
xor U3645 (N_3645,In_2244,In_1225);
xnor U3646 (N_3646,In_686,In_4594);
or U3647 (N_3647,In_3117,In_4785);
xor U3648 (N_3648,In_2919,In_1533);
xnor U3649 (N_3649,In_3408,In_4071);
xor U3650 (N_3650,In_3092,In_1712);
or U3651 (N_3651,In_293,In_1469);
nor U3652 (N_3652,In_3296,In_3393);
nand U3653 (N_3653,In_2479,In_4128);
xor U3654 (N_3654,In_1146,In_3118);
nand U3655 (N_3655,In_4876,In_4053);
or U3656 (N_3656,In_360,In_752);
and U3657 (N_3657,In_1394,In_2203);
nand U3658 (N_3658,In_286,In_2237);
nand U3659 (N_3659,In_1999,In_2848);
and U3660 (N_3660,In_737,In_3259);
nand U3661 (N_3661,In_2897,In_1447);
xor U3662 (N_3662,In_4590,In_3335);
xor U3663 (N_3663,In_1002,In_4763);
nand U3664 (N_3664,In_138,In_164);
xnor U3665 (N_3665,In_3876,In_3309);
xnor U3666 (N_3666,In_2852,In_1692);
xor U3667 (N_3667,In_3758,In_4002);
and U3668 (N_3668,In_1788,In_2468);
or U3669 (N_3669,In_1957,In_4854);
or U3670 (N_3670,In_4758,In_3037);
xor U3671 (N_3671,In_1283,In_2523);
nor U3672 (N_3672,In_1094,In_1159);
and U3673 (N_3673,In_4541,In_1331);
and U3674 (N_3674,In_3444,In_2326);
nor U3675 (N_3675,In_2489,In_2420);
xor U3676 (N_3676,In_2824,In_4214);
or U3677 (N_3677,In_3485,In_4885);
or U3678 (N_3678,In_4127,In_2177);
and U3679 (N_3679,In_4584,In_3835);
nor U3680 (N_3680,In_2796,In_48);
nor U3681 (N_3681,In_1069,In_1978);
xnor U3682 (N_3682,In_93,In_3225);
nand U3683 (N_3683,In_2506,In_1391);
nand U3684 (N_3684,In_2033,In_65);
or U3685 (N_3685,In_4919,In_3585);
xnor U3686 (N_3686,In_2997,In_4034);
and U3687 (N_3687,In_2685,In_3296);
xor U3688 (N_3688,In_120,In_2561);
nor U3689 (N_3689,In_625,In_2533);
and U3690 (N_3690,In_3283,In_1545);
nor U3691 (N_3691,In_2734,In_1213);
nor U3692 (N_3692,In_3924,In_4080);
and U3693 (N_3693,In_4802,In_4287);
nor U3694 (N_3694,In_1770,In_4298);
nor U3695 (N_3695,In_39,In_731);
nand U3696 (N_3696,In_380,In_4739);
or U3697 (N_3697,In_203,In_997);
and U3698 (N_3698,In_174,In_4022);
xnor U3699 (N_3699,In_4080,In_3233);
or U3700 (N_3700,In_3688,In_453);
or U3701 (N_3701,In_4073,In_2656);
xor U3702 (N_3702,In_3197,In_1833);
nor U3703 (N_3703,In_1881,In_1463);
or U3704 (N_3704,In_856,In_3537);
and U3705 (N_3705,In_3956,In_3960);
nand U3706 (N_3706,In_2145,In_3029);
nand U3707 (N_3707,In_3801,In_1339);
nor U3708 (N_3708,In_558,In_2352);
nand U3709 (N_3709,In_4740,In_3052);
xor U3710 (N_3710,In_2104,In_4730);
xnor U3711 (N_3711,In_3483,In_4932);
or U3712 (N_3712,In_3354,In_2876);
xnor U3713 (N_3713,In_2789,In_1590);
xor U3714 (N_3714,In_2311,In_2881);
xor U3715 (N_3715,In_125,In_3957);
xnor U3716 (N_3716,In_1169,In_4936);
nand U3717 (N_3717,In_3087,In_701);
and U3718 (N_3718,In_3674,In_1356);
and U3719 (N_3719,In_4191,In_4510);
and U3720 (N_3720,In_3702,In_1041);
or U3721 (N_3721,In_2851,In_3477);
and U3722 (N_3722,In_4615,In_3852);
or U3723 (N_3723,In_3914,In_2230);
and U3724 (N_3724,In_2370,In_1699);
or U3725 (N_3725,In_411,In_1108);
or U3726 (N_3726,In_2454,In_3526);
or U3727 (N_3727,In_3215,In_2487);
xnor U3728 (N_3728,In_3100,In_702);
nand U3729 (N_3729,In_1779,In_3187);
or U3730 (N_3730,In_3914,In_1492);
or U3731 (N_3731,In_3893,In_3384);
nor U3732 (N_3732,In_4113,In_722);
or U3733 (N_3733,In_4245,In_1961);
or U3734 (N_3734,In_840,In_1650);
nand U3735 (N_3735,In_1283,In_1938);
nand U3736 (N_3736,In_4772,In_912);
nor U3737 (N_3737,In_2876,In_3177);
or U3738 (N_3738,In_257,In_3584);
nor U3739 (N_3739,In_222,In_1973);
and U3740 (N_3740,In_2408,In_3277);
or U3741 (N_3741,In_1159,In_3781);
nor U3742 (N_3742,In_1087,In_4667);
or U3743 (N_3743,In_4756,In_2710);
or U3744 (N_3744,In_4853,In_3800);
and U3745 (N_3745,In_1078,In_4894);
and U3746 (N_3746,In_4062,In_2029);
or U3747 (N_3747,In_1933,In_4810);
nor U3748 (N_3748,In_882,In_772);
nor U3749 (N_3749,In_2210,In_1805);
or U3750 (N_3750,In_3147,In_4001);
nor U3751 (N_3751,In_956,In_3336);
xnor U3752 (N_3752,In_4719,In_2883);
nand U3753 (N_3753,In_993,In_1725);
nor U3754 (N_3754,In_4155,In_2906);
and U3755 (N_3755,In_399,In_2118);
nor U3756 (N_3756,In_2435,In_4899);
and U3757 (N_3757,In_870,In_3463);
nor U3758 (N_3758,In_662,In_240);
or U3759 (N_3759,In_1292,In_3765);
or U3760 (N_3760,In_1465,In_2779);
xor U3761 (N_3761,In_4223,In_2973);
xnor U3762 (N_3762,In_3089,In_1709);
nand U3763 (N_3763,In_3062,In_4873);
nor U3764 (N_3764,In_3416,In_854);
nand U3765 (N_3765,In_559,In_1100);
or U3766 (N_3766,In_713,In_3991);
and U3767 (N_3767,In_4350,In_836);
and U3768 (N_3768,In_2311,In_42);
nor U3769 (N_3769,In_3620,In_3086);
and U3770 (N_3770,In_3171,In_3974);
or U3771 (N_3771,In_596,In_1500);
or U3772 (N_3772,In_2974,In_4546);
or U3773 (N_3773,In_4176,In_1852);
xor U3774 (N_3774,In_1713,In_1024);
or U3775 (N_3775,In_4607,In_962);
and U3776 (N_3776,In_3582,In_521);
nand U3777 (N_3777,In_93,In_2595);
or U3778 (N_3778,In_3528,In_2613);
nand U3779 (N_3779,In_475,In_1326);
xnor U3780 (N_3780,In_221,In_3902);
or U3781 (N_3781,In_1170,In_3699);
or U3782 (N_3782,In_3868,In_4747);
nor U3783 (N_3783,In_2819,In_61);
and U3784 (N_3784,In_2686,In_4100);
nand U3785 (N_3785,In_714,In_2335);
nor U3786 (N_3786,In_4658,In_3356);
xnor U3787 (N_3787,In_3362,In_1341);
xor U3788 (N_3788,In_4463,In_4737);
and U3789 (N_3789,In_336,In_4464);
nand U3790 (N_3790,In_3463,In_4691);
xor U3791 (N_3791,In_3450,In_1738);
nor U3792 (N_3792,In_4944,In_3973);
nand U3793 (N_3793,In_3095,In_4097);
or U3794 (N_3794,In_2362,In_1743);
nor U3795 (N_3795,In_1971,In_236);
nand U3796 (N_3796,In_1621,In_3489);
or U3797 (N_3797,In_3909,In_3802);
xnor U3798 (N_3798,In_3279,In_2279);
nand U3799 (N_3799,In_1974,In_4588);
nor U3800 (N_3800,In_1118,In_4405);
nand U3801 (N_3801,In_2433,In_4358);
nand U3802 (N_3802,In_1955,In_2267);
nor U3803 (N_3803,In_2870,In_1780);
nor U3804 (N_3804,In_3358,In_882);
and U3805 (N_3805,In_1904,In_397);
or U3806 (N_3806,In_2085,In_1051);
nor U3807 (N_3807,In_2174,In_603);
or U3808 (N_3808,In_328,In_1041);
and U3809 (N_3809,In_4287,In_639);
nand U3810 (N_3810,In_365,In_4859);
and U3811 (N_3811,In_1357,In_224);
and U3812 (N_3812,In_156,In_676);
or U3813 (N_3813,In_3427,In_1813);
and U3814 (N_3814,In_3122,In_2689);
and U3815 (N_3815,In_4753,In_3830);
or U3816 (N_3816,In_2395,In_1533);
nor U3817 (N_3817,In_1848,In_1248);
and U3818 (N_3818,In_3466,In_3562);
nor U3819 (N_3819,In_867,In_2979);
and U3820 (N_3820,In_3647,In_3312);
nor U3821 (N_3821,In_1662,In_2474);
nor U3822 (N_3822,In_1437,In_1287);
nor U3823 (N_3823,In_2322,In_755);
or U3824 (N_3824,In_2517,In_2987);
and U3825 (N_3825,In_4111,In_2920);
nor U3826 (N_3826,In_3153,In_4211);
nand U3827 (N_3827,In_3210,In_1578);
xnor U3828 (N_3828,In_2864,In_4839);
nor U3829 (N_3829,In_4558,In_712);
nand U3830 (N_3830,In_2330,In_4094);
nand U3831 (N_3831,In_3689,In_4536);
xnor U3832 (N_3832,In_1717,In_2783);
or U3833 (N_3833,In_2948,In_2592);
or U3834 (N_3834,In_761,In_3096);
nand U3835 (N_3835,In_1429,In_914);
nor U3836 (N_3836,In_3545,In_3975);
nand U3837 (N_3837,In_4711,In_1913);
xnor U3838 (N_3838,In_4566,In_4749);
nor U3839 (N_3839,In_4062,In_3461);
and U3840 (N_3840,In_3593,In_4062);
nor U3841 (N_3841,In_225,In_2384);
and U3842 (N_3842,In_2135,In_1608);
xor U3843 (N_3843,In_3901,In_3037);
nand U3844 (N_3844,In_4391,In_4746);
and U3845 (N_3845,In_3785,In_2405);
nand U3846 (N_3846,In_2490,In_2459);
and U3847 (N_3847,In_4790,In_4374);
and U3848 (N_3848,In_2237,In_3126);
xor U3849 (N_3849,In_4103,In_1123);
or U3850 (N_3850,In_668,In_1100);
and U3851 (N_3851,In_2758,In_4374);
nor U3852 (N_3852,In_1324,In_2566);
nor U3853 (N_3853,In_4480,In_504);
or U3854 (N_3854,In_2754,In_752);
nand U3855 (N_3855,In_4772,In_4484);
or U3856 (N_3856,In_2028,In_576);
nand U3857 (N_3857,In_2429,In_2821);
and U3858 (N_3858,In_333,In_937);
nand U3859 (N_3859,In_3354,In_380);
or U3860 (N_3860,In_4235,In_3158);
nand U3861 (N_3861,In_1606,In_3501);
nand U3862 (N_3862,In_1912,In_643);
or U3863 (N_3863,In_4547,In_2366);
nor U3864 (N_3864,In_564,In_4468);
nand U3865 (N_3865,In_4172,In_1574);
and U3866 (N_3866,In_1503,In_1860);
and U3867 (N_3867,In_1454,In_1432);
xor U3868 (N_3868,In_2367,In_4060);
and U3869 (N_3869,In_2726,In_3073);
or U3870 (N_3870,In_4154,In_732);
xor U3871 (N_3871,In_138,In_2808);
xnor U3872 (N_3872,In_4326,In_100);
xor U3873 (N_3873,In_2651,In_2475);
nand U3874 (N_3874,In_3441,In_435);
nor U3875 (N_3875,In_942,In_4134);
nand U3876 (N_3876,In_191,In_1559);
xnor U3877 (N_3877,In_4636,In_2671);
nor U3878 (N_3878,In_2210,In_3580);
and U3879 (N_3879,In_2674,In_4004);
or U3880 (N_3880,In_978,In_4073);
xnor U3881 (N_3881,In_1809,In_1850);
nand U3882 (N_3882,In_21,In_1371);
nand U3883 (N_3883,In_100,In_3651);
or U3884 (N_3884,In_3668,In_2646);
nor U3885 (N_3885,In_1181,In_1801);
or U3886 (N_3886,In_863,In_816);
nor U3887 (N_3887,In_4887,In_1074);
xnor U3888 (N_3888,In_401,In_3068);
nand U3889 (N_3889,In_657,In_1287);
xnor U3890 (N_3890,In_1493,In_1032);
nor U3891 (N_3891,In_465,In_1701);
xor U3892 (N_3892,In_2619,In_4039);
or U3893 (N_3893,In_1818,In_3066);
nor U3894 (N_3894,In_2293,In_3821);
nand U3895 (N_3895,In_2287,In_124);
nor U3896 (N_3896,In_858,In_4486);
xnor U3897 (N_3897,In_2004,In_560);
nor U3898 (N_3898,In_427,In_1205);
xnor U3899 (N_3899,In_2657,In_1044);
xnor U3900 (N_3900,In_138,In_1298);
nor U3901 (N_3901,In_486,In_1668);
nand U3902 (N_3902,In_521,In_2300);
or U3903 (N_3903,In_1451,In_3757);
xnor U3904 (N_3904,In_4313,In_104);
nand U3905 (N_3905,In_773,In_320);
nor U3906 (N_3906,In_4898,In_3143);
and U3907 (N_3907,In_2527,In_357);
and U3908 (N_3908,In_4582,In_2439);
nor U3909 (N_3909,In_168,In_1798);
and U3910 (N_3910,In_3779,In_4836);
nand U3911 (N_3911,In_4218,In_197);
and U3912 (N_3912,In_2587,In_538);
nor U3913 (N_3913,In_2753,In_2741);
nand U3914 (N_3914,In_3248,In_2330);
and U3915 (N_3915,In_1252,In_1967);
and U3916 (N_3916,In_4821,In_4871);
or U3917 (N_3917,In_2130,In_3256);
and U3918 (N_3918,In_2333,In_1939);
xnor U3919 (N_3919,In_4716,In_3135);
xnor U3920 (N_3920,In_3937,In_4122);
xor U3921 (N_3921,In_1172,In_4030);
and U3922 (N_3922,In_2699,In_4286);
or U3923 (N_3923,In_4429,In_2173);
nor U3924 (N_3924,In_2892,In_2619);
xor U3925 (N_3925,In_1491,In_3259);
and U3926 (N_3926,In_4588,In_4108);
nand U3927 (N_3927,In_2713,In_4779);
or U3928 (N_3928,In_4905,In_203);
nand U3929 (N_3929,In_85,In_1421);
and U3930 (N_3930,In_3410,In_1124);
nand U3931 (N_3931,In_2043,In_2511);
nand U3932 (N_3932,In_1639,In_217);
nor U3933 (N_3933,In_3114,In_3035);
xor U3934 (N_3934,In_497,In_3031);
or U3935 (N_3935,In_4671,In_1689);
nor U3936 (N_3936,In_2937,In_1487);
or U3937 (N_3937,In_4864,In_1312);
or U3938 (N_3938,In_14,In_204);
nand U3939 (N_3939,In_45,In_3052);
and U3940 (N_3940,In_1092,In_2257);
or U3941 (N_3941,In_2939,In_2052);
and U3942 (N_3942,In_4461,In_4850);
xor U3943 (N_3943,In_105,In_2365);
nand U3944 (N_3944,In_4296,In_2877);
xor U3945 (N_3945,In_2477,In_1751);
nor U3946 (N_3946,In_3303,In_3905);
and U3947 (N_3947,In_1207,In_178);
or U3948 (N_3948,In_2883,In_3947);
nand U3949 (N_3949,In_3507,In_3998);
nor U3950 (N_3950,In_344,In_4515);
or U3951 (N_3951,In_4832,In_2752);
xnor U3952 (N_3952,In_1722,In_4040);
nor U3953 (N_3953,In_3832,In_1136);
nor U3954 (N_3954,In_1993,In_3748);
and U3955 (N_3955,In_102,In_4158);
or U3956 (N_3956,In_1417,In_4314);
and U3957 (N_3957,In_2709,In_830);
nand U3958 (N_3958,In_2757,In_3223);
or U3959 (N_3959,In_3581,In_3182);
nand U3960 (N_3960,In_1559,In_2197);
or U3961 (N_3961,In_1453,In_3968);
xnor U3962 (N_3962,In_4409,In_1946);
nand U3963 (N_3963,In_1329,In_1418);
xnor U3964 (N_3964,In_800,In_2464);
nand U3965 (N_3965,In_4209,In_2133);
and U3966 (N_3966,In_2769,In_1915);
or U3967 (N_3967,In_3765,In_2699);
nor U3968 (N_3968,In_384,In_3319);
nand U3969 (N_3969,In_313,In_3489);
nand U3970 (N_3970,In_3205,In_393);
nor U3971 (N_3971,In_122,In_1312);
xnor U3972 (N_3972,In_2354,In_2296);
and U3973 (N_3973,In_184,In_92);
or U3974 (N_3974,In_4984,In_4596);
or U3975 (N_3975,In_3575,In_3491);
and U3976 (N_3976,In_1352,In_4039);
and U3977 (N_3977,In_2264,In_2073);
nand U3978 (N_3978,In_4195,In_1110);
xnor U3979 (N_3979,In_2902,In_3050);
or U3980 (N_3980,In_2345,In_36);
nor U3981 (N_3981,In_3266,In_3475);
and U3982 (N_3982,In_1557,In_3108);
nand U3983 (N_3983,In_4855,In_3470);
or U3984 (N_3984,In_3900,In_3981);
nor U3985 (N_3985,In_2960,In_3062);
nand U3986 (N_3986,In_2588,In_1586);
xnor U3987 (N_3987,In_1092,In_1994);
and U3988 (N_3988,In_2922,In_2251);
xor U3989 (N_3989,In_362,In_1799);
and U3990 (N_3990,In_1464,In_1301);
nor U3991 (N_3991,In_681,In_4406);
xor U3992 (N_3992,In_4525,In_1610);
nand U3993 (N_3993,In_4488,In_4635);
or U3994 (N_3994,In_1193,In_1764);
nand U3995 (N_3995,In_2102,In_4903);
nand U3996 (N_3996,In_4575,In_1914);
and U3997 (N_3997,In_1894,In_2063);
nor U3998 (N_3998,In_4610,In_69);
xor U3999 (N_3999,In_3444,In_539);
nor U4000 (N_4000,In_796,In_4547);
and U4001 (N_4001,In_1797,In_4151);
and U4002 (N_4002,In_3511,In_598);
nor U4003 (N_4003,In_1153,In_411);
nand U4004 (N_4004,In_1172,In_1099);
xnor U4005 (N_4005,In_409,In_942);
nand U4006 (N_4006,In_4743,In_3269);
nand U4007 (N_4007,In_936,In_1205);
and U4008 (N_4008,In_257,In_555);
xnor U4009 (N_4009,In_4624,In_4183);
nor U4010 (N_4010,In_2102,In_973);
xnor U4011 (N_4011,In_3402,In_3217);
xor U4012 (N_4012,In_1956,In_4790);
and U4013 (N_4013,In_4506,In_462);
and U4014 (N_4014,In_2462,In_1672);
xor U4015 (N_4015,In_754,In_1325);
or U4016 (N_4016,In_1653,In_3610);
and U4017 (N_4017,In_3480,In_924);
or U4018 (N_4018,In_3531,In_4301);
or U4019 (N_4019,In_2835,In_4402);
and U4020 (N_4020,In_2384,In_4472);
and U4021 (N_4021,In_3028,In_3865);
nand U4022 (N_4022,In_3837,In_4682);
nand U4023 (N_4023,In_1141,In_1036);
nor U4024 (N_4024,In_2438,In_1042);
nand U4025 (N_4025,In_90,In_1798);
nand U4026 (N_4026,In_3093,In_2680);
and U4027 (N_4027,In_2373,In_3266);
nand U4028 (N_4028,In_2932,In_1135);
and U4029 (N_4029,In_2072,In_3941);
xor U4030 (N_4030,In_4313,In_1871);
nor U4031 (N_4031,In_3398,In_1345);
nand U4032 (N_4032,In_2247,In_416);
or U4033 (N_4033,In_992,In_4457);
nor U4034 (N_4034,In_1540,In_4509);
and U4035 (N_4035,In_613,In_853);
and U4036 (N_4036,In_1748,In_2914);
nor U4037 (N_4037,In_4809,In_3546);
xnor U4038 (N_4038,In_3939,In_209);
nor U4039 (N_4039,In_2780,In_4694);
nand U4040 (N_4040,In_3690,In_1461);
or U4041 (N_4041,In_3520,In_496);
nand U4042 (N_4042,In_3722,In_2265);
nand U4043 (N_4043,In_56,In_1360);
xor U4044 (N_4044,In_2392,In_4011);
nand U4045 (N_4045,In_2464,In_897);
or U4046 (N_4046,In_3117,In_2690);
nand U4047 (N_4047,In_3400,In_4480);
xor U4048 (N_4048,In_2046,In_3652);
and U4049 (N_4049,In_2445,In_3590);
xor U4050 (N_4050,In_624,In_379);
or U4051 (N_4051,In_4681,In_4809);
and U4052 (N_4052,In_2213,In_600);
and U4053 (N_4053,In_4066,In_425);
xnor U4054 (N_4054,In_1943,In_4129);
or U4055 (N_4055,In_4922,In_4634);
nand U4056 (N_4056,In_2865,In_1165);
nor U4057 (N_4057,In_695,In_1615);
or U4058 (N_4058,In_548,In_569);
or U4059 (N_4059,In_2940,In_1250);
xor U4060 (N_4060,In_3010,In_3601);
or U4061 (N_4061,In_2519,In_3600);
nand U4062 (N_4062,In_3631,In_100);
or U4063 (N_4063,In_645,In_4549);
xnor U4064 (N_4064,In_2194,In_1583);
or U4065 (N_4065,In_3859,In_686);
nor U4066 (N_4066,In_1694,In_4593);
and U4067 (N_4067,In_1284,In_2401);
and U4068 (N_4068,In_2315,In_3066);
nor U4069 (N_4069,In_1252,In_726);
nand U4070 (N_4070,In_1398,In_3340);
xnor U4071 (N_4071,In_1499,In_622);
and U4072 (N_4072,In_524,In_4616);
and U4073 (N_4073,In_2908,In_272);
xnor U4074 (N_4074,In_3757,In_984);
or U4075 (N_4075,In_2501,In_2152);
and U4076 (N_4076,In_4907,In_4156);
and U4077 (N_4077,In_4063,In_233);
xnor U4078 (N_4078,In_4829,In_4);
and U4079 (N_4079,In_1001,In_2620);
xor U4080 (N_4080,In_4772,In_447);
nand U4081 (N_4081,In_3160,In_648);
or U4082 (N_4082,In_3687,In_2577);
and U4083 (N_4083,In_1423,In_2748);
nand U4084 (N_4084,In_4429,In_4931);
nor U4085 (N_4085,In_174,In_2420);
or U4086 (N_4086,In_546,In_1236);
or U4087 (N_4087,In_3982,In_747);
nor U4088 (N_4088,In_0,In_1798);
and U4089 (N_4089,In_894,In_963);
nor U4090 (N_4090,In_3854,In_4973);
xnor U4091 (N_4091,In_2483,In_4148);
or U4092 (N_4092,In_2394,In_3534);
and U4093 (N_4093,In_391,In_2159);
or U4094 (N_4094,In_2983,In_2052);
and U4095 (N_4095,In_1509,In_2068);
nor U4096 (N_4096,In_1641,In_1374);
xnor U4097 (N_4097,In_3906,In_1512);
xnor U4098 (N_4098,In_2869,In_3718);
nand U4099 (N_4099,In_3472,In_4190);
or U4100 (N_4100,In_1652,In_75);
nand U4101 (N_4101,In_4805,In_4022);
nor U4102 (N_4102,In_2595,In_1822);
or U4103 (N_4103,In_1896,In_3419);
or U4104 (N_4104,In_3164,In_4351);
nand U4105 (N_4105,In_3382,In_3664);
xnor U4106 (N_4106,In_2959,In_3962);
nand U4107 (N_4107,In_3924,In_1888);
nand U4108 (N_4108,In_2465,In_1404);
and U4109 (N_4109,In_3036,In_2879);
or U4110 (N_4110,In_3001,In_1602);
xnor U4111 (N_4111,In_1065,In_501);
nand U4112 (N_4112,In_2498,In_770);
xnor U4113 (N_4113,In_4994,In_2656);
xor U4114 (N_4114,In_3663,In_3894);
xor U4115 (N_4115,In_1473,In_1231);
or U4116 (N_4116,In_259,In_1282);
and U4117 (N_4117,In_479,In_4941);
xor U4118 (N_4118,In_2931,In_467);
and U4119 (N_4119,In_851,In_4595);
nor U4120 (N_4120,In_198,In_4374);
nand U4121 (N_4121,In_4777,In_3315);
nor U4122 (N_4122,In_2080,In_4176);
or U4123 (N_4123,In_4032,In_1723);
nand U4124 (N_4124,In_4988,In_2632);
xnor U4125 (N_4125,In_130,In_3519);
or U4126 (N_4126,In_638,In_759);
nand U4127 (N_4127,In_4044,In_2348);
nand U4128 (N_4128,In_4829,In_4277);
nand U4129 (N_4129,In_1570,In_314);
nand U4130 (N_4130,In_3346,In_2316);
xnor U4131 (N_4131,In_4937,In_25);
and U4132 (N_4132,In_2454,In_3664);
or U4133 (N_4133,In_4613,In_1972);
and U4134 (N_4134,In_2785,In_3716);
nand U4135 (N_4135,In_3935,In_2590);
and U4136 (N_4136,In_4012,In_421);
or U4137 (N_4137,In_2913,In_3731);
or U4138 (N_4138,In_2685,In_2516);
nor U4139 (N_4139,In_4460,In_2925);
or U4140 (N_4140,In_1888,In_2386);
xnor U4141 (N_4141,In_2205,In_2936);
nor U4142 (N_4142,In_4113,In_211);
nor U4143 (N_4143,In_1215,In_490);
xor U4144 (N_4144,In_1902,In_3035);
or U4145 (N_4145,In_3350,In_2194);
xor U4146 (N_4146,In_1122,In_4344);
nor U4147 (N_4147,In_3120,In_420);
nor U4148 (N_4148,In_3703,In_3531);
nor U4149 (N_4149,In_248,In_1715);
or U4150 (N_4150,In_4604,In_306);
nor U4151 (N_4151,In_3336,In_4337);
nand U4152 (N_4152,In_2902,In_2144);
nand U4153 (N_4153,In_4011,In_3549);
xor U4154 (N_4154,In_2778,In_504);
nand U4155 (N_4155,In_1646,In_4873);
and U4156 (N_4156,In_2794,In_2211);
nor U4157 (N_4157,In_4033,In_3413);
or U4158 (N_4158,In_2274,In_3394);
or U4159 (N_4159,In_4566,In_551);
xor U4160 (N_4160,In_317,In_4590);
nor U4161 (N_4161,In_911,In_2097);
or U4162 (N_4162,In_4158,In_755);
nor U4163 (N_4163,In_3146,In_2461);
or U4164 (N_4164,In_4849,In_4553);
and U4165 (N_4165,In_2282,In_3331);
or U4166 (N_4166,In_4625,In_4323);
nand U4167 (N_4167,In_805,In_2812);
or U4168 (N_4168,In_4281,In_599);
or U4169 (N_4169,In_1395,In_3648);
and U4170 (N_4170,In_4738,In_216);
xor U4171 (N_4171,In_841,In_1667);
xnor U4172 (N_4172,In_3880,In_1950);
xor U4173 (N_4173,In_2707,In_23);
xnor U4174 (N_4174,In_940,In_4919);
and U4175 (N_4175,In_2641,In_4926);
nand U4176 (N_4176,In_3448,In_112);
nor U4177 (N_4177,In_795,In_4396);
xor U4178 (N_4178,In_549,In_1925);
and U4179 (N_4179,In_3138,In_3056);
nand U4180 (N_4180,In_408,In_1904);
nor U4181 (N_4181,In_897,In_1214);
xnor U4182 (N_4182,In_4759,In_4232);
or U4183 (N_4183,In_902,In_3141);
nand U4184 (N_4184,In_3993,In_4233);
and U4185 (N_4185,In_2078,In_1090);
nand U4186 (N_4186,In_91,In_4275);
xor U4187 (N_4187,In_2263,In_190);
nand U4188 (N_4188,In_4625,In_1820);
and U4189 (N_4189,In_1646,In_3943);
nor U4190 (N_4190,In_1507,In_2075);
nand U4191 (N_4191,In_3261,In_2970);
nor U4192 (N_4192,In_3792,In_2589);
or U4193 (N_4193,In_4490,In_2270);
xnor U4194 (N_4194,In_2790,In_4376);
nand U4195 (N_4195,In_712,In_2682);
or U4196 (N_4196,In_502,In_2481);
xnor U4197 (N_4197,In_653,In_1409);
xor U4198 (N_4198,In_2410,In_712);
xor U4199 (N_4199,In_3281,In_4354);
nor U4200 (N_4200,In_3407,In_1334);
and U4201 (N_4201,In_845,In_4576);
xor U4202 (N_4202,In_1407,In_503);
nor U4203 (N_4203,In_3099,In_4843);
xnor U4204 (N_4204,In_2101,In_3982);
and U4205 (N_4205,In_3969,In_2228);
xor U4206 (N_4206,In_3181,In_2852);
and U4207 (N_4207,In_2203,In_994);
nand U4208 (N_4208,In_1558,In_4424);
and U4209 (N_4209,In_2103,In_4152);
or U4210 (N_4210,In_1589,In_777);
or U4211 (N_4211,In_1804,In_1483);
or U4212 (N_4212,In_4916,In_3620);
or U4213 (N_4213,In_3016,In_252);
nor U4214 (N_4214,In_3172,In_4514);
or U4215 (N_4215,In_674,In_3901);
and U4216 (N_4216,In_1496,In_3202);
or U4217 (N_4217,In_2608,In_2223);
nor U4218 (N_4218,In_4991,In_1804);
nor U4219 (N_4219,In_3850,In_4533);
or U4220 (N_4220,In_1653,In_996);
nand U4221 (N_4221,In_19,In_433);
and U4222 (N_4222,In_3264,In_3795);
and U4223 (N_4223,In_1246,In_793);
and U4224 (N_4224,In_2410,In_4530);
xnor U4225 (N_4225,In_666,In_615);
xnor U4226 (N_4226,In_4759,In_2221);
and U4227 (N_4227,In_877,In_871);
or U4228 (N_4228,In_4131,In_85);
xor U4229 (N_4229,In_356,In_3436);
nand U4230 (N_4230,In_1986,In_4006);
nand U4231 (N_4231,In_2816,In_467);
and U4232 (N_4232,In_1428,In_1295);
nor U4233 (N_4233,In_3962,In_2270);
xor U4234 (N_4234,In_1671,In_254);
xor U4235 (N_4235,In_4830,In_3043);
nor U4236 (N_4236,In_4903,In_3518);
or U4237 (N_4237,In_4393,In_3570);
nand U4238 (N_4238,In_2447,In_1933);
or U4239 (N_4239,In_1779,In_1404);
and U4240 (N_4240,In_461,In_4270);
and U4241 (N_4241,In_2842,In_4460);
nor U4242 (N_4242,In_3037,In_2770);
nand U4243 (N_4243,In_296,In_84);
nand U4244 (N_4244,In_4338,In_215);
or U4245 (N_4245,In_3644,In_3697);
nand U4246 (N_4246,In_3315,In_551);
or U4247 (N_4247,In_4496,In_2565);
nor U4248 (N_4248,In_4860,In_1440);
nand U4249 (N_4249,In_3076,In_220);
nor U4250 (N_4250,In_1056,In_145);
and U4251 (N_4251,In_4441,In_2899);
or U4252 (N_4252,In_4570,In_686);
xor U4253 (N_4253,In_796,In_301);
and U4254 (N_4254,In_512,In_3355);
nand U4255 (N_4255,In_913,In_4236);
xnor U4256 (N_4256,In_1420,In_566);
nand U4257 (N_4257,In_4155,In_2034);
xnor U4258 (N_4258,In_4620,In_4214);
nand U4259 (N_4259,In_2691,In_167);
xor U4260 (N_4260,In_1714,In_843);
nand U4261 (N_4261,In_21,In_1393);
xnor U4262 (N_4262,In_4536,In_4854);
nand U4263 (N_4263,In_13,In_1713);
nor U4264 (N_4264,In_4935,In_1720);
xnor U4265 (N_4265,In_1614,In_665);
or U4266 (N_4266,In_2786,In_3595);
nand U4267 (N_4267,In_3258,In_366);
nand U4268 (N_4268,In_2146,In_4984);
or U4269 (N_4269,In_2108,In_163);
nor U4270 (N_4270,In_2474,In_3382);
and U4271 (N_4271,In_4139,In_4718);
xor U4272 (N_4272,In_137,In_2590);
nor U4273 (N_4273,In_1506,In_4793);
xnor U4274 (N_4274,In_3599,In_1275);
and U4275 (N_4275,In_859,In_38);
or U4276 (N_4276,In_2760,In_1888);
xnor U4277 (N_4277,In_2053,In_584);
nand U4278 (N_4278,In_4161,In_4395);
and U4279 (N_4279,In_2764,In_4291);
xnor U4280 (N_4280,In_2814,In_2838);
and U4281 (N_4281,In_627,In_3353);
xor U4282 (N_4282,In_4074,In_1476);
nor U4283 (N_4283,In_3261,In_2542);
nor U4284 (N_4284,In_4062,In_649);
xnor U4285 (N_4285,In_3018,In_3813);
nand U4286 (N_4286,In_362,In_2670);
nand U4287 (N_4287,In_2353,In_1152);
and U4288 (N_4288,In_1226,In_167);
nand U4289 (N_4289,In_2252,In_1132);
nor U4290 (N_4290,In_2230,In_4229);
xor U4291 (N_4291,In_2264,In_3846);
or U4292 (N_4292,In_3968,In_2405);
nor U4293 (N_4293,In_3021,In_3690);
nand U4294 (N_4294,In_1428,In_4896);
or U4295 (N_4295,In_2792,In_848);
nor U4296 (N_4296,In_2343,In_1851);
and U4297 (N_4297,In_157,In_2119);
and U4298 (N_4298,In_4272,In_3989);
and U4299 (N_4299,In_3191,In_1712);
or U4300 (N_4300,In_866,In_3715);
xor U4301 (N_4301,In_1837,In_18);
and U4302 (N_4302,In_3721,In_1865);
and U4303 (N_4303,In_3271,In_211);
xnor U4304 (N_4304,In_3099,In_957);
or U4305 (N_4305,In_2234,In_1836);
and U4306 (N_4306,In_1528,In_554);
nand U4307 (N_4307,In_4224,In_937);
xor U4308 (N_4308,In_776,In_83);
nor U4309 (N_4309,In_2799,In_3764);
xnor U4310 (N_4310,In_3035,In_2902);
nor U4311 (N_4311,In_3767,In_1208);
and U4312 (N_4312,In_953,In_3995);
nor U4313 (N_4313,In_487,In_1291);
xor U4314 (N_4314,In_4244,In_1362);
xor U4315 (N_4315,In_247,In_1292);
and U4316 (N_4316,In_630,In_3297);
xnor U4317 (N_4317,In_2929,In_2630);
nor U4318 (N_4318,In_95,In_1715);
nor U4319 (N_4319,In_3404,In_1586);
and U4320 (N_4320,In_1041,In_26);
or U4321 (N_4321,In_1960,In_3472);
and U4322 (N_4322,In_4543,In_4523);
xor U4323 (N_4323,In_1067,In_2982);
xor U4324 (N_4324,In_206,In_1812);
xor U4325 (N_4325,In_4330,In_3517);
nor U4326 (N_4326,In_207,In_1572);
xor U4327 (N_4327,In_707,In_131);
nor U4328 (N_4328,In_2882,In_3190);
nor U4329 (N_4329,In_2011,In_2573);
or U4330 (N_4330,In_3545,In_4006);
nand U4331 (N_4331,In_673,In_2711);
nand U4332 (N_4332,In_70,In_3649);
nor U4333 (N_4333,In_2239,In_3793);
or U4334 (N_4334,In_953,In_2906);
nor U4335 (N_4335,In_1334,In_3729);
nor U4336 (N_4336,In_3982,In_993);
xor U4337 (N_4337,In_3683,In_558);
xor U4338 (N_4338,In_3609,In_3749);
nand U4339 (N_4339,In_1064,In_1521);
or U4340 (N_4340,In_1111,In_4193);
or U4341 (N_4341,In_4066,In_3146);
nor U4342 (N_4342,In_2905,In_4712);
nor U4343 (N_4343,In_1045,In_2888);
xor U4344 (N_4344,In_764,In_2092);
or U4345 (N_4345,In_4730,In_2279);
nor U4346 (N_4346,In_3269,In_640);
nand U4347 (N_4347,In_64,In_2209);
nand U4348 (N_4348,In_4737,In_1521);
and U4349 (N_4349,In_1120,In_959);
xor U4350 (N_4350,In_2253,In_2663);
nor U4351 (N_4351,In_3943,In_4401);
or U4352 (N_4352,In_25,In_3389);
and U4353 (N_4353,In_4732,In_575);
or U4354 (N_4354,In_207,In_441);
xor U4355 (N_4355,In_2005,In_888);
nor U4356 (N_4356,In_2277,In_387);
xnor U4357 (N_4357,In_2028,In_2049);
and U4358 (N_4358,In_720,In_4401);
or U4359 (N_4359,In_206,In_1621);
xnor U4360 (N_4360,In_3396,In_3374);
nand U4361 (N_4361,In_3834,In_4301);
xnor U4362 (N_4362,In_2284,In_3162);
nand U4363 (N_4363,In_2216,In_3827);
nand U4364 (N_4364,In_479,In_2356);
or U4365 (N_4365,In_4142,In_1897);
nand U4366 (N_4366,In_2250,In_2018);
xor U4367 (N_4367,In_176,In_672);
nor U4368 (N_4368,In_1954,In_1468);
or U4369 (N_4369,In_3601,In_2477);
xnor U4370 (N_4370,In_2725,In_121);
and U4371 (N_4371,In_4756,In_2241);
or U4372 (N_4372,In_2491,In_1812);
or U4373 (N_4373,In_888,In_4447);
or U4374 (N_4374,In_1541,In_4046);
nor U4375 (N_4375,In_4506,In_242);
nor U4376 (N_4376,In_2403,In_339);
nor U4377 (N_4377,In_2419,In_623);
xnor U4378 (N_4378,In_2335,In_671);
xor U4379 (N_4379,In_1839,In_1276);
nand U4380 (N_4380,In_1012,In_4716);
or U4381 (N_4381,In_2633,In_2543);
nor U4382 (N_4382,In_4520,In_4880);
nor U4383 (N_4383,In_4595,In_470);
nand U4384 (N_4384,In_1179,In_572);
and U4385 (N_4385,In_3088,In_556);
or U4386 (N_4386,In_3556,In_3283);
xnor U4387 (N_4387,In_4681,In_1441);
xnor U4388 (N_4388,In_2803,In_85);
nor U4389 (N_4389,In_13,In_1501);
or U4390 (N_4390,In_2435,In_4809);
nor U4391 (N_4391,In_1482,In_2306);
and U4392 (N_4392,In_3330,In_3448);
nor U4393 (N_4393,In_4845,In_276);
xnor U4394 (N_4394,In_1318,In_1196);
nor U4395 (N_4395,In_4836,In_3518);
nand U4396 (N_4396,In_436,In_2976);
and U4397 (N_4397,In_4381,In_3673);
nor U4398 (N_4398,In_945,In_4352);
xor U4399 (N_4399,In_1392,In_4260);
nand U4400 (N_4400,In_4053,In_1643);
or U4401 (N_4401,In_3397,In_299);
and U4402 (N_4402,In_2557,In_3963);
xor U4403 (N_4403,In_4081,In_1993);
nor U4404 (N_4404,In_1629,In_4730);
nand U4405 (N_4405,In_648,In_2847);
nor U4406 (N_4406,In_622,In_2256);
nor U4407 (N_4407,In_1960,In_4753);
xnor U4408 (N_4408,In_1355,In_2670);
nand U4409 (N_4409,In_3059,In_2244);
or U4410 (N_4410,In_1019,In_2452);
or U4411 (N_4411,In_1996,In_3686);
or U4412 (N_4412,In_322,In_2135);
nor U4413 (N_4413,In_1495,In_2113);
nor U4414 (N_4414,In_65,In_2684);
xnor U4415 (N_4415,In_1718,In_3004);
nor U4416 (N_4416,In_2574,In_1545);
and U4417 (N_4417,In_1414,In_2672);
xor U4418 (N_4418,In_1436,In_2235);
nand U4419 (N_4419,In_741,In_1878);
nand U4420 (N_4420,In_363,In_711);
or U4421 (N_4421,In_299,In_3064);
nor U4422 (N_4422,In_4911,In_574);
xor U4423 (N_4423,In_1287,In_444);
nor U4424 (N_4424,In_2689,In_3461);
nand U4425 (N_4425,In_1388,In_2665);
xnor U4426 (N_4426,In_1087,In_3577);
nand U4427 (N_4427,In_3891,In_1638);
xnor U4428 (N_4428,In_1772,In_1822);
nor U4429 (N_4429,In_276,In_4993);
xnor U4430 (N_4430,In_4144,In_300);
and U4431 (N_4431,In_3268,In_4896);
and U4432 (N_4432,In_4333,In_2815);
or U4433 (N_4433,In_2718,In_4088);
or U4434 (N_4434,In_1672,In_2019);
xor U4435 (N_4435,In_4389,In_311);
and U4436 (N_4436,In_3257,In_406);
nor U4437 (N_4437,In_903,In_3366);
or U4438 (N_4438,In_3770,In_3761);
and U4439 (N_4439,In_1552,In_927);
xor U4440 (N_4440,In_4788,In_604);
nand U4441 (N_4441,In_4327,In_3231);
and U4442 (N_4442,In_2950,In_3013);
nor U4443 (N_4443,In_4910,In_3547);
nor U4444 (N_4444,In_146,In_3897);
nor U4445 (N_4445,In_883,In_2296);
nor U4446 (N_4446,In_1951,In_3536);
nor U4447 (N_4447,In_193,In_2766);
and U4448 (N_4448,In_540,In_363);
or U4449 (N_4449,In_4931,In_2071);
or U4450 (N_4450,In_3440,In_719);
and U4451 (N_4451,In_4307,In_717);
xnor U4452 (N_4452,In_812,In_4376);
nor U4453 (N_4453,In_2836,In_4884);
or U4454 (N_4454,In_2951,In_191);
xnor U4455 (N_4455,In_4688,In_2294);
nand U4456 (N_4456,In_3281,In_1);
and U4457 (N_4457,In_212,In_369);
and U4458 (N_4458,In_780,In_3844);
and U4459 (N_4459,In_750,In_877);
nor U4460 (N_4460,In_4309,In_975);
and U4461 (N_4461,In_1663,In_2784);
or U4462 (N_4462,In_554,In_4463);
or U4463 (N_4463,In_846,In_241);
or U4464 (N_4464,In_3912,In_1113);
or U4465 (N_4465,In_416,In_4370);
and U4466 (N_4466,In_422,In_2243);
or U4467 (N_4467,In_267,In_606);
and U4468 (N_4468,In_1491,In_2210);
or U4469 (N_4469,In_4383,In_1500);
xnor U4470 (N_4470,In_4218,In_1753);
nand U4471 (N_4471,In_4374,In_2235);
nor U4472 (N_4472,In_1321,In_3067);
xor U4473 (N_4473,In_850,In_420);
xor U4474 (N_4474,In_2999,In_4803);
and U4475 (N_4475,In_2503,In_4394);
and U4476 (N_4476,In_360,In_1992);
xnor U4477 (N_4477,In_1008,In_1881);
nor U4478 (N_4478,In_2803,In_4609);
nand U4479 (N_4479,In_2939,In_3788);
or U4480 (N_4480,In_2682,In_1790);
nand U4481 (N_4481,In_4617,In_1834);
nor U4482 (N_4482,In_498,In_4454);
and U4483 (N_4483,In_3626,In_1131);
and U4484 (N_4484,In_830,In_1441);
xnor U4485 (N_4485,In_362,In_4233);
nand U4486 (N_4486,In_2818,In_3820);
nand U4487 (N_4487,In_1196,In_1919);
or U4488 (N_4488,In_2356,In_301);
nor U4489 (N_4489,In_4590,In_3473);
or U4490 (N_4490,In_1624,In_3046);
or U4491 (N_4491,In_2078,In_2427);
xnor U4492 (N_4492,In_4874,In_4347);
xnor U4493 (N_4493,In_851,In_1847);
nand U4494 (N_4494,In_4018,In_3562);
and U4495 (N_4495,In_1079,In_1505);
xnor U4496 (N_4496,In_2542,In_2546);
and U4497 (N_4497,In_939,In_923);
nor U4498 (N_4498,In_3230,In_7);
xor U4499 (N_4499,In_2590,In_605);
xor U4500 (N_4500,In_296,In_4288);
nor U4501 (N_4501,In_999,In_3451);
nor U4502 (N_4502,In_4856,In_2933);
nand U4503 (N_4503,In_319,In_2332);
or U4504 (N_4504,In_2553,In_2347);
nor U4505 (N_4505,In_2064,In_94);
nand U4506 (N_4506,In_1741,In_4154);
nand U4507 (N_4507,In_379,In_2183);
nand U4508 (N_4508,In_687,In_27);
or U4509 (N_4509,In_1253,In_2380);
and U4510 (N_4510,In_4715,In_3164);
nor U4511 (N_4511,In_1518,In_2563);
and U4512 (N_4512,In_970,In_4060);
or U4513 (N_4513,In_4967,In_857);
xnor U4514 (N_4514,In_3843,In_3749);
xor U4515 (N_4515,In_4287,In_2426);
or U4516 (N_4516,In_2273,In_3066);
xor U4517 (N_4517,In_2148,In_3429);
and U4518 (N_4518,In_2063,In_688);
and U4519 (N_4519,In_3585,In_3947);
or U4520 (N_4520,In_3025,In_2239);
xnor U4521 (N_4521,In_560,In_860);
xor U4522 (N_4522,In_2073,In_1054);
or U4523 (N_4523,In_495,In_2937);
nand U4524 (N_4524,In_366,In_220);
or U4525 (N_4525,In_522,In_2752);
nor U4526 (N_4526,In_2022,In_1470);
xnor U4527 (N_4527,In_1641,In_4246);
xor U4528 (N_4528,In_1680,In_286);
and U4529 (N_4529,In_4735,In_3701);
xnor U4530 (N_4530,In_4620,In_1605);
nor U4531 (N_4531,In_1843,In_1497);
or U4532 (N_4532,In_2162,In_2068);
xnor U4533 (N_4533,In_3955,In_2667);
or U4534 (N_4534,In_1908,In_2163);
xor U4535 (N_4535,In_3555,In_4095);
xnor U4536 (N_4536,In_2026,In_4757);
nand U4537 (N_4537,In_3016,In_2872);
nand U4538 (N_4538,In_1867,In_125);
xor U4539 (N_4539,In_4644,In_236);
or U4540 (N_4540,In_4441,In_1322);
and U4541 (N_4541,In_3256,In_1253);
or U4542 (N_4542,In_3096,In_1667);
nor U4543 (N_4543,In_4725,In_3491);
xnor U4544 (N_4544,In_2657,In_1972);
nand U4545 (N_4545,In_4082,In_1176);
nand U4546 (N_4546,In_4170,In_2738);
nand U4547 (N_4547,In_1633,In_2504);
or U4548 (N_4548,In_2989,In_2524);
and U4549 (N_4549,In_2884,In_3337);
and U4550 (N_4550,In_713,In_4673);
or U4551 (N_4551,In_4037,In_1837);
and U4552 (N_4552,In_3333,In_4309);
or U4553 (N_4553,In_2907,In_1849);
and U4554 (N_4554,In_1670,In_4052);
xnor U4555 (N_4555,In_2105,In_217);
and U4556 (N_4556,In_2332,In_3422);
nand U4557 (N_4557,In_3526,In_978);
and U4558 (N_4558,In_4259,In_3892);
nand U4559 (N_4559,In_1517,In_4425);
or U4560 (N_4560,In_919,In_4501);
xor U4561 (N_4561,In_3940,In_3058);
and U4562 (N_4562,In_3525,In_1560);
nor U4563 (N_4563,In_4165,In_151);
or U4564 (N_4564,In_48,In_1609);
nor U4565 (N_4565,In_1518,In_3698);
or U4566 (N_4566,In_384,In_3569);
xor U4567 (N_4567,In_2610,In_4331);
and U4568 (N_4568,In_2865,In_4046);
and U4569 (N_4569,In_2411,In_4850);
nor U4570 (N_4570,In_3146,In_2123);
or U4571 (N_4571,In_2588,In_3923);
and U4572 (N_4572,In_3058,In_3000);
or U4573 (N_4573,In_249,In_2294);
and U4574 (N_4574,In_2398,In_4145);
xnor U4575 (N_4575,In_4107,In_3182);
or U4576 (N_4576,In_1260,In_1691);
nand U4577 (N_4577,In_4470,In_4355);
and U4578 (N_4578,In_3434,In_202);
and U4579 (N_4579,In_4772,In_6);
and U4580 (N_4580,In_4077,In_294);
and U4581 (N_4581,In_4864,In_1374);
nor U4582 (N_4582,In_3668,In_4423);
nand U4583 (N_4583,In_1334,In_4760);
xnor U4584 (N_4584,In_688,In_2133);
and U4585 (N_4585,In_4869,In_753);
or U4586 (N_4586,In_1939,In_2894);
nand U4587 (N_4587,In_2300,In_17);
xnor U4588 (N_4588,In_2700,In_470);
nand U4589 (N_4589,In_2081,In_935);
xor U4590 (N_4590,In_3062,In_1349);
nand U4591 (N_4591,In_1891,In_4721);
xnor U4592 (N_4592,In_1843,In_1005);
or U4593 (N_4593,In_4999,In_4282);
xor U4594 (N_4594,In_2382,In_2792);
nand U4595 (N_4595,In_3663,In_4659);
and U4596 (N_4596,In_3531,In_4764);
nand U4597 (N_4597,In_4811,In_3793);
nand U4598 (N_4598,In_421,In_2453);
xor U4599 (N_4599,In_4555,In_1116);
xnor U4600 (N_4600,In_2463,In_1321);
or U4601 (N_4601,In_3941,In_1956);
and U4602 (N_4602,In_80,In_4325);
xnor U4603 (N_4603,In_2518,In_2937);
nand U4604 (N_4604,In_4705,In_289);
or U4605 (N_4605,In_3555,In_1389);
or U4606 (N_4606,In_153,In_4291);
nor U4607 (N_4607,In_4973,In_4350);
or U4608 (N_4608,In_3579,In_1105);
nor U4609 (N_4609,In_2843,In_4308);
or U4610 (N_4610,In_4638,In_3860);
nor U4611 (N_4611,In_2076,In_2241);
or U4612 (N_4612,In_3530,In_4798);
xor U4613 (N_4613,In_3183,In_2800);
and U4614 (N_4614,In_305,In_4591);
nand U4615 (N_4615,In_4533,In_1071);
xnor U4616 (N_4616,In_4292,In_4235);
or U4617 (N_4617,In_2307,In_2534);
or U4618 (N_4618,In_3923,In_183);
nor U4619 (N_4619,In_4032,In_4899);
xor U4620 (N_4620,In_4750,In_537);
xor U4621 (N_4621,In_3276,In_3839);
or U4622 (N_4622,In_4116,In_4982);
or U4623 (N_4623,In_3703,In_1904);
nand U4624 (N_4624,In_752,In_1829);
nand U4625 (N_4625,In_3060,In_4977);
and U4626 (N_4626,In_101,In_1776);
xnor U4627 (N_4627,In_3781,In_4530);
nor U4628 (N_4628,In_1446,In_1886);
or U4629 (N_4629,In_1653,In_1766);
xor U4630 (N_4630,In_3714,In_4471);
xnor U4631 (N_4631,In_1578,In_1938);
or U4632 (N_4632,In_1700,In_4872);
and U4633 (N_4633,In_3441,In_180);
xor U4634 (N_4634,In_4350,In_1909);
nor U4635 (N_4635,In_3872,In_3752);
and U4636 (N_4636,In_3035,In_2487);
or U4637 (N_4637,In_516,In_2957);
nor U4638 (N_4638,In_62,In_4237);
xnor U4639 (N_4639,In_2901,In_1873);
nand U4640 (N_4640,In_202,In_436);
or U4641 (N_4641,In_3188,In_212);
nor U4642 (N_4642,In_2402,In_582);
nand U4643 (N_4643,In_3985,In_1909);
nand U4644 (N_4644,In_123,In_2320);
nand U4645 (N_4645,In_1063,In_4927);
or U4646 (N_4646,In_1121,In_4989);
nor U4647 (N_4647,In_3726,In_3472);
or U4648 (N_4648,In_1430,In_2945);
and U4649 (N_4649,In_2359,In_3113);
and U4650 (N_4650,In_4754,In_3896);
nand U4651 (N_4651,In_2082,In_688);
nand U4652 (N_4652,In_2820,In_1870);
and U4653 (N_4653,In_4059,In_4029);
or U4654 (N_4654,In_96,In_1343);
nand U4655 (N_4655,In_4436,In_4552);
xnor U4656 (N_4656,In_4761,In_2251);
and U4657 (N_4657,In_3931,In_4777);
nor U4658 (N_4658,In_2017,In_4955);
nand U4659 (N_4659,In_4095,In_2732);
and U4660 (N_4660,In_457,In_1595);
and U4661 (N_4661,In_1446,In_1825);
or U4662 (N_4662,In_1170,In_4340);
xnor U4663 (N_4663,In_2622,In_4172);
nor U4664 (N_4664,In_3498,In_3485);
nand U4665 (N_4665,In_4492,In_4477);
xnor U4666 (N_4666,In_3415,In_782);
nand U4667 (N_4667,In_1199,In_1749);
nand U4668 (N_4668,In_4497,In_1679);
and U4669 (N_4669,In_1050,In_1222);
or U4670 (N_4670,In_188,In_609);
or U4671 (N_4671,In_2380,In_4031);
nor U4672 (N_4672,In_4568,In_3702);
nor U4673 (N_4673,In_3153,In_4704);
nand U4674 (N_4674,In_2339,In_369);
or U4675 (N_4675,In_2455,In_1);
nor U4676 (N_4676,In_1413,In_883);
or U4677 (N_4677,In_497,In_951);
xnor U4678 (N_4678,In_2761,In_2843);
nand U4679 (N_4679,In_1180,In_697);
nand U4680 (N_4680,In_18,In_3997);
xor U4681 (N_4681,In_2925,In_3576);
nor U4682 (N_4682,In_3136,In_277);
nor U4683 (N_4683,In_4678,In_1709);
nand U4684 (N_4684,In_1372,In_2342);
nor U4685 (N_4685,In_676,In_3395);
nor U4686 (N_4686,In_4604,In_4964);
xnor U4687 (N_4687,In_2363,In_2747);
or U4688 (N_4688,In_2239,In_4550);
or U4689 (N_4689,In_4012,In_4810);
and U4690 (N_4690,In_598,In_3559);
or U4691 (N_4691,In_940,In_2602);
xnor U4692 (N_4692,In_4883,In_4689);
and U4693 (N_4693,In_3362,In_4868);
or U4694 (N_4694,In_631,In_2834);
and U4695 (N_4695,In_1581,In_3855);
nand U4696 (N_4696,In_4486,In_2164);
or U4697 (N_4697,In_4525,In_302);
nor U4698 (N_4698,In_578,In_1644);
xor U4699 (N_4699,In_1966,In_4691);
xor U4700 (N_4700,In_4997,In_304);
nand U4701 (N_4701,In_1755,In_871);
xnor U4702 (N_4702,In_4698,In_4887);
nor U4703 (N_4703,In_2925,In_2432);
xor U4704 (N_4704,In_1781,In_2651);
or U4705 (N_4705,In_4986,In_2781);
and U4706 (N_4706,In_4286,In_1796);
and U4707 (N_4707,In_1066,In_1311);
and U4708 (N_4708,In_4977,In_4920);
xnor U4709 (N_4709,In_2281,In_1731);
nand U4710 (N_4710,In_2858,In_156);
nor U4711 (N_4711,In_3869,In_2996);
nor U4712 (N_4712,In_3315,In_3754);
nand U4713 (N_4713,In_3253,In_1342);
and U4714 (N_4714,In_4197,In_1619);
xor U4715 (N_4715,In_133,In_4811);
or U4716 (N_4716,In_1780,In_4557);
and U4717 (N_4717,In_1577,In_4991);
nor U4718 (N_4718,In_3739,In_1977);
nand U4719 (N_4719,In_4826,In_2712);
nor U4720 (N_4720,In_4766,In_36);
and U4721 (N_4721,In_21,In_2814);
nor U4722 (N_4722,In_4663,In_3307);
nor U4723 (N_4723,In_3566,In_4750);
xnor U4724 (N_4724,In_4226,In_1710);
nor U4725 (N_4725,In_1223,In_85);
or U4726 (N_4726,In_2260,In_1855);
nand U4727 (N_4727,In_175,In_4565);
or U4728 (N_4728,In_4140,In_230);
nand U4729 (N_4729,In_1211,In_3864);
xor U4730 (N_4730,In_4469,In_4677);
or U4731 (N_4731,In_3292,In_2074);
and U4732 (N_4732,In_3185,In_4058);
or U4733 (N_4733,In_1074,In_2813);
xor U4734 (N_4734,In_1443,In_3069);
nor U4735 (N_4735,In_618,In_1427);
or U4736 (N_4736,In_4990,In_4311);
xnor U4737 (N_4737,In_2749,In_3056);
xnor U4738 (N_4738,In_1870,In_4757);
nor U4739 (N_4739,In_1828,In_4802);
and U4740 (N_4740,In_3516,In_385);
xor U4741 (N_4741,In_4782,In_2735);
and U4742 (N_4742,In_1169,In_3839);
nand U4743 (N_4743,In_4776,In_1807);
or U4744 (N_4744,In_4309,In_2922);
nand U4745 (N_4745,In_1773,In_2951);
nor U4746 (N_4746,In_1334,In_2874);
xor U4747 (N_4747,In_1767,In_4638);
nand U4748 (N_4748,In_1038,In_1356);
or U4749 (N_4749,In_4611,In_2739);
or U4750 (N_4750,In_1493,In_3108);
nor U4751 (N_4751,In_3318,In_378);
xor U4752 (N_4752,In_4419,In_2116);
nand U4753 (N_4753,In_0,In_3058);
nor U4754 (N_4754,In_3653,In_1816);
nand U4755 (N_4755,In_824,In_4009);
and U4756 (N_4756,In_1024,In_4924);
nor U4757 (N_4757,In_553,In_2490);
nand U4758 (N_4758,In_2277,In_2393);
and U4759 (N_4759,In_3931,In_3859);
and U4760 (N_4760,In_4509,In_110);
and U4761 (N_4761,In_769,In_4966);
nand U4762 (N_4762,In_2863,In_4435);
and U4763 (N_4763,In_1136,In_4871);
xnor U4764 (N_4764,In_4899,In_3330);
nor U4765 (N_4765,In_3550,In_4049);
xor U4766 (N_4766,In_4260,In_2025);
xor U4767 (N_4767,In_3929,In_2811);
nand U4768 (N_4768,In_1372,In_1607);
nand U4769 (N_4769,In_4950,In_1966);
or U4770 (N_4770,In_3426,In_3070);
nand U4771 (N_4771,In_2542,In_541);
and U4772 (N_4772,In_591,In_50);
nor U4773 (N_4773,In_4750,In_4695);
nand U4774 (N_4774,In_1529,In_1556);
nor U4775 (N_4775,In_1755,In_2338);
and U4776 (N_4776,In_4154,In_4153);
nor U4777 (N_4777,In_325,In_4444);
nor U4778 (N_4778,In_3666,In_2528);
xor U4779 (N_4779,In_1363,In_2405);
xor U4780 (N_4780,In_2619,In_315);
and U4781 (N_4781,In_608,In_4279);
nand U4782 (N_4782,In_3086,In_2101);
and U4783 (N_4783,In_3919,In_985);
and U4784 (N_4784,In_1815,In_3833);
and U4785 (N_4785,In_2315,In_4324);
nand U4786 (N_4786,In_2769,In_840);
nor U4787 (N_4787,In_2290,In_1370);
nand U4788 (N_4788,In_4246,In_4939);
or U4789 (N_4789,In_4827,In_3026);
nor U4790 (N_4790,In_1683,In_4904);
nand U4791 (N_4791,In_483,In_139);
nor U4792 (N_4792,In_488,In_2394);
and U4793 (N_4793,In_3284,In_679);
nor U4794 (N_4794,In_2984,In_225);
or U4795 (N_4795,In_3309,In_2942);
and U4796 (N_4796,In_4973,In_1761);
nand U4797 (N_4797,In_4862,In_4143);
xor U4798 (N_4798,In_1627,In_4069);
and U4799 (N_4799,In_1259,In_3284);
nand U4800 (N_4800,In_1273,In_4402);
and U4801 (N_4801,In_4434,In_2130);
xor U4802 (N_4802,In_1173,In_574);
or U4803 (N_4803,In_4399,In_3855);
xor U4804 (N_4804,In_1746,In_1448);
and U4805 (N_4805,In_2852,In_4612);
nor U4806 (N_4806,In_4450,In_3685);
nand U4807 (N_4807,In_1058,In_3219);
xor U4808 (N_4808,In_3037,In_4126);
nand U4809 (N_4809,In_4451,In_2294);
nand U4810 (N_4810,In_1661,In_2776);
nor U4811 (N_4811,In_1059,In_621);
or U4812 (N_4812,In_598,In_2205);
nor U4813 (N_4813,In_159,In_3699);
nand U4814 (N_4814,In_559,In_3056);
xnor U4815 (N_4815,In_3005,In_2747);
xnor U4816 (N_4816,In_4745,In_3810);
xor U4817 (N_4817,In_2342,In_4645);
and U4818 (N_4818,In_1761,In_2343);
nor U4819 (N_4819,In_1452,In_143);
or U4820 (N_4820,In_4728,In_3005);
xnor U4821 (N_4821,In_1581,In_468);
nor U4822 (N_4822,In_3469,In_4528);
xnor U4823 (N_4823,In_2631,In_3179);
or U4824 (N_4824,In_4937,In_1483);
nand U4825 (N_4825,In_3412,In_4320);
xnor U4826 (N_4826,In_573,In_4208);
nand U4827 (N_4827,In_655,In_3856);
nand U4828 (N_4828,In_3017,In_4559);
and U4829 (N_4829,In_3356,In_3900);
xnor U4830 (N_4830,In_3239,In_467);
nor U4831 (N_4831,In_3332,In_2925);
or U4832 (N_4832,In_158,In_1126);
nor U4833 (N_4833,In_4805,In_2402);
nor U4834 (N_4834,In_4463,In_1765);
nand U4835 (N_4835,In_4794,In_1905);
and U4836 (N_4836,In_2125,In_1425);
nor U4837 (N_4837,In_4736,In_4633);
nand U4838 (N_4838,In_2703,In_3272);
xor U4839 (N_4839,In_4259,In_306);
and U4840 (N_4840,In_3053,In_4110);
and U4841 (N_4841,In_2864,In_2201);
or U4842 (N_4842,In_3982,In_4009);
and U4843 (N_4843,In_852,In_2743);
xnor U4844 (N_4844,In_689,In_2517);
nand U4845 (N_4845,In_2248,In_1751);
nor U4846 (N_4846,In_360,In_138);
or U4847 (N_4847,In_807,In_112);
nand U4848 (N_4848,In_981,In_2333);
or U4849 (N_4849,In_1129,In_2895);
and U4850 (N_4850,In_4520,In_669);
xnor U4851 (N_4851,In_4427,In_3903);
and U4852 (N_4852,In_4386,In_1760);
or U4853 (N_4853,In_3752,In_2165);
xor U4854 (N_4854,In_4503,In_2747);
and U4855 (N_4855,In_4085,In_1918);
xor U4856 (N_4856,In_1656,In_1654);
nand U4857 (N_4857,In_195,In_903);
and U4858 (N_4858,In_3838,In_4635);
nand U4859 (N_4859,In_4053,In_1243);
or U4860 (N_4860,In_2792,In_2089);
and U4861 (N_4861,In_3342,In_4095);
xor U4862 (N_4862,In_2081,In_1230);
nor U4863 (N_4863,In_4215,In_4863);
and U4864 (N_4864,In_866,In_4275);
nand U4865 (N_4865,In_2353,In_3838);
xnor U4866 (N_4866,In_3772,In_4927);
or U4867 (N_4867,In_209,In_3004);
nor U4868 (N_4868,In_4745,In_2807);
xnor U4869 (N_4869,In_989,In_1939);
or U4870 (N_4870,In_2967,In_664);
nor U4871 (N_4871,In_2384,In_1248);
and U4872 (N_4872,In_233,In_1029);
xor U4873 (N_4873,In_2370,In_2274);
nor U4874 (N_4874,In_3971,In_0);
nor U4875 (N_4875,In_1494,In_1190);
nor U4876 (N_4876,In_2863,In_931);
or U4877 (N_4877,In_1097,In_2283);
or U4878 (N_4878,In_1764,In_3579);
or U4879 (N_4879,In_3860,In_3303);
nand U4880 (N_4880,In_2720,In_2017);
nand U4881 (N_4881,In_3586,In_2449);
and U4882 (N_4882,In_140,In_374);
nand U4883 (N_4883,In_2989,In_2149);
nand U4884 (N_4884,In_4488,In_1707);
and U4885 (N_4885,In_4976,In_587);
or U4886 (N_4886,In_1428,In_1451);
nand U4887 (N_4887,In_751,In_821);
xnor U4888 (N_4888,In_2948,In_2088);
nand U4889 (N_4889,In_4077,In_2701);
nor U4890 (N_4890,In_4524,In_4447);
nand U4891 (N_4891,In_1711,In_1013);
nand U4892 (N_4892,In_2606,In_807);
nand U4893 (N_4893,In_1005,In_2457);
nand U4894 (N_4894,In_4283,In_2330);
and U4895 (N_4895,In_4396,In_255);
and U4896 (N_4896,In_2129,In_258);
or U4897 (N_4897,In_3692,In_375);
xnor U4898 (N_4898,In_4515,In_81);
or U4899 (N_4899,In_1768,In_2269);
nand U4900 (N_4900,In_4435,In_3735);
nor U4901 (N_4901,In_1531,In_1463);
and U4902 (N_4902,In_3470,In_2664);
or U4903 (N_4903,In_305,In_958);
nand U4904 (N_4904,In_3704,In_1060);
or U4905 (N_4905,In_1745,In_912);
or U4906 (N_4906,In_2076,In_1253);
or U4907 (N_4907,In_3865,In_4506);
nor U4908 (N_4908,In_4953,In_4949);
nand U4909 (N_4909,In_4642,In_121);
or U4910 (N_4910,In_1267,In_676);
or U4911 (N_4911,In_1012,In_3917);
and U4912 (N_4912,In_3911,In_2967);
xnor U4913 (N_4913,In_2522,In_4228);
nor U4914 (N_4914,In_2983,In_2970);
xnor U4915 (N_4915,In_4003,In_1080);
nor U4916 (N_4916,In_990,In_3354);
nand U4917 (N_4917,In_2079,In_2694);
or U4918 (N_4918,In_1916,In_226);
and U4919 (N_4919,In_3748,In_2914);
xnor U4920 (N_4920,In_4656,In_3339);
nor U4921 (N_4921,In_3480,In_3069);
and U4922 (N_4922,In_1921,In_953);
and U4923 (N_4923,In_1151,In_3471);
xor U4924 (N_4924,In_833,In_4900);
nor U4925 (N_4925,In_2376,In_4534);
nor U4926 (N_4926,In_2296,In_2791);
or U4927 (N_4927,In_3381,In_1712);
and U4928 (N_4928,In_2559,In_2985);
nand U4929 (N_4929,In_4232,In_4525);
and U4930 (N_4930,In_1322,In_3945);
xnor U4931 (N_4931,In_3499,In_4661);
xnor U4932 (N_4932,In_4801,In_3067);
nand U4933 (N_4933,In_3403,In_4240);
or U4934 (N_4934,In_2217,In_1198);
xor U4935 (N_4935,In_4815,In_3883);
and U4936 (N_4936,In_1927,In_704);
nor U4937 (N_4937,In_1185,In_4808);
nand U4938 (N_4938,In_4540,In_1459);
nor U4939 (N_4939,In_1221,In_2088);
and U4940 (N_4940,In_1491,In_904);
and U4941 (N_4941,In_407,In_2534);
or U4942 (N_4942,In_1051,In_25);
and U4943 (N_4943,In_3876,In_1096);
xnor U4944 (N_4944,In_1916,In_2998);
and U4945 (N_4945,In_459,In_3354);
xor U4946 (N_4946,In_3358,In_2669);
nand U4947 (N_4947,In_781,In_2316);
and U4948 (N_4948,In_2563,In_3128);
and U4949 (N_4949,In_3679,In_3048);
nand U4950 (N_4950,In_3684,In_4102);
nand U4951 (N_4951,In_427,In_4307);
nor U4952 (N_4952,In_3555,In_1524);
or U4953 (N_4953,In_526,In_4614);
or U4954 (N_4954,In_3921,In_3919);
or U4955 (N_4955,In_1346,In_2858);
and U4956 (N_4956,In_2281,In_1257);
xnor U4957 (N_4957,In_4258,In_3500);
or U4958 (N_4958,In_4248,In_4681);
and U4959 (N_4959,In_830,In_3554);
nor U4960 (N_4960,In_615,In_805);
nand U4961 (N_4961,In_2399,In_3446);
and U4962 (N_4962,In_4650,In_1989);
nor U4963 (N_4963,In_2603,In_1574);
nor U4964 (N_4964,In_4069,In_3969);
and U4965 (N_4965,In_2762,In_2889);
and U4966 (N_4966,In_104,In_263);
xor U4967 (N_4967,In_100,In_3058);
xnor U4968 (N_4968,In_617,In_3274);
nor U4969 (N_4969,In_1491,In_2325);
nor U4970 (N_4970,In_4559,In_2918);
xor U4971 (N_4971,In_997,In_2401);
xor U4972 (N_4972,In_1953,In_3950);
and U4973 (N_4973,In_4888,In_2064);
nand U4974 (N_4974,In_1169,In_2531);
nor U4975 (N_4975,In_4004,In_419);
nand U4976 (N_4976,In_3662,In_4018);
or U4977 (N_4977,In_419,In_3270);
and U4978 (N_4978,In_4015,In_4856);
nor U4979 (N_4979,In_3355,In_3559);
or U4980 (N_4980,In_3657,In_3738);
xor U4981 (N_4981,In_820,In_2354);
nor U4982 (N_4982,In_1741,In_2037);
xor U4983 (N_4983,In_4814,In_2565);
and U4984 (N_4984,In_4653,In_1216);
or U4985 (N_4985,In_1860,In_4597);
nand U4986 (N_4986,In_1691,In_3300);
xor U4987 (N_4987,In_4782,In_2212);
nand U4988 (N_4988,In_1400,In_2126);
and U4989 (N_4989,In_1790,In_2913);
and U4990 (N_4990,In_2469,In_3508);
xnor U4991 (N_4991,In_343,In_3455);
nor U4992 (N_4992,In_2576,In_950);
nand U4993 (N_4993,In_1114,In_1062);
xor U4994 (N_4994,In_1260,In_2284);
or U4995 (N_4995,In_1362,In_862);
and U4996 (N_4996,In_4311,In_2995);
or U4997 (N_4997,In_1124,In_3310);
and U4998 (N_4998,In_1374,In_1077);
and U4999 (N_4999,In_3966,In_624);
nor U5000 (N_5000,N_4128,N_928);
or U5001 (N_5001,N_4789,N_2770);
or U5002 (N_5002,N_1015,N_1801);
xnor U5003 (N_5003,N_3397,N_4020);
nand U5004 (N_5004,N_761,N_4536);
or U5005 (N_5005,N_4451,N_4774);
xnor U5006 (N_5006,N_2602,N_289);
nand U5007 (N_5007,N_631,N_867);
or U5008 (N_5008,N_4659,N_489);
and U5009 (N_5009,N_4094,N_3120);
nor U5010 (N_5010,N_4405,N_1521);
and U5011 (N_5011,N_4655,N_2195);
nand U5012 (N_5012,N_2817,N_2329);
nor U5013 (N_5013,N_4191,N_3053);
and U5014 (N_5014,N_4423,N_2284);
and U5015 (N_5015,N_3785,N_1459);
nor U5016 (N_5016,N_1298,N_2234);
nor U5017 (N_5017,N_4845,N_3270);
and U5018 (N_5018,N_3230,N_2975);
nand U5019 (N_5019,N_4573,N_4647);
xor U5020 (N_5020,N_1297,N_4061);
nand U5021 (N_5021,N_1181,N_104);
nand U5022 (N_5022,N_1689,N_4348);
nor U5023 (N_5023,N_4673,N_1940);
nor U5024 (N_5024,N_2398,N_1619);
nor U5025 (N_5025,N_4228,N_2368);
xnor U5026 (N_5026,N_3472,N_1887);
and U5027 (N_5027,N_849,N_2695);
or U5028 (N_5028,N_973,N_471);
or U5029 (N_5029,N_2105,N_2137);
and U5030 (N_5030,N_4723,N_703);
nor U5031 (N_5031,N_3014,N_4392);
and U5032 (N_5032,N_4415,N_3551);
nand U5033 (N_5033,N_2045,N_2459);
or U5034 (N_5034,N_4565,N_4034);
or U5035 (N_5035,N_2856,N_3231);
nor U5036 (N_5036,N_2675,N_921);
xnor U5037 (N_5037,N_4317,N_1236);
xor U5038 (N_5038,N_4920,N_3870);
nand U5039 (N_5039,N_589,N_4242);
or U5040 (N_5040,N_2692,N_3089);
nor U5041 (N_5041,N_157,N_4626);
nor U5042 (N_5042,N_887,N_3914);
nand U5043 (N_5043,N_2120,N_4289);
or U5044 (N_5044,N_2269,N_2507);
and U5045 (N_5045,N_1379,N_252);
or U5046 (N_5046,N_3070,N_4460);
xor U5047 (N_5047,N_4106,N_3916);
nand U5048 (N_5048,N_2025,N_894);
or U5049 (N_5049,N_3498,N_4780);
nor U5050 (N_5050,N_698,N_1874);
nand U5051 (N_5051,N_430,N_109);
nor U5052 (N_5052,N_4428,N_4422);
and U5053 (N_5053,N_1764,N_689);
xor U5054 (N_5054,N_2651,N_1515);
nor U5055 (N_5055,N_4874,N_1660);
or U5056 (N_5056,N_2781,N_3692);
and U5057 (N_5057,N_400,N_1734);
or U5058 (N_5058,N_1749,N_1659);
xnor U5059 (N_5059,N_1322,N_2630);
nor U5060 (N_5060,N_3359,N_3437);
or U5061 (N_5061,N_1520,N_13);
nand U5062 (N_5062,N_4346,N_1434);
nand U5063 (N_5063,N_4892,N_1216);
nor U5064 (N_5064,N_251,N_2057);
or U5065 (N_5065,N_4986,N_4374);
or U5066 (N_5066,N_614,N_3325);
or U5067 (N_5067,N_4999,N_48);
nor U5068 (N_5068,N_263,N_2967);
nor U5069 (N_5069,N_4375,N_2657);
xnor U5070 (N_5070,N_2422,N_904);
nor U5071 (N_5071,N_1074,N_3180);
nand U5072 (N_5072,N_4746,N_1321);
nor U5073 (N_5073,N_3453,N_2176);
xor U5074 (N_5074,N_4104,N_3224);
xor U5075 (N_5075,N_3521,N_2166);
and U5076 (N_5076,N_1138,N_356);
nor U5077 (N_5077,N_4599,N_490);
nand U5078 (N_5078,N_1964,N_3335);
nand U5079 (N_5079,N_84,N_1990);
nor U5080 (N_5080,N_4617,N_2155);
and U5081 (N_5081,N_2158,N_4881);
xor U5082 (N_5082,N_4581,N_999);
and U5083 (N_5083,N_3966,N_818);
and U5084 (N_5084,N_1227,N_3164);
nand U5085 (N_5085,N_2172,N_3924);
nor U5086 (N_5086,N_685,N_4880);
or U5087 (N_5087,N_4725,N_4591);
and U5088 (N_5088,N_4563,N_154);
or U5089 (N_5089,N_143,N_1451);
or U5090 (N_5090,N_971,N_2421);
nand U5091 (N_5091,N_2959,N_2793);
or U5092 (N_5092,N_3479,N_3087);
nor U5093 (N_5093,N_4463,N_2382);
xor U5094 (N_5094,N_142,N_1192);
xnor U5095 (N_5095,N_1108,N_4509);
or U5096 (N_5096,N_2849,N_1654);
nand U5097 (N_5097,N_1334,N_4437);
and U5098 (N_5098,N_3592,N_3755);
nor U5099 (N_5099,N_60,N_2525);
nor U5100 (N_5100,N_2191,N_2788);
or U5101 (N_5101,N_2992,N_483);
nand U5102 (N_5102,N_1413,N_372);
and U5103 (N_5103,N_2659,N_1026);
nand U5104 (N_5104,N_2464,N_2117);
nand U5105 (N_5105,N_3513,N_3375);
xnor U5106 (N_5106,N_4871,N_3999);
and U5107 (N_5107,N_385,N_1507);
nor U5108 (N_5108,N_2409,N_2691);
or U5109 (N_5109,N_353,N_457);
nand U5110 (N_5110,N_923,N_375);
and U5111 (N_5111,N_3403,N_4692);
and U5112 (N_5112,N_3042,N_1273);
nand U5113 (N_5113,N_3394,N_4164);
xnor U5114 (N_5114,N_995,N_358);
nand U5115 (N_5115,N_4328,N_4544);
nand U5116 (N_5116,N_3439,N_1748);
nor U5117 (N_5117,N_2118,N_4301);
nand U5118 (N_5118,N_2873,N_2211);
nor U5119 (N_5119,N_1137,N_3222);
or U5120 (N_5120,N_3787,N_2365);
xor U5121 (N_5121,N_2955,N_61);
xor U5122 (N_5122,N_2109,N_3866);
nor U5123 (N_5123,N_3322,N_2958);
nor U5124 (N_5124,N_1633,N_1928);
xnor U5125 (N_5125,N_2946,N_2820);
nor U5126 (N_5126,N_4395,N_2361);
and U5127 (N_5127,N_113,N_4635);
and U5128 (N_5128,N_3185,N_4434);
nor U5129 (N_5129,N_795,N_1866);
nand U5130 (N_5130,N_1057,N_4997);
and U5131 (N_5131,N_3991,N_2640);
nand U5132 (N_5132,N_139,N_3243);
nor U5133 (N_5133,N_2373,N_3057);
nor U5134 (N_5134,N_1552,N_256);
nand U5135 (N_5135,N_1541,N_1881);
or U5136 (N_5136,N_3434,N_1981);
xnor U5137 (N_5137,N_1369,N_1551);
nand U5138 (N_5138,N_519,N_3934);
or U5139 (N_5139,N_269,N_344);
nor U5140 (N_5140,N_4934,N_331);
xor U5141 (N_5141,N_718,N_3738);
nand U5142 (N_5142,N_997,N_722);
xnor U5143 (N_5143,N_4837,N_440);
nand U5144 (N_5144,N_4925,N_4417);
and U5145 (N_5145,N_3074,N_3552);
nor U5146 (N_5146,N_4715,N_2564);
nor U5147 (N_5147,N_3500,N_4476);
xor U5148 (N_5148,N_525,N_3491);
nand U5149 (N_5149,N_441,N_858);
xnor U5150 (N_5150,N_3109,N_1182);
nor U5151 (N_5151,N_2775,N_2543);
or U5152 (N_5152,N_4987,N_3876);
xnor U5153 (N_5153,N_4053,N_1078);
nand U5154 (N_5154,N_1781,N_686);
or U5155 (N_5155,N_527,N_2981);
and U5156 (N_5156,N_2486,N_950);
nor U5157 (N_5157,N_2713,N_4564);
and U5158 (N_5158,N_3220,N_3277);
or U5159 (N_5159,N_4446,N_1729);
nand U5160 (N_5160,N_1937,N_3218);
xor U5161 (N_5161,N_1669,N_2064);
nand U5162 (N_5162,N_2749,N_4452);
and U5163 (N_5163,N_4649,N_955);
nor U5164 (N_5164,N_1152,N_526);
xor U5165 (N_5165,N_1492,N_337);
nor U5166 (N_5166,N_4033,N_1514);
nand U5167 (N_5167,N_4268,N_2816);
xor U5168 (N_5168,N_3568,N_1106);
and U5169 (N_5169,N_1315,N_1096);
nor U5170 (N_5170,N_1376,N_1031);
xor U5171 (N_5171,N_2810,N_173);
nand U5172 (N_5172,N_1891,N_4199);
xor U5173 (N_5173,N_357,N_1696);
nand U5174 (N_5174,N_55,N_4201);
xor U5175 (N_5175,N_4225,N_574);
nand U5176 (N_5176,N_3715,N_128);
or U5177 (N_5177,N_2047,N_4220);
nor U5178 (N_5178,N_339,N_2554);
and U5179 (N_5179,N_968,N_3878);
nand U5180 (N_5180,N_437,N_962);
nand U5181 (N_5181,N_3826,N_122);
and U5182 (N_5182,N_2467,N_102);
nand U5183 (N_5183,N_4802,N_4148);
nor U5184 (N_5184,N_1076,N_4279);
nor U5185 (N_5185,N_2567,N_3152);
nor U5186 (N_5186,N_4505,N_107);
xnor U5187 (N_5187,N_2646,N_3832);
nor U5188 (N_5188,N_1428,N_4841);
or U5189 (N_5189,N_3194,N_3674);
and U5190 (N_5190,N_1204,N_521);
and U5191 (N_5191,N_1538,N_4895);
and U5192 (N_5192,N_4963,N_577);
nand U5193 (N_5193,N_463,N_468);
and U5194 (N_5194,N_936,N_1288);
nor U5195 (N_5195,N_3825,N_3353);
xor U5196 (N_5196,N_3219,N_4413);
nand U5197 (N_5197,N_351,N_1494);
and U5198 (N_5198,N_1848,N_3763);
and U5199 (N_5199,N_1884,N_1957);
xor U5200 (N_5200,N_346,N_1364);
and U5201 (N_5201,N_1247,N_563);
nand U5202 (N_5202,N_1120,N_623);
or U5203 (N_5203,N_3780,N_1859);
or U5204 (N_5204,N_2104,N_692);
nand U5205 (N_5205,N_1502,N_3233);
or U5206 (N_5206,N_4869,N_1454);
and U5207 (N_5207,N_2380,N_2574);
and U5208 (N_5208,N_3179,N_3962);
and U5209 (N_5209,N_546,N_1398);
and U5210 (N_5210,N_1030,N_2208);
nand U5211 (N_5211,N_3009,N_1287);
xnor U5212 (N_5212,N_2178,N_4896);
nand U5213 (N_5213,N_4632,N_2678);
nor U5214 (N_5214,N_4523,N_4322);
nand U5215 (N_5215,N_4889,N_3203);
or U5216 (N_5216,N_4876,N_1738);
or U5217 (N_5217,N_2994,N_1215);
xor U5218 (N_5218,N_2845,N_1537);
nand U5219 (N_5219,N_18,N_2026);
nor U5220 (N_5220,N_424,N_4064);
and U5221 (N_5221,N_3901,N_4705);
nand U5222 (N_5222,N_725,N_3974);
nor U5223 (N_5223,N_1042,N_3919);
nand U5224 (N_5224,N_4827,N_4271);
xnor U5225 (N_5225,N_4399,N_2613);
xor U5226 (N_5226,N_126,N_1797);
nand U5227 (N_5227,N_3871,N_2868);
xor U5228 (N_5228,N_2111,N_3603);
xnor U5229 (N_5229,N_594,N_4818);
nor U5230 (N_5230,N_2081,N_359);
xor U5231 (N_5231,N_3560,N_3376);
xnor U5232 (N_5232,N_4989,N_389);
or U5233 (N_5233,N_2795,N_2902);
xor U5234 (N_5234,N_404,N_4024);
or U5235 (N_5235,N_3310,N_838);
nor U5236 (N_5236,N_2689,N_2332);
xnor U5237 (N_5237,N_1680,N_2779);
or U5238 (N_5238,N_132,N_3405);
nand U5239 (N_5239,N_4238,N_2592);
nand U5240 (N_5240,N_4656,N_1690);
xor U5241 (N_5241,N_1979,N_2700);
nor U5242 (N_5242,N_2844,N_4479);
nor U5243 (N_5243,N_1718,N_1499);
nor U5244 (N_5244,N_1661,N_3160);
or U5245 (N_5245,N_835,N_4085);
nor U5246 (N_5246,N_2731,N_4254);
or U5247 (N_5247,N_4010,N_4894);
and U5248 (N_5248,N_629,N_1005);
nor U5249 (N_5249,N_3732,N_816);
xor U5250 (N_5250,N_343,N_4716);
nand U5251 (N_5251,N_2476,N_4249);
nand U5252 (N_5252,N_2846,N_1067);
and U5253 (N_5253,N_1133,N_1943);
and U5254 (N_5254,N_658,N_1773);
xnor U5255 (N_5255,N_3944,N_3019);
xnor U5256 (N_5256,N_2393,N_1007);
nand U5257 (N_5257,N_3884,N_1355);
nor U5258 (N_5258,N_4110,N_3468);
nor U5259 (N_5259,N_4490,N_3309);
nor U5260 (N_5260,N_2426,N_1121);
or U5261 (N_5261,N_2511,N_4051);
nand U5262 (N_5262,N_2535,N_1854);
and U5263 (N_5263,N_1542,N_2314);
xnor U5264 (N_5264,N_3840,N_4442);
nand U5265 (N_5265,N_595,N_1130);
xnor U5266 (N_5266,N_341,N_1550);
and U5267 (N_5267,N_2462,N_4043);
xor U5268 (N_5268,N_2067,N_204);
nand U5269 (N_5269,N_3128,N_1561);
nand U5270 (N_5270,N_4398,N_1612);
nor U5271 (N_5271,N_609,N_338);
or U5272 (N_5272,N_2229,N_1857);
nand U5273 (N_5273,N_2214,N_1176);
xor U5274 (N_5274,N_1424,N_73);
or U5275 (N_5275,N_2228,N_4764);
or U5276 (N_5276,N_1628,N_573);
nand U5277 (N_5277,N_2253,N_662);
and U5278 (N_5278,N_1305,N_4843);
and U5279 (N_5279,N_4385,N_4458);
xor U5280 (N_5280,N_4341,N_306);
xor U5281 (N_5281,N_4561,N_2552);
and U5282 (N_5282,N_488,N_1109);
xor U5283 (N_5283,N_1190,N_1480);
or U5284 (N_5284,N_1260,N_2008);
nand U5285 (N_5285,N_2582,N_4281);
nor U5286 (N_5286,N_607,N_3794);
and U5287 (N_5287,N_4585,N_4791);
or U5288 (N_5288,N_3234,N_323);
nand U5289 (N_5289,N_2962,N_2468);
xnor U5290 (N_5290,N_2907,N_3044);
and U5291 (N_5291,N_4886,N_1731);
xnor U5292 (N_5292,N_1582,N_3656);
nand U5293 (N_5293,N_4763,N_2685);
xnor U5294 (N_5294,N_2362,N_1702);
or U5295 (N_5295,N_1564,N_1302);
and U5296 (N_5296,N_1638,N_2059);
nor U5297 (N_5297,N_4500,N_4244);
xor U5298 (N_5298,N_3023,N_4605);
or U5299 (N_5299,N_1039,N_1463);
nand U5300 (N_5300,N_2197,N_2363);
or U5301 (N_5301,N_3446,N_2355);
nand U5302 (N_5302,N_1224,N_4263);
xnor U5303 (N_5303,N_2069,N_1617);
and U5304 (N_5304,N_1372,N_3389);
or U5305 (N_5305,N_3428,N_3346);
xnor U5306 (N_5306,N_1706,N_4616);
or U5307 (N_5307,N_2027,N_2055);
or U5308 (N_5308,N_285,N_2478);
nand U5309 (N_5309,N_4652,N_4803);
xor U5310 (N_5310,N_125,N_799);
nand U5311 (N_5311,N_3415,N_1501);
nand U5312 (N_5312,N_2805,N_976);
or U5313 (N_5313,N_1545,N_2903);
xor U5314 (N_5314,N_1019,N_4132);
and U5315 (N_5315,N_4361,N_560);
xnor U5316 (N_5316,N_4900,N_1301);
or U5317 (N_5317,N_151,N_946);
xor U5318 (N_5318,N_1594,N_1168);
nor U5319 (N_5319,N_1524,N_924);
or U5320 (N_5320,N_2206,N_4157);
xnor U5321 (N_5321,N_2599,N_2391);
xnor U5322 (N_5322,N_3132,N_3192);
or U5323 (N_5323,N_2668,N_2869);
nor U5324 (N_5324,N_4000,N_4663);
nand U5325 (N_5325,N_3525,N_4910);
nor U5326 (N_5326,N_2219,N_2889);
nor U5327 (N_5327,N_2121,N_3010);
nor U5328 (N_5328,N_2251,N_1615);
or U5329 (N_5329,N_50,N_1104);
nor U5330 (N_5330,N_4750,N_4670);
xnor U5331 (N_5331,N_4823,N_4717);
nand U5332 (N_5332,N_2839,N_166);
and U5333 (N_5333,N_993,N_393);
nand U5334 (N_5334,N_749,N_1035);
xnor U5335 (N_5335,N_4362,N_1179);
nor U5336 (N_5336,N_4976,N_221);
xnor U5337 (N_5337,N_2450,N_1665);
nand U5338 (N_5338,N_1445,N_879);
or U5339 (N_5339,N_2237,N_179);
nor U5340 (N_5340,N_3701,N_4642);
and U5341 (N_5341,N_3212,N_2082);
and U5342 (N_5342,N_1698,N_4060);
nor U5343 (N_5343,N_4660,N_3822);
and U5344 (N_5344,N_4911,N_3723);
and U5345 (N_5345,N_1256,N_3361);
nor U5346 (N_5346,N_4069,N_3499);
nand U5347 (N_5347,N_466,N_1711);
and U5348 (N_5348,N_4410,N_2402);
nand U5349 (N_5349,N_3287,N_2407);
and U5350 (N_5350,N_2550,N_3381);
nand U5351 (N_5351,N_3323,N_2758);
nand U5352 (N_5352,N_1716,N_499);
nor U5353 (N_5353,N_3267,N_2860);
nand U5354 (N_5354,N_701,N_1739);
or U5355 (N_5355,N_3471,N_4137);
and U5356 (N_5356,N_2796,N_796);
nand U5357 (N_5357,N_2446,N_2679);
nor U5358 (N_5358,N_4352,N_2192);
or U5359 (N_5359,N_3569,N_3802);
nor U5360 (N_5360,N_4693,N_556);
xnor U5361 (N_5361,N_3550,N_2414);
nor U5362 (N_5362,N_3949,N_2800);
or U5363 (N_5363,N_897,N_1624);
or U5364 (N_5364,N_4344,N_354);
or U5365 (N_5365,N_1897,N_2641);
and U5366 (N_5366,N_1578,N_2972);
nand U5367 (N_5367,N_3842,N_1983);
xor U5368 (N_5368,N_3427,N_3043);
nor U5369 (N_5369,N_2763,N_33);
nor U5370 (N_5370,N_2207,N_1085);
nor U5371 (N_5371,N_1388,N_4411);
nand U5372 (N_5372,N_3990,N_1126);
nand U5373 (N_5373,N_1052,N_1004);
nand U5374 (N_5374,N_3331,N_875);
and U5375 (N_5375,N_2419,N_105);
or U5376 (N_5376,N_954,N_1154);
and U5377 (N_5377,N_1913,N_1946);
xor U5378 (N_5378,N_568,N_1905);
nand U5379 (N_5379,N_2993,N_1294);
or U5380 (N_5380,N_4482,N_2502);
xnor U5381 (N_5381,N_3302,N_1471);
and U5382 (N_5382,N_1324,N_4808);
nand U5383 (N_5383,N_2017,N_4497);
and U5384 (N_5384,N_2619,N_869);
nand U5385 (N_5385,N_4507,N_1318);
xor U5386 (N_5386,N_294,N_3720);
nand U5387 (N_5387,N_756,N_3808);
and U5388 (N_5388,N_186,N_4721);
xor U5389 (N_5389,N_4338,N_1519);
xor U5390 (N_5390,N_3638,N_1725);
nand U5391 (N_5391,N_3947,N_4908);
nor U5392 (N_5392,N_590,N_1784);
xnor U5393 (N_5393,N_461,N_156);
nand U5394 (N_5394,N_399,N_633);
nor U5395 (N_5395,N_947,N_4518);
or U5396 (N_5396,N_2703,N_1783);
and U5397 (N_5397,N_3905,N_1647);
nor U5398 (N_5398,N_446,N_2273);
nor U5399 (N_5399,N_605,N_3460);
or U5400 (N_5400,N_3239,N_2275);
or U5401 (N_5401,N_510,N_2544);
or U5402 (N_5402,N_4683,N_4286);
and U5403 (N_5403,N_3561,N_3426);
and U5404 (N_5404,N_774,N_1629);
and U5405 (N_5405,N_3669,N_2825);
nor U5406 (N_5406,N_4601,N_240);
nor U5407 (N_5407,N_3305,N_3844);
nand U5408 (N_5408,N_2415,N_4508);
or U5409 (N_5409,N_493,N_2074);
nand U5410 (N_5410,N_2987,N_1370);
and U5411 (N_5411,N_1525,N_3216);
or U5412 (N_5412,N_1481,N_329);
and U5413 (N_5413,N_1311,N_579);
or U5414 (N_5414,N_2693,N_3400);
and U5415 (N_5415,N_941,N_846);
nand U5416 (N_5416,N_295,N_3077);
or U5417 (N_5417,N_1207,N_626);
nor U5418 (N_5418,N_788,N_3659);
nand U5419 (N_5419,N_3859,N_1470);
xor U5420 (N_5420,N_286,N_3156);
or U5421 (N_5421,N_704,N_4521);
xor U5422 (N_5422,N_4108,N_1081);
and U5423 (N_5423,N_2034,N_3184);
nor U5424 (N_5424,N_2037,N_801);
or U5425 (N_5425,N_1479,N_2381);
xnor U5426 (N_5426,N_274,N_2935);
and U5427 (N_5427,N_2428,N_2737);
nand U5428 (N_5428,N_316,N_4114);
and U5429 (N_5429,N_3485,N_4555);
xnor U5430 (N_5430,N_4498,N_3547);
nor U5431 (N_5431,N_1834,N_368);
nor U5432 (N_5432,N_624,N_4756);
nor U5433 (N_5433,N_2855,N_3241);
and U5434 (N_5434,N_4968,N_3791);
or U5435 (N_5435,N_69,N_1625);
and U5436 (N_5436,N_789,N_1387);
xnor U5437 (N_5437,N_2186,N_2359);
xnor U5438 (N_5438,N_2549,N_2126);
nor U5439 (N_5439,N_2568,N_4133);
nor U5440 (N_5440,N_860,N_4884);
or U5441 (N_5441,N_1832,N_1143);
or U5442 (N_5442,N_4676,N_4772);
or U5443 (N_5443,N_4621,N_79);
nand U5444 (N_5444,N_970,N_4560);
and U5445 (N_5445,N_1354,N_4532);
xor U5446 (N_5446,N_1200,N_1603);
xor U5447 (N_5447,N_3504,N_1510);
nor U5448 (N_5448,N_12,N_4255);
xor U5449 (N_5449,N_2614,N_4124);
or U5450 (N_5450,N_1780,N_2270);
and U5451 (N_5451,N_3249,N_1458);
and U5452 (N_5452,N_2130,N_2201);
nor U5453 (N_5453,N_3758,N_227);
nor U5454 (N_5454,N_3888,N_593);
and U5455 (N_5455,N_779,N_212);
or U5456 (N_5456,N_1575,N_2073);
nor U5457 (N_5457,N_3040,N_1054);
and U5458 (N_5458,N_2033,N_3745);
or U5459 (N_5459,N_1930,N_3668);
and U5460 (N_5460,N_454,N_1566);
nor U5461 (N_5461,N_4027,N_1319);
or U5462 (N_5462,N_1485,N_3803);
and U5463 (N_5463,N_3103,N_1487);
and U5464 (N_5464,N_885,N_3242);
and U5465 (N_5465,N_2920,N_888);
and U5466 (N_5466,N_4607,N_4455);
xnor U5467 (N_5467,N_3165,N_4813);
xor U5468 (N_5468,N_2798,N_1068);
or U5469 (N_5469,N_2811,N_3574);
nor U5470 (N_5470,N_4431,N_2533);
or U5471 (N_5471,N_2910,N_4877);
or U5472 (N_5472,N_308,N_258);
xnor U5473 (N_5473,N_3125,N_318);
nand U5474 (N_5474,N_2089,N_3262);
or U5475 (N_5475,N_2872,N_2255);
xor U5476 (N_5476,N_3025,N_3162);
or U5477 (N_5477,N_2386,N_1572);
nor U5478 (N_5478,N_1061,N_1977);
and U5479 (N_5479,N_2056,N_690);
nor U5480 (N_5480,N_3885,N_397);
nand U5481 (N_5481,N_4951,N_4001);
or U5482 (N_5482,N_4002,N_4834);
nand U5483 (N_5483,N_3251,N_4);
or U5484 (N_5484,N_729,N_1535);
and U5485 (N_5485,N_678,N_1044);
nand U5486 (N_5486,N_1942,N_3131);
and U5487 (N_5487,N_367,N_2420);
or U5488 (N_5488,N_4857,N_3367);
nand U5489 (N_5489,N_823,N_4454);
nand U5490 (N_5490,N_4144,N_4214);
and U5491 (N_5491,N_1113,N_2099);
nor U5492 (N_5492,N_3831,N_4210);
or U5493 (N_5493,N_634,N_3761);
xor U5494 (N_5494,N_2470,N_1300);
or U5495 (N_5495,N_1291,N_1095);
and U5496 (N_5496,N_4628,N_4576);
nor U5497 (N_5497,N_4526,N_724);
or U5498 (N_5498,N_218,N_1733);
and U5499 (N_5499,N_2327,N_1909);
and U5500 (N_5500,N_1444,N_3407);
or U5501 (N_5501,N_2569,N_983);
nor U5502 (N_5502,N_2175,N_161);
xor U5503 (N_5503,N_163,N_3862);
xnor U5504 (N_5504,N_4731,N_4749);
or U5505 (N_5505,N_2773,N_2617);
nor U5506 (N_5506,N_1598,N_412);
or U5507 (N_5507,N_655,N_2699);
nand U5508 (N_5508,N_3462,N_1565);
nand U5509 (N_5509,N_3716,N_3334);
nor U5510 (N_5510,N_3801,N_3406);
or U5511 (N_5511,N_3898,N_1949);
xnor U5512 (N_5512,N_1790,N_2317);
or U5513 (N_5513,N_253,N_881);
xor U5514 (N_5514,N_22,N_4216);
and U5515 (N_5515,N_500,N_4597);
nor U5516 (N_5516,N_133,N_1837);
nor U5517 (N_5517,N_4931,N_2300);
or U5518 (N_5518,N_3833,N_1678);
xor U5519 (N_5519,N_429,N_3636);
or U5520 (N_5520,N_2677,N_1681);
nand U5521 (N_5521,N_3983,N_1533);
or U5522 (N_5522,N_2751,N_2638);
nand U5523 (N_5523,N_3279,N_1345);
and U5524 (N_5524,N_3943,N_4666);
nand U5525 (N_5525,N_2898,N_2282);
and U5526 (N_5526,N_2727,N_4325);
nor U5527 (N_5527,N_3495,N_438);
nor U5528 (N_5528,N_4487,N_4612);
nor U5529 (N_5529,N_1577,N_2469);
and U5530 (N_5530,N_4269,N_4620);
and U5531 (N_5531,N_4019,N_4083);
xor U5532 (N_5532,N_1346,N_1093);
nand U5533 (N_5533,N_3411,N_964);
xnor U5534 (N_5534,N_3729,N_3188);
and U5535 (N_5535,N_829,N_3824);
nand U5536 (N_5536,N_2633,N_1540);
xor U5537 (N_5537,N_1410,N_3211);
nand U5538 (N_5538,N_3049,N_2545);
xnor U5539 (N_5539,N_3686,N_961);
nor U5540 (N_5540,N_1226,N_391);
or U5541 (N_5541,N_3474,N_2537);
or U5542 (N_5542,N_1870,N_2303);
nand U5543 (N_5543,N_2670,N_3790);
nor U5544 (N_5544,N_1850,N_2927);
nor U5545 (N_5545,N_1889,N_4420);
nor U5546 (N_5546,N_3478,N_3214);
and U5547 (N_5547,N_4218,N_2092);
nor U5548 (N_5548,N_3178,N_1916);
or U5549 (N_5549,N_4516,N_1954);
nand U5550 (N_5550,N_4719,N_1852);
or U5551 (N_5551,N_3110,N_2);
nor U5552 (N_5552,N_4308,N_3750);
and U5553 (N_5553,N_4688,N_2923);
nand U5554 (N_5554,N_2310,N_4119);
and U5555 (N_5555,N_112,N_2833);
and U5556 (N_5556,N_2909,N_3047);
nand U5557 (N_5557,N_586,N_868);
and U5558 (N_5558,N_1998,N_1159);
nor U5559 (N_5559,N_2116,N_2922);
or U5560 (N_5560,N_3443,N_1597);
or U5561 (N_5561,N_4980,N_3829);
xor U5562 (N_5562,N_1484,N_3283);
xnor U5563 (N_5563,N_3284,N_4697);
nand U5564 (N_5564,N_4792,N_492);
and U5565 (N_5565,N_4155,N_449);
nand U5566 (N_5566,N_2114,N_3069);
or U5567 (N_5567,N_3597,N_4197);
or U5568 (N_5568,N_1555,N_2039);
nor U5569 (N_5569,N_3951,N_3810);
nor U5570 (N_5570,N_2937,N_592);
and U5571 (N_5571,N_4883,N_4456);
xor U5572 (N_5572,N_2021,N_2103);
xnor U5573 (N_5573,N_4329,N_4868);
xor U5574 (N_5574,N_2560,N_931);
and U5575 (N_5575,N_854,N_1420);
nor U5576 (N_5576,N_2007,N_2517);
xnor U5577 (N_5577,N_4972,N_4638);
xnor U5578 (N_5578,N_1380,N_952);
and U5579 (N_5579,N_2809,N_2652);
and U5580 (N_5580,N_1556,N_217);
xor U5581 (N_5581,N_1639,N_3118);
or U5582 (N_5582,N_2250,N_4135);
or U5583 (N_5583,N_3017,N_4287);
xor U5584 (N_5584,N_504,N_3065);
or U5585 (N_5585,N_4113,N_1099);
nor U5586 (N_5586,N_2991,N_4179);
and U5587 (N_5587,N_3319,N_4761);
nand U5588 (N_5588,N_2260,N_1693);
and U5589 (N_5589,N_3090,N_1841);
or U5590 (N_5590,N_1580,N_721);
xnor U5591 (N_5591,N_4425,N_3865);
or U5592 (N_5592,N_303,N_4641);
and U5593 (N_5593,N_2353,N_2510);
nor U5594 (N_5594,N_3002,N_4766);
or U5595 (N_5595,N_3213,N_3463);
nand U5596 (N_5596,N_44,N_822);
nor U5597 (N_5597,N_1071,N_37);
nand U5598 (N_5598,N_2906,N_3609);
nor U5599 (N_5599,N_538,N_2085);
or U5600 (N_5600,N_4073,N_3997);
nand U5601 (N_5601,N_4513,N_3864);
and U5602 (N_5602,N_2291,N_3587);
or U5603 (N_5603,N_106,N_1238);
or U5604 (N_5604,N_3628,N_2307);
xnor U5605 (N_5605,N_141,N_4657);
and U5606 (N_5606,N_1409,N_4252);
xnor U5607 (N_5607,N_4474,N_4753);
nand U5608 (N_5608,N_1877,N_3911);
or U5609 (N_5609,N_3067,N_988);
nand U5610 (N_5610,N_4501,N_3036);
nor U5611 (N_5611,N_1105,N_3425);
xnor U5612 (N_5612,N_3631,N_2351);
or U5613 (N_5613,N_3027,N_1464);
nand U5614 (N_5614,N_1193,N_245);
and U5615 (N_5615,N_2254,N_4942);
or U5616 (N_5616,N_4769,N_4822);
xor U5617 (N_5617,N_1344,N_3170);
nand U5618 (N_5618,N_1114,N_1468);
xnor U5619 (N_5619,N_1060,N_1996);
nand U5620 (N_5620,N_747,N_2792);
nor U5621 (N_5621,N_3895,N_4762);
xor U5622 (N_5622,N_1232,N_896);
and U5623 (N_5623,N_2708,N_2011);
nor U5624 (N_5624,N_611,N_4469);
nor U5625 (N_5625,N_3994,N_2122);
and U5626 (N_5626,N_241,N_3817);
nand U5627 (N_5627,N_1974,N_750);
nand U5628 (N_5628,N_873,N_3932);
nand U5629 (N_5629,N_160,N_496);
nand U5630 (N_5630,N_3108,N_2973);
nor U5631 (N_5631,N_3390,N_3264);
nor U5632 (N_5632,N_755,N_3321);
nand U5633 (N_5633,N_1472,N_4812);
and U5634 (N_5634,N_4117,N_3259);
and U5635 (N_5635,N_3646,N_1225);
nor U5636 (N_5636,N_434,N_3436);
or U5637 (N_5637,N_518,N_4459);
nand U5638 (N_5638,N_3972,N_1164);
and U5639 (N_5639,N_207,N_2760);
nor U5640 (N_5640,N_693,N_3324);
nor U5641 (N_5641,N_3041,N_3505);
and U5642 (N_5642,N_2497,N_503);
or U5643 (N_5643,N_3343,N_189);
and U5644 (N_5644,N_480,N_2536);
nor U5645 (N_5645,N_456,N_3655);
or U5646 (N_5646,N_114,N_2051);
nand U5647 (N_5647,N_1325,N_812);
nor U5648 (N_5648,N_3289,N_3948);
xor U5649 (N_5649,N_1732,N_1978);
nor U5650 (N_5650,N_4321,N_2726);
xnor U5651 (N_5651,N_4842,N_1631);
xnor U5652 (N_5652,N_4187,N_2406);
xor U5653 (N_5653,N_384,N_4397);
or U5654 (N_5654,N_1656,N_2952);
nand U5655 (N_5655,N_845,N_2505);
and U5656 (N_5656,N_1363,N_4596);
nor U5657 (N_5657,N_1777,N_1788);
xor U5658 (N_5658,N_2862,N_3258);
and U5659 (N_5659,N_4933,N_469);
nor U5660 (N_5660,N_4855,N_763);
and U5661 (N_5661,N_1087,N_4172);
xor U5662 (N_5662,N_4477,N_1136);
nand U5663 (N_5663,N_96,N_4736);
or U5664 (N_5664,N_1205,N_545);
xor U5665 (N_5665,N_4031,N_1103);
or U5666 (N_5666,N_3466,N_1266);
or U5667 (N_5667,N_1213,N_2451);
or U5668 (N_5668,N_3821,N_3080);
nor U5669 (N_5669,N_4327,N_4627);
nand U5670 (N_5670,N_3508,N_275);
nor U5671 (N_5671,N_101,N_883);
xor U5672 (N_5672,N_2824,N_559);
xnor U5673 (N_5673,N_2344,N_4018);
nand U5674 (N_5674,N_949,N_4703);
and U5675 (N_5675,N_3208,N_1508);
and U5676 (N_5676,N_2383,N_1611);
nand U5677 (N_5677,N_2479,N_1237);
nor U5678 (N_5678,N_3621,N_4165);
nor U5679 (N_5679,N_279,N_3136);
or U5680 (N_5680,N_477,N_1993);
nand U5681 (N_5681,N_4930,N_1056);
nand U5682 (N_5682,N_4940,N_1161);
or U5683 (N_5683,N_937,N_1304);
nand U5684 (N_5684,N_4378,N_2506);
nand U5685 (N_5685,N_2857,N_4139);
nand U5686 (N_5686,N_3940,N_1416);
xor U5687 (N_5687,N_4578,N_2925);
xor U5688 (N_5688,N_4872,N_1469);
and U5689 (N_5689,N_1820,N_2458);
and U5690 (N_5690,N_824,N_612);
xnor U5691 (N_5691,N_4533,N_3416);
nor U5692 (N_5692,N_1373,N_2480);
xnor U5693 (N_5693,N_193,N_1101);
nor U5694 (N_5694,N_2483,N_3384);
nand U5695 (N_5695,N_1635,N_2366);
and U5696 (N_5696,N_4974,N_2891);
or U5697 (N_5697,N_1139,N_2153);
nand U5698 (N_5698,N_977,N_3417);
xnor U5699 (N_5699,N_3534,N_2784);
and U5700 (N_5700,N_4696,N_2672);
or U5701 (N_5701,N_1562,N_585);
nand U5702 (N_5702,N_4195,N_2894);
nand U5703 (N_5703,N_3788,N_4292);
and U5704 (N_5704,N_3526,N_575);
nand U5705 (N_5705,N_2541,N_4864);
nand U5706 (N_5706,N_1880,N_3925);
nor U5707 (N_5707,N_4849,N_4491);
and U5708 (N_5708,N_2002,N_1717);
and U5709 (N_5709,N_4926,N_1008);
or U5710 (N_5710,N_4419,N_3658);
nand U5711 (N_5711,N_3584,N_4551);
xnor U5712 (N_5712,N_1768,N_4319);
nand U5713 (N_5713,N_4875,N_2410);
nand U5714 (N_5714,N_2520,N_3351);
and U5715 (N_5715,N_4256,N_3451);
or U5716 (N_5716,N_2030,N_1233);
nor U5717 (N_5717,N_2583,N_4595);
nor U5718 (N_5718,N_3388,N_2014);
xnor U5719 (N_5719,N_3736,N_4025);
xnor U5720 (N_5720,N_2547,N_3869);
xor U5721 (N_5721,N_4674,N_4260);
nand U5722 (N_5722,N_4961,N_982);
or U5723 (N_5723,N_4472,N_2046);
nor U5724 (N_5724,N_3094,N_2078);
xnor U5725 (N_5725,N_819,N_2887);
nor U5726 (N_5726,N_1994,N_2850);
nor U5727 (N_5727,N_4517,N_4966);
nor U5728 (N_5728,N_2799,N_3698);
and U5729 (N_5729,N_2225,N_3168);
xor U5730 (N_5730,N_2224,N_728);
nor U5731 (N_5731,N_299,N_1769);
xnor U5732 (N_5732,N_1634,N_3570);
nor U5733 (N_5733,N_4105,N_4427);
nand U5734 (N_5734,N_4677,N_3358);
xnor U5735 (N_5735,N_598,N_3374);
nor U5736 (N_5736,N_4251,N_1426);
and U5737 (N_5737,N_2006,N_4939);
or U5738 (N_5738,N_3877,N_3671);
or U5739 (N_5739,N_3256,N_4151);
nor U5740 (N_5740,N_2701,N_4204);
nand U5741 (N_5741,N_3112,N_90);
xnor U5742 (N_5742,N_1055,N_1323);
nor U5743 (N_5743,N_2957,N_2735);
or U5744 (N_5744,N_773,N_1853);
nor U5745 (N_5745,N_4646,N_158);
and U5746 (N_5746,N_3754,N_3487);
xnor U5747 (N_5747,N_3345,N_2753);
or U5748 (N_5748,N_4261,N_4690);
xnor U5749 (N_5749,N_1965,N_1212);
xnor U5750 (N_5750,N_2742,N_2341);
xor U5751 (N_5751,N_4947,N_2236);
and U5752 (N_5752,N_620,N_1116);
nand U5753 (N_5753,N_3744,N_4944);
xnor U5754 (N_5754,N_1079,N_3613);
or U5755 (N_5755,N_2842,N_651);
or U5756 (N_5756,N_1024,N_70);
and U5757 (N_5757,N_2509,N_3913);
nand U5758 (N_5758,N_246,N_4340);
nor U5759 (N_5759,N_3385,N_588);
nand U5760 (N_5760,N_2164,N_513);
nand U5761 (N_5761,N_2518,N_557);
and U5762 (N_5762,N_2643,N_1186);
nand U5763 (N_5763,N_1529,N_2215);
and U5764 (N_5764,N_2739,N_619);
nand U5765 (N_5765,N_3281,N_40);
nand U5766 (N_5766,N_3610,N_706);
or U5767 (N_5767,N_2580,N_382);
nor U5768 (N_5768,N_2942,N_4744);
nor U5769 (N_5769,N_1794,N_512);
nor U5770 (N_5770,N_313,N_572);
and U5771 (N_5771,N_3278,N_2871);
or U5772 (N_5772,N_3751,N_2305);
and U5773 (N_5773,N_4861,N_2247);
xor U5774 (N_5774,N_401,N_293);
nand U5775 (N_5775,N_1330,N_726);
nand U5776 (N_5776,N_39,N_1228);
and U5777 (N_5777,N_4468,N_4182);
nand U5778 (N_5778,N_4380,N_1906);
or U5779 (N_5779,N_1257,N_1879);
or U5780 (N_5780,N_2606,N_1506);
and U5781 (N_5781,N_1559,N_4531);
xnor U5782 (N_5782,N_4602,N_2135);
and U5783 (N_5783,N_1209,N_4360);
nand U5784 (N_5784,N_1483,N_1886);
and U5785 (N_5785,N_4496,N_1595);
xnor U5786 (N_5786,N_1196,N_957);
and U5787 (N_5787,N_3740,N_1536);
xor U5788 (N_5788,N_1527,N_4021);
nand U5789 (N_5789,N_2323,N_876);
nand U5790 (N_5790,N_566,N_4439);
nand U5791 (N_5791,N_2984,N_3596);
or U5792 (N_5792,N_4807,N_3282);
or U5793 (N_5793,N_3921,N_3835);
nor U5794 (N_5794,N_3640,N_4786);
or U5795 (N_5795,N_757,N_3183);
and U5796 (N_5796,N_536,N_4258);
and U5797 (N_5797,N_3029,N_2401);
nor U5798 (N_5798,N_3236,N_1763);
xor U5799 (N_5799,N_4433,N_1037);
xor U5800 (N_5800,N_1695,N_4237);
nor U5801 (N_5801,N_2819,N_2884);
xor U5802 (N_5802,N_3461,N_4023);
nor U5803 (N_5803,N_3511,N_1846);
xor U5804 (N_5804,N_1662,N_1526);
nor U5805 (N_5805,N_3915,N_2526);
or U5806 (N_5806,N_3679,N_2575);
nand U5807 (N_5807,N_4928,N_3910);
and U5808 (N_5808,N_4200,N_135);
or U5809 (N_5809,N_1110,N_3617);
xnor U5810 (N_5810,N_4495,N_1821);
and U5811 (N_5811,N_2299,N_1018);
and U5812 (N_5812,N_1918,N_4389);
and U5813 (N_5813,N_1295,N_3903);
and U5814 (N_5814,N_4473,N_3699);
or U5815 (N_5815,N_940,N_4959);
nor U5816 (N_5816,N_1332,N_302);
nor U5817 (N_5817,N_684,N_2378);
or U5818 (N_5818,N_899,N_458);
nand U5819 (N_5819,N_2822,N_2943);
or U5820 (N_5820,N_200,N_1162);
or U5821 (N_5821,N_874,N_715);
and U5822 (N_5822,N_170,N_739);
nand U5823 (N_5823,N_2501,N_2471);
xnor U5824 (N_5824,N_2492,N_2804);
nor U5825 (N_5825,N_960,N_1010);
or U5826 (N_5826,N_2977,N_922);
or U5827 (N_5827,N_3253,N_2744);
or U5828 (N_5828,N_3799,N_4609);
and U5829 (N_5829,N_3377,N_1263);
and U5830 (N_5830,N_406,N_4709);
and U5831 (N_5831,N_3291,N_2968);
nor U5832 (N_5832,N_3123,N_4826);
and U5833 (N_5833,N_1144,N_4358);
nor U5834 (N_5834,N_476,N_4624);
nor U5835 (N_5835,N_138,N_4554);
or U5836 (N_5836,N_4209,N_497);
or U5837 (N_5837,N_2690,N_439);
xnor U5838 (N_5838,N_1912,N_2764);
nand U5839 (N_5839,N_1489,N_679);
nand U5840 (N_5840,N_3672,N_2985);
nand U5841 (N_5841,N_3767,N_4099);
nor U5842 (N_5842,N_3928,N_4098);
nand U5843 (N_5843,N_3226,N_1956);
or U5844 (N_5844,N_4679,N_1677);
nand U5845 (N_5845,N_326,N_3667);
xor U5846 (N_5846,N_3268,N_2088);
or U5847 (N_5847,N_2724,N_1252);
or U5848 (N_5848,N_4227,N_1327);
nor U5849 (N_5849,N_4831,N_4461);
nor U5850 (N_5850,N_2585,N_1460);
xnor U5851 (N_5851,N_1310,N_129);
or U5852 (N_5852,N_4668,N_3247);
nand U5853 (N_5853,N_27,N_3779);
nor U5854 (N_5854,N_1579,N_4687);
nor U5855 (N_5855,N_2311,N_328);
xor U5856 (N_5856,N_2596,N_3248);
nor U5857 (N_5857,N_3366,N_2877);
nand U5858 (N_5858,N_3827,N_2785);
xnor U5859 (N_5859,N_547,N_2148);
nand U5860 (N_5860,N_3992,N_3429);
nand U5861 (N_5861,N_564,N_3819);
xor U5862 (N_5862,N_4123,N_3737);
xnor U5863 (N_5863,N_4492,N_3602);
nand U5864 (N_5864,N_4799,N_927);
or U5865 (N_5865,N_2755,N_3015);
and U5866 (N_5866,N_2556,N_998);
nor U5867 (N_5867,N_3937,N_4825);
and U5868 (N_5868,N_713,N_2221);
xor U5869 (N_5869,N_3688,N_2312);
or U5870 (N_5870,N_2190,N_2587);
or U5871 (N_5871,N_3741,N_347);
and U5872 (N_5872,N_3055,N_1830);
nand U5873 (N_5873,N_467,N_2892);
or U5874 (N_5874,N_1505,N_1418);
nand U5875 (N_5875,N_710,N_0);
or U5876 (N_5876,N_2806,N_250);
nor U5877 (N_5877,N_4590,N_4185);
and U5878 (N_5878,N_1676,N_3008);
and U5879 (N_5879,N_2783,N_1307);
nor U5880 (N_5880,N_2847,N_195);
nor U5881 (N_5881,N_229,N_2664);
xor U5882 (N_5882,N_3576,N_1606);
nand U5883 (N_5883,N_3387,N_1249);
nand U5884 (N_5884,N_1075,N_3629);
xnor U5885 (N_5885,N_3382,N_3056);
nor U5886 (N_5886,N_805,N_4847);
xnor U5887 (N_5887,N_811,N_3815);
nand U5888 (N_5888,N_943,N_4373);
nand U5889 (N_5889,N_1960,N_2597);
xor U5890 (N_5890,N_2604,N_3364);
or U5891 (N_5891,N_214,N_1856);
nor U5892 (N_5892,N_4049,N_4453);
or U5893 (N_5893,N_432,N_2258);
nand U5894 (N_5894,N_4759,N_3465);
or U5895 (N_5895,N_2174,N_932);
nor U5896 (N_5896,N_1197,N_1453);
and U5897 (N_5897,N_7,N_2474);
or U5898 (N_5898,N_2455,N_1591);
nor U5899 (N_5899,N_4798,N_3517);
or U5900 (N_5900,N_3703,N_4529);
xnor U5901 (N_5901,N_2436,N_929);
or U5902 (N_5902,N_1032,N_509);
and U5903 (N_5903,N_1292,N_3035);
and U5904 (N_5904,N_445,N_2660);
or U5905 (N_5905,N_4093,N_4740);
nor U5906 (N_5906,N_852,N_3151);
xnor U5907 (N_5907,N_2438,N_3099);
or U5908 (N_5908,N_3618,N_209);
and U5909 (N_5909,N_4953,N_4927);
xnor U5910 (N_5910,N_3227,N_4387);
xnor U5911 (N_5911,N_4745,N_3772);
and U5912 (N_5912,N_3393,N_3623);
nor U5913 (N_5913,N_2100,N_4457);
nand U5914 (N_5914,N_3875,N_4074);
or U5915 (N_5915,N_4991,N_1745);
xnor U5916 (N_5916,N_2005,N_17);
or U5917 (N_5917,N_419,N_4773);
xnor U5918 (N_5918,N_958,N_3169);
nor U5919 (N_5919,N_3626,N_1123);
and U5920 (N_5920,N_3633,N_410);
or U5921 (N_5921,N_3728,N_2449);
and U5922 (N_5922,N_1396,N_2086);
xor U5923 (N_5923,N_3143,N_1642);
nor U5924 (N_5924,N_3543,N_98);
nor U5925 (N_5925,N_1911,N_1645);
nand U5926 (N_5926,N_863,N_124);
or U5927 (N_5927,N_407,N_3770);
and U5928 (N_5928,N_1828,N_3982);
xor U5929 (N_5929,N_1920,N_2995);
nor U5930 (N_5930,N_1618,N_242);
and U5931 (N_5931,N_1673,N_2863);
nand U5932 (N_5932,N_3900,N_4776);
nor U5933 (N_5933,N_4181,N_4176);
nor U5934 (N_5934,N_4704,N_4919);
or U5935 (N_5935,N_4006,N_3542);
nand U5936 (N_5936,N_748,N_1737);
xnor U5937 (N_5937,N_4240,N_2508);
or U5938 (N_5938,N_4770,N_666);
nand U5939 (N_5939,N_1243,N_3747);
and U5940 (N_5940,N_1394,N_1254);
nand U5941 (N_5941,N_1268,N_282);
nor U5942 (N_5942,N_383,N_2188);
or U5943 (N_5943,N_4421,N_3532);
and U5944 (N_5944,N_1888,N_1498);
nand U5945 (N_5945,N_3467,N_4056);
or U5946 (N_5946,N_314,N_4052);
nand U5947 (N_5947,N_324,N_3858);
nor U5948 (N_5948,N_311,N_36);
xor U5949 (N_5949,N_10,N_4637);
xnor U5950 (N_5950,N_3365,N_4401);
nor U5951 (N_5951,N_3726,N_3506);
xnor U5952 (N_5952,N_364,N_2210);
nor U5953 (N_5953,N_3438,N_1150);
nor U5954 (N_5954,N_3193,N_3555);
nand U5955 (N_5955,N_2048,N_3320);
or U5956 (N_5956,N_4747,N_4905);
xor U5957 (N_5957,N_3489,N_1819);
nand U5958 (N_5958,N_2220,N_3204);
nand U5959 (N_5959,N_1833,N_1778);
nand U5960 (N_5960,N_3689,N_4264);
or U5961 (N_5961,N_4571,N_2465);
or U5962 (N_5962,N_3003,N_3066);
or U5963 (N_5963,N_953,N_3402);
xor U5964 (N_5964,N_4600,N_2736);
xnor U5965 (N_5965,N_2418,N_1824);
and U5966 (N_5966,N_1630,N_591);
and U5967 (N_5967,N_3993,N_374);
or U5968 (N_5968,N_505,N_211);
xor U5969 (N_5969,N_1584,N_4794);
nor U5970 (N_5970,N_3725,N_191);
xnor U5971 (N_5971,N_1814,N_3697);
nor U5972 (N_5972,N_19,N_4120);
xnor U5973 (N_5973,N_4424,N_1493);
and U5974 (N_5974,N_1815,N_3084);
nor U5975 (N_5975,N_702,N_2801);
nor U5976 (N_5976,N_2620,N_3535);
xnor U5977 (N_5977,N_956,N_1174);
or U5978 (N_5978,N_3848,N_3483);
nor U5979 (N_5979,N_4732,N_1720);
or U5980 (N_5980,N_1511,N_3868);
xnor U5981 (N_5981,N_1063,N_3624);
and U5982 (N_5982,N_206,N_4550);
and U5983 (N_5983,N_4178,N_4464);
nand U5984 (N_5984,N_2566,N_4589);
xor U5985 (N_5985,N_2940,N_301);
nand U5986 (N_5986,N_2590,N_355);
or U5987 (N_5987,N_4226,N_34);
nor U5988 (N_5988,N_3590,N_2837);
nand U5989 (N_5989,N_300,N_3598);
or U5990 (N_5990,N_26,N_2914);
or U5991 (N_5991,N_2430,N_2761);
nor U5992 (N_5992,N_2669,N_3857);
nand U5993 (N_5993,N_877,N_1522);
nand U5994 (N_5994,N_1264,N_4613);
or U5995 (N_5995,N_3458,N_700);
nor U5996 (N_5996,N_2068,N_2149);
xnor U5997 (N_5997,N_1423,N_3976);
nor U5998 (N_5998,N_1750,N_534);
or U5999 (N_5999,N_4409,N_35);
nand U6000 (N_6000,N_479,N_322);
nand U6001 (N_6001,N_3139,N_1167);
nor U6002 (N_6002,N_4821,N_4836);
nand U6003 (N_6003,N_238,N_2709);
xnor U6004 (N_6004,N_1129,N_3435);
nor U6005 (N_6005,N_1574,N_3422);
nand U6006 (N_6006,N_2187,N_2360);
nor U6007 (N_6007,N_4904,N_2976);
or U6008 (N_6008,N_4898,N_3593);
nand U6009 (N_6009,N_4323,N_2684);
nand U6010 (N_6010,N_4838,N_4276);
and U6011 (N_6011,N_1795,N_1320);
xnor U6012 (N_6012,N_4993,N_136);
or U6013 (N_6013,N_411,N_3033);
nand U6014 (N_6014,N_1899,N_975);
xor U6015 (N_6015,N_3691,N_3980);
xor U6016 (N_6016,N_1664,N_3988);
and U6017 (N_6017,N_3317,N_1208);
nor U6018 (N_6018,N_2287,N_482);
or U6019 (N_6019,N_2009,N_2666);
nor U6020 (N_6020,N_4365,N_74);
xnor U6021 (N_6021,N_906,N_333);
and U6022 (N_6022,N_3150,N_3295);
nor U6023 (N_6023,N_3906,N_2080);
and U6024 (N_6024,N_1206,N_1932);
or U6025 (N_6025,N_3849,N_2948);
xor U6026 (N_6026,N_2232,N_4440);
nand U6027 (N_6027,N_2233,N_2803);
nand U6028 (N_6028,N_4314,N_532);
nand U6029 (N_6029,N_576,N_772);
and U6030 (N_6030,N_4556,N_268);
xor U6031 (N_6031,N_453,N_4815);
or U6032 (N_6032,N_3595,N_4050);
and U6033 (N_6033,N_3158,N_4755);
nand U6034 (N_6034,N_3743,N_2144);
nor U6035 (N_6035,N_3149,N_910);
and U6036 (N_6036,N_1811,N_2165);
xnor U6037 (N_6037,N_464,N_3931);
nand U6038 (N_6038,N_373,N_4443);
xnor U6039 (N_6039,N_3909,N_2444);
xor U6040 (N_6040,N_4107,N_3052);
nor U6041 (N_6041,N_288,N_1184);
and U6042 (N_6042,N_2729,N_507);
nand U6043 (N_6043,N_2832,N_3565);
and U6044 (N_6044,N_3215,N_4333);
and U6045 (N_6045,N_1082,N_1742);
nor U6046 (N_6046,N_1309,N_717);
xnor U6047 (N_6047,N_562,N_3704);
nand U6048 (N_6048,N_1586,N_3034);
nor U6049 (N_6049,N_4619,N_865);
nor U6050 (N_6050,N_1962,N_1000);
nand U6051 (N_6051,N_3048,N_1829);
or U6052 (N_6052,N_266,N_1350);
or U6053 (N_6053,N_3886,N_47);
nand U6054 (N_6054,N_415,N_2859);
and U6055 (N_6055,N_1476,N_257);
nor U6056 (N_6056,N_1199,N_1655);
nor U6057 (N_6057,N_4681,N_30);
and U6058 (N_6058,N_2061,N_72);
nand U6059 (N_6059,N_2901,N_1371);
nand U6060 (N_6060,N_2589,N_1646);
xor U6061 (N_6061,N_1020,N_1663);
or U6062 (N_6062,N_15,N_1553);
or U6063 (N_6063,N_3409,N_220);
and U6064 (N_6064,N_3031,N_3161);
xor U6065 (N_6065,N_4949,N_1437);
and U6066 (N_6066,N_2756,N_4970);
nand U6067 (N_6067,N_2392,N_2888);
nor U6068 (N_6068,N_4912,N_3544);
nand U6069 (N_6069,N_1961,N_2272);
xnor U6070 (N_6070,N_1455,N_1984);
and U6071 (N_6071,N_3978,N_1908);
or U6072 (N_6072,N_2108,N_2870);
and U6073 (N_6073,N_3600,N_4958);
nor U6074 (N_6074,N_3255,N_2826);
or U6075 (N_6075,N_4852,N_3493);
nor U6076 (N_6076,N_4462,N_4937);
nand U6077 (N_6077,N_3294,N_3328);
nor U6078 (N_6078,N_2649,N_2090);
or U6079 (N_6079,N_4840,N_4639);
nand U6080 (N_6080,N_3348,N_4559);
nor U6081 (N_6081,N_4783,N_2667);
and U6082 (N_6082,N_648,N_1900);
nor U6083 (N_6083,N_3037,N_1356);
and U6084 (N_6084,N_4206,N_2263);
nand U6085 (N_6085,N_3696,N_1976);
or U6086 (N_6086,N_3018,N_3719);
nand U6087 (N_6087,N_1040,N_2023);
and U6088 (N_6088,N_861,N_558);
nor U6089 (N_6089,N_1147,N_1855);
or U6090 (N_6090,N_1111,N_1792);
nor U6091 (N_6091,N_1975,N_4520);
or U6092 (N_6092,N_1951,N_2454);
nand U6093 (N_6093,N_3177,N_3746);
xnor U6094 (N_6094,N_2283,N_2213);
nand U6095 (N_6095,N_4130,N_1626);
xnor U6096 (N_6096,N_3769,N_4219);
xor U6097 (N_6097,N_695,N_1377);
nand U6098 (N_6098,N_1775,N_2308);
nor U6099 (N_6099,N_450,N_1684);
and U6100 (N_6100,N_4078,N_1649);
or U6101 (N_6101,N_1995,N_3141);
xnor U6102 (N_6102,N_2905,N_4720);
and U6103 (N_6103,N_3424,N_4205);
and U6104 (N_6104,N_4694,N_4684);
nand U6105 (N_6105,N_4275,N_3573);
nor U6106 (N_6106,N_1157,N_2298);
nor U6107 (N_6107,N_3967,N_4418);
nor U6108 (N_6108,N_3530,N_80);
nand U6109 (N_6109,N_683,N_2274);
nor U6110 (N_6110,N_714,N_4109);
nor U6111 (N_6111,N_2354,N_4315);
xnor U6112 (N_6112,N_3115,N_4879);
nand U6113 (N_6113,N_4580,N_1560);
and U6114 (N_6114,N_4615,N_1546);
nand U6115 (N_6115,N_2066,N_2999);
nand U6116 (N_6116,N_2881,N_3662);
or U6117 (N_6117,N_1567,N_996);
xnor U6118 (N_6118,N_2496,N_2096);
or U6119 (N_6119,N_3516,N_3386);
nand U6120 (N_6120,N_2591,N_3134);
xnor U6121 (N_6121,N_1798,N_2028);
nand U6122 (N_6122,N_3225,N_137);
nor U6123 (N_6123,N_2834,N_2941);
or U6124 (N_6124,N_925,N_4631);
nand U6125 (N_6125,N_3789,N_2576);
xnor U6126 (N_6126,N_2697,N_3904);
xor U6127 (N_6127,N_2623,N_4534);
and U6128 (N_6128,N_2823,N_2954);
nand U6129 (N_6129,N_388,N_1195);
or U6130 (N_6130,N_352,N_1803);
xnor U6131 (N_6131,N_2712,N_2070);
and U6132 (N_6132,N_1904,N_3181);
and U6133 (N_6133,N_1862,N_1967);
nand U6134 (N_6134,N_3481,N_3396);
nand U6135 (N_6135,N_4633,N_4524);
xnor U6136 (N_6136,N_4689,N_4973);
nand U6137 (N_6137,N_4866,N_1528);
nand U6138 (N_6138,N_4022,N_1011);
nor U6139 (N_6139,N_4994,N_312);
and U6140 (N_6140,N_1048,N_1092);
xor U6141 (N_6141,N_2538,N_187);
or U6142 (N_6142,N_3199,N_2746);
xnor U6143 (N_6143,N_1923,N_4005);
nand U6144 (N_6144,N_3874,N_1158);
and U6145 (N_6145,N_2316,N_3845);
nor U6146 (N_6146,N_2493,N_3159);
and U6147 (N_6147,N_3714,N_4175);
nor U6148 (N_6148,N_2012,N_4388);
xor U6149 (N_6149,N_310,N_800);
nor U6150 (N_6150,N_1898,N_4095);
xor U6151 (N_6151,N_2647,N_413);
nand U6152 (N_6152,N_1721,N_1589);
nor U6153 (N_6153,N_3246,N_3501);
or U6154 (N_6154,N_2482,N_4170);
nand U6155 (N_6155,N_1169,N_2377);
and U6156 (N_6156,N_2400,N_4248);
xnor U6157 (N_6157,N_422,N_1674);
nand U6158 (N_6158,N_4080,N_834);
nor U6159 (N_6159,N_942,N_3298);
and U6160 (N_6160,N_4239,N_3768);
or U6161 (N_6161,N_4407,N_1581);
nor U6162 (N_6162,N_1286,N_4213);
and U6163 (N_6163,N_828,N_3313);
and U6164 (N_6164,N_1171,N_4549);
and U6165 (N_6165,N_88,N_1650);
nand U6166 (N_6166,N_3970,N_2815);
nor U6167 (N_6167,N_524,N_1028);
and U6168 (N_6168,N_1627,N_4801);
xor U6169 (N_6169,N_2754,N_870);
nand U6170 (N_6170,N_3773,N_3421);
nor U6171 (N_6171,N_793,N_420);
xnor U6172 (N_6172,N_1385,N_857);
and U6173 (N_6173,N_2179,N_1490);
or U6174 (N_6174,N_4538,N_1435);
and U6175 (N_6175,N_4707,N_3022);
or U6176 (N_6176,N_65,N_262);
and U6177 (N_6177,N_465,N_4081);
nand U6178 (N_6178,N_2930,N_4235);
and U6179 (N_6179,N_674,N_1175);
nand U6180 (N_6180,N_3205,N_2553);
nor U6181 (N_6181,N_2318,N_641);
nand U6182 (N_6182,N_4318,N_320);
nand U6183 (N_6183,N_148,N_4781);
nor U6184 (N_6184,N_951,N_298);
nor U6185 (N_6185,N_661,N_4775);
nand U6186 (N_6186,N_4921,N_2904);
or U6187 (N_6187,N_2199,N_3687);
and U6188 (N_6188,N_4293,N_3793);
nand U6189 (N_6189,N_3572,N_1276);
xnor U6190 (N_6190,N_1864,N_3664);
or U6191 (N_6191,N_1686,N_4787);
nand U6192 (N_6192,N_4332,N_4950);
and U6193 (N_6193,N_4494,N_3670);
nand U6194 (N_6194,N_2874,N_1735);
nor U6195 (N_6195,N_83,N_3372);
nor U6196 (N_6196,N_4167,N_672);
nor U6197 (N_6197,N_1329,N_2618);
nand U6198 (N_6198,N_746,N_3887);
xnor U6199 (N_6199,N_920,N_1876);
xnor U6200 (N_6200,N_2880,N_3408);
and U6201 (N_6201,N_4039,N_255);
or U6202 (N_6202,N_2725,N_1488);
and U6203 (N_6203,N_1382,N_847);
nor U6204 (N_6204,N_4339,N_1442);
nor U6205 (N_6205,N_3378,N_4250);
nor U6206 (N_6206,N_4089,N_1107);
nor U6207 (N_6207,N_3202,N_2079);
xnor U6208 (N_6208,N_1800,N_4804);
nor U6209 (N_6209,N_4351,N_3581);
nand U6210 (N_6210,N_185,N_1813);
xnor U6211 (N_6211,N_2168,N_1843);
or U6212 (N_6212,N_3563,N_3391);
xor U6213 (N_6213,N_1825,N_4145);
or U6214 (N_6214,N_46,N_3163);
xor U6215 (N_6215,N_3707,N_3583);
xor U6216 (N_6216,N_165,N_4648);
nand U6217 (N_6217,N_3333,N_325);
nand U6218 (N_6218,N_3930,N_4134);
or U6219 (N_6219,N_646,N_259);
and U6220 (N_6220,N_4511,N_130);
and U6221 (N_6221,N_3148,N_2835);
nor U6222 (N_6222,N_4514,N_3250);
xnor U6223 (N_6223,N_3286,N_2481);
or U6224 (N_6224,N_4077,N_1335);
or U6225 (N_6225,N_2577,N_3559);
xnor U6226 (N_6226,N_3615,N_1707);
and U6227 (N_6227,N_912,N_414);
nor U6228 (N_6228,N_771,N_2429);
or U6229 (N_6229,N_4396,N_1945);
nor U6230 (N_6230,N_91,N_694);
nand U6231 (N_6231,N_1277,N_3955);
nand U6232 (N_6232,N_3853,N_3956);
and U6233 (N_6233,N_1919,N_2403);
nor U6234 (N_6234,N_2217,N_1741);
nand U6235 (N_6235,N_2000,N_3370);
nand U6236 (N_6236,N_1012,N_3038);
and U6237 (N_6237,N_2280,N_4742);
xor U6238 (N_6238,N_3734,N_2371);
and U6239 (N_6239,N_1446,N_506);
nand U6240 (N_6240,N_4587,N_4070);
nand U6241 (N_6241,N_765,N_2908);
xnor U6242 (N_6242,N_3059,N_280);
nand U6243 (N_6243,N_3058,N_2399);
nand U6244 (N_6244,N_4183,N_4795);
xnor U6245 (N_6245,N_3644,N_4984);
nor U6246 (N_6246,N_1744,N_2603);
nand U6247 (N_6247,N_4586,N_4941);
xnor U6248 (N_6248,N_3173,N_2110);
nand U6249 (N_6249,N_4988,N_1997);
and U6250 (N_6250,N_778,N_1336);
or U6251 (N_6251,N_4754,N_2790);
xnor U6252 (N_6252,N_2528,N_1675);
or U6253 (N_6253,N_775,N_1235);
nand U6254 (N_6254,N_4429,N_4685);
xor U6255 (N_6255,N_4347,N_4414);
and U6256 (N_6256,N_1714,N_4403);
nand U6257 (N_6257,N_1929,N_1089);
xnor U6258 (N_6258,N_2494,N_1314);
and U6259 (N_6259,N_3731,N_3585);
xnor U6260 (N_6260,N_2720,N_2719);
or U6261 (N_6261,N_3238,N_804);
or U6262 (N_6262,N_840,N_1383);
nor U6263 (N_6263,N_4100,N_3195);
xor U6264 (N_6264,N_455,N_487);
nand U6265 (N_6265,N_1156,N_2083);
xor U6266 (N_6266,N_1160,N_1359);
and U6267 (N_6267,N_769,N_1934);
xnor U6268 (N_6268,N_4733,N_4611);
nand U6269 (N_6269,N_4543,N_4512);
and U6270 (N_6270,N_3649,N_309);
and U6271 (N_6271,N_4288,N_2504);
or U6272 (N_6272,N_501,N_1303);
nor U6273 (N_6273,N_4186,N_4141);
or U6274 (N_6274,N_891,N_3920);
nor U6275 (N_6275,N_3786,N_4221);
nand U6276 (N_6276,N_905,N_31);
and U6277 (N_6277,N_1229,N_2297);
xnor U6278 (N_6278,N_277,N_1816);
nand U6279 (N_6279,N_2350,N_2594);
and U6280 (N_6280,N_3252,N_2319);
nand U6281 (N_6281,N_802,N_3318);
and U6282 (N_6282,N_991,N_2807);
xnor U6283 (N_6283,N_3894,N_2938);
nand U6284 (N_6284,N_3601,N_4669);
nor U6285 (N_6285,N_1970,N_1938);
nand U6286 (N_6286,N_4779,N_3232);
or U6287 (N_6287,N_4234,N_535);
xnor U6288 (N_6288,N_2584,N_3523);
nand U6289 (N_6289,N_4862,N_1475);
nand U6290 (N_6290,N_3564,N_205);
nand U6291 (N_6291,N_3001,N_1290);
xor U6292 (N_6292,N_1415,N_3700);
nand U6293 (N_6293,N_215,N_601);
xnor U6294 (N_6294,N_4192,N_4028);
nand U6295 (N_6295,N_3546,N_3430);
xor U6296 (N_6296,N_2445,N_4118);
xnor U6297 (N_6297,N_4406,N_2338);
and U6298 (N_6298,N_2683,N_821);
nor U6299 (N_6299,N_4160,N_2448);
or U6300 (N_6300,N_1094,N_4253);
or U6301 (N_6301,N_3958,N_123);
and U6302 (N_6302,N_4007,N_3454);
nand U6303 (N_6303,N_2185,N_4810);
nor U6304 (N_6304,N_1441,N_719);
nand U6305 (N_6305,N_554,N_1875);
nor U6306 (N_6306,N_348,N_791);
nor U6307 (N_6307,N_2013,N_2829);
and U6308 (N_6308,N_720,N_2031);
and U6309 (N_6309,N_3541,N_2516);
or U6310 (N_6310,N_884,N_2598);
or U6311 (N_6311,N_643,N_1861);
or U6312 (N_6312,N_3625,N_4309);
or U6313 (N_6313,N_3710,N_4486);
nor U6314 (N_6314,N_4445,N_1986);
xnor U6315 (N_6315,N_2326,N_978);
nor U6316 (N_6316,N_2095,N_1827);
xor U6317 (N_6317,N_3712,N_4510);
nand U6318 (N_6318,N_1712,N_1341);
nand U6319 (N_6319,N_447,N_2953);
or U6320 (N_6320,N_640,N_2658);
and U6321 (N_6321,N_4466,N_2688);
and U6322 (N_6322,N_742,N_900);
nor U6323 (N_6323,N_3735,N_3071);
or U6324 (N_6324,N_4079,N_4087);
xor U6325 (N_6325,N_844,N_1786);
nor U6326 (N_6326,N_3776,N_1462);
nor U6327 (N_6327,N_1188,N_4381);
or U6328 (N_6328,N_1532,N_1936);
nand U6329 (N_6329,N_3362,N_1807);
or U6330 (N_6330,N_1842,N_3538);
and U6331 (N_6331,N_2890,N_4805);
or U6332 (N_6332,N_1610,N_2838);
and U6333 (N_6333,N_1882,N_2732);
or U6334 (N_6334,N_760,N_4488);
xor U6335 (N_6335,N_3682,N_4163);
nor U6336 (N_6336,N_4046,N_4036);
and U6337 (N_6337,N_3757,N_3823);
xnor U6338 (N_6338,N_2413,N_3533);
nand U6339 (N_6339,N_3113,N_3085);
nor U6340 (N_6340,N_766,N_3855);
or U6341 (N_6341,N_3981,N_417);
xor U6342 (N_6342,N_898,N_3418);
xnor U6343 (N_6343,N_2379,N_2087);
or U6344 (N_6344,N_486,N_1244);
and U6345 (N_6345,N_3814,N_2369);
nand U6346 (N_6346,N_735,N_2563);
and U6347 (N_6347,N_625,N_2851);
nor U6348 (N_6348,N_2170,N_4946);
nand U6349 (N_6349,N_1808,N_3207);
or U6350 (N_6350,N_1173,N_4700);
or U6351 (N_6351,N_2883,N_4193);
xor U6352 (N_6352,N_377,N_3137);
xor U6353 (N_6353,N_3300,N_4680);
xor U6354 (N_6354,N_2169,N_1421);
nand U6355 (N_6355,N_4835,N_3063);
xnor U6356 (N_6356,N_56,N_2632);
nor U6357 (N_6357,N_1516,N_878);
nand U6358 (N_6358,N_926,N_1003);
nor U6359 (N_6359,N_3196,N_1883);
nor U6360 (N_6360,N_1220,N_3880);
nand U6361 (N_6361,N_4121,N_4996);
or U6362 (N_6362,N_1102,N_474);
xnor U6363 (N_6363,N_2947,N_4828);
nand U6364 (N_6364,N_2306,N_2242);
xor U6365 (N_6365,N_2861,N_1255);
nand U6366 (N_6366,N_1705,N_2439);
nand U6367 (N_6367,N_3834,N_25);
nand U6368 (N_6368,N_1366,N_531);
xnor U6369 (N_6369,N_4122,N_3337);
xnor U6370 (N_6370,N_63,N_174);
nand U6371 (N_6371,N_543,N_1347);
nor U6372 (N_6372,N_3312,N_1316);
nand U6373 (N_6373,N_4465,N_1941);
and U6374 (N_6374,N_3846,N_2789);
xor U6375 (N_6375,N_3580,N_1002);
and U6376 (N_6376,N_2740,N_1648);
or U6377 (N_6377,N_405,N_4645);
nand U6378 (N_6378,N_2128,N_4009);
nand U6379 (N_6379,N_198,N_1340);
nor U6380 (N_6380,N_3545,N_315);
xnor U6381 (N_6381,N_2551,N_4146);
xor U6382 (N_6382,N_1823,N_3540);
xnor U6383 (N_6383,N_4992,N_1384);
nor U6384 (N_6384,N_2966,N_859);
nor U6385 (N_6385,N_3571,N_1270);
nand U6386 (N_6386,N_4575,N_52);
and U6387 (N_6387,N_744,N_4377);
xor U6388 (N_6388,N_3124,N_1064);
nor U6389 (N_6389,N_2257,N_4797);
nand U6390 (N_6390,N_862,N_3718);
nor U6391 (N_6391,N_3784,N_2238);
nor U6392 (N_6392,N_1447,N_730);
and U6393 (N_6393,N_381,N_2778);
nor U6394 (N_6394,N_3327,N_1709);
nand U6395 (N_6395,N_855,N_2133);
or U6396 (N_6396,N_270,N_738);
and U6397 (N_6397,N_3,N_3419);
nor U6398 (N_6398,N_2472,N_213);
and U6399 (N_6399,N_553,N_786);
and U6400 (N_6400,N_394,N_3144);
or U6401 (N_6401,N_4044,N_2337);
xor U6402 (N_6402,N_1153,N_4887);
or U6403 (N_6403,N_3079,N_752);
and U6404 (N_6404,N_3775,N_2924);
nor U6405 (N_6405,N_2741,N_1959);
nor U6406 (N_6406,N_3155,N_4588);
nand U6407 (N_6407,N_3721,N_2477);
nor U6408 (N_6408,N_3797,N_2348);
xnor U6409 (N_6409,N_3717,N_426);
and U6410 (N_6410,N_4860,N_1590);
nor U6411 (N_6411,N_2707,N_1452);
and U6412 (N_6412,N_3260,N_4636);
xnor U6413 (N_6413,N_1231,N_1337);
or U6414 (N_6414,N_3635,N_1172);
nand U6415 (N_6415,N_3153,N_3455);
nand U6416 (N_6416,N_2093,N_4408);
nand U6417 (N_6417,N_2180,N_2065);
nand U6418 (N_6418,N_3579,N_4935);
or U6419 (N_6419,N_4436,N_2728);
and U6420 (N_6420,N_4067,N_1267);
nor U6421 (N_6421,N_1041,N_2189);
nand U6422 (N_6422,N_3760,N_2457);
and U6423 (N_6423,N_1544,N_2163);
or U6424 (N_6424,N_271,N_3945);
nor U6425 (N_6425,N_787,N_2125);
xor U6426 (N_6426,N_284,N_2226);
or U6427 (N_6427,N_872,N_2916);
and U6428 (N_6428,N_3082,N_261);
nand U6429 (N_6429,N_3675,N_3665);
or U6430 (N_6430,N_1869,N_4978);
and U6431 (N_6431,N_2900,N_3528);
nor U6432 (N_6432,N_2131,N_386);
and U6433 (N_6433,N_4300,N_3828);
nor U6434 (N_6434,N_1972,N_3412);
nand U6435 (N_6435,N_3130,N_3708);
or U6436 (N_6436,N_155,N_1592);
and U6437 (N_6437,N_444,N_882);
and U6438 (N_6438,N_2432,N_1793);
or U6439 (N_6439,N_3509,N_4088);
and U6440 (N_6440,N_990,N_4037);
or U6441 (N_6441,N_4290,N_677);
or U6442 (N_6442,N_1151,N_1146);
xor U6443 (N_6443,N_427,N_3809);
or U6444 (N_6444,N_2608,N_2370);
nor U6445 (N_6445,N_4357,N_2245);
and U6446 (N_6446,N_3582,N_1033);
nor U6447 (N_6447,N_92,N_4354);
and U6448 (N_6448,N_2058,N_2777);
xor U6449 (N_6449,N_1571,N_3554);
and U6450 (N_6450,N_4447,N_4817);
nor U6451 (N_6451,N_4102,N_4614);
nand U6452 (N_6452,N_3269,N_798);
nand U6453 (N_6453,N_4502,N_4302);
nand U6454 (N_6454,N_4233,N_4751);
xnor U6455 (N_6455,N_502,N_4131);
and U6456 (N_6456,N_3781,N_2060);
nor U6457 (N_6457,N_621,N_670);
nor U6458 (N_6458,N_1043,N_2094);
xor U6459 (N_6459,N_2498,N_3605);
or U6460 (N_6460,N_2356,N_1246);
nand U6461 (N_6461,N_2996,N_3694);
and U6462 (N_6462,N_3122,N_1166);
nor U6463 (N_6463,N_817,N_1036);
and U6464 (N_6464,N_4236,N_2540);
nor U6465 (N_6465,N_4416,N_1988);
and U6466 (N_6466,N_1895,N_4653);
and U6467 (N_6467,N_1165,N_2989);
xnor U6468 (N_6468,N_1530,N_537);
nand U6469 (N_6469,N_1687,N_4567);
and U6470 (N_6470,N_4735,N_1804);
nor U6471 (N_6471,N_3998,N_2827);
nand U6472 (N_6472,N_3836,N_2288);
or U6473 (N_6473,N_233,N_1399);
xor U6474 (N_6474,N_3206,N_1001);
or U6475 (N_6475,N_3648,N_4557);
nand U6476 (N_6476,N_4914,N_2202);
nor U6477 (N_6477,N_2372,N_342);
nor U6478 (N_6478,N_436,N_3575);
xor U6479 (N_6479,N_831,N_1491);
and U6480 (N_6480,N_3586,N_2102);
or U6481 (N_6481,N_2320,N_2395);
xnor U6482 (N_6482,N_4954,N_3373);
xnor U6483 (N_6483,N_4712,N_944);
or U6484 (N_6484,N_669,N_4312);
xnor U6485 (N_6485,N_1397,N_1403);
nor U6486 (N_6486,N_3011,N_3311);
and U6487 (N_6487,N_969,N_1658);
xor U6488 (N_6488,N_2152,N_1407);
xor U6489 (N_6489,N_3316,N_712);
or U6490 (N_6490,N_813,N_396);
xor U6491 (N_6491,N_2557,N_3985);
nor U6492 (N_6492,N_4809,N_3315);
nor U6493 (N_6493,N_2244,N_4846);
nor U6494 (N_6494,N_2292,N_768);
or U6495 (N_6495,N_1148,N_3486);
nor U6496 (N_6496,N_1831,N_478);
and U6497 (N_6497,N_4202,N_4865);
nor U6498 (N_6498,N_3371,N_1027);
or U6499 (N_6499,N_1353,N_2266);
nor U6500 (N_6500,N_3759,N_4820);
nand U6501 (N_6501,N_2581,N_4979);
and U6502 (N_6502,N_1903,N_4691);
nand U6503 (N_6503,N_3350,N_62);
nand U6504 (N_6504,N_673,N_1799);
nand U6505 (N_6505,N_4558,N_1921);
nor U6506 (N_6506,N_71,N_3841);
nor U6507 (N_6507,N_2216,N_4065);
xor U6508 (N_6508,N_1683,N_2840);
xnor U6509 (N_6509,N_283,N_4142);
nand U6510 (N_6510,N_3081,N_3607);
or U6511 (N_6511,N_1736,N_291);
nor U6512 (N_6512,N_4382,N_4708);
xnor U6513 (N_6513,N_783,N_2521);
or U6514 (N_6514,N_2374,N_2926);
nor U6515 (N_6515,N_837,N_1952);
and U6516 (N_6516,N_54,N_907);
nand U6517 (N_6517,N_85,N_4758);
and U6518 (N_6518,N_583,N_599);
or U6519 (N_6519,N_550,N_4304);
or U6520 (N_6520,N_1726,N_2911);
or U6521 (N_6521,N_4311,N_4741);
or U6522 (N_6522,N_4063,N_2808);
xnor U6523 (N_6523,N_4072,N_2335);
nor U6524 (N_6524,N_3138,N_2530);
nand U6525 (N_6525,N_1433,N_1299);
and U6526 (N_6526,N_815,N_2016);
or U6527 (N_6527,N_2140,N_4833);
nor U6528 (N_6528,N_29,N_1378);
nor U6529 (N_6529,N_2427,N_1872);
nor U6530 (N_6530,N_530,N_3519);
or U6531 (N_6531,N_1392,N_3890);
nor U6532 (N_6532,N_555,N_4326);
or U6533 (N_6533,N_716,N_108);
or U6534 (N_6534,N_842,N_2631);
or U6535 (N_6535,N_2198,N_839);
nand U6536 (N_6536,N_1809,N_2072);
nand U6537 (N_6537,N_2294,N_1534);
xor U6538 (N_6538,N_2572,N_880);
xor U6539 (N_6539,N_3977,N_4675);
nand U6540 (N_6540,N_3680,N_3028);
or U6541 (N_6541,N_751,N_287);
or U6542 (N_6542,N_1142,N_3459);
nand U6543 (N_6543,N_1873,N_2246);
and U6544 (N_6544,N_1802,N_508);
nor U6545 (N_6545,N_3093,N_21);
or U6546 (N_6546,N_3395,N_3266);
and U6547 (N_6547,N_4730,N_3457);
and U6548 (N_6548,N_4334,N_3392);
nor U6549 (N_6549,N_1118,N_2716);
nand U6550 (N_6550,N_248,N_2588);
xnor U6551 (N_6551,N_691,N_2858);
or U6552 (N_6552,N_1467,N_4610);
or U6553 (N_6553,N_4404,N_4330);
nor U6554 (N_6554,N_1576,N_4916);
and U6555 (N_6555,N_1066,N_4983);
nand U6556 (N_6556,N_1563,N_4353);
or U6557 (N_6557,N_743,N_2913);
and U6558 (N_6558,N_1822,N_4923);
nor U6559 (N_6559,N_1730,N_3711);
or U6560 (N_6560,N_3961,N_4115);
xor U6561 (N_6561,N_3492,N_2980);
and U6562 (N_6562,N_4280,N_2864);
nor U6563 (N_6563,N_1289,N_144);
nand U6564 (N_6564,N_203,N_2004);
xor U6565 (N_6565,N_4156,N_2304);
and U6566 (N_6566,N_2752,N_4277);
xor U6567 (N_6567,N_4478,N_3953);
nor U6568 (N_6568,N_2205,N_1474);
and U6569 (N_6569,N_494,N_1568);
nand U6570 (N_6570,N_2532,N_3752);
nand U6571 (N_6571,N_4727,N_2193);
xnor U6572 (N_6572,N_2610,N_4714);
and U6573 (N_6573,N_3497,N_4960);
and U6574 (N_6574,N_1955,N_3073);
xnor U6575 (N_6575,N_2519,N_1518);
and U6576 (N_6576,N_967,N_4695);
xor U6577 (N_6577,N_965,N_1939);
xor U6578 (N_6578,N_484,N_4748);
nand U6579 (N_6579,N_581,N_3529);
xor U6580 (N_6580,N_3197,N_4548);
or U6581 (N_6581,N_4082,N_1767);
xnor U6582 (N_6582,N_1326,N_4320);
nor U6583 (N_6583,N_4702,N_1023);
xor U6584 (N_6584,N_1381,N_4844);
or U6585 (N_6585,N_3296,N_145);
nor U6586 (N_6586,N_327,N_3713);
xor U6587 (N_6587,N_3957,N_2714);
and U6588 (N_6588,N_2301,N_3024);
nand U6589 (N_6589,N_1072,N_2042);
and U6590 (N_6590,N_3191,N_638);
nand U6591 (N_6591,N_3730,N_1293);
nand U6592 (N_6592,N_2841,N_42);
nand U6593 (N_6593,N_1761,N_587);
xor U6594 (N_6594,N_2050,N_3847);
nor U6595 (N_6595,N_4356,N_3005);
and U6596 (N_6596,N_1457,N_1112);
nor U6597 (N_6597,N_2527,N_979);
xnor U6598 (N_6598,N_2071,N_617);
nor U6599 (N_6599,N_4651,N_1836);
and U6600 (N_6600,N_4998,N_2612);
xor U6601 (N_6601,N_4066,N_4349);
xor U6602 (N_6602,N_2706,N_121);
nor U6603 (N_6603,N_514,N_188);
nand U6604 (N_6604,N_606,N_3369);
or U6605 (N_6605,N_2616,N_4014);
xor U6606 (N_6606,N_515,N_3273);
or U6607 (N_6607,N_3198,N_1155);
xnor U6608 (N_6608,N_615,N_3627);
nand U6609 (N_6609,N_4918,N_3863);
nor U6610 (N_6610,N_2434,N_1915);
nor U6611 (N_6611,N_1573,N_1349);
or U6612 (N_6612,N_1558,N_1127);
or U6613 (N_6613,N_2893,N_2503);
or U6614 (N_6614,N_4671,N_159);
nand U6615 (N_6615,N_1258,N_3588);
and U6616 (N_6616,N_2285,N_4071);
nor U6617 (N_6617,N_664,N_475);
or U6618 (N_6618,N_2686,N_3007);
and U6619 (N_6619,N_1971,N_3653);
or U6620 (N_6620,N_2440,N_856);
nand U6621 (N_6621,N_1620,N_235);
xnor U6622 (N_6622,N_2579,N_2035);
xor U6623 (N_6623,N_4310,N_3456);
nor U6624 (N_6624,N_1296,N_1583);
nand U6625 (N_6625,N_2687,N_4230);
nand U6626 (N_6626,N_1062,N_2605);
and U6627 (N_6627,N_4177,N_99);
xnor U6628 (N_6628,N_2412,N_3490);
nor U6629 (N_6629,N_2146,N_3000);
xor U6630 (N_6630,N_2015,N_2636);
xor U6631 (N_6631,N_2443,N_935);
or U6632 (N_6632,N_903,N_2313);
nand U6633 (N_6633,N_1787,N_3097);
nor U6634 (N_6634,N_4535,N_567);
and U6635 (N_6635,N_3795,N_4112);
xor U6636 (N_6636,N_4962,N_2917);
nor U6637 (N_6637,N_1740,N_3748);
xor U6638 (N_6638,N_4103,N_3092);
nor U6639 (N_6639,N_4664,N_4577);
xnor U6640 (N_6640,N_1605,N_4259);
nand U6641 (N_6641,N_3072,N_278);
or U6642 (N_6642,N_1760,N_4045);
and U6643 (N_6643,N_945,N_4444);
nor U6644 (N_6644,N_3762,N_3117);
or U6645 (N_6645,N_3637,N_4658);
nand U6646 (N_6646,N_230,N_3330);
xor U6647 (N_6647,N_3329,N_2865);
nor U6648 (N_6648,N_3660,N_2049);
nand U6649 (N_6649,N_4729,N_2661);
and U6650 (N_6650,N_3301,N_336);
or U6651 (N_6651,N_4572,N_3114);
and U6652 (N_6652,N_371,N_2347);
nor U6653 (N_6653,N_2375,N_2573);
or U6654 (N_6654,N_1279,N_3950);
nor U6655 (N_6655,N_1351,N_1754);
or U6656 (N_6656,N_1429,N_4291);
nand U6657 (N_6657,N_2928,N_841);
and U6658 (N_6658,N_2123,N_627);
nand U6659 (N_6659,N_3244,N_784);
nand U6660 (N_6660,N_985,N_2762);
xor U6661 (N_6661,N_1614,N_4568);
or U6662 (N_6662,N_2249,N_1779);
or U6663 (N_6663,N_470,N_4369);
nand U6664 (N_6664,N_3706,N_2848);
or U6665 (N_6665,N_2376,N_390);
nor U6666 (N_6666,N_2698,N_2141);
or U6667 (N_6667,N_2524,N_3933);
or U6668 (N_6668,N_1924,N_66);
or U6669 (N_6669,N_4662,N_4324);
and U6670 (N_6670,N_2853,N_232);
or U6671 (N_6671,N_239,N_1);
xnor U6672 (N_6672,N_4546,N_4870);
or U6673 (N_6673,N_539,N_111);
nor U6674 (N_6674,N_2812,N_3952);
nand U6675 (N_6675,N_2931,N_4355);
and U6676 (N_6676,N_832,N_152);
and U6677 (N_6677,N_4952,N_3494);
and U6678 (N_6678,N_3502,N_4977);
nor U6679 (N_6679,N_2933,N_64);
or U6680 (N_6680,N_3702,N_2293);
nor U6681 (N_6681,N_1812,N_2279);
or U6682 (N_6682,N_3942,N_3941);
nor U6683 (N_6683,N_2223,N_1601);
or U6684 (N_6684,N_2797,N_4040);
and U6685 (N_6685,N_4699,N_4598);
and U6686 (N_6686,N_3308,N_1966);
or U6687 (N_6687,N_3433,N_1539);
nand U6688 (N_6688,N_3292,N_1038);
or U6689 (N_6689,N_3676,N_234);
or U6690 (N_6690,N_2934,N_2655);
or U6691 (N_6691,N_1240,N_365);
nor U6692 (N_6692,N_4698,N_2101);
nand U6693 (N_6693,N_3299,N_2578);
and U6694 (N_6694,N_4116,N_2648);
and U6695 (N_6695,N_4625,N_8);
and U6696 (N_6696,N_4390,N_959);
or U6697 (N_6697,N_540,N_3954);
xor U6698 (N_6698,N_994,N_3774);
and U6699 (N_6699,N_93,N_1602);
or U6700 (N_6700,N_202,N_733);
xnor U6701 (N_6701,N_3306,N_2433);
nand U6702 (N_6702,N_4217,N_4603);
xor U6703 (N_6703,N_1710,N_3332);
or U6704 (N_6704,N_1272,N_1419);
and U6705 (N_6705,N_243,N_604);
xor U6706 (N_6706,N_4640,N_2982);
nand U6707 (N_6707,N_516,N_4015);
xor U6708 (N_6708,N_16,N_807);
nor U6709 (N_6709,N_1401,N_1045);
and U6710 (N_6710,N_2802,N_1688);
xor U6711 (N_6711,N_1466,N_723);
nand U6712 (N_6712,N_4367,N_3030);
xnor U6713 (N_6713,N_1439,N_3647);
or U6714 (N_6714,N_4412,N_1503);
and U6715 (N_6715,N_4995,N_4350);
and U6716 (N_6716,N_304,N_3167);
nor U6717 (N_6717,N_3101,N_3176);
or U6718 (N_6718,N_2278,N_2705);
or U6719 (N_6719,N_4777,N_4111);
xor U6720 (N_6720,N_2818,N_78);
or U6721 (N_6721,N_1058,N_1367);
xnor U6722 (N_6722,N_4296,N_2694);
xnor U6723 (N_6723,N_76,N_2624);
or U6724 (N_6724,N_1025,N_4785);
nor U6725 (N_6725,N_2956,N_2171);
nand U6726 (N_6726,N_2160,N_276);
nor U6727 (N_6727,N_709,N_3360);
or U6728 (N_6728,N_3145,N_4485);
and U6729 (N_6729,N_797,N_4718);
or U6730 (N_6730,N_32,N_2622);
or U6731 (N_6731,N_3908,N_340);
and U6732 (N_6732,N_2084,N_2404);
and U6733 (N_6733,N_4848,N_653);
xnor U6734 (N_6734,N_4129,N_3641);
nor U6735 (N_6735,N_4274,N_3442);
xor U6736 (N_6736,N_4368,N_236);
xnor U6737 (N_6737,N_820,N_2240);
nor U6738 (N_6738,N_3064,N_1281);
nor U6739 (N_6739,N_2334,N_4215);
or U6740 (N_6740,N_2734,N_2921);
or U6741 (N_6741,N_1191,N_2336);
xor U6742 (N_6742,N_3539,N_3918);
or U6743 (N_6743,N_2040,N_3673);
or U6744 (N_6744,N_2461,N_3987);
nor U6745 (N_6745,N_1910,N_4743);
nor U6746 (N_6746,N_3872,N_3959);
or U6747 (N_6747,N_939,N_4956);
and U6748 (N_6748,N_3733,N_2063);
nor U6749 (N_6749,N_3254,N_1414);
nand U6750 (N_6750,N_3632,N_4173);
and U6751 (N_6751,N_2154,N_1925);
nand U6752 (N_6752,N_4391,N_1838);
and U6753 (N_6753,N_1328,N_853);
or U6754 (N_6754,N_4644,N_622);
or U6755 (N_6755,N_707,N_1640);
xor U6756 (N_6756,N_2019,N_425);
nand U6757 (N_6757,N_2349,N_3892);
nor U6758 (N_6758,N_3091,N_4481);
or U6759 (N_6759,N_58,N_2621);
and U6760 (N_6760,N_2408,N_3800);
or U6761 (N_6761,N_2230,N_1963);
nand U6762 (N_6762,N_1119,N_2611);
nor U6763 (N_6763,N_4528,N_2730);
or U6764 (N_6764,N_95,N_3410);
nor U6765 (N_6765,N_688,N_1776);
nor U6766 (N_6766,N_110,N_472);
xnor U6767 (N_6767,N_4278,N_2867);
and U6768 (N_6768,N_637,N_4222);
or U6769 (N_6769,N_4136,N_2936);
and U6770 (N_6770,N_2878,N_1543);
nand U6771 (N_6771,N_2325,N_3347);
nor U6772 (N_6772,N_57,N_181);
nor U6773 (N_6773,N_705,N_184);
xnor U6774 (N_6774,N_1722,N_2261);
nor U6775 (N_6775,N_2680,N_43);
and U6776 (N_6776,N_565,N_3796);
xor U6777 (N_6777,N_4682,N_2290);
nand U6778 (N_6778,N_4284,N_1284);
nor U6779 (N_6779,N_2986,N_3383);
xnor U6780 (N_6780,N_1080,N_3297);
xor U6781 (N_6781,N_172,N_1358);
nor U6782 (N_6782,N_4029,N_2671);
xor U6783 (N_6783,N_4041,N_803);
xnor U6784 (N_6784,N_4713,N_4127);
nor U6785 (N_6785,N_4343,N_2515);
and U6786 (N_6786,N_208,N_1083);
or U6787 (N_6787,N_2212,N_3304);
xnor U6788 (N_6788,N_4569,N_3140);
xor U6789 (N_6789,N_3548,N_4493);
xnor U6790 (N_6790,N_1871,N_3837);
nor U6791 (N_6791,N_1791,N_3816);
nand U6792 (N_6792,N_4162,N_4058);
nand U6793 (N_6793,N_460,N_4932);
nand U6794 (N_6794,N_1588,N_3742);
nand U6795 (N_6795,N_3599,N_2276);
and U6796 (N_6796,N_2231,N_596);
nand U6797 (N_6797,N_4964,N_4038);
and U6798 (N_6798,N_2243,N_1643);
nand U6799 (N_6799,N_4885,N_3146);
or U6800 (N_6800,N_3782,N_3261);
and U6801 (N_6801,N_4552,N_3051);
and U6802 (N_6802,N_2513,N_785);
nand U6803 (N_6803,N_2388,N_3926);
or U6804 (N_6804,N_1013,N_3075);
nand U6805 (N_6805,N_2139,N_3399);
xor U6806 (N_6806,N_3363,N_23);
nor U6807 (N_6807,N_1425,N_3186);
nor U6808 (N_6808,N_3006,N_395);
nor U6809 (N_6809,N_2437,N_473);
xor U6810 (N_6810,N_1890,N_3756);
nand U6811 (N_6811,N_833,N_915);
or U6812 (N_6812,N_3813,N_3879);
xor U6813 (N_6813,N_224,N_1393);
xnor U6814 (N_6814,N_4584,N_569);
xor U6815 (N_6815,N_3111,N_2358);
or U6816 (N_6816,N_223,N_1743);
or U6817 (N_6817,N_162,N_3515);
and U6818 (N_6818,N_2425,N_1097);
or U6819 (N_6819,N_370,N_727);
and U6820 (N_6820,N_2157,N_3922);
nand U6821 (N_6821,N_529,N_164);
nor U6822 (N_6822,N_3096,N_2183);
xor U6823 (N_6823,N_1265,N_548);
nor U6824 (N_6824,N_2352,N_3927);
nor U6825 (N_6825,N_190,N_2150);
xnor U6826 (N_6826,N_3820,N_3338);
xor U6827 (N_6827,N_2456,N_3060);
nand U6828 (N_6828,N_618,N_2463);
and U6829 (N_6829,N_2912,N_3778);
nor U6830 (N_6830,N_1622,N_6);
xnor U6831 (N_6831,N_4530,N_1132);
and U6832 (N_6832,N_4618,N_2774);
nor U6833 (N_6833,N_827,N_1752);
nor U6834 (N_6834,N_2151,N_4824);
and U6835 (N_6835,N_1134,N_1386);
nand U6836 (N_6836,N_1333,N_1342);
xnor U6837 (N_6837,N_4450,N_3965);
xnor U6838 (N_6838,N_3996,N_1014);
xnor U6839 (N_6839,N_103,N_4048);
or U6840 (N_6840,N_231,N_4297);
and U6841 (N_6841,N_2499,N_4153);
and U6842 (N_6842,N_919,N_4856);
xnor U6843 (N_6843,N_1183,N_1269);
xor U6844 (N_6844,N_4814,N_1948);
nand U6845 (N_6845,N_578,N_1607);
xor U6846 (N_6846,N_2836,N_4448);
nand U6847 (N_6847,N_987,N_4055);
and U6848 (N_6848,N_2345,N_4030);
or U6849 (N_6849,N_770,N_3142);
or U6850 (N_6850,N_4194,N_1189);
nand U6851 (N_6851,N_708,N_4957);
nor U6852 (N_6852,N_3245,N_3963);
nor U6853 (N_6853,N_764,N_2983);
nor U6854 (N_6854,N_387,N_741);
xnor U6855 (N_6855,N_4035,N_409);
nand U6856 (N_6856,N_4265,N_3946);
and U6857 (N_6857,N_4757,N_183);
and U6858 (N_6858,N_4839,N_1217);
or U6859 (N_6859,N_2147,N_3449);
or U6860 (N_6860,N_914,N_1651);
or U6861 (N_6861,N_2442,N_1361);
xnor U6862 (N_6862,N_2053,N_1953);
or U6863 (N_6863,N_1691,N_2718);
nor U6864 (N_6864,N_1587,N_2682);
or U6865 (N_6865,N_2032,N_2394);
and U6866 (N_6866,N_4313,N_1613);
xor U6867 (N_6867,N_4811,N_1747);
and U6868 (N_6868,N_4166,N_67);
nand U6869 (N_6869,N_4372,N_3171);
and U6870 (N_6870,N_2441,N_4710);
and U6871 (N_6871,N_4402,N_1274);
nor U6872 (N_6872,N_1810,N_1892);
xor U6873 (N_6873,N_642,N_2001);
or U6874 (N_6874,N_3355,N_2194);
and U6875 (N_6875,N_2562,N_4017);
and U6876 (N_6876,N_4097,N_652);
xor U6877 (N_6877,N_2453,N_2077);
and U6878 (N_6878,N_2988,N_376);
nor U6879 (N_6879,N_1666,N_131);
nand U6880 (N_6880,N_2854,N_3620);
xnor U6881 (N_6881,N_225,N_4158);
xor U6882 (N_6882,N_4147,N_1950);
nand U6883 (N_6883,N_4475,N_3830);
xor U6884 (N_6884,N_2969,N_4540);
nand U6885 (N_6885,N_1513,N_3107);
and U6886 (N_6886,N_1653,N_4734);
nor U6887 (N_6887,N_2665,N_1682);
and U6888 (N_6888,N_378,N_216);
or U6889 (N_6889,N_4897,N_3016);
or U6890 (N_6890,N_1865,N_4867);
xor U6891 (N_6891,N_963,N_636);
or U6892 (N_6892,N_53,N_4042);
nand U6893 (N_6893,N_1999,N_4830);
xnor U6894 (N_6894,N_1557,N_4982);
nor U6895 (N_6895,N_3200,N_4606);
xor U6896 (N_6896,N_4196,N_671);
nand U6897 (N_6897,N_2340,N_3867);
or U6898 (N_6898,N_4901,N_4016);
xnor U6899 (N_6899,N_3119,N_4706);
and U6900 (N_6900,N_4853,N_1935);
xor U6901 (N_6901,N_1222,N_4608);
xor U6902 (N_6902,N_930,N_864);
and U6903 (N_6903,N_1070,N_448);
and U6904 (N_6904,N_2876,N_2145);
nand U6905 (N_6905,N_1907,N_4229);
or U6906 (N_6906,N_2184,N_3510);
nand U6907 (N_6907,N_1395,N_2043);
nor U6908 (N_6908,N_3556,N_423);
xnor U6909 (N_6909,N_2010,N_3061);
and U6910 (N_6910,N_3341,N_1128);
nand U6911 (N_6911,N_4971,N_4816);
or U6912 (N_6912,N_3899,N_4026);
xnor U6913 (N_6913,N_1504,N_4515);
and U6914 (N_6914,N_3480,N_3013);
xor U6915 (N_6915,N_1391,N_2113);
and U6916 (N_6916,N_3106,N_4223);
and U6917 (N_6917,N_3518,N_830);
or U6918 (N_6918,N_4579,N_1636);
nand U6919 (N_6919,N_3705,N_4728);
and U6920 (N_6920,N_254,N_3201);
xnor U6921 (N_6921,N_2038,N_918);
xnor U6922 (N_6922,N_2843,N_4303);
nand U6923 (N_6923,N_4891,N_1817);
or U6924 (N_6924,N_826,N_4211);
nand U6925 (N_6925,N_2607,N_177);
nor U6926 (N_6926,N_4542,N_1016);
or U6927 (N_6927,N_2262,N_2949);
or U6928 (N_6928,N_1091,N_3088);
nand U6929 (N_6929,N_1194,N_4282);
or U6930 (N_6930,N_681,N_1933);
and U6931 (N_6931,N_2286,N_4075);
nand U6932 (N_6932,N_321,N_194);
nor U6933 (N_6933,N_2558,N_1239);
nor U6934 (N_6934,N_4266,N_2364);
nand U6935 (N_6935,N_2710,N_4316);
nor U6936 (N_6936,N_3882,N_2343);
or U6937 (N_6937,N_2828,N_2650);
nor U6938 (N_6938,N_1755,N_3604);
nor U6939 (N_6939,N_38,N_2548);
nor U6940 (N_6940,N_4863,N_1317);
or U6941 (N_6941,N_2529,N_4969);
and U6942 (N_6942,N_1762,N_1512);
or U6943 (N_6943,N_1242,N_3045);
and U6944 (N_6944,N_3121,N_3098);
and U6945 (N_6945,N_731,N_3619);
or U6946 (N_6946,N_3818,N_3522);
or U6947 (N_6947,N_4566,N_1616);
and U6948 (N_6948,N_3929,N_676);
nand U6949 (N_6949,N_362,N_4672);
nand U6950 (N_6950,N_3157,N_4047);
xor U6951 (N_6951,N_613,N_1389);
nor U6952 (N_6952,N_4435,N_1547);
nor U6953 (N_6953,N_4212,N_3854);
nand U6954 (N_6954,N_549,N_408);
or U6955 (N_6955,N_4630,N_1719);
and U6956 (N_6956,N_199,N_265);
nand U6957 (N_6957,N_848,N_3135);
and U6958 (N_6958,N_2676,N_4376);
and U6959 (N_6959,N_4126,N_3764);
and U6960 (N_6960,N_1427,N_4143);
and U6961 (N_6961,N_4654,N_2267);
xnor U6962 (N_6962,N_1312,N_4917);
xnor U6963 (N_6963,N_24,N_3432);
nand U6964 (N_6964,N_3897,N_4859);
nand U6965 (N_6965,N_3263,N_1728);
nand U6966 (N_6966,N_2052,N_3643);
nor U6967 (N_6967,N_4851,N_1348);
and U6968 (N_6968,N_659,N_1753);
nor U6969 (N_6969,N_1069,N_392);
or U6970 (N_6970,N_2765,N_3228);
or U6971 (N_6971,N_790,N_3303);
and U6972 (N_6972,N_1548,N_2264);
xor U6973 (N_6973,N_4782,N_697);
or U6974 (N_6974,N_2814,N_2776);
nor U6975 (N_6975,N_1115,N_1211);
nand U6976 (N_6976,N_4432,N_1757);
nor U6977 (N_6977,N_1593,N_305);
or U6978 (N_6978,N_3531,N_3902);
or U6979 (N_6979,N_600,N_1408);
nand U6980 (N_6980,N_3272,N_4541);
xnor U6981 (N_6981,N_3549,N_3860);
nor U6982 (N_6982,N_4307,N_4337);
nor U6983 (N_6983,N_2107,N_1343);
or U6984 (N_6984,N_1672,N_3630);
xor U6985 (N_6985,N_1785,N_781);
or U6986 (N_6986,N_1262,N_4553);
nand U6987 (N_6987,N_1412,N_4686);
xor U6988 (N_6988,N_349,N_2534);
nand U6989 (N_6989,N_603,N_4184);
xor U6990 (N_6990,N_86,N_3851);
nand U6991 (N_6991,N_1250,N_4484);
nor U6992 (N_6992,N_5,N_1641);
or U6993 (N_6993,N_2586,N_1404);
xor U6994 (N_6994,N_3257,N_97);
nand U6995 (N_6995,N_3235,N_1170);
xnor U6996 (N_6996,N_4057,N_2960);
or U6997 (N_6997,N_1241,N_428);
xor U6998 (N_6998,N_3861,N_3777);
xnor U6999 (N_6999,N_3102,N_4915);
nor U7000 (N_7000,N_1411,N_2405);
nor U7001 (N_7001,N_4370,N_1198);
xnor U7002 (N_7002,N_4174,N_4335);
and U7003 (N_7003,N_2162,N_1402);
nor U7004 (N_7004,N_2963,N_2626);
nand U7005 (N_7005,N_668,N_1443);
nand U7006 (N_7006,N_2156,N_3765);
nor U7007 (N_7007,N_3986,N_2733);
or U7008 (N_7008,N_3326,N_1140);
nand U7009 (N_7009,N_4062,N_1500);
and U7010 (N_7010,N_2639,N_3068);
or U7011 (N_7011,N_4888,N_1652);
nor U7012 (N_7012,N_4092,N_3749);
nor U7013 (N_7013,N_1245,N_3577);
xnor U7014 (N_7014,N_431,N_4593);
and U7015 (N_7015,N_1839,N_4470);
xnor U7016 (N_7016,N_3166,N_2003);
and U7017 (N_7017,N_4522,N_4519);
and U7018 (N_7018,N_2723,N_2416);
nor U7019 (N_7019,N_2460,N_1163);
and U7020 (N_7020,N_178,N_3936);
and U7021 (N_7021,N_1086,N_4788);
nand U7022 (N_7022,N_1009,N_116);
nand U7023 (N_7023,N_1724,N_4231);
and U7024 (N_7024,N_3562,N_4506);
xor U7025 (N_7025,N_4384,N_2715);
and U7026 (N_7026,N_4902,N_2076);
nand U7027 (N_7027,N_2821,N_2333);
nand U7028 (N_7028,N_3307,N_4929);
and U7029 (N_7029,N_3512,N_4975);
and U7030 (N_7030,N_4906,N_244);
and U7031 (N_7031,N_3187,N_3843);
nor U7032 (N_7032,N_3172,N_3223);
nor U7033 (N_7033,N_4643,N_1234);
nor U7034 (N_7034,N_4345,N_14);
or U7035 (N_7035,N_2791,N_523);
or U7036 (N_7036,N_1623,N_561);
nor U7037 (N_7037,N_4873,N_2609);
nor U7038 (N_7038,N_4622,N_3340);
and U7039 (N_7039,N_2271,N_4965);
xnor U7040 (N_7040,N_2495,N_175);
xnor U7041 (N_7041,N_3514,N_2978);
xor U7042 (N_7042,N_4154,N_150);
and U7043 (N_7043,N_120,N_2227);
nor U7044 (N_7044,N_3046,N_4503);
nor U7045 (N_7045,N_4948,N_2044);
xnor U7046 (N_7046,N_1958,N_2559);
nor U7047 (N_7047,N_630,N_4430);
xor U7048 (N_7048,N_890,N_1922);
nand U7049 (N_7049,N_319,N_4913);
nand U7050 (N_7050,N_1968,N_2239);
and U7051 (N_7051,N_2143,N_4295);
and U7052 (N_7052,N_4924,N_699);
and U7053 (N_7053,N_1671,N_1944);
nor U7054 (N_7054,N_4738,N_3344);
xor U7055 (N_7055,N_2974,N_2466);
nand U7056 (N_7056,N_3616,N_2106);
and U7057 (N_7057,N_1088,N_2235);
and U7058 (N_7058,N_2896,N_481);
or U7059 (N_7059,N_4739,N_2915);
xnor U7060 (N_7060,N_1219,N_3989);
xor U7061 (N_7061,N_2396,N_171);
xnor U7062 (N_7062,N_1149,N_4068);
xnor U7063 (N_7063,N_20,N_2561);
nor U7064 (N_7064,N_1230,N_2417);
or U7065 (N_7065,N_1050,N_2473);
xor U7066 (N_7066,N_317,N_825);
or U7067 (N_7067,N_3368,N_3591);
and U7068 (N_7068,N_4262,N_1599);
xnor U7069 (N_7069,N_3839,N_754);
nor U7070 (N_7070,N_4004,N_2091);
or U7071 (N_7071,N_1604,N_4283);
or U7072 (N_7072,N_2786,N_1449);
or U7073 (N_7073,N_421,N_2134);
or U7074 (N_7074,N_2645,N_3469);
nor U7075 (N_7075,N_2124,N_117);
xor U7076 (N_7076,N_398,N_2321);
xnor U7077 (N_7077,N_1818,N_4943);
and U7078 (N_7078,N_459,N_4800);
nor U7079 (N_7079,N_1448,N_3503);
nand U7080 (N_7080,N_675,N_2897);
xor U7081 (N_7081,N_3126,N_656);
and U7082 (N_7082,N_4246,N_711);
nor U7083 (N_7083,N_4449,N_4701);
nor U7084 (N_7084,N_94,N_201);
nor U7085 (N_7085,N_2484,N_2615);
nor U7086 (N_7086,N_1893,N_1405);
and U7087 (N_7087,N_2036,N_3642);
xnor U7088 (N_7088,N_1926,N_1845);
nand U7089 (N_7089,N_1283,N_4394);
and U7090 (N_7090,N_192,N_2384);
nor U7091 (N_7091,N_2830,N_938);
or U7092 (N_7092,N_2794,N_1644);
or U7093 (N_7093,N_402,N_11);
nand U7094 (N_7094,N_3175,N_1049);
and U7095 (N_7095,N_871,N_2555);
nand U7096 (N_7096,N_1796,N_2961);
and U7097 (N_7097,N_2780,N_1331);
xor U7098 (N_7098,N_3352,N_4650);
nand U7099 (N_7099,N_2022,N_1770);
or U7100 (N_7100,N_1947,N_4091);
or U7101 (N_7101,N_1694,N_451);
xnor U7102 (N_7102,N_4480,N_2342);
and U7103 (N_7103,N_645,N_2875);
nor U7104 (N_7104,N_4400,N_2029);
nor U7105 (N_7105,N_81,N_1621);
nand U7106 (N_7106,N_222,N_2662);
nor U7107 (N_7107,N_4086,N_1059);
xnor U7108 (N_7108,N_2522,N_2950);
or U7109 (N_7109,N_2879,N_2097);
and U7110 (N_7110,N_660,N_4990);
or U7111 (N_7111,N_3979,N_4188);
nand U7112 (N_7112,N_1282,N_551);
nand U7113 (N_7113,N_127,N_1973);
or U7114 (N_7114,N_134,N_45);
and U7115 (N_7115,N_4441,N_3634);
nor U7116 (N_7116,N_2965,N_1017);
nor U7117 (N_7117,N_4765,N_1670);
nor U7118 (N_7118,N_4359,N_3380);
nor U7119 (N_7119,N_3452,N_2385);
or U7120 (N_7120,N_3969,N_889);
and U7121 (N_7121,N_2324,N_3975);
nand U7122 (N_7122,N_3537,N_3271);
nand U7123 (N_7123,N_3917,N_418);
and U7124 (N_7124,N_1486,N_4180);
xnor U7125 (N_7125,N_443,N_2721);
nand U7126 (N_7126,N_4545,N_1896);
nor U7127 (N_7127,N_759,N_1338);
nor U7128 (N_7128,N_51,N_616);
nand U7129 (N_7129,N_2745,N_1901);
nor U7130 (N_7130,N_917,N_4806);
or U7131 (N_7131,N_3488,N_3210);
nand U7132 (N_7132,N_1177,N_4562);
nand U7133 (N_7133,N_3614,N_2132);
or U7134 (N_7134,N_1390,N_2487);
and U7135 (N_7135,N_2452,N_498);
nand U7136 (N_7136,N_2435,N_635);
xor U7137 (N_7137,N_3805,N_146);
nand U7138 (N_7138,N_762,N_628);
xnor U7139 (N_7139,N_3798,N_3507);
and U7140 (N_7140,N_657,N_2939);
xor U7141 (N_7141,N_4890,N_3004);
and U7142 (N_7142,N_82,N_4570);
and U7143 (N_7143,N_2295,N_602);
nand U7144 (N_7144,N_4878,N_1826);
or U7145 (N_7145,N_3050,N_1847);
and U7146 (N_7146,N_644,N_1440);
xor U7147 (N_7147,N_663,N_3104);
xnor U7148 (N_7148,N_632,N_901);
and U7149 (N_7149,N_4076,N_1685);
nand U7150 (N_7150,N_2054,N_3654);
xnor U7151 (N_7151,N_1982,N_1034);
xor U7152 (N_7152,N_814,N_3677);
and U7153 (N_7153,N_1980,N_1840);
or U7154 (N_7154,N_782,N_2769);
and U7155 (N_7155,N_1117,N_2173);
or U7156 (N_7156,N_2971,N_745);
nor U7157 (N_7157,N_3971,N_758);
and U7158 (N_7158,N_1360,N_1851);
nor U7159 (N_7159,N_4331,N_2653);
and U7160 (N_7160,N_1365,N_75);
nand U7161 (N_7161,N_2411,N_3026);
xnor U7162 (N_7162,N_1554,N_1600);
and U7163 (N_7163,N_736,N_984);
nor U7164 (N_7164,N_520,N_4241);
or U7165 (N_7165,N_491,N_2782);
or U7166 (N_7166,N_433,N_2771);
or U7167 (N_7167,N_2182,N_3448);
and U7168 (N_7168,N_780,N_4793);
xnor U7169 (N_7169,N_3116,N_1090);
or U7170 (N_7170,N_3960,N_3221);
nand U7171 (N_7171,N_4547,N_737);
or U7172 (N_7172,N_1368,N_1523);
and U7173 (N_7173,N_2512,N_2674);
and U7174 (N_7174,N_3520,N_1477);
nand U7175 (N_7175,N_1178,N_2750);
xor U7176 (N_7176,N_4298,N_2644);
xnor U7177 (N_7177,N_2020,N_1766);
nand U7178 (N_7178,N_2595,N_2895);
nand U7179 (N_7179,N_267,N_3413);
nor U7180 (N_7180,N_3275,N_3431);
or U7181 (N_7181,N_1699,N_1051);
and U7182 (N_7182,N_3608,N_3288);
xnor U7183 (N_7183,N_4138,N_1782);
and U7184 (N_7184,N_4726,N_654);
xnor U7185 (N_7185,N_992,N_2629);
or U7186 (N_7186,N_3527,N_3891);
nand U7187 (N_7187,N_687,N_2748);
nand U7188 (N_7188,N_4938,N_379);
and U7189 (N_7189,N_2531,N_1700);
and U7190 (N_7190,N_1758,N_3217);
xor U7191 (N_7191,N_734,N_2944);
nor U7192 (N_7192,N_3379,N_2637);
and U7193 (N_7193,N_4245,N_3681);
xnor U7194 (N_7194,N_1456,N_1253);
or U7195 (N_7195,N_4724,N_4722);
nand U7196 (N_7196,N_4945,N_3881);
or U7197 (N_7197,N_3856,N_3804);
nor U7198 (N_7198,N_2722,N_1756);
xnor U7199 (N_7199,N_2932,N_2514);
nand U7200 (N_7200,N_3476,N_366);
and U7201 (N_7201,N_4168,N_2628);
nor U7202 (N_7202,N_1436,N_4471);
nand U7203 (N_7203,N_3807,N_2431);
and U7204 (N_7204,N_296,N_4152);
and U7205 (N_7205,N_916,N_3727);
xor U7206 (N_7206,N_2268,N_2990);
or U7207 (N_7207,N_2997,N_3722);
xor U7208 (N_7208,N_2929,N_570);
and U7209 (N_7209,N_3414,N_3792);
xor U7210 (N_7210,N_2696,N_753);
nand U7211 (N_7211,N_3606,N_580);
xnor U7212 (N_7212,N_989,N_3896);
nor U7213 (N_7213,N_639,N_4371);
nand U7214 (N_7214,N_264,N_1708);
or U7215 (N_7215,N_680,N_2423);
nand U7216 (N_7216,N_4767,N_4752);
xor U7217 (N_7217,N_335,N_1084);
xor U7218 (N_7218,N_3182,N_3639);
or U7219 (N_7219,N_1275,N_4882);
nor U7220 (N_7220,N_1609,N_4294);
and U7221 (N_7221,N_3907,N_228);
or U7222 (N_7222,N_2490,N_4539);
or U7223 (N_7223,N_2542,N_3062);
or U7224 (N_7224,N_810,N_2767);
and U7225 (N_7225,N_3678,N_4243);
nor U7226 (N_7226,N_2593,N_3553);
xnor U7227 (N_7227,N_361,N_777);
or U7228 (N_7228,N_4383,N_1789);
nor U7229 (N_7229,N_3420,N_3021);
xnor U7230 (N_7230,N_3695,N_4760);
nor U7231 (N_7231,N_2831,N_2704);
xor U7232 (N_7232,N_1570,N_3939);
nor U7233 (N_7233,N_3684,N_4832);
xnor U7234 (N_7234,N_4955,N_4525);
or U7235 (N_7235,N_196,N_1450);
or U7236 (N_7236,N_1917,N_3724);
nor U7237 (N_7237,N_902,N_3209);
and U7238 (N_7238,N_1727,N_2743);
and U7239 (N_7239,N_1218,N_541);
and U7240 (N_7240,N_1125,N_1141);
nand U7241 (N_7241,N_4032,N_2136);
xnor U7242 (N_7242,N_2200,N_1100);
nand U7243 (N_7243,N_2945,N_2475);
and U7244 (N_7244,N_3912,N_3293);
nand U7245 (N_7245,N_4096,N_808);
nor U7246 (N_7246,N_2489,N_1863);
nand U7247 (N_7247,N_895,N_4665);
nand U7248 (N_7248,N_1180,N_1053);
xnor U7249 (N_7249,N_4011,N_2642);
xor U7250 (N_7250,N_909,N_1478);
nor U7251 (N_7251,N_649,N_4737);
or U7252 (N_7252,N_4273,N_1668);
and U7253 (N_7253,N_3683,N_2277);
nand U7254 (N_7254,N_3274,N_3645);
and U7255 (N_7255,N_1844,N_3806);
xor U7256 (N_7256,N_4247,N_2882);
or U7257 (N_7257,N_4850,N_3964);
nor U7258 (N_7258,N_153,N_2500);
nand U7259 (N_7259,N_334,N_1765);
nand U7260 (N_7260,N_210,N_3783);
or U7261 (N_7261,N_4504,N_4796);
or U7262 (N_7262,N_4537,N_966);
nand U7263 (N_7263,N_2918,N_4342);
nor U7264 (N_7264,N_4582,N_4778);
or U7265 (N_7265,N_740,N_3475);
and U7266 (N_7266,N_416,N_1400);
nand U7267 (N_7267,N_4207,N_972);
xnor U7268 (N_7268,N_2951,N_1223);
xnor U7269 (N_7269,N_1703,N_292);
xor U7270 (N_7270,N_2673,N_350);
or U7271 (N_7271,N_794,N_2161);
nor U7272 (N_7272,N_2787,N_3753);
nor U7273 (N_7273,N_511,N_2119);
xor U7274 (N_7274,N_3404,N_1202);
nand U7275 (N_7275,N_4967,N_1569);
xnor U7276 (N_7276,N_4059,N_3464);
and U7277 (N_7277,N_908,N_3612);
nor U7278 (N_7278,N_1517,N_1098);
or U7279 (N_7279,N_59,N_2979);
and U7280 (N_7280,N_4829,N_4149);
nand U7281 (N_7281,N_4985,N_2523);
nand U7282 (N_7282,N_442,N_330);
and U7283 (N_7283,N_582,N_4150);
nor U7284 (N_7284,N_2203,N_197);
nand U7285 (N_7285,N_1465,N_1406);
xnor U7286 (N_7286,N_3650,N_4364);
nand U7287 (N_7287,N_4467,N_1858);
xnor U7288 (N_7288,N_4623,N_1122);
or U7289 (N_7289,N_3524,N_1280);
xor U7290 (N_7290,N_3349,N_2919);
or U7291 (N_7291,N_3709,N_3973);
and U7292 (N_7292,N_1751,N_272);
xor U7293 (N_7293,N_68,N_49);
nor U7294 (N_7294,N_2491,N_118);
and U7295 (N_7295,N_3083,N_2885);
nand U7296 (N_7296,N_9,N_4171);
nand U7297 (N_7297,N_696,N_3285);
or U7298 (N_7298,N_1849,N_3938);
and U7299 (N_7299,N_4819,N_77);
or U7300 (N_7300,N_2367,N_28);
xnor U7301 (N_7301,N_219,N_4489);
nand U7302 (N_7302,N_3968,N_3470);
and U7303 (N_7303,N_1715,N_3314);
or U7304 (N_7304,N_610,N_2302);
xor U7305 (N_7305,N_1549,N_4336);
or U7306 (N_7306,N_2600,N_3012);
and U7307 (N_7307,N_140,N_4936);
nor U7308 (N_7308,N_650,N_4013);
nand U7309 (N_7309,N_1374,N_2024);
and U7310 (N_7310,N_273,N_2663);
or U7311 (N_7311,N_4198,N_893);
nand U7312 (N_7312,N_4438,N_3923);
nor U7313 (N_7313,N_3133,N_4003);
and U7314 (N_7314,N_2331,N_986);
nand U7315 (N_7315,N_1497,N_495);
nand U7316 (N_7316,N_4592,N_1885);
and U7317 (N_7317,N_1221,N_3594);
nand U7318 (N_7318,N_2964,N_933);
or U7319 (N_7319,N_2248,N_297);
nand U7320 (N_7320,N_1987,N_4667);
and U7321 (N_7321,N_2485,N_2259);
nor U7322 (N_7322,N_3852,N_809);
or U7323 (N_7323,N_1308,N_1692);
or U7324 (N_7324,N_87,N_281);
nor U7325 (N_7325,N_3482,N_3496);
nor U7326 (N_7326,N_3078,N_2289);
nand U7327 (N_7327,N_260,N_1596);
nor U7328 (N_7328,N_2766,N_2018);
or U7329 (N_7329,N_3423,N_3812);
nand U7330 (N_7330,N_2866,N_1047);
or U7331 (N_7331,N_3445,N_1430);
nand U7332 (N_7332,N_2702,N_4661);
nand U7333 (N_7333,N_1285,N_3265);
or U7334 (N_7334,N_3578,N_3339);
nor U7335 (N_7335,N_1806,N_2546);
and U7336 (N_7336,N_3484,N_776);
nor U7337 (N_7337,N_792,N_4854);
nand U7338 (N_7338,N_1251,N_4054);
nor U7339 (N_7339,N_843,N_2181);
xnor U7340 (N_7340,N_1135,N_4907);
nor U7341 (N_7341,N_974,N_3154);
nand U7342 (N_7342,N_2635,N_3342);
xnor U7343 (N_7343,N_2222,N_552);
nand U7344 (N_7344,N_2177,N_1073);
nor U7345 (N_7345,N_544,N_851);
or U7346 (N_7346,N_462,N_1131);
or U7347 (N_7347,N_1860,N_3105);
and U7348 (N_7348,N_4299,N_176);
xnor U7349 (N_7349,N_1772,N_3873);
nand U7350 (N_7350,N_2681,N_307);
or U7351 (N_7351,N_2129,N_1006);
nor U7352 (N_7352,N_1697,N_1278);
nor U7353 (N_7353,N_4768,N_2447);
nand U7354 (N_7354,N_2424,N_533);
nor U7355 (N_7355,N_2322,N_2634);
and U7356 (N_7356,N_380,N_1531);
nand U7357 (N_7357,N_1992,N_4366);
nand U7358 (N_7358,N_1187,N_1914);
or U7359 (N_7359,N_2296,N_1482);
and U7360 (N_7360,N_1362,N_2138);
nand U7361 (N_7361,N_3401,N_2397);
and U7362 (N_7362,N_2041,N_1927);
or U7363 (N_7363,N_3054,N_1352);
nand U7364 (N_7364,N_1759,N_369);
nor U7365 (N_7365,N_4169,N_3076);
and U7366 (N_7366,N_1496,N_4189);
nand U7367 (N_7367,N_1313,N_3190);
xnor U7368 (N_7368,N_4499,N_3685);
and U7369 (N_7369,N_1201,N_3661);
nor U7370 (N_7370,N_2112,N_4903);
nor U7371 (N_7371,N_1306,N_2209);
nand U7372 (N_7372,N_2328,N_4771);
nor U7373 (N_7373,N_3883,N_3850);
xnor U7374 (N_7374,N_3567,N_517);
or U7375 (N_7375,N_167,N_3657);
nor U7376 (N_7376,N_3356,N_1473);
and U7377 (N_7377,N_3557,N_2970);
or U7378 (N_7378,N_2389,N_2656);
or U7379 (N_7379,N_1713,N_2813);
or U7380 (N_7380,N_4594,N_3147);
nand U7381 (N_7381,N_1585,N_1021);
and U7382 (N_7382,N_2241,N_182);
nor U7383 (N_7383,N_4272,N_1805);
nor U7384 (N_7384,N_571,N_836);
nand U7385 (N_7385,N_3032,N_2772);
and U7386 (N_7386,N_3129,N_1771);
nand U7387 (N_7387,N_3447,N_1835);
nor U7388 (N_7388,N_4634,N_4084);
and U7389 (N_7389,N_3589,N_147);
xnor U7390 (N_7390,N_2539,N_3240);
or U7391 (N_7391,N_237,N_1701);
and U7392 (N_7392,N_4527,N_2315);
xor U7393 (N_7393,N_2768,N_1259);
or U7394 (N_7394,N_850,N_180);
or U7395 (N_7395,N_4257,N_3357);
or U7396 (N_7396,N_3354,N_2759);
or U7397 (N_7397,N_1878,N_4270);
nor U7398 (N_7398,N_4858,N_1509);
and U7399 (N_7399,N_4711,N_3039);
xnor U7400 (N_7400,N_3477,N_1357);
xnor U7401 (N_7401,N_1422,N_2309);
or U7402 (N_7402,N_247,N_934);
and U7403 (N_7403,N_3100,N_2357);
or U7404 (N_7404,N_1261,N_1667);
nor U7405 (N_7405,N_911,N_981);
or U7406 (N_7406,N_345,N_2062);
or U7407 (N_7407,N_3536,N_3935);
xor U7408 (N_7408,N_2115,N_249);
xor U7409 (N_7409,N_4008,N_892);
nand U7410 (N_7410,N_1637,N_4140);
and U7411 (N_7411,N_1022,N_3127);
and U7412 (N_7412,N_3440,N_2265);
and U7413 (N_7413,N_2899,N_3450);
and U7414 (N_7414,N_1214,N_3889);
or U7415 (N_7415,N_3984,N_1046);
xnor U7416 (N_7416,N_2159,N_363);
xnor U7417 (N_7417,N_4101,N_4363);
nand U7418 (N_7418,N_3622,N_3651);
nor U7419 (N_7419,N_4306,N_1029);
nand U7420 (N_7420,N_913,N_2256);
or U7421 (N_7421,N_2570,N_3771);
and U7422 (N_7422,N_4090,N_1375);
nand U7423 (N_7423,N_2565,N_3838);
or U7424 (N_7424,N_3995,N_149);
nand U7425 (N_7425,N_3237,N_3811);
xnor U7426 (N_7426,N_2387,N_4267);
xnor U7427 (N_7427,N_3473,N_732);
and U7428 (N_7428,N_4893,N_3893);
nor U7429 (N_7429,N_2625,N_3086);
and U7430 (N_7430,N_1894,N_3652);
nor U7431 (N_7431,N_866,N_2757);
xnor U7432 (N_7432,N_3095,N_1679);
nor U7433 (N_7433,N_332,N_4583);
nor U7434 (N_7434,N_1431,N_4012);
nor U7435 (N_7435,N_3611,N_1746);
xor U7436 (N_7436,N_1461,N_1077);
and U7437 (N_7437,N_2098,N_4285);
nand U7438 (N_7438,N_1248,N_1203);
and U7439 (N_7439,N_4678,N_542);
and U7440 (N_7440,N_980,N_3020);
nor U7441 (N_7441,N_3663,N_4232);
nand U7442 (N_7442,N_608,N_2281);
xnor U7443 (N_7443,N_3280,N_4790);
nand U7444 (N_7444,N_1124,N_89);
or U7445 (N_7445,N_4393,N_2488);
and U7446 (N_7446,N_4981,N_452);
and U7447 (N_7447,N_4379,N_290);
or U7448 (N_7448,N_4574,N_435);
nor U7449 (N_7449,N_2127,N_647);
or U7450 (N_7450,N_169,N_1774);
nand U7451 (N_7451,N_522,N_3690);
or U7452 (N_7452,N_3336,N_2252);
nor U7453 (N_7453,N_115,N_1902);
or U7454 (N_7454,N_2738,N_4159);
or U7455 (N_7455,N_4161,N_3174);
and U7456 (N_7456,N_667,N_1185);
nand U7457 (N_7457,N_3441,N_1931);
or U7458 (N_7458,N_1432,N_1723);
or U7459 (N_7459,N_2218,N_2204);
nand U7460 (N_7460,N_4386,N_806);
nor U7461 (N_7461,N_2142,N_1989);
nand U7462 (N_7462,N_665,N_1210);
and U7463 (N_7463,N_2339,N_3189);
or U7464 (N_7464,N_682,N_3290);
xnor U7465 (N_7465,N_4922,N_1867);
or U7466 (N_7466,N_3558,N_4125);
and U7467 (N_7467,N_1495,N_4899);
nor U7468 (N_7468,N_403,N_4203);
nand U7469 (N_7469,N_2654,N_2196);
nand U7470 (N_7470,N_1438,N_2390);
or U7471 (N_7471,N_41,N_1985);
xor U7472 (N_7472,N_948,N_2852);
and U7473 (N_7473,N_100,N_3739);
nor U7474 (N_7474,N_2998,N_4305);
xnor U7475 (N_7475,N_2711,N_3666);
nand U7476 (N_7476,N_360,N_4224);
xnor U7477 (N_7477,N_2601,N_886);
and U7478 (N_7478,N_3276,N_2330);
nor U7479 (N_7479,N_2717,N_2627);
nand U7480 (N_7480,N_3444,N_2571);
nor U7481 (N_7481,N_1065,N_2747);
nor U7482 (N_7482,N_119,N_3229);
or U7483 (N_7483,N_767,N_2167);
nor U7484 (N_7484,N_1657,N_2075);
and U7485 (N_7485,N_168,N_3566);
or U7486 (N_7486,N_528,N_1145);
and U7487 (N_7487,N_4629,N_597);
and U7488 (N_7488,N_485,N_1271);
nand U7489 (N_7489,N_584,N_1969);
nor U7490 (N_7490,N_4909,N_1868);
nand U7491 (N_7491,N_4426,N_3766);
and U7492 (N_7492,N_4208,N_4190);
xor U7493 (N_7493,N_2886,N_4483);
and U7494 (N_7494,N_2346,N_1704);
xnor U7495 (N_7495,N_4784,N_3398);
or U7496 (N_7496,N_1991,N_4604);
nor U7497 (N_7497,N_226,N_1632);
nor U7498 (N_7498,N_3693,N_1417);
xnor U7499 (N_7499,N_1608,N_1339);
or U7500 (N_7500,N_4590,N_3896);
nand U7501 (N_7501,N_4226,N_4427);
nand U7502 (N_7502,N_4133,N_3498);
nor U7503 (N_7503,N_2292,N_430);
nand U7504 (N_7504,N_4439,N_4267);
nand U7505 (N_7505,N_4171,N_3833);
and U7506 (N_7506,N_1613,N_2066);
and U7507 (N_7507,N_4933,N_2347);
and U7508 (N_7508,N_1861,N_3641);
xor U7509 (N_7509,N_3370,N_1813);
and U7510 (N_7510,N_3368,N_4499);
nor U7511 (N_7511,N_2975,N_2470);
nand U7512 (N_7512,N_4400,N_1449);
nor U7513 (N_7513,N_3440,N_4403);
and U7514 (N_7514,N_3713,N_3732);
or U7515 (N_7515,N_2765,N_472);
nand U7516 (N_7516,N_2667,N_920);
nand U7517 (N_7517,N_1087,N_3215);
or U7518 (N_7518,N_138,N_4410);
xor U7519 (N_7519,N_1433,N_785);
nand U7520 (N_7520,N_3224,N_4230);
xnor U7521 (N_7521,N_2745,N_1226);
or U7522 (N_7522,N_3166,N_4205);
and U7523 (N_7523,N_341,N_3350);
nor U7524 (N_7524,N_2874,N_2);
nor U7525 (N_7525,N_850,N_1365);
or U7526 (N_7526,N_77,N_18);
nand U7527 (N_7527,N_3287,N_2620);
and U7528 (N_7528,N_2064,N_3317);
xor U7529 (N_7529,N_2505,N_2639);
nor U7530 (N_7530,N_2330,N_3998);
or U7531 (N_7531,N_2202,N_2532);
and U7532 (N_7532,N_4797,N_3839);
nand U7533 (N_7533,N_4545,N_3772);
xor U7534 (N_7534,N_4372,N_392);
xor U7535 (N_7535,N_2221,N_3354);
xor U7536 (N_7536,N_354,N_792);
xor U7537 (N_7537,N_4215,N_1169);
xnor U7538 (N_7538,N_3058,N_1668);
nand U7539 (N_7539,N_1106,N_4100);
and U7540 (N_7540,N_3281,N_2890);
or U7541 (N_7541,N_2011,N_571);
or U7542 (N_7542,N_4539,N_4283);
or U7543 (N_7543,N_3578,N_1269);
nor U7544 (N_7544,N_1968,N_401);
or U7545 (N_7545,N_3644,N_3278);
nor U7546 (N_7546,N_317,N_758);
or U7547 (N_7547,N_1113,N_3692);
nor U7548 (N_7548,N_3144,N_2808);
nor U7549 (N_7549,N_2723,N_169);
or U7550 (N_7550,N_3068,N_3089);
xnor U7551 (N_7551,N_4260,N_1014);
nand U7552 (N_7552,N_4237,N_545);
nor U7553 (N_7553,N_649,N_2620);
xnor U7554 (N_7554,N_585,N_4513);
nor U7555 (N_7555,N_1815,N_74);
xor U7556 (N_7556,N_2597,N_489);
and U7557 (N_7557,N_781,N_4114);
xor U7558 (N_7558,N_368,N_1298);
and U7559 (N_7559,N_3368,N_3056);
nand U7560 (N_7560,N_2923,N_3165);
nor U7561 (N_7561,N_1268,N_1679);
xnor U7562 (N_7562,N_2281,N_163);
or U7563 (N_7563,N_4569,N_523);
nand U7564 (N_7564,N_2354,N_1256);
nor U7565 (N_7565,N_749,N_234);
and U7566 (N_7566,N_2855,N_2303);
nor U7567 (N_7567,N_933,N_1656);
nor U7568 (N_7568,N_537,N_130);
nor U7569 (N_7569,N_3858,N_3952);
nor U7570 (N_7570,N_1423,N_4673);
or U7571 (N_7571,N_2556,N_4109);
nand U7572 (N_7572,N_4754,N_4315);
xor U7573 (N_7573,N_707,N_2660);
or U7574 (N_7574,N_2832,N_2932);
or U7575 (N_7575,N_581,N_3098);
xor U7576 (N_7576,N_3419,N_4057);
or U7577 (N_7577,N_3896,N_1096);
and U7578 (N_7578,N_2243,N_2209);
xor U7579 (N_7579,N_1921,N_2851);
nor U7580 (N_7580,N_4093,N_1348);
nor U7581 (N_7581,N_2704,N_5);
or U7582 (N_7582,N_999,N_1808);
xor U7583 (N_7583,N_3648,N_2157);
and U7584 (N_7584,N_57,N_1973);
and U7585 (N_7585,N_4795,N_1774);
or U7586 (N_7586,N_2373,N_4617);
xnor U7587 (N_7587,N_4874,N_3107);
or U7588 (N_7588,N_3622,N_2750);
nand U7589 (N_7589,N_4586,N_3410);
xor U7590 (N_7590,N_171,N_561);
nand U7591 (N_7591,N_4538,N_2937);
nor U7592 (N_7592,N_627,N_3767);
nand U7593 (N_7593,N_3275,N_3712);
nand U7594 (N_7594,N_4124,N_4610);
xnor U7595 (N_7595,N_1270,N_605);
nor U7596 (N_7596,N_4856,N_1886);
xor U7597 (N_7597,N_786,N_2360);
and U7598 (N_7598,N_4752,N_4481);
or U7599 (N_7599,N_386,N_4759);
nor U7600 (N_7600,N_2641,N_3966);
and U7601 (N_7601,N_1883,N_2506);
nand U7602 (N_7602,N_585,N_3469);
nor U7603 (N_7603,N_2071,N_409);
nand U7604 (N_7604,N_2109,N_1058);
xor U7605 (N_7605,N_4751,N_3525);
and U7606 (N_7606,N_480,N_2014);
nor U7607 (N_7607,N_453,N_2362);
and U7608 (N_7608,N_3083,N_90);
and U7609 (N_7609,N_4693,N_3804);
xor U7610 (N_7610,N_2452,N_4732);
or U7611 (N_7611,N_2943,N_1762);
or U7612 (N_7612,N_512,N_4241);
or U7613 (N_7613,N_4387,N_2337);
or U7614 (N_7614,N_4396,N_901);
xor U7615 (N_7615,N_1433,N_2134);
nor U7616 (N_7616,N_3028,N_1534);
xnor U7617 (N_7617,N_4271,N_1784);
nand U7618 (N_7618,N_3982,N_4705);
nand U7619 (N_7619,N_2430,N_2557);
or U7620 (N_7620,N_2839,N_2181);
nor U7621 (N_7621,N_2333,N_2744);
xnor U7622 (N_7622,N_4081,N_459);
nor U7623 (N_7623,N_1836,N_4920);
nand U7624 (N_7624,N_2586,N_3917);
or U7625 (N_7625,N_3285,N_4900);
or U7626 (N_7626,N_4886,N_1035);
xnor U7627 (N_7627,N_3491,N_1233);
nor U7628 (N_7628,N_2343,N_1351);
and U7629 (N_7629,N_4544,N_860);
xnor U7630 (N_7630,N_2975,N_1880);
xor U7631 (N_7631,N_35,N_3960);
and U7632 (N_7632,N_3263,N_566);
nor U7633 (N_7633,N_4796,N_2250);
and U7634 (N_7634,N_3461,N_3553);
nor U7635 (N_7635,N_2693,N_2730);
and U7636 (N_7636,N_4094,N_4752);
or U7637 (N_7637,N_379,N_2641);
nand U7638 (N_7638,N_4095,N_2942);
nor U7639 (N_7639,N_12,N_4400);
xor U7640 (N_7640,N_3144,N_771);
or U7641 (N_7641,N_659,N_2344);
nor U7642 (N_7642,N_1302,N_4643);
or U7643 (N_7643,N_530,N_2806);
xor U7644 (N_7644,N_4489,N_2570);
nor U7645 (N_7645,N_2659,N_582);
or U7646 (N_7646,N_877,N_248);
and U7647 (N_7647,N_1260,N_1243);
nand U7648 (N_7648,N_61,N_3790);
nor U7649 (N_7649,N_4893,N_2148);
and U7650 (N_7650,N_4138,N_1585);
xor U7651 (N_7651,N_4494,N_1414);
nor U7652 (N_7652,N_1356,N_2717);
nor U7653 (N_7653,N_1530,N_3187);
nor U7654 (N_7654,N_633,N_1719);
and U7655 (N_7655,N_4503,N_3432);
xor U7656 (N_7656,N_692,N_439);
and U7657 (N_7657,N_2622,N_4019);
and U7658 (N_7658,N_444,N_2510);
xnor U7659 (N_7659,N_852,N_2542);
xor U7660 (N_7660,N_2429,N_768);
nand U7661 (N_7661,N_2902,N_105);
or U7662 (N_7662,N_4622,N_1104);
xnor U7663 (N_7663,N_1418,N_913);
and U7664 (N_7664,N_1771,N_3684);
or U7665 (N_7665,N_3766,N_4823);
nand U7666 (N_7666,N_247,N_3750);
nand U7667 (N_7667,N_1587,N_88);
or U7668 (N_7668,N_3383,N_4813);
and U7669 (N_7669,N_4726,N_1728);
and U7670 (N_7670,N_1097,N_1598);
nand U7671 (N_7671,N_1560,N_134);
nand U7672 (N_7672,N_289,N_4147);
and U7673 (N_7673,N_4155,N_843);
or U7674 (N_7674,N_3399,N_3740);
or U7675 (N_7675,N_1213,N_4837);
nor U7676 (N_7676,N_4703,N_1107);
or U7677 (N_7677,N_13,N_157);
nand U7678 (N_7678,N_42,N_3237);
nor U7679 (N_7679,N_3959,N_4744);
nand U7680 (N_7680,N_2681,N_2078);
and U7681 (N_7681,N_1563,N_428);
and U7682 (N_7682,N_4823,N_4606);
xor U7683 (N_7683,N_4456,N_3784);
and U7684 (N_7684,N_1667,N_3625);
xor U7685 (N_7685,N_1349,N_1201);
nand U7686 (N_7686,N_4092,N_3047);
nor U7687 (N_7687,N_1384,N_2269);
xor U7688 (N_7688,N_4615,N_85);
or U7689 (N_7689,N_82,N_2282);
and U7690 (N_7690,N_1745,N_1048);
xnor U7691 (N_7691,N_1036,N_3398);
and U7692 (N_7692,N_2994,N_10);
xnor U7693 (N_7693,N_4184,N_1668);
xnor U7694 (N_7694,N_18,N_1523);
or U7695 (N_7695,N_1650,N_2828);
and U7696 (N_7696,N_4431,N_1467);
or U7697 (N_7697,N_1055,N_278);
or U7698 (N_7698,N_2105,N_875);
nand U7699 (N_7699,N_4711,N_2596);
nand U7700 (N_7700,N_1098,N_1371);
and U7701 (N_7701,N_3201,N_1923);
nand U7702 (N_7702,N_4454,N_3410);
xnor U7703 (N_7703,N_3944,N_1774);
nand U7704 (N_7704,N_1427,N_1620);
nand U7705 (N_7705,N_2543,N_1627);
nand U7706 (N_7706,N_1004,N_448);
xnor U7707 (N_7707,N_2330,N_4605);
or U7708 (N_7708,N_3248,N_2321);
xor U7709 (N_7709,N_3901,N_3635);
or U7710 (N_7710,N_4736,N_3813);
or U7711 (N_7711,N_2416,N_2150);
nand U7712 (N_7712,N_4155,N_1799);
nand U7713 (N_7713,N_1259,N_1219);
nand U7714 (N_7714,N_1924,N_4325);
or U7715 (N_7715,N_1265,N_4263);
and U7716 (N_7716,N_3787,N_2346);
and U7717 (N_7717,N_1272,N_1728);
or U7718 (N_7718,N_359,N_1149);
xnor U7719 (N_7719,N_1697,N_258);
nor U7720 (N_7720,N_712,N_2377);
xnor U7721 (N_7721,N_865,N_2698);
xor U7722 (N_7722,N_3882,N_250);
and U7723 (N_7723,N_2587,N_3636);
or U7724 (N_7724,N_4954,N_2834);
xor U7725 (N_7725,N_126,N_2000);
nand U7726 (N_7726,N_3454,N_1858);
xnor U7727 (N_7727,N_4835,N_3558);
nor U7728 (N_7728,N_4927,N_2079);
and U7729 (N_7729,N_4400,N_4887);
nand U7730 (N_7730,N_4352,N_4648);
nand U7731 (N_7731,N_3399,N_3374);
nand U7732 (N_7732,N_2112,N_2423);
or U7733 (N_7733,N_1720,N_1613);
nand U7734 (N_7734,N_4343,N_3456);
nand U7735 (N_7735,N_1344,N_3708);
and U7736 (N_7736,N_3049,N_4088);
or U7737 (N_7737,N_4776,N_1112);
xor U7738 (N_7738,N_1542,N_1797);
nor U7739 (N_7739,N_1323,N_3779);
xor U7740 (N_7740,N_4677,N_3957);
nor U7741 (N_7741,N_2979,N_3183);
xor U7742 (N_7742,N_1981,N_152);
and U7743 (N_7743,N_3952,N_3899);
and U7744 (N_7744,N_4846,N_583);
nor U7745 (N_7745,N_3789,N_2555);
and U7746 (N_7746,N_2021,N_2794);
or U7747 (N_7747,N_237,N_1523);
and U7748 (N_7748,N_1947,N_614);
and U7749 (N_7749,N_4441,N_3499);
and U7750 (N_7750,N_2525,N_3848);
or U7751 (N_7751,N_3669,N_783);
nand U7752 (N_7752,N_3968,N_517);
and U7753 (N_7753,N_3891,N_2376);
xor U7754 (N_7754,N_3719,N_4867);
and U7755 (N_7755,N_3375,N_4295);
xor U7756 (N_7756,N_1137,N_135);
and U7757 (N_7757,N_653,N_2149);
and U7758 (N_7758,N_3368,N_408);
or U7759 (N_7759,N_2779,N_1257);
xor U7760 (N_7760,N_3499,N_4438);
nor U7761 (N_7761,N_4067,N_2988);
and U7762 (N_7762,N_111,N_143);
nor U7763 (N_7763,N_3134,N_382);
or U7764 (N_7764,N_4195,N_1852);
xor U7765 (N_7765,N_2306,N_2966);
nand U7766 (N_7766,N_4640,N_3850);
or U7767 (N_7767,N_2360,N_3724);
xor U7768 (N_7768,N_3323,N_1448);
xor U7769 (N_7769,N_1675,N_3325);
xnor U7770 (N_7770,N_2261,N_1179);
nand U7771 (N_7771,N_157,N_2187);
nor U7772 (N_7772,N_3140,N_3263);
nor U7773 (N_7773,N_3158,N_3316);
xnor U7774 (N_7774,N_113,N_3487);
nand U7775 (N_7775,N_2018,N_2185);
nand U7776 (N_7776,N_3942,N_4491);
nor U7777 (N_7777,N_2871,N_2575);
nor U7778 (N_7778,N_2292,N_4249);
nor U7779 (N_7779,N_3902,N_3244);
xor U7780 (N_7780,N_1843,N_4505);
xnor U7781 (N_7781,N_3205,N_31);
or U7782 (N_7782,N_381,N_801);
nor U7783 (N_7783,N_4680,N_3289);
and U7784 (N_7784,N_4310,N_71);
nand U7785 (N_7785,N_924,N_1737);
nor U7786 (N_7786,N_4873,N_2801);
nand U7787 (N_7787,N_3373,N_594);
nand U7788 (N_7788,N_2425,N_4164);
nor U7789 (N_7789,N_3877,N_2862);
xor U7790 (N_7790,N_1774,N_4881);
nand U7791 (N_7791,N_276,N_1897);
xnor U7792 (N_7792,N_860,N_1202);
xor U7793 (N_7793,N_3912,N_2137);
or U7794 (N_7794,N_203,N_4353);
or U7795 (N_7795,N_1463,N_1036);
nand U7796 (N_7796,N_1143,N_267);
or U7797 (N_7797,N_849,N_583);
nor U7798 (N_7798,N_1513,N_3839);
xor U7799 (N_7799,N_4997,N_1265);
xor U7800 (N_7800,N_3326,N_3726);
or U7801 (N_7801,N_1166,N_4851);
xnor U7802 (N_7802,N_2299,N_2134);
or U7803 (N_7803,N_1348,N_3856);
nand U7804 (N_7804,N_134,N_2292);
or U7805 (N_7805,N_3832,N_4369);
nor U7806 (N_7806,N_1941,N_1078);
or U7807 (N_7807,N_3383,N_2676);
and U7808 (N_7808,N_2623,N_2612);
nand U7809 (N_7809,N_707,N_3434);
nand U7810 (N_7810,N_4024,N_3326);
xnor U7811 (N_7811,N_2097,N_2561);
and U7812 (N_7812,N_279,N_3168);
or U7813 (N_7813,N_2985,N_656);
nor U7814 (N_7814,N_2518,N_3241);
xor U7815 (N_7815,N_2464,N_2904);
and U7816 (N_7816,N_3052,N_4344);
nand U7817 (N_7817,N_2117,N_210);
xor U7818 (N_7818,N_1857,N_509);
and U7819 (N_7819,N_154,N_2862);
nor U7820 (N_7820,N_658,N_3353);
nor U7821 (N_7821,N_906,N_3338);
and U7822 (N_7822,N_1687,N_321);
xnor U7823 (N_7823,N_3403,N_728);
xnor U7824 (N_7824,N_847,N_3607);
nand U7825 (N_7825,N_65,N_1189);
nand U7826 (N_7826,N_3945,N_477);
xor U7827 (N_7827,N_1044,N_3329);
nor U7828 (N_7828,N_1738,N_645);
nor U7829 (N_7829,N_3799,N_1395);
xnor U7830 (N_7830,N_2637,N_1274);
xor U7831 (N_7831,N_1548,N_2279);
nor U7832 (N_7832,N_3589,N_3106);
and U7833 (N_7833,N_639,N_3815);
and U7834 (N_7834,N_146,N_3398);
or U7835 (N_7835,N_1922,N_76);
and U7836 (N_7836,N_579,N_424);
nand U7837 (N_7837,N_2023,N_567);
nor U7838 (N_7838,N_3523,N_3039);
nand U7839 (N_7839,N_4807,N_3414);
and U7840 (N_7840,N_1240,N_627);
nand U7841 (N_7841,N_2328,N_1793);
or U7842 (N_7842,N_445,N_935);
nand U7843 (N_7843,N_1249,N_1509);
nor U7844 (N_7844,N_2831,N_3993);
xor U7845 (N_7845,N_4433,N_331);
nand U7846 (N_7846,N_2663,N_3645);
xnor U7847 (N_7847,N_2141,N_3091);
nand U7848 (N_7848,N_502,N_891);
xnor U7849 (N_7849,N_2342,N_292);
nand U7850 (N_7850,N_4626,N_847);
xnor U7851 (N_7851,N_2386,N_1197);
nor U7852 (N_7852,N_3117,N_3737);
xnor U7853 (N_7853,N_1532,N_3437);
nand U7854 (N_7854,N_1333,N_731);
nor U7855 (N_7855,N_52,N_4770);
nand U7856 (N_7856,N_4519,N_4155);
xor U7857 (N_7857,N_2461,N_1738);
nor U7858 (N_7858,N_1806,N_2442);
and U7859 (N_7859,N_2033,N_1171);
or U7860 (N_7860,N_727,N_645);
nor U7861 (N_7861,N_4708,N_4256);
and U7862 (N_7862,N_4455,N_2290);
nand U7863 (N_7863,N_4335,N_2426);
nor U7864 (N_7864,N_821,N_407);
nand U7865 (N_7865,N_1737,N_4282);
or U7866 (N_7866,N_1960,N_2678);
nand U7867 (N_7867,N_1034,N_182);
nand U7868 (N_7868,N_367,N_4457);
or U7869 (N_7869,N_3074,N_3492);
or U7870 (N_7870,N_129,N_4559);
nand U7871 (N_7871,N_47,N_4269);
or U7872 (N_7872,N_2154,N_2317);
nand U7873 (N_7873,N_1374,N_3546);
and U7874 (N_7874,N_2565,N_2667);
and U7875 (N_7875,N_631,N_1099);
nor U7876 (N_7876,N_1485,N_1962);
nand U7877 (N_7877,N_362,N_2899);
nor U7878 (N_7878,N_4588,N_1799);
or U7879 (N_7879,N_2287,N_2529);
or U7880 (N_7880,N_3645,N_365);
or U7881 (N_7881,N_888,N_4474);
or U7882 (N_7882,N_270,N_376);
nand U7883 (N_7883,N_2204,N_2287);
nor U7884 (N_7884,N_1900,N_4206);
nor U7885 (N_7885,N_2372,N_4921);
nand U7886 (N_7886,N_4174,N_1451);
nor U7887 (N_7887,N_4753,N_4339);
nand U7888 (N_7888,N_4093,N_1877);
xor U7889 (N_7889,N_4003,N_4393);
and U7890 (N_7890,N_588,N_2041);
nor U7891 (N_7891,N_2415,N_237);
or U7892 (N_7892,N_1393,N_2120);
nor U7893 (N_7893,N_1861,N_218);
nor U7894 (N_7894,N_2416,N_454);
nor U7895 (N_7895,N_1709,N_2350);
nor U7896 (N_7896,N_1590,N_3096);
xor U7897 (N_7897,N_4837,N_3199);
or U7898 (N_7898,N_887,N_4341);
xor U7899 (N_7899,N_484,N_15);
xnor U7900 (N_7900,N_2732,N_3042);
and U7901 (N_7901,N_2561,N_1383);
and U7902 (N_7902,N_1369,N_4587);
xor U7903 (N_7903,N_3059,N_407);
nor U7904 (N_7904,N_3333,N_2292);
and U7905 (N_7905,N_1987,N_1202);
nand U7906 (N_7906,N_533,N_2378);
and U7907 (N_7907,N_2540,N_669);
nor U7908 (N_7908,N_4114,N_2438);
xnor U7909 (N_7909,N_3058,N_4049);
and U7910 (N_7910,N_404,N_2738);
nor U7911 (N_7911,N_3421,N_2483);
xnor U7912 (N_7912,N_4491,N_4890);
xor U7913 (N_7913,N_1336,N_1846);
nor U7914 (N_7914,N_2988,N_1015);
nor U7915 (N_7915,N_2963,N_4616);
xor U7916 (N_7916,N_739,N_308);
or U7917 (N_7917,N_3934,N_4494);
or U7918 (N_7918,N_292,N_1014);
xor U7919 (N_7919,N_773,N_1063);
nor U7920 (N_7920,N_904,N_3507);
and U7921 (N_7921,N_4069,N_1334);
and U7922 (N_7922,N_3468,N_3197);
nor U7923 (N_7923,N_4511,N_4108);
xor U7924 (N_7924,N_2744,N_4562);
and U7925 (N_7925,N_4132,N_4237);
nor U7926 (N_7926,N_1734,N_1784);
xnor U7927 (N_7927,N_3825,N_314);
xor U7928 (N_7928,N_4273,N_2667);
nor U7929 (N_7929,N_1137,N_4317);
and U7930 (N_7930,N_4289,N_3282);
or U7931 (N_7931,N_1229,N_122);
xnor U7932 (N_7932,N_1559,N_164);
xor U7933 (N_7933,N_819,N_3233);
xor U7934 (N_7934,N_4606,N_2131);
and U7935 (N_7935,N_2590,N_2266);
nor U7936 (N_7936,N_4715,N_1665);
xnor U7937 (N_7937,N_4695,N_483);
xnor U7938 (N_7938,N_1001,N_2750);
xor U7939 (N_7939,N_4121,N_754);
and U7940 (N_7940,N_2242,N_4783);
xnor U7941 (N_7941,N_3903,N_4141);
or U7942 (N_7942,N_1434,N_4372);
and U7943 (N_7943,N_2216,N_3931);
or U7944 (N_7944,N_115,N_705);
nor U7945 (N_7945,N_3073,N_4086);
and U7946 (N_7946,N_375,N_2636);
nor U7947 (N_7947,N_2809,N_361);
or U7948 (N_7948,N_3489,N_285);
xor U7949 (N_7949,N_447,N_2753);
xnor U7950 (N_7950,N_2597,N_1536);
xor U7951 (N_7951,N_3729,N_48);
or U7952 (N_7952,N_121,N_1790);
and U7953 (N_7953,N_4770,N_3159);
xnor U7954 (N_7954,N_325,N_1752);
and U7955 (N_7955,N_1540,N_1422);
nor U7956 (N_7956,N_1289,N_2612);
nand U7957 (N_7957,N_2490,N_1370);
nor U7958 (N_7958,N_617,N_1988);
or U7959 (N_7959,N_754,N_4388);
nor U7960 (N_7960,N_2275,N_464);
or U7961 (N_7961,N_1530,N_2345);
and U7962 (N_7962,N_1458,N_4390);
nand U7963 (N_7963,N_1646,N_567);
nand U7964 (N_7964,N_3456,N_2457);
and U7965 (N_7965,N_3441,N_3356);
xor U7966 (N_7966,N_4807,N_4666);
xor U7967 (N_7967,N_2877,N_993);
nor U7968 (N_7968,N_695,N_4161);
and U7969 (N_7969,N_3939,N_3206);
xnor U7970 (N_7970,N_4728,N_2100);
xor U7971 (N_7971,N_806,N_3750);
xnor U7972 (N_7972,N_824,N_807);
nor U7973 (N_7973,N_4715,N_3681);
xor U7974 (N_7974,N_3223,N_3443);
xnor U7975 (N_7975,N_2970,N_4046);
xnor U7976 (N_7976,N_2017,N_3145);
and U7977 (N_7977,N_1385,N_2300);
nor U7978 (N_7978,N_4389,N_4371);
nor U7979 (N_7979,N_2338,N_2911);
nand U7980 (N_7980,N_4930,N_3900);
nand U7981 (N_7981,N_3194,N_1807);
nor U7982 (N_7982,N_1539,N_2237);
nand U7983 (N_7983,N_957,N_928);
nor U7984 (N_7984,N_1048,N_4232);
nor U7985 (N_7985,N_2144,N_226);
or U7986 (N_7986,N_2895,N_286);
nand U7987 (N_7987,N_1260,N_2510);
and U7988 (N_7988,N_3355,N_195);
xor U7989 (N_7989,N_2181,N_3073);
nor U7990 (N_7990,N_2266,N_4290);
or U7991 (N_7991,N_2720,N_2779);
nand U7992 (N_7992,N_4450,N_981);
and U7993 (N_7993,N_4920,N_4310);
nor U7994 (N_7994,N_4758,N_171);
and U7995 (N_7995,N_4191,N_144);
or U7996 (N_7996,N_3057,N_1639);
nand U7997 (N_7997,N_4535,N_4543);
nor U7998 (N_7998,N_3079,N_878);
xnor U7999 (N_7999,N_1193,N_2823);
or U8000 (N_8000,N_1629,N_3554);
nor U8001 (N_8001,N_4286,N_2357);
and U8002 (N_8002,N_1331,N_1177);
nor U8003 (N_8003,N_4102,N_3739);
or U8004 (N_8004,N_3925,N_2203);
nor U8005 (N_8005,N_3359,N_2514);
nor U8006 (N_8006,N_735,N_2528);
xor U8007 (N_8007,N_1897,N_3933);
nand U8008 (N_8008,N_160,N_2841);
xor U8009 (N_8009,N_2226,N_1191);
nand U8010 (N_8010,N_2288,N_1940);
xnor U8011 (N_8011,N_394,N_4337);
and U8012 (N_8012,N_2262,N_2279);
and U8013 (N_8013,N_660,N_4357);
nand U8014 (N_8014,N_506,N_4323);
nor U8015 (N_8015,N_1635,N_843);
or U8016 (N_8016,N_2771,N_498);
and U8017 (N_8017,N_91,N_2913);
or U8018 (N_8018,N_3729,N_1994);
nand U8019 (N_8019,N_4584,N_1301);
xor U8020 (N_8020,N_4461,N_2505);
or U8021 (N_8021,N_1871,N_3546);
or U8022 (N_8022,N_4473,N_1586);
or U8023 (N_8023,N_2276,N_1194);
and U8024 (N_8024,N_4807,N_4457);
nor U8025 (N_8025,N_696,N_1425);
or U8026 (N_8026,N_3098,N_2465);
nor U8027 (N_8027,N_196,N_1298);
xnor U8028 (N_8028,N_3024,N_2335);
nand U8029 (N_8029,N_1222,N_870);
or U8030 (N_8030,N_1636,N_691);
nand U8031 (N_8031,N_4603,N_2732);
and U8032 (N_8032,N_4468,N_2610);
nor U8033 (N_8033,N_572,N_3916);
xor U8034 (N_8034,N_1482,N_1729);
or U8035 (N_8035,N_4449,N_1343);
nand U8036 (N_8036,N_52,N_3816);
or U8037 (N_8037,N_3247,N_720);
nand U8038 (N_8038,N_1515,N_2457);
xor U8039 (N_8039,N_2001,N_3891);
and U8040 (N_8040,N_1966,N_3643);
and U8041 (N_8041,N_1813,N_4626);
xor U8042 (N_8042,N_3809,N_850);
nor U8043 (N_8043,N_821,N_836);
and U8044 (N_8044,N_1836,N_4932);
and U8045 (N_8045,N_1565,N_1390);
or U8046 (N_8046,N_1159,N_3114);
xor U8047 (N_8047,N_1917,N_568);
or U8048 (N_8048,N_4086,N_3982);
or U8049 (N_8049,N_4706,N_4159);
and U8050 (N_8050,N_1369,N_3344);
xor U8051 (N_8051,N_2400,N_1517);
nand U8052 (N_8052,N_3762,N_2918);
nand U8053 (N_8053,N_2386,N_1438);
and U8054 (N_8054,N_3555,N_3900);
nand U8055 (N_8055,N_4081,N_2153);
nor U8056 (N_8056,N_3703,N_3562);
xor U8057 (N_8057,N_3127,N_1482);
or U8058 (N_8058,N_2815,N_3981);
nor U8059 (N_8059,N_1121,N_2520);
or U8060 (N_8060,N_3308,N_636);
xnor U8061 (N_8061,N_3296,N_3521);
or U8062 (N_8062,N_4632,N_1860);
or U8063 (N_8063,N_351,N_4255);
and U8064 (N_8064,N_4528,N_1982);
nand U8065 (N_8065,N_2994,N_2563);
and U8066 (N_8066,N_1136,N_2436);
or U8067 (N_8067,N_2709,N_2427);
nor U8068 (N_8068,N_4423,N_3962);
or U8069 (N_8069,N_2258,N_2406);
nand U8070 (N_8070,N_1279,N_4130);
nor U8071 (N_8071,N_501,N_1473);
nor U8072 (N_8072,N_5,N_4225);
nor U8073 (N_8073,N_1902,N_3254);
or U8074 (N_8074,N_3720,N_2720);
nor U8075 (N_8075,N_1242,N_626);
or U8076 (N_8076,N_440,N_2879);
nor U8077 (N_8077,N_346,N_2298);
nand U8078 (N_8078,N_3569,N_2373);
or U8079 (N_8079,N_1162,N_658);
or U8080 (N_8080,N_4568,N_3163);
nand U8081 (N_8081,N_125,N_3993);
xor U8082 (N_8082,N_3907,N_2835);
nor U8083 (N_8083,N_4285,N_1091);
or U8084 (N_8084,N_1125,N_3648);
nand U8085 (N_8085,N_3859,N_2668);
or U8086 (N_8086,N_2616,N_4724);
nand U8087 (N_8087,N_2792,N_2762);
and U8088 (N_8088,N_4483,N_1328);
xnor U8089 (N_8089,N_3811,N_655);
nand U8090 (N_8090,N_4296,N_266);
xor U8091 (N_8091,N_311,N_3126);
nand U8092 (N_8092,N_4714,N_3048);
xor U8093 (N_8093,N_1752,N_651);
xor U8094 (N_8094,N_1213,N_1957);
xor U8095 (N_8095,N_1999,N_2363);
xnor U8096 (N_8096,N_3078,N_2590);
nand U8097 (N_8097,N_4568,N_2361);
xor U8098 (N_8098,N_1878,N_1348);
xnor U8099 (N_8099,N_3891,N_4465);
xnor U8100 (N_8100,N_2148,N_2144);
xnor U8101 (N_8101,N_853,N_3837);
and U8102 (N_8102,N_4979,N_4913);
xnor U8103 (N_8103,N_3993,N_2572);
or U8104 (N_8104,N_2551,N_3539);
nand U8105 (N_8105,N_1961,N_995);
or U8106 (N_8106,N_2064,N_2765);
xnor U8107 (N_8107,N_894,N_3680);
and U8108 (N_8108,N_3013,N_4603);
or U8109 (N_8109,N_1832,N_4917);
xnor U8110 (N_8110,N_4016,N_3618);
nor U8111 (N_8111,N_4570,N_4482);
or U8112 (N_8112,N_2638,N_3429);
and U8113 (N_8113,N_2817,N_1682);
and U8114 (N_8114,N_1213,N_349);
or U8115 (N_8115,N_4169,N_2108);
and U8116 (N_8116,N_2197,N_3403);
xor U8117 (N_8117,N_497,N_3237);
xor U8118 (N_8118,N_4493,N_2586);
nor U8119 (N_8119,N_4404,N_1385);
and U8120 (N_8120,N_4932,N_196);
or U8121 (N_8121,N_3424,N_3809);
nand U8122 (N_8122,N_3836,N_1371);
nand U8123 (N_8123,N_3991,N_2372);
or U8124 (N_8124,N_4332,N_2303);
nor U8125 (N_8125,N_128,N_3654);
nand U8126 (N_8126,N_762,N_1842);
nand U8127 (N_8127,N_1186,N_1077);
nor U8128 (N_8128,N_3205,N_199);
nor U8129 (N_8129,N_377,N_219);
nand U8130 (N_8130,N_2653,N_148);
and U8131 (N_8131,N_4790,N_2491);
xor U8132 (N_8132,N_4469,N_1940);
or U8133 (N_8133,N_453,N_2080);
and U8134 (N_8134,N_2285,N_484);
and U8135 (N_8135,N_3292,N_1128);
and U8136 (N_8136,N_4589,N_195);
or U8137 (N_8137,N_3266,N_4558);
or U8138 (N_8138,N_4046,N_3781);
nand U8139 (N_8139,N_4040,N_3524);
xnor U8140 (N_8140,N_2454,N_1518);
nor U8141 (N_8141,N_4363,N_2462);
or U8142 (N_8142,N_1314,N_3479);
and U8143 (N_8143,N_4796,N_4420);
nand U8144 (N_8144,N_3240,N_2476);
or U8145 (N_8145,N_933,N_2317);
nand U8146 (N_8146,N_3178,N_453);
and U8147 (N_8147,N_2640,N_404);
nand U8148 (N_8148,N_3973,N_4208);
nand U8149 (N_8149,N_885,N_4332);
nand U8150 (N_8150,N_661,N_3478);
xnor U8151 (N_8151,N_724,N_3856);
xnor U8152 (N_8152,N_645,N_1774);
or U8153 (N_8153,N_4028,N_2543);
xnor U8154 (N_8154,N_3853,N_133);
nand U8155 (N_8155,N_4200,N_2972);
nand U8156 (N_8156,N_374,N_2454);
xor U8157 (N_8157,N_3026,N_4450);
and U8158 (N_8158,N_3523,N_1765);
or U8159 (N_8159,N_185,N_728);
or U8160 (N_8160,N_254,N_4190);
nand U8161 (N_8161,N_553,N_3138);
and U8162 (N_8162,N_1250,N_4126);
nor U8163 (N_8163,N_942,N_902);
nand U8164 (N_8164,N_1945,N_3754);
nor U8165 (N_8165,N_307,N_1136);
xor U8166 (N_8166,N_727,N_2158);
nand U8167 (N_8167,N_3629,N_467);
xnor U8168 (N_8168,N_4450,N_1025);
and U8169 (N_8169,N_343,N_4894);
xor U8170 (N_8170,N_4019,N_3520);
nor U8171 (N_8171,N_3122,N_3563);
nor U8172 (N_8172,N_1103,N_312);
or U8173 (N_8173,N_2542,N_3974);
nor U8174 (N_8174,N_3036,N_4251);
nor U8175 (N_8175,N_1731,N_3655);
nand U8176 (N_8176,N_3325,N_4382);
nor U8177 (N_8177,N_3570,N_1265);
or U8178 (N_8178,N_4354,N_505);
xnor U8179 (N_8179,N_3739,N_760);
nand U8180 (N_8180,N_3591,N_1262);
and U8181 (N_8181,N_3137,N_4418);
nor U8182 (N_8182,N_4982,N_4804);
xnor U8183 (N_8183,N_2314,N_4730);
nor U8184 (N_8184,N_3734,N_4245);
and U8185 (N_8185,N_4738,N_4920);
or U8186 (N_8186,N_3375,N_535);
and U8187 (N_8187,N_1141,N_766);
nand U8188 (N_8188,N_4365,N_2681);
nor U8189 (N_8189,N_2805,N_3756);
nand U8190 (N_8190,N_3059,N_3331);
nor U8191 (N_8191,N_710,N_869);
or U8192 (N_8192,N_3810,N_302);
nand U8193 (N_8193,N_926,N_4159);
nor U8194 (N_8194,N_981,N_3970);
xnor U8195 (N_8195,N_2420,N_4873);
and U8196 (N_8196,N_2790,N_4598);
nor U8197 (N_8197,N_2039,N_3783);
xor U8198 (N_8198,N_3334,N_3469);
and U8199 (N_8199,N_4109,N_217);
nand U8200 (N_8200,N_160,N_4909);
and U8201 (N_8201,N_2828,N_3524);
and U8202 (N_8202,N_1199,N_1983);
xnor U8203 (N_8203,N_2302,N_1055);
and U8204 (N_8204,N_747,N_3229);
or U8205 (N_8205,N_3539,N_1429);
nand U8206 (N_8206,N_1165,N_3708);
nand U8207 (N_8207,N_3406,N_4631);
or U8208 (N_8208,N_1733,N_4707);
or U8209 (N_8209,N_1714,N_4943);
or U8210 (N_8210,N_385,N_1922);
xnor U8211 (N_8211,N_3398,N_1233);
nand U8212 (N_8212,N_4099,N_4938);
nand U8213 (N_8213,N_3920,N_2754);
and U8214 (N_8214,N_3098,N_110);
nand U8215 (N_8215,N_1666,N_4641);
nand U8216 (N_8216,N_121,N_3128);
xnor U8217 (N_8217,N_2977,N_683);
nor U8218 (N_8218,N_684,N_1950);
nand U8219 (N_8219,N_1358,N_3017);
and U8220 (N_8220,N_673,N_3083);
xnor U8221 (N_8221,N_2262,N_106);
nor U8222 (N_8222,N_2152,N_43);
nand U8223 (N_8223,N_1934,N_2164);
or U8224 (N_8224,N_4904,N_1069);
or U8225 (N_8225,N_2907,N_4334);
or U8226 (N_8226,N_3912,N_3951);
nor U8227 (N_8227,N_3919,N_3312);
or U8228 (N_8228,N_4344,N_3005);
nor U8229 (N_8229,N_562,N_3918);
nor U8230 (N_8230,N_466,N_1952);
nor U8231 (N_8231,N_4442,N_365);
and U8232 (N_8232,N_2727,N_1977);
nor U8233 (N_8233,N_1070,N_4972);
and U8234 (N_8234,N_1781,N_3333);
nor U8235 (N_8235,N_3366,N_1852);
and U8236 (N_8236,N_1562,N_2088);
and U8237 (N_8237,N_4813,N_1147);
and U8238 (N_8238,N_753,N_4600);
or U8239 (N_8239,N_4614,N_3434);
xor U8240 (N_8240,N_3744,N_995);
and U8241 (N_8241,N_4991,N_2064);
xor U8242 (N_8242,N_3410,N_467);
nand U8243 (N_8243,N_1366,N_2968);
nor U8244 (N_8244,N_200,N_2926);
and U8245 (N_8245,N_1776,N_2672);
xor U8246 (N_8246,N_3947,N_1888);
nand U8247 (N_8247,N_537,N_4333);
nor U8248 (N_8248,N_1685,N_3851);
nor U8249 (N_8249,N_1312,N_1608);
nand U8250 (N_8250,N_1637,N_2680);
xor U8251 (N_8251,N_131,N_2876);
or U8252 (N_8252,N_3252,N_2525);
nand U8253 (N_8253,N_1746,N_1706);
and U8254 (N_8254,N_1041,N_2308);
nand U8255 (N_8255,N_289,N_1221);
xor U8256 (N_8256,N_1576,N_355);
nor U8257 (N_8257,N_3837,N_3201);
nor U8258 (N_8258,N_2533,N_3100);
xor U8259 (N_8259,N_3474,N_2913);
nor U8260 (N_8260,N_4367,N_4406);
xnor U8261 (N_8261,N_4381,N_2771);
nor U8262 (N_8262,N_3517,N_1812);
or U8263 (N_8263,N_1653,N_3935);
and U8264 (N_8264,N_2073,N_3683);
nor U8265 (N_8265,N_2980,N_677);
nor U8266 (N_8266,N_1464,N_3049);
and U8267 (N_8267,N_4108,N_2381);
xor U8268 (N_8268,N_501,N_2850);
nor U8269 (N_8269,N_1146,N_1294);
or U8270 (N_8270,N_2372,N_724);
or U8271 (N_8271,N_624,N_161);
nand U8272 (N_8272,N_4838,N_2145);
nor U8273 (N_8273,N_4219,N_3497);
nand U8274 (N_8274,N_2972,N_4318);
nand U8275 (N_8275,N_4419,N_4964);
nor U8276 (N_8276,N_4236,N_4068);
nand U8277 (N_8277,N_3146,N_4535);
xor U8278 (N_8278,N_1840,N_3521);
xnor U8279 (N_8279,N_4808,N_430);
xor U8280 (N_8280,N_3330,N_2082);
nand U8281 (N_8281,N_490,N_4131);
and U8282 (N_8282,N_3383,N_3496);
nand U8283 (N_8283,N_2140,N_2430);
nand U8284 (N_8284,N_3003,N_4384);
nand U8285 (N_8285,N_622,N_3373);
nor U8286 (N_8286,N_4673,N_4724);
nand U8287 (N_8287,N_391,N_706);
nand U8288 (N_8288,N_868,N_4500);
or U8289 (N_8289,N_4717,N_2723);
nand U8290 (N_8290,N_3236,N_768);
xor U8291 (N_8291,N_2447,N_2464);
or U8292 (N_8292,N_4755,N_3991);
nand U8293 (N_8293,N_182,N_3321);
nor U8294 (N_8294,N_753,N_560);
or U8295 (N_8295,N_509,N_412);
xnor U8296 (N_8296,N_2982,N_2324);
nor U8297 (N_8297,N_1975,N_1618);
nand U8298 (N_8298,N_3119,N_406);
or U8299 (N_8299,N_2005,N_4668);
or U8300 (N_8300,N_133,N_4970);
nor U8301 (N_8301,N_228,N_2838);
and U8302 (N_8302,N_4242,N_641);
nand U8303 (N_8303,N_69,N_3354);
nand U8304 (N_8304,N_4907,N_2109);
and U8305 (N_8305,N_1726,N_2496);
nor U8306 (N_8306,N_4165,N_172);
nor U8307 (N_8307,N_2661,N_502);
nor U8308 (N_8308,N_3088,N_3351);
nor U8309 (N_8309,N_1316,N_3634);
nand U8310 (N_8310,N_2734,N_3292);
xnor U8311 (N_8311,N_2316,N_1458);
or U8312 (N_8312,N_2274,N_2517);
nor U8313 (N_8313,N_3597,N_4837);
or U8314 (N_8314,N_1966,N_1826);
or U8315 (N_8315,N_922,N_4249);
and U8316 (N_8316,N_311,N_156);
or U8317 (N_8317,N_4480,N_143);
and U8318 (N_8318,N_3286,N_2379);
and U8319 (N_8319,N_1946,N_4742);
and U8320 (N_8320,N_2951,N_2476);
nand U8321 (N_8321,N_655,N_947);
nand U8322 (N_8322,N_797,N_325);
nand U8323 (N_8323,N_1798,N_882);
and U8324 (N_8324,N_3622,N_1082);
or U8325 (N_8325,N_1736,N_1914);
nor U8326 (N_8326,N_59,N_3329);
or U8327 (N_8327,N_1229,N_3869);
nor U8328 (N_8328,N_4214,N_1600);
nand U8329 (N_8329,N_1844,N_4647);
nor U8330 (N_8330,N_4369,N_4241);
or U8331 (N_8331,N_1559,N_4973);
nand U8332 (N_8332,N_405,N_3787);
xor U8333 (N_8333,N_3901,N_137);
or U8334 (N_8334,N_3519,N_4533);
and U8335 (N_8335,N_4261,N_1130);
nand U8336 (N_8336,N_2558,N_4781);
or U8337 (N_8337,N_4953,N_565);
or U8338 (N_8338,N_1121,N_2528);
nand U8339 (N_8339,N_3660,N_220);
and U8340 (N_8340,N_1815,N_2595);
or U8341 (N_8341,N_2084,N_2506);
nand U8342 (N_8342,N_34,N_4657);
and U8343 (N_8343,N_122,N_4986);
nand U8344 (N_8344,N_2333,N_4560);
and U8345 (N_8345,N_177,N_2008);
or U8346 (N_8346,N_241,N_319);
xnor U8347 (N_8347,N_1278,N_2280);
xnor U8348 (N_8348,N_3141,N_1312);
or U8349 (N_8349,N_1905,N_3036);
or U8350 (N_8350,N_3112,N_2139);
nand U8351 (N_8351,N_3718,N_1532);
or U8352 (N_8352,N_3974,N_4226);
xnor U8353 (N_8353,N_1633,N_1214);
and U8354 (N_8354,N_1296,N_4534);
xor U8355 (N_8355,N_3970,N_2611);
nand U8356 (N_8356,N_2974,N_2754);
and U8357 (N_8357,N_852,N_3233);
and U8358 (N_8358,N_926,N_3446);
or U8359 (N_8359,N_1013,N_4490);
and U8360 (N_8360,N_166,N_3026);
nor U8361 (N_8361,N_918,N_83);
nand U8362 (N_8362,N_2190,N_975);
nor U8363 (N_8363,N_1656,N_3500);
xnor U8364 (N_8364,N_2253,N_1556);
nor U8365 (N_8365,N_709,N_16);
xnor U8366 (N_8366,N_2963,N_4009);
and U8367 (N_8367,N_4402,N_248);
nor U8368 (N_8368,N_272,N_2892);
and U8369 (N_8369,N_571,N_2873);
and U8370 (N_8370,N_2085,N_243);
xor U8371 (N_8371,N_3513,N_1321);
and U8372 (N_8372,N_4375,N_271);
nor U8373 (N_8373,N_936,N_4237);
nand U8374 (N_8374,N_2860,N_4976);
or U8375 (N_8375,N_4912,N_2352);
xnor U8376 (N_8376,N_846,N_3179);
or U8377 (N_8377,N_78,N_492);
or U8378 (N_8378,N_4513,N_521);
and U8379 (N_8379,N_3092,N_1007);
nand U8380 (N_8380,N_4327,N_1847);
xor U8381 (N_8381,N_695,N_19);
xnor U8382 (N_8382,N_41,N_1057);
nand U8383 (N_8383,N_4855,N_970);
or U8384 (N_8384,N_486,N_780);
nor U8385 (N_8385,N_2143,N_1668);
nor U8386 (N_8386,N_4278,N_4281);
nand U8387 (N_8387,N_1688,N_1065);
and U8388 (N_8388,N_3564,N_1812);
nor U8389 (N_8389,N_3494,N_507);
and U8390 (N_8390,N_2701,N_3553);
nor U8391 (N_8391,N_1784,N_574);
and U8392 (N_8392,N_314,N_1744);
nor U8393 (N_8393,N_1250,N_1238);
nor U8394 (N_8394,N_1374,N_4892);
xor U8395 (N_8395,N_874,N_3295);
nand U8396 (N_8396,N_549,N_4380);
nor U8397 (N_8397,N_3208,N_2044);
nand U8398 (N_8398,N_2883,N_3304);
xor U8399 (N_8399,N_2681,N_595);
nor U8400 (N_8400,N_3559,N_3392);
and U8401 (N_8401,N_3147,N_2174);
nor U8402 (N_8402,N_2833,N_2696);
nand U8403 (N_8403,N_281,N_3693);
and U8404 (N_8404,N_819,N_4372);
nand U8405 (N_8405,N_3680,N_1776);
nor U8406 (N_8406,N_3184,N_665);
and U8407 (N_8407,N_1359,N_3478);
xor U8408 (N_8408,N_465,N_4610);
xnor U8409 (N_8409,N_3139,N_2471);
nor U8410 (N_8410,N_1295,N_4859);
and U8411 (N_8411,N_3347,N_191);
and U8412 (N_8412,N_2531,N_3414);
and U8413 (N_8413,N_2444,N_3264);
or U8414 (N_8414,N_3868,N_2525);
nand U8415 (N_8415,N_2602,N_13);
or U8416 (N_8416,N_3324,N_3506);
nand U8417 (N_8417,N_3448,N_3181);
xnor U8418 (N_8418,N_2614,N_1372);
and U8419 (N_8419,N_2631,N_3528);
or U8420 (N_8420,N_201,N_2813);
xnor U8421 (N_8421,N_4608,N_4125);
or U8422 (N_8422,N_3037,N_3371);
nand U8423 (N_8423,N_4411,N_1235);
nor U8424 (N_8424,N_1889,N_978);
or U8425 (N_8425,N_4664,N_1179);
xnor U8426 (N_8426,N_2300,N_3508);
nor U8427 (N_8427,N_2650,N_1904);
or U8428 (N_8428,N_2276,N_3730);
or U8429 (N_8429,N_3627,N_1436);
xor U8430 (N_8430,N_1403,N_1487);
xor U8431 (N_8431,N_4510,N_3422);
or U8432 (N_8432,N_2513,N_2640);
xnor U8433 (N_8433,N_268,N_4002);
nand U8434 (N_8434,N_2140,N_2588);
or U8435 (N_8435,N_389,N_3259);
or U8436 (N_8436,N_48,N_1161);
nor U8437 (N_8437,N_2568,N_1708);
nor U8438 (N_8438,N_1102,N_2399);
nor U8439 (N_8439,N_2324,N_1075);
or U8440 (N_8440,N_1320,N_4322);
nor U8441 (N_8441,N_4191,N_1018);
nand U8442 (N_8442,N_3066,N_1677);
or U8443 (N_8443,N_1519,N_2887);
nand U8444 (N_8444,N_4780,N_4251);
nand U8445 (N_8445,N_342,N_2744);
or U8446 (N_8446,N_1563,N_2609);
and U8447 (N_8447,N_1318,N_1272);
nor U8448 (N_8448,N_160,N_1164);
nand U8449 (N_8449,N_2140,N_3920);
xnor U8450 (N_8450,N_3291,N_457);
and U8451 (N_8451,N_2855,N_4501);
or U8452 (N_8452,N_1494,N_4210);
nand U8453 (N_8453,N_1387,N_2827);
nor U8454 (N_8454,N_3742,N_1948);
or U8455 (N_8455,N_3342,N_4755);
nor U8456 (N_8456,N_2018,N_4494);
or U8457 (N_8457,N_896,N_3683);
nor U8458 (N_8458,N_4198,N_2025);
nand U8459 (N_8459,N_4135,N_3560);
or U8460 (N_8460,N_1173,N_2599);
or U8461 (N_8461,N_4565,N_1717);
nand U8462 (N_8462,N_1399,N_4660);
xnor U8463 (N_8463,N_2954,N_1458);
or U8464 (N_8464,N_3330,N_742);
xor U8465 (N_8465,N_4626,N_4114);
xnor U8466 (N_8466,N_4604,N_230);
nor U8467 (N_8467,N_4322,N_1205);
or U8468 (N_8468,N_4808,N_2822);
nor U8469 (N_8469,N_2479,N_4660);
and U8470 (N_8470,N_4575,N_4108);
and U8471 (N_8471,N_2641,N_1724);
xnor U8472 (N_8472,N_4188,N_4063);
nand U8473 (N_8473,N_3391,N_4673);
and U8474 (N_8474,N_2649,N_2976);
nor U8475 (N_8475,N_542,N_4469);
nor U8476 (N_8476,N_1351,N_133);
nor U8477 (N_8477,N_1374,N_3195);
and U8478 (N_8478,N_3704,N_3393);
or U8479 (N_8479,N_1103,N_3252);
nand U8480 (N_8480,N_4858,N_1833);
xor U8481 (N_8481,N_193,N_4437);
and U8482 (N_8482,N_3381,N_671);
nor U8483 (N_8483,N_802,N_3075);
nor U8484 (N_8484,N_2239,N_4249);
nand U8485 (N_8485,N_1169,N_4606);
nand U8486 (N_8486,N_3754,N_1617);
and U8487 (N_8487,N_2679,N_824);
or U8488 (N_8488,N_4860,N_4104);
nor U8489 (N_8489,N_2437,N_1318);
xor U8490 (N_8490,N_4407,N_3280);
xnor U8491 (N_8491,N_653,N_127);
or U8492 (N_8492,N_2138,N_3885);
nand U8493 (N_8493,N_3174,N_4860);
xor U8494 (N_8494,N_2001,N_4812);
xor U8495 (N_8495,N_2593,N_906);
nor U8496 (N_8496,N_2494,N_927);
or U8497 (N_8497,N_4537,N_4090);
xor U8498 (N_8498,N_2725,N_2466);
and U8499 (N_8499,N_1363,N_2358);
xor U8500 (N_8500,N_37,N_3409);
or U8501 (N_8501,N_61,N_3560);
nand U8502 (N_8502,N_4080,N_4811);
xor U8503 (N_8503,N_1753,N_2964);
xor U8504 (N_8504,N_3380,N_4870);
nand U8505 (N_8505,N_228,N_1621);
or U8506 (N_8506,N_2071,N_4002);
and U8507 (N_8507,N_4285,N_797);
nand U8508 (N_8508,N_2149,N_4613);
nor U8509 (N_8509,N_1735,N_1229);
or U8510 (N_8510,N_4803,N_2549);
nand U8511 (N_8511,N_1494,N_2773);
xnor U8512 (N_8512,N_1512,N_2292);
nor U8513 (N_8513,N_3442,N_705);
and U8514 (N_8514,N_857,N_3738);
or U8515 (N_8515,N_1056,N_3332);
nand U8516 (N_8516,N_1456,N_4340);
and U8517 (N_8517,N_1309,N_790);
and U8518 (N_8518,N_2568,N_1669);
and U8519 (N_8519,N_3967,N_1609);
or U8520 (N_8520,N_192,N_3923);
or U8521 (N_8521,N_727,N_4161);
nor U8522 (N_8522,N_3989,N_4960);
or U8523 (N_8523,N_2162,N_1114);
and U8524 (N_8524,N_895,N_2407);
nor U8525 (N_8525,N_1533,N_1608);
nor U8526 (N_8526,N_4243,N_2546);
xnor U8527 (N_8527,N_634,N_2263);
nand U8528 (N_8528,N_1793,N_4266);
nor U8529 (N_8529,N_3321,N_1860);
nand U8530 (N_8530,N_2257,N_971);
and U8531 (N_8531,N_2952,N_2121);
or U8532 (N_8532,N_2081,N_175);
nand U8533 (N_8533,N_1902,N_226);
and U8534 (N_8534,N_850,N_198);
nor U8535 (N_8535,N_3932,N_4409);
nand U8536 (N_8536,N_2540,N_171);
nor U8537 (N_8537,N_4152,N_3045);
and U8538 (N_8538,N_3482,N_1766);
or U8539 (N_8539,N_3561,N_1265);
xnor U8540 (N_8540,N_4111,N_1739);
xnor U8541 (N_8541,N_1464,N_3727);
or U8542 (N_8542,N_2988,N_4945);
or U8543 (N_8543,N_1569,N_2873);
xor U8544 (N_8544,N_1348,N_716);
xor U8545 (N_8545,N_2066,N_3961);
nand U8546 (N_8546,N_2377,N_2540);
xnor U8547 (N_8547,N_1621,N_2564);
xnor U8548 (N_8548,N_627,N_1740);
nand U8549 (N_8549,N_1132,N_4330);
nor U8550 (N_8550,N_1057,N_3049);
nor U8551 (N_8551,N_4191,N_3034);
xnor U8552 (N_8552,N_4695,N_2793);
xor U8553 (N_8553,N_994,N_2860);
nand U8554 (N_8554,N_2613,N_4885);
nor U8555 (N_8555,N_4242,N_1275);
or U8556 (N_8556,N_4519,N_2811);
nor U8557 (N_8557,N_200,N_3063);
or U8558 (N_8558,N_4895,N_4810);
nand U8559 (N_8559,N_1671,N_1637);
nand U8560 (N_8560,N_1626,N_3186);
or U8561 (N_8561,N_3284,N_4858);
xor U8562 (N_8562,N_3095,N_3683);
xnor U8563 (N_8563,N_169,N_2587);
or U8564 (N_8564,N_3704,N_4516);
nand U8565 (N_8565,N_3488,N_3838);
nand U8566 (N_8566,N_1223,N_40);
xnor U8567 (N_8567,N_1357,N_2298);
or U8568 (N_8568,N_574,N_2280);
or U8569 (N_8569,N_799,N_3019);
xnor U8570 (N_8570,N_1977,N_4365);
or U8571 (N_8571,N_611,N_607);
xor U8572 (N_8572,N_4012,N_2854);
xnor U8573 (N_8573,N_1834,N_3813);
xor U8574 (N_8574,N_2379,N_3071);
and U8575 (N_8575,N_525,N_974);
nor U8576 (N_8576,N_2179,N_1118);
nor U8577 (N_8577,N_4473,N_2416);
and U8578 (N_8578,N_2862,N_3277);
xor U8579 (N_8579,N_4019,N_2351);
or U8580 (N_8580,N_4049,N_1116);
nor U8581 (N_8581,N_2804,N_718);
and U8582 (N_8582,N_2785,N_2861);
and U8583 (N_8583,N_3297,N_2478);
nor U8584 (N_8584,N_2514,N_4828);
xor U8585 (N_8585,N_1427,N_2813);
and U8586 (N_8586,N_994,N_3105);
and U8587 (N_8587,N_2570,N_1341);
nand U8588 (N_8588,N_524,N_597);
nand U8589 (N_8589,N_3722,N_4048);
nand U8590 (N_8590,N_1243,N_3840);
and U8591 (N_8591,N_2984,N_2781);
xnor U8592 (N_8592,N_3929,N_4825);
xnor U8593 (N_8593,N_53,N_2455);
xor U8594 (N_8594,N_3878,N_769);
nand U8595 (N_8595,N_3789,N_2839);
and U8596 (N_8596,N_1947,N_3335);
nand U8597 (N_8597,N_4764,N_992);
nand U8598 (N_8598,N_148,N_3595);
or U8599 (N_8599,N_3471,N_1038);
xnor U8600 (N_8600,N_2408,N_537);
and U8601 (N_8601,N_1533,N_1884);
xnor U8602 (N_8602,N_3526,N_2178);
nor U8603 (N_8603,N_3188,N_2335);
nor U8604 (N_8604,N_815,N_921);
nand U8605 (N_8605,N_1698,N_27);
xor U8606 (N_8606,N_2469,N_697);
nand U8607 (N_8607,N_4532,N_2189);
and U8608 (N_8608,N_2910,N_1202);
or U8609 (N_8609,N_2754,N_2807);
nand U8610 (N_8610,N_4108,N_2267);
and U8611 (N_8611,N_2140,N_3568);
nor U8612 (N_8612,N_3807,N_1742);
xnor U8613 (N_8613,N_2746,N_3038);
or U8614 (N_8614,N_872,N_3964);
nor U8615 (N_8615,N_1783,N_946);
and U8616 (N_8616,N_1,N_4975);
xnor U8617 (N_8617,N_4891,N_2956);
or U8618 (N_8618,N_4317,N_1172);
and U8619 (N_8619,N_3531,N_4509);
and U8620 (N_8620,N_4801,N_629);
nand U8621 (N_8621,N_3064,N_4568);
or U8622 (N_8622,N_2723,N_4812);
xor U8623 (N_8623,N_3445,N_2485);
and U8624 (N_8624,N_2756,N_773);
and U8625 (N_8625,N_2437,N_969);
or U8626 (N_8626,N_3263,N_4103);
nor U8627 (N_8627,N_455,N_4502);
or U8628 (N_8628,N_1062,N_3855);
or U8629 (N_8629,N_2508,N_3980);
and U8630 (N_8630,N_733,N_1118);
xnor U8631 (N_8631,N_4935,N_1874);
nor U8632 (N_8632,N_516,N_1320);
nand U8633 (N_8633,N_3805,N_3002);
xnor U8634 (N_8634,N_3036,N_2498);
nand U8635 (N_8635,N_4008,N_4272);
and U8636 (N_8636,N_4097,N_3225);
nor U8637 (N_8637,N_4069,N_2105);
or U8638 (N_8638,N_4074,N_2098);
nor U8639 (N_8639,N_658,N_4437);
nand U8640 (N_8640,N_3108,N_1967);
nand U8641 (N_8641,N_3115,N_436);
nand U8642 (N_8642,N_2992,N_2347);
nand U8643 (N_8643,N_138,N_390);
and U8644 (N_8644,N_827,N_1426);
nand U8645 (N_8645,N_1846,N_1250);
nand U8646 (N_8646,N_1088,N_1494);
nand U8647 (N_8647,N_1008,N_4426);
nand U8648 (N_8648,N_4058,N_4198);
or U8649 (N_8649,N_1995,N_2447);
or U8650 (N_8650,N_4543,N_3686);
xor U8651 (N_8651,N_1001,N_3087);
and U8652 (N_8652,N_1499,N_2755);
or U8653 (N_8653,N_4898,N_3140);
and U8654 (N_8654,N_1579,N_1429);
xor U8655 (N_8655,N_679,N_4452);
xnor U8656 (N_8656,N_68,N_3187);
xnor U8657 (N_8657,N_1834,N_2976);
xnor U8658 (N_8658,N_751,N_2036);
xor U8659 (N_8659,N_1184,N_210);
nor U8660 (N_8660,N_4419,N_2044);
and U8661 (N_8661,N_879,N_1864);
nand U8662 (N_8662,N_4059,N_1447);
nand U8663 (N_8663,N_3007,N_2247);
and U8664 (N_8664,N_2379,N_80);
nand U8665 (N_8665,N_1312,N_2743);
nand U8666 (N_8666,N_28,N_1309);
nor U8667 (N_8667,N_764,N_3374);
nor U8668 (N_8668,N_4077,N_4733);
and U8669 (N_8669,N_2468,N_1953);
nand U8670 (N_8670,N_1555,N_4643);
nand U8671 (N_8671,N_4035,N_891);
xor U8672 (N_8672,N_2641,N_3373);
and U8673 (N_8673,N_2691,N_3080);
or U8674 (N_8674,N_3062,N_424);
or U8675 (N_8675,N_2229,N_1208);
or U8676 (N_8676,N_1105,N_1214);
nand U8677 (N_8677,N_768,N_3447);
nor U8678 (N_8678,N_2509,N_1246);
xnor U8679 (N_8679,N_2210,N_631);
nor U8680 (N_8680,N_4866,N_3748);
xnor U8681 (N_8681,N_2249,N_2439);
nor U8682 (N_8682,N_4181,N_2797);
or U8683 (N_8683,N_4709,N_2785);
and U8684 (N_8684,N_1873,N_4443);
xor U8685 (N_8685,N_734,N_3602);
and U8686 (N_8686,N_2316,N_2412);
and U8687 (N_8687,N_2415,N_3553);
and U8688 (N_8688,N_700,N_3365);
xor U8689 (N_8689,N_1597,N_1505);
xor U8690 (N_8690,N_2915,N_1478);
and U8691 (N_8691,N_2157,N_349);
or U8692 (N_8692,N_3967,N_3815);
nor U8693 (N_8693,N_1805,N_4581);
nand U8694 (N_8694,N_536,N_1273);
nand U8695 (N_8695,N_4341,N_2213);
nand U8696 (N_8696,N_3746,N_3795);
nor U8697 (N_8697,N_4927,N_1181);
and U8698 (N_8698,N_1379,N_1667);
nor U8699 (N_8699,N_4831,N_266);
nand U8700 (N_8700,N_639,N_1850);
nor U8701 (N_8701,N_688,N_795);
xnor U8702 (N_8702,N_2352,N_3105);
or U8703 (N_8703,N_3074,N_1407);
xor U8704 (N_8704,N_3979,N_711);
xnor U8705 (N_8705,N_1727,N_1969);
xor U8706 (N_8706,N_1040,N_2260);
nor U8707 (N_8707,N_849,N_3268);
xnor U8708 (N_8708,N_2216,N_4992);
xor U8709 (N_8709,N_4976,N_965);
nand U8710 (N_8710,N_717,N_4172);
nand U8711 (N_8711,N_4915,N_3336);
nor U8712 (N_8712,N_4423,N_239);
nor U8713 (N_8713,N_4858,N_3785);
nor U8714 (N_8714,N_3302,N_1445);
and U8715 (N_8715,N_3576,N_4660);
or U8716 (N_8716,N_522,N_3137);
nand U8717 (N_8717,N_4427,N_2073);
nand U8718 (N_8718,N_403,N_3016);
xor U8719 (N_8719,N_955,N_353);
nor U8720 (N_8720,N_4603,N_4337);
or U8721 (N_8721,N_785,N_1072);
nand U8722 (N_8722,N_4240,N_4203);
nor U8723 (N_8723,N_4050,N_2471);
nand U8724 (N_8724,N_240,N_1895);
nor U8725 (N_8725,N_281,N_248);
and U8726 (N_8726,N_1565,N_2784);
or U8727 (N_8727,N_2331,N_1872);
xor U8728 (N_8728,N_1182,N_1285);
xor U8729 (N_8729,N_1605,N_2819);
or U8730 (N_8730,N_1056,N_2097);
nand U8731 (N_8731,N_4578,N_707);
nand U8732 (N_8732,N_4713,N_134);
nand U8733 (N_8733,N_2306,N_2435);
xnor U8734 (N_8734,N_2469,N_3220);
and U8735 (N_8735,N_81,N_26);
nor U8736 (N_8736,N_4791,N_1724);
nor U8737 (N_8737,N_183,N_2128);
nor U8738 (N_8738,N_2338,N_2645);
or U8739 (N_8739,N_622,N_967);
and U8740 (N_8740,N_3926,N_3822);
or U8741 (N_8741,N_4429,N_4265);
nor U8742 (N_8742,N_400,N_3999);
xor U8743 (N_8743,N_1324,N_3251);
and U8744 (N_8744,N_636,N_1664);
nand U8745 (N_8745,N_4812,N_1022);
or U8746 (N_8746,N_4625,N_4073);
or U8747 (N_8747,N_731,N_1178);
or U8748 (N_8748,N_4849,N_2149);
nand U8749 (N_8749,N_3987,N_1743);
and U8750 (N_8750,N_4511,N_1352);
or U8751 (N_8751,N_2689,N_1850);
xnor U8752 (N_8752,N_3772,N_3640);
and U8753 (N_8753,N_222,N_2041);
nor U8754 (N_8754,N_2676,N_3860);
or U8755 (N_8755,N_939,N_4065);
and U8756 (N_8756,N_1528,N_1898);
xnor U8757 (N_8757,N_255,N_3075);
nor U8758 (N_8758,N_2709,N_3131);
nor U8759 (N_8759,N_3138,N_418);
nor U8760 (N_8760,N_1511,N_3481);
or U8761 (N_8761,N_1860,N_1735);
and U8762 (N_8762,N_1689,N_2846);
nor U8763 (N_8763,N_1200,N_3923);
nor U8764 (N_8764,N_1952,N_1848);
nor U8765 (N_8765,N_2759,N_1627);
xor U8766 (N_8766,N_3747,N_936);
xnor U8767 (N_8767,N_2011,N_693);
nand U8768 (N_8768,N_2640,N_2692);
nor U8769 (N_8769,N_377,N_4083);
xor U8770 (N_8770,N_4772,N_1657);
or U8771 (N_8771,N_3459,N_2084);
or U8772 (N_8772,N_436,N_3665);
xnor U8773 (N_8773,N_2314,N_3654);
and U8774 (N_8774,N_3997,N_1747);
nor U8775 (N_8775,N_2434,N_808);
or U8776 (N_8776,N_2344,N_2318);
nor U8777 (N_8777,N_1038,N_2022);
xor U8778 (N_8778,N_2825,N_1941);
nand U8779 (N_8779,N_1284,N_2396);
xor U8780 (N_8780,N_3672,N_3223);
and U8781 (N_8781,N_3704,N_1980);
xnor U8782 (N_8782,N_3547,N_4901);
or U8783 (N_8783,N_541,N_258);
and U8784 (N_8784,N_186,N_3860);
nand U8785 (N_8785,N_4007,N_1575);
nand U8786 (N_8786,N_518,N_3006);
nor U8787 (N_8787,N_3964,N_4976);
or U8788 (N_8788,N_3935,N_1290);
and U8789 (N_8789,N_1584,N_313);
xnor U8790 (N_8790,N_3757,N_246);
nor U8791 (N_8791,N_4889,N_3634);
and U8792 (N_8792,N_1017,N_2757);
nor U8793 (N_8793,N_4458,N_340);
xor U8794 (N_8794,N_1739,N_3995);
or U8795 (N_8795,N_3834,N_799);
or U8796 (N_8796,N_1416,N_4304);
xnor U8797 (N_8797,N_2063,N_4900);
and U8798 (N_8798,N_65,N_2992);
or U8799 (N_8799,N_3090,N_4023);
nand U8800 (N_8800,N_3321,N_4148);
or U8801 (N_8801,N_1414,N_3023);
nand U8802 (N_8802,N_786,N_1618);
or U8803 (N_8803,N_2445,N_3628);
xor U8804 (N_8804,N_1133,N_3999);
nor U8805 (N_8805,N_2976,N_2163);
nand U8806 (N_8806,N_3188,N_1913);
or U8807 (N_8807,N_661,N_3544);
or U8808 (N_8808,N_987,N_3672);
or U8809 (N_8809,N_1779,N_362);
and U8810 (N_8810,N_1351,N_4246);
nor U8811 (N_8811,N_436,N_3496);
or U8812 (N_8812,N_3408,N_625);
and U8813 (N_8813,N_2290,N_3072);
nor U8814 (N_8814,N_325,N_2712);
nor U8815 (N_8815,N_2882,N_1798);
nor U8816 (N_8816,N_165,N_2613);
or U8817 (N_8817,N_528,N_4106);
or U8818 (N_8818,N_748,N_4012);
and U8819 (N_8819,N_4133,N_2839);
nand U8820 (N_8820,N_129,N_1077);
and U8821 (N_8821,N_3355,N_2301);
nor U8822 (N_8822,N_423,N_2082);
xnor U8823 (N_8823,N_2499,N_3523);
nand U8824 (N_8824,N_3190,N_4704);
or U8825 (N_8825,N_3594,N_1781);
nand U8826 (N_8826,N_4799,N_570);
nand U8827 (N_8827,N_690,N_4714);
xor U8828 (N_8828,N_3478,N_4238);
and U8829 (N_8829,N_3877,N_2650);
xor U8830 (N_8830,N_1408,N_3467);
and U8831 (N_8831,N_567,N_2511);
nor U8832 (N_8832,N_2049,N_3283);
nor U8833 (N_8833,N_2644,N_4754);
and U8834 (N_8834,N_3425,N_2564);
xnor U8835 (N_8835,N_2039,N_105);
nand U8836 (N_8836,N_3226,N_4917);
nor U8837 (N_8837,N_2743,N_651);
and U8838 (N_8838,N_1810,N_849);
or U8839 (N_8839,N_1742,N_2598);
xnor U8840 (N_8840,N_311,N_1803);
and U8841 (N_8841,N_3245,N_1913);
nand U8842 (N_8842,N_3585,N_3845);
nor U8843 (N_8843,N_3347,N_4352);
and U8844 (N_8844,N_3464,N_4782);
or U8845 (N_8845,N_1905,N_2533);
or U8846 (N_8846,N_324,N_1524);
and U8847 (N_8847,N_408,N_1537);
nand U8848 (N_8848,N_4502,N_2931);
and U8849 (N_8849,N_1527,N_3006);
nor U8850 (N_8850,N_3469,N_1494);
nand U8851 (N_8851,N_2991,N_1922);
or U8852 (N_8852,N_3524,N_1986);
nor U8853 (N_8853,N_3752,N_2874);
and U8854 (N_8854,N_4064,N_1613);
and U8855 (N_8855,N_4475,N_1756);
xor U8856 (N_8856,N_3842,N_664);
nor U8857 (N_8857,N_1792,N_4046);
nor U8858 (N_8858,N_3512,N_1917);
and U8859 (N_8859,N_1731,N_4745);
xor U8860 (N_8860,N_67,N_3688);
xor U8861 (N_8861,N_3279,N_3010);
and U8862 (N_8862,N_3918,N_3603);
nor U8863 (N_8863,N_2265,N_48);
nor U8864 (N_8864,N_1516,N_3685);
xor U8865 (N_8865,N_2454,N_195);
nand U8866 (N_8866,N_1253,N_3309);
nor U8867 (N_8867,N_4832,N_4442);
or U8868 (N_8868,N_2923,N_903);
or U8869 (N_8869,N_231,N_2215);
and U8870 (N_8870,N_3784,N_31);
and U8871 (N_8871,N_1624,N_755);
and U8872 (N_8872,N_674,N_4615);
xor U8873 (N_8873,N_2697,N_3590);
nor U8874 (N_8874,N_772,N_746);
xor U8875 (N_8875,N_1944,N_3613);
xnor U8876 (N_8876,N_3375,N_4981);
nand U8877 (N_8877,N_3590,N_2499);
nor U8878 (N_8878,N_1910,N_343);
nand U8879 (N_8879,N_165,N_2853);
nand U8880 (N_8880,N_581,N_4487);
xor U8881 (N_8881,N_3201,N_4237);
xnor U8882 (N_8882,N_4030,N_2607);
and U8883 (N_8883,N_635,N_935);
nor U8884 (N_8884,N_2471,N_2587);
or U8885 (N_8885,N_2692,N_1432);
or U8886 (N_8886,N_1536,N_83);
nor U8887 (N_8887,N_3013,N_2394);
or U8888 (N_8888,N_2993,N_4050);
nand U8889 (N_8889,N_362,N_714);
nor U8890 (N_8890,N_3685,N_2106);
or U8891 (N_8891,N_2075,N_362);
nor U8892 (N_8892,N_4520,N_1307);
xor U8893 (N_8893,N_3943,N_702);
xor U8894 (N_8894,N_4876,N_3569);
or U8895 (N_8895,N_118,N_4689);
xor U8896 (N_8896,N_450,N_558);
nor U8897 (N_8897,N_1196,N_4031);
or U8898 (N_8898,N_532,N_2153);
or U8899 (N_8899,N_1481,N_2597);
and U8900 (N_8900,N_546,N_2395);
xnor U8901 (N_8901,N_2983,N_1059);
nand U8902 (N_8902,N_574,N_1282);
and U8903 (N_8903,N_632,N_4326);
or U8904 (N_8904,N_2594,N_4333);
and U8905 (N_8905,N_3507,N_529);
nor U8906 (N_8906,N_742,N_4414);
and U8907 (N_8907,N_2627,N_772);
and U8908 (N_8908,N_1622,N_3656);
nand U8909 (N_8909,N_3175,N_2244);
xor U8910 (N_8910,N_694,N_2804);
nor U8911 (N_8911,N_4650,N_1859);
nand U8912 (N_8912,N_2496,N_1946);
nor U8913 (N_8913,N_734,N_2715);
nand U8914 (N_8914,N_2732,N_2566);
xnor U8915 (N_8915,N_1984,N_703);
nor U8916 (N_8916,N_3673,N_4364);
or U8917 (N_8917,N_3885,N_2307);
nand U8918 (N_8918,N_1990,N_3021);
or U8919 (N_8919,N_524,N_2248);
xor U8920 (N_8920,N_3957,N_1549);
or U8921 (N_8921,N_1131,N_868);
xnor U8922 (N_8922,N_617,N_1318);
or U8923 (N_8923,N_4629,N_3728);
nor U8924 (N_8924,N_161,N_2078);
nor U8925 (N_8925,N_4180,N_310);
or U8926 (N_8926,N_667,N_3292);
nand U8927 (N_8927,N_4491,N_180);
or U8928 (N_8928,N_4137,N_4235);
and U8929 (N_8929,N_977,N_3677);
xnor U8930 (N_8930,N_402,N_4380);
nand U8931 (N_8931,N_684,N_2246);
xor U8932 (N_8932,N_986,N_346);
and U8933 (N_8933,N_3476,N_1006);
nor U8934 (N_8934,N_1573,N_381);
or U8935 (N_8935,N_577,N_585);
or U8936 (N_8936,N_1444,N_3718);
nand U8937 (N_8937,N_4944,N_529);
nand U8938 (N_8938,N_3910,N_1005);
or U8939 (N_8939,N_394,N_4502);
nand U8940 (N_8940,N_3980,N_2777);
nor U8941 (N_8941,N_4485,N_1583);
or U8942 (N_8942,N_2990,N_3945);
nand U8943 (N_8943,N_3875,N_3547);
and U8944 (N_8944,N_1486,N_4542);
nand U8945 (N_8945,N_4847,N_4268);
xnor U8946 (N_8946,N_1555,N_2497);
nor U8947 (N_8947,N_3458,N_1081);
and U8948 (N_8948,N_3232,N_259);
nand U8949 (N_8949,N_3232,N_990);
nand U8950 (N_8950,N_2886,N_2390);
and U8951 (N_8951,N_1208,N_2713);
or U8952 (N_8952,N_1250,N_3765);
xor U8953 (N_8953,N_193,N_4393);
or U8954 (N_8954,N_2308,N_43);
nor U8955 (N_8955,N_2941,N_673);
or U8956 (N_8956,N_183,N_3149);
nor U8957 (N_8957,N_3503,N_3631);
nand U8958 (N_8958,N_3649,N_4005);
xor U8959 (N_8959,N_4999,N_4088);
xor U8960 (N_8960,N_215,N_421);
nand U8961 (N_8961,N_3529,N_148);
nand U8962 (N_8962,N_1532,N_3465);
and U8963 (N_8963,N_1714,N_534);
nor U8964 (N_8964,N_1584,N_413);
or U8965 (N_8965,N_168,N_1028);
nor U8966 (N_8966,N_1981,N_4688);
nand U8967 (N_8967,N_1786,N_3585);
or U8968 (N_8968,N_813,N_1267);
nor U8969 (N_8969,N_2610,N_1563);
nor U8970 (N_8970,N_2296,N_4252);
or U8971 (N_8971,N_454,N_725);
nor U8972 (N_8972,N_1415,N_2955);
nand U8973 (N_8973,N_3305,N_714);
xnor U8974 (N_8974,N_207,N_4827);
nor U8975 (N_8975,N_3547,N_600);
nor U8976 (N_8976,N_3335,N_835);
or U8977 (N_8977,N_4256,N_4092);
nand U8978 (N_8978,N_33,N_2303);
xnor U8979 (N_8979,N_1406,N_3531);
or U8980 (N_8980,N_4753,N_905);
xor U8981 (N_8981,N_2607,N_4109);
and U8982 (N_8982,N_1161,N_3029);
nor U8983 (N_8983,N_383,N_3339);
or U8984 (N_8984,N_3900,N_4385);
and U8985 (N_8985,N_4617,N_3884);
nor U8986 (N_8986,N_2578,N_1071);
and U8987 (N_8987,N_694,N_3747);
nand U8988 (N_8988,N_371,N_3444);
nor U8989 (N_8989,N_2568,N_1462);
xor U8990 (N_8990,N_2663,N_3317);
xor U8991 (N_8991,N_958,N_3128);
nor U8992 (N_8992,N_2325,N_3332);
nor U8993 (N_8993,N_1122,N_4117);
and U8994 (N_8994,N_3402,N_57);
and U8995 (N_8995,N_1333,N_2610);
xor U8996 (N_8996,N_4723,N_3692);
or U8997 (N_8997,N_2861,N_1532);
nand U8998 (N_8998,N_625,N_2836);
nand U8999 (N_8999,N_143,N_4209);
xor U9000 (N_9000,N_2126,N_3571);
xnor U9001 (N_9001,N_3481,N_3278);
xnor U9002 (N_9002,N_3941,N_2390);
nand U9003 (N_9003,N_4417,N_2058);
and U9004 (N_9004,N_4106,N_803);
or U9005 (N_9005,N_1261,N_574);
xor U9006 (N_9006,N_4133,N_1405);
xnor U9007 (N_9007,N_1752,N_3042);
and U9008 (N_9008,N_4955,N_1919);
nor U9009 (N_9009,N_2741,N_2483);
xnor U9010 (N_9010,N_4854,N_959);
nor U9011 (N_9011,N_2853,N_3512);
and U9012 (N_9012,N_1976,N_576);
nand U9013 (N_9013,N_268,N_3945);
or U9014 (N_9014,N_4887,N_2826);
xnor U9015 (N_9015,N_3329,N_685);
xor U9016 (N_9016,N_714,N_3916);
xor U9017 (N_9017,N_2519,N_1768);
xor U9018 (N_9018,N_3350,N_2889);
xnor U9019 (N_9019,N_3802,N_899);
nor U9020 (N_9020,N_2437,N_1563);
or U9021 (N_9021,N_2088,N_4574);
nand U9022 (N_9022,N_3412,N_1198);
or U9023 (N_9023,N_1180,N_1628);
and U9024 (N_9024,N_3294,N_4295);
nor U9025 (N_9025,N_4863,N_3331);
and U9026 (N_9026,N_2605,N_4252);
nor U9027 (N_9027,N_3952,N_1179);
xnor U9028 (N_9028,N_2630,N_3132);
nand U9029 (N_9029,N_624,N_2876);
nor U9030 (N_9030,N_4444,N_2752);
nand U9031 (N_9031,N_788,N_2623);
and U9032 (N_9032,N_2280,N_1396);
and U9033 (N_9033,N_4270,N_3043);
nand U9034 (N_9034,N_2726,N_1065);
and U9035 (N_9035,N_1949,N_4480);
or U9036 (N_9036,N_1413,N_4260);
xnor U9037 (N_9037,N_3020,N_1317);
nand U9038 (N_9038,N_288,N_2720);
nor U9039 (N_9039,N_3451,N_4682);
nand U9040 (N_9040,N_2549,N_3952);
xor U9041 (N_9041,N_4362,N_659);
xor U9042 (N_9042,N_4386,N_4510);
or U9043 (N_9043,N_4294,N_2119);
and U9044 (N_9044,N_4458,N_3418);
nor U9045 (N_9045,N_2669,N_4108);
or U9046 (N_9046,N_4200,N_143);
nor U9047 (N_9047,N_2675,N_146);
nor U9048 (N_9048,N_175,N_2263);
nor U9049 (N_9049,N_70,N_2924);
and U9050 (N_9050,N_816,N_620);
xor U9051 (N_9051,N_761,N_562);
nor U9052 (N_9052,N_2488,N_4889);
nand U9053 (N_9053,N_1295,N_61);
and U9054 (N_9054,N_2544,N_1752);
or U9055 (N_9055,N_3690,N_3502);
and U9056 (N_9056,N_2432,N_2624);
xnor U9057 (N_9057,N_340,N_228);
xnor U9058 (N_9058,N_4762,N_3882);
and U9059 (N_9059,N_1479,N_1913);
xor U9060 (N_9060,N_1557,N_2696);
nand U9061 (N_9061,N_3717,N_1635);
nor U9062 (N_9062,N_2338,N_1088);
or U9063 (N_9063,N_4689,N_855);
nor U9064 (N_9064,N_3814,N_4037);
xor U9065 (N_9065,N_4577,N_2551);
xor U9066 (N_9066,N_4001,N_585);
nor U9067 (N_9067,N_3410,N_2724);
or U9068 (N_9068,N_3440,N_4856);
or U9069 (N_9069,N_3395,N_4262);
or U9070 (N_9070,N_4950,N_724);
and U9071 (N_9071,N_305,N_705);
or U9072 (N_9072,N_1246,N_1213);
nand U9073 (N_9073,N_3955,N_1061);
nand U9074 (N_9074,N_2666,N_2122);
xor U9075 (N_9075,N_2562,N_1403);
nand U9076 (N_9076,N_3398,N_3548);
nor U9077 (N_9077,N_1664,N_1877);
nand U9078 (N_9078,N_2516,N_4873);
nand U9079 (N_9079,N_2348,N_775);
or U9080 (N_9080,N_754,N_3261);
and U9081 (N_9081,N_4814,N_1587);
xnor U9082 (N_9082,N_563,N_2865);
nor U9083 (N_9083,N_4752,N_4571);
nor U9084 (N_9084,N_4007,N_275);
nor U9085 (N_9085,N_2564,N_3225);
xor U9086 (N_9086,N_2268,N_4743);
or U9087 (N_9087,N_4451,N_4324);
or U9088 (N_9088,N_1090,N_27);
nand U9089 (N_9089,N_1932,N_3687);
xor U9090 (N_9090,N_2431,N_2423);
nor U9091 (N_9091,N_3303,N_3204);
nor U9092 (N_9092,N_3391,N_4964);
and U9093 (N_9093,N_2337,N_1293);
nor U9094 (N_9094,N_1032,N_2841);
or U9095 (N_9095,N_154,N_655);
nand U9096 (N_9096,N_2360,N_1029);
xor U9097 (N_9097,N_265,N_4021);
nor U9098 (N_9098,N_3542,N_264);
and U9099 (N_9099,N_1841,N_1210);
nor U9100 (N_9100,N_3752,N_1621);
nand U9101 (N_9101,N_3156,N_4380);
xor U9102 (N_9102,N_1088,N_3143);
and U9103 (N_9103,N_2063,N_4541);
and U9104 (N_9104,N_2908,N_2195);
nor U9105 (N_9105,N_4672,N_3669);
nor U9106 (N_9106,N_2896,N_4229);
and U9107 (N_9107,N_646,N_4672);
xor U9108 (N_9108,N_387,N_3153);
and U9109 (N_9109,N_3305,N_1005);
xnor U9110 (N_9110,N_157,N_4250);
and U9111 (N_9111,N_4007,N_2458);
nand U9112 (N_9112,N_4648,N_765);
and U9113 (N_9113,N_1673,N_3632);
or U9114 (N_9114,N_2907,N_1945);
nor U9115 (N_9115,N_2760,N_4794);
xnor U9116 (N_9116,N_123,N_2277);
nor U9117 (N_9117,N_3517,N_3701);
nand U9118 (N_9118,N_3967,N_4200);
nor U9119 (N_9119,N_4758,N_4978);
nor U9120 (N_9120,N_3784,N_2499);
xnor U9121 (N_9121,N_1967,N_1473);
nor U9122 (N_9122,N_4502,N_2067);
xnor U9123 (N_9123,N_4472,N_3003);
nor U9124 (N_9124,N_494,N_3448);
xnor U9125 (N_9125,N_2850,N_1070);
or U9126 (N_9126,N_636,N_4815);
nor U9127 (N_9127,N_1328,N_4765);
xor U9128 (N_9128,N_1007,N_580);
nor U9129 (N_9129,N_3158,N_98);
nand U9130 (N_9130,N_3163,N_3004);
and U9131 (N_9131,N_2358,N_82);
or U9132 (N_9132,N_1441,N_4205);
xor U9133 (N_9133,N_1386,N_283);
or U9134 (N_9134,N_2116,N_3416);
xor U9135 (N_9135,N_2407,N_1802);
or U9136 (N_9136,N_3682,N_1080);
nor U9137 (N_9137,N_1656,N_4169);
and U9138 (N_9138,N_4787,N_1075);
and U9139 (N_9139,N_2997,N_3122);
nor U9140 (N_9140,N_2612,N_1326);
nand U9141 (N_9141,N_1375,N_1688);
or U9142 (N_9142,N_4021,N_405);
or U9143 (N_9143,N_1498,N_1832);
nor U9144 (N_9144,N_3756,N_4347);
nor U9145 (N_9145,N_1375,N_3933);
and U9146 (N_9146,N_1699,N_4409);
nand U9147 (N_9147,N_4839,N_8);
nor U9148 (N_9148,N_1946,N_4967);
nor U9149 (N_9149,N_3947,N_1914);
nor U9150 (N_9150,N_2932,N_3879);
xnor U9151 (N_9151,N_3195,N_2449);
or U9152 (N_9152,N_1972,N_772);
and U9153 (N_9153,N_2140,N_2209);
and U9154 (N_9154,N_494,N_4006);
nand U9155 (N_9155,N_2209,N_4562);
or U9156 (N_9156,N_2679,N_435);
nand U9157 (N_9157,N_999,N_1619);
or U9158 (N_9158,N_4660,N_2923);
xor U9159 (N_9159,N_1364,N_1274);
and U9160 (N_9160,N_1325,N_1993);
xnor U9161 (N_9161,N_967,N_267);
or U9162 (N_9162,N_4247,N_1526);
nor U9163 (N_9163,N_1823,N_315);
or U9164 (N_9164,N_3316,N_520);
or U9165 (N_9165,N_1599,N_938);
and U9166 (N_9166,N_4459,N_1266);
nand U9167 (N_9167,N_802,N_2465);
and U9168 (N_9168,N_2454,N_3629);
nor U9169 (N_9169,N_4343,N_504);
nor U9170 (N_9170,N_2746,N_235);
and U9171 (N_9171,N_1175,N_1535);
nor U9172 (N_9172,N_2291,N_1748);
and U9173 (N_9173,N_787,N_1416);
nor U9174 (N_9174,N_2680,N_443);
or U9175 (N_9175,N_1574,N_4518);
nand U9176 (N_9176,N_543,N_20);
nor U9177 (N_9177,N_4355,N_2271);
or U9178 (N_9178,N_3490,N_4949);
xor U9179 (N_9179,N_3187,N_3182);
and U9180 (N_9180,N_3979,N_2768);
nor U9181 (N_9181,N_3821,N_1311);
nor U9182 (N_9182,N_2025,N_3731);
nand U9183 (N_9183,N_244,N_3728);
xnor U9184 (N_9184,N_4950,N_4348);
xnor U9185 (N_9185,N_2511,N_113);
or U9186 (N_9186,N_840,N_3822);
nor U9187 (N_9187,N_2515,N_3927);
nand U9188 (N_9188,N_348,N_3208);
and U9189 (N_9189,N_2515,N_3296);
nor U9190 (N_9190,N_1551,N_4040);
or U9191 (N_9191,N_3267,N_3909);
xor U9192 (N_9192,N_3510,N_2482);
nor U9193 (N_9193,N_1423,N_4078);
or U9194 (N_9194,N_3332,N_4343);
nor U9195 (N_9195,N_3198,N_2257);
or U9196 (N_9196,N_3890,N_794);
or U9197 (N_9197,N_2378,N_1174);
and U9198 (N_9198,N_798,N_3296);
nor U9199 (N_9199,N_4275,N_51);
xnor U9200 (N_9200,N_3450,N_451);
xnor U9201 (N_9201,N_897,N_4130);
and U9202 (N_9202,N_1988,N_3831);
nor U9203 (N_9203,N_1136,N_968);
xnor U9204 (N_9204,N_4141,N_2773);
nor U9205 (N_9205,N_2356,N_2632);
nand U9206 (N_9206,N_4289,N_1083);
nand U9207 (N_9207,N_3746,N_525);
nand U9208 (N_9208,N_726,N_603);
xor U9209 (N_9209,N_3223,N_4385);
xor U9210 (N_9210,N_98,N_3053);
nand U9211 (N_9211,N_4767,N_2411);
and U9212 (N_9212,N_3326,N_4700);
and U9213 (N_9213,N_1056,N_1812);
xnor U9214 (N_9214,N_334,N_1677);
nand U9215 (N_9215,N_677,N_1499);
or U9216 (N_9216,N_3684,N_3917);
nor U9217 (N_9217,N_490,N_2189);
or U9218 (N_9218,N_3621,N_4070);
nand U9219 (N_9219,N_2425,N_4836);
xor U9220 (N_9220,N_2533,N_4744);
nand U9221 (N_9221,N_3984,N_1757);
nor U9222 (N_9222,N_1981,N_3124);
xnor U9223 (N_9223,N_2201,N_2719);
or U9224 (N_9224,N_2567,N_4101);
xor U9225 (N_9225,N_719,N_2730);
nand U9226 (N_9226,N_1527,N_3042);
and U9227 (N_9227,N_1646,N_3603);
and U9228 (N_9228,N_4814,N_4739);
nor U9229 (N_9229,N_4562,N_3523);
nor U9230 (N_9230,N_2159,N_857);
xnor U9231 (N_9231,N_2920,N_693);
nand U9232 (N_9232,N_3370,N_2759);
nor U9233 (N_9233,N_142,N_3925);
nor U9234 (N_9234,N_3649,N_2822);
or U9235 (N_9235,N_3966,N_187);
nand U9236 (N_9236,N_1504,N_269);
nor U9237 (N_9237,N_2943,N_4058);
or U9238 (N_9238,N_1098,N_4643);
xnor U9239 (N_9239,N_172,N_1482);
nor U9240 (N_9240,N_4156,N_2925);
xor U9241 (N_9241,N_2772,N_1063);
nand U9242 (N_9242,N_4360,N_3213);
xnor U9243 (N_9243,N_3938,N_4214);
nor U9244 (N_9244,N_1006,N_1101);
nand U9245 (N_9245,N_115,N_4409);
nand U9246 (N_9246,N_1821,N_337);
and U9247 (N_9247,N_4583,N_905);
or U9248 (N_9248,N_4568,N_487);
xnor U9249 (N_9249,N_587,N_756);
nor U9250 (N_9250,N_1694,N_3632);
or U9251 (N_9251,N_742,N_547);
or U9252 (N_9252,N_3047,N_4381);
nand U9253 (N_9253,N_3153,N_2224);
nor U9254 (N_9254,N_1694,N_1175);
or U9255 (N_9255,N_14,N_4619);
nand U9256 (N_9256,N_3900,N_2051);
or U9257 (N_9257,N_770,N_1044);
nor U9258 (N_9258,N_352,N_3055);
xor U9259 (N_9259,N_2176,N_3486);
and U9260 (N_9260,N_3802,N_560);
or U9261 (N_9261,N_4463,N_3700);
xor U9262 (N_9262,N_4345,N_635);
and U9263 (N_9263,N_103,N_2913);
nand U9264 (N_9264,N_3328,N_1344);
xor U9265 (N_9265,N_4090,N_664);
xnor U9266 (N_9266,N_3801,N_1604);
nor U9267 (N_9267,N_2618,N_72);
xnor U9268 (N_9268,N_3150,N_3278);
and U9269 (N_9269,N_2211,N_961);
and U9270 (N_9270,N_728,N_2099);
nor U9271 (N_9271,N_4577,N_3444);
xnor U9272 (N_9272,N_2291,N_1597);
xnor U9273 (N_9273,N_3324,N_3168);
xor U9274 (N_9274,N_925,N_1912);
nand U9275 (N_9275,N_562,N_3398);
nand U9276 (N_9276,N_3672,N_3937);
nand U9277 (N_9277,N_3473,N_562);
and U9278 (N_9278,N_4635,N_3818);
nor U9279 (N_9279,N_1484,N_3863);
and U9280 (N_9280,N_4208,N_1990);
nand U9281 (N_9281,N_1542,N_312);
or U9282 (N_9282,N_3057,N_4740);
nand U9283 (N_9283,N_1598,N_4213);
and U9284 (N_9284,N_3195,N_1366);
nand U9285 (N_9285,N_664,N_1094);
xnor U9286 (N_9286,N_2064,N_1227);
xnor U9287 (N_9287,N_232,N_1457);
or U9288 (N_9288,N_3481,N_111);
or U9289 (N_9289,N_804,N_1413);
xnor U9290 (N_9290,N_2628,N_2896);
or U9291 (N_9291,N_4101,N_3400);
nor U9292 (N_9292,N_206,N_3100);
nor U9293 (N_9293,N_2324,N_4882);
nand U9294 (N_9294,N_1320,N_737);
or U9295 (N_9295,N_4555,N_3261);
nor U9296 (N_9296,N_2427,N_470);
nor U9297 (N_9297,N_2940,N_1103);
or U9298 (N_9298,N_1491,N_265);
or U9299 (N_9299,N_4890,N_3834);
xnor U9300 (N_9300,N_1069,N_878);
nand U9301 (N_9301,N_68,N_3537);
and U9302 (N_9302,N_137,N_363);
nand U9303 (N_9303,N_1747,N_1758);
and U9304 (N_9304,N_3528,N_1879);
nand U9305 (N_9305,N_150,N_584);
and U9306 (N_9306,N_1364,N_1101);
and U9307 (N_9307,N_4102,N_276);
nor U9308 (N_9308,N_4488,N_3718);
nand U9309 (N_9309,N_3690,N_3150);
and U9310 (N_9310,N_3769,N_4157);
xor U9311 (N_9311,N_1053,N_1877);
xnor U9312 (N_9312,N_1975,N_4249);
xor U9313 (N_9313,N_818,N_2769);
and U9314 (N_9314,N_2680,N_3715);
or U9315 (N_9315,N_815,N_716);
or U9316 (N_9316,N_213,N_2093);
and U9317 (N_9317,N_2798,N_1832);
xnor U9318 (N_9318,N_2364,N_896);
nor U9319 (N_9319,N_3937,N_1607);
nand U9320 (N_9320,N_413,N_3782);
nand U9321 (N_9321,N_2654,N_2276);
and U9322 (N_9322,N_4020,N_200);
xnor U9323 (N_9323,N_4356,N_2676);
nand U9324 (N_9324,N_2868,N_3569);
and U9325 (N_9325,N_3725,N_126);
xor U9326 (N_9326,N_1736,N_4129);
and U9327 (N_9327,N_3926,N_2449);
xnor U9328 (N_9328,N_3482,N_139);
nand U9329 (N_9329,N_242,N_462);
nand U9330 (N_9330,N_364,N_1939);
and U9331 (N_9331,N_4426,N_797);
or U9332 (N_9332,N_701,N_1246);
xor U9333 (N_9333,N_2143,N_3848);
xnor U9334 (N_9334,N_1794,N_4037);
and U9335 (N_9335,N_2409,N_1565);
xnor U9336 (N_9336,N_2413,N_4766);
xor U9337 (N_9337,N_1695,N_2253);
and U9338 (N_9338,N_77,N_2141);
nand U9339 (N_9339,N_2726,N_138);
and U9340 (N_9340,N_3119,N_1436);
nand U9341 (N_9341,N_4935,N_1829);
nand U9342 (N_9342,N_472,N_4861);
xor U9343 (N_9343,N_3223,N_3790);
and U9344 (N_9344,N_1726,N_3904);
and U9345 (N_9345,N_1105,N_561);
and U9346 (N_9346,N_2401,N_4472);
or U9347 (N_9347,N_4343,N_3464);
and U9348 (N_9348,N_2508,N_232);
xnor U9349 (N_9349,N_546,N_4910);
xor U9350 (N_9350,N_873,N_2155);
xnor U9351 (N_9351,N_2573,N_926);
or U9352 (N_9352,N_1964,N_2202);
xnor U9353 (N_9353,N_168,N_3893);
and U9354 (N_9354,N_339,N_4478);
or U9355 (N_9355,N_3147,N_3506);
xor U9356 (N_9356,N_2476,N_780);
nor U9357 (N_9357,N_461,N_521);
and U9358 (N_9358,N_2407,N_467);
nand U9359 (N_9359,N_3524,N_4198);
nand U9360 (N_9360,N_302,N_3413);
nand U9361 (N_9361,N_4313,N_1316);
nor U9362 (N_9362,N_1408,N_4511);
xnor U9363 (N_9363,N_2070,N_1873);
nand U9364 (N_9364,N_3141,N_3492);
and U9365 (N_9365,N_2730,N_854);
xnor U9366 (N_9366,N_3256,N_1136);
and U9367 (N_9367,N_2289,N_4267);
xor U9368 (N_9368,N_799,N_4754);
nor U9369 (N_9369,N_2630,N_3799);
nor U9370 (N_9370,N_4765,N_3283);
nor U9371 (N_9371,N_1570,N_3001);
nand U9372 (N_9372,N_4099,N_3033);
xnor U9373 (N_9373,N_3780,N_1499);
or U9374 (N_9374,N_5,N_3972);
nor U9375 (N_9375,N_4302,N_3734);
nor U9376 (N_9376,N_1522,N_3088);
or U9377 (N_9377,N_3135,N_362);
xor U9378 (N_9378,N_3628,N_2485);
nand U9379 (N_9379,N_1169,N_3696);
or U9380 (N_9380,N_4556,N_1775);
xor U9381 (N_9381,N_1458,N_2294);
and U9382 (N_9382,N_3523,N_2073);
nand U9383 (N_9383,N_4839,N_3340);
xor U9384 (N_9384,N_3974,N_767);
or U9385 (N_9385,N_3966,N_1583);
xor U9386 (N_9386,N_1538,N_1704);
xnor U9387 (N_9387,N_1478,N_4831);
nand U9388 (N_9388,N_729,N_2958);
nor U9389 (N_9389,N_1286,N_2343);
nor U9390 (N_9390,N_1970,N_1117);
nand U9391 (N_9391,N_4035,N_3620);
and U9392 (N_9392,N_2686,N_2110);
or U9393 (N_9393,N_52,N_4806);
or U9394 (N_9394,N_4306,N_205);
or U9395 (N_9395,N_3224,N_4863);
or U9396 (N_9396,N_4488,N_4767);
and U9397 (N_9397,N_3586,N_2690);
or U9398 (N_9398,N_438,N_727);
nor U9399 (N_9399,N_3940,N_3581);
nand U9400 (N_9400,N_4721,N_3144);
nand U9401 (N_9401,N_3925,N_3551);
or U9402 (N_9402,N_3555,N_1573);
nor U9403 (N_9403,N_591,N_257);
or U9404 (N_9404,N_574,N_4875);
and U9405 (N_9405,N_2903,N_98);
nor U9406 (N_9406,N_178,N_3794);
nand U9407 (N_9407,N_4224,N_4946);
or U9408 (N_9408,N_2613,N_4842);
xor U9409 (N_9409,N_2509,N_1221);
xnor U9410 (N_9410,N_105,N_2807);
nand U9411 (N_9411,N_3573,N_4869);
and U9412 (N_9412,N_1631,N_3329);
or U9413 (N_9413,N_4340,N_292);
or U9414 (N_9414,N_678,N_79);
or U9415 (N_9415,N_301,N_1109);
and U9416 (N_9416,N_4921,N_3793);
xnor U9417 (N_9417,N_3286,N_4953);
nor U9418 (N_9418,N_351,N_4414);
nor U9419 (N_9419,N_907,N_3489);
or U9420 (N_9420,N_2699,N_983);
and U9421 (N_9421,N_2825,N_3115);
nor U9422 (N_9422,N_3003,N_141);
nor U9423 (N_9423,N_4691,N_1164);
nor U9424 (N_9424,N_4741,N_598);
nand U9425 (N_9425,N_4494,N_1570);
nand U9426 (N_9426,N_2412,N_1523);
nand U9427 (N_9427,N_4966,N_4774);
nor U9428 (N_9428,N_2623,N_4426);
and U9429 (N_9429,N_1522,N_45);
nor U9430 (N_9430,N_4457,N_3951);
nor U9431 (N_9431,N_2085,N_259);
nor U9432 (N_9432,N_1636,N_4146);
nand U9433 (N_9433,N_3940,N_3708);
and U9434 (N_9434,N_1761,N_4399);
and U9435 (N_9435,N_4556,N_4360);
nand U9436 (N_9436,N_3212,N_4167);
or U9437 (N_9437,N_4105,N_1677);
nor U9438 (N_9438,N_3939,N_1503);
and U9439 (N_9439,N_3252,N_4238);
xnor U9440 (N_9440,N_3736,N_529);
and U9441 (N_9441,N_911,N_3321);
xnor U9442 (N_9442,N_2682,N_902);
nand U9443 (N_9443,N_1752,N_8);
or U9444 (N_9444,N_232,N_1948);
nor U9445 (N_9445,N_1890,N_1514);
or U9446 (N_9446,N_3449,N_4835);
nand U9447 (N_9447,N_36,N_3048);
or U9448 (N_9448,N_4488,N_287);
xnor U9449 (N_9449,N_2453,N_2722);
xor U9450 (N_9450,N_4058,N_4804);
nor U9451 (N_9451,N_1395,N_1785);
and U9452 (N_9452,N_1632,N_2704);
or U9453 (N_9453,N_4575,N_3746);
and U9454 (N_9454,N_4041,N_4717);
and U9455 (N_9455,N_3319,N_4438);
xnor U9456 (N_9456,N_4088,N_2900);
xor U9457 (N_9457,N_3784,N_4784);
xnor U9458 (N_9458,N_4966,N_2260);
nand U9459 (N_9459,N_2458,N_2643);
and U9460 (N_9460,N_3720,N_629);
xnor U9461 (N_9461,N_1037,N_3112);
nor U9462 (N_9462,N_3232,N_4083);
or U9463 (N_9463,N_2477,N_4188);
xor U9464 (N_9464,N_1470,N_1756);
nand U9465 (N_9465,N_248,N_802);
nand U9466 (N_9466,N_1554,N_4110);
nor U9467 (N_9467,N_4199,N_1473);
nand U9468 (N_9468,N_2172,N_460);
nand U9469 (N_9469,N_482,N_3652);
nor U9470 (N_9470,N_1041,N_3225);
or U9471 (N_9471,N_3889,N_3587);
xnor U9472 (N_9472,N_2858,N_3685);
or U9473 (N_9473,N_1274,N_3446);
and U9474 (N_9474,N_3229,N_2370);
nor U9475 (N_9475,N_544,N_2430);
xor U9476 (N_9476,N_3234,N_3724);
and U9477 (N_9477,N_4296,N_1641);
nor U9478 (N_9478,N_753,N_1412);
and U9479 (N_9479,N_561,N_1665);
and U9480 (N_9480,N_4328,N_4563);
nor U9481 (N_9481,N_1492,N_3296);
nor U9482 (N_9482,N_1488,N_211);
and U9483 (N_9483,N_2872,N_95);
nor U9484 (N_9484,N_4666,N_4929);
nor U9485 (N_9485,N_126,N_1788);
or U9486 (N_9486,N_3909,N_2469);
or U9487 (N_9487,N_2428,N_3560);
nand U9488 (N_9488,N_4788,N_4564);
and U9489 (N_9489,N_3393,N_2963);
nand U9490 (N_9490,N_3259,N_4683);
nor U9491 (N_9491,N_1154,N_3411);
and U9492 (N_9492,N_2582,N_3305);
nand U9493 (N_9493,N_2226,N_1905);
or U9494 (N_9494,N_4129,N_4957);
and U9495 (N_9495,N_1173,N_4106);
nor U9496 (N_9496,N_2045,N_3835);
nor U9497 (N_9497,N_581,N_1445);
nand U9498 (N_9498,N_1296,N_937);
xnor U9499 (N_9499,N_3340,N_1445);
nand U9500 (N_9500,N_370,N_3531);
xor U9501 (N_9501,N_3778,N_2904);
nor U9502 (N_9502,N_4879,N_320);
nand U9503 (N_9503,N_2156,N_2748);
or U9504 (N_9504,N_4156,N_3494);
nand U9505 (N_9505,N_2612,N_3945);
xor U9506 (N_9506,N_1933,N_4205);
or U9507 (N_9507,N_2064,N_2406);
xor U9508 (N_9508,N_2016,N_2174);
nor U9509 (N_9509,N_3285,N_895);
nor U9510 (N_9510,N_4350,N_1016);
or U9511 (N_9511,N_137,N_1999);
and U9512 (N_9512,N_3165,N_1614);
or U9513 (N_9513,N_1574,N_710);
and U9514 (N_9514,N_1234,N_1487);
and U9515 (N_9515,N_3720,N_2925);
and U9516 (N_9516,N_1454,N_4323);
and U9517 (N_9517,N_1124,N_4469);
xor U9518 (N_9518,N_1746,N_3931);
and U9519 (N_9519,N_3291,N_2491);
nand U9520 (N_9520,N_1875,N_3947);
nor U9521 (N_9521,N_2644,N_3018);
or U9522 (N_9522,N_3079,N_3779);
xnor U9523 (N_9523,N_3258,N_1949);
xor U9524 (N_9524,N_4773,N_2557);
and U9525 (N_9525,N_4042,N_449);
xor U9526 (N_9526,N_2032,N_946);
nand U9527 (N_9527,N_177,N_3742);
xnor U9528 (N_9528,N_1403,N_3383);
nor U9529 (N_9529,N_2548,N_1029);
or U9530 (N_9530,N_4525,N_4130);
nand U9531 (N_9531,N_2718,N_3854);
and U9532 (N_9532,N_523,N_1924);
nand U9533 (N_9533,N_1001,N_4193);
nand U9534 (N_9534,N_1395,N_4346);
nor U9535 (N_9535,N_4649,N_4908);
nand U9536 (N_9536,N_1176,N_2027);
or U9537 (N_9537,N_2871,N_3584);
or U9538 (N_9538,N_4089,N_3722);
nor U9539 (N_9539,N_1477,N_1141);
nand U9540 (N_9540,N_2118,N_285);
or U9541 (N_9541,N_839,N_4927);
nor U9542 (N_9542,N_116,N_2809);
nand U9543 (N_9543,N_2736,N_4267);
xor U9544 (N_9544,N_1890,N_2795);
xor U9545 (N_9545,N_3548,N_3687);
and U9546 (N_9546,N_434,N_4999);
nor U9547 (N_9547,N_3771,N_169);
or U9548 (N_9548,N_1379,N_2632);
nand U9549 (N_9549,N_74,N_846);
xor U9550 (N_9550,N_1690,N_4965);
and U9551 (N_9551,N_3514,N_2419);
or U9552 (N_9552,N_691,N_4810);
or U9553 (N_9553,N_4560,N_2459);
xor U9554 (N_9554,N_1805,N_2068);
or U9555 (N_9555,N_1718,N_4466);
and U9556 (N_9556,N_261,N_398);
and U9557 (N_9557,N_2989,N_316);
nor U9558 (N_9558,N_2152,N_4660);
nand U9559 (N_9559,N_2505,N_368);
and U9560 (N_9560,N_2208,N_991);
and U9561 (N_9561,N_3299,N_4518);
nor U9562 (N_9562,N_2957,N_3199);
nand U9563 (N_9563,N_3881,N_551);
nor U9564 (N_9564,N_3725,N_3205);
xor U9565 (N_9565,N_3159,N_2718);
xnor U9566 (N_9566,N_4909,N_481);
nor U9567 (N_9567,N_1736,N_3131);
nand U9568 (N_9568,N_538,N_3800);
nand U9569 (N_9569,N_468,N_4157);
xnor U9570 (N_9570,N_3587,N_3030);
xor U9571 (N_9571,N_1666,N_3561);
and U9572 (N_9572,N_2589,N_4243);
or U9573 (N_9573,N_4113,N_4522);
nand U9574 (N_9574,N_218,N_4548);
and U9575 (N_9575,N_3794,N_1577);
or U9576 (N_9576,N_341,N_3564);
xor U9577 (N_9577,N_2089,N_1230);
or U9578 (N_9578,N_923,N_1847);
nand U9579 (N_9579,N_4684,N_2201);
nand U9580 (N_9580,N_1483,N_63);
nand U9581 (N_9581,N_3172,N_4166);
nand U9582 (N_9582,N_4747,N_4892);
xor U9583 (N_9583,N_1453,N_4371);
nor U9584 (N_9584,N_2896,N_1575);
xor U9585 (N_9585,N_3024,N_4839);
nor U9586 (N_9586,N_1602,N_3352);
nor U9587 (N_9587,N_2385,N_3191);
nand U9588 (N_9588,N_3807,N_62);
or U9589 (N_9589,N_1352,N_1616);
or U9590 (N_9590,N_217,N_2219);
xor U9591 (N_9591,N_4357,N_3894);
xor U9592 (N_9592,N_4263,N_1809);
and U9593 (N_9593,N_1299,N_1555);
nand U9594 (N_9594,N_4574,N_408);
xnor U9595 (N_9595,N_1259,N_3912);
nor U9596 (N_9596,N_1082,N_1371);
or U9597 (N_9597,N_862,N_3695);
nor U9598 (N_9598,N_66,N_3083);
and U9599 (N_9599,N_685,N_1259);
nand U9600 (N_9600,N_3046,N_4316);
nand U9601 (N_9601,N_754,N_3765);
xor U9602 (N_9602,N_4668,N_4934);
xor U9603 (N_9603,N_4171,N_1687);
nor U9604 (N_9604,N_4356,N_4775);
and U9605 (N_9605,N_4517,N_3541);
nor U9606 (N_9606,N_3980,N_3939);
nand U9607 (N_9607,N_3000,N_3475);
nor U9608 (N_9608,N_4341,N_2917);
nor U9609 (N_9609,N_3443,N_491);
and U9610 (N_9610,N_1725,N_737);
xnor U9611 (N_9611,N_1312,N_4268);
nand U9612 (N_9612,N_4762,N_1600);
nand U9613 (N_9613,N_1987,N_104);
nand U9614 (N_9614,N_4668,N_1751);
xor U9615 (N_9615,N_4019,N_3233);
or U9616 (N_9616,N_4982,N_257);
nor U9617 (N_9617,N_3260,N_2722);
nor U9618 (N_9618,N_1071,N_3859);
nand U9619 (N_9619,N_1774,N_454);
and U9620 (N_9620,N_2378,N_1629);
and U9621 (N_9621,N_1211,N_4344);
or U9622 (N_9622,N_2188,N_2354);
and U9623 (N_9623,N_3583,N_1337);
and U9624 (N_9624,N_3772,N_3638);
or U9625 (N_9625,N_1884,N_961);
nand U9626 (N_9626,N_1724,N_1757);
nor U9627 (N_9627,N_2135,N_3128);
nand U9628 (N_9628,N_829,N_571);
and U9629 (N_9629,N_2357,N_935);
nand U9630 (N_9630,N_1070,N_4156);
or U9631 (N_9631,N_3520,N_4482);
or U9632 (N_9632,N_4211,N_4206);
nand U9633 (N_9633,N_4976,N_3739);
and U9634 (N_9634,N_25,N_1239);
nor U9635 (N_9635,N_3116,N_2444);
and U9636 (N_9636,N_495,N_3279);
and U9637 (N_9637,N_2400,N_3370);
and U9638 (N_9638,N_4461,N_3575);
nand U9639 (N_9639,N_4830,N_1108);
xnor U9640 (N_9640,N_1933,N_3562);
or U9641 (N_9641,N_63,N_138);
and U9642 (N_9642,N_892,N_4511);
and U9643 (N_9643,N_2565,N_3472);
xnor U9644 (N_9644,N_2872,N_2327);
nand U9645 (N_9645,N_1950,N_2075);
or U9646 (N_9646,N_4075,N_448);
nand U9647 (N_9647,N_2791,N_4601);
xor U9648 (N_9648,N_3622,N_976);
xnor U9649 (N_9649,N_4630,N_3296);
or U9650 (N_9650,N_1157,N_1646);
xnor U9651 (N_9651,N_78,N_2104);
nand U9652 (N_9652,N_3305,N_4958);
nand U9653 (N_9653,N_2751,N_2261);
nor U9654 (N_9654,N_448,N_4440);
or U9655 (N_9655,N_1937,N_239);
or U9656 (N_9656,N_1813,N_2767);
and U9657 (N_9657,N_2961,N_3172);
and U9658 (N_9658,N_2265,N_3021);
and U9659 (N_9659,N_159,N_1586);
or U9660 (N_9660,N_726,N_2944);
xor U9661 (N_9661,N_3160,N_4667);
xnor U9662 (N_9662,N_1719,N_4374);
nand U9663 (N_9663,N_2164,N_4856);
nor U9664 (N_9664,N_2778,N_1889);
xor U9665 (N_9665,N_364,N_3174);
xnor U9666 (N_9666,N_4530,N_3261);
and U9667 (N_9667,N_131,N_4010);
xor U9668 (N_9668,N_3873,N_4556);
or U9669 (N_9669,N_2599,N_2237);
or U9670 (N_9670,N_418,N_948);
and U9671 (N_9671,N_3883,N_1771);
and U9672 (N_9672,N_1815,N_3125);
and U9673 (N_9673,N_4708,N_3047);
and U9674 (N_9674,N_3010,N_1628);
nor U9675 (N_9675,N_1806,N_1880);
nand U9676 (N_9676,N_2505,N_4019);
or U9677 (N_9677,N_1325,N_2662);
xnor U9678 (N_9678,N_1354,N_4213);
nand U9679 (N_9679,N_72,N_81);
nand U9680 (N_9680,N_3935,N_1500);
xor U9681 (N_9681,N_4479,N_1523);
or U9682 (N_9682,N_2906,N_530);
and U9683 (N_9683,N_1811,N_1852);
and U9684 (N_9684,N_4878,N_334);
nand U9685 (N_9685,N_3757,N_1335);
and U9686 (N_9686,N_4279,N_1125);
xnor U9687 (N_9687,N_4750,N_1505);
nor U9688 (N_9688,N_2022,N_2449);
or U9689 (N_9689,N_4051,N_3568);
nor U9690 (N_9690,N_933,N_3784);
xor U9691 (N_9691,N_2475,N_2342);
nand U9692 (N_9692,N_2094,N_2632);
or U9693 (N_9693,N_1747,N_2800);
nand U9694 (N_9694,N_2797,N_348);
nand U9695 (N_9695,N_2239,N_1951);
xnor U9696 (N_9696,N_3511,N_1607);
nor U9697 (N_9697,N_3199,N_3813);
nor U9698 (N_9698,N_4122,N_219);
nand U9699 (N_9699,N_944,N_1843);
and U9700 (N_9700,N_4239,N_1127);
or U9701 (N_9701,N_4852,N_1964);
or U9702 (N_9702,N_3174,N_4189);
and U9703 (N_9703,N_1532,N_1802);
and U9704 (N_9704,N_2323,N_366);
nor U9705 (N_9705,N_716,N_4154);
nand U9706 (N_9706,N_3518,N_551);
and U9707 (N_9707,N_1462,N_196);
nand U9708 (N_9708,N_1488,N_3183);
nand U9709 (N_9709,N_1807,N_1255);
and U9710 (N_9710,N_1023,N_4167);
xor U9711 (N_9711,N_2826,N_2336);
and U9712 (N_9712,N_2348,N_4009);
or U9713 (N_9713,N_2749,N_4929);
or U9714 (N_9714,N_4024,N_3679);
or U9715 (N_9715,N_1487,N_1956);
or U9716 (N_9716,N_2819,N_2767);
and U9717 (N_9717,N_4965,N_4145);
nand U9718 (N_9718,N_520,N_2162);
nor U9719 (N_9719,N_3523,N_432);
and U9720 (N_9720,N_978,N_2333);
nand U9721 (N_9721,N_1237,N_1058);
and U9722 (N_9722,N_4375,N_520);
and U9723 (N_9723,N_2997,N_650);
or U9724 (N_9724,N_1308,N_2638);
xor U9725 (N_9725,N_188,N_1655);
and U9726 (N_9726,N_3384,N_2782);
xnor U9727 (N_9727,N_3402,N_1091);
nor U9728 (N_9728,N_2991,N_2689);
xor U9729 (N_9729,N_1583,N_3187);
or U9730 (N_9730,N_931,N_1853);
or U9731 (N_9731,N_2637,N_4976);
or U9732 (N_9732,N_2195,N_1976);
nand U9733 (N_9733,N_1424,N_2509);
and U9734 (N_9734,N_921,N_3124);
or U9735 (N_9735,N_1678,N_3100);
and U9736 (N_9736,N_2354,N_1926);
nor U9737 (N_9737,N_1285,N_3960);
or U9738 (N_9738,N_4277,N_3001);
nor U9739 (N_9739,N_4446,N_4852);
or U9740 (N_9740,N_838,N_3509);
nor U9741 (N_9741,N_4712,N_1180);
xor U9742 (N_9742,N_3046,N_4565);
nand U9743 (N_9743,N_876,N_3035);
or U9744 (N_9744,N_1572,N_3224);
or U9745 (N_9745,N_4174,N_3800);
xor U9746 (N_9746,N_4889,N_4623);
and U9747 (N_9747,N_2338,N_4573);
or U9748 (N_9748,N_2310,N_3360);
and U9749 (N_9749,N_1821,N_583);
and U9750 (N_9750,N_4863,N_4419);
nor U9751 (N_9751,N_1399,N_174);
and U9752 (N_9752,N_1086,N_875);
nor U9753 (N_9753,N_2792,N_2362);
and U9754 (N_9754,N_1152,N_2453);
nor U9755 (N_9755,N_2951,N_2919);
and U9756 (N_9756,N_4598,N_3681);
nand U9757 (N_9757,N_406,N_1140);
and U9758 (N_9758,N_4011,N_3040);
nor U9759 (N_9759,N_799,N_889);
nand U9760 (N_9760,N_1989,N_1587);
and U9761 (N_9761,N_1318,N_2275);
and U9762 (N_9762,N_1609,N_3036);
or U9763 (N_9763,N_412,N_1395);
nand U9764 (N_9764,N_4497,N_3154);
and U9765 (N_9765,N_480,N_2300);
and U9766 (N_9766,N_780,N_3379);
nor U9767 (N_9767,N_2686,N_69);
or U9768 (N_9768,N_4245,N_4474);
and U9769 (N_9769,N_3169,N_4660);
nand U9770 (N_9770,N_3557,N_3401);
nor U9771 (N_9771,N_2021,N_931);
or U9772 (N_9772,N_4520,N_1952);
nor U9773 (N_9773,N_4779,N_2168);
and U9774 (N_9774,N_3403,N_2112);
and U9775 (N_9775,N_4155,N_2839);
nand U9776 (N_9776,N_1851,N_4262);
nor U9777 (N_9777,N_3119,N_852);
nand U9778 (N_9778,N_1618,N_25);
or U9779 (N_9779,N_723,N_1791);
or U9780 (N_9780,N_2387,N_3172);
or U9781 (N_9781,N_4144,N_3764);
or U9782 (N_9782,N_1112,N_4915);
and U9783 (N_9783,N_4338,N_4298);
xnor U9784 (N_9784,N_3492,N_1552);
and U9785 (N_9785,N_3178,N_2194);
xnor U9786 (N_9786,N_2745,N_3344);
nor U9787 (N_9787,N_2665,N_1495);
or U9788 (N_9788,N_1313,N_1186);
nor U9789 (N_9789,N_3359,N_3606);
and U9790 (N_9790,N_3273,N_4378);
or U9791 (N_9791,N_2764,N_3687);
nor U9792 (N_9792,N_2399,N_4248);
or U9793 (N_9793,N_126,N_2944);
nand U9794 (N_9794,N_2124,N_3206);
nand U9795 (N_9795,N_1727,N_661);
or U9796 (N_9796,N_2450,N_2036);
and U9797 (N_9797,N_2842,N_4442);
and U9798 (N_9798,N_237,N_1754);
or U9799 (N_9799,N_246,N_1237);
xnor U9800 (N_9800,N_1854,N_3220);
nand U9801 (N_9801,N_1486,N_1904);
nand U9802 (N_9802,N_902,N_1999);
nand U9803 (N_9803,N_3905,N_3268);
nor U9804 (N_9804,N_2989,N_2126);
nor U9805 (N_9805,N_2568,N_733);
and U9806 (N_9806,N_1792,N_300);
nor U9807 (N_9807,N_1174,N_1297);
or U9808 (N_9808,N_40,N_2437);
xor U9809 (N_9809,N_907,N_1723);
nand U9810 (N_9810,N_2475,N_3505);
xnor U9811 (N_9811,N_3605,N_150);
nor U9812 (N_9812,N_1521,N_3565);
xor U9813 (N_9813,N_3087,N_2830);
xor U9814 (N_9814,N_4303,N_3114);
nor U9815 (N_9815,N_445,N_3734);
nor U9816 (N_9816,N_4068,N_1019);
nand U9817 (N_9817,N_2020,N_1648);
and U9818 (N_9818,N_115,N_4147);
and U9819 (N_9819,N_3707,N_3093);
xor U9820 (N_9820,N_3882,N_169);
xor U9821 (N_9821,N_4428,N_4682);
nor U9822 (N_9822,N_2151,N_2218);
nor U9823 (N_9823,N_4188,N_3049);
xnor U9824 (N_9824,N_2044,N_4135);
or U9825 (N_9825,N_1643,N_1760);
or U9826 (N_9826,N_2046,N_4335);
nand U9827 (N_9827,N_3168,N_4689);
xor U9828 (N_9828,N_3149,N_204);
or U9829 (N_9829,N_2881,N_1385);
nor U9830 (N_9830,N_1067,N_3642);
or U9831 (N_9831,N_3564,N_3186);
nor U9832 (N_9832,N_4543,N_4874);
or U9833 (N_9833,N_1192,N_2180);
xnor U9834 (N_9834,N_4479,N_467);
or U9835 (N_9835,N_2234,N_3691);
or U9836 (N_9836,N_370,N_2162);
nand U9837 (N_9837,N_1915,N_1456);
and U9838 (N_9838,N_2327,N_2991);
and U9839 (N_9839,N_4772,N_4990);
nand U9840 (N_9840,N_1121,N_2305);
and U9841 (N_9841,N_4097,N_2106);
nand U9842 (N_9842,N_3848,N_87);
and U9843 (N_9843,N_118,N_2214);
and U9844 (N_9844,N_3477,N_2662);
or U9845 (N_9845,N_4730,N_4266);
nor U9846 (N_9846,N_2871,N_763);
nor U9847 (N_9847,N_2077,N_1874);
nor U9848 (N_9848,N_458,N_2245);
xnor U9849 (N_9849,N_292,N_2807);
or U9850 (N_9850,N_4346,N_4866);
nand U9851 (N_9851,N_4904,N_4906);
nor U9852 (N_9852,N_3692,N_4233);
nor U9853 (N_9853,N_563,N_3758);
or U9854 (N_9854,N_4532,N_3587);
nor U9855 (N_9855,N_2830,N_2144);
and U9856 (N_9856,N_42,N_3641);
or U9857 (N_9857,N_4483,N_3436);
nor U9858 (N_9858,N_4935,N_4458);
nand U9859 (N_9859,N_3583,N_3171);
and U9860 (N_9860,N_1239,N_2384);
or U9861 (N_9861,N_78,N_4243);
and U9862 (N_9862,N_1654,N_4532);
xor U9863 (N_9863,N_4059,N_1905);
nand U9864 (N_9864,N_2149,N_2587);
nor U9865 (N_9865,N_856,N_3860);
nand U9866 (N_9866,N_1092,N_1159);
nand U9867 (N_9867,N_4051,N_4440);
or U9868 (N_9868,N_4133,N_781);
nand U9869 (N_9869,N_739,N_3796);
nand U9870 (N_9870,N_3276,N_3981);
or U9871 (N_9871,N_2265,N_400);
nand U9872 (N_9872,N_2436,N_610);
nand U9873 (N_9873,N_843,N_3151);
or U9874 (N_9874,N_741,N_3470);
nor U9875 (N_9875,N_3749,N_4266);
nor U9876 (N_9876,N_1969,N_1614);
or U9877 (N_9877,N_2452,N_1434);
xor U9878 (N_9878,N_3948,N_522);
nor U9879 (N_9879,N_4920,N_155);
xor U9880 (N_9880,N_4191,N_411);
nor U9881 (N_9881,N_1461,N_4832);
or U9882 (N_9882,N_2810,N_4631);
and U9883 (N_9883,N_590,N_2740);
nand U9884 (N_9884,N_555,N_1481);
xor U9885 (N_9885,N_1530,N_828);
or U9886 (N_9886,N_4417,N_1216);
xnor U9887 (N_9887,N_1324,N_4663);
nand U9888 (N_9888,N_4281,N_1354);
or U9889 (N_9889,N_1666,N_2424);
and U9890 (N_9890,N_3472,N_840);
xnor U9891 (N_9891,N_703,N_3921);
or U9892 (N_9892,N_805,N_825);
nand U9893 (N_9893,N_3615,N_161);
xor U9894 (N_9894,N_4467,N_4733);
nor U9895 (N_9895,N_356,N_3812);
and U9896 (N_9896,N_4283,N_232);
or U9897 (N_9897,N_3082,N_2847);
xor U9898 (N_9898,N_1463,N_1555);
or U9899 (N_9899,N_725,N_4623);
nor U9900 (N_9900,N_2364,N_3260);
nand U9901 (N_9901,N_652,N_4220);
and U9902 (N_9902,N_1223,N_3542);
and U9903 (N_9903,N_3719,N_1347);
or U9904 (N_9904,N_4339,N_4816);
xnor U9905 (N_9905,N_2381,N_4068);
or U9906 (N_9906,N_1830,N_4387);
and U9907 (N_9907,N_1662,N_610);
nand U9908 (N_9908,N_4562,N_243);
and U9909 (N_9909,N_2493,N_1596);
nand U9910 (N_9910,N_4183,N_281);
or U9911 (N_9911,N_1894,N_1461);
nand U9912 (N_9912,N_3247,N_2334);
and U9913 (N_9913,N_298,N_218);
nor U9914 (N_9914,N_735,N_4414);
or U9915 (N_9915,N_2045,N_415);
nand U9916 (N_9916,N_3949,N_895);
xor U9917 (N_9917,N_1319,N_1073);
and U9918 (N_9918,N_3347,N_2719);
nand U9919 (N_9919,N_3994,N_4519);
nand U9920 (N_9920,N_194,N_759);
and U9921 (N_9921,N_3706,N_3935);
and U9922 (N_9922,N_464,N_2939);
and U9923 (N_9923,N_1487,N_3766);
or U9924 (N_9924,N_3945,N_2706);
nand U9925 (N_9925,N_608,N_2477);
or U9926 (N_9926,N_1327,N_2023);
or U9927 (N_9927,N_2188,N_3802);
and U9928 (N_9928,N_1769,N_4935);
nor U9929 (N_9929,N_580,N_2814);
and U9930 (N_9930,N_3257,N_4612);
or U9931 (N_9931,N_190,N_4005);
and U9932 (N_9932,N_3938,N_4484);
and U9933 (N_9933,N_1723,N_4670);
xnor U9934 (N_9934,N_4887,N_1657);
nor U9935 (N_9935,N_3356,N_2455);
xor U9936 (N_9936,N_4684,N_2332);
or U9937 (N_9937,N_2385,N_3180);
xor U9938 (N_9938,N_568,N_3193);
nor U9939 (N_9939,N_4742,N_428);
and U9940 (N_9940,N_3122,N_958);
xnor U9941 (N_9941,N_1522,N_1319);
and U9942 (N_9942,N_3227,N_2617);
nor U9943 (N_9943,N_1976,N_1167);
nor U9944 (N_9944,N_581,N_1962);
nor U9945 (N_9945,N_2717,N_2023);
and U9946 (N_9946,N_2613,N_4944);
or U9947 (N_9947,N_4362,N_2363);
or U9948 (N_9948,N_700,N_1629);
or U9949 (N_9949,N_375,N_1135);
and U9950 (N_9950,N_830,N_4035);
or U9951 (N_9951,N_1609,N_3655);
nor U9952 (N_9952,N_542,N_3887);
nor U9953 (N_9953,N_1644,N_3544);
nand U9954 (N_9954,N_4843,N_2436);
and U9955 (N_9955,N_3917,N_948);
or U9956 (N_9956,N_973,N_1259);
or U9957 (N_9957,N_1049,N_174);
and U9958 (N_9958,N_3874,N_1979);
nor U9959 (N_9959,N_4562,N_1128);
nand U9960 (N_9960,N_3628,N_3958);
or U9961 (N_9961,N_2526,N_2736);
nand U9962 (N_9962,N_433,N_3719);
xnor U9963 (N_9963,N_4655,N_2941);
and U9964 (N_9964,N_1258,N_2822);
nor U9965 (N_9965,N_2804,N_4811);
or U9966 (N_9966,N_4069,N_4490);
nand U9967 (N_9967,N_4028,N_1945);
nor U9968 (N_9968,N_3917,N_1823);
xnor U9969 (N_9969,N_4535,N_4473);
nor U9970 (N_9970,N_4374,N_1913);
xor U9971 (N_9971,N_2491,N_1725);
xor U9972 (N_9972,N_4006,N_4290);
or U9973 (N_9973,N_3114,N_923);
or U9974 (N_9974,N_4285,N_3195);
nand U9975 (N_9975,N_4188,N_3062);
or U9976 (N_9976,N_3935,N_3162);
or U9977 (N_9977,N_2017,N_2561);
or U9978 (N_9978,N_4374,N_4767);
nor U9979 (N_9979,N_4314,N_2920);
xnor U9980 (N_9980,N_1787,N_4894);
nor U9981 (N_9981,N_4710,N_4395);
xor U9982 (N_9982,N_4456,N_2542);
and U9983 (N_9983,N_4978,N_3189);
and U9984 (N_9984,N_2895,N_4325);
and U9985 (N_9985,N_1730,N_3002);
xnor U9986 (N_9986,N_2389,N_2127);
xor U9987 (N_9987,N_3272,N_1272);
or U9988 (N_9988,N_3094,N_4149);
or U9989 (N_9989,N_1837,N_473);
nor U9990 (N_9990,N_559,N_2291);
xor U9991 (N_9991,N_3070,N_1464);
xor U9992 (N_9992,N_572,N_2855);
or U9993 (N_9993,N_2695,N_2255);
or U9994 (N_9994,N_614,N_3228);
nand U9995 (N_9995,N_3993,N_993);
xnor U9996 (N_9996,N_1500,N_4604);
and U9997 (N_9997,N_1614,N_3942);
nand U9998 (N_9998,N_2794,N_2132);
and U9999 (N_9999,N_3293,N_296);
and U10000 (N_10000,N_6225,N_5000);
nor U10001 (N_10001,N_7527,N_6246);
nand U10002 (N_10002,N_5499,N_7016);
or U10003 (N_10003,N_7511,N_9396);
xor U10004 (N_10004,N_7610,N_5542);
nand U10005 (N_10005,N_7187,N_9167);
nand U10006 (N_10006,N_9412,N_5174);
or U10007 (N_10007,N_8291,N_6650);
and U10008 (N_10008,N_7532,N_9054);
nand U10009 (N_10009,N_7025,N_6054);
or U10010 (N_10010,N_9707,N_9518);
xor U10011 (N_10011,N_6792,N_8537);
nand U10012 (N_10012,N_8315,N_9478);
xnor U10013 (N_10013,N_5705,N_9304);
nand U10014 (N_10014,N_7769,N_5994);
nand U10015 (N_10015,N_6907,N_8087);
nor U10016 (N_10016,N_6090,N_5795);
nand U10017 (N_10017,N_6699,N_9076);
xor U10018 (N_10018,N_7036,N_6071);
nor U10019 (N_10019,N_8363,N_9634);
or U10020 (N_10020,N_6053,N_8621);
nor U10021 (N_10021,N_9460,N_6689);
xnor U10022 (N_10022,N_8675,N_7596);
or U10023 (N_10023,N_7560,N_9057);
nand U10024 (N_10024,N_9116,N_9899);
nand U10025 (N_10025,N_6942,N_6450);
or U10026 (N_10026,N_5647,N_8521);
nand U10027 (N_10027,N_8000,N_7108);
nor U10028 (N_10028,N_8443,N_8078);
and U10029 (N_10029,N_7185,N_5677);
nor U10030 (N_10030,N_9719,N_9286);
xor U10031 (N_10031,N_7049,N_8891);
and U10032 (N_10032,N_8049,N_5361);
xnor U10033 (N_10033,N_6295,N_9986);
nor U10034 (N_10034,N_5833,N_6874);
nor U10035 (N_10035,N_5044,N_8316);
and U10036 (N_10036,N_6336,N_9061);
nor U10037 (N_10037,N_9356,N_6515);
nor U10038 (N_10038,N_5513,N_6543);
nor U10039 (N_10039,N_7396,N_9758);
xor U10040 (N_10040,N_7044,N_7363);
or U10041 (N_10041,N_8089,N_6341);
xnor U10042 (N_10042,N_7866,N_9547);
nand U10043 (N_10043,N_9425,N_5024);
and U10044 (N_10044,N_9801,N_9436);
and U10045 (N_10045,N_9000,N_6372);
nand U10046 (N_10046,N_7197,N_7010);
nand U10047 (N_10047,N_8310,N_5548);
and U10048 (N_10048,N_6769,N_6241);
xnor U10049 (N_10049,N_5657,N_6023);
nand U10050 (N_10050,N_9843,N_6891);
and U10051 (N_10051,N_7570,N_8102);
nor U10052 (N_10052,N_7736,N_8012);
nand U10053 (N_10053,N_9643,N_9528);
nor U10054 (N_10054,N_5124,N_6832);
nor U10055 (N_10055,N_6464,N_9946);
nand U10056 (N_10056,N_6229,N_5557);
and U10057 (N_10057,N_9674,N_5093);
or U10058 (N_10058,N_6919,N_7141);
xor U10059 (N_10059,N_6320,N_8014);
and U10060 (N_10060,N_6974,N_8511);
nand U10061 (N_10061,N_7754,N_5637);
xor U10062 (N_10062,N_6644,N_9560);
or U10063 (N_10063,N_8506,N_8736);
or U10064 (N_10064,N_7882,N_6763);
or U10065 (N_10065,N_8331,N_9533);
or U10066 (N_10066,N_8913,N_6161);
or U10067 (N_10067,N_5570,N_6804);
nand U10068 (N_10068,N_8903,N_8971);
and U10069 (N_10069,N_7526,N_8759);
nand U10070 (N_10070,N_8898,N_7340);
nor U10071 (N_10071,N_8026,N_5720);
nand U10072 (N_10072,N_6685,N_6022);
or U10073 (N_10073,N_9979,N_9174);
and U10074 (N_10074,N_8941,N_5263);
or U10075 (N_10075,N_9339,N_6383);
nand U10076 (N_10076,N_5250,N_6684);
and U10077 (N_10077,N_7784,N_6790);
and U10078 (N_10078,N_8622,N_8356);
nor U10079 (N_10079,N_8646,N_6553);
or U10080 (N_10080,N_5514,N_8803);
nor U10081 (N_10081,N_5804,N_8233);
nand U10082 (N_10082,N_7216,N_9866);
nor U10083 (N_10083,N_5006,N_9820);
and U10084 (N_10084,N_5281,N_5616);
nor U10085 (N_10085,N_5672,N_7382);
nor U10086 (N_10086,N_8387,N_7004);
nand U10087 (N_10087,N_7297,N_5107);
nor U10088 (N_10088,N_5929,N_6042);
nand U10089 (N_10089,N_5908,N_8836);
nor U10090 (N_10090,N_7895,N_9583);
xnor U10091 (N_10091,N_6806,N_6932);
or U10092 (N_10092,N_9814,N_6351);
or U10093 (N_10093,N_5734,N_7224);
xnor U10094 (N_10094,N_5111,N_9012);
xor U10095 (N_10095,N_7559,N_7376);
xnor U10096 (N_10096,N_7426,N_8340);
xor U10097 (N_10097,N_9661,N_7764);
xor U10098 (N_10098,N_9324,N_5416);
nand U10099 (N_10099,N_5079,N_8307);
nand U10100 (N_10100,N_5597,N_6688);
nand U10101 (N_10101,N_5354,N_6875);
nand U10102 (N_10102,N_8961,N_6014);
nor U10103 (N_10103,N_6619,N_9744);
or U10104 (N_10104,N_7674,N_7354);
and U10105 (N_10105,N_8351,N_7473);
nor U10106 (N_10106,N_6902,N_7497);
nor U10107 (N_10107,N_5751,N_6477);
and U10108 (N_10108,N_5138,N_5539);
and U10109 (N_10109,N_9085,N_7208);
or U10110 (N_10110,N_6539,N_9865);
nor U10111 (N_10111,N_8042,N_6368);
or U10112 (N_10112,N_5625,N_7673);
and U10113 (N_10113,N_7359,N_7186);
nand U10114 (N_10114,N_7849,N_5295);
nor U10115 (N_10115,N_9739,N_9751);
nand U10116 (N_10116,N_7465,N_9181);
nor U10117 (N_10117,N_5309,N_9546);
or U10118 (N_10118,N_9123,N_6583);
nor U10119 (N_10119,N_5709,N_5817);
or U10120 (N_10120,N_6597,N_7593);
and U10121 (N_10121,N_7933,N_6995);
nand U10122 (N_10122,N_8477,N_5075);
xor U10123 (N_10123,N_9694,N_5988);
and U10124 (N_10124,N_5066,N_7577);
and U10125 (N_10125,N_5633,N_9168);
and U10126 (N_10126,N_6065,N_8981);
or U10127 (N_10127,N_8261,N_5879);
nand U10128 (N_10128,N_5293,N_8928);
nand U10129 (N_10129,N_9972,N_8203);
xnor U10130 (N_10130,N_9235,N_5171);
or U10131 (N_10131,N_9691,N_8910);
nand U10132 (N_10132,N_8999,N_5134);
nand U10133 (N_10133,N_5407,N_7615);
and U10134 (N_10134,N_9182,N_7647);
or U10135 (N_10135,N_8894,N_7496);
or U10136 (N_10136,N_8714,N_5648);
or U10137 (N_10137,N_6214,N_5193);
and U10138 (N_10138,N_6937,N_9483);
or U10139 (N_10139,N_5360,N_9535);
xor U10140 (N_10140,N_9937,N_7361);
and U10141 (N_10141,N_9156,N_9921);
nor U10142 (N_10142,N_5797,N_5957);
nor U10143 (N_10143,N_9296,N_9203);
nor U10144 (N_10144,N_5646,N_6044);
xor U10145 (N_10145,N_7232,N_9112);
xnor U10146 (N_10146,N_8332,N_7694);
nor U10147 (N_10147,N_6510,N_6513);
and U10148 (N_10148,N_8962,N_5356);
xor U10149 (N_10149,N_6289,N_6439);
and U10150 (N_10150,N_9141,N_7468);
xnor U10151 (N_10151,N_6716,N_9936);
and U10152 (N_10152,N_7196,N_6869);
nand U10153 (N_10153,N_6871,N_8755);
xnor U10154 (N_10154,N_9432,N_6112);
nand U10155 (N_10155,N_7734,N_9733);
or U10156 (N_10156,N_7793,N_8181);
nand U10157 (N_10157,N_5924,N_7977);
nor U10158 (N_10158,N_9851,N_8439);
and U10159 (N_10159,N_5213,N_7225);
or U10160 (N_10160,N_6444,N_7791);
nor U10161 (N_10161,N_6984,N_5338);
nor U10162 (N_10162,N_7198,N_9512);
and U10163 (N_10163,N_9603,N_6549);
or U10164 (N_10164,N_6658,N_5890);
xnor U10165 (N_10165,N_9928,N_7774);
nor U10166 (N_10166,N_5381,N_8769);
or U10167 (N_10167,N_6627,N_9294);
nand U10168 (N_10168,N_9420,N_5023);
or U10169 (N_10169,N_7427,N_6475);
nand U10170 (N_10170,N_5915,N_6774);
xnor U10171 (N_10171,N_7257,N_6133);
nor U10172 (N_10172,N_6537,N_7029);
or U10173 (N_10173,N_9514,N_5313);
and U10174 (N_10174,N_7488,N_7444);
nand U10175 (N_10175,N_5078,N_5554);
xnor U10176 (N_10176,N_6200,N_6777);
nand U10177 (N_10177,N_5184,N_9492);
or U10178 (N_10178,N_7850,N_8508);
and U10179 (N_10179,N_9569,N_8562);
nand U10180 (N_10180,N_7301,N_7242);
or U10181 (N_10181,N_6279,N_7751);
and U10182 (N_10182,N_5605,N_9242);
and U10183 (N_10183,N_7909,N_6409);
or U10184 (N_10184,N_9151,N_7438);
xor U10185 (N_10185,N_7403,N_8818);
xnor U10186 (N_10186,N_8832,N_8745);
and U10187 (N_10187,N_9407,N_9943);
nor U10188 (N_10188,N_9735,N_6296);
and U10189 (N_10189,N_6945,N_9025);
or U10190 (N_10190,N_7926,N_6518);
and U10191 (N_10191,N_8826,N_7355);
xor U10192 (N_10192,N_8733,N_8752);
or U10193 (N_10193,N_9374,N_7262);
xor U10194 (N_10194,N_9708,N_8044);
nor U10195 (N_10195,N_5087,N_7210);
nand U10196 (N_10196,N_7495,N_5277);
and U10197 (N_10197,N_9393,N_6394);
or U10198 (N_10198,N_5673,N_7084);
nor U10199 (N_10199,N_7041,N_9490);
and U10200 (N_10200,N_8636,N_5242);
or U10201 (N_10201,N_8209,N_9976);
or U10202 (N_10202,N_9952,N_9699);
xnor U10203 (N_10203,N_8187,N_5674);
xor U10204 (N_10204,N_5246,N_8976);
nand U10205 (N_10205,N_6753,N_9347);
nor U10206 (N_10206,N_7170,N_5463);
or U10207 (N_10207,N_6025,N_9780);
xor U10208 (N_10208,N_9981,N_6460);
nor U10209 (N_10209,N_8041,N_9348);
nand U10210 (N_10210,N_7020,N_7556);
and U10211 (N_10211,N_9785,N_5712);
nor U10212 (N_10212,N_5930,N_8608);
nor U10213 (N_10213,N_8278,N_9344);
nor U10214 (N_10214,N_5995,N_6916);
xnor U10215 (N_10215,N_8334,N_9874);
nand U10216 (N_10216,N_7443,N_8220);
nor U10217 (N_10217,N_7146,N_8101);
xnor U10218 (N_10218,N_7147,N_7890);
xnor U10219 (N_10219,N_5442,N_6138);
or U10220 (N_10220,N_5469,N_9641);
or U10221 (N_10221,N_7879,N_6507);
nand U10222 (N_10222,N_9137,N_8716);
or U10223 (N_10223,N_7578,N_5651);
or U10224 (N_10224,N_5280,N_9280);
and U10225 (N_10225,N_6135,N_9971);
nand U10226 (N_10226,N_5460,N_6365);
nor U10227 (N_10227,N_5900,N_7489);
or U10228 (N_10228,N_8343,N_7436);
and U10229 (N_10229,N_9748,N_7070);
xnor U10230 (N_10230,N_5653,N_5229);
and U10231 (N_10231,N_6980,N_6099);
and U10232 (N_10232,N_5088,N_7737);
or U10233 (N_10233,N_7843,N_8066);
and U10234 (N_10234,N_8448,N_7523);
and U10235 (N_10235,N_9718,N_6678);
or U10236 (N_10236,N_7291,N_8839);
or U10237 (N_10237,N_5287,N_9760);
and U10238 (N_10238,N_6795,N_6242);
nand U10239 (N_10239,N_8699,N_6631);
nand U10240 (N_10240,N_8657,N_8442);
nor U10241 (N_10241,N_7904,N_9951);
xnor U10242 (N_10242,N_7117,N_9292);
nor U10243 (N_10243,N_6292,N_6814);
nand U10244 (N_10244,N_6393,N_6330);
xor U10245 (N_10245,N_8647,N_9225);
nand U10246 (N_10246,N_6441,N_6963);
or U10247 (N_10247,N_5738,N_8995);
xor U10248 (N_10248,N_9004,N_5468);
or U10249 (N_10249,N_5113,N_7475);
and U10250 (N_10250,N_8449,N_7357);
or U10251 (N_10251,N_5163,N_7370);
nor U10252 (N_10252,N_9369,N_5319);
xor U10253 (N_10253,N_8170,N_9013);
and U10254 (N_10254,N_7928,N_6883);
or U10255 (N_10255,N_9045,N_5665);
nand U10256 (N_10256,N_7255,N_5100);
nand U10257 (N_10257,N_9966,N_9403);
xor U10258 (N_10258,N_5549,N_8269);
and U10259 (N_10259,N_8611,N_9998);
nand U10260 (N_10260,N_8500,N_7077);
or U10261 (N_10261,N_5116,N_5009);
nor U10262 (N_10262,N_8814,N_5562);
nand U10263 (N_10263,N_9754,N_8128);
nand U10264 (N_10264,N_8824,N_8746);
nand U10265 (N_10265,N_7252,N_9611);
xnor U10266 (N_10266,N_7964,N_5528);
nor U10267 (N_10267,N_5253,N_5551);
nor U10268 (N_10268,N_9269,N_5636);
and U10269 (N_10269,N_8045,N_6183);
and U10270 (N_10270,N_6208,N_9632);
nand U10271 (N_10271,N_9633,N_8303);
xnor U10272 (N_10272,N_7995,N_7305);
and U10273 (N_10273,N_7639,N_5214);
and U10274 (N_10274,N_6666,N_9160);
or U10275 (N_10275,N_8244,N_6234);
and U10276 (N_10276,N_7931,N_7585);
or U10277 (N_10277,N_5224,N_5004);
nor U10278 (N_10278,N_8034,N_8282);
and U10279 (N_10279,N_6352,N_5257);
nor U10280 (N_10280,N_8205,N_6864);
nand U10281 (N_10281,N_7299,N_9246);
xnor U10282 (N_10282,N_6749,N_7899);
and U10283 (N_10283,N_5571,N_8707);
nor U10284 (N_10284,N_5807,N_5225);
nor U10285 (N_10285,N_5103,N_5221);
or U10286 (N_10286,N_5486,N_7499);
nand U10287 (N_10287,N_7708,N_8112);
and U10288 (N_10288,N_5559,N_7810);
xor U10289 (N_10289,N_9591,N_8724);
xnor U10290 (N_10290,N_9671,N_6975);
or U10291 (N_10291,N_9620,N_7812);
and U10292 (N_10292,N_8531,N_6509);
nor U10293 (N_10293,N_5201,N_7459);
nand U10294 (N_10294,N_5129,N_6554);
nor U10295 (N_10295,N_9383,N_7422);
nor U10296 (N_10296,N_9254,N_7212);
and U10297 (N_10297,N_9322,N_8830);
or U10298 (N_10298,N_8262,N_7770);
and U10299 (N_10299,N_6645,N_8377);
nand U10300 (N_10300,N_8599,N_5148);
nor U10301 (N_10301,N_7115,N_9639);
and U10302 (N_10302,N_6056,N_7019);
or U10303 (N_10303,N_5052,N_6487);
and U10304 (N_10304,N_9549,N_6113);
nand U10305 (N_10305,N_6656,N_8079);
or U10306 (N_10306,N_7125,N_8149);
and U10307 (N_10307,N_5268,N_8854);
or U10308 (N_10308,N_9400,N_7592);
nand U10309 (N_10309,N_8749,N_8238);
and U10310 (N_10310,N_6519,N_8989);
nor U10311 (N_10311,N_8865,N_5901);
and U10312 (N_10312,N_6207,N_6194);
nand U10313 (N_10313,N_7380,N_8974);
and U10314 (N_10314,N_7285,N_5683);
and U10315 (N_10315,N_8541,N_5439);
or U10316 (N_10316,N_9266,N_9204);
and U10317 (N_10317,N_6280,N_6411);
nor U10318 (N_10318,N_6471,N_9404);
nand U10319 (N_10319,N_9609,N_8929);
and U10320 (N_10320,N_6377,N_6596);
nand U10321 (N_10321,N_7097,N_7913);
nand U10322 (N_10322,N_5808,N_7270);
nor U10323 (N_10323,N_6924,N_7545);
nor U10324 (N_10324,N_8402,N_9454);
and U10325 (N_10325,N_5679,N_6436);
nand U10326 (N_10326,N_7867,N_6074);
or U10327 (N_10327,N_7725,N_5306);
and U10328 (N_10328,N_7169,N_9781);
and U10329 (N_10329,N_8862,N_9342);
xnor U10330 (N_10330,N_7395,N_9202);
nand U10331 (N_10331,N_6350,N_9062);
or U10332 (N_10332,N_5623,N_5726);
nand U10333 (N_10333,N_9883,N_6116);
nand U10334 (N_10334,N_9250,N_7109);
or U10335 (N_10335,N_7709,N_5656);
nand U10336 (N_10336,N_9836,N_8417);
or U10337 (N_10337,N_5602,N_6081);
nor U10338 (N_10338,N_8888,N_5058);
and U10339 (N_10339,N_8174,N_8080);
or U10340 (N_10340,N_6859,N_8185);
xor U10341 (N_10341,N_7287,N_9568);
or U10342 (N_10342,N_7298,N_5691);
or U10343 (N_10343,N_7732,N_7798);
or U10344 (N_10344,N_7534,N_5925);
and U10345 (N_10345,N_9389,N_7521);
xnor U10346 (N_10346,N_8290,N_7956);
xnor U10347 (N_10347,N_8543,N_7872);
xor U10348 (N_10348,N_7851,N_8420);
and U10349 (N_10349,N_8147,N_8492);
or U10350 (N_10350,N_5286,N_7719);
nand U10351 (N_10351,N_7759,N_7309);
nand U10352 (N_10352,N_9665,N_7978);
nor U10353 (N_10353,N_6822,N_7447);
or U10354 (N_10354,N_9877,N_5788);
nor U10355 (N_10355,N_5535,N_7093);
and U10356 (N_10356,N_5466,N_8392);
and U10357 (N_10357,N_9714,N_5881);
nand U10358 (N_10358,N_7460,N_7790);
and U10359 (N_10359,N_6816,N_5408);
and U10360 (N_10360,N_9846,N_6258);
and U10361 (N_10361,N_9053,N_9684);
or U10362 (N_10362,N_6223,N_7183);
nor U10363 (N_10363,N_8011,N_9955);
xor U10364 (N_10364,N_9486,N_9232);
or U10365 (N_10365,N_8982,N_9152);
or U10366 (N_10366,N_7157,N_5098);
nor U10367 (N_10367,N_9906,N_9521);
and U10368 (N_10368,N_8844,N_9598);
nor U10369 (N_10369,N_5332,N_8081);
xor U10370 (N_10370,N_8969,N_9150);
and U10371 (N_10371,N_5326,N_5708);
nor U10372 (N_10372,N_8216,N_5456);
nand U10373 (N_10373,N_6717,N_9502);
nor U10374 (N_10374,N_6679,N_8513);
and U10375 (N_10375,N_7827,N_8243);
nand U10376 (N_10376,N_8538,N_7520);
xor U10377 (N_10377,N_5136,N_6903);
nor U10378 (N_10378,N_5060,N_8029);
nor U10379 (N_10379,N_9120,N_6879);
and U10380 (N_10380,N_9497,N_8878);
nand U10381 (N_10381,N_7388,N_9871);
nor U10382 (N_10382,N_8237,N_5713);
nand U10383 (N_10383,N_5167,N_8390);
xnor U10384 (N_10384,N_8375,N_6641);
nand U10385 (N_10385,N_7750,N_9066);
xnor U10386 (N_10386,N_5234,N_7180);
nor U10387 (N_10387,N_5706,N_8326);
and U10388 (N_10388,N_5343,N_8100);
and U10389 (N_10389,N_5311,N_6185);
and U10390 (N_10390,N_8594,N_6849);
or U10391 (N_10391,N_9752,N_5830);
xnor U10392 (N_10392,N_7903,N_8587);
nand U10393 (N_10393,N_9930,N_9849);
and U10394 (N_10394,N_7567,N_9175);
xor U10395 (N_10395,N_6881,N_5482);
or U10396 (N_10396,N_5906,N_6488);
nand U10397 (N_10397,N_6747,N_8718);
or U10398 (N_10398,N_6156,N_6779);
or U10399 (N_10399,N_7957,N_7937);
nor U10400 (N_10400,N_9376,N_8478);
xnor U10401 (N_10401,N_5851,N_8848);
nor U10402 (N_10402,N_7986,N_6270);
or U10403 (N_10403,N_7908,N_7996);
nor U10404 (N_10404,N_8131,N_8965);
nand U10405 (N_10405,N_5765,N_7568);
nor U10406 (N_10406,N_9402,N_8005);
or U10407 (N_10407,N_9985,N_8321);
xor U10408 (N_10408,N_6310,N_8108);
nor U10409 (N_10409,N_9216,N_8428);
nor U10410 (N_10410,N_7189,N_6429);
xnor U10411 (N_10411,N_7675,N_8722);
and U10412 (N_10412,N_8890,N_7048);
nor U10413 (N_10413,N_5318,N_9869);
nand U10414 (N_10414,N_7431,N_8719);
and U10415 (N_10415,N_5447,N_8681);
nor U10416 (N_10416,N_6829,N_9970);
and U10417 (N_10417,N_5770,N_8528);
xnor U10418 (N_10418,N_9783,N_5379);
nand U10419 (N_10419,N_6705,N_7923);
and U10420 (N_10420,N_5130,N_6134);
nand U10421 (N_10421,N_5086,N_7102);
nor U10422 (N_10422,N_8958,N_5818);
xor U10423 (N_10423,N_9625,N_6061);
nand U10424 (N_10424,N_8906,N_6900);
nand U10425 (N_10425,N_5815,N_5870);
or U10426 (N_10426,N_7893,N_7419);
and U10427 (N_10427,N_8480,N_8404);
nand U10428 (N_10428,N_5761,N_6407);
nor U10429 (N_10429,N_8937,N_7229);
nand U10430 (N_10430,N_6101,N_8588);
or U10431 (N_10431,N_9029,N_9476);
nor U10432 (N_10432,N_8602,N_9720);
nand U10433 (N_10433,N_8612,N_5394);
nor U10434 (N_10434,N_5474,N_5315);
nor U10435 (N_10435,N_8204,N_7244);
and U10436 (N_10436,N_9142,N_9862);
or U10437 (N_10437,N_5349,N_7151);
or U10438 (N_10438,N_5158,N_8977);
nor U10439 (N_10439,N_5462,N_9678);
xor U10440 (N_10440,N_5337,N_5898);
xor U10441 (N_10441,N_7690,N_9272);
xor U10442 (N_10442,N_7181,N_7341);
or U10443 (N_10443,N_6427,N_6754);
xnor U10444 (N_10444,N_9165,N_5388);
and U10445 (N_10445,N_9954,N_7930);
xor U10446 (N_10446,N_6836,N_7949);
and U10447 (N_10447,N_9046,N_8771);
nor U10448 (N_10448,N_6178,N_9071);
nor U10449 (N_10449,N_5176,N_9230);
nand U10450 (N_10450,N_6718,N_7152);
nor U10451 (N_10451,N_8273,N_7074);
xnor U10452 (N_10452,N_5137,N_8737);
and U10453 (N_10453,N_6415,N_5283);
or U10454 (N_10454,N_6286,N_6338);
nand U10455 (N_10455,N_5596,N_7544);
or U10456 (N_10456,N_9014,N_9145);
and U10457 (N_10457,N_9787,N_7481);
xnor U10458 (N_10458,N_8772,N_6181);
nand U10459 (N_10459,N_8407,N_6815);
nor U10460 (N_10460,N_5036,N_7491);
or U10461 (N_10461,N_7007,N_8490);
or U10462 (N_10462,N_8115,N_5072);
xnor U10463 (N_10463,N_8936,N_7235);
or U10464 (N_10464,N_5639,N_9140);
or U10465 (N_10465,N_6648,N_9829);
and U10466 (N_10466,N_6837,N_8176);
or U10467 (N_10467,N_7050,N_9188);
nand U10468 (N_10468,N_8415,N_8498);
nand U10469 (N_10469,N_6985,N_7462);
xor U10470 (N_10470,N_8200,N_8884);
or U10471 (N_10471,N_6870,N_9179);
or U10472 (N_10472,N_6896,N_9401);
nor U10473 (N_10473,N_5125,N_8869);
nor U10474 (N_10474,N_7024,N_8674);
and U10475 (N_10475,N_8514,N_6760);
nor U10476 (N_10476,N_8438,N_5013);
xor U10477 (N_10477,N_8082,N_5586);
nand U10478 (N_10478,N_8361,N_6991);
and U10479 (N_10479,N_6316,N_6574);
nor U10480 (N_10480,N_7800,N_5628);
and U10481 (N_10481,N_9571,N_6793);
nand U10482 (N_10482,N_8740,N_6008);
and U10483 (N_10483,N_8834,N_5371);
xnor U10484 (N_10484,N_7013,N_5392);
and U10485 (N_10485,N_8441,N_6233);
xnor U10486 (N_10486,N_6326,N_8355);
and U10487 (N_10487,N_8137,N_6398);
or U10488 (N_10488,N_5374,N_8685);
nor U10489 (N_10489,N_8347,N_6148);
nand U10490 (N_10490,N_7143,N_9517);
or U10491 (N_10491,N_8314,N_9010);
and U10492 (N_10492,N_8654,N_5493);
xnor U10493 (N_10493,N_6511,N_7135);
nand U10494 (N_10494,N_7449,N_5428);
nor U10495 (N_10495,N_7717,N_7295);
and U10496 (N_10496,N_7494,N_8135);
nand U10497 (N_10497,N_6697,N_6702);
nor U10498 (N_10498,N_8923,N_8394);
xnor U10499 (N_10499,N_7705,N_5832);
or U10500 (N_10500,N_8136,N_9595);
nor U10501 (N_10501,N_8882,N_6506);
nand U10502 (N_10502,N_8468,N_8412);
xor U10503 (N_10503,N_5630,N_7665);
or U10504 (N_10504,N_5219,N_5750);
xor U10505 (N_10505,N_9685,N_5635);
nor U10506 (N_10506,N_5838,N_9080);
nor U10507 (N_10507,N_8246,N_7154);
xor U10508 (N_10508,N_6033,N_9200);
xnor U10509 (N_10509,N_7367,N_5569);
or U10510 (N_10510,N_6734,N_8800);
and U10511 (N_10511,N_5316,N_9637);
nor U10512 (N_10512,N_9351,N_9885);
and U10513 (N_10513,N_6560,N_7680);
and U10514 (N_10514,N_5395,N_7306);
nor U10515 (N_10515,N_9565,N_7952);
xnor U10516 (N_10516,N_8994,N_7948);
or U10517 (N_10517,N_5578,N_7535);
nand U10518 (N_10518,N_7066,N_5265);
nand U10519 (N_10519,N_6910,N_6027);
nor U10520 (N_10520,N_7078,N_6098);
or U10521 (N_10521,N_9548,N_7599);
nor U10522 (N_10522,N_6992,N_6823);
and U10523 (N_10523,N_9224,N_9527);
nor U10524 (N_10524,N_6567,N_6143);
or U10525 (N_10525,N_6887,N_9666);
nor U10526 (N_10526,N_5579,N_8895);
nand U10527 (N_10527,N_9159,N_7113);
or U10528 (N_10528,N_7221,N_9467);
or U10529 (N_10529,N_5357,N_8279);
and U10530 (N_10530,N_9026,N_9353);
and U10531 (N_10531,N_8463,N_6926);
nor U10532 (N_10532,N_8535,N_7259);
nor U10533 (N_10533,N_6818,N_5108);
xor U10534 (N_10534,N_5441,N_5975);
xnor U10535 (N_10535,N_8388,N_6969);
xnor U10536 (N_10536,N_9001,N_5654);
or U10537 (N_10537,N_7889,N_7549);
nor U10538 (N_10538,N_8350,N_9312);
nand U10539 (N_10539,N_8085,N_7988);
and U10540 (N_10540,N_8575,N_6681);
nand U10541 (N_10541,N_7932,N_9960);
xnor U10542 (N_10542,N_5198,N_8284);
nor U10543 (N_10543,N_5231,N_9493);
and U10544 (N_10544,N_9414,N_9385);
and U10545 (N_10545,N_8838,N_7809);
nand U10546 (N_10546,N_5415,N_8337);
and U10547 (N_10547,N_7631,N_6158);
nor U10548 (N_10548,N_8324,N_7947);
xnor U10549 (N_10549,N_5330,N_7440);
xnor U10550 (N_10550,N_9087,N_7683);
nand U10551 (N_10551,N_8306,N_5525);
or U10552 (N_10552,N_8519,N_9146);
nor U10553 (N_10553,N_9069,N_6604);
xor U10554 (N_10554,N_5444,N_7653);
xnor U10555 (N_10555,N_8452,N_9249);
and U10556 (N_10556,N_9429,N_9271);
xor U10557 (N_10557,N_5802,N_6387);
nor U10558 (N_10558,N_5055,N_5889);
or U10559 (N_10559,N_7959,N_6558);
nand U10560 (N_10560,N_9148,N_9287);
or U10561 (N_10561,N_6660,N_8107);
and U10562 (N_10562,N_9044,N_6709);
xnor U10563 (N_10563,N_7786,N_8360);
and U10564 (N_10564,N_7612,N_7057);
nor U10565 (N_10565,N_6247,N_6278);
and U10566 (N_10566,N_9949,N_6755);
and U10567 (N_10567,N_6126,N_6727);
nand U10568 (N_10568,N_6585,N_8121);
nand U10569 (N_10569,N_7442,N_5854);
nand U10570 (N_10570,N_7248,N_8686);
xnor U10571 (N_10571,N_7327,N_5771);
xnor U10572 (N_10572,N_5012,N_6227);
or U10573 (N_10573,N_8353,N_6226);
nand U10574 (N_10574,N_5577,N_9555);
or U10575 (N_10575,N_8250,N_8055);
nor U10576 (N_10576,N_7153,N_5966);
nand U10577 (N_10577,N_5798,N_6742);
nor U10578 (N_10578,N_9349,N_6993);
nand U10579 (N_10579,N_5341,N_9355);
and U10580 (N_10580,N_5160,N_6322);
and U10581 (N_10581,N_8631,N_7421);
and U10582 (N_10582,N_6414,N_5776);
or U10583 (N_10583,N_5969,N_8051);
and U10584 (N_10584,N_9931,N_6582);
xnor U10585 (N_10585,N_5576,N_8127);
or U10586 (N_10586,N_6346,N_6540);
nand U10587 (N_10587,N_5347,N_5285);
nand U10588 (N_10588,N_6391,N_9487);
xor U10589 (N_10589,N_9100,N_8601);
and U10590 (N_10590,N_5047,N_7624);
and U10591 (N_10591,N_5585,N_8159);
or U10592 (N_10592,N_6007,N_7399);
nor U10593 (N_10593,N_8195,N_9988);
or U10594 (N_10594,N_6695,N_5553);
and U10595 (N_10595,N_8031,N_7763);
xor U10596 (N_10596,N_6384,N_6848);
nor U10597 (N_10597,N_6844,N_5711);
and U10598 (N_10598,N_7519,N_8985);
nand U10599 (N_10599,N_7630,N_7407);
nor U10600 (N_10600,N_6899,N_8172);
and U10601 (N_10601,N_6004,N_5420);
or U10602 (N_10602,N_9068,N_7608);
xor U10603 (N_10603,N_8979,N_8544);
or U10604 (N_10604,N_5521,N_9757);
nand U10605 (N_10605,N_9466,N_9969);
and U10606 (N_10606,N_8453,N_9161);
nor U10607 (N_10607,N_5199,N_5719);
and U10608 (N_10608,N_7245,N_8605);
xor U10609 (N_10609,N_9870,N_7124);
nor U10610 (N_10610,N_9992,N_5296);
nor U10611 (N_10611,N_6947,N_6842);
nand U10612 (N_10612,N_5135,N_8886);
or U10613 (N_10613,N_6087,N_9631);
or U10614 (N_10614,N_6917,N_9275);
nand U10615 (N_10615,N_7003,N_8305);
and U10616 (N_10616,N_5117,N_5418);
nor U10617 (N_10617,N_7318,N_5155);
xor U10618 (N_10618,N_8827,N_7283);
nor U10619 (N_10619,N_8373,N_6773);
or U10620 (N_10620,N_9734,N_7161);
nand U10621 (N_10621,N_5206,N_7051);
and U10622 (N_10622,N_6039,N_9798);
nor U10623 (N_10623,N_7640,N_5558);
xnor U10624 (N_10624,N_8240,N_8239);
nor U10625 (N_10625,N_8348,N_8821);
nor U10626 (N_10626,N_9330,N_8156);
nand U10627 (N_10627,N_5104,N_6867);
and U10628 (N_10628,N_6335,N_7312);
nand U10629 (N_10629,N_7091,N_8713);
nor U10630 (N_10630,N_5650,N_5397);
nand U10631 (N_10631,N_5941,N_5262);
and U10632 (N_10632,N_9696,N_7940);
nor U10633 (N_10633,N_7525,N_7678);
or U10634 (N_10634,N_8294,N_8596);
nor U10635 (N_10635,N_6677,N_6502);
nor U10636 (N_10636,N_9205,N_8008);
and U10637 (N_10637,N_9624,N_6264);
nand U10638 (N_10638,N_5840,N_7813);
nand U10639 (N_10639,N_7338,N_5422);
nand U10640 (N_10640,N_6606,N_6521);
xnor U10641 (N_10641,N_5839,N_6382);
xor U10642 (N_10642,N_5928,N_8432);
xnor U10643 (N_10643,N_9890,N_5624);
xor U10644 (N_10644,N_5603,N_5477);
nor U10645 (N_10645,N_7512,N_8257);
nand U10646 (N_10646,N_5744,N_7658);
nand U10647 (N_10647,N_8625,N_8649);
and U10648 (N_10648,N_5409,N_9842);
xnor U10649 (N_10649,N_7776,N_9452);
nor U10650 (N_10650,N_5062,N_6221);
xnor U10651 (N_10651,N_8125,N_6714);
xnor U10652 (N_10652,N_5254,N_7580);
or U10653 (N_10653,N_6858,N_9673);
or U10654 (N_10654,N_7972,N_5519);
nor U10655 (N_10655,N_9722,N_5986);
xnor U10656 (N_10656,N_5412,N_9654);
nor U10657 (N_10657,N_7984,N_5492);
or U10658 (N_10658,N_9642,N_6798);
nor U10659 (N_10659,N_6796,N_5896);
xnor U10660 (N_10660,N_5173,N_8162);
nor U10661 (N_10661,N_5340,N_9856);
xnor U10662 (N_10662,N_6751,N_5096);
and U10663 (N_10663,N_7182,N_9105);
and U10664 (N_10664,N_7017,N_9333);
nor U10665 (N_10665,N_5220,N_7945);
nor U10666 (N_10666,N_5999,N_8329);
and U10667 (N_10667,N_9668,N_5517);
or U10668 (N_10668,N_8369,N_5512);
and U10669 (N_10669,N_8446,N_8557);
nand U10670 (N_10670,N_7303,N_7569);
or U10671 (N_10671,N_6389,N_7504);
nor U10672 (N_10672,N_6535,N_7748);
nor U10673 (N_10673,N_6657,N_6452);
nand U10674 (N_10674,N_8518,N_6674);
or U10675 (N_10675,N_6328,N_5526);
nand U10676 (N_10676,N_6110,N_7818);
and U10677 (N_10677,N_7122,N_9426);
nand U10678 (N_10678,N_5681,N_5511);
or U10679 (N_10679,N_7574,N_8883);
nor U10680 (N_10680,N_8880,N_7939);
and U10681 (N_10681,N_9413,N_7749);
xor U10682 (N_10682,N_5695,N_7533);
nor U10683 (N_10683,N_5692,N_7429);
nor U10684 (N_10684,N_7423,N_5967);
or U10685 (N_10685,N_6342,N_9117);
xor U10686 (N_10686,N_8617,N_9037);
and U10687 (N_10687,N_8754,N_8267);
or U10688 (N_10688,N_8098,N_5613);
xor U10689 (N_10689,N_6381,N_8778);
nand U10690 (N_10690,N_8122,N_6371);
nand U10691 (N_10691,N_8828,N_6220);
nand U10692 (N_10692,N_9826,N_8474);
xor U10693 (N_10693,N_7992,N_5368);
xnor U10694 (N_10694,N_8119,N_9552);
and U10695 (N_10695,N_5450,N_5631);
nand U10696 (N_10696,N_9370,N_9570);
and U10697 (N_10697,N_7156,N_8228);
or U10698 (N_10698,N_7120,N_6047);
xor U10699 (N_10699,N_9346,N_5165);
and U10700 (N_10700,N_9582,N_7246);
xor U10701 (N_10701,N_5594,N_6137);
xnor U10702 (N_10702,N_9910,N_7935);
xnor U10703 (N_10703,N_5714,N_8427);
or U10704 (N_10704,N_5475,N_7401);
or U10705 (N_10705,N_5976,N_6029);
nand U10706 (N_10706,N_6484,N_9586);
and U10707 (N_10707,N_7649,N_8871);
or U10708 (N_10708,N_6981,N_8623);
or U10709 (N_10709,N_8059,N_6201);
xnor U10710 (N_10710,N_7901,N_5943);
and U10711 (N_10711,N_6165,N_7272);
or U10712 (N_10712,N_7014,N_5581);
nand U10713 (N_10713,N_7377,N_9154);
and U10714 (N_10714,N_6933,N_5025);
nor U10715 (N_10715,N_6620,N_7970);
nand U10716 (N_10716,N_6334,N_8760);
nor U10717 (N_10717,N_7636,N_5972);
and U10718 (N_10718,N_8577,N_9940);
or U10719 (N_10719,N_6962,N_5520);
or U10720 (N_10720,N_6825,N_6465);
nand U10721 (N_10721,N_9381,N_6493);
xor U10722 (N_10722,N_5997,N_5588);
and U10723 (N_10723,N_9830,N_5687);
and U10724 (N_10724,N_9278,N_9525);
xnor U10725 (N_10725,N_6416,N_5754);
nor U10726 (N_10726,N_9326,N_9114);
and U10727 (N_10727,N_7238,N_9816);
nand U10728 (N_10728,N_9675,N_7562);
nor U10729 (N_10729,N_8464,N_8286);
xnor U10730 (N_10730,N_5842,N_6425);
nand U10731 (N_10731,N_7538,N_8167);
or U10732 (N_10732,N_7752,N_8712);
nand U10733 (N_10733,N_5865,N_9164);
nand U10734 (N_10734,N_7375,N_5038);
nor U10735 (N_10735,N_8992,N_8723);
and U10736 (N_10736,N_6989,N_6164);
or U10737 (N_10737,N_9544,N_7203);
and U10738 (N_10738,N_6230,N_7042);
or U10739 (N_10739,N_6592,N_9896);
nand U10740 (N_10740,N_8214,N_8970);
or U10741 (N_10741,N_8401,N_9975);
or U10742 (N_10742,N_6833,N_5859);
xor U10743 (N_10743,N_5856,N_6546);
nor U10744 (N_10744,N_9669,N_6118);
nor U10745 (N_10745,N_6557,N_8680);
or U10746 (N_10746,N_5834,N_7542);
and U10747 (N_10747,N_8986,N_6281);
and U10748 (N_10748,N_6069,N_6504);
and U10749 (N_10749,N_8276,N_6262);
nand U10750 (N_10750,N_7981,N_6252);
nand U10751 (N_10751,N_7137,N_8489);
nand U10752 (N_10752,N_6812,N_7464);
nand U10753 (N_10753,N_6649,N_6359);
and U10754 (N_10754,N_8050,N_9063);
nand U10755 (N_10755,N_7967,N_8226);
nand U10756 (N_10756,N_6482,N_9894);
nor U10757 (N_10757,N_6895,N_9127);
and U10758 (N_10758,N_6277,N_6999);
nor U10759 (N_10759,N_5077,N_8738);
or U10760 (N_10760,N_8510,N_9314);
nor U10761 (N_10761,N_5950,N_8311);
nand U10762 (N_10762,N_7755,N_9875);
and U10763 (N_10763,N_9613,N_6269);
nor U10764 (N_10764,N_8990,N_6257);
nor U10765 (N_10765,N_7563,N_9615);
nand U10766 (N_10766,N_9268,N_6497);
or U10767 (N_10767,N_9968,N_9759);
xor U10768 (N_10768,N_6145,N_9448);
nor U10769 (N_10769,N_6267,N_6423);
nand U10770 (N_10770,N_6402,N_9392);
or U10771 (N_10771,N_6049,N_9513);
nand U10772 (N_10772,N_5406,N_9107);
or U10773 (N_10773,N_8413,N_7110);
and U10774 (N_10774,N_7858,N_5736);
or U10775 (N_10775,N_9815,N_9494);
xnor U10776 (N_10776,N_8781,N_9102);
nand U10777 (N_10777,N_6813,N_6408);
or U10778 (N_10778,N_8365,N_6348);
nor U10779 (N_10779,N_5161,N_9768);
xnor U10780 (N_10780,N_9808,N_8497);
or U10781 (N_10781,N_6096,N_9925);
nor U10782 (N_10782,N_7470,N_9409);
or U10783 (N_10783,N_9599,N_7493);
or U10784 (N_10784,N_8318,N_5880);
nand U10785 (N_10785,N_6140,N_8473);
nand U10786 (N_10786,N_9410,N_7771);
and U10787 (N_10787,N_5638,N_9662);
and U10788 (N_10788,N_7938,N_7779);
or U10789 (N_10789,N_6799,N_7894);
nor U10790 (N_10790,N_8440,N_5615);
nand U10791 (N_10791,N_6122,N_7643);
and U10792 (N_10792,N_7188,N_7046);
nand U10793 (N_10793,N_6501,N_9186);
xor U10794 (N_10794,N_7289,N_8777);
or U10795 (N_10795,N_5479,N_5933);
or U10796 (N_10796,N_9770,N_5236);
or U10797 (N_10797,N_8720,N_5495);
nand U10798 (N_10798,N_9450,N_6189);
nor U10799 (N_10799,N_5048,N_8730);
and U10800 (N_10800,N_6959,N_5405);
nor U10801 (N_10801,N_8659,N_6299);
and U10802 (N_10802,N_5041,N_7159);
nand U10803 (N_10803,N_9581,N_7976);
or U10804 (N_10804,N_6196,N_9185);
nand U10805 (N_10805,N_8624,N_5484);
and U10806 (N_10806,N_5868,N_8567);
nor U10807 (N_10807,N_5164,N_6055);
nand U10808 (N_10808,N_8922,N_6807);
and U10809 (N_10809,N_6544,N_6706);
and U10810 (N_10810,N_8481,N_6591);
or U10811 (N_10811,N_9422,N_8944);
and U10812 (N_10812,N_9260,N_5404);
nand U10813 (N_10813,N_8833,N_9766);
or U10814 (N_10814,N_8218,N_9649);
xor U10815 (N_10815,N_5501,N_6160);
or U10816 (N_10816,N_9811,N_7079);
and U10817 (N_10817,N_9991,N_8173);
xor U10818 (N_10818,N_5769,N_6720);
and U10819 (N_10819,N_6668,N_8391);
or U10820 (N_10820,N_7974,N_8765);
nand U10821 (N_10821,N_6001,N_7747);
or U10822 (N_10822,N_8217,N_7551);
and U10823 (N_10823,N_5912,N_8146);
nand U10824 (N_10824,N_5704,N_6037);
nor U10825 (N_10825,N_7023,N_5448);
and U10826 (N_10826,N_9608,N_8806);
nor U10827 (N_10827,N_6534,N_5796);
or U10828 (N_10828,N_7065,N_8234);
nor U10829 (N_10829,N_6472,N_9593);
xor U10830 (N_10830,N_9723,N_9867);
and U10831 (N_10831,N_8134,N_9805);
nor U10832 (N_10832,N_5949,N_6791);
or U10833 (N_10833,N_5888,N_6093);
xnor U10834 (N_10834,N_6811,N_7603);
xor U10835 (N_10835,N_8256,N_8924);
nand U10836 (N_10836,N_6780,N_8656);
xor U10837 (N_10837,N_8184,N_8589);
xor U10838 (N_10838,N_7728,N_9226);
or U10839 (N_10839,N_6528,N_7651);
and U10840 (N_10840,N_9861,N_9559);
xnor U10841 (N_10841,N_9178,N_8456);
and U10842 (N_10842,N_8843,N_9365);
or U10843 (N_10843,N_9267,N_9545);
or U10844 (N_10844,N_8123,N_7479);
nor U10845 (N_10845,N_9698,N_9373);
nand U10846 (N_10846,N_9504,N_7253);
and U10847 (N_10847,N_8938,N_7015);
or U10848 (N_10848,N_9055,N_8088);
nand U10849 (N_10849,N_7616,N_6765);
nor U10850 (N_10850,N_5232,N_9380);
nand U10851 (N_10851,N_5333,N_7950);
nor U10852 (N_10852,N_7398,N_5755);
and U10853 (N_10853,N_6272,N_8018);
or U10854 (N_10854,N_6430,N_5611);
nand U10855 (N_10855,N_6901,N_6897);
nand U10856 (N_10856,N_5153,N_9602);
or U10857 (N_10857,N_6147,N_6480);
or U10858 (N_10858,N_6440,N_5867);
or U10859 (N_10859,N_6982,N_6058);
and U10860 (N_10860,N_6130,N_5866);
and U10861 (N_10861,N_5678,N_8630);
xnor U10862 (N_10862,N_5186,N_6428);
and U10863 (N_10863,N_8301,N_7987);
or U10864 (N_10864,N_9364,N_5223);
and U10865 (N_10865,N_8583,N_9819);
nand U10866 (N_10866,N_7762,N_5689);
nand U10867 (N_10867,N_6573,N_8444);
nand U10868 (N_10868,N_8052,N_9075);
nand U10869 (N_10869,N_6514,N_8275);
nand U10870 (N_10870,N_7558,N_8545);
nand U10871 (N_10871,N_5476,N_9860);
nand U10872 (N_10872,N_8183,N_7379);
and U10873 (N_10873,N_7069,N_8287);
nor U10874 (N_10874,N_9804,N_9455);
nor U10875 (N_10875,N_6139,N_5269);
nor U10876 (N_10876,N_6020,N_5342);
nor U10877 (N_10877,N_8919,N_7346);
and U10878 (N_10878,N_6939,N_7211);
xor U10879 (N_10879,N_7269,N_7679);
nor U10880 (N_10880,N_7735,N_9139);
nor U10881 (N_10881,N_9532,N_8117);
nand U10882 (N_10882,N_8110,N_5276);
nand U10883 (N_10883,N_5378,N_8225);
and U10884 (N_10884,N_7173,N_8140);
xor U10885 (N_10885,N_9984,N_6520);
xnor U10886 (N_10886,N_8068,N_6675);
nor U10887 (N_10887,N_6863,N_5454);
nand U10888 (N_10888,N_8915,N_8876);
xnor U10889 (N_10889,N_9750,N_8914);
and U10890 (N_10890,N_6726,N_7971);
nand U10891 (N_10891,N_7339,N_5288);
xnor U10892 (N_10892,N_7826,N_8539);
nor U10893 (N_10893,N_7857,N_9096);
and U10894 (N_10894,N_7273,N_6576);
xor U10895 (N_10895,N_9441,N_8679);
xnor U10896 (N_10896,N_8930,N_9999);
or U10897 (N_10897,N_8753,N_8352);
and U10898 (N_10898,N_9371,N_6360);
or U10899 (N_10899,N_5601,N_6032);
nand U10900 (N_10900,N_7284,N_6994);
nand U10901 (N_10901,N_5582,N_6224);
xnor U10902 (N_10902,N_5189,N_7333);
xnor U10903 (N_10903,N_5339,N_5707);
and U10904 (N_10904,N_9082,N_6547);
and U10905 (N_10905,N_9705,N_6759);
or U10906 (N_10906,N_8560,N_5660);
nand U10907 (N_10907,N_8083,N_5774);
or U10908 (N_10908,N_5955,N_8870);
nand U10909 (N_10909,N_7134,N_5964);
xnor U10910 (N_10910,N_9658,N_9039);
and U10911 (N_10911,N_8555,N_5266);
xor U10912 (N_10912,N_9073,N_6854);
and U10913 (N_10913,N_7635,N_7260);
nand U10914 (N_10914,N_9737,N_8773);
nand U10915 (N_10915,N_6613,N_9446);
xnor U10916 (N_10916,N_9813,N_9741);
nor U10917 (N_10917,N_6291,N_7450);
or U10918 (N_10918,N_9688,N_6454);
nand U10919 (N_10919,N_7076,N_9746);
xnor U10920 (N_10920,N_9097,N_5112);
nand U10921 (N_10921,N_8030,N_9406);
and U10922 (N_10922,N_6715,N_8411);
or U10923 (N_10923,N_8399,N_6638);
xnor U10924 (N_10924,N_8454,N_8124);
or U10925 (N_10925,N_6378,N_9270);
xnor U10926 (N_10926,N_5875,N_8874);
xor U10927 (N_10927,N_9309,N_5688);
or U10928 (N_10928,N_8455,N_9032);
xnor U10929 (N_10929,N_5216,N_7413);
or U10930 (N_10930,N_5543,N_6498);
nor U10931 (N_10931,N_7011,N_9822);
and U10932 (N_10932,N_5377,N_5893);
xnor U10933 (N_10933,N_7418,N_8744);
nand U10934 (N_10934,N_6581,N_7960);
nand U10935 (N_10935,N_8168,N_5973);
nor U10936 (N_10936,N_5723,N_6123);
xnor U10937 (N_10937,N_6655,N_9656);
nand U10938 (N_10938,N_5279,N_5752);
nand U10939 (N_10939,N_5204,N_9927);
or U10940 (N_10940,N_9218,N_5156);
and U10941 (N_10941,N_5358,N_7575);
and U10942 (N_10942,N_6703,N_8302);
nor U10943 (N_10943,N_5095,N_8221);
xnor U10944 (N_10944,N_5449,N_9795);
and U10945 (N_10945,N_8585,N_8179);
nor U10946 (N_10946,N_7308,N_6282);
xor U10947 (N_10947,N_8726,N_9835);
nor U10948 (N_10948,N_5127,N_7620);
nor U10949 (N_10949,N_8434,N_8775);
xor U10950 (N_10950,N_5836,N_6626);
and U10951 (N_10951,N_8296,N_9745);
xor U10952 (N_10952,N_6707,N_9317);
nand U10953 (N_10953,N_7480,N_5375);
or U10954 (N_10954,N_7618,N_6297);
xor U10955 (N_10955,N_5690,N_8808);
or U10956 (N_10956,N_7794,N_5344);
xor U10957 (N_10957,N_8948,N_5015);
or U10958 (N_10958,N_5364,N_7430);
xor U10959 (N_10959,N_9498,N_9118);
nor U10960 (N_10960,N_6752,N_8036);
xnor U10961 (N_10961,N_6155,N_8540);
nor U10962 (N_10962,N_5150,N_9458);
or U10963 (N_10963,N_5233,N_6362);
or U10964 (N_10964,N_5367,N_6228);
nor U10965 (N_10965,N_8281,N_8857);
or U10966 (N_10966,N_5676,N_8939);
or U10967 (N_10967,N_8570,N_7405);
nor U10968 (N_10968,N_7804,N_7953);
nand U10969 (N_10969,N_8934,N_9884);
nor U10970 (N_10970,N_8748,N_9807);
or U10971 (N_10971,N_9101,N_8357);
nor U10972 (N_10972,N_5816,N_6575);
and U10973 (N_10973,N_7095,N_8408);
nand U10974 (N_10974,N_8253,N_6723);
nand U10975 (N_10975,N_6672,N_7830);
or U10976 (N_10976,N_9967,N_8715);
nor U10977 (N_10977,N_9702,N_8342);
or U10978 (N_10978,N_7150,N_5238);
nor U10979 (N_10979,N_8009,N_5937);
or U10980 (N_10980,N_6026,N_5436);
and U10981 (N_10981,N_6970,N_5106);
or U10982 (N_10982,N_9732,N_6132);
nor U10983 (N_10983,N_6486,N_5620);
or U10984 (N_10984,N_5413,N_8792);
xor U10985 (N_10985,N_6456,N_9284);
and U10986 (N_10986,N_7233,N_6323);
nand U10987 (N_10987,N_5824,N_9897);
nand U10988 (N_10988,N_7206,N_5931);
nor U10989 (N_10989,N_6724,N_7254);
or U10990 (N_10990,N_6625,N_9784);
or U10991 (N_10991,N_7887,N_6345);
nor U10992 (N_10992,N_5978,N_6663);
xnor U10993 (N_10993,N_5118,N_8634);
nand U10994 (N_10994,N_5019,N_5191);
and U10995 (N_10995,N_8887,N_9651);
nand U10996 (N_10996,N_5350,N_8371);
xnor U10997 (N_10997,N_6083,N_8751);
nor U10998 (N_10998,N_6128,N_6319);
or U10999 (N_10999,N_5366,N_5640);
xnor U11000 (N_11000,N_9630,N_5121);
nor U11001 (N_11001,N_7342,N_6904);
nand U11002 (N_11002,N_5497,N_8109);
or U11003 (N_11003,N_7032,N_5151);
xnor U11004 (N_11004,N_6632,N_5390);
or U11005 (N_11005,N_8046,N_8770);
nor U11006 (N_11006,N_5938,N_8152);
or U11007 (N_11007,N_6686,N_8133);
xnor U11008 (N_11008,N_9193,N_6928);
nand U11009 (N_11009,N_8258,N_8437);
xor U11010 (N_11010,N_8633,N_5790);
and U11011 (N_11011,N_9206,N_5981);
and U11012 (N_11012,N_8932,N_5758);
or U11013 (N_11013,N_5573,N_7865);
nor U11014 (N_11014,N_7581,N_6593);
xor U11015 (N_11015,N_9686,N_5954);
nor U11016 (N_11016,N_7081,N_5682);
or U11017 (N_11017,N_9111,N_7710);
nand U11018 (N_11018,N_6447,N_6432);
or U11019 (N_11019,N_7121,N_9341);
and U11020 (N_11020,N_5853,N_5823);
xnor U11021 (N_11021,N_7034,N_5721);
nor U11022 (N_11022,N_8526,N_6021);
and U11023 (N_11023,N_9786,N_6925);
nor U11024 (N_11024,N_6894,N_9712);
or U11025 (N_11025,N_5452,N_9098);
xor U11026 (N_11026,N_6240,N_6249);
nor U11027 (N_11027,N_8676,N_7989);
xnor U11028 (N_11028,N_7432,N_8551);
xor U11029 (N_11029,N_8696,N_7980);
xor U11030 (N_11030,N_8867,N_7408);
and U11031 (N_11031,N_8422,N_9038);
and U11032 (N_11032,N_7364,N_9888);
nor U11033 (N_11033,N_8141,N_7571);
nand U11034 (N_11034,N_7875,N_7446);
and U11035 (N_11035,N_5195,N_9077);
or U11036 (N_11036,N_9468,N_8040);
nor U11037 (N_11037,N_9853,N_5820);
and U11038 (N_11038,N_9180,N_8762);
or U11039 (N_11039,N_6490,N_9334);
nor U11040 (N_11040,N_5686,N_6150);
xor U11041 (N_11041,N_7508,N_5789);
xor U11042 (N_11042,N_7317,N_8479);
nor U11043 (N_11043,N_9913,N_5458);
nor U11044 (N_11044,N_7410,N_7600);
xor U11045 (N_11045,N_5606,N_9310);
and U11046 (N_11046,N_7803,N_6298);
or U11047 (N_11047,N_5304,N_8683);
nor U11048 (N_11048,N_5490,N_9143);
and U11049 (N_11049,N_8774,N_9792);
or U11050 (N_11050,N_9394,N_5414);
and U11051 (N_11051,N_6308,N_7514);
or U11052 (N_11052,N_5197,N_8786);
nor U11053 (N_11053,N_5716,N_6781);
xnor U11054 (N_11054,N_9214,N_6966);
nand U11055 (N_11055,N_9338,N_6516);
or U11056 (N_11056,N_9879,N_7455);
and U11057 (N_11057,N_5322,N_8171);
or U11058 (N_11058,N_8527,N_9464);
nand U11059 (N_11059,N_8758,N_7251);
and U11060 (N_11060,N_8158,N_6210);
xnor U11061 (N_11061,N_5119,N_5852);
nor U11062 (N_11062,N_5927,N_8988);
and U11063 (N_11063,N_8166,N_8734);
and U11064 (N_11064,N_9667,N_7332);
nand U11065 (N_11065,N_9424,N_6064);
and U11066 (N_11066,N_5314,N_6294);
nand U11067 (N_11067,N_6102,N_6141);
nor U11068 (N_11068,N_8235,N_5494);
and U11069 (N_11069,N_9993,N_5764);
nor U11070 (N_11070,N_6500,N_6590);
or U11071 (N_11071,N_6287,N_5508);
or U11072 (N_11072,N_8013,N_6929);
and U11073 (N_11073,N_8433,N_8946);
xor U11074 (N_11074,N_5403,N_8664);
xnor U11075 (N_11075,N_7745,N_5670);
nand U11076 (N_11076,N_6045,N_9477);
or U11077 (N_11077,N_5207,N_5819);
xor U11078 (N_11078,N_9438,N_6696);
xor U11079 (N_11079,N_6512,N_9605);
or U11080 (N_11080,N_7929,N_8073);
or U11081 (N_11081,N_9484,N_7905);
nand U11082 (N_11082,N_7082,N_9405);
and U11083 (N_11083,N_9378,N_7368);
xnor U11084 (N_11084,N_5084,N_8426);
and U11085 (N_11085,N_6344,N_6997);
or U11086 (N_11086,N_8629,N_8835);
or U11087 (N_11087,N_8466,N_9059);
nand U11088 (N_11088,N_7315,N_7743);
nand U11089 (N_11089,N_7214,N_6478);
nor U11090 (N_11090,N_7582,N_9199);
nor U11091 (N_11091,N_8668,N_9276);
and U11092 (N_11092,N_9375,N_9223);
nand U11093 (N_11093,N_9574,N_5031);
nor U11094 (N_11094,N_6986,N_9511);
xnor U11095 (N_11095,N_5473,N_7787);
or U11096 (N_11096,N_6159,N_5323);
or U11097 (N_11097,N_9245,N_6157);
or U11098 (N_11098,N_7993,N_7373);
nand U11099 (N_11099,N_9361,N_8548);
or U11100 (N_11100,N_9626,N_5417);
nand U11101 (N_11101,N_8955,N_7148);
and U11102 (N_11102,N_8202,N_5053);
nor U11103 (N_11103,N_6803,N_6129);
nand U11104 (N_11104,N_8071,N_8702);
or U11105 (N_11105,N_5760,N_7386);
and U11106 (N_11106,N_6168,N_5090);
nand U11107 (N_11107,N_9905,N_8616);
nor U11108 (N_11108,N_9231,N_5046);
and U11109 (N_11109,N_8520,N_7144);
and U11110 (N_11110,N_9743,N_5622);
and U11111 (N_11111,N_5627,N_6339);
and U11112 (N_11112,N_9584,N_6783);
nand U11113 (N_11113,N_6721,N_8191);
or U11114 (N_11114,N_9453,N_6048);
xor U11115 (N_11115,N_7766,N_8090);
xor U11116 (N_11116,N_5961,N_5730);
xor U11117 (N_11117,N_9771,N_6217);
xor U11118 (N_11118,N_5218,N_7687);
or U11119 (N_11119,N_7712,N_9818);
or U11120 (N_11120,N_7841,N_8389);
nor U11121 (N_11121,N_6167,N_6944);
or U11122 (N_11122,N_6579,N_5252);
and U11123 (N_11123,N_5728,N_5245);
nor U11124 (N_11124,N_7132,N_7358);
xor U11125 (N_11125,N_9474,N_6204);
xor U11126 (N_11126,N_7811,N_9289);
xor U11127 (N_11127,N_7268,N_9109);
xor U11128 (N_11128,N_7669,N_6964);
or U11129 (N_11129,N_8805,N_7644);
or U11130 (N_11130,N_9834,N_9419);
and U11131 (N_11131,N_6354,N_7343);
or U11132 (N_11132,N_8957,N_6898);
or U11133 (N_11133,N_9790,N_5629);
nand U11134 (N_11134,N_6598,N_5376);
or U11135 (N_11135,N_7829,N_7632);
and U11136 (N_11136,N_5369,N_5022);
nand U11137 (N_11137,N_5061,N_8603);
and U11138 (N_11138,N_6361,N_7009);
nand U11139 (N_11139,N_7411,N_8065);
and U11140 (N_11140,N_9196,N_5659);
and U11141 (N_11141,N_9354,N_8120);
xnor U11142 (N_11142,N_5987,N_9471);
nand U11143 (N_11143,N_7345,N_6809);
and U11144 (N_11144,N_8829,N_7704);
nor U11145 (N_11145,N_5081,N_6564);
xor U11146 (N_11146,N_6733,N_5786);
xnor U11147 (N_11147,N_6802,N_5334);
and U11148 (N_11148,N_8248,N_8378);
nand U11149 (N_11149,N_9755,N_7595);
xnor U11150 (N_11150,N_8328,N_6005);
nor U11151 (N_11151,N_9601,N_5181);
and U11152 (N_11152,N_8728,N_7584);
nand U11153 (N_11153,N_7424,N_8802);
nand U11154 (N_11154,N_5398,N_8590);
nor U11155 (N_11155,N_6778,N_6011);
and U11156 (N_11156,N_6379,N_8255);
xor U11157 (N_11157,N_5434,N_7529);
or U11158 (N_11158,N_9579,N_8750);
and U11159 (N_11159,N_6095,N_7662);
nand U11160 (N_11160,N_8445,N_6107);
nand U11161 (N_11161,N_5655,N_6434);
xnor U11162 (N_11162,N_7622,N_6317);
nand U11163 (N_11163,N_7412,N_6082);
or U11164 (N_11164,N_8691,N_9716);
nand U11165 (N_11165,N_5825,N_5604);
or U11166 (N_11166,N_9529,N_5033);
nor U11167 (N_11167,N_5259,N_5251);
and U11168 (N_11168,N_5465,N_8998);
and U11169 (N_11169,N_9749,N_6555);
nor U11170 (N_11170,N_9265,N_7098);
nor U11171 (N_11171,N_5183,N_8554);
nand U11172 (N_11172,N_5430,N_5909);
and U11173 (N_11173,N_7096,N_5290);
or U11174 (N_11174,N_6757,N_9473);
or U11175 (N_11175,N_6301,N_7839);
nand U11176 (N_11176,N_9537,N_6405);
nor U11177 (N_11177,N_6314,N_7129);
nor U11178 (N_11178,N_7397,N_8613);
nand U11179 (N_11179,N_7292,N_6420);
nor U11180 (N_11180,N_8346,N_8972);
nand U11181 (N_11181,N_6103,N_5074);
or U11182 (N_11182,N_8529,N_7614);
nor U11183 (N_11183,N_6700,N_5099);
xor U11184 (N_11184,N_8245,N_9907);
nand U11185 (N_11185,N_5560,N_8154);
or U11186 (N_11186,N_7816,N_8229);
and U11187 (N_11187,N_8637,N_9617);
and U11188 (N_11188,N_5827,N_6831);
or U11189 (N_11189,N_8297,N_9881);
nand U11190 (N_11190,N_9033,N_9515);
nor U11191 (N_11191,N_9797,N_8571);
or U11192 (N_11192,N_6358,N_5264);
or U11193 (N_11193,N_8354,N_5437);
xor U11194 (N_11194,N_6847,N_6468);
nor U11195 (N_11195,N_6691,N_8021);
xor U11196 (N_11196,N_6594,N_5563);
xnor U11197 (N_11197,N_7043,N_5609);
xnor U11198 (N_11198,N_6495,N_8484);
or U11199 (N_11199,N_8701,N_7164);
nand U11200 (N_11200,N_9091,N_9980);
nor U11201 (N_11201,N_6105,N_5391);
nand U11202 (N_11202,N_7103,N_5564);
xnor U11203 (N_11203,N_6311,N_9336);
xor U11204 (N_11204,N_8211,N_7222);
nand U11205 (N_11205,N_8987,N_7457);
xor U11206 (N_11206,N_9241,N_5675);
and U11207 (N_11207,N_9983,N_8072);
or U11208 (N_11208,N_6740,N_6088);
and U11209 (N_11209,N_6422,N_8732);
xor U11210 (N_11210,N_5863,N_6016);
nand U11211 (N_11211,N_5826,N_5575);
nor U11212 (N_11212,N_5810,N_6035);
and U11213 (N_11213,N_7702,N_6374);
and U11214 (N_11214,N_9763,N_7140);
nand U11215 (N_11215,N_7546,N_7884);
or U11216 (N_11216,N_9129,N_7006);
nand U11217 (N_11217,N_6417,N_7195);
or U11218 (N_11218,N_9657,N_9228);
or U11219 (N_11219,N_9839,N_5984);
nor U11220 (N_11220,N_7985,N_9399);
xnor U11221 (N_11221,N_7123,N_9390);
or U11222 (N_11222,N_5989,N_6787);
nor U11223 (N_11223,N_8542,N_6860);
and U11224 (N_11224,N_9562,N_5443);
nand U11225 (N_11225,N_7040,N_7707);
nor U11226 (N_11226,N_5718,N_5032);
or U11227 (N_11227,N_5102,N_8935);
and U11228 (N_11228,N_5782,N_8024);
xor U11229 (N_11229,N_6698,N_9440);
and U11230 (N_11230,N_9501,N_7092);
and U11231 (N_11231,N_6024,N_6998);
or U11232 (N_11232,N_6412,N_7820);
and U11233 (N_11233,N_6236,N_5270);
or U11234 (N_11234,N_6673,N_7825);
and U11235 (N_11235,N_6922,N_8607);
and U11236 (N_11236,N_5014,N_8942);
nor U11237 (N_11237,N_7856,N_7900);
or U11238 (N_11238,N_6146,N_9769);
and U11239 (N_11239,N_8954,N_8698);
nand U11240 (N_11240,N_9982,N_5947);
nand U11241 (N_11241,N_7664,N_5862);
xor U11242 (N_11242,N_6327,N_8662);
or U11243 (N_11243,N_7838,N_5923);
nor U11244 (N_11244,N_9747,N_8485);
nand U11245 (N_11245,N_5336,N_5534);
xnor U11246 (N_11246,N_7767,N_9238);
and U11247 (N_11247,N_5531,N_7686);
or U11248 (N_11248,N_9132,N_5411);
and U11249 (N_11249,N_9496,N_9695);
or U11250 (N_11250,N_9016,N_9350);
and U11251 (N_11251,N_7347,N_7437);
or U11252 (N_11252,N_9171,N_6057);
and U11253 (N_11253,N_7484,N_8384);
nor U11254 (N_11254,N_5383,N_7324);
nand U11255 (N_11255,N_5168,N_7834);
and U11256 (N_11256,N_6878,N_8597);
nor U11257 (N_11257,N_9428,N_9844);
nor U11258 (N_11258,N_5886,N_5982);
xor U11259 (N_11259,N_7381,N_9978);
and U11260 (N_11260,N_7746,N_7055);
nor U11261 (N_11261,N_6395,N_9130);
nor U11262 (N_11262,N_5299,N_9646);
and U11263 (N_11263,N_9209,N_7968);
nor U11264 (N_11264,N_5763,N_5662);
and U11265 (N_11265,N_5274,N_9195);
or U11266 (N_11266,N_6467,N_8866);
nor U11267 (N_11267,N_7142,N_9482);
and U11268 (N_11268,N_9838,N_6905);
nor U11269 (N_11269,N_8598,N_6355);
or U11270 (N_11270,N_9153,N_6885);
or U11271 (N_11271,N_6884,N_9635);
nand U11272 (N_11272,N_7428,N_8182);
xnor U11273 (N_11273,N_8787,N_5003);
nor U11274 (N_11274,N_8020,N_7814);
or U11275 (N_11275,N_7344,N_5194);
nor U11276 (N_11276,N_9416,N_7886);
nand U11277 (N_11277,N_7881,N_9531);
or U11278 (N_11278,N_5203,N_6556);
and U11279 (N_11279,N_9520,N_9215);
nor U11280 (N_11280,N_9809,N_7573);
or U11281 (N_11281,N_9648,N_6442);
xnor U11282 (N_11282,N_6216,N_6100);
and U11283 (N_11283,N_7163,N_9064);
or U11284 (N_11284,N_8431,N_8242);
nand U11285 (N_11285,N_6683,N_8797);
or U11286 (N_11286,N_6694,N_9290);
xor U11287 (N_11287,N_6080,N_5803);
xnor U11288 (N_11288,N_5874,N_7174);
nand U11289 (N_11289,N_7217,N_6971);
or U11290 (N_11290,N_7116,N_7000);
xnor U11291 (N_11291,N_9043,N_5566);
or U11292 (N_11292,N_9285,N_5402);
nand U11293 (N_11293,N_7799,N_8706);
xnor U11294 (N_11294,N_7524,N_7249);
and U11295 (N_11295,N_9935,N_7335);
nand U11296 (N_11296,N_5643,N_5793);
nand U11297 (N_11297,N_9299,N_6332);
or U11298 (N_11298,N_9924,N_9923);
nor U11299 (N_11299,N_5869,N_5217);
nand U11300 (N_11300,N_5910,N_6127);
and U11301 (N_11301,N_8313,N_6215);
or U11302 (N_11302,N_8074,N_9522);
xnor U11303 (N_11303,N_5180,N_9240);
nor U11304 (N_11304,N_5727,N_5983);
or U11305 (N_11305,N_9892,N_8093);
nor U11306 (N_11306,N_9663,N_6750);
nand U11307 (N_11307,N_8670,N_8153);
and U11308 (N_11308,N_5085,N_7539);
nand U11309 (N_11309,N_6850,N_7469);
and U11310 (N_11310,N_8779,N_7565);
or U11311 (N_11311,N_5064,N_8213);
or U11312 (N_11312,N_7676,N_9944);
and U11313 (N_11313,N_8761,N_7693);
nand U11314 (N_11314,N_7962,N_5702);
nand U11315 (N_11315,N_8254,N_5152);
xor U11316 (N_11316,N_9664,N_6060);
nor U11317 (N_11317,N_8499,N_7209);
xor U11318 (N_11318,N_9128,N_5694);
and U11319 (N_11319,N_9918,N_9895);
nor U11320 (N_11320,N_8028,N_8215);
nand U11321 (N_11321,N_7202,N_8532);
and U11322 (N_11322,N_6629,N_8075);
xnor U11323 (N_11323,N_5011,N_9573);
xnor U11324 (N_11324,N_9782,N_5980);
nand U11325 (N_11325,N_7352,N_5946);
and U11326 (N_11326,N_9388,N_7561);
nor U11327 (N_11327,N_6651,N_6084);
and U11328 (N_11328,N_8048,N_9878);
or U11329 (N_11329,N_7922,N_5261);
nor U11330 (N_11330,N_9081,N_7806);
or U11331 (N_11331,N_9040,N_6988);
nand U11332 (N_11332,N_6735,N_5487);
nor U11333 (N_11333,N_9730,N_5346);
and U11334 (N_11334,N_5873,N_7247);
or U11335 (N_11335,N_8552,N_5115);
nand U11336 (N_11336,N_6508,N_6302);
nand U11337 (N_11337,N_9086,N_7656);
xor U11338 (N_11338,N_9793,N_7158);
nor U11339 (N_11339,N_7296,N_8902);
and U11340 (N_11340,N_7192,N_7319);
xnor U11341 (N_11341,N_9219,N_9277);
and U11342 (N_11342,N_6153,N_6461);
and U11343 (N_11343,N_6455,N_7281);
nor U11344 (N_11344,N_7760,N_5105);
nand U11345 (N_11345,N_5308,N_5425);
or U11346 (N_11346,N_5883,N_6040);
and U11347 (N_11347,N_9261,N_7833);
xnor U11348 (N_11348,N_5222,N_8086);
xnor U11349 (N_11349,N_9938,N_6636);
and U11350 (N_11350,N_9379,N_7650);
nor U11351 (N_11351,N_5256,N_7869);
or U11352 (N_11352,N_5537,N_6483);
and U11353 (N_11353,N_8370,N_5312);
or U11354 (N_11354,N_9281,N_5960);
nand U11355 (N_11355,N_7492,N_6621);
and U11356 (N_11356,N_5159,N_8410);
nand U11357 (N_11357,N_7389,N_6211);
nor U11358 (N_11358,N_7112,N_6404);
nor U11359 (N_11359,N_8896,N_8374);
nand U11360 (N_11360,N_6010,N_5812);
nand U11361 (N_11361,N_5552,N_8904);
or U11362 (N_11362,N_7414,N_8925);
nor U11363 (N_11363,N_5491,N_5380);
xor U11364 (N_11364,N_8096,N_9491);
or U11365 (N_11365,N_7392,N_7552);
or U11366 (N_11366,N_8677,N_6453);
nor U11367 (N_11367,N_8486,N_7107);
or U11368 (N_11368,N_9693,N_9610);
and U11369 (N_11369,N_7840,N_8817);
or U11370 (N_11370,N_8578,N_6253);
and U11371 (N_11371,N_8694,N_6729);
or U11372 (N_11372,N_7537,N_5272);
or U11373 (N_11373,N_6886,N_7848);
and U11374 (N_11374,N_9600,N_6318);
or U11375 (N_11375,N_7916,N_6866);
nand U11376 (N_11376,N_8155,N_8339);
xor U11377 (N_11377,N_5809,N_9074);
and U11378 (N_11378,N_7119,N_9806);
nand U11379 (N_11379,N_8280,N_8553);
xnor U11380 (N_11380,N_9764,N_8409);
nand U11381 (N_11381,N_5940,N_8644);
xor U11382 (N_11382,N_7369,N_8010);
xnor U11383 (N_11383,N_6094,N_8224);
nand U11384 (N_11384,N_8763,N_6076);
or U11385 (N_11385,N_5359,N_5680);
xnor U11386 (N_11386,N_6179,N_6548);
and U11387 (N_11387,N_5056,N_7409);
nor U11388 (N_11388,N_7300,N_5205);
nor U11389 (N_11389,N_6771,N_6908);
nand U11390 (N_11390,N_5488,N_5590);
and U11391 (N_11391,N_8574,N_8908);
nor U11392 (N_11392,N_9236,N_8796);
and U11393 (N_11393,N_5685,N_7425);
nand U11394 (N_11394,N_7775,N_9868);
nor U11395 (N_11395,N_9953,N_8091);
and U11396 (N_11396,N_9147,N_5393);
and U11397 (N_11397,N_5029,N_9257);
or U11398 (N_11398,N_6936,N_9616);
nor U11399 (N_11399,N_6331,N_8768);
xnor U11400 (N_11400,N_6068,N_9036);
nor U11401 (N_11401,N_8022,N_8980);
nand U11402 (N_11402,N_7700,N_5903);
or U11403 (N_11403,N_8709,N_9796);
nor U11404 (N_11404,N_6761,N_5008);
or U11405 (N_11405,N_9451,N_7722);
and U11406 (N_11406,N_9872,N_5904);
nor U11407 (N_11407,N_6182,N_6458);
nand U11408 (N_11408,N_7773,N_8186);
or U11409 (N_11409,N_9550,N_8956);
nand U11410 (N_11410,N_8859,N_5784);
or U11411 (N_11411,N_5845,N_9480);
or U11412 (N_11412,N_8812,N_5396);
nor U11413 (N_11413,N_8628,N_9557);
nand U11414 (N_11414,N_7100,N_8951);
xor U11415 (N_11415,N_9489,N_8688);
xor U11416 (N_11416,N_6313,N_8151);
and U11417 (N_11417,N_5007,N_5701);
and U11418 (N_11418,N_7543,N_6661);
nand U11419 (N_11419,N_6446,N_5239);
and U11420 (N_11420,N_9125,N_9670);
or U11421 (N_11421,N_6800,N_5327);
xnor U11422 (N_11422,N_6186,N_9523);
nor U11423 (N_11423,N_9472,N_5045);
nor U11424 (N_11424,N_9288,N_8580);
and U11425 (N_11425,N_6736,N_9212);
nor U11426 (N_11426,N_6003,N_8690);
or U11427 (N_11427,N_7498,N_5699);
xor U11428 (N_11428,N_8230,N_8227);
nand U11429 (N_11429,N_9915,N_7184);
and U11430 (N_11430,N_6218,N_6680);
xnor U11431 (N_11431,N_8573,N_6188);
nand U11432 (N_11432,N_9417,N_9510);
nor U11433 (N_11433,N_9558,N_5743);
or U11434 (N_11434,N_6012,N_6013);
xor U11435 (N_11435,N_9538,N_7888);
xnor U11436 (N_11436,N_6375,N_8249);
nor U11437 (N_11437,N_7540,N_7969);
xnor U11438 (N_11438,N_7175,N_8198);
xnor U11439 (N_11439,N_9395,N_9421);
and U11440 (N_11440,N_7954,N_9377);
or U11441 (N_11441,N_5255,N_7621);
or U11442 (N_11442,N_5128,N_5432);
xnor U11443 (N_11443,N_5506,N_5114);
nor U11444 (N_11444,N_8909,N_6789);
or U11445 (N_11445,N_8710,N_6276);
xor U11446 (N_11446,N_9183,N_5020);
nor U11447 (N_11447,N_7677,N_8132);
nor U11448 (N_11448,N_7223,N_6347);
nand U11449 (N_11449,N_5595,N_8820);
xnor U11450 (N_11450,N_5438,N_7490);
xor U11451 (N_11451,N_5027,N_8642);
or U11452 (N_11452,N_9572,N_7885);
and U11453 (N_11453,N_5192,N_5732);
nor U11454 (N_11454,N_5370,N_8609);
nand U11455 (N_11455,N_6476,N_6205);
nand U11456 (N_11456,N_5483,N_8451);
and U11457 (N_11457,N_7605,N_9689);
xor U11458 (N_11458,N_6914,N_9325);
and U11459 (N_11459,N_6325,N_8960);
and U11460 (N_11460,N_6303,N_9959);
nor U11461 (N_11461,N_9449,N_8672);
or U11462 (N_11462,N_9916,N_6923);
xnor U11463 (N_11463,N_6562,N_5435);
nor U11464 (N_11464,N_5814,N_5540);
xnor U11465 (N_11465,N_5384,N_8330);
or U11466 (N_11466,N_5212,N_5421);
nand U11467 (N_11467,N_6584,N_8536);
or U11468 (N_11468,N_8523,N_6882);
xor U11469 (N_11469,N_6957,N_7416);
nor U11470 (N_11470,N_8658,N_5600);
and U11471 (N_11471,N_8558,N_7028);
and U11472 (N_11472,N_9756,N_8471);
xor U11473 (N_11473,N_5747,N_5892);
and U11474 (N_11474,N_5729,N_9711);
nor U11475 (N_11475,N_6687,N_6756);
nor U11476 (N_11476,N_6893,N_9357);
xnor U11477 (N_11477,N_6349,N_9901);
or U11478 (N_11478,N_8207,N_6170);
xnor U11479 (N_11479,N_9252,N_6363);
xnor U11480 (N_11480,N_8266,N_6396);
nor U11481 (N_11481,N_9239,N_7067);
or U11482 (N_11482,N_6570,N_6826);
nor U11483 (N_11483,N_7453,N_7638);
xnor U11484 (N_11484,N_6212,N_8150);
nor U11485 (N_11485,N_7177,N_9306);
or U11486 (N_11486,N_8457,N_5050);
and U11487 (N_11487,N_7966,N_7126);
nand U11488 (N_11488,N_9926,N_6492);
and U11489 (N_11489,N_7086,N_9672);
or U11490 (N_11490,N_7870,N_7038);
nand U11491 (N_11491,N_7027,N_5541);
nand U11492 (N_11492,N_8841,N_8054);
nor U11493 (N_11493,N_6144,N_9912);
xor U11494 (N_11494,N_7516,N_5028);
xnor U11495 (N_11495,N_9134,N_6768);
nand U11496 (N_11496,N_6586,N_7149);
nand U11497 (N_11497,N_6271,N_9803);
or U11498 (N_11498,N_9721,N_6152);
nor U11499 (N_11499,N_9358,N_7611);
nor U11500 (N_11500,N_7321,N_5952);
nand U11501 (N_11501,N_5145,N_7898);
nand U11502 (N_11502,N_8400,N_8002);
nor U11503 (N_11503,N_5139,N_6784);
nor U11504 (N_11504,N_6704,N_9679);
nor U11505 (N_11505,N_8247,N_8811);
nor U11506 (N_11506,N_6149,N_6861);
and U11507 (N_11507,N_7554,N_6603);
xor U11508 (N_11508,N_6433,N_5172);
and U11509 (N_11509,N_6426,N_7231);
nand U11510 (N_11510,N_6403,N_7064);
xor U11511 (N_11511,N_8047,N_7434);
xnor U11512 (N_11512,N_8103,N_6356);
and U11513 (N_11513,N_7951,N_9052);
or U11514 (N_11514,N_9837,N_9832);
xor U11515 (N_11515,N_8860,N_7030);
nand U11516 (N_11516,N_5026,N_8461);
xnor U11517 (N_11517,N_7128,N_5132);
and U11518 (N_11518,N_5914,N_6739);
nand U11519 (N_11519,N_9996,N_9201);
or U11520 (N_11520,N_6187,N_6256);
nand U11521 (N_11521,N_7234,N_7824);
nor U11522 (N_11522,N_9876,N_6523);
or U11523 (N_11523,N_8565,N_9051);
or U11524 (N_11524,N_6643,N_5320);
and U11525 (N_11525,N_6830,N_8663);
or U11526 (N_11526,N_5446,N_6243);
nand U11527 (N_11527,N_5496,N_7911);
nand U11528 (N_11528,N_6572,N_5944);
and U11529 (N_11529,N_6260,N_6671);
xnor U11530 (N_11530,N_8317,N_7155);
and U11531 (N_11531,N_5568,N_8964);
xor U11532 (N_11532,N_5829,N_5301);
or U11533 (N_11533,N_9682,N_7350);
nand U11534 (N_11534,N_7685,N_6941);
xnor U11535 (N_11535,N_5948,N_9854);
or U11536 (N_11536,N_6424,N_7226);
nand U11537 (N_11537,N_8199,N_9311);
nand U11538 (N_11538,N_8739,N_8386);
and U11539 (N_11539,N_8507,N_7566);
nor U11540 (N_11540,N_9788,N_9828);
or U11541 (N_11541,N_6956,N_8655);
nor U11542 (N_11542,N_8525,N_7506);
nor U11543 (N_11543,N_9084,N_7261);
xor U11544 (N_11544,N_8300,N_9279);
and U11545 (N_11545,N_7001,N_9315);
and U11546 (N_11546,N_9776,N_7265);
nor U11547 (N_11547,N_5457,N_5652);
nor U11548 (N_11548,N_5431,N_6835);
nand U11549 (N_11549,N_7240,N_6960);
nand U11550 (N_11550,N_7837,N_8143);
or U11551 (N_11551,N_8333,N_9433);
nor U11552 (N_11552,N_8327,N_6124);
xor U11553 (N_11553,N_6640,N_7768);
or U11554 (N_11554,N_9282,N_7946);
nand U11555 (N_11555,N_6108,N_5498);
nor U11556 (N_11556,N_9778,N_7924);
nor U11557 (N_11557,N_5503,N_7393);
xnor U11558 (N_11558,N_5182,N_6743);
nand U11559 (N_11559,N_7323,N_8062);
and U11560 (N_11560,N_9298,N_8007);
nand U11561 (N_11561,N_5076,N_8210);
or U11562 (N_11562,N_9220,N_9442);
nor U11563 (N_11563,N_8362,N_7633);
nand U11564 (N_11564,N_9810,N_5968);
nand U11565 (N_11565,N_8819,N_7374);
nand U11566 (N_11566,N_7629,N_9690);
and U11567 (N_11567,N_5037,N_7597);
nand U11568 (N_11568,N_5227,N_5267);
or U11569 (N_11569,N_5310,N_8038);
nand U11570 (N_11570,N_5424,N_9941);
and U11571 (N_11571,N_5471,N_6785);
nand U11572 (N_11572,N_5303,N_5527);
and U11573 (N_11573,N_9622,N_7975);
or U11574 (N_11574,N_6288,N_6474);
xor U11575 (N_11575,N_8687,N_6169);
nand U11576 (N_11576,N_5419,N_7167);
nor U11577 (N_11577,N_8118,N_9681);
and U11578 (N_11578,N_7845,N_7733);
xnor U11579 (N_11579,N_9418,N_8177);
nor U11580 (N_11580,N_7853,N_6565);
and U11581 (N_11581,N_5963,N_8084);
nor U11582 (N_11582,N_8501,N_5884);
nor U11583 (N_11583,N_9687,N_8165);
nor U11584 (N_11584,N_6872,N_9841);
nand U11585 (N_11585,N_5895,N_7783);
nand U11586 (N_11586,N_6067,N_7550);
nor U11587 (N_11587,N_8192,N_8581);
nand U11588 (N_11588,N_5919,N_6222);
xnor U11589 (N_11589,N_7058,N_9500);
and U11590 (N_11590,N_6306,N_8138);
nor U11591 (N_11591,N_7880,N_7789);
nand U11592 (N_11592,N_6889,N_8705);
xor U11593 (N_11593,N_9655,N_6616);
nand U11594 (N_11594,N_6935,N_7613);
nor U11595 (N_11595,N_7458,N_5522);
xnor U11596 (N_11596,N_5572,N_6943);
nand U11597 (N_11597,N_9319,N_6950);
or U11598 (N_11598,N_6092,N_6503);
and U11599 (N_11599,N_6983,N_8920);
nor U11600 (N_11600,N_5282,N_5043);
nor U11601 (N_11601,N_8858,N_8435);
nor U11602 (N_11602,N_9564,N_7862);
nand U11603 (N_11603,N_7127,N_6737);
and U11604 (N_11604,N_9293,N_8516);
nor U11605 (N_11605,N_7063,N_9950);
nor U11606 (N_11606,N_8689,N_6491);
or U11607 (N_11607,N_6239,N_7914);
or U11608 (N_11608,N_8921,N_6009);
xor U11609 (N_11609,N_8983,N_6633);
or U11610 (N_11610,N_5089,N_8695);
nand U11611 (N_11611,N_7741,N_9176);
or U11612 (N_11612,N_9524,N_9398);
nand U11613 (N_11613,N_5240,N_6340);
xnor U11614 (N_11614,N_7176,N_8236);
xor U11615 (N_11615,N_5202,N_8077);
xnor U11616 (N_11616,N_7061,N_5200);
and U11617 (N_11617,N_5131,N_9767);
nand U11618 (N_11618,N_5669,N_7723);
nor U11619 (N_11619,N_7056,N_7406);
and U11620 (N_11620,N_6525,N_5858);
xor U11621 (N_11621,N_9873,N_7619);
or U11622 (N_11622,N_7271,N_8070);
and U11623 (N_11623,N_8201,N_9166);
or U11624 (N_11624,N_9099,N_6104);
nand U11625 (N_11625,N_9742,N_7452);
and U11626 (N_11626,N_8731,N_6622);
nand U11627 (N_11627,N_8785,N_7720);
nand U11628 (N_11628,N_7868,N_7031);
xor U11629 (N_11629,N_5529,N_5399);
nor U11630 (N_11630,N_7290,N_7726);
xnor U11631 (N_11631,N_6266,N_6846);
nand U11632 (N_11632,N_9363,N_7590);
nor U11633 (N_11633,N_7689,N_8372);
xnor U11634 (N_11634,N_9479,N_8092);
and U11635 (N_11635,N_9007,N_9475);
xor U11636 (N_11636,N_7823,N_7390);
or U11637 (N_11637,N_8142,N_8966);
nand U11638 (N_11638,N_9352,N_8852);
xnor U11639 (N_11639,N_9882,N_7351);
xor U11640 (N_11640,N_7179,N_9162);
nand U11641 (N_11641,N_9234,N_6976);
nand U11642 (N_11642,N_8949,N_9244);
nand U11643 (N_11643,N_5632,N_8704);
and U11644 (N_11644,N_8566,N_9652);
or U11645 (N_11645,N_7528,N_7310);
and U11646 (N_11646,N_9640,N_7012);
nor U11647 (N_11647,N_7772,N_7691);
or U11648 (N_11648,N_8877,N_8359);
xor U11649 (N_11649,N_7476,N_7384);
xnor U11650 (N_11650,N_5746,N_6062);
nor U11651 (N_11651,N_5504,N_9461);
nor U11652 (N_11652,N_6788,N_7696);
xor U11653 (N_11653,N_8114,N_9088);
xor U11654 (N_11654,N_5932,N_9443);
and U11655 (N_11655,N_7227,N_7576);
and U11656 (N_11656,N_6485,N_7731);
and U11657 (N_11657,N_5618,N_8459);
or U11658 (N_11658,N_7053,N_6097);
nor U11659 (N_11659,N_8345,N_5335);
or U11660 (N_11660,N_9553,N_7730);
nand U11661 (N_11661,N_8606,N_5010);
nand U11662 (N_11662,N_7955,N_8196);
xor U11663 (N_11663,N_7852,N_7266);
or U11664 (N_11664,N_9210,N_7472);
and U11665 (N_11665,N_7162,N_5530);
nor U11666 (N_11666,N_5472,N_7087);
and U11667 (N_11667,N_6530,N_5956);
nor U11668 (N_11668,N_6231,N_5767);
or U11669 (N_11669,N_7628,N_6979);
or U11670 (N_11670,N_9908,N_8423);
xnor U11671 (N_11671,N_9863,N_9095);
or U11672 (N_11672,N_6857,N_9172);
nor U11673 (N_11673,N_6722,N_8309);
or U11674 (N_11674,N_7594,N_9597);
xnor U11675 (N_11675,N_7500,N_5766);
nor U11676 (N_11676,N_8175,N_9948);
and U11677 (N_11677,N_8035,N_9563);
nor U11678 (N_11678,N_7441,N_6996);
nor U11679 (N_11679,N_9002,N_9556);
nor U11680 (N_11680,N_5547,N_6364);
nand U11681 (N_11681,N_9367,N_8320);
nand U11682 (N_11682,N_8952,N_7831);
or U11683 (N_11683,N_5453,N_7714);
or U11684 (N_11684,N_9540,N_8231);
or U11685 (N_11685,N_5524,N_5773);
xor U11686 (N_11686,N_7999,N_8060);
nor U11687 (N_11687,N_7842,N_7052);
or U11688 (N_11688,N_7802,N_5536);
nand U11689 (N_11689,N_5772,N_9300);
xnor U11690 (N_11690,N_5953,N_6174);
xor U11691 (N_11691,N_5049,N_8193);
nand U11692 (N_11692,N_6209,N_8223);
or U11693 (N_11693,N_9382,N_8197);
nor U11694 (N_11694,N_9169,N_9078);
and U11695 (N_11695,N_8364,N_6527);
xnor U11696 (N_11696,N_6154,N_8169);
xor U11697 (N_11697,N_6968,N_8917);
nor U11698 (N_11698,N_5035,N_5209);
xor U11699 (N_11699,N_8783,N_5284);
and U11700 (N_11700,N_7663,N_7934);
and U11701 (N_11701,N_5757,N_5258);
or U11702 (N_11702,N_5612,N_6321);
xor U11703 (N_11703,N_8549,N_7213);
nand U11704 (N_11704,N_7360,N_8163);
nor U11705 (N_11705,N_8916,N_5325);
or U11706 (N_11706,N_9773,N_5478);
or U11707 (N_11707,N_6580,N_9283);
nor U11708 (N_11708,N_9251,N_8164);
nand U11709 (N_11709,N_5958,N_8799);
nand U11710 (N_11710,N_9825,N_6566);
and U11711 (N_11711,N_9144,N_7583);
nor U11712 (N_11712,N_6577,N_5226);
and U11713 (N_11713,N_7085,N_7655);
xor U11714 (N_11714,N_8595,N_7781);
and U11715 (N_11715,N_9612,N_9308);
nand U11716 (N_11716,N_7404,N_8180);
and U11717 (N_11717,N_7877,N_7941);
nand U11718 (N_11718,N_7609,N_8323);
and U11719 (N_11719,N_7670,N_5664);
nor U11720 (N_11720,N_7008,N_9227);
and U11721 (N_11721,N_9917,N_9465);
or U11722 (N_11722,N_5237,N_9110);
xor U11723 (N_11723,N_6343,N_7304);
nor U11724 (N_11724,N_8592,N_7715);
nor U11725 (N_11725,N_6841,N_8488);
nand U11726 (N_11726,N_7925,N_9628);
and U11727 (N_11727,N_7331,N_8842);
or U11728 (N_11728,N_8627,N_9343);
or U11729 (N_11729,N_9301,N_9530);
xor U11730 (N_11730,N_6693,N_6066);
or U11731 (N_11731,N_5001,N_7160);
and U11732 (N_11732,N_7927,N_6177);
nor U11733 (N_11733,N_7139,N_8973);
nor U11734 (N_11734,N_7711,N_8645);
or U11735 (N_11735,N_6667,N_7243);
xnor U11736 (N_11736,N_5291,N_8414);
or U11737 (N_11737,N_6953,N_7973);
or U11738 (N_11738,N_6921,N_7919);
nor U11739 (N_11739,N_8757,N_7604);
xor U11740 (N_11740,N_5070,N_5831);
xnor U11741 (N_11741,N_6052,N_5208);
xnor U11742 (N_11742,N_8503,N_7294);
nor U11743 (N_11743,N_7062,N_6091);
nand U11744 (N_11744,N_5843,N_6532);
xnor U11745 (N_11745,N_7420,N_8795);
nor U11746 (N_11746,N_8472,N_7531);
nor U11747 (N_11747,N_9725,N_7871);
nor U11748 (N_11748,N_7256,N_6738);
xor U11749 (N_11749,N_9964,N_9852);
nor U11750 (N_11750,N_8735,N_6438);
and U11751 (N_11751,N_9434,N_5144);
or U11752 (N_11752,N_6701,N_8667);
xnor U11753 (N_11753,N_6470,N_7391);
nand U11754 (N_11754,N_8632,N_9208);
and U11755 (N_11755,N_8801,N_8747);
and U11756 (N_11756,N_8494,N_9318);
or U11757 (N_11757,N_7316,N_9041);
or U11758 (N_11758,N_8861,N_7983);
nor U11759 (N_11759,N_6615,N_9093);
nand U11760 (N_11760,N_7263,N_6385);
xnor U11761 (N_11761,N_6913,N_7902);
and U11762 (N_11762,N_6710,N_8462);
xnor U11763 (N_11763,N_6180,N_9089);
nor U11764 (N_11764,N_6059,N_5545);
nor U11765 (N_11765,N_9700,N_5822);
nand U11766 (N_11766,N_5385,N_6595);
nor U11767 (N_11767,N_9415,N_6333);
xnor U11768 (N_11768,N_9728,N_9435);
or U11769 (N_11769,N_7666,N_5109);
nand U11770 (N_11770,N_7617,N_8794);
nand U11771 (N_11771,N_9303,N_5860);
and U11772 (N_11772,N_9561,N_6940);
nor U11773 (N_11773,N_5724,N_8776);
or U11774 (N_11774,N_8729,N_8893);
and U11775 (N_11775,N_9079,N_8789);
nand U11776 (N_11776,N_8265,N_7713);
nand U11777 (N_11777,N_8766,N_6646);
and U11778 (N_11778,N_9237,N_9914);
and U11779 (N_11779,N_8271,N_7075);
and U11780 (N_11780,N_5891,N_9459);
and U11781 (N_11781,N_6473,N_7483);
xor U11782 (N_11782,N_5538,N_7796);
xnor U11783 (N_11783,N_9855,N_6952);
nor U11784 (N_11784,N_8380,N_7274);
xor U11785 (N_11785,N_7394,N_6772);
nand U11786 (N_11786,N_9680,N_9065);
and U11787 (N_11787,N_7547,N_8393);
xor U11788 (N_11788,N_7387,N_7607);
or U11789 (N_11789,N_7088,N_8639);
and U11790 (N_11790,N_5799,N_9022);
nor U11791 (N_11791,N_8788,N_5550);
nand U11792 (N_11792,N_5243,N_7530);
nor U11793 (N_11793,N_9122,N_8341);
nor U11794 (N_11794,N_7807,N_9857);
or U11795 (N_11795,N_9590,N_8270);
nor U11796 (N_11796,N_9994,N_8299);
or U11797 (N_11797,N_6876,N_9880);
and U11798 (N_11798,N_8465,N_9431);
or U11799 (N_11799,N_7659,N_5926);
xor U11800 (N_11800,N_7433,N_6542);
xnor U11801 (N_11801,N_6967,N_9957);
xor U11802 (N_11802,N_5178,N_6911);
nor U11803 (N_11803,N_6533,N_7250);
or U11804 (N_11804,N_6642,N_8502);
and U11805 (N_11805,N_7515,N_9619);
and U11806 (N_11806,N_7805,N_5779);
xor U11807 (N_11807,N_6692,N_9503);
nor U11808 (N_11808,N_6906,N_8483);
nand U11809 (N_11809,N_7336,N_9072);
xor U11810 (N_11810,N_9207,N_9701);
xnor U11811 (N_11811,N_9677,N_5837);
or U11812 (N_11812,N_6834,N_5768);
and U11813 (N_11813,N_6290,N_6824);
xor U11814 (N_11814,N_6324,N_9709);
nand U11815 (N_11815,N_7286,N_6449);
xnor U11816 (N_11816,N_7912,N_7230);
nand U11817 (N_11817,N_6072,N_5661);
nand U11818 (N_11818,N_8593,N_8130);
and U11819 (N_11819,N_6973,N_5977);
xor U11820 (N_11820,N_6036,N_8430);
or U11821 (N_11821,N_5080,N_7758);
xor U11822 (N_11822,N_8798,N_6708);
or U11823 (N_11823,N_9090,N_8099);
or U11824 (N_11824,N_5123,N_6954);
nor U11825 (N_11825,N_7228,N_9596);
and U11826 (N_11826,N_5593,N_6235);
nor U11827 (N_11827,N_9893,N_6285);
xor U11828 (N_11828,N_5057,N_9329);
xor U11829 (N_11829,N_9187,N_6030);
xnor U11830 (N_11830,N_6283,N_7936);
nand U11831 (N_11831,N_6265,N_8784);
and U11832 (N_11832,N_9821,N_5429);
or U11833 (N_11833,N_9903,N_8491);
xor U11834 (N_11834,N_9011,N_8743);
xor U11835 (N_11835,N_7101,N_6172);
nor U11836 (N_11836,N_5510,N_7353);
or U11837 (N_11837,N_7757,N_7505);
xnor U11838 (N_11838,N_9104,N_5591);
xnor U11839 (N_11839,N_6367,N_7557);
nand U11840 (N_11840,N_7200,N_6263);
nand U11841 (N_11841,N_6443,N_7703);
or U11842 (N_11842,N_6767,N_5785);
xnor U11843 (N_11843,N_6410,N_7788);
or U11844 (N_11844,N_8496,N_9217);
or U11845 (N_11845,N_6370,N_5644);
or U11846 (N_11846,N_6406,N_5777);
and U11847 (N_11847,N_9106,N_7487);
and U11848 (N_11848,N_7131,N_5324);
or U11849 (N_11849,N_8831,N_9727);
nand U11850 (N_11850,N_8023,N_6219);
nor U11851 (N_11851,N_5971,N_7997);
or U11852 (N_11852,N_7199,N_5617);
nand U11853 (N_11853,N_7587,N_8061);
and U11854 (N_11854,N_8997,N_9295);
and U11855 (N_11855,N_5696,N_6268);
or U11856 (N_11856,N_9659,N_9543);
xnor U11857 (N_11857,N_8840,N_6397);
nor U11858 (N_11858,N_5042,N_7625);
nor U11859 (N_11859,N_9386,N_5693);
or U11860 (N_11860,N_8863,N_6609);
and U11861 (N_11861,N_7815,N_7906);
xnor U11862 (N_11862,N_8139,N_7753);
or U11863 (N_11863,N_5363,N_7738);
or U11864 (N_11864,N_9297,N_7366);
or U11865 (N_11865,N_9567,N_9902);
nand U11866 (N_11866,N_9904,N_8996);
nand U11867 (N_11867,N_5317,N_5733);
xor U11868 (N_11868,N_7130,N_6786);
nor U11869 (N_11869,N_5423,N_8847);
and U11870 (N_11870,N_7166,N_8984);
and U11871 (N_11871,N_9802,N_9149);
xnor U11872 (N_11872,N_9942,N_5668);
and U11873 (N_11873,N_5352,N_7461);
and U11874 (N_11874,N_8660,N_7402);
nand U11875 (N_11875,N_8015,N_5353);
and U11876 (N_11876,N_6046,N_6958);
nor U11877 (N_11877,N_9124,N_8006);
nand U11878 (N_11878,N_9211,N_9067);
or U11879 (N_11879,N_5140,N_6605);
nand U11880 (N_11880,N_6909,N_9585);
xnor U11881 (N_11881,N_9864,N_8476);
nor U11882 (N_11882,N_9305,N_5608);
nor U11883 (N_11883,N_9594,N_9898);
or U11884 (N_11884,N_9627,N_7026);
or U11885 (N_11885,N_9660,N_9430);
xor U11886 (N_11886,N_8804,N_5228);
nor U11887 (N_11887,N_8241,N_6070);
nand U11888 (N_11888,N_6670,N_7378);
or U11889 (N_11889,N_7626,N_9850);
or U11890 (N_11890,N_8756,N_5878);
nor U11891 (N_11891,N_9247,N_5489);
nand U11892 (N_11892,N_5067,N_8222);
or U11893 (N_11893,N_7699,N_7606);
nor U11894 (N_11894,N_9606,N_9779);
and U11895 (N_11895,N_9886,N_5592);
nor U11896 (N_11896,N_7832,N_8845);
xnor U11897 (N_11897,N_9194,N_9485);
xnor U11898 (N_11898,N_5005,N_5351);
nand U11899 (N_11899,N_9789,N_6115);
and U11900 (N_11900,N_7671,N_5791);
or U11901 (N_11901,N_9155,N_7439);
xor U11902 (N_11902,N_6106,N_8853);
and U11903 (N_11903,N_7792,N_9047);
nand U11904 (N_11904,N_7859,N_8019);
xnor U11905 (N_11905,N_5082,N_7536);
nand U11906 (N_11906,N_7204,N_6006);
xor U11907 (N_11907,N_9715,N_6762);
nand U11908 (N_11908,N_9929,N_6197);
nor U11909 (N_11909,N_9031,N_6758);
nand U11910 (N_11910,N_7961,N_8661);
and U11911 (N_11911,N_5244,N_6653);
nand U11912 (N_11912,N_8482,N_7509);
xnor U11913 (N_11913,N_5844,N_6002);
xnor U11914 (N_11914,N_8322,N_7701);
xnor U11915 (N_11915,N_6232,N_7445);
nor U11916 (N_11916,N_7471,N_9623);
or U11917 (N_11917,N_5847,N_6623);
nor U11918 (N_11918,N_8697,N_5481);
or U11919 (N_11919,N_5533,N_6712);
or U11920 (N_11920,N_7136,N_5876);
xor U11921 (N_11921,N_6828,N_9554);
xor U11922 (N_11922,N_7623,N_7267);
xnor U11923 (N_11923,N_6466,N_9932);
and U11924 (N_11924,N_6481,N_9542);
nand U11925 (N_11925,N_6244,N_5373);
and U11926 (N_11926,N_5642,N_5039);
and U11927 (N_11927,N_7883,N_6413);
or U11928 (N_11928,N_7910,N_7334);
nor U11929 (N_11929,N_6817,N_5885);
and U11930 (N_11930,N_5480,N_6571);
nor U11931 (N_11931,N_6776,N_6307);
and U11932 (N_11932,N_5897,N_5857);
nand U11933 (N_11933,N_5273,N_5962);
nor U11934 (N_11934,N_9505,N_9340);
or U11935 (N_11935,N_5464,N_8582);
or U11936 (N_11936,N_7349,N_9008);
or U11937 (N_11937,N_6801,N_5902);
xnor U11938 (N_11938,N_8383,N_6373);
or U11939 (N_11939,N_5505,N_8851);
and U11940 (N_11940,N_9947,N_8095);
nor U11941 (N_11941,N_6662,N_5051);
nand U11942 (N_11942,N_9717,N_7896);
and U11943 (N_11943,N_5905,N_8721);
xor U11944 (N_11944,N_5990,N_8682);
or U11945 (N_11945,N_9158,N_7337);
and U11946 (N_11946,N_5780,N_6972);
xor U11947 (N_11947,N_8764,N_8398);
xnor U11948 (N_11948,N_7400,N_9048);
nand U11949 (N_11949,N_9575,N_9397);
nor U11950 (N_11950,N_5305,N_6171);
and U11951 (N_11951,N_6628,N_8419);
nand U11952 (N_11952,N_7073,N_9922);
xor U11953 (N_11953,N_7220,N_7873);
or U11954 (N_11954,N_7264,N_5260);
nor U11955 (N_11955,N_9962,N_8161);
nor U11956 (N_11956,N_5120,N_9173);
nor U11957 (N_11957,N_6731,N_6151);
nor U11958 (N_11958,N_9163,N_6732);
nand U11959 (N_11959,N_8298,N_7313);
or U11960 (N_11960,N_8559,N_9965);
xor U11961 (N_11961,N_8447,N_8666);
or U11962 (N_11962,N_7518,N_6745);
xor U11963 (N_11963,N_9958,N_8424);
nor U11964 (N_11964,N_6445,N_7876);
nor U11965 (N_11965,N_5778,N_8652);
and U11966 (N_11966,N_6125,N_6078);
and U11967 (N_11967,N_6206,N_7486);
nand U11968 (N_11968,N_5389,N_7218);
nor U11969 (N_11969,N_6192,N_9676);
nor U11970 (N_11970,N_8782,N_7688);
nand U11971 (N_11971,N_6353,N_6390);
xnor U11972 (N_11972,N_9845,N_9724);
nand U11973 (N_11973,N_9034,N_8105);
and U11974 (N_11974,N_7942,N_8358);
nand U11975 (N_11975,N_8067,N_9362);
xor U11976 (N_11976,N_8850,N_7282);
xor U11977 (N_11977,N_7897,N_5154);
xnor U11978 (N_11978,N_6018,N_7365);
nor U11979 (N_11979,N_5289,N_5427);
nor U11980 (N_11980,N_6920,N_7645);
and U11981 (N_11981,N_9706,N_9103);
or U11982 (N_11982,N_8504,N_8584);
nor U11983 (N_11983,N_9488,N_8568);
or U11984 (N_11984,N_6890,N_6827);
and U11985 (N_11985,N_9042,N_5300);
and U11986 (N_11986,N_6191,N_5759);
nand U11987 (N_11987,N_8405,N_7456);
or U11988 (N_11988,N_9050,N_7944);
or U11989 (N_11989,N_7071,N_5671);
xnor U11990 (N_11990,N_5907,N_8615);
xor U11991 (N_11991,N_6524,N_7191);
xor U11992 (N_11992,N_6782,N_6376);
xnor U11993 (N_11993,N_8547,N_6840);
or U11994 (N_11994,N_9049,N_9121);
and U11995 (N_11995,N_8991,N_8470);
or U11996 (N_11996,N_5500,N_6551);
nor U11997 (N_11997,N_5561,N_7328);
nand U11998 (N_11998,N_5913,N_7991);
and U11999 (N_11999,N_6202,N_6293);
or U12000 (N_12000,N_5626,N_7682);
xor U12001 (N_12001,N_5386,N_5248);
xnor U12002 (N_12002,N_9263,N_8126);
and U12003 (N_12003,N_7507,N_8406);
nor U12004 (N_12004,N_9017,N_6386);
xnor U12005 (N_12005,N_9956,N_5297);
xor U12006 (N_12006,N_7047,N_7684);
or U12007 (N_12007,N_7314,N_7965);
and U12008 (N_12008,N_7706,N_7777);
nand U12009 (N_12009,N_7039,N_8638);
nor U12010 (N_12010,N_6865,N_6600);
nand U12011 (N_12011,N_8610,N_6079);
nand U12012 (N_12012,N_8978,N_7005);
xnor U12013 (N_12013,N_8897,N_6114);
nor U12014 (N_12014,N_9009,N_5666);
nor U12015 (N_12015,N_8263,N_9911);
or U12016 (N_12016,N_7522,N_5855);
nand U12017 (N_12017,N_8767,N_9588);
or U12018 (N_12018,N_7037,N_6463);
xor U12019 (N_12019,N_7021,N_5331);
nand U12020 (N_12020,N_9274,N_9900);
or U12021 (N_12021,N_7118,N_9934);
xor U12022 (N_12022,N_8825,N_6337);
and U12023 (N_12023,N_6121,N_6305);
or U12024 (N_12024,N_8889,N_5149);
nand U12025 (N_12025,N_7326,N_7114);
and U12026 (N_12026,N_8900,N_7588);
nor U12027 (N_12027,N_5722,N_9462);
xor U12028 (N_12028,N_8892,N_5210);
xnor U12029 (N_12029,N_7510,N_6746);
xor U12030 (N_12030,N_6190,N_9191);
nor U12031 (N_12031,N_9495,N_6399);
nand U12032 (N_12032,N_5147,N_6852);
or U12033 (N_12033,N_9427,N_8875);
or U12034 (N_12034,N_7572,N_7920);
and U12035 (N_12035,N_9713,N_6868);
or U12036 (N_12036,N_9638,N_7778);
nand U12037 (N_12037,N_6421,N_9587);
and U12038 (N_12038,N_9255,N_7417);
nor U12039 (N_12039,N_6748,N_8308);
or U12040 (N_12040,N_6775,N_8517);
nor U12041 (N_12041,N_9258,N_6810);
nand U12042 (N_12042,N_5546,N_9697);
xor U12043 (N_12043,N_6166,N_9509);
nand U12044 (N_12044,N_8780,N_9463);
and U12045 (N_12045,N_7054,N_6400);
nand U12046 (N_12046,N_7642,N_6618);
xor U12047 (N_12047,N_8094,N_5974);
xor U12048 (N_12048,N_8823,N_7943);
nand U12049 (N_12049,N_5587,N_9213);
xnor U12050 (N_12050,N_5740,N_9177);
nor U12051 (N_12051,N_8381,N_6730);
and U12052 (N_12052,N_8586,N_5911);
or U12053 (N_12053,N_6043,N_6435);
and U12054 (N_12054,N_5841,N_9113);
nor U12055 (N_12055,N_5016,N_5249);
nand U12056 (N_12056,N_5584,N_5936);
nor U12057 (N_12057,N_5518,N_9253);
and U12058 (N_12058,N_9331,N_7698);
nor U12059 (N_12059,N_5142,N_5583);
or U12060 (N_12060,N_8868,N_6451);
and U12061 (N_12061,N_5922,N_5996);
or U12062 (N_12062,N_6820,N_7863);
and U12063 (N_12063,N_6853,N_8905);
nand U12064 (N_12064,N_9027,N_8968);
and U12065 (N_12065,N_5515,N_6173);
nor U12066 (N_12066,N_9138,N_8004);
nand U12067 (N_12067,N_7385,N_6862);
and U12068 (N_12068,N_8907,N_7022);
and U12069 (N_12069,N_8619,N_6077);
xor U12070 (N_12070,N_7724,N_8017);
xnor U12071 (N_12071,N_5619,N_5979);
nor U12072 (N_12072,N_8671,N_7035);
nor U12073 (N_12073,N_8846,N_9321);
xnor U12074 (N_12074,N_8397,N_7915);
nand U12075 (N_12075,N_5021,N_7727);
and U12076 (N_12076,N_7917,N_9909);
or U12077 (N_12077,N_5663,N_8113);
and U12078 (N_12078,N_5365,N_8344);
xor U12079 (N_12079,N_6821,N_5507);
or U12080 (N_12080,N_7172,N_6329);
or U12081 (N_12081,N_7448,N_5710);
nor U12082 (N_12082,N_7756,N_7652);
and U12083 (N_12083,N_8063,N_9990);
nand U12084 (N_12084,N_7133,N_7090);
or U12085 (N_12085,N_7847,N_8550);
xnor U12086 (N_12086,N_5861,N_6839);
nand U12087 (N_12087,N_5805,N_6000);
or U12088 (N_12088,N_7860,N_9775);
or U12089 (N_12089,N_7892,N_6608);
xor U12090 (N_12090,N_8703,N_9499);
nand U12091 (N_12091,N_7721,N_8911);
or U12092 (N_12092,N_6255,N_9170);
or U12093 (N_12093,N_8678,N_6457);
nand U12094 (N_12094,N_9526,N_6652);
xor U12095 (N_12095,N_9262,N_8458);
nor U12096 (N_12096,N_8272,N_8252);
nand U12097 (N_12097,N_9812,N_8918);
xor U12098 (N_12098,N_7302,N_5749);
nor U12099 (N_12099,N_8064,N_9444);
or U12100 (N_12100,N_9481,N_8368);
xnor U12101 (N_12101,N_9536,N_5697);
nor U12102 (N_12102,N_5030,N_6617);
and U12103 (N_12103,N_7854,N_9977);
or U12104 (N_12104,N_6038,N_7485);
nand U12105 (N_12105,N_8684,N_7278);
nor U12106 (N_12106,N_5059,N_5991);
xor U12107 (N_12107,N_6019,N_9094);
or U12108 (N_12108,N_7739,N_7780);
and U12109 (N_12109,N_7835,N_7383);
nor U12110 (N_12110,N_9578,N_8822);
and U12111 (N_12111,N_6017,N_5951);
or U12112 (N_12112,N_8469,N_7190);
and U12113 (N_12113,N_8436,N_6669);
and U12114 (N_12114,N_7193,N_9447);
nand U12115 (N_12115,N_7165,N_5658);
and U12116 (N_12116,N_7785,N_5387);
xor U12117 (N_12117,N_6599,N_9135);
nand U12118 (N_12118,N_6612,N_7602);
or U12119 (N_12119,N_8069,N_5850);
nor U12120 (N_12120,N_8104,N_5792);
and U12121 (N_12121,N_9133,N_6531);
and U12122 (N_12122,N_9273,N_5445);
or U12123 (N_12123,N_5992,N_5745);
nand U12124 (N_12124,N_9023,N_9840);
or U12125 (N_12125,N_9058,N_5211);
and U12126 (N_12126,N_6041,N_7145);
and U12127 (N_12127,N_5166,N_5065);
xor U12128 (N_12128,N_9576,N_7288);
or U12129 (N_12129,N_6892,N_7668);
nand U12130 (N_12130,N_7765,N_5607);
or U12131 (N_12131,N_6770,N_9683);
and U12132 (N_12132,N_8692,N_5872);
nand U12133 (N_12133,N_5882,N_8268);
or U12134 (N_12134,N_8742,N_9157);
or U12135 (N_12135,N_9887,N_6015);
xnor U12136 (N_12136,N_7660,N_9817);
nand U12137 (N_12137,N_9345,N_8959);
xnor U12138 (N_12138,N_9313,N_6051);
nor U12139 (N_12139,N_5190,N_7219);
or U12140 (N_12140,N_6086,N_6955);
xnor U12141 (N_12141,N_6938,N_7836);
nand U12142 (N_12142,N_8899,N_6654);
xnor U12143 (N_12143,N_5348,N_7207);
xor U12144 (N_12144,N_8967,N_6392);
nand U12145 (N_12145,N_5877,N_8933);
nor U12146 (N_12146,N_6639,N_5756);
xnor U12147 (N_12147,N_7060,N_9015);
xnor U12148 (N_12148,N_8993,N_6529);
nor U12149 (N_12149,N_8157,N_5092);
or U12150 (N_12150,N_9997,N_6559);
nand U12151 (N_12151,N_7828,N_9307);
and U12152 (N_12152,N_7579,N_8396);
or U12153 (N_12153,N_7846,N_9762);
xnor U12154 (N_12154,N_9987,N_8403);
nand U12155 (N_12155,N_6951,N_8116);
and U12156 (N_12156,N_8467,N_6764);
xnor U12157 (N_12157,N_6563,N_8056);
or U12158 (N_12158,N_8807,N_9372);
and U12159 (N_12159,N_8727,N_5071);
xor U12160 (N_12160,N_5645,N_8416);
or U12161 (N_12161,N_6089,N_6977);
and U12162 (N_12162,N_8815,N_9320);
nand U12163 (N_12163,N_6578,N_7692);
or U12164 (N_12164,N_5433,N_8251);
or U12165 (N_12165,N_8148,N_7555);
nor U12166 (N_12166,N_5018,N_6401);
nand U12167 (N_12167,N_5717,N_7478);
nand U12168 (N_12168,N_5942,N_8963);
or U12169 (N_12169,N_7553,N_8145);
nand U12170 (N_12170,N_9259,N_8003);
nand U12171 (N_12171,N_5641,N_8206);
nor U12172 (N_12172,N_9387,N_6489);
and U12173 (N_12173,N_7275,N_8129);
or U12174 (N_12174,N_9248,N_9753);
and U12175 (N_12175,N_7258,N_5455);
or U12176 (N_12176,N_8534,N_7002);
nor U12177 (N_12177,N_5278,N_5846);
xor U12178 (N_12178,N_6851,N_7138);
or U12179 (N_12179,N_6744,N_6522);
nand U12180 (N_12180,N_6946,N_8385);
nor U12181 (N_12181,N_7797,N_5574);
xnor U12182 (N_12182,N_7648,N_7994);
nor U12183 (N_12183,N_5610,N_5742);
nand U12184 (N_12184,N_9411,N_9198);
nand U12185 (N_12185,N_9580,N_8260);
xnor U12186 (N_12186,N_8741,N_8881);
nand U12187 (N_12187,N_9291,N_9445);
nand U12188 (N_12188,N_6496,N_9184);
or U12189 (N_12189,N_6843,N_7627);
and U12190 (N_12190,N_7168,N_6517);
xnor U12191 (N_12191,N_6713,N_6309);
nor U12192 (N_12192,N_6659,N_5945);
xor U12193 (N_12193,N_9229,N_9629);
or U12194 (N_12194,N_8367,N_9774);
nor U12195 (N_12195,N_6366,N_8190);
and U12196 (N_12196,N_7372,N_8650);
and U12197 (N_12197,N_5762,N_9831);
xnor U12198 (N_12198,N_6541,N_9729);
or U12199 (N_12199,N_9316,N_6766);
or U12200 (N_12200,N_5372,N_9794);
or U12201 (N_12201,N_6357,N_5196);
and U12202 (N_12202,N_5177,N_8515);
nor U12203 (N_12203,N_7548,N_5470);
xor U12204 (N_12204,N_5700,N_9920);
and U12205 (N_12205,N_5275,N_7018);
and U12206 (N_12206,N_9233,N_5741);
nor U12207 (N_12207,N_6248,N_7998);
nor U12208 (N_12208,N_9192,N_6961);
nor U12209 (N_12209,N_9859,N_6741);
and U12210 (N_12210,N_7801,N_8178);
and U12211 (N_12211,N_7716,N_9614);
xnor U12212 (N_12212,N_9731,N_9221);
and U12213 (N_12213,N_5599,N_9366);
or U12214 (N_12214,N_6728,N_6479);
or U12215 (N_12215,N_5141,N_9653);
xnor U12216 (N_12216,N_9222,N_6203);
nand U12217 (N_12217,N_7654,N_8790);
nor U12218 (N_12218,N_9799,N_9703);
xor U12219 (N_12219,N_8564,N_8304);
nand U12220 (N_12220,N_8648,N_7541);
xnor U12221 (N_12221,N_9508,N_6690);
or U12222 (N_12222,N_9589,N_8626);
nand U12223 (N_12223,N_7068,N_5162);
and U12224 (N_12224,N_8295,N_7104);
nor U12225 (N_12225,N_7477,N_8032);
xnor U12226 (N_12226,N_5871,N_9710);
nor U12227 (N_12227,N_6819,N_9108);
xor U12228 (N_12228,N_6184,N_7178);
or U12229 (N_12229,N_5781,N_5775);
or U12230 (N_12230,N_8873,N_5122);
nand U12231 (N_12231,N_8953,N_5735);
nand U12232 (N_12232,N_9126,N_8043);
or U12233 (N_12233,N_7415,N_8057);
and U12234 (N_12234,N_9645,N_9131);
and U12235 (N_12235,N_9019,N_9060);
nor U12236 (N_12236,N_6380,N_7205);
or U12237 (N_12237,N_7293,N_9963);
and U12238 (N_12238,N_6163,N_7982);
nor U12239 (N_12239,N_7821,N_7744);
xor U12240 (N_12240,N_5828,N_6459);
nor U12241 (N_12241,N_6419,N_5811);
and U12242 (N_12242,N_7598,N_5294);
and U12243 (N_12243,N_9621,N_6915);
or U12244 (N_12244,N_6624,N_7463);
nor U12245 (N_12245,N_5298,N_5083);
and U12246 (N_12246,N_9243,N_7864);
nor U12247 (N_12247,N_7311,N_5698);
nand U12248 (N_12248,N_9006,N_8725);
or U12249 (N_12249,N_5649,N_8879);
nor U12250 (N_12250,N_6610,N_8816);
xor U12251 (N_12251,N_6448,N_6388);
nand U12252 (N_12252,N_9704,N_6131);
nor U12253 (N_12253,N_7239,N_9119);
and U12254 (N_12254,N_5993,N_8864);
nand U12255 (N_12255,N_7990,N_7072);
or U12256 (N_12256,N_5235,N_5821);
and U12257 (N_12257,N_7280,N_8219);
xnor U12258 (N_12258,N_7891,N_5565);
and U12259 (N_12259,N_5271,N_6505);
and U12260 (N_12260,N_6050,N_5097);
nor U12261 (N_12261,N_6469,N_8872);
nand U12262 (N_12262,N_8493,N_7236);
xnor U12263 (N_12263,N_8495,N_7661);
xnor U12264 (N_12264,N_5307,N_5703);
nand U12265 (N_12265,N_7105,N_6237);
xor U12266 (N_12266,N_9534,N_6369);
nand U12267 (N_12267,N_7111,N_6978);
xor U12268 (N_12268,N_6665,N_8849);
nor U12269 (N_12269,N_7695,N_9777);
or U12270 (N_12270,N_6259,N_9551);
nand U12271 (N_12271,N_7466,N_6949);
nand U12272 (N_12272,N_7681,N_9327);
nand U12273 (N_12273,N_9391,N_5230);
nand U12274 (N_12274,N_8349,N_5894);
and U12275 (N_12275,N_8418,N_5509);
and U12276 (N_12276,N_7277,N_8283);
nand U12277 (N_12277,N_5787,N_5170);
xor U12278 (N_12278,N_6676,N_6918);
nand U12279 (N_12279,N_5918,N_6418);
nor U12280 (N_12280,N_9824,N_8614);
nand U12281 (N_12281,N_6109,N_7080);
or U12282 (N_12282,N_9692,N_6987);
and U12283 (N_12283,N_9256,N_5739);
or U12284 (N_12284,N_6873,N_8487);
nor U12285 (N_12285,N_5068,N_6545);
and U12286 (N_12286,N_7878,N_9827);
xnor U12287 (N_12287,N_7718,N_6437);
or U12288 (N_12288,N_6120,N_5321);
or U12289 (N_12289,N_5731,N_6614);
nor U12290 (N_12290,N_7742,N_9469);
nor U12291 (N_12291,N_6931,N_5101);
or U12292 (N_12292,N_5146,N_8293);
or U12293 (N_12293,N_6877,N_6808);
or U12294 (N_12294,N_5813,N_7194);
xnor U12295 (N_12295,N_8277,N_8312);
and U12296 (N_12296,N_9848,N_7201);
nor U12297 (N_12297,N_8717,N_5935);
or U12298 (N_12298,N_8194,N_7918);
and U12299 (N_12299,N_8546,N_6805);
xor U12300 (N_12300,N_8576,N_5169);
and U12301 (N_12301,N_8097,N_9092);
xor U12302 (N_12302,N_8926,N_5002);
nor U12303 (N_12303,N_9592,N_5017);
or U12304 (N_12304,N_9919,N_9457);
nor U12305 (N_12305,N_9190,N_5382);
xnor U12306 (N_12306,N_8144,N_5959);
nand U12307 (N_12307,N_8643,N_7819);
or U12308 (N_12308,N_8600,N_9189);
nor U12309 (N_12309,N_8319,N_9335);
and U12310 (N_12310,N_6238,N_6965);
nand U12311 (N_12311,N_7517,N_5302);
and U12312 (N_12312,N_9833,N_8673);
or U12313 (N_12313,N_8325,N_7276);
xor U12314 (N_12314,N_6273,N_6085);
xnor U12315 (N_12315,N_6536,N_8813);
xor U12316 (N_12316,N_5921,N_9636);
and U12317 (N_12317,N_6250,N_8285);
or U12318 (N_12318,N_8232,N_8940);
and U12319 (N_12319,N_9264,N_5400);
xnor U12320 (N_12320,N_8569,N_6312);
xor U12321 (N_12321,N_5848,N_5800);
or U12322 (N_12322,N_8208,N_5069);
xnor U12323 (N_12323,N_6725,N_8641);
nand U12324 (N_12324,N_6199,N_8530);
xnor U12325 (N_12325,N_8665,N_9056);
nor U12326 (N_12326,N_8711,N_5806);
nor U12327 (N_12327,N_9761,N_9650);
nand U12328 (N_12328,N_5887,N_7171);
or U12329 (N_12329,N_9791,N_5965);
nor U12330 (N_12330,N_9506,N_5580);
xor U12331 (N_12331,N_5614,N_6028);
or U12332 (N_12332,N_5970,N_8001);
and U12333 (N_12333,N_8700,N_9368);
and U12334 (N_12334,N_6856,N_5801);
nand U12335 (N_12335,N_8579,N_6637);
and U12336 (N_12336,N_5715,N_8460);
or U12337 (N_12337,N_7564,N_6031);
nand U12338 (N_12338,N_6664,N_8259);
xor U12339 (N_12339,N_5917,N_9823);
xnor U12340 (N_12340,N_8793,N_9384);
nor U12341 (N_12341,N_9516,N_7362);
nor U12342 (N_12342,N_7795,N_5187);
nand U12343 (N_12343,N_6119,N_6195);
xor U12344 (N_12344,N_8640,N_8931);
and U12345 (N_12345,N_5467,N_9070);
nand U12346 (N_12346,N_9889,N_5920);
xnor U12347 (N_12347,N_8912,N_8111);
nor U12348 (N_12348,N_8336,N_9456);
or U12349 (N_12349,N_9197,N_7241);
or U12350 (N_12350,N_9003,N_5899);
and U12351 (N_12351,N_9328,N_6261);
nand U12352 (N_12352,N_7861,N_6431);
or U12353 (N_12353,N_8274,N_6797);
nand U12354 (N_12354,N_9083,N_6251);
and U12355 (N_12355,N_8651,N_7435);
and U12356 (N_12356,N_6304,N_7356);
nor U12357 (N_12357,N_5179,N_8604);
or U12358 (N_12358,N_9018,N_9332);
xnor U12359 (N_12359,N_7501,N_6073);
nor U12360 (N_12360,N_7322,N_9136);
xor U12361 (N_12361,N_5835,N_8160);
xnor U12362 (N_12362,N_5555,N_7646);
xor U12363 (N_12363,N_6176,N_8039);
nand U12364 (N_12364,N_9736,N_9740);
or U12365 (N_12365,N_6611,N_8810);
and U12366 (N_12366,N_6075,N_9519);
and U12367 (N_12367,N_9961,N_7482);
and U12368 (N_12368,N_8076,N_9360);
nand U12369 (N_12369,N_8376,N_8950);
nand U12370 (N_12370,N_5034,N_7237);
or U12371 (N_12371,N_8027,N_9995);
xnor U12372 (N_12372,N_7907,N_5523);
nand U12373 (N_12373,N_6719,N_9989);
or U12374 (N_12374,N_5939,N_8856);
or U12375 (N_12375,N_7979,N_7641);
and U12376 (N_12376,N_8425,N_9021);
xnor U12377 (N_12377,N_5063,N_6794);
xnor U12378 (N_12378,N_5532,N_6838);
nand U12379 (N_12379,N_8693,N_7083);
xor U12380 (N_12380,N_5589,N_8058);
xnor U12381 (N_12381,N_8421,N_7094);
nor U12382 (N_12382,N_5567,N_6602);
xor U12383 (N_12383,N_7667,N_7822);
nor U12384 (N_12384,N_6601,N_5362);
or U12385 (N_12385,N_6111,N_9115);
nand U12386 (N_12386,N_6634,N_8885);
nand U12387 (N_12387,N_9604,N_7307);
and U12388 (N_12388,N_7634,N_8927);
xor U12389 (N_12389,N_7502,N_5410);
and U12390 (N_12390,N_7844,N_5091);
xnor U12391 (N_12391,N_6682,N_5157);
nor U12392 (N_12392,N_5329,N_5516);
and U12393 (N_12393,N_9974,N_5621);
nor U12394 (N_12394,N_8947,N_5934);
nor U12395 (N_12395,N_8379,N_9035);
or U12396 (N_12396,N_8366,N_7099);
nor U12397 (N_12397,N_8505,N_6063);
and U12398 (N_12398,N_5185,N_5783);
and U12399 (N_12399,N_6245,N_9423);
nor U12400 (N_12400,N_6162,N_8335);
nor U12401 (N_12401,N_8053,N_8945);
nand U12402 (N_12402,N_8653,N_7045);
or U12403 (N_12403,N_7697,N_5544);
or U12404 (N_12404,N_6630,N_5916);
nor U12405 (N_12405,N_7330,N_8533);
xnor U12406 (N_12406,N_8382,N_8635);
xnor U12407 (N_12407,N_8837,N_5110);
nand U12408 (N_12408,N_9945,N_5328);
nand U12409 (N_12409,N_6462,N_9028);
and U12410 (N_12410,N_8809,N_9541);
or U12411 (N_12411,N_6711,N_8522);
and U12412 (N_12412,N_5215,N_7215);
nor U12413 (N_12413,N_7586,N_9765);
or U12414 (N_12414,N_9607,N_5461);
xnor U12415 (N_12415,N_8264,N_8037);
or U12416 (N_12416,N_9439,N_7855);
nand U12417 (N_12417,N_6034,N_5175);
and U12418 (N_12418,N_8512,N_6136);
nor U12419 (N_12419,N_8429,N_5247);
or U12420 (N_12420,N_5040,N_6912);
nor U12421 (N_12421,N_8708,N_6934);
nor U12422 (N_12422,N_9030,N_5094);
nand U12423 (N_12423,N_7454,N_9507);
or U12424 (N_12424,N_6930,N_5725);
or U12425 (N_12425,N_7325,N_9847);
nor U12426 (N_12426,N_7371,N_6948);
or U12427 (N_12427,N_7320,N_7761);
and U12428 (N_12428,N_6315,N_5684);
nand U12429 (N_12429,N_8556,N_8901);
nand U12430 (N_12430,N_8025,N_7740);
and U12431 (N_12431,N_8524,N_5598);
nand U12432 (N_12432,N_6845,N_7921);
and U12433 (N_12433,N_9772,N_6589);
xnor U12434 (N_12434,N_6927,N_7808);
xor U12435 (N_12435,N_9005,N_9858);
or U12436 (N_12436,N_8561,N_5292);
nor U12437 (N_12437,N_6635,N_9647);
nand U12438 (N_12438,N_7601,N_9359);
xor U12439 (N_12439,N_8033,N_6587);
or U12440 (N_12440,N_7958,N_6193);
xor U12441 (N_12441,N_5459,N_8189);
nor U12442 (N_12442,N_8618,N_7467);
or U12443 (N_12443,N_5241,N_6117);
xnor U12444 (N_12444,N_6284,N_6550);
nor U12445 (N_12445,N_8620,N_5667);
or U12446 (N_12446,N_5451,N_9566);
nor U12447 (N_12447,N_6538,N_7451);
and U12448 (N_12448,N_6607,N_7059);
nor U12449 (N_12449,N_5188,N_9323);
or U12450 (N_12450,N_9337,N_9618);
xor U12451 (N_12451,N_7589,N_8475);
or U12452 (N_12452,N_7657,N_6499);
nor U12453 (N_12453,N_6275,N_5133);
or U12454 (N_12454,N_6568,N_8016);
nand U12455 (N_12455,N_7729,N_7089);
nand U12456 (N_12456,N_9539,N_9408);
xor U12457 (N_12457,N_7329,N_6880);
nand U12458 (N_12458,N_7503,N_7963);
nor U12459 (N_12459,N_8338,N_5440);
nor U12460 (N_12460,N_8855,N_7874);
nor U12461 (N_12461,N_9577,N_9437);
nor U12462 (N_12462,N_7348,N_5426);
nand U12463 (N_12463,N_8188,N_8106);
nor U12464 (N_12464,N_5054,N_5485);
xnor U12465 (N_12465,N_6274,N_9020);
nor U12466 (N_12466,N_7106,N_6647);
xnor U12467 (N_12467,N_6990,N_9024);
nand U12468 (N_12468,N_6198,N_7817);
and U12469 (N_12469,N_8292,N_7033);
nand U12470 (N_12470,N_5073,N_9738);
nor U12471 (N_12471,N_7591,N_6300);
nand U12472 (N_12472,N_9726,N_8212);
nor U12473 (N_12473,N_7782,N_6552);
nand U12474 (N_12474,N_5849,N_6855);
nand U12475 (N_12475,N_6494,N_5556);
or U12476 (N_12476,N_5502,N_9800);
xnor U12477 (N_12477,N_8669,N_6254);
nand U12478 (N_12478,N_8791,N_5345);
nor U12479 (N_12479,N_8289,N_7637);
nand U12480 (N_12480,N_6526,N_7513);
xnor U12481 (N_12481,N_8591,N_9973);
xnor U12482 (N_12482,N_8509,N_8288);
xor U12483 (N_12483,N_9933,N_8572);
nand U12484 (N_12484,N_8395,N_8975);
nor U12485 (N_12485,N_5401,N_5634);
nand U12486 (N_12486,N_8943,N_9470);
and U12487 (N_12487,N_7672,N_6588);
and U12488 (N_12488,N_5864,N_5998);
and U12489 (N_12489,N_9891,N_9644);
nand U12490 (N_12490,N_5794,N_7279);
nor U12491 (N_12491,N_5143,N_6142);
nor U12492 (N_12492,N_9302,N_5985);
or U12493 (N_12493,N_6888,N_9939);
and U12494 (N_12494,N_5126,N_5753);
xor U12495 (N_12495,N_6213,N_6175);
or U12496 (N_12496,N_6561,N_5355);
and U12497 (N_12497,N_5748,N_8563);
nand U12498 (N_12498,N_7474,N_6569);
nand U12499 (N_12499,N_5737,N_8450);
nor U12500 (N_12500,N_9286,N_6501);
nor U12501 (N_12501,N_8355,N_9192);
nor U12502 (N_12502,N_5552,N_8520);
or U12503 (N_12503,N_8830,N_6440);
nand U12504 (N_12504,N_5687,N_9876);
or U12505 (N_12505,N_9654,N_5438);
xnor U12506 (N_12506,N_5962,N_5983);
xnor U12507 (N_12507,N_5952,N_7318);
xor U12508 (N_12508,N_5548,N_7784);
nand U12509 (N_12509,N_7164,N_8470);
and U12510 (N_12510,N_9762,N_6186);
nor U12511 (N_12511,N_5883,N_9044);
and U12512 (N_12512,N_8295,N_9727);
and U12513 (N_12513,N_7340,N_8894);
or U12514 (N_12514,N_9395,N_8191);
and U12515 (N_12515,N_6275,N_8333);
or U12516 (N_12516,N_7617,N_9206);
nand U12517 (N_12517,N_8676,N_9859);
xor U12518 (N_12518,N_5420,N_8166);
and U12519 (N_12519,N_9381,N_5525);
nor U12520 (N_12520,N_5449,N_7337);
nand U12521 (N_12521,N_7410,N_9125);
xor U12522 (N_12522,N_6803,N_6865);
or U12523 (N_12523,N_9200,N_9863);
xnor U12524 (N_12524,N_7877,N_5454);
nor U12525 (N_12525,N_8819,N_5732);
nor U12526 (N_12526,N_8264,N_5343);
or U12527 (N_12527,N_6754,N_9454);
nor U12528 (N_12528,N_6755,N_8991);
and U12529 (N_12529,N_6006,N_9854);
xor U12530 (N_12530,N_8147,N_9331);
xor U12531 (N_12531,N_9265,N_5788);
and U12532 (N_12532,N_7144,N_9376);
and U12533 (N_12533,N_9154,N_5682);
xor U12534 (N_12534,N_6493,N_5997);
xor U12535 (N_12535,N_5998,N_6925);
xnor U12536 (N_12536,N_8264,N_6092);
nand U12537 (N_12537,N_5026,N_8884);
xnor U12538 (N_12538,N_5806,N_6536);
and U12539 (N_12539,N_5273,N_9344);
nor U12540 (N_12540,N_8730,N_9295);
xor U12541 (N_12541,N_5402,N_5269);
nand U12542 (N_12542,N_5217,N_6404);
or U12543 (N_12543,N_8696,N_6833);
nor U12544 (N_12544,N_6918,N_5308);
xnor U12545 (N_12545,N_7877,N_5540);
and U12546 (N_12546,N_9463,N_8145);
and U12547 (N_12547,N_7496,N_9176);
nand U12548 (N_12548,N_5929,N_6199);
nor U12549 (N_12549,N_6915,N_6303);
xnor U12550 (N_12550,N_9956,N_6279);
nor U12551 (N_12551,N_7027,N_8805);
nand U12552 (N_12552,N_6231,N_7612);
nand U12553 (N_12553,N_7973,N_9559);
nor U12554 (N_12554,N_7679,N_6277);
or U12555 (N_12555,N_7277,N_6479);
or U12556 (N_12556,N_9534,N_6036);
nor U12557 (N_12557,N_9466,N_9879);
nand U12558 (N_12558,N_8820,N_9865);
and U12559 (N_12559,N_8517,N_5943);
nand U12560 (N_12560,N_5157,N_8966);
and U12561 (N_12561,N_8244,N_6965);
xor U12562 (N_12562,N_5361,N_9454);
nor U12563 (N_12563,N_6618,N_6580);
or U12564 (N_12564,N_6158,N_9269);
and U12565 (N_12565,N_5562,N_9196);
nand U12566 (N_12566,N_9088,N_6521);
nor U12567 (N_12567,N_7246,N_9981);
nand U12568 (N_12568,N_9568,N_8188);
nor U12569 (N_12569,N_8095,N_6105);
nor U12570 (N_12570,N_9050,N_5287);
nor U12571 (N_12571,N_8404,N_9783);
and U12572 (N_12572,N_6204,N_6210);
nand U12573 (N_12573,N_7437,N_9003);
nor U12574 (N_12574,N_7479,N_5020);
or U12575 (N_12575,N_5571,N_6120);
and U12576 (N_12576,N_5235,N_7056);
nor U12577 (N_12577,N_9774,N_7550);
nand U12578 (N_12578,N_9623,N_5755);
xnor U12579 (N_12579,N_9329,N_8615);
nand U12580 (N_12580,N_7603,N_6141);
nor U12581 (N_12581,N_5022,N_5882);
xnor U12582 (N_12582,N_5211,N_8290);
or U12583 (N_12583,N_6510,N_5394);
xnor U12584 (N_12584,N_6580,N_6680);
nand U12585 (N_12585,N_8384,N_7496);
nand U12586 (N_12586,N_9073,N_5304);
and U12587 (N_12587,N_5009,N_7964);
or U12588 (N_12588,N_5063,N_6285);
and U12589 (N_12589,N_8369,N_6661);
or U12590 (N_12590,N_9998,N_6967);
and U12591 (N_12591,N_6538,N_5483);
nor U12592 (N_12592,N_7860,N_5224);
and U12593 (N_12593,N_7835,N_6172);
and U12594 (N_12594,N_5549,N_9917);
or U12595 (N_12595,N_8136,N_7381);
and U12596 (N_12596,N_6868,N_5627);
or U12597 (N_12597,N_6230,N_8514);
and U12598 (N_12598,N_8437,N_7426);
nand U12599 (N_12599,N_9880,N_9175);
nand U12600 (N_12600,N_6907,N_8186);
nor U12601 (N_12601,N_5275,N_7221);
or U12602 (N_12602,N_7941,N_8841);
xor U12603 (N_12603,N_9849,N_5987);
or U12604 (N_12604,N_6325,N_9769);
nand U12605 (N_12605,N_7645,N_5006);
and U12606 (N_12606,N_7419,N_8332);
nor U12607 (N_12607,N_9729,N_5716);
nand U12608 (N_12608,N_7185,N_6348);
and U12609 (N_12609,N_8596,N_6525);
nand U12610 (N_12610,N_6756,N_5354);
and U12611 (N_12611,N_8127,N_7730);
nand U12612 (N_12612,N_6957,N_6217);
xor U12613 (N_12613,N_7536,N_5156);
or U12614 (N_12614,N_6234,N_9127);
xnor U12615 (N_12615,N_8925,N_9214);
xnor U12616 (N_12616,N_6409,N_5598);
nor U12617 (N_12617,N_5310,N_5691);
and U12618 (N_12618,N_7458,N_6406);
and U12619 (N_12619,N_7369,N_5508);
nand U12620 (N_12620,N_9567,N_6471);
xor U12621 (N_12621,N_6441,N_7098);
nor U12622 (N_12622,N_5250,N_7731);
nor U12623 (N_12623,N_9544,N_5440);
nor U12624 (N_12624,N_7921,N_9020);
or U12625 (N_12625,N_6668,N_8633);
or U12626 (N_12626,N_6542,N_7960);
and U12627 (N_12627,N_7484,N_6418);
nand U12628 (N_12628,N_8853,N_7681);
or U12629 (N_12629,N_6907,N_9575);
nor U12630 (N_12630,N_7377,N_8397);
xnor U12631 (N_12631,N_6380,N_7499);
nand U12632 (N_12632,N_6687,N_8439);
xor U12633 (N_12633,N_5879,N_9635);
nor U12634 (N_12634,N_5017,N_7241);
nor U12635 (N_12635,N_5788,N_8342);
nand U12636 (N_12636,N_7892,N_5769);
nor U12637 (N_12637,N_9781,N_9900);
nand U12638 (N_12638,N_7586,N_9921);
nor U12639 (N_12639,N_7051,N_6803);
nand U12640 (N_12640,N_6387,N_5986);
or U12641 (N_12641,N_7592,N_8420);
and U12642 (N_12642,N_7649,N_8796);
nor U12643 (N_12643,N_7339,N_5460);
nor U12644 (N_12644,N_5693,N_7607);
and U12645 (N_12645,N_7526,N_5442);
nor U12646 (N_12646,N_9896,N_9248);
or U12647 (N_12647,N_7853,N_6511);
nand U12648 (N_12648,N_8005,N_6582);
nand U12649 (N_12649,N_7102,N_8463);
and U12650 (N_12650,N_6741,N_8015);
and U12651 (N_12651,N_5023,N_7823);
nand U12652 (N_12652,N_8932,N_5211);
xnor U12653 (N_12653,N_5217,N_6778);
xnor U12654 (N_12654,N_5964,N_7503);
or U12655 (N_12655,N_8646,N_8725);
nand U12656 (N_12656,N_7627,N_8406);
or U12657 (N_12657,N_8810,N_8179);
nand U12658 (N_12658,N_7208,N_5351);
or U12659 (N_12659,N_5442,N_8215);
nor U12660 (N_12660,N_7081,N_7382);
nand U12661 (N_12661,N_7775,N_5502);
and U12662 (N_12662,N_6239,N_7705);
or U12663 (N_12663,N_7089,N_8506);
nand U12664 (N_12664,N_9250,N_5609);
nand U12665 (N_12665,N_6556,N_6137);
nor U12666 (N_12666,N_6057,N_7911);
nand U12667 (N_12667,N_6642,N_8941);
or U12668 (N_12668,N_5071,N_7604);
nor U12669 (N_12669,N_7785,N_6643);
or U12670 (N_12670,N_8780,N_5574);
and U12671 (N_12671,N_8240,N_9802);
xnor U12672 (N_12672,N_9226,N_7044);
and U12673 (N_12673,N_7449,N_7349);
xnor U12674 (N_12674,N_5295,N_9170);
or U12675 (N_12675,N_7446,N_9015);
nand U12676 (N_12676,N_7807,N_9408);
xor U12677 (N_12677,N_9524,N_8853);
or U12678 (N_12678,N_5492,N_5221);
nand U12679 (N_12679,N_6157,N_9895);
and U12680 (N_12680,N_7294,N_6667);
nor U12681 (N_12681,N_8157,N_5814);
xnor U12682 (N_12682,N_8050,N_9053);
xor U12683 (N_12683,N_9658,N_9576);
nor U12684 (N_12684,N_8472,N_8884);
nor U12685 (N_12685,N_5955,N_9457);
nor U12686 (N_12686,N_8804,N_5567);
and U12687 (N_12687,N_6169,N_8657);
nand U12688 (N_12688,N_7477,N_5602);
or U12689 (N_12689,N_8460,N_6695);
and U12690 (N_12690,N_9196,N_9083);
nor U12691 (N_12691,N_7477,N_9475);
and U12692 (N_12692,N_8279,N_7564);
or U12693 (N_12693,N_8280,N_8380);
nand U12694 (N_12694,N_5181,N_7800);
nand U12695 (N_12695,N_7437,N_9438);
nand U12696 (N_12696,N_9373,N_8477);
nor U12697 (N_12697,N_9516,N_8188);
or U12698 (N_12698,N_6366,N_5232);
nor U12699 (N_12699,N_5451,N_8321);
xor U12700 (N_12700,N_7817,N_7724);
xor U12701 (N_12701,N_8817,N_8581);
or U12702 (N_12702,N_6574,N_5058);
nand U12703 (N_12703,N_8242,N_6168);
nor U12704 (N_12704,N_6342,N_9646);
or U12705 (N_12705,N_6499,N_5249);
nor U12706 (N_12706,N_6433,N_7054);
and U12707 (N_12707,N_7896,N_6532);
nor U12708 (N_12708,N_8574,N_7726);
xor U12709 (N_12709,N_8916,N_6709);
nor U12710 (N_12710,N_9802,N_8650);
xnor U12711 (N_12711,N_9404,N_5748);
nand U12712 (N_12712,N_7243,N_6788);
nor U12713 (N_12713,N_5673,N_9312);
and U12714 (N_12714,N_9133,N_6839);
nor U12715 (N_12715,N_7952,N_5238);
or U12716 (N_12716,N_8875,N_6320);
xor U12717 (N_12717,N_5460,N_9606);
xnor U12718 (N_12718,N_6114,N_7124);
and U12719 (N_12719,N_6036,N_8508);
nand U12720 (N_12720,N_5139,N_6861);
or U12721 (N_12721,N_6144,N_7679);
and U12722 (N_12722,N_5311,N_7204);
or U12723 (N_12723,N_6246,N_8389);
nand U12724 (N_12724,N_9036,N_9659);
and U12725 (N_12725,N_5527,N_9581);
and U12726 (N_12726,N_6224,N_5517);
nor U12727 (N_12727,N_8843,N_6446);
xor U12728 (N_12728,N_6590,N_8339);
nor U12729 (N_12729,N_5164,N_5435);
nand U12730 (N_12730,N_9535,N_9867);
or U12731 (N_12731,N_5919,N_5920);
nand U12732 (N_12732,N_9770,N_9745);
or U12733 (N_12733,N_7204,N_5780);
nand U12734 (N_12734,N_8576,N_6781);
xor U12735 (N_12735,N_7427,N_9115);
nand U12736 (N_12736,N_6297,N_9444);
and U12737 (N_12737,N_9413,N_7512);
or U12738 (N_12738,N_9842,N_8720);
nand U12739 (N_12739,N_9821,N_7325);
nor U12740 (N_12740,N_7407,N_8139);
and U12741 (N_12741,N_6155,N_9513);
nor U12742 (N_12742,N_5311,N_6818);
xor U12743 (N_12743,N_9604,N_5164);
and U12744 (N_12744,N_8985,N_6235);
nand U12745 (N_12745,N_5398,N_7421);
nor U12746 (N_12746,N_5229,N_7360);
or U12747 (N_12747,N_8566,N_6836);
nor U12748 (N_12748,N_9186,N_5893);
xor U12749 (N_12749,N_8367,N_6932);
and U12750 (N_12750,N_6526,N_6982);
xnor U12751 (N_12751,N_5518,N_5871);
nand U12752 (N_12752,N_7876,N_9382);
or U12753 (N_12753,N_6491,N_8199);
xnor U12754 (N_12754,N_9807,N_9990);
or U12755 (N_12755,N_6895,N_8582);
xnor U12756 (N_12756,N_8347,N_5394);
nor U12757 (N_12757,N_9991,N_5816);
or U12758 (N_12758,N_7467,N_9946);
nand U12759 (N_12759,N_8308,N_8020);
and U12760 (N_12760,N_9405,N_9663);
or U12761 (N_12761,N_7086,N_9624);
or U12762 (N_12762,N_5045,N_9551);
and U12763 (N_12763,N_6500,N_5671);
and U12764 (N_12764,N_5567,N_9417);
and U12765 (N_12765,N_7631,N_9909);
or U12766 (N_12766,N_8356,N_6859);
nand U12767 (N_12767,N_6456,N_9192);
and U12768 (N_12768,N_8344,N_6640);
or U12769 (N_12769,N_5235,N_7740);
and U12770 (N_12770,N_6180,N_9115);
and U12771 (N_12771,N_7200,N_7070);
xnor U12772 (N_12772,N_8076,N_5807);
and U12773 (N_12773,N_9239,N_6711);
and U12774 (N_12774,N_9804,N_6879);
nand U12775 (N_12775,N_7334,N_9638);
and U12776 (N_12776,N_5612,N_9957);
or U12777 (N_12777,N_8379,N_8720);
and U12778 (N_12778,N_9656,N_6632);
nor U12779 (N_12779,N_8136,N_6854);
and U12780 (N_12780,N_6693,N_8669);
nand U12781 (N_12781,N_7227,N_6393);
xnor U12782 (N_12782,N_8208,N_5709);
nor U12783 (N_12783,N_6980,N_6969);
nor U12784 (N_12784,N_8449,N_7197);
xor U12785 (N_12785,N_5892,N_9073);
xor U12786 (N_12786,N_6935,N_9157);
nor U12787 (N_12787,N_7391,N_7620);
and U12788 (N_12788,N_7530,N_9970);
xnor U12789 (N_12789,N_7975,N_8067);
nor U12790 (N_12790,N_7947,N_5374);
nor U12791 (N_12791,N_8905,N_5502);
or U12792 (N_12792,N_7079,N_6964);
nor U12793 (N_12793,N_6359,N_8043);
and U12794 (N_12794,N_6240,N_7076);
nor U12795 (N_12795,N_5429,N_8014);
or U12796 (N_12796,N_6743,N_7159);
nand U12797 (N_12797,N_7019,N_6178);
xor U12798 (N_12798,N_6360,N_7605);
and U12799 (N_12799,N_8206,N_8683);
or U12800 (N_12800,N_5751,N_6968);
nor U12801 (N_12801,N_8581,N_9090);
nand U12802 (N_12802,N_8311,N_5346);
and U12803 (N_12803,N_5463,N_5384);
and U12804 (N_12804,N_6482,N_7046);
nor U12805 (N_12805,N_8573,N_8601);
nand U12806 (N_12806,N_6008,N_9704);
nor U12807 (N_12807,N_8701,N_5674);
nand U12808 (N_12808,N_6517,N_9386);
nor U12809 (N_12809,N_7295,N_7223);
and U12810 (N_12810,N_5408,N_6382);
nor U12811 (N_12811,N_9454,N_6092);
or U12812 (N_12812,N_5661,N_8455);
nor U12813 (N_12813,N_7979,N_8744);
nor U12814 (N_12814,N_7602,N_7262);
nor U12815 (N_12815,N_7612,N_5226);
and U12816 (N_12816,N_6059,N_5576);
nand U12817 (N_12817,N_8768,N_6833);
nor U12818 (N_12818,N_9594,N_6440);
nor U12819 (N_12819,N_5219,N_8382);
xor U12820 (N_12820,N_8517,N_9090);
and U12821 (N_12821,N_7313,N_6524);
nor U12822 (N_12822,N_8398,N_6737);
or U12823 (N_12823,N_6110,N_9195);
and U12824 (N_12824,N_5937,N_7199);
xor U12825 (N_12825,N_6279,N_5363);
or U12826 (N_12826,N_9753,N_9656);
or U12827 (N_12827,N_7169,N_7059);
nand U12828 (N_12828,N_6479,N_5161);
and U12829 (N_12829,N_7180,N_6742);
xor U12830 (N_12830,N_7186,N_8317);
or U12831 (N_12831,N_9371,N_5863);
and U12832 (N_12832,N_9874,N_6374);
nand U12833 (N_12833,N_5617,N_9457);
xnor U12834 (N_12834,N_9570,N_6585);
and U12835 (N_12835,N_9806,N_5337);
and U12836 (N_12836,N_9159,N_7297);
nand U12837 (N_12837,N_8636,N_9192);
xor U12838 (N_12838,N_8757,N_6731);
xor U12839 (N_12839,N_9826,N_9832);
and U12840 (N_12840,N_8983,N_9251);
or U12841 (N_12841,N_9272,N_9994);
nor U12842 (N_12842,N_8819,N_6574);
and U12843 (N_12843,N_6126,N_6106);
and U12844 (N_12844,N_6625,N_7876);
xor U12845 (N_12845,N_9909,N_5735);
and U12846 (N_12846,N_6446,N_7585);
or U12847 (N_12847,N_5889,N_6951);
and U12848 (N_12848,N_8613,N_9115);
nand U12849 (N_12849,N_7799,N_9068);
and U12850 (N_12850,N_7829,N_8226);
nand U12851 (N_12851,N_7370,N_8863);
and U12852 (N_12852,N_8959,N_8439);
and U12853 (N_12853,N_5688,N_6683);
and U12854 (N_12854,N_7917,N_9337);
nand U12855 (N_12855,N_9878,N_8099);
xnor U12856 (N_12856,N_6997,N_5500);
nor U12857 (N_12857,N_6104,N_6441);
nand U12858 (N_12858,N_5439,N_9151);
xnor U12859 (N_12859,N_7663,N_7551);
or U12860 (N_12860,N_5707,N_9151);
nor U12861 (N_12861,N_7059,N_8928);
nand U12862 (N_12862,N_9226,N_6105);
or U12863 (N_12863,N_7864,N_6074);
xnor U12864 (N_12864,N_7110,N_6155);
xor U12865 (N_12865,N_9875,N_5699);
nand U12866 (N_12866,N_8139,N_6433);
or U12867 (N_12867,N_8080,N_7160);
xor U12868 (N_12868,N_5905,N_6438);
xnor U12869 (N_12869,N_9885,N_8241);
xnor U12870 (N_12870,N_5929,N_8577);
xnor U12871 (N_12871,N_7490,N_6852);
nand U12872 (N_12872,N_8804,N_7074);
and U12873 (N_12873,N_7748,N_6353);
nand U12874 (N_12874,N_7726,N_9232);
or U12875 (N_12875,N_7723,N_6013);
nand U12876 (N_12876,N_9320,N_6119);
xnor U12877 (N_12877,N_5843,N_8423);
nor U12878 (N_12878,N_8338,N_9749);
nand U12879 (N_12879,N_5498,N_5371);
and U12880 (N_12880,N_9413,N_5739);
xnor U12881 (N_12881,N_7589,N_8467);
and U12882 (N_12882,N_9698,N_6531);
nor U12883 (N_12883,N_7829,N_7400);
or U12884 (N_12884,N_5548,N_6836);
nor U12885 (N_12885,N_5953,N_9210);
nor U12886 (N_12886,N_7706,N_6917);
and U12887 (N_12887,N_7687,N_5648);
or U12888 (N_12888,N_6930,N_9515);
nor U12889 (N_12889,N_5600,N_5481);
nand U12890 (N_12890,N_9696,N_9851);
nor U12891 (N_12891,N_6866,N_9243);
nand U12892 (N_12892,N_8351,N_9617);
xor U12893 (N_12893,N_7063,N_6314);
xor U12894 (N_12894,N_9026,N_5598);
xor U12895 (N_12895,N_5613,N_7692);
or U12896 (N_12896,N_9274,N_6898);
nand U12897 (N_12897,N_7515,N_8774);
or U12898 (N_12898,N_9167,N_6911);
nand U12899 (N_12899,N_8874,N_7316);
nor U12900 (N_12900,N_8970,N_8275);
or U12901 (N_12901,N_9704,N_6630);
nand U12902 (N_12902,N_7961,N_5770);
and U12903 (N_12903,N_9636,N_7922);
and U12904 (N_12904,N_5967,N_7392);
nor U12905 (N_12905,N_6710,N_8732);
xnor U12906 (N_12906,N_9316,N_7642);
or U12907 (N_12907,N_9381,N_6733);
xnor U12908 (N_12908,N_7206,N_8736);
nand U12909 (N_12909,N_9711,N_7191);
nand U12910 (N_12910,N_9707,N_8253);
or U12911 (N_12911,N_7212,N_9014);
xnor U12912 (N_12912,N_8939,N_9633);
nand U12913 (N_12913,N_6490,N_7226);
nor U12914 (N_12914,N_7942,N_5860);
nand U12915 (N_12915,N_5216,N_5072);
nand U12916 (N_12916,N_6435,N_8720);
nor U12917 (N_12917,N_6472,N_6873);
xor U12918 (N_12918,N_7751,N_7924);
and U12919 (N_12919,N_9417,N_6732);
and U12920 (N_12920,N_8353,N_7888);
or U12921 (N_12921,N_9335,N_5709);
nor U12922 (N_12922,N_9970,N_5955);
nor U12923 (N_12923,N_8773,N_8314);
xor U12924 (N_12924,N_9912,N_8864);
nor U12925 (N_12925,N_9549,N_9643);
xor U12926 (N_12926,N_8198,N_5879);
nand U12927 (N_12927,N_7674,N_7572);
nand U12928 (N_12928,N_8146,N_7629);
and U12929 (N_12929,N_8702,N_9209);
or U12930 (N_12930,N_5104,N_5716);
nor U12931 (N_12931,N_5531,N_5409);
nand U12932 (N_12932,N_8102,N_9177);
or U12933 (N_12933,N_9950,N_7557);
nor U12934 (N_12934,N_7286,N_8372);
nor U12935 (N_12935,N_7946,N_5388);
or U12936 (N_12936,N_6910,N_9952);
or U12937 (N_12937,N_7274,N_8836);
xor U12938 (N_12938,N_6719,N_7235);
nand U12939 (N_12939,N_8957,N_5542);
or U12940 (N_12940,N_9353,N_9708);
xnor U12941 (N_12941,N_6482,N_9805);
nand U12942 (N_12942,N_9013,N_8166);
nand U12943 (N_12943,N_5711,N_7236);
nor U12944 (N_12944,N_9459,N_8798);
and U12945 (N_12945,N_6093,N_9589);
xor U12946 (N_12946,N_5684,N_8548);
nand U12947 (N_12947,N_9670,N_6696);
xnor U12948 (N_12948,N_8999,N_8195);
nor U12949 (N_12949,N_9932,N_6641);
xnor U12950 (N_12950,N_6778,N_9358);
or U12951 (N_12951,N_9216,N_8309);
or U12952 (N_12952,N_8617,N_6424);
or U12953 (N_12953,N_8191,N_9440);
and U12954 (N_12954,N_5291,N_9422);
and U12955 (N_12955,N_5621,N_9568);
or U12956 (N_12956,N_9644,N_8716);
xnor U12957 (N_12957,N_7941,N_9589);
nand U12958 (N_12958,N_7784,N_5864);
or U12959 (N_12959,N_6570,N_6919);
and U12960 (N_12960,N_8223,N_9195);
nor U12961 (N_12961,N_9852,N_7673);
nor U12962 (N_12962,N_7205,N_8940);
or U12963 (N_12963,N_9428,N_7840);
and U12964 (N_12964,N_8903,N_7184);
and U12965 (N_12965,N_5238,N_6245);
or U12966 (N_12966,N_8769,N_9249);
xnor U12967 (N_12967,N_6082,N_5014);
nor U12968 (N_12968,N_9336,N_9294);
nand U12969 (N_12969,N_8264,N_6870);
xnor U12970 (N_12970,N_9684,N_9607);
or U12971 (N_12971,N_7129,N_8351);
nor U12972 (N_12972,N_9080,N_9143);
and U12973 (N_12973,N_7423,N_7016);
or U12974 (N_12974,N_9800,N_9725);
and U12975 (N_12975,N_8530,N_5591);
and U12976 (N_12976,N_9879,N_5427);
or U12977 (N_12977,N_5921,N_6397);
and U12978 (N_12978,N_9233,N_9721);
nand U12979 (N_12979,N_7615,N_5477);
nor U12980 (N_12980,N_5030,N_7672);
or U12981 (N_12981,N_7014,N_7670);
xnor U12982 (N_12982,N_9748,N_6179);
or U12983 (N_12983,N_5698,N_6466);
xnor U12984 (N_12984,N_9094,N_6641);
and U12985 (N_12985,N_5903,N_6786);
xnor U12986 (N_12986,N_9370,N_8291);
or U12987 (N_12987,N_7170,N_9839);
nand U12988 (N_12988,N_6672,N_5058);
and U12989 (N_12989,N_9633,N_8633);
and U12990 (N_12990,N_5230,N_9701);
nor U12991 (N_12991,N_7190,N_9897);
nand U12992 (N_12992,N_5563,N_6335);
and U12993 (N_12993,N_9943,N_6923);
nor U12994 (N_12994,N_9674,N_7608);
nand U12995 (N_12995,N_5362,N_9438);
and U12996 (N_12996,N_8335,N_8180);
and U12997 (N_12997,N_6067,N_5229);
or U12998 (N_12998,N_9750,N_7675);
or U12999 (N_12999,N_5652,N_8893);
xnor U13000 (N_13000,N_8093,N_6971);
nor U13001 (N_13001,N_9859,N_8495);
xnor U13002 (N_13002,N_7892,N_7236);
nand U13003 (N_13003,N_9116,N_7166);
xnor U13004 (N_13004,N_7769,N_7235);
nand U13005 (N_13005,N_7360,N_8752);
or U13006 (N_13006,N_5603,N_8302);
xnor U13007 (N_13007,N_5285,N_7265);
nor U13008 (N_13008,N_6325,N_9754);
and U13009 (N_13009,N_5872,N_7925);
and U13010 (N_13010,N_5232,N_8407);
or U13011 (N_13011,N_8416,N_5991);
nor U13012 (N_13012,N_5393,N_5854);
xnor U13013 (N_13013,N_5606,N_7117);
nand U13014 (N_13014,N_6649,N_6580);
nand U13015 (N_13015,N_7239,N_6371);
nand U13016 (N_13016,N_5085,N_9530);
nand U13017 (N_13017,N_8014,N_5856);
nand U13018 (N_13018,N_5007,N_9266);
nor U13019 (N_13019,N_9499,N_6256);
or U13020 (N_13020,N_9281,N_6225);
nor U13021 (N_13021,N_9341,N_8465);
nor U13022 (N_13022,N_5613,N_5570);
or U13023 (N_13023,N_6096,N_9678);
or U13024 (N_13024,N_8051,N_7651);
and U13025 (N_13025,N_5378,N_9222);
xnor U13026 (N_13026,N_8926,N_7514);
and U13027 (N_13027,N_8548,N_9070);
xor U13028 (N_13028,N_8956,N_5524);
and U13029 (N_13029,N_9852,N_8294);
and U13030 (N_13030,N_6125,N_6043);
nand U13031 (N_13031,N_7153,N_7169);
nor U13032 (N_13032,N_7632,N_9297);
nor U13033 (N_13033,N_6198,N_9996);
or U13034 (N_13034,N_7030,N_7199);
or U13035 (N_13035,N_6401,N_8170);
and U13036 (N_13036,N_5206,N_5577);
xor U13037 (N_13037,N_7315,N_7979);
or U13038 (N_13038,N_6499,N_6073);
nand U13039 (N_13039,N_9788,N_5405);
nand U13040 (N_13040,N_9230,N_6260);
nand U13041 (N_13041,N_5857,N_9800);
nor U13042 (N_13042,N_6607,N_7481);
nor U13043 (N_13043,N_6247,N_5972);
nor U13044 (N_13044,N_7421,N_6080);
nand U13045 (N_13045,N_5493,N_6839);
xor U13046 (N_13046,N_6536,N_5899);
xnor U13047 (N_13047,N_9105,N_6605);
and U13048 (N_13048,N_5678,N_7615);
xor U13049 (N_13049,N_6274,N_5658);
nand U13050 (N_13050,N_8120,N_7818);
nand U13051 (N_13051,N_6853,N_7369);
nor U13052 (N_13052,N_8592,N_6330);
or U13053 (N_13053,N_6793,N_9459);
nor U13054 (N_13054,N_5813,N_7412);
nand U13055 (N_13055,N_5952,N_5457);
and U13056 (N_13056,N_8726,N_8210);
xor U13057 (N_13057,N_8056,N_7001);
xor U13058 (N_13058,N_7758,N_5442);
or U13059 (N_13059,N_7455,N_7439);
and U13060 (N_13060,N_8143,N_8217);
and U13061 (N_13061,N_6350,N_6086);
nand U13062 (N_13062,N_6224,N_5953);
xnor U13063 (N_13063,N_5194,N_7001);
and U13064 (N_13064,N_8875,N_8293);
nand U13065 (N_13065,N_8476,N_5050);
nor U13066 (N_13066,N_8649,N_9353);
xnor U13067 (N_13067,N_6804,N_5681);
nand U13068 (N_13068,N_6227,N_7984);
and U13069 (N_13069,N_8584,N_7322);
or U13070 (N_13070,N_9091,N_6384);
xor U13071 (N_13071,N_7685,N_9108);
nor U13072 (N_13072,N_7454,N_6169);
nand U13073 (N_13073,N_9496,N_6529);
nor U13074 (N_13074,N_5565,N_5395);
and U13075 (N_13075,N_9540,N_9847);
or U13076 (N_13076,N_8631,N_6908);
nor U13077 (N_13077,N_7880,N_9693);
or U13078 (N_13078,N_8940,N_9458);
nand U13079 (N_13079,N_6211,N_8750);
nand U13080 (N_13080,N_9691,N_7564);
or U13081 (N_13081,N_6994,N_9323);
nor U13082 (N_13082,N_9750,N_8366);
or U13083 (N_13083,N_7384,N_6072);
and U13084 (N_13084,N_7157,N_8189);
xor U13085 (N_13085,N_5868,N_6290);
nor U13086 (N_13086,N_9098,N_7574);
nand U13087 (N_13087,N_5608,N_7932);
nor U13088 (N_13088,N_8943,N_6577);
nor U13089 (N_13089,N_9311,N_6157);
nand U13090 (N_13090,N_5534,N_5761);
and U13091 (N_13091,N_5652,N_8667);
or U13092 (N_13092,N_8595,N_7645);
and U13093 (N_13093,N_5785,N_7925);
xor U13094 (N_13094,N_5242,N_8935);
xor U13095 (N_13095,N_9361,N_9443);
nand U13096 (N_13096,N_9102,N_6248);
or U13097 (N_13097,N_7177,N_9204);
xnor U13098 (N_13098,N_9008,N_6218);
nand U13099 (N_13099,N_5435,N_5347);
or U13100 (N_13100,N_8420,N_5142);
nand U13101 (N_13101,N_9804,N_8866);
nand U13102 (N_13102,N_7682,N_9049);
xor U13103 (N_13103,N_5494,N_7526);
nor U13104 (N_13104,N_9686,N_6618);
nor U13105 (N_13105,N_8323,N_7727);
or U13106 (N_13106,N_6431,N_5606);
or U13107 (N_13107,N_7036,N_7350);
xor U13108 (N_13108,N_8585,N_9576);
nor U13109 (N_13109,N_9750,N_6921);
and U13110 (N_13110,N_8251,N_7010);
xor U13111 (N_13111,N_9891,N_7110);
nand U13112 (N_13112,N_8628,N_5355);
and U13113 (N_13113,N_9061,N_8635);
and U13114 (N_13114,N_6484,N_6721);
nor U13115 (N_13115,N_8116,N_7335);
nor U13116 (N_13116,N_6992,N_8153);
or U13117 (N_13117,N_5495,N_7522);
xnor U13118 (N_13118,N_6367,N_7233);
nor U13119 (N_13119,N_7953,N_8495);
nand U13120 (N_13120,N_8970,N_6355);
and U13121 (N_13121,N_7055,N_7217);
or U13122 (N_13122,N_8181,N_9928);
nor U13123 (N_13123,N_9457,N_5774);
and U13124 (N_13124,N_6499,N_6096);
nor U13125 (N_13125,N_6632,N_8155);
nor U13126 (N_13126,N_7124,N_9416);
and U13127 (N_13127,N_7641,N_7800);
or U13128 (N_13128,N_7855,N_5705);
xnor U13129 (N_13129,N_5456,N_5539);
nor U13130 (N_13130,N_6468,N_8697);
or U13131 (N_13131,N_6467,N_6698);
xor U13132 (N_13132,N_5892,N_8335);
nor U13133 (N_13133,N_5690,N_9823);
xor U13134 (N_13134,N_5385,N_6348);
or U13135 (N_13135,N_5597,N_5747);
xor U13136 (N_13136,N_6108,N_6627);
nand U13137 (N_13137,N_8086,N_6425);
nor U13138 (N_13138,N_8646,N_9077);
xor U13139 (N_13139,N_8188,N_7857);
nand U13140 (N_13140,N_9534,N_8021);
and U13141 (N_13141,N_6208,N_7180);
nor U13142 (N_13142,N_6423,N_6584);
and U13143 (N_13143,N_5329,N_5642);
or U13144 (N_13144,N_7790,N_8714);
xnor U13145 (N_13145,N_6169,N_5269);
and U13146 (N_13146,N_7183,N_7444);
nor U13147 (N_13147,N_8772,N_9637);
or U13148 (N_13148,N_8331,N_7533);
nor U13149 (N_13149,N_7008,N_8054);
nand U13150 (N_13150,N_6431,N_8827);
xor U13151 (N_13151,N_8628,N_5498);
and U13152 (N_13152,N_8100,N_6004);
xor U13153 (N_13153,N_7144,N_8302);
nand U13154 (N_13154,N_7879,N_6607);
nand U13155 (N_13155,N_5586,N_6535);
nor U13156 (N_13156,N_9632,N_5405);
nor U13157 (N_13157,N_7378,N_9798);
and U13158 (N_13158,N_8416,N_7498);
and U13159 (N_13159,N_8908,N_7259);
or U13160 (N_13160,N_5901,N_9004);
nor U13161 (N_13161,N_7356,N_5358);
and U13162 (N_13162,N_5650,N_9788);
xnor U13163 (N_13163,N_5738,N_7191);
or U13164 (N_13164,N_8575,N_6255);
or U13165 (N_13165,N_6970,N_7637);
and U13166 (N_13166,N_6941,N_5279);
and U13167 (N_13167,N_7257,N_7868);
nand U13168 (N_13168,N_7222,N_6877);
nand U13169 (N_13169,N_8569,N_7707);
nand U13170 (N_13170,N_8873,N_6881);
and U13171 (N_13171,N_5065,N_8978);
and U13172 (N_13172,N_5420,N_8793);
or U13173 (N_13173,N_5450,N_5904);
nand U13174 (N_13174,N_5322,N_7894);
xor U13175 (N_13175,N_6773,N_5559);
xor U13176 (N_13176,N_8577,N_5998);
or U13177 (N_13177,N_9490,N_6433);
and U13178 (N_13178,N_8915,N_7120);
and U13179 (N_13179,N_7740,N_8328);
or U13180 (N_13180,N_5503,N_5519);
xnor U13181 (N_13181,N_8117,N_8883);
nor U13182 (N_13182,N_5999,N_8481);
nand U13183 (N_13183,N_7846,N_9907);
nand U13184 (N_13184,N_5247,N_7748);
xor U13185 (N_13185,N_9808,N_6286);
or U13186 (N_13186,N_5946,N_6696);
nor U13187 (N_13187,N_7643,N_8133);
nand U13188 (N_13188,N_5080,N_6097);
and U13189 (N_13189,N_7436,N_9484);
nor U13190 (N_13190,N_9787,N_7385);
nor U13191 (N_13191,N_5163,N_5406);
xor U13192 (N_13192,N_9956,N_8547);
xnor U13193 (N_13193,N_7503,N_7533);
nand U13194 (N_13194,N_9239,N_6578);
nand U13195 (N_13195,N_8224,N_5629);
nor U13196 (N_13196,N_7215,N_7584);
nand U13197 (N_13197,N_6355,N_8709);
nor U13198 (N_13198,N_9108,N_5960);
or U13199 (N_13199,N_7830,N_6578);
and U13200 (N_13200,N_6993,N_7122);
nand U13201 (N_13201,N_6077,N_9623);
xnor U13202 (N_13202,N_9312,N_6944);
nor U13203 (N_13203,N_7137,N_8718);
or U13204 (N_13204,N_5155,N_8323);
nand U13205 (N_13205,N_7642,N_5424);
xor U13206 (N_13206,N_8096,N_8751);
nand U13207 (N_13207,N_7139,N_8694);
nor U13208 (N_13208,N_8347,N_8684);
xnor U13209 (N_13209,N_7174,N_6372);
or U13210 (N_13210,N_7977,N_8946);
xnor U13211 (N_13211,N_7850,N_5704);
or U13212 (N_13212,N_9455,N_9410);
nand U13213 (N_13213,N_8629,N_5447);
or U13214 (N_13214,N_7511,N_7785);
or U13215 (N_13215,N_7071,N_9091);
or U13216 (N_13216,N_6179,N_5773);
nor U13217 (N_13217,N_8937,N_6249);
nand U13218 (N_13218,N_9978,N_6959);
xor U13219 (N_13219,N_8633,N_7641);
nand U13220 (N_13220,N_6529,N_5873);
or U13221 (N_13221,N_5964,N_5977);
nor U13222 (N_13222,N_9544,N_9566);
xnor U13223 (N_13223,N_7378,N_6189);
or U13224 (N_13224,N_6985,N_5156);
xnor U13225 (N_13225,N_5101,N_7795);
xor U13226 (N_13226,N_5212,N_9026);
or U13227 (N_13227,N_9902,N_6983);
and U13228 (N_13228,N_5509,N_9553);
and U13229 (N_13229,N_7163,N_6974);
or U13230 (N_13230,N_7976,N_7985);
nand U13231 (N_13231,N_7839,N_6485);
and U13232 (N_13232,N_7745,N_5065);
and U13233 (N_13233,N_6867,N_7716);
nor U13234 (N_13234,N_9487,N_7832);
xor U13235 (N_13235,N_6983,N_9433);
or U13236 (N_13236,N_9010,N_9714);
nor U13237 (N_13237,N_7178,N_6493);
and U13238 (N_13238,N_6987,N_5975);
nor U13239 (N_13239,N_5637,N_6958);
nor U13240 (N_13240,N_8714,N_7159);
xor U13241 (N_13241,N_8562,N_8244);
nand U13242 (N_13242,N_5755,N_5951);
or U13243 (N_13243,N_8838,N_6713);
nor U13244 (N_13244,N_6410,N_6677);
nor U13245 (N_13245,N_5222,N_7627);
and U13246 (N_13246,N_7849,N_8359);
or U13247 (N_13247,N_6490,N_9443);
xor U13248 (N_13248,N_7092,N_8623);
and U13249 (N_13249,N_5682,N_7308);
xnor U13250 (N_13250,N_9992,N_7141);
nor U13251 (N_13251,N_7513,N_7307);
or U13252 (N_13252,N_9808,N_9385);
or U13253 (N_13253,N_8940,N_9304);
xor U13254 (N_13254,N_7490,N_8982);
and U13255 (N_13255,N_8215,N_5110);
or U13256 (N_13256,N_5730,N_6179);
xnor U13257 (N_13257,N_8158,N_5714);
or U13258 (N_13258,N_8222,N_7380);
or U13259 (N_13259,N_9328,N_6375);
nand U13260 (N_13260,N_5040,N_5643);
xnor U13261 (N_13261,N_6785,N_9200);
nor U13262 (N_13262,N_6938,N_7393);
or U13263 (N_13263,N_8825,N_8762);
or U13264 (N_13264,N_5753,N_5565);
nand U13265 (N_13265,N_8135,N_8766);
or U13266 (N_13266,N_7331,N_8756);
or U13267 (N_13267,N_7366,N_9565);
nor U13268 (N_13268,N_8289,N_6056);
nor U13269 (N_13269,N_6845,N_9183);
or U13270 (N_13270,N_8643,N_9750);
xor U13271 (N_13271,N_6355,N_6277);
nor U13272 (N_13272,N_5925,N_9482);
xnor U13273 (N_13273,N_5682,N_7844);
xor U13274 (N_13274,N_9260,N_6796);
and U13275 (N_13275,N_8409,N_6361);
or U13276 (N_13276,N_6647,N_6059);
or U13277 (N_13277,N_5570,N_6194);
xnor U13278 (N_13278,N_8312,N_5028);
and U13279 (N_13279,N_7372,N_5757);
or U13280 (N_13280,N_9632,N_7982);
and U13281 (N_13281,N_6030,N_7257);
nand U13282 (N_13282,N_8157,N_5771);
and U13283 (N_13283,N_7449,N_9105);
and U13284 (N_13284,N_6926,N_8390);
and U13285 (N_13285,N_8833,N_7963);
nor U13286 (N_13286,N_7789,N_8254);
and U13287 (N_13287,N_5791,N_5227);
xor U13288 (N_13288,N_7243,N_8015);
xor U13289 (N_13289,N_8843,N_7920);
xnor U13290 (N_13290,N_5750,N_6030);
nand U13291 (N_13291,N_5220,N_8218);
nand U13292 (N_13292,N_8032,N_6099);
nand U13293 (N_13293,N_6078,N_9836);
or U13294 (N_13294,N_8381,N_7933);
and U13295 (N_13295,N_7509,N_5485);
xnor U13296 (N_13296,N_8745,N_7883);
nor U13297 (N_13297,N_5799,N_8040);
or U13298 (N_13298,N_9210,N_9163);
nor U13299 (N_13299,N_9584,N_7495);
nor U13300 (N_13300,N_8526,N_9894);
or U13301 (N_13301,N_9671,N_9440);
nand U13302 (N_13302,N_9304,N_9176);
nor U13303 (N_13303,N_5191,N_6237);
and U13304 (N_13304,N_8394,N_9913);
or U13305 (N_13305,N_5383,N_5827);
nand U13306 (N_13306,N_5323,N_7831);
xor U13307 (N_13307,N_5019,N_9094);
nand U13308 (N_13308,N_7143,N_6725);
or U13309 (N_13309,N_6620,N_9390);
xor U13310 (N_13310,N_9743,N_9878);
and U13311 (N_13311,N_6944,N_6241);
nand U13312 (N_13312,N_8251,N_6413);
and U13313 (N_13313,N_9366,N_7011);
and U13314 (N_13314,N_6486,N_8525);
nand U13315 (N_13315,N_9619,N_9922);
nor U13316 (N_13316,N_9634,N_5506);
nor U13317 (N_13317,N_6034,N_6411);
or U13318 (N_13318,N_5742,N_6715);
or U13319 (N_13319,N_7402,N_8411);
nor U13320 (N_13320,N_7998,N_9603);
nor U13321 (N_13321,N_6069,N_7535);
xor U13322 (N_13322,N_6195,N_7946);
nor U13323 (N_13323,N_9638,N_8304);
nand U13324 (N_13324,N_6718,N_5206);
nand U13325 (N_13325,N_5495,N_7218);
nor U13326 (N_13326,N_5116,N_9818);
nand U13327 (N_13327,N_7004,N_9474);
xnor U13328 (N_13328,N_5568,N_8205);
nand U13329 (N_13329,N_9660,N_9360);
xnor U13330 (N_13330,N_9361,N_7518);
xnor U13331 (N_13331,N_9274,N_9684);
nor U13332 (N_13332,N_7744,N_8611);
or U13333 (N_13333,N_9143,N_5910);
nand U13334 (N_13334,N_5032,N_8326);
nand U13335 (N_13335,N_8289,N_7821);
xor U13336 (N_13336,N_7280,N_7089);
nor U13337 (N_13337,N_6799,N_9237);
or U13338 (N_13338,N_8194,N_6282);
nand U13339 (N_13339,N_6483,N_6568);
nor U13340 (N_13340,N_8738,N_5960);
nor U13341 (N_13341,N_8437,N_8156);
xor U13342 (N_13342,N_8991,N_8472);
nor U13343 (N_13343,N_7369,N_7221);
xor U13344 (N_13344,N_6668,N_5947);
nor U13345 (N_13345,N_8070,N_5472);
nand U13346 (N_13346,N_8100,N_6100);
nand U13347 (N_13347,N_6736,N_9058);
xor U13348 (N_13348,N_5108,N_9729);
nor U13349 (N_13349,N_7565,N_5950);
and U13350 (N_13350,N_6167,N_9206);
and U13351 (N_13351,N_7394,N_9802);
and U13352 (N_13352,N_5503,N_8163);
xor U13353 (N_13353,N_9830,N_6142);
nand U13354 (N_13354,N_9413,N_9516);
xor U13355 (N_13355,N_5895,N_5959);
nand U13356 (N_13356,N_5447,N_8614);
and U13357 (N_13357,N_6283,N_7515);
xor U13358 (N_13358,N_5128,N_8672);
or U13359 (N_13359,N_7098,N_6819);
nor U13360 (N_13360,N_6092,N_7563);
or U13361 (N_13361,N_7838,N_7496);
xor U13362 (N_13362,N_7366,N_9666);
or U13363 (N_13363,N_6628,N_9177);
or U13364 (N_13364,N_9954,N_5113);
xor U13365 (N_13365,N_8726,N_6678);
or U13366 (N_13366,N_5721,N_7623);
or U13367 (N_13367,N_9198,N_9919);
nor U13368 (N_13368,N_8737,N_6285);
xnor U13369 (N_13369,N_9228,N_5827);
or U13370 (N_13370,N_7650,N_7856);
and U13371 (N_13371,N_8142,N_6386);
nor U13372 (N_13372,N_8181,N_5176);
or U13373 (N_13373,N_7213,N_7742);
and U13374 (N_13374,N_9514,N_7444);
nand U13375 (N_13375,N_8987,N_5850);
nand U13376 (N_13376,N_8917,N_7394);
or U13377 (N_13377,N_6130,N_8518);
xnor U13378 (N_13378,N_8703,N_9640);
xnor U13379 (N_13379,N_6425,N_6898);
xnor U13380 (N_13380,N_5099,N_5692);
nor U13381 (N_13381,N_5994,N_9331);
xnor U13382 (N_13382,N_7171,N_6981);
nor U13383 (N_13383,N_8966,N_7611);
or U13384 (N_13384,N_8582,N_7175);
and U13385 (N_13385,N_6575,N_9774);
or U13386 (N_13386,N_6303,N_9519);
and U13387 (N_13387,N_9210,N_7288);
nand U13388 (N_13388,N_9125,N_6954);
nor U13389 (N_13389,N_9102,N_5587);
nor U13390 (N_13390,N_9549,N_8536);
xor U13391 (N_13391,N_7216,N_5296);
xnor U13392 (N_13392,N_6526,N_7887);
nand U13393 (N_13393,N_6542,N_5292);
and U13394 (N_13394,N_6487,N_9393);
nand U13395 (N_13395,N_9160,N_5610);
xor U13396 (N_13396,N_9699,N_6559);
nand U13397 (N_13397,N_5166,N_7346);
or U13398 (N_13398,N_7784,N_6544);
and U13399 (N_13399,N_7343,N_7874);
xor U13400 (N_13400,N_7319,N_9224);
and U13401 (N_13401,N_8385,N_5885);
nand U13402 (N_13402,N_9072,N_6426);
xnor U13403 (N_13403,N_7407,N_7821);
or U13404 (N_13404,N_6369,N_7985);
and U13405 (N_13405,N_8130,N_7427);
and U13406 (N_13406,N_9668,N_5377);
nor U13407 (N_13407,N_8640,N_5877);
xor U13408 (N_13408,N_6710,N_5093);
nand U13409 (N_13409,N_5764,N_5784);
and U13410 (N_13410,N_5025,N_8782);
or U13411 (N_13411,N_7478,N_8721);
xor U13412 (N_13412,N_8785,N_8796);
nand U13413 (N_13413,N_6214,N_7451);
nand U13414 (N_13414,N_5698,N_8756);
or U13415 (N_13415,N_7431,N_5452);
xor U13416 (N_13416,N_8559,N_9854);
nor U13417 (N_13417,N_6067,N_7498);
nor U13418 (N_13418,N_6694,N_9314);
and U13419 (N_13419,N_5595,N_5141);
nor U13420 (N_13420,N_5602,N_8281);
xor U13421 (N_13421,N_6207,N_9667);
and U13422 (N_13422,N_9841,N_5759);
xnor U13423 (N_13423,N_8355,N_5612);
or U13424 (N_13424,N_9592,N_8029);
nor U13425 (N_13425,N_6928,N_5777);
nor U13426 (N_13426,N_9835,N_8668);
nor U13427 (N_13427,N_8210,N_8067);
and U13428 (N_13428,N_9612,N_5634);
nor U13429 (N_13429,N_7621,N_9971);
nor U13430 (N_13430,N_9920,N_6993);
or U13431 (N_13431,N_8051,N_9832);
nand U13432 (N_13432,N_5481,N_5410);
xnor U13433 (N_13433,N_8936,N_9885);
or U13434 (N_13434,N_6287,N_9543);
xor U13435 (N_13435,N_9562,N_5718);
xor U13436 (N_13436,N_5078,N_5927);
nand U13437 (N_13437,N_6894,N_8690);
xor U13438 (N_13438,N_9897,N_5068);
nor U13439 (N_13439,N_6989,N_8091);
xor U13440 (N_13440,N_7354,N_9443);
nand U13441 (N_13441,N_5416,N_7605);
nand U13442 (N_13442,N_8314,N_7767);
nand U13443 (N_13443,N_5372,N_7539);
and U13444 (N_13444,N_9315,N_5763);
nor U13445 (N_13445,N_9110,N_7853);
nor U13446 (N_13446,N_6683,N_9806);
nor U13447 (N_13447,N_6724,N_8409);
or U13448 (N_13448,N_6983,N_7931);
nand U13449 (N_13449,N_7095,N_5414);
or U13450 (N_13450,N_8056,N_9550);
and U13451 (N_13451,N_7576,N_6997);
nand U13452 (N_13452,N_9836,N_8787);
nor U13453 (N_13453,N_8464,N_5346);
nor U13454 (N_13454,N_7174,N_5838);
and U13455 (N_13455,N_6304,N_6330);
nor U13456 (N_13456,N_7851,N_5336);
nor U13457 (N_13457,N_6876,N_5443);
or U13458 (N_13458,N_9310,N_9047);
nand U13459 (N_13459,N_6576,N_9703);
and U13460 (N_13460,N_9761,N_8935);
nor U13461 (N_13461,N_9908,N_9705);
nand U13462 (N_13462,N_5450,N_5955);
xor U13463 (N_13463,N_9062,N_5300);
nor U13464 (N_13464,N_9076,N_9513);
nor U13465 (N_13465,N_8568,N_8628);
and U13466 (N_13466,N_9883,N_6718);
or U13467 (N_13467,N_7954,N_6105);
or U13468 (N_13468,N_9798,N_7050);
nor U13469 (N_13469,N_9644,N_5513);
nand U13470 (N_13470,N_5195,N_8620);
nor U13471 (N_13471,N_9698,N_7881);
or U13472 (N_13472,N_5121,N_6450);
nor U13473 (N_13473,N_7991,N_7872);
xor U13474 (N_13474,N_6788,N_7959);
xnor U13475 (N_13475,N_7617,N_7464);
xor U13476 (N_13476,N_8775,N_6505);
nor U13477 (N_13477,N_7371,N_8279);
and U13478 (N_13478,N_6638,N_5030);
nor U13479 (N_13479,N_9800,N_9807);
xnor U13480 (N_13480,N_7452,N_8952);
nor U13481 (N_13481,N_6727,N_8242);
nand U13482 (N_13482,N_7857,N_7020);
xor U13483 (N_13483,N_9422,N_5510);
and U13484 (N_13484,N_8336,N_5149);
nor U13485 (N_13485,N_9082,N_9479);
or U13486 (N_13486,N_9546,N_7190);
nand U13487 (N_13487,N_8586,N_7209);
nand U13488 (N_13488,N_6215,N_9482);
or U13489 (N_13489,N_9050,N_5381);
nor U13490 (N_13490,N_8582,N_8133);
xnor U13491 (N_13491,N_8446,N_7907);
or U13492 (N_13492,N_8104,N_8200);
nand U13493 (N_13493,N_8339,N_7684);
nor U13494 (N_13494,N_5328,N_8717);
xor U13495 (N_13495,N_8941,N_6202);
and U13496 (N_13496,N_8770,N_8743);
and U13497 (N_13497,N_7190,N_6513);
and U13498 (N_13498,N_6854,N_8904);
xor U13499 (N_13499,N_6321,N_7821);
nor U13500 (N_13500,N_5840,N_8049);
nand U13501 (N_13501,N_7715,N_9092);
and U13502 (N_13502,N_8991,N_7287);
nor U13503 (N_13503,N_7189,N_7877);
xnor U13504 (N_13504,N_7552,N_9150);
xnor U13505 (N_13505,N_6837,N_5229);
nor U13506 (N_13506,N_5631,N_5872);
and U13507 (N_13507,N_7493,N_5312);
nor U13508 (N_13508,N_8566,N_6520);
nor U13509 (N_13509,N_6126,N_8632);
nand U13510 (N_13510,N_9249,N_6736);
and U13511 (N_13511,N_8286,N_5402);
or U13512 (N_13512,N_9888,N_6319);
nor U13513 (N_13513,N_5210,N_8932);
nor U13514 (N_13514,N_8386,N_9742);
nand U13515 (N_13515,N_5310,N_8388);
and U13516 (N_13516,N_6500,N_8941);
or U13517 (N_13517,N_8212,N_8747);
xnor U13518 (N_13518,N_9584,N_7523);
xnor U13519 (N_13519,N_8811,N_7195);
or U13520 (N_13520,N_7184,N_9037);
nand U13521 (N_13521,N_8583,N_7189);
and U13522 (N_13522,N_7529,N_9502);
or U13523 (N_13523,N_8717,N_7171);
and U13524 (N_13524,N_5804,N_6586);
and U13525 (N_13525,N_7181,N_8326);
xor U13526 (N_13526,N_8737,N_8405);
nor U13527 (N_13527,N_5820,N_8876);
or U13528 (N_13528,N_7997,N_9230);
nor U13529 (N_13529,N_5614,N_5735);
nand U13530 (N_13530,N_7435,N_9343);
and U13531 (N_13531,N_8105,N_7163);
nand U13532 (N_13532,N_8538,N_8747);
nor U13533 (N_13533,N_6873,N_9306);
xnor U13534 (N_13534,N_8070,N_8335);
nand U13535 (N_13535,N_7080,N_5347);
or U13536 (N_13536,N_8974,N_8510);
nand U13537 (N_13537,N_5125,N_9365);
xnor U13538 (N_13538,N_8402,N_8011);
or U13539 (N_13539,N_8336,N_8151);
or U13540 (N_13540,N_9470,N_8201);
or U13541 (N_13541,N_5866,N_8115);
and U13542 (N_13542,N_5571,N_7194);
xnor U13543 (N_13543,N_6903,N_8778);
nand U13544 (N_13544,N_7601,N_5570);
and U13545 (N_13545,N_9075,N_8485);
nand U13546 (N_13546,N_8393,N_5775);
and U13547 (N_13547,N_9896,N_6510);
nor U13548 (N_13548,N_5698,N_8864);
nand U13549 (N_13549,N_6887,N_7496);
xor U13550 (N_13550,N_7379,N_7896);
and U13551 (N_13551,N_8433,N_7325);
or U13552 (N_13552,N_7655,N_8918);
or U13553 (N_13553,N_8846,N_8820);
or U13554 (N_13554,N_9521,N_7587);
and U13555 (N_13555,N_6651,N_5994);
nand U13556 (N_13556,N_8144,N_5136);
xor U13557 (N_13557,N_6457,N_5167);
nand U13558 (N_13558,N_5730,N_9479);
nor U13559 (N_13559,N_9950,N_5883);
nor U13560 (N_13560,N_6050,N_5609);
nand U13561 (N_13561,N_8555,N_7604);
xor U13562 (N_13562,N_5647,N_9964);
xor U13563 (N_13563,N_5624,N_9761);
nand U13564 (N_13564,N_6959,N_5800);
or U13565 (N_13565,N_8740,N_9711);
nand U13566 (N_13566,N_7144,N_5994);
xor U13567 (N_13567,N_8357,N_8303);
or U13568 (N_13568,N_8731,N_7858);
nand U13569 (N_13569,N_6758,N_6584);
xnor U13570 (N_13570,N_5059,N_6310);
xnor U13571 (N_13571,N_9813,N_9942);
and U13572 (N_13572,N_7301,N_5023);
or U13573 (N_13573,N_8153,N_7468);
xor U13574 (N_13574,N_9755,N_7250);
and U13575 (N_13575,N_8186,N_8500);
nor U13576 (N_13576,N_7549,N_9479);
nand U13577 (N_13577,N_5816,N_7118);
nor U13578 (N_13578,N_9164,N_5175);
or U13579 (N_13579,N_8961,N_6355);
xnor U13580 (N_13580,N_8855,N_6437);
xnor U13581 (N_13581,N_7261,N_5226);
and U13582 (N_13582,N_7007,N_6780);
xnor U13583 (N_13583,N_8994,N_7175);
or U13584 (N_13584,N_7822,N_9576);
nand U13585 (N_13585,N_7227,N_6115);
or U13586 (N_13586,N_9271,N_7522);
xnor U13587 (N_13587,N_9084,N_8612);
and U13588 (N_13588,N_5328,N_5330);
and U13589 (N_13589,N_6652,N_6374);
or U13590 (N_13590,N_7185,N_9063);
xor U13591 (N_13591,N_7376,N_8798);
and U13592 (N_13592,N_5600,N_8188);
or U13593 (N_13593,N_6302,N_5918);
nand U13594 (N_13594,N_9991,N_7146);
nand U13595 (N_13595,N_7024,N_5793);
or U13596 (N_13596,N_5344,N_5533);
nor U13597 (N_13597,N_7979,N_5454);
xor U13598 (N_13598,N_5982,N_8989);
or U13599 (N_13599,N_8669,N_8874);
and U13600 (N_13600,N_6549,N_5455);
xor U13601 (N_13601,N_8162,N_8042);
and U13602 (N_13602,N_9993,N_8459);
nand U13603 (N_13603,N_5736,N_9061);
nand U13604 (N_13604,N_9227,N_6717);
or U13605 (N_13605,N_9842,N_8183);
or U13606 (N_13606,N_6072,N_7280);
or U13607 (N_13607,N_5528,N_5202);
and U13608 (N_13608,N_9129,N_9641);
nand U13609 (N_13609,N_6099,N_5765);
nand U13610 (N_13610,N_9098,N_9620);
nand U13611 (N_13611,N_7758,N_9952);
and U13612 (N_13612,N_9425,N_5655);
nor U13613 (N_13613,N_9916,N_7572);
nand U13614 (N_13614,N_5234,N_8209);
and U13615 (N_13615,N_9294,N_6301);
nor U13616 (N_13616,N_8304,N_6409);
nor U13617 (N_13617,N_5462,N_7765);
or U13618 (N_13618,N_5176,N_9750);
or U13619 (N_13619,N_5532,N_8194);
nand U13620 (N_13620,N_9997,N_7378);
nor U13621 (N_13621,N_9704,N_5980);
and U13622 (N_13622,N_6998,N_6226);
xor U13623 (N_13623,N_6081,N_8855);
and U13624 (N_13624,N_7358,N_6746);
nand U13625 (N_13625,N_6922,N_8439);
nor U13626 (N_13626,N_8842,N_7086);
xnor U13627 (N_13627,N_5361,N_7629);
xor U13628 (N_13628,N_5121,N_7436);
xnor U13629 (N_13629,N_9475,N_9806);
xnor U13630 (N_13630,N_9924,N_7559);
nand U13631 (N_13631,N_7109,N_5107);
nand U13632 (N_13632,N_8295,N_8160);
xnor U13633 (N_13633,N_8671,N_7391);
nand U13634 (N_13634,N_5762,N_5718);
xor U13635 (N_13635,N_7000,N_8734);
xor U13636 (N_13636,N_6982,N_5846);
xnor U13637 (N_13637,N_7564,N_6245);
and U13638 (N_13638,N_7996,N_9123);
xor U13639 (N_13639,N_5791,N_8891);
nor U13640 (N_13640,N_8310,N_8983);
nand U13641 (N_13641,N_6285,N_6144);
nand U13642 (N_13642,N_6966,N_8309);
xnor U13643 (N_13643,N_6548,N_7352);
nand U13644 (N_13644,N_7871,N_6920);
nand U13645 (N_13645,N_6612,N_5683);
or U13646 (N_13646,N_7323,N_8304);
xor U13647 (N_13647,N_7051,N_7303);
or U13648 (N_13648,N_9870,N_9936);
xor U13649 (N_13649,N_6250,N_8210);
or U13650 (N_13650,N_5544,N_9875);
and U13651 (N_13651,N_7150,N_6126);
or U13652 (N_13652,N_8979,N_9641);
nor U13653 (N_13653,N_7278,N_8390);
and U13654 (N_13654,N_8234,N_8842);
xnor U13655 (N_13655,N_5924,N_7749);
xor U13656 (N_13656,N_8061,N_5029);
or U13657 (N_13657,N_8490,N_5096);
nand U13658 (N_13658,N_6436,N_5534);
nand U13659 (N_13659,N_5718,N_9343);
or U13660 (N_13660,N_6542,N_6850);
nor U13661 (N_13661,N_9046,N_5836);
xnor U13662 (N_13662,N_9151,N_9056);
xor U13663 (N_13663,N_5211,N_5330);
xor U13664 (N_13664,N_8086,N_6370);
xnor U13665 (N_13665,N_5272,N_9542);
and U13666 (N_13666,N_9779,N_8047);
or U13667 (N_13667,N_7649,N_8060);
nor U13668 (N_13668,N_9158,N_7548);
nand U13669 (N_13669,N_7116,N_8431);
or U13670 (N_13670,N_8529,N_7344);
xnor U13671 (N_13671,N_9870,N_5121);
and U13672 (N_13672,N_8435,N_8198);
nand U13673 (N_13673,N_5433,N_8972);
nand U13674 (N_13674,N_7124,N_6629);
nand U13675 (N_13675,N_6787,N_7207);
xnor U13676 (N_13676,N_8756,N_6083);
xnor U13677 (N_13677,N_6483,N_8547);
nor U13678 (N_13678,N_6848,N_5841);
nor U13679 (N_13679,N_9124,N_9665);
and U13680 (N_13680,N_6095,N_6917);
nor U13681 (N_13681,N_6884,N_7686);
xor U13682 (N_13682,N_7200,N_5858);
and U13683 (N_13683,N_9739,N_7824);
nor U13684 (N_13684,N_6945,N_9916);
xnor U13685 (N_13685,N_7312,N_6146);
xor U13686 (N_13686,N_8659,N_5850);
or U13687 (N_13687,N_8403,N_6901);
or U13688 (N_13688,N_7878,N_7592);
and U13689 (N_13689,N_9303,N_7664);
nand U13690 (N_13690,N_8784,N_5045);
xor U13691 (N_13691,N_8577,N_8785);
nand U13692 (N_13692,N_9231,N_9954);
and U13693 (N_13693,N_9446,N_8805);
or U13694 (N_13694,N_5075,N_9722);
and U13695 (N_13695,N_8811,N_8640);
and U13696 (N_13696,N_8651,N_6584);
or U13697 (N_13697,N_6057,N_5419);
and U13698 (N_13698,N_6878,N_6961);
nor U13699 (N_13699,N_9407,N_5803);
xor U13700 (N_13700,N_7973,N_6672);
nand U13701 (N_13701,N_6107,N_6120);
nor U13702 (N_13702,N_5219,N_9884);
xnor U13703 (N_13703,N_7063,N_5443);
nand U13704 (N_13704,N_5444,N_7253);
and U13705 (N_13705,N_8311,N_7033);
xnor U13706 (N_13706,N_9205,N_8914);
or U13707 (N_13707,N_9871,N_5711);
and U13708 (N_13708,N_8229,N_8809);
and U13709 (N_13709,N_6182,N_9237);
nor U13710 (N_13710,N_9424,N_9121);
xor U13711 (N_13711,N_5393,N_7416);
nand U13712 (N_13712,N_7356,N_8978);
or U13713 (N_13713,N_6743,N_6149);
and U13714 (N_13714,N_6438,N_7496);
xnor U13715 (N_13715,N_8544,N_8909);
nor U13716 (N_13716,N_8342,N_7692);
xnor U13717 (N_13717,N_5256,N_8653);
nor U13718 (N_13718,N_8404,N_9196);
and U13719 (N_13719,N_8755,N_6285);
or U13720 (N_13720,N_7421,N_6560);
xnor U13721 (N_13721,N_5215,N_6557);
xor U13722 (N_13722,N_6754,N_7162);
or U13723 (N_13723,N_9039,N_9398);
and U13724 (N_13724,N_7023,N_9868);
nor U13725 (N_13725,N_8007,N_8491);
xor U13726 (N_13726,N_7914,N_6220);
xor U13727 (N_13727,N_6017,N_8136);
xnor U13728 (N_13728,N_8194,N_5388);
and U13729 (N_13729,N_5359,N_6787);
or U13730 (N_13730,N_7667,N_5769);
xor U13731 (N_13731,N_8181,N_9420);
nand U13732 (N_13732,N_6109,N_9062);
nor U13733 (N_13733,N_6681,N_6817);
nor U13734 (N_13734,N_6065,N_9864);
nor U13735 (N_13735,N_6374,N_9274);
xnor U13736 (N_13736,N_9391,N_9273);
and U13737 (N_13737,N_5184,N_8198);
nor U13738 (N_13738,N_5988,N_7638);
xor U13739 (N_13739,N_7663,N_7140);
xor U13740 (N_13740,N_5295,N_8970);
or U13741 (N_13741,N_6725,N_5247);
xor U13742 (N_13742,N_9658,N_7157);
nand U13743 (N_13743,N_8641,N_6056);
nand U13744 (N_13744,N_6159,N_9307);
or U13745 (N_13745,N_9401,N_8216);
nand U13746 (N_13746,N_8592,N_9013);
or U13747 (N_13747,N_5364,N_5970);
xor U13748 (N_13748,N_9998,N_9857);
and U13749 (N_13749,N_5385,N_7616);
nand U13750 (N_13750,N_8904,N_9975);
nand U13751 (N_13751,N_6383,N_8528);
and U13752 (N_13752,N_5625,N_9713);
nor U13753 (N_13753,N_8086,N_8376);
xor U13754 (N_13754,N_6444,N_7923);
nand U13755 (N_13755,N_9357,N_7009);
nor U13756 (N_13756,N_8587,N_8273);
xor U13757 (N_13757,N_5214,N_7874);
and U13758 (N_13758,N_7337,N_6781);
and U13759 (N_13759,N_9575,N_7445);
or U13760 (N_13760,N_6030,N_8128);
or U13761 (N_13761,N_7299,N_8666);
xor U13762 (N_13762,N_8172,N_9282);
nand U13763 (N_13763,N_7733,N_7181);
nand U13764 (N_13764,N_5489,N_9540);
or U13765 (N_13765,N_8446,N_6701);
nor U13766 (N_13766,N_8929,N_5022);
nor U13767 (N_13767,N_7514,N_7565);
nor U13768 (N_13768,N_8849,N_7013);
xor U13769 (N_13769,N_9503,N_8198);
nor U13770 (N_13770,N_7996,N_7061);
nand U13771 (N_13771,N_9903,N_7806);
and U13772 (N_13772,N_9332,N_9326);
and U13773 (N_13773,N_6116,N_6410);
and U13774 (N_13774,N_7785,N_9481);
or U13775 (N_13775,N_7357,N_6039);
nand U13776 (N_13776,N_6631,N_6268);
and U13777 (N_13777,N_9636,N_6702);
xor U13778 (N_13778,N_8472,N_6161);
or U13779 (N_13779,N_9384,N_9686);
nand U13780 (N_13780,N_5531,N_6727);
nand U13781 (N_13781,N_6541,N_8625);
xor U13782 (N_13782,N_5538,N_7662);
or U13783 (N_13783,N_8068,N_7414);
nand U13784 (N_13784,N_6032,N_7324);
nand U13785 (N_13785,N_7909,N_7676);
or U13786 (N_13786,N_5839,N_6541);
nand U13787 (N_13787,N_9994,N_9806);
and U13788 (N_13788,N_9855,N_6408);
and U13789 (N_13789,N_8676,N_7306);
xor U13790 (N_13790,N_6639,N_5382);
nand U13791 (N_13791,N_5305,N_6548);
xor U13792 (N_13792,N_6854,N_8152);
and U13793 (N_13793,N_7691,N_7957);
nand U13794 (N_13794,N_5292,N_9654);
nor U13795 (N_13795,N_9886,N_5683);
xor U13796 (N_13796,N_7113,N_5868);
xnor U13797 (N_13797,N_5174,N_6665);
or U13798 (N_13798,N_5949,N_6402);
and U13799 (N_13799,N_6020,N_6981);
nor U13800 (N_13800,N_8915,N_6762);
and U13801 (N_13801,N_6868,N_6780);
xor U13802 (N_13802,N_8388,N_9168);
or U13803 (N_13803,N_5550,N_6139);
xnor U13804 (N_13804,N_7251,N_5398);
and U13805 (N_13805,N_7853,N_9205);
or U13806 (N_13806,N_6537,N_7733);
or U13807 (N_13807,N_9003,N_6625);
and U13808 (N_13808,N_6467,N_9531);
and U13809 (N_13809,N_8428,N_5832);
xnor U13810 (N_13810,N_6877,N_7643);
and U13811 (N_13811,N_9615,N_9674);
nor U13812 (N_13812,N_9645,N_5715);
and U13813 (N_13813,N_5043,N_5308);
and U13814 (N_13814,N_5370,N_8025);
and U13815 (N_13815,N_7470,N_5412);
or U13816 (N_13816,N_5182,N_7841);
xnor U13817 (N_13817,N_6347,N_8520);
nand U13818 (N_13818,N_7869,N_5529);
or U13819 (N_13819,N_7128,N_6530);
xor U13820 (N_13820,N_5596,N_5944);
xor U13821 (N_13821,N_8977,N_8273);
nand U13822 (N_13822,N_9837,N_6688);
nor U13823 (N_13823,N_8295,N_6804);
nand U13824 (N_13824,N_7227,N_6525);
nor U13825 (N_13825,N_8760,N_7409);
nor U13826 (N_13826,N_7856,N_8332);
and U13827 (N_13827,N_9472,N_6652);
nor U13828 (N_13828,N_8519,N_5332);
and U13829 (N_13829,N_8147,N_7462);
and U13830 (N_13830,N_6806,N_7086);
nand U13831 (N_13831,N_5593,N_6731);
xor U13832 (N_13832,N_8041,N_6470);
nand U13833 (N_13833,N_5244,N_9945);
xor U13834 (N_13834,N_8516,N_8730);
xor U13835 (N_13835,N_8546,N_5969);
or U13836 (N_13836,N_9653,N_9637);
xnor U13837 (N_13837,N_6894,N_8513);
or U13838 (N_13838,N_5938,N_8262);
nand U13839 (N_13839,N_7603,N_9580);
nor U13840 (N_13840,N_8456,N_6893);
nor U13841 (N_13841,N_6197,N_6850);
nor U13842 (N_13842,N_7634,N_9778);
nand U13843 (N_13843,N_7940,N_5984);
nor U13844 (N_13844,N_5958,N_9235);
nor U13845 (N_13845,N_9735,N_7105);
or U13846 (N_13846,N_8655,N_5165);
or U13847 (N_13847,N_5755,N_6638);
nor U13848 (N_13848,N_5237,N_8413);
xnor U13849 (N_13849,N_8946,N_5267);
and U13850 (N_13850,N_6486,N_6062);
xor U13851 (N_13851,N_5806,N_7866);
nor U13852 (N_13852,N_5068,N_9882);
nand U13853 (N_13853,N_8159,N_7168);
or U13854 (N_13854,N_5103,N_9747);
or U13855 (N_13855,N_9383,N_7463);
or U13856 (N_13856,N_6788,N_8772);
xnor U13857 (N_13857,N_8777,N_5186);
nor U13858 (N_13858,N_5839,N_9657);
xnor U13859 (N_13859,N_5617,N_9224);
nor U13860 (N_13860,N_8468,N_9835);
nand U13861 (N_13861,N_7590,N_7172);
and U13862 (N_13862,N_9196,N_5115);
xnor U13863 (N_13863,N_9543,N_7684);
or U13864 (N_13864,N_8965,N_5540);
nor U13865 (N_13865,N_9378,N_8420);
nor U13866 (N_13866,N_7885,N_7759);
and U13867 (N_13867,N_6502,N_7309);
nand U13868 (N_13868,N_8327,N_8935);
or U13869 (N_13869,N_7249,N_7664);
or U13870 (N_13870,N_8700,N_9181);
and U13871 (N_13871,N_5264,N_9035);
nor U13872 (N_13872,N_7888,N_7653);
or U13873 (N_13873,N_6641,N_5697);
and U13874 (N_13874,N_8027,N_6942);
or U13875 (N_13875,N_5591,N_8020);
or U13876 (N_13876,N_8425,N_7513);
and U13877 (N_13877,N_9302,N_6160);
nor U13878 (N_13878,N_5390,N_8659);
nand U13879 (N_13879,N_9341,N_8296);
nand U13880 (N_13880,N_9693,N_6072);
or U13881 (N_13881,N_7546,N_7621);
and U13882 (N_13882,N_5749,N_5566);
and U13883 (N_13883,N_6509,N_5563);
and U13884 (N_13884,N_6831,N_8241);
nand U13885 (N_13885,N_6630,N_8728);
or U13886 (N_13886,N_7934,N_9623);
nor U13887 (N_13887,N_8878,N_6058);
xor U13888 (N_13888,N_6420,N_7183);
or U13889 (N_13889,N_8666,N_9247);
and U13890 (N_13890,N_7749,N_6593);
nor U13891 (N_13891,N_5430,N_7348);
xor U13892 (N_13892,N_8216,N_9544);
or U13893 (N_13893,N_9438,N_5431);
or U13894 (N_13894,N_7001,N_8175);
nor U13895 (N_13895,N_9501,N_7978);
or U13896 (N_13896,N_7673,N_6409);
xor U13897 (N_13897,N_9705,N_7385);
or U13898 (N_13898,N_7459,N_8735);
xor U13899 (N_13899,N_9114,N_5541);
or U13900 (N_13900,N_5481,N_7116);
nand U13901 (N_13901,N_6080,N_8406);
and U13902 (N_13902,N_5598,N_7769);
xor U13903 (N_13903,N_5806,N_7978);
or U13904 (N_13904,N_8184,N_8001);
or U13905 (N_13905,N_5945,N_5867);
nor U13906 (N_13906,N_5080,N_6448);
or U13907 (N_13907,N_7109,N_9281);
nand U13908 (N_13908,N_5681,N_6620);
or U13909 (N_13909,N_8346,N_8084);
and U13910 (N_13910,N_5679,N_6899);
or U13911 (N_13911,N_6407,N_7806);
or U13912 (N_13912,N_9110,N_8506);
nand U13913 (N_13913,N_5773,N_8593);
nor U13914 (N_13914,N_6812,N_6633);
or U13915 (N_13915,N_8464,N_7982);
or U13916 (N_13916,N_7856,N_9409);
or U13917 (N_13917,N_9047,N_9191);
nor U13918 (N_13918,N_5554,N_5862);
or U13919 (N_13919,N_7504,N_8312);
xor U13920 (N_13920,N_5605,N_6041);
or U13921 (N_13921,N_7190,N_6359);
or U13922 (N_13922,N_9751,N_8485);
xnor U13923 (N_13923,N_6762,N_7062);
nor U13924 (N_13924,N_7497,N_6211);
or U13925 (N_13925,N_5563,N_7524);
nor U13926 (N_13926,N_6314,N_6790);
nand U13927 (N_13927,N_8863,N_9611);
nor U13928 (N_13928,N_5166,N_8770);
xor U13929 (N_13929,N_9304,N_6192);
nand U13930 (N_13930,N_8894,N_8441);
or U13931 (N_13931,N_5960,N_8143);
nor U13932 (N_13932,N_5786,N_8982);
nand U13933 (N_13933,N_5207,N_5214);
and U13934 (N_13934,N_8631,N_5882);
xor U13935 (N_13935,N_6029,N_9219);
nand U13936 (N_13936,N_9044,N_5463);
and U13937 (N_13937,N_6419,N_5710);
xor U13938 (N_13938,N_9060,N_9712);
or U13939 (N_13939,N_6869,N_9856);
and U13940 (N_13940,N_7915,N_8422);
and U13941 (N_13941,N_9882,N_5705);
nor U13942 (N_13942,N_6234,N_8930);
xor U13943 (N_13943,N_5320,N_9324);
nand U13944 (N_13944,N_6553,N_8848);
or U13945 (N_13945,N_6862,N_5848);
xor U13946 (N_13946,N_7525,N_7295);
or U13947 (N_13947,N_5181,N_9344);
and U13948 (N_13948,N_7463,N_7286);
or U13949 (N_13949,N_6773,N_6314);
nand U13950 (N_13950,N_8001,N_5668);
and U13951 (N_13951,N_6732,N_5527);
or U13952 (N_13952,N_6520,N_9095);
and U13953 (N_13953,N_5771,N_9230);
or U13954 (N_13954,N_7888,N_6230);
xor U13955 (N_13955,N_5965,N_7322);
nor U13956 (N_13956,N_6540,N_7828);
or U13957 (N_13957,N_8233,N_6035);
and U13958 (N_13958,N_5346,N_9301);
or U13959 (N_13959,N_9686,N_8122);
and U13960 (N_13960,N_5346,N_9543);
nand U13961 (N_13961,N_9064,N_8296);
nand U13962 (N_13962,N_9757,N_6482);
nand U13963 (N_13963,N_8840,N_5489);
and U13964 (N_13964,N_9644,N_6313);
nor U13965 (N_13965,N_9960,N_5143);
and U13966 (N_13966,N_7674,N_7011);
xnor U13967 (N_13967,N_7424,N_6382);
xnor U13968 (N_13968,N_9095,N_6213);
or U13969 (N_13969,N_5133,N_6562);
nand U13970 (N_13970,N_6885,N_5741);
or U13971 (N_13971,N_6713,N_8232);
nor U13972 (N_13972,N_9984,N_9837);
or U13973 (N_13973,N_7736,N_9176);
nor U13974 (N_13974,N_5651,N_8282);
xnor U13975 (N_13975,N_7332,N_7153);
nor U13976 (N_13976,N_8560,N_7014);
and U13977 (N_13977,N_8275,N_5013);
or U13978 (N_13978,N_9394,N_7663);
nor U13979 (N_13979,N_9619,N_6703);
nand U13980 (N_13980,N_6443,N_9075);
nor U13981 (N_13981,N_7329,N_8831);
or U13982 (N_13982,N_9699,N_6708);
and U13983 (N_13983,N_6365,N_8175);
or U13984 (N_13984,N_6449,N_6693);
nor U13985 (N_13985,N_7979,N_8005);
nor U13986 (N_13986,N_6702,N_6352);
nor U13987 (N_13987,N_6125,N_8020);
and U13988 (N_13988,N_5400,N_6259);
xor U13989 (N_13989,N_9464,N_8594);
nor U13990 (N_13990,N_9451,N_5028);
nand U13991 (N_13991,N_6387,N_8971);
and U13992 (N_13992,N_8505,N_7842);
and U13993 (N_13993,N_9666,N_6839);
xor U13994 (N_13994,N_9287,N_7322);
nand U13995 (N_13995,N_5050,N_5168);
or U13996 (N_13996,N_8270,N_7992);
and U13997 (N_13997,N_6111,N_7372);
or U13998 (N_13998,N_9839,N_8398);
xnor U13999 (N_13999,N_6384,N_9510);
nor U14000 (N_14000,N_8267,N_6797);
nor U14001 (N_14001,N_6277,N_5005);
or U14002 (N_14002,N_5951,N_8524);
and U14003 (N_14003,N_9378,N_5416);
nor U14004 (N_14004,N_6052,N_8494);
or U14005 (N_14005,N_5102,N_7947);
nand U14006 (N_14006,N_9213,N_9122);
xnor U14007 (N_14007,N_6989,N_6498);
and U14008 (N_14008,N_5712,N_6137);
xnor U14009 (N_14009,N_9930,N_8655);
xor U14010 (N_14010,N_9572,N_7647);
xnor U14011 (N_14011,N_8663,N_8683);
xnor U14012 (N_14012,N_8480,N_5653);
or U14013 (N_14013,N_7180,N_7400);
and U14014 (N_14014,N_8461,N_8880);
or U14015 (N_14015,N_9953,N_8695);
nor U14016 (N_14016,N_5440,N_7770);
nor U14017 (N_14017,N_9804,N_6105);
or U14018 (N_14018,N_8101,N_6369);
or U14019 (N_14019,N_9124,N_7990);
and U14020 (N_14020,N_9546,N_6905);
xor U14021 (N_14021,N_7590,N_7564);
nand U14022 (N_14022,N_8143,N_9992);
xor U14023 (N_14023,N_9657,N_7705);
and U14024 (N_14024,N_9210,N_8452);
or U14025 (N_14025,N_9020,N_8714);
nand U14026 (N_14026,N_8050,N_7271);
nor U14027 (N_14027,N_6633,N_9017);
nor U14028 (N_14028,N_8361,N_8197);
or U14029 (N_14029,N_7521,N_6062);
and U14030 (N_14030,N_7915,N_7254);
or U14031 (N_14031,N_5653,N_6498);
and U14032 (N_14032,N_7308,N_7817);
nor U14033 (N_14033,N_9419,N_9846);
nor U14034 (N_14034,N_5390,N_9385);
nand U14035 (N_14035,N_9680,N_6137);
nor U14036 (N_14036,N_9957,N_9796);
nand U14037 (N_14037,N_6945,N_7574);
nor U14038 (N_14038,N_5718,N_5128);
nand U14039 (N_14039,N_6451,N_5709);
nor U14040 (N_14040,N_5886,N_7026);
xnor U14041 (N_14041,N_8482,N_5348);
nor U14042 (N_14042,N_6779,N_6183);
nand U14043 (N_14043,N_7412,N_8517);
and U14044 (N_14044,N_7626,N_8427);
xor U14045 (N_14045,N_7675,N_9375);
nor U14046 (N_14046,N_8767,N_6356);
xor U14047 (N_14047,N_7672,N_8479);
and U14048 (N_14048,N_6689,N_9016);
or U14049 (N_14049,N_5570,N_5793);
nor U14050 (N_14050,N_9794,N_8145);
nor U14051 (N_14051,N_7991,N_7626);
or U14052 (N_14052,N_7813,N_5861);
and U14053 (N_14053,N_8215,N_6802);
xnor U14054 (N_14054,N_6248,N_6312);
nand U14055 (N_14055,N_8719,N_5058);
nand U14056 (N_14056,N_6177,N_5075);
nand U14057 (N_14057,N_7725,N_7253);
nand U14058 (N_14058,N_6147,N_5396);
and U14059 (N_14059,N_6574,N_6179);
and U14060 (N_14060,N_9995,N_7338);
or U14061 (N_14061,N_7686,N_7967);
nand U14062 (N_14062,N_5826,N_6841);
or U14063 (N_14063,N_6024,N_9931);
xor U14064 (N_14064,N_5012,N_5602);
xor U14065 (N_14065,N_9084,N_5042);
nor U14066 (N_14066,N_9630,N_6444);
nand U14067 (N_14067,N_8338,N_8372);
and U14068 (N_14068,N_6851,N_8075);
nor U14069 (N_14069,N_6285,N_6459);
and U14070 (N_14070,N_6343,N_6127);
nand U14071 (N_14071,N_6366,N_5962);
xor U14072 (N_14072,N_9852,N_5883);
nand U14073 (N_14073,N_7464,N_8119);
or U14074 (N_14074,N_7569,N_7059);
nand U14075 (N_14075,N_8874,N_8022);
or U14076 (N_14076,N_8006,N_6418);
and U14077 (N_14077,N_8134,N_5927);
nor U14078 (N_14078,N_6900,N_5490);
xnor U14079 (N_14079,N_7388,N_6082);
and U14080 (N_14080,N_6151,N_9351);
nand U14081 (N_14081,N_9505,N_5786);
xnor U14082 (N_14082,N_7308,N_6907);
xor U14083 (N_14083,N_6235,N_6355);
and U14084 (N_14084,N_7676,N_8160);
and U14085 (N_14085,N_9065,N_9529);
nor U14086 (N_14086,N_5178,N_8091);
or U14087 (N_14087,N_5790,N_7272);
and U14088 (N_14088,N_6238,N_8924);
xor U14089 (N_14089,N_9621,N_6106);
or U14090 (N_14090,N_9122,N_8002);
nor U14091 (N_14091,N_8282,N_8010);
xor U14092 (N_14092,N_8739,N_8141);
nor U14093 (N_14093,N_6563,N_6576);
and U14094 (N_14094,N_7834,N_8910);
nand U14095 (N_14095,N_7341,N_6729);
xnor U14096 (N_14096,N_8643,N_6963);
nand U14097 (N_14097,N_8166,N_8614);
xor U14098 (N_14098,N_9907,N_8431);
xor U14099 (N_14099,N_6456,N_8888);
nand U14100 (N_14100,N_6260,N_7092);
xnor U14101 (N_14101,N_7096,N_6612);
xor U14102 (N_14102,N_9694,N_7345);
or U14103 (N_14103,N_6014,N_9994);
or U14104 (N_14104,N_9952,N_9405);
and U14105 (N_14105,N_9409,N_8940);
nand U14106 (N_14106,N_6933,N_7017);
and U14107 (N_14107,N_5110,N_9364);
nor U14108 (N_14108,N_5510,N_9331);
xnor U14109 (N_14109,N_9129,N_5799);
xnor U14110 (N_14110,N_5597,N_8071);
xnor U14111 (N_14111,N_5815,N_6793);
nor U14112 (N_14112,N_9642,N_9075);
nor U14113 (N_14113,N_7610,N_9828);
and U14114 (N_14114,N_7973,N_5625);
and U14115 (N_14115,N_8246,N_9663);
xor U14116 (N_14116,N_5019,N_6054);
xnor U14117 (N_14117,N_5291,N_8272);
and U14118 (N_14118,N_5286,N_7320);
or U14119 (N_14119,N_5132,N_8079);
xor U14120 (N_14120,N_8566,N_7388);
nor U14121 (N_14121,N_5436,N_7942);
or U14122 (N_14122,N_7167,N_9994);
xnor U14123 (N_14123,N_6292,N_7739);
xor U14124 (N_14124,N_8771,N_8427);
nor U14125 (N_14125,N_5885,N_8881);
nand U14126 (N_14126,N_8294,N_6983);
xnor U14127 (N_14127,N_8144,N_7105);
xnor U14128 (N_14128,N_6784,N_9420);
or U14129 (N_14129,N_7897,N_6404);
and U14130 (N_14130,N_9636,N_7028);
nor U14131 (N_14131,N_9192,N_5948);
or U14132 (N_14132,N_7733,N_7967);
nor U14133 (N_14133,N_7904,N_8221);
xor U14134 (N_14134,N_8159,N_7848);
or U14135 (N_14135,N_9138,N_8312);
nand U14136 (N_14136,N_7172,N_8506);
or U14137 (N_14137,N_6546,N_7988);
nand U14138 (N_14138,N_8318,N_5040);
nor U14139 (N_14139,N_5358,N_8820);
xor U14140 (N_14140,N_6868,N_8595);
nor U14141 (N_14141,N_5411,N_6062);
and U14142 (N_14142,N_9262,N_7224);
or U14143 (N_14143,N_5388,N_7712);
nor U14144 (N_14144,N_8251,N_7904);
nor U14145 (N_14145,N_8261,N_5986);
nor U14146 (N_14146,N_8452,N_6019);
nor U14147 (N_14147,N_9357,N_9278);
or U14148 (N_14148,N_8160,N_5175);
or U14149 (N_14149,N_7499,N_8886);
or U14150 (N_14150,N_6938,N_8233);
and U14151 (N_14151,N_8947,N_8372);
nor U14152 (N_14152,N_8661,N_9579);
or U14153 (N_14153,N_8796,N_8958);
nand U14154 (N_14154,N_9173,N_6559);
nor U14155 (N_14155,N_6278,N_6360);
and U14156 (N_14156,N_5057,N_7895);
or U14157 (N_14157,N_7785,N_5039);
xor U14158 (N_14158,N_9107,N_9825);
xor U14159 (N_14159,N_7027,N_7406);
nand U14160 (N_14160,N_8721,N_8894);
xnor U14161 (N_14161,N_5701,N_6114);
and U14162 (N_14162,N_6267,N_8807);
nand U14163 (N_14163,N_6548,N_8050);
xnor U14164 (N_14164,N_7666,N_8250);
nand U14165 (N_14165,N_6889,N_5541);
nand U14166 (N_14166,N_6920,N_6641);
xor U14167 (N_14167,N_5624,N_7276);
nand U14168 (N_14168,N_6807,N_6966);
and U14169 (N_14169,N_8820,N_9085);
nand U14170 (N_14170,N_9192,N_6110);
nor U14171 (N_14171,N_6774,N_8316);
nor U14172 (N_14172,N_7003,N_8786);
xor U14173 (N_14173,N_7908,N_7867);
or U14174 (N_14174,N_7429,N_7029);
and U14175 (N_14175,N_5303,N_9664);
nor U14176 (N_14176,N_8905,N_9005);
nor U14177 (N_14177,N_7221,N_8058);
nor U14178 (N_14178,N_6129,N_9393);
or U14179 (N_14179,N_6474,N_9379);
nor U14180 (N_14180,N_9981,N_6875);
xnor U14181 (N_14181,N_8303,N_5710);
xnor U14182 (N_14182,N_7757,N_6614);
or U14183 (N_14183,N_8942,N_6524);
xor U14184 (N_14184,N_8191,N_9236);
nor U14185 (N_14185,N_9433,N_8001);
xnor U14186 (N_14186,N_7323,N_6368);
xor U14187 (N_14187,N_5625,N_8975);
nand U14188 (N_14188,N_9193,N_9858);
xnor U14189 (N_14189,N_6875,N_9104);
or U14190 (N_14190,N_6768,N_6684);
nor U14191 (N_14191,N_6215,N_6185);
or U14192 (N_14192,N_7547,N_9270);
and U14193 (N_14193,N_6529,N_8575);
or U14194 (N_14194,N_9795,N_6596);
nand U14195 (N_14195,N_5335,N_5786);
xor U14196 (N_14196,N_5754,N_7408);
nand U14197 (N_14197,N_7245,N_8785);
nor U14198 (N_14198,N_6806,N_6799);
nor U14199 (N_14199,N_8596,N_8713);
and U14200 (N_14200,N_9514,N_6639);
and U14201 (N_14201,N_5845,N_6012);
xnor U14202 (N_14202,N_8042,N_8202);
nand U14203 (N_14203,N_6011,N_8208);
or U14204 (N_14204,N_9868,N_8725);
nor U14205 (N_14205,N_7587,N_6423);
and U14206 (N_14206,N_6892,N_5200);
or U14207 (N_14207,N_5569,N_7428);
and U14208 (N_14208,N_5509,N_6692);
or U14209 (N_14209,N_8944,N_6409);
nand U14210 (N_14210,N_9912,N_9462);
xor U14211 (N_14211,N_6468,N_7171);
nand U14212 (N_14212,N_9912,N_9843);
nor U14213 (N_14213,N_8932,N_8360);
xor U14214 (N_14214,N_5702,N_6130);
nand U14215 (N_14215,N_7813,N_7634);
xor U14216 (N_14216,N_9581,N_6159);
nand U14217 (N_14217,N_9797,N_7443);
and U14218 (N_14218,N_9591,N_6243);
or U14219 (N_14219,N_7458,N_5306);
or U14220 (N_14220,N_9630,N_6560);
or U14221 (N_14221,N_9449,N_7227);
or U14222 (N_14222,N_6895,N_6021);
or U14223 (N_14223,N_8346,N_6885);
and U14224 (N_14224,N_8263,N_7315);
nand U14225 (N_14225,N_5235,N_7807);
nor U14226 (N_14226,N_7251,N_8459);
nor U14227 (N_14227,N_8268,N_5482);
and U14228 (N_14228,N_8509,N_7415);
nor U14229 (N_14229,N_5563,N_5155);
or U14230 (N_14230,N_5380,N_5239);
xor U14231 (N_14231,N_8517,N_7385);
nand U14232 (N_14232,N_9927,N_8776);
xor U14233 (N_14233,N_7918,N_7229);
nand U14234 (N_14234,N_6849,N_7835);
and U14235 (N_14235,N_8355,N_6070);
or U14236 (N_14236,N_5766,N_9364);
nor U14237 (N_14237,N_7555,N_9853);
or U14238 (N_14238,N_6592,N_8552);
xnor U14239 (N_14239,N_7050,N_5768);
or U14240 (N_14240,N_9421,N_7974);
and U14241 (N_14241,N_6616,N_5600);
and U14242 (N_14242,N_6461,N_6085);
and U14243 (N_14243,N_7158,N_7160);
and U14244 (N_14244,N_8764,N_9281);
or U14245 (N_14245,N_6160,N_5898);
and U14246 (N_14246,N_8406,N_9421);
xor U14247 (N_14247,N_8302,N_5199);
nand U14248 (N_14248,N_6947,N_5519);
or U14249 (N_14249,N_5552,N_7874);
nor U14250 (N_14250,N_6998,N_6348);
and U14251 (N_14251,N_9325,N_5933);
nand U14252 (N_14252,N_7707,N_7721);
and U14253 (N_14253,N_5211,N_9045);
nor U14254 (N_14254,N_8676,N_6310);
xor U14255 (N_14255,N_5449,N_6871);
nor U14256 (N_14256,N_8787,N_7297);
nand U14257 (N_14257,N_7504,N_5702);
nor U14258 (N_14258,N_8868,N_9069);
and U14259 (N_14259,N_8380,N_8911);
nand U14260 (N_14260,N_9997,N_7518);
or U14261 (N_14261,N_9035,N_6529);
nor U14262 (N_14262,N_8917,N_9925);
xor U14263 (N_14263,N_5353,N_6958);
nor U14264 (N_14264,N_8519,N_9357);
nor U14265 (N_14265,N_8682,N_7957);
xnor U14266 (N_14266,N_5234,N_6111);
nand U14267 (N_14267,N_5550,N_7670);
xnor U14268 (N_14268,N_6188,N_7037);
nor U14269 (N_14269,N_5065,N_9235);
and U14270 (N_14270,N_8285,N_9053);
nor U14271 (N_14271,N_8552,N_9087);
nor U14272 (N_14272,N_6792,N_6357);
nand U14273 (N_14273,N_7785,N_7481);
or U14274 (N_14274,N_8620,N_9947);
or U14275 (N_14275,N_8678,N_5060);
and U14276 (N_14276,N_7469,N_7597);
and U14277 (N_14277,N_5428,N_6979);
and U14278 (N_14278,N_8594,N_7358);
or U14279 (N_14279,N_6418,N_5522);
xnor U14280 (N_14280,N_9976,N_9402);
nor U14281 (N_14281,N_5466,N_6232);
xnor U14282 (N_14282,N_9828,N_5961);
nor U14283 (N_14283,N_7936,N_8963);
nand U14284 (N_14284,N_7715,N_7804);
xor U14285 (N_14285,N_5023,N_6200);
nor U14286 (N_14286,N_8057,N_5181);
nand U14287 (N_14287,N_5413,N_5960);
and U14288 (N_14288,N_6967,N_8504);
or U14289 (N_14289,N_9950,N_6425);
nor U14290 (N_14290,N_7743,N_8353);
and U14291 (N_14291,N_6274,N_8741);
or U14292 (N_14292,N_8649,N_5787);
and U14293 (N_14293,N_8069,N_9577);
nor U14294 (N_14294,N_5519,N_8204);
or U14295 (N_14295,N_7879,N_5713);
nor U14296 (N_14296,N_5795,N_9244);
nor U14297 (N_14297,N_9642,N_7305);
xor U14298 (N_14298,N_8362,N_7959);
or U14299 (N_14299,N_9306,N_5434);
nand U14300 (N_14300,N_8784,N_8013);
or U14301 (N_14301,N_6847,N_8316);
and U14302 (N_14302,N_7183,N_7717);
xnor U14303 (N_14303,N_9163,N_5478);
xor U14304 (N_14304,N_9092,N_8202);
nor U14305 (N_14305,N_9205,N_9846);
and U14306 (N_14306,N_6551,N_9780);
and U14307 (N_14307,N_8888,N_8616);
nor U14308 (N_14308,N_7759,N_5105);
xor U14309 (N_14309,N_6114,N_8358);
and U14310 (N_14310,N_8150,N_9437);
nand U14311 (N_14311,N_9424,N_7433);
and U14312 (N_14312,N_6897,N_9064);
nand U14313 (N_14313,N_5702,N_5001);
xnor U14314 (N_14314,N_9891,N_8922);
and U14315 (N_14315,N_7405,N_7746);
or U14316 (N_14316,N_7365,N_7997);
nand U14317 (N_14317,N_8509,N_9720);
nor U14318 (N_14318,N_8516,N_5654);
and U14319 (N_14319,N_5058,N_6906);
nand U14320 (N_14320,N_8132,N_8698);
and U14321 (N_14321,N_9804,N_9346);
or U14322 (N_14322,N_8264,N_8826);
nor U14323 (N_14323,N_7636,N_9695);
nor U14324 (N_14324,N_6738,N_8603);
nor U14325 (N_14325,N_9752,N_5946);
and U14326 (N_14326,N_5854,N_9137);
or U14327 (N_14327,N_8761,N_8182);
nor U14328 (N_14328,N_7099,N_7126);
or U14329 (N_14329,N_7876,N_7729);
nand U14330 (N_14330,N_6429,N_6124);
nor U14331 (N_14331,N_6086,N_7383);
nor U14332 (N_14332,N_5311,N_5680);
and U14333 (N_14333,N_9202,N_5598);
nand U14334 (N_14334,N_7559,N_7783);
nor U14335 (N_14335,N_5360,N_6975);
nand U14336 (N_14336,N_7223,N_5445);
nand U14337 (N_14337,N_8763,N_7783);
xor U14338 (N_14338,N_9274,N_6020);
nand U14339 (N_14339,N_8395,N_9918);
and U14340 (N_14340,N_7169,N_7277);
nor U14341 (N_14341,N_6488,N_9577);
xnor U14342 (N_14342,N_9370,N_9645);
xnor U14343 (N_14343,N_7631,N_9163);
or U14344 (N_14344,N_5066,N_7513);
xnor U14345 (N_14345,N_8233,N_7544);
nand U14346 (N_14346,N_5001,N_6775);
nand U14347 (N_14347,N_5330,N_8705);
nor U14348 (N_14348,N_7461,N_8177);
nor U14349 (N_14349,N_5977,N_8970);
and U14350 (N_14350,N_8277,N_8643);
or U14351 (N_14351,N_7780,N_7441);
nor U14352 (N_14352,N_5494,N_5118);
nand U14353 (N_14353,N_7334,N_7198);
xnor U14354 (N_14354,N_6114,N_9323);
or U14355 (N_14355,N_5500,N_7077);
and U14356 (N_14356,N_9884,N_6499);
xor U14357 (N_14357,N_8417,N_7946);
and U14358 (N_14358,N_6774,N_5613);
and U14359 (N_14359,N_9858,N_8271);
nand U14360 (N_14360,N_9188,N_9279);
nand U14361 (N_14361,N_8342,N_5547);
nand U14362 (N_14362,N_9117,N_8635);
nand U14363 (N_14363,N_9311,N_5433);
or U14364 (N_14364,N_9634,N_7880);
nand U14365 (N_14365,N_5790,N_6183);
or U14366 (N_14366,N_7191,N_8559);
nor U14367 (N_14367,N_6573,N_6151);
nor U14368 (N_14368,N_5618,N_7987);
nor U14369 (N_14369,N_8128,N_6778);
nand U14370 (N_14370,N_9862,N_9740);
xnor U14371 (N_14371,N_6883,N_5926);
and U14372 (N_14372,N_6085,N_8323);
or U14373 (N_14373,N_5342,N_7779);
and U14374 (N_14374,N_8538,N_5017);
or U14375 (N_14375,N_7435,N_5321);
or U14376 (N_14376,N_8218,N_7612);
or U14377 (N_14377,N_7637,N_7675);
nand U14378 (N_14378,N_5126,N_5778);
xnor U14379 (N_14379,N_6713,N_5093);
or U14380 (N_14380,N_5701,N_8896);
or U14381 (N_14381,N_9310,N_9851);
nand U14382 (N_14382,N_8079,N_9814);
xor U14383 (N_14383,N_7588,N_9888);
and U14384 (N_14384,N_7869,N_6499);
nor U14385 (N_14385,N_7391,N_9088);
nand U14386 (N_14386,N_9608,N_6707);
nand U14387 (N_14387,N_8749,N_9503);
or U14388 (N_14388,N_7202,N_7792);
nand U14389 (N_14389,N_8868,N_5466);
and U14390 (N_14390,N_6573,N_6869);
nand U14391 (N_14391,N_8929,N_8573);
and U14392 (N_14392,N_5994,N_7901);
and U14393 (N_14393,N_7899,N_5888);
nor U14394 (N_14394,N_8974,N_6148);
and U14395 (N_14395,N_8690,N_8502);
or U14396 (N_14396,N_7416,N_6371);
nor U14397 (N_14397,N_6122,N_5299);
and U14398 (N_14398,N_8820,N_8729);
or U14399 (N_14399,N_9253,N_7117);
or U14400 (N_14400,N_6659,N_8820);
xnor U14401 (N_14401,N_5041,N_9954);
nor U14402 (N_14402,N_8397,N_8805);
xor U14403 (N_14403,N_5968,N_6641);
nand U14404 (N_14404,N_5624,N_6805);
xor U14405 (N_14405,N_9830,N_9465);
nand U14406 (N_14406,N_9403,N_7376);
nand U14407 (N_14407,N_8363,N_9791);
nor U14408 (N_14408,N_9356,N_8903);
xnor U14409 (N_14409,N_8202,N_8663);
and U14410 (N_14410,N_8669,N_5419);
xor U14411 (N_14411,N_9450,N_7264);
xor U14412 (N_14412,N_9348,N_7886);
or U14413 (N_14413,N_5609,N_6894);
nor U14414 (N_14414,N_9381,N_7408);
and U14415 (N_14415,N_8795,N_9670);
nor U14416 (N_14416,N_6440,N_9122);
nor U14417 (N_14417,N_7360,N_9731);
xor U14418 (N_14418,N_9078,N_6783);
and U14419 (N_14419,N_8033,N_5845);
or U14420 (N_14420,N_9545,N_6928);
and U14421 (N_14421,N_9739,N_9923);
nand U14422 (N_14422,N_9288,N_8139);
or U14423 (N_14423,N_8098,N_7957);
nand U14424 (N_14424,N_6736,N_6626);
nand U14425 (N_14425,N_6798,N_6319);
xnor U14426 (N_14426,N_8174,N_5517);
xor U14427 (N_14427,N_7180,N_8844);
nor U14428 (N_14428,N_7095,N_8371);
and U14429 (N_14429,N_5329,N_5371);
and U14430 (N_14430,N_7343,N_5411);
nand U14431 (N_14431,N_5963,N_8422);
nand U14432 (N_14432,N_5759,N_6649);
or U14433 (N_14433,N_8621,N_6165);
or U14434 (N_14434,N_9637,N_7678);
and U14435 (N_14435,N_6251,N_9410);
nor U14436 (N_14436,N_7874,N_5922);
and U14437 (N_14437,N_7451,N_9482);
or U14438 (N_14438,N_7189,N_9421);
or U14439 (N_14439,N_5826,N_9319);
or U14440 (N_14440,N_6834,N_8080);
and U14441 (N_14441,N_6432,N_7398);
nor U14442 (N_14442,N_8216,N_7634);
xor U14443 (N_14443,N_5252,N_9109);
xor U14444 (N_14444,N_8245,N_6836);
or U14445 (N_14445,N_5428,N_7726);
and U14446 (N_14446,N_9726,N_5960);
or U14447 (N_14447,N_6134,N_5504);
nor U14448 (N_14448,N_5049,N_5282);
and U14449 (N_14449,N_5588,N_5782);
or U14450 (N_14450,N_5101,N_5171);
nand U14451 (N_14451,N_7935,N_6006);
or U14452 (N_14452,N_5772,N_7118);
nor U14453 (N_14453,N_8984,N_9698);
nor U14454 (N_14454,N_5242,N_5314);
nor U14455 (N_14455,N_6784,N_8075);
nand U14456 (N_14456,N_6245,N_7207);
xnor U14457 (N_14457,N_6202,N_7443);
xor U14458 (N_14458,N_8056,N_6633);
and U14459 (N_14459,N_8942,N_8722);
xor U14460 (N_14460,N_6581,N_6341);
xnor U14461 (N_14461,N_6886,N_6425);
nand U14462 (N_14462,N_9455,N_9542);
or U14463 (N_14463,N_7980,N_5398);
nand U14464 (N_14464,N_7939,N_9590);
xnor U14465 (N_14465,N_5469,N_9986);
and U14466 (N_14466,N_7109,N_6808);
nor U14467 (N_14467,N_5993,N_8178);
nor U14468 (N_14468,N_5041,N_9664);
nand U14469 (N_14469,N_9082,N_9021);
nand U14470 (N_14470,N_6921,N_7448);
nand U14471 (N_14471,N_5378,N_9118);
or U14472 (N_14472,N_9667,N_5666);
nor U14473 (N_14473,N_5971,N_8138);
or U14474 (N_14474,N_5909,N_9431);
nor U14475 (N_14475,N_6412,N_9270);
xor U14476 (N_14476,N_8682,N_5386);
or U14477 (N_14477,N_6402,N_5874);
xnor U14478 (N_14478,N_6519,N_5553);
and U14479 (N_14479,N_9927,N_6748);
nor U14480 (N_14480,N_6283,N_7756);
nand U14481 (N_14481,N_6409,N_9789);
xor U14482 (N_14482,N_5547,N_5532);
or U14483 (N_14483,N_5741,N_6048);
or U14484 (N_14484,N_8006,N_5801);
nor U14485 (N_14485,N_5903,N_7218);
nor U14486 (N_14486,N_5975,N_9485);
nor U14487 (N_14487,N_9697,N_9513);
and U14488 (N_14488,N_5292,N_5620);
nand U14489 (N_14489,N_9882,N_6471);
and U14490 (N_14490,N_7661,N_9158);
nor U14491 (N_14491,N_6395,N_9133);
xnor U14492 (N_14492,N_9587,N_8869);
xor U14493 (N_14493,N_7296,N_7975);
or U14494 (N_14494,N_5334,N_7235);
xor U14495 (N_14495,N_7645,N_9397);
nand U14496 (N_14496,N_7087,N_6705);
xor U14497 (N_14497,N_7929,N_6195);
nor U14498 (N_14498,N_5077,N_7988);
nand U14499 (N_14499,N_9986,N_9917);
nand U14500 (N_14500,N_5696,N_8961);
or U14501 (N_14501,N_7417,N_7640);
xnor U14502 (N_14502,N_7580,N_6495);
nand U14503 (N_14503,N_9540,N_7571);
nand U14504 (N_14504,N_7924,N_7177);
or U14505 (N_14505,N_7427,N_8757);
nor U14506 (N_14506,N_9023,N_5760);
nand U14507 (N_14507,N_8357,N_8783);
nand U14508 (N_14508,N_7546,N_7647);
and U14509 (N_14509,N_9936,N_7685);
nor U14510 (N_14510,N_9628,N_9830);
nor U14511 (N_14511,N_6922,N_5899);
nand U14512 (N_14512,N_9864,N_8814);
or U14513 (N_14513,N_5185,N_8673);
or U14514 (N_14514,N_9310,N_6564);
xnor U14515 (N_14515,N_8155,N_7055);
xnor U14516 (N_14516,N_5244,N_6196);
or U14517 (N_14517,N_5602,N_6508);
and U14518 (N_14518,N_6785,N_5795);
xnor U14519 (N_14519,N_5873,N_5441);
xnor U14520 (N_14520,N_7924,N_6147);
and U14521 (N_14521,N_8328,N_6509);
nand U14522 (N_14522,N_5878,N_7386);
or U14523 (N_14523,N_9338,N_6980);
nand U14524 (N_14524,N_7829,N_5571);
and U14525 (N_14525,N_6164,N_9393);
nand U14526 (N_14526,N_6454,N_7482);
nor U14527 (N_14527,N_9644,N_6503);
xor U14528 (N_14528,N_9722,N_6229);
nor U14529 (N_14529,N_9412,N_9978);
xnor U14530 (N_14530,N_7209,N_7963);
nor U14531 (N_14531,N_7274,N_5149);
nand U14532 (N_14532,N_9838,N_6408);
and U14533 (N_14533,N_6941,N_6160);
nor U14534 (N_14534,N_8710,N_7762);
or U14535 (N_14535,N_7568,N_5767);
nand U14536 (N_14536,N_5511,N_7973);
and U14537 (N_14537,N_6418,N_9807);
or U14538 (N_14538,N_8499,N_9287);
xor U14539 (N_14539,N_8425,N_9385);
or U14540 (N_14540,N_9040,N_7008);
xor U14541 (N_14541,N_9520,N_9783);
and U14542 (N_14542,N_8137,N_9347);
nand U14543 (N_14543,N_7137,N_6405);
and U14544 (N_14544,N_6694,N_7183);
xnor U14545 (N_14545,N_5930,N_6365);
or U14546 (N_14546,N_8494,N_7249);
xnor U14547 (N_14547,N_8834,N_8490);
xnor U14548 (N_14548,N_7718,N_9533);
nor U14549 (N_14549,N_5238,N_5040);
nand U14550 (N_14550,N_7777,N_9597);
nand U14551 (N_14551,N_8527,N_5773);
xor U14552 (N_14552,N_7051,N_6402);
nand U14553 (N_14553,N_9111,N_6892);
nand U14554 (N_14554,N_8891,N_5738);
or U14555 (N_14555,N_5099,N_6108);
or U14556 (N_14556,N_6465,N_6461);
nor U14557 (N_14557,N_5493,N_6991);
nand U14558 (N_14558,N_9629,N_8279);
and U14559 (N_14559,N_9207,N_8636);
and U14560 (N_14560,N_7530,N_9228);
or U14561 (N_14561,N_7849,N_8400);
or U14562 (N_14562,N_8558,N_6931);
or U14563 (N_14563,N_7902,N_6974);
nor U14564 (N_14564,N_5884,N_8032);
or U14565 (N_14565,N_8998,N_9982);
nor U14566 (N_14566,N_7084,N_5066);
xnor U14567 (N_14567,N_6293,N_8590);
or U14568 (N_14568,N_9846,N_8067);
nand U14569 (N_14569,N_9485,N_7065);
nand U14570 (N_14570,N_5807,N_9906);
nor U14571 (N_14571,N_7508,N_9910);
nand U14572 (N_14572,N_7924,N_9466);
and U14573 (N_14573,N_5334,N_5176);
or U14574 (N_14574,N_9298,N_5114);
nand U14575 (N_14575,N_9898,N_5964);
nor U14576 (N_14576,N_9860,N_6137);
nand U14577 (N_14577,N_5921,N_5291);
or U14578 (N_14578,N_5588,N_9511);
nor U14579 (N_14579,N_8937,N_8651);
nor U14580 (N_14580,N_5477,N_5914);
nor U14581 (N_14581,N_7125,N_9760);
nor U14582 (N_14582,N_7439,N_5034);
and U14583 (N_14583,N_5593,N_6407);
nand U14584 (N_14584,N_9190,N_8998);
and U14585 (N_14585,N_9547,N_5982);
and U14586 (N_14586,N_5180,N_9006);
and U14587 (N_14587,N_5025,N_9524);
nand U14588 (N_14588,N_5257,N_6276);
and U14589 (N_14589,N_9576,N_9420);
or U14590 (N_14590,N_6525,N_6585);
or U14591 (N_14591,N_7704,N_7329);
nand U14592 (N_14592,N_5259,N_5311);
xor U14593 (N_14593,N_5902,N_9188);
and U14594 (N_14594,N_8074,N_5079);
and U14595 (N_14595,N_5307,N_8413);
or U14596 (N_14596,N_6314,N_7412);
xnor U14597 (N_14597,N_5487,N_7011);
and U14598 (N_14598,N_7416,N_7037);
xnor U14599 (N_14599,N_7699,N_6588);
xor U14600 (N_14600,N_5100,N_5042);
or U14601 (N_14601,N_8617,N_5386);
nand U14602 (N_14602,N_5449,N_5305);
or U14603 (N_14603,N_9603,N_9103);
xnor U14604 (N_14604,N_8949,N_8221);
nor U14605 (N_14605,N_8766,N_8857);
or U14606 (N_14606,N_9248,N_5198);
and U14607 (N_14607,N_9686,N_6927);
xor U14608 (N_14608,N_5890,N_5420);
xnor U14609 (N_14609,N_6508,N_5884);
nor U14610 (N_14610,N_8323,N_7451);
and U14611 (N_14611,N_9518,N_9878);
or U14612 (N_14612,N_7354,N_7279);
or U14613 (N_14613,N_7265,N_5708);
or U14614 (N_14614,N_7147,N_5958);
or U14615 (N_14615,N_7709,N_8352);
nor U14616 (N_14616,N_7991,N_8259);
and U14617 (N_14617,N_9484,N_8118);
nor U14618 (N_14618,N_7806,N_7139);
xnor U14619 (N_14619,N_9395,N_9339);
or U14620 (N_14620,N_8108,N_5410);
and U14621 (N_14621,N_6929,N_8499);
xor U14622 (N_14622,N_9522,N_5640);
xor U14623 (N_14623,N_5094,N_6160);
or U14624 (N_14624,N_7257,N_6446);
or U14625 (N_14625,N_6568,N_8140);
and U14626 (N_14626,N_9546,N_7914);
nand U14627 (N_14627,N_8610,N_7818);
nand U14628 (N_14628,N_8886,N_6051);
xnor U14629 (N_14629,N_9171,N_7366);
or U14630 (N_14630,N_6710,N_7257);
nor U14631 (N_14631,N_8136,N_7837);
nand U14632 (N_14632,N_7038,N_5465);
and U14633 (N_14633,N_7486,N_6188);
nand U14634 (N_14634,N_5624,N_5381);
nand U14635 (N_14635,N_8814,N_6517);
xnor U14636 (N_14636,N_7063,N_6778);
or U14637 (N_14637,N_6790,N_6952);
nand U14638 (N_14638,N_8037,N_9188);
nand U14639 (N_14639,N_9603,N_8914);
and U14640 (N_14640,N_7992,N_5893);
and U14641 (N_14641,N_8226,N_7915);
nand U14642 (N_14642,N_5574,N_8384);
and U14643 (N_14643,N_7298,N_7348);
and U14644 (N_14644,N_5452,N_6577);
and U14645 (N_14645,N_5919,N_9956);
and U14646 (N_14646,N_6492,N_9648);
xor U14647 (N_14647,N_8629,N_6005);
nor U14648 (N_14648,N_5780,N_6673);
nor U14649 (N_14649,N_6331,N_7183);
and U14650 (N_14650,N_6359,N_7386);
xor U14651 (N_14651,N_6088,N_7686);
nor U14652 (N_14652,N_9748,N_7502);
or U14653 (N_14653,N_8367,N_9153);
xnor U14654 (N_14654,N_9911,N_6853);
nor U14655 (N_14655,N_9505,N_6846);
or U14656 (N_14656,N_8850,N_7552);
nand U14657 (N_14657,N_9609,N_8375);
xnor U14658 (N_14658,N_6625,N_5276);
and U14659 (N_14659,N_9404,N_6400);
nor U14660 (N_14660,N_6632,N_5250);
or U14661 (N_14661,N_6332,N_7692);
nor U14662 (N_14662,N_8203,N_7900);
xor U14663 (N_14663,N_5396,N_6053);
nor U14664 (N_14664,N_8134,N_7197);
or U14665 (N_14665,N_6494,N_7319);
xor U14666 (N_14666,N_7879,N_6712);
nand U14667 (N_14667,N_7252,N_9645);
nand U14668 (N_14668,N_5657,N_6573);
or U14669 (N_14669,N_9446,N_9573);
or U14670 (N_14670,N_7592,N_8973);
xnor U14671 (N_14671,N_6794,N_5052);
xor U14672 (N_14672,N_8089,N_6373);
or U14673 (N_14673,N_5492,N_7865);
nor U14674 (N_14674,N_8607,N_6352);
or U14675 (N_14675,N_9805,N_5238);
nor U14676 (N_14676,N_5562,N_8334);
nand U14677 (N_14677,N_5225,N_9217);
and U14678 (N_14678,N_5090,N_9850);
and U14679 (N_14679,N_8997,N_9582);
nand U14680 (N_14680,N_9830,N_5873);
nand U14681 (N_14681,N_5692,N_5372);
nor U14682 (N_14682,N_6134,N_6650);
nor U14683 (N_14683,N_5259,N_6298);
nor U14684 (N_14684,N_9413,N_8078);
and U14685 (N_14685,N_6642,N_9960);
nor U14686 (N_14686,N_7901,N_6110);
or U14687 (N_14687,N_7206,N_8791);
xnor U14688 (N_14688,N_9778,N_7602);
xnor U14689 (N_14689,N_9977,N_8325);
or U14690 (N_14690,N_7498,N_9447);
xnor U14691 (N_14691,N_7798,N_7994);
nand U14692 (N_14692,N_5367,N_9752);
and U14693 (N_14693,N_6710,N_5977);
or U14694 (N_14694,N_9219,N_8306);
nand U14695 (N_14695,N_5098,N_9219);
nand U14696 (N_14696,N_8607,N_8437);
nor U14697 (N_14697,N_7060,N_8045);
xor U14698 (N_14698,N_7413,N_7689);
xor U14699 (N_14699,N_8119,N_5387);
nor U14700 (N_14700,N_8931,N_9348);
nand U14701 (N_14701,N_8443,N_6205);
nor U14702 (N_14702,N_7495,N_6225);
nor U14703 (N_14703,N_6709,N_9951);
or U14704 (N_14704,N_8978,N_6890);
xnor U14705 (N_14705,N_6150,N_9833);
nor U14706 (N_14706,N_5189,N_6465);
xor U14707 (N_14707,N_5336,N_6444);
nor U14708 (N_14708,N_6147,N_8654);
or U14709 (N_14709,N_5601,N_5514);
and U14710 (N_14710,N_5630,N_5531);
or U14711 (N_14711,N_6038,N_8942);
nor U14712 (N_14712,N_9947,N_5478);
or U14713 (N_14713,N_6220,N_5258);
and U14714 (N_14714,N_9777,N_9186);
xnor U14715 (N_14715,N_6239,N_9301);
nand U14716 (N_14716,N_5629,N_6565);
nor U14717 (N_14717,N_6612,N_5825);
or U14718 (N_14718,N_5270,N_9714);
and U14719 (N_14719,N_6571,N_7012);
nand U14720 (N_14720,N_9619,N_7589);
and U14721 (N_14721,N_9992,N_9900);
nand U14722 (N_14722,N_9003,N_8596);
nor U14723 (N_14723,N_6633,N_7103);
and U14724 (N_14724,N_7825,N_8650);
nor U14725 (N_14725,N_8780,N_8273);
nand U14726 (N_14726,N_9211,N_6450);
xnor U14727 (N_14727,N_9304,N_5582);
and U14728 (N_14728,N_6268,N_7587);
or U14729 (N_14729,N_6592,N_8020);
and U14730 (N_14730,N_5022,N_7071);
and U14731 (N_14731,N_9827,N_5735);
and U14732 (N_14732,N_9192,N_6802);
and U14733 (N_14733,N_6060,N_9542);
nor U14734 (N_14734,N_9287,N_6602);
and U14735 (N_14735,N_5692,N_6978);
nor U14736 (N_14736,N_8511,N_9322);
nand U14737 (N_14737,N_8972,N_8154);
and U14738 (N_14738,N_6733,N_9245);
nand U14739 (N_14739,N_5848,N_5117);
and U14740 (N_14740,N_6338,N_7312);
nor U14741 (N_14741,N_6881,N_6196);
and U14742 (N_14742,N_9941,N_7324);
nor U14743 (N_14743,N_8317,N_5381);
nand U14744 (N_14744,N_9854,N_6554);
or U14745 (N_14745,N_8933,N_7616);
nor U14746 (N_14746,N_8687,N_7802);
and U14747 (N_14747,N_5335,N_5546);
or U14748 (N_14748,N_6934,N_9653);
and U14749 (N_14749,N_5960,N_8400);
or U14750 (N_14750,N_5052,N_6440);
or U14751 (N_14751,N_9979,N_5029);
or U14752 (N_14752,N_7435,N_9463);
xor U14753 (N_14753,N_9751,N_6350);
or U14754 (N_14754,N_9913,N_9058);
nor U14755 (N_14755,N_9121,N_8608);
and U14756 (N_14756,N_7504,N_8939);
and U14757 (N_14757,N_7710,N_9208);
or U14758 (N_14758,N_8700,N_6531);
nand U14759 (N_14759,N_7010,N_7408);
or U14760 (N_14760,N_5022,N_5676);
xor U14761 (N_14761,N_9662,N_8921);
nor U14762 (N_14762,N_8391,N_9382);
xor U14763 (N_14763,N_7869,N_7172);
or U14764 (N_14764,N_8531,N_5671);
and U14765 (N_14765,N_8564,N_8886);
nand U14766 (N_14766,N_5397,N_5659);
and U14767 (N_14767,N_7352,N_5441);
or U14768 (N_14768,N_6746,N_7562);
or U14769 (N_14769,N_5711,N_8496);
and U14770 (N_14770,N_6017,N_5453);
xnor U14771 (N_14771,N_5266,N_5175);
nor U14772 (N_14772,N_5506,N_7261);
xnor U14773 (N_14773,N_5051,N_8985);
or U14774 (N_14774,N_9472,N_7764);
or U14775 (N_14775,N_7837,N_5364);
nand U14776 (N_14776,N_8377,N_7026);
and U14777 (N_14777,N_8699,N_6950);
xor U14778 (N_14778,N_7281,N_5850);
nor U14779 (N_14779,N_6623,N_7324);
nor U14780 (N_14780,N_5586,N_8994);
or U14781 (N_14781,N_6146,N_5079);
nand U14782 (N_14782,N_5382,N_8060);
and U14783 (N_14783,N_6302,N_7796);
nor U14784 (N_14784,N_8636,N_5089);
xnor U14785 (N_14785,N_9819,N_6325);
nand U14786 (N_14786,N_5556,N_5912);
and U14787 (N_14787,N_6470,N_9391);
xnor U14788 (N_14788,N_5996,N_8038);
nand U14789 (N_14789,N_8276,N_5005);
or U14790 (N_14790,N_6501,N_5869);
nor U14791 (N_14791,N_7040,N_9326);
nor U14792 (N_14792,N_6110,N_7003);
nand U14793 (N_14793,N_5107,N_7762);
nor U14794 (N_14794,N_7524,N_9453);
and U14795 (N_14795,N_6854,N_5051);
nand U14796 (N_14796,N_7022,N_5187);
and U14797 (N_14797,N_5029,N_8831);
xnor U14798 (N_14798,N_6908,N_8033);
and U14799 (N_14799,N_5065,N_8297);
xnor U14800 (N_14800,N_7194,N_8338);
nor U14801 (N_14801,N_7357,N_6851);
xnor U14802 (N_14802,N_5365,N_8772);
or U14803 (N_14803,N_6105,N_6980);
xor U14804 (N_14804,N_5845,N_9282);
or U14805 (N_14805,N_8014,N_8576);
nor U14806 (N_14806,N_6071,N_9656);
and U14807 (N_14807,N_7882,N_5788);
and U14808 (N_14808,N_9324,N_9446);
nand U14809 (N_14809,N_5129,N_5100);
xnor U14810 (N_14810,N_6077,N_9753);
nand U14811 (N_14811,N_6975,N_6780);
xor U14812 (N_14812,N_5886,N_5643);
nand U14813 (N_14813,N_9081,N_6322);
xor U14814 (N_14814,N_6208,N_5491);
or U14815 (N_14815,N_6025,N_7297);
or U14816 (N_14816,N_6165,N_7673);
nor U14817 (N_14817,N_5441,N_9427);
nor U14818 (N_14818,N_6959,N_6086);
xor U14819 (N_14819,N_8416,N_5155);
nand U14820 (N_14820,N_6538,N_5488);
or U14821 (N_14821,N_6107,N_6381);
nand U14822 (N_14822,N_7882,N_9649);
nor U14823 (N_14823,N_6359,N_5518);
xnor U14824 (N_14824,N_8872,N_6737);
or U14825 (N_14825,N_5346,N_9633);
or U14826 (N_14826,N_5407,N_9162);
xor U14827 (N_14827,N_7662,N_9230);
nand U14828 (N_14828,N_5548,N_8824);
or U14829 (N_14829,N_9773,N_9698);
nor U14830 (N_14830,N_5050,N_5944);
nand U14831 (N_14831,N_6153,N_5070);
and U14832 (N_14832,N_9195,N_5197);
and U14833 (N_14833,N_6936,N_8063);
xnor U14834 (N_14834,N_7241,N_8002);
and U14835 (N_14835,N_5779,N_9938);
xnor U14836 (N_14836,N_5363,N_5920);
and U14837 (N_14837,N_8790,N_7189);
xnor U14838 (N_14838,N_8097,N_7705);
xor U14839 (N_14839,N_5028,N_6540);
nor U14840 (N_14840,N_7811,N_9770);
nand U14841 (N_14841,N_5455,N_8681);
xnor U14842 (N_14842,N_8733,N_9859);
nand U14843 (N_14843,N_7875,N_8359);
nor U14844 (N_14844,N_5275,N_7218);
xnor U14845 (N_14845,N_8126,N_7816);
and U14846 (N_14846,N_9993,N_9738);
or U14847 (N_14847,N_6776,N_6888);
nand U14848 (N_14848,N_8412,N_6367);
or U14849 (N_14849,N_6648,N_7552);
and U14850 (N_14850,N_6644,N_7925);
nor U14851 (N_14851,N_5689,N_5760);
or U14852 (N_14852,N_7440,N_7047);
nor U14853 (N_14853,N_6378,N_8776);
xnor U14854 (N_14854,N_8046,N_5671);
nor U14855 (N_14855,N_6393,N_9498);
or U14856 (N_14856,N_5304,N_6255);
and U14857 (N_14857,N_6281,N_7214);
and U14858 (N_14858,N_9751,N_9672);
nor U14859 (N_14859,N_6485,N_7276);
or U14860 (N_14860,N_9498,N_7481);
nor U14861 (N_14861,N_9800,N_5449);
or U14862 (N_14862,N_6245,N_5170);
or U14863 (N_14863,N_7750,N_9086);
or U14864 (N_14864,N_5416,N_8150);
and U14865 (N_14865,N_6984,N_7350);
and U14866 (N_14866,N_9249,N_8130);
nor U14867 (N_14867,N_9562,N_7930);
and U14868 (N_14868,N_5099,N_7224);
nor U14869 (N_14869,N_8366,N_5133);
or U14870 (N_14870,N_9773,N_8373);
nor U14871 (N_14871,N_9840,N_8131);
nand U14872 (N_14872,N_7152,N_5569);
or U14873 (N_14873,N_9789,N_9500);
xor U14874 (N_14874,N_7086,N_9974);
nand U14875 (N_14875,N_9879,N_9796);
and U14876 (N_14876,N_5903,N_6859);
or U14877 (N_14877,N_8249,N_9645);
and U14878 (N_14878,N_6531,N_9299);
and U14879 (N_14879,N_8153,N_5798);
nand U14880 (N_14880,N_5144,N_7328);
or U14881 (N_14881,N_7377,N_8720);
nor U14882 (N_14882,N_5028,N_9036);
and U14883 (N_14883,N_9279,N_6671);
or U14884 (N_14884,N_8536,N_8989);
and U14885 (N_14885,N_8547,N_5612);
and U14886 (N_14886,N_7309,N_8821);
and U14887 (N_14887,N_7394,N_8953);
xnor U14888 (N_14888,N_7782,N_9932);
nor U14889 (N_14889,N_8180,N_9236);
or U14890 (N_14890,N_9254,N_9957);
nand U14891 (N_14891,N_5170,N_5819);
nand U14892 (N_14892,N_6087,N_8879);
and U14893 (N_14893,N_6694,N_5949);
nor U14894 (N_14894,N_5407,N_8866);
nor U14895 (N_14895,N_9200,N_9974);
xnor U14896 (N_14896,N_7130,N_8844);
or U14897 (N_14897,N_8372,N_7741);
nand U14898 (N_14898,N_8364,N_7000);
xor U14899 (N_14899,N_5740,N_8838);
nand U14900 (N_14900,N_6687,N_6139);
and U14901 (N_14901,N_5337,N_7613);
and U14902 (N_14902,N_9401,N_7142);
xor U14903 (N_14903,N_6206,N_7640);
nor U14904 (N_14904,N_7160,N_5511);
nor U14905 (N_14905,N_5481,N_7919);
and U14906 (N_14906,N_8852,N_7512);
nor U14907 (N_14907,N_6128,N_5195);
nor U14908 (N_14908,N_7651,N_5759);
nor U14909 (N_14909,N_9947,N_8183);
xnor U14910 (N_14910,N_5362,N_5611);
or U14911 (N_14911,N_9170,N_6185);
or U14912 (N_14912,N_7784,N_9765);
nor U14913 (N_14913,N_7652,N_6902);
xor U14914 (N_14914,N_5524,N_8960);
nor U14915 (N_14915,N_5308,N_9786);
nor U14916 (N_14916,N_7442,N_5930);
and U14917 (N_14917,N_5992,N_5324);
nor U14918 (N_14918,N_8901,N_5816);
xor U14919 (N_14919,N_9531,N_8890);
xor U14920 (N_14920,N_9105,N_8208);
nand U14921 (N_14921,N_6536,N_6366);
xor U14922 (N_14922,N_5871,N_5478);
nand U14923 (N_14923,N_6527,N_5831);
or U14924 (N_14924,N_6901,N_9051);
or U14925 (N_14925,N_8663,N_6949);
nor U14926 (N_14926,N_9657,N_5212);
nor U14927 (N_14927,N_7782,N_6706);
nand U14928 (N_14928,N_7575,N_5516);
xnor U14929 (N_14929,N_8610,N_6302);
xnor U14930 (N_14930,N_9492,N_6108);
or U14931 (N_14931,N_5969,N_5461);
nor U14932 (N_14932,N_9894,N_5470);
or U14933 (N_14933,N_5829,N_7404);
nand U14934 (N_14934,N_5722,N_5878);
or U14935 (N_14935,N_9872,N_5712);
xor U14936 (N_14936,N_7275,N_6851);
nand U14937 (N_14937,N_8750,N_9326);
nor U14938 (N_14938,N_5826,N_5991);
nand U14939 (N_14939,N_7741,N_9427);
or U14940 (N_14940,N_9503,N_8932);
xor U14941 (N_14941,N_5389,N_6061);
xor U14942 (N_14942,N_9599,N_7568);
or U14943 (N_14943,N_5521,N_8188);
or U14944 (N_14944,N_6470,N_6266);
nand U14945 (N_14945,N_8031,N_8984);
xnor U14946 (N_14946,N_5386,N_6533);
nand U14947 (N_14947,N_7505,N_5202);
nor U14948 (N_14948,N_7437,N_6264);
or U14949 (N_14949,N_5700,N_7928);
or U14950 (N_14950,N_5571,N_9920);
and U14951 (N_14951,N_8346,N_9957);
or U14952 (N_14952,N_5085,N_6955);
and U14953 (N_14953,N_8492,N_9409);
nor U14954 (N_14954,N_6860,N_8754);
and U14955 (N_14955,N_9863,N_7256);
nor U14956 (N_14956,N_7140,N_8596);
xnor U14957 (N_14957,N_6730,N_6045);
nand U14958 (N_14958,N_8595,N_9419);
or U14959 (N_14959,N_9122,N_7505);
nand U14960 (N_14960,N_9067,N_6711);
xor U14961 (N_14961,N_5806,N_8743);
nand U14962 (N_14962,N_7361,N_8627);
nor U14963 (N_14963,N_7229,N_8661);
nor U14964 (N_14964,N_6015,N_7026);
or U14965 (N_14965,N_5623,N_7442);
and U14966 (N_14966,N_7741,N_7709);
nand U14967 (N_14967,N_6874,N_6279);
or U14968 (N_14968,N_8809,N_8466);
xor U14969 (N_14969,N_6230,N_6460);
nand U14970 (N_14970,N_6966,N_9444);
or U14971 (N_14971,N_6406,N_6144);
xnor U14972 (N_14972,N_5661,N_9794);
or U14973 (N_14973,N_8140,N_9379);
or U14974 (N_14974,N_5439,N_8446);
or U14975 (N_14975,N_8704,N_9710);
xor U14976 (N_14976,N_8499,N_5792);
nor U14977 (N_14977,N_7225,N_6745);
nand U14978 (N_14978,N_6103,N_7963);
nor U14979 (N_14979,N_8102,N_9641);
xnor U14980 (N_14980,N_9043,N_8182);
or U14981 (N_14981,N_7559,N_8658);
xnor U14982 (N_14982,N_7940,N_7742);
and U14983 (N_14983,N_7744,N_6742);
nand U14984 (N_14984,N_7406,N_8176);
xnor U14985 (N_14985,N_5423,N_9544);
nand U14986 (N_14986,N_7669,N_8561);
and U14987 (N_14987,N_9106,N_5555);
and U14988 (N_14988,N_5137,N_6687);
xor U14989 (N_14989,N_5083,N_7437);
xor U14990 (N_14990,N_9373,N_8792);
nor U14991 (N_14991,N_7201,N_5815);
and U14992 (N_14992,N_8976,N_5218);
nor U14993 (N_14993,N_8890,N_6452);
or U14994 (N_14994,N_5164,N_9406);
or U14995 (N_14995,N_8065,N_6046);
and U14996 (N_14996,N_8463,N_9065);
nand U14997 (N_14997,N_7893,N_6595);
and U14998 (N_14998,N_7343,N_5352);
xnor U14999 (N_14999,N_5580,N_6153);
and U15000 (N_15000,N_10756,N_13843);
nor U15001 (N_15001,N_10885,N_13709);
xor U15002 (N_15002,N_10351,N_14583);
and U15003 (N_15003,N_13463,N_12199);
xnor U15004 (N_15004,N_10370,N_11771);
nor U15005 (N_15005,N_12063,N_14021);
and U15006 (N_15006,N_14491,N_13179);
and U15007 (N_15007,N_11182,N_10889);
nand U15008 (N_15008,N_13110,N_10219);
and U15009 (N_15009,N_12369,N_13829);
xor U15010 (N_15010,N_10625,N_13538);
nor U15011 (N_15011,N_12992,N_11782);
xnor U15012 (N_15012,N_14991,N_14635);
nand U15013 (N_15013,N_13044,N_13899);
nor U15014 (N_15014,N_13532,N_14143);
nand U15015 (N_15015,N_14729,N_13125);
nand U15016 (N_15016,N_14405,N_11750);
nor U15017 (N_15017,N_13957,N_10311);
nor U15018 (N_15018,N_13119,N_14339);
xor U15019 (N_15019,N_11339,N_14736);
nand U15020 (N_15020,N_14528,N_10528);
or U15021 (N_15021,N_11699,N_11094);
or U15022 (N_15022,N_13702,N_12153);
xor U15023 (N_15023,N_11131,N_11362);
or U15024 (N_15024,N_10613,N_13336);
nor U15025 (N_15025,N_14937,N_10247);
or U15026 (N_15026,N_12714,N_10531);
nor U15027 (N_15027,N_12514,N_11395);
or U15028 (N_15028,N_12581,N_12543);
nor U15029 (N_15029,N_10192,N_10439);
or U15030 (N_15030,N_12549,N_13235);
xnor U15031 (N_15031,N_12462,N_11388);
xnor U15032 (N_15032,N_14778,N_11296);
nand U15033 (N_15033,N_14306,N_10884);
nand U15034 (N_15034,N_10555,N_10113);
and U15035 (N_15035,N_11817,N_13672);
or U15036 (N_15036,N_13715,N_11382);
and U15037 (N_15037,N_10600,N_14199);
nor U15038 (N_15038,N_10206,N_10424);
nand U15039 (N_15039,N_10903,N_11040);
nand U15040 (N_15040,N_11862,N_11334);
nor U15041 (N_15041,N_12646,N_13258);
xor U15042 (N_15042,N_10389,N_13846);
or U15043 (N_15043,N_14412,N_14332);
nor U15044 (N_15044,N_11289,N_14803);
xnor U15045 (N_15045,N_12840,N_13568);
nand U15046 (N_15046,N_14419,N_10794);
or U15047 (N_15047,N_10569,N_13601);
or U15048 (N_15048,N_12511,N_11744);
or U15049 (N_15049,N_14890,N_12558);
xor U15050 (N_15050,N_11082,N_11530);
and U15051 (N_15051,N_14426,N_11555);
and U15052 (N_15052,N_14063,N_13143);
or U15053 (N_15053,N_10190,N_14791);
xor U15054 (N_15054,N_14741,N_11413);
or U15055 (N_15055,N_12267,N_14107);
and U15056 (N_15056,N_12134,N_14847);
xnor U15057 (N_15057,N_13060,N_12707);
nor U15058 (N_15058,N_14660,N_13832);
nor U15059 (N_15059,N_13640,N_14216);
and U15060 (N_15060,N_13885,N_10633);
nor U15061 (N_15061,N_12172,N_13091);
xnor U15062 (N_15062,N_13623,N_12455);
and U15063 (N_15063,N_11251,N_14866);
nand U15064 (N_15064,N_14254,N_14687);
nor U15065 (N_15065,N_12734,N_10754);
nand U15066 (N_15066,N_10287,N_14919);
xnor U15067 (N_15067,N_11481,N_12588);
nor U15068 (N_15068,N_11735,N_12784);
xnor U15069 (N_15069,N_10760,N_13276);
xnor U15070 (N_15070,N_12483,N_14764);
and U15071 (N_15071,N_13561,N_10355);
xnor U15072 (N_15072,N_13114,N_12246);
or U15073 (N_15073,N_13969,N_11150);
and U15074 (N_15074,N_10014,N_10841);
xor U15075 (N_15075,N_14158,N_11820);
or U15076 (N_15076,N_11965,N_11090);
xor U15077 (N_15077,N_14353,N_14561);
or U15078 (N_15078,N_10980,N_12421);
xor U15079 (N_15079,N_12275,N_10874);
xor U15080 (N_15080,N_12896,N_10144);
or U15081 (N_15081,N_11327,N_12539);
or U15082 (N_15082,N_11857,N_11297);
xor U15083 (N_15083,N_14577,N_13577);
nand U15084 (N_15084,N_14886,N_13901);
nor U15085 (N_15085,N_11140,N_11153);
nand U15086 (N_15086,N_14206,N_13933);
xnor U15087 (N_15087,N_13854,N_10791);
nor U15088 (N_15088,N_11147,N_13196);
nand U15089 (N_15089,N_11952,N_11762);
xor U15090 (N_15090,N_12047,N_10130);
xor U15091 (N_15091,N_10267,N_13612);
xnor U15092 (N_15092,N_12485,N_13681);
nor U15093 (N_15093,N_12092,N_11126);
nor U15094 (N_15094,N_13663,N_12750);
nand U15095 (N_15095,N_13657,N_14275);
nor U15096 (N_15096,N_11637,N_12264);
nand U15097 (N_15097,N_13037,N_14065);
xor U15098 (N_15098,N_10111,N_10009);
xor U15099 (N_15099,N_13820,N_12522);
or U15100 (N_15100,N_14915,N_13491);
nor U15101 (N_15101,N_12472,N_10728);
and U15102 (N_15102,N_14361,N_13948);
and U15103 (N_15103,N_14105,N_14551);
or U15104 (N_15104,N_13708,N_12062);
or U15105 (N_15105,N_13731,N_13874);
nand U15106 (N_15106,N_14864,N_13941);
or U15107 (N_15107,N_14467,N_11397);
nand U15108 (N_15108,N_11989,N_13878);
xor U15109 (N_15109,N_13231,N_11770);
nand U15110 (N_15110,N_12351,N_10087);
or U15111 (N_15111,N_11858,N_12510);
nor U15112 (N_15112,N_11874,N_10145);
xnor U15113 (N_15113,N_12247,N_13599);
or U15114 (N_15114,N_14322,N_14940);
and U15115 (N_15115,N_12290,N_12139);
nand U15116 (N_15116,N_12637,N_10747);
or U15117 (N_15117,N_14975,N_14670);
xnor U15118 (N_15118,N_14544,N_10753);
or U15119 (N_15119,N_10392,N_10184);
or U15120 (N_15120,N_13747,N_10844);
nand U15121 (N_15121,N_14377,N_10133);
and U15122 (N_15122,N_12097,N_14389);
and U15123 (N_15123,N_12829,N_14028);
nand U15124 (N_15124,N_13081,N_13535);
nand U15125 (N_15125,N_10007,N_10979);
nor U15126 (N_15126,N_10568,N_10049);
or U15127 (N_15127,N_12778,N_14747);
nand U15128 (N_15128,N_12149,N_10292);
and U15129 (N_15129,N_14235,N_14617);
nand U15130 (N_15130,N_12959,N_14448);
nand U15131 (N_15131,N_10989,N_10000);
nor U15132 (N_15132,N_13668,N_13860);
nor U15133 (N_15133,N_10615,N_11706);
and U15134 (N_15134,N_14769,N_11093);
or U15135 (N_15135,N_13790,N_10911);
nor U15136 (N_15136,N_13513,N_12739);
nor U15137 (N_15137,N_12673,N_12403);
and U15138 (N_15138,N_10935,N_10254);
or U15139 (N_15139,N_14980,N_11004);
nor U15140 (N_15140,N_11642,N_12001);
xnor U15141 (N_15141,N_14304,N_13711);
xnor U15142 (N_15142,N_12185,N_14809);
nand U15143 (N_15143,N_11423,N_14329);
and U15144 (N_15144,N_10385,N_13457);
nor U15145 (N_15145,N_13597,N_14810);
nor U15146 (N_15146,N_14030,N_14900);
nor U15147 (N_15147,N_13862,N_12426);
nand U15148 (N_15148,N_13682,N_11483);
nand U15149 (N_15149,N_10800,N_12453);
xor U15150 (N_15150,N_13382,N_13685);
xor U15151 (N_15151,N_14870,N_12947);
nand U15152 (N_15152,N_10418,N_10153);
nand U15153 (N_15153,N_11134,N_11578);
or U15154 (N_15154,N_12123,N_13507);
nor U15155 (N_15155,N_10922,N_11176);
or U15156 (N_15156,N_13321,N_13815);
and U15157 (N_15157,N_11472,N_13710);
nand U15158 (N_15158,N_12838,N_10458);
and U15159 (N_15159,N_10305,N_12442);
and U15160 (N_15160,N_13281,N_10624);
xnor U15161 (N_15161,N_14058,N_14050);
nand U15162 (N_15162,N_13920,N_14044);
nand U15163 (N_15163,N_14182,N_12484);
or U15164 (N_15164,N_13480,N_12361);
nor U15165 (N_15165,N_10450,N_12937);
xor U15166 (N_15166,N_13377,N_14618);
nor U15167 (N_15167,N_11677,N_12336);
nand U15168 (N_15168,N_12254,N_14212);
and U15169 (N_15169,N_14923,N_12690);
or U15170 (N_15170,N_10508,N_12265);
nor U15171 (N_15171,N_12043,N_14625);
and U15172 (N_15172,N_10557,N_10428);
nor U15173 (N_15173,N_14939,N_14394);
or U15174 (N_15174,N_13869,N_14409);
nor U15175 (N_15175,N_10805,N_14424);
and U15176 (N_15176,N_10835,N_14961);
or U15177 (N_15177,N_10647,N_11162);
nor U15178 (N_15178,N_11737,N_12632);
and U15179 (N_15179,N_12626,N_10606);
or U15180 (N_15180,N_12732,N_11001);
nand U15181 (N_15181,N_13550,N_13900);
nand U15182 (N_15182,N_10224,N_14237);
xor U15183 (N_15183,N_13266,N_13922);
or U15184 (N_15184,N_10100,N_13896);
or U15185 (N_15185,N_13588,N_14090);
nor U15186 (N_15186,N_14689,N_14996);
nand U15187 (N_15187,N_12885,N_12441);
nand U15188 (N_15188,N_10055,N_11166);
and U15189 (N_15189,N_10533,N_13230);
xnor U15190 (N_15190,N_10988,N_11864);
or U15191 (N_15191,N_13775,N_13355);
xnor U15192 (N_15192,N_10412,N_10630);
nor U15193 (N_15193,N_14250,N_11047);
or U15194 (N_15194,N_13489,N_12644);
or U15195 (N_15195,N_12533,N_13012);
nand U15196 (N_15196,N_13564,N_14648);
nor U15197 (N_15197,N_12180,N_14624);
nor U15198 (N_15198,N_14367,N_13644);
and U15199 (N_15199,N_11235,N_13741);
nor U15200 (N_15200,N_11003,N_14166);
or U15201 (N_15201,N_14461,N_11427);
xor U15202 (N_15202,N_12866,N_12924);
and U15203 (N_15203,N_12518,N_12119);
xnor U15204 (N_15204,N_11139,N_11630);
xor U15205 (N_15205,N_13593,N_13186);
xnor U15206 (N_15206,N_11037,N_13939);
nand U15207 (N_15207,N_10715,N_13079);
nand U15208 (N_15208,N_11160,N_13793);
xnor U15209 (N_15209,N_11676,N_11077);
nor U15210 (N_15210,N_14234,N_13766);
xnor U15211 (N_15211,N_14944,N_14278);
and U15212 (N_15212,N_13773,N_12118);
nand U15213 (N_15213,N_11211,N_14557);
or U15214 (N_15214,N_10442,N_13866);
and U15215 (N_15215,N_13157,N_13462);
nor U15216 (N_15216,N_13581,N_11400);
xor U15217 (N_15217,N_13752,N_10478);
nor U15218 (N_15218,N_13032,N_14533);
nand U15219 (N_15219,N_10675,N_12691);
and U15220 (N_15220,N_11100,N_11880);
or U15221 (N_15221,N_11316,N_12024);
xor U15222 (N_15222,N_12033,N_11931);
nand U15223 (N_15223,N_14117,N_14153);
and U15224 (N_15224,N_10829,N_11691);
nor U15225 (N_15225,N_10086,N_10734);
xor U15226 (N_15226,N_13147,N_11405);
nor U15227 (N_15227,N_13592,N_13774);
xnor U15228 (N_15228,N_13048,N_13465);
and U15229 (N_15229,N_14674,N_13019);
xnor U15230 (N_15230,N_11921,N_13995);
and U15231 (N_15231,N_10063,N_13735);
nand U15232 (N_15232,N_11967,N_13097);
xor U15233 (N_15233,N_12210,N_10899);
or U15234 (N_15234,N_14497,N_12125);
xor U15235 (N_15235,N_13796,N_14756);
and U15236 (N_15236,N_14362,N_12618);
xnor U15237 (N_15237,N_13436,N_10107);
nor U15238 (N_15238,N_14701,N_14602);
nand U15239 (N_15239,N_11407,N_10880);
nand U15240 (N_15240,N_13460,N_14694);
nand U15241 (N_15241,N_14225,N_12716);
xor U15242 (N_15242,N_13646,N_11070);
or U15243 (N_15243,N_10148,N_13419);
and U15244 (N_15244,N_13971,N_14507);
nand U15245 (N_15245,N_13270,N_11018);
or U15246 (N_15246,N_10785,N_10214);
nor U15247 (N_15247,N_12585,N_14502);
or U15248 (N_15248,N_10310,N_11611);
xnor U15249 (N_15249,N_14781,N_10853);
nor U15250 (N_15250,N_14043,N_11071);
or U15251 (N_15251,N_14775,N_14321);
nor U15252 (N_15252,N_11619,N_14675);
nand U15253 (N_15253,N_11463,N_13030);
and U15254 (N_15254,N_13686,N_13596);
nor U15255 (N_15255,N_10406,N_11268);
and U15256 (N_15256,N_11743,N_13403);
or U15257 (N_15257,N_13085,N_14818);
nor U15258 (N_15258,N_11475,N_12622);
nand U15259 (N_15259,N_11519,N_10912);
nor U15260 (N_15260,N_14718,N_10462);
nand U15261 (N_15261,N_12423,N_14435);
and U15262 (N_15262,N_13968,N_13442);
and U15263 (N_15263,N_13853,N_14941);
nand U15264 (N_15264,N_12635,N_13055);
nor U15265 (N_15265,N_13805,N_14655);
and U15266 (N_15266,N_13603,N_13637);
xnor U15267 (N_15267,N_10187,N_13486);
and U15268 (N_15268,N_13456,N_11261);
nand U15269 (N_15269,N_12771,N_10875);
and U15270 (N_15270,N_12841,N_11119);
nand U15271 (N_15271,N_11640,N_10654);
nand U15272 (N_15272,N_13046,N_11972);
nor U15273 (N_15273,N_10347,N_14416);
nand U15274 (N_15274,N_11133,N_10270);
or U15275 (N_15275,N_12542,N_12295);
xor U15276 (N_15276,N_11746,N_14100);
nand U15277 (N_15277,N_14956,N_12934);
xnor U15278 (N_15278,N_14962,N_12531);
xor U15279 (N_15279,N_12650,N_13988);
or U15280 (N_15280,N_13958,N_10317);
and U15281 (N_15281,N_11883,N_12861);
xnor U15282 (N_15282,N_11391,N_11184);
xnor U15283 (N_15283,N_12002,N_11513);
and U15284 (N_15284,N_13387,N_10601);
nand U15285 (N_15285,N_11249,N_11204);
xor U15286 (N_15286,N_11978,N_13288);
nand U15287 (N_15287,N_14516,N_12614);
or U15288 (N_15288,N_12174,N_10904);
nor U15289 (N_15289,N_10376,N_13673);
nor U15290 (N_15290,N_14280,N_14536);
or U15291 (N_15291,N_12687,N_13575);
or U15292 (N_15292,N_10906,N_10264);
or U15293 (N_15293,N_14372,N_10393);
nor U15294 (N_15294,N_10871,N_13088);
or U15295 (N_15295,N_14464,N_14255);
and U15296 (N_15296,N_14925,N_14802);
nand U15297 (N_15297,N_10650,N_14668);
nand U15298 (N_15298,N_12479,N_13689);
xnor U15299 (N_15299,N_10218,N_11084);
nand U15300 (N_15300,N_10030,N_14676);
xor U15301 (N_15301,N_14553,N_14401);
nand U15302 (N_15302,N_12516,N_10188);
or U15303 (N_15303,N_10448,N_10474);
nor U15304 (N_15304,N_12034,N_13608);
xnor U15305 (N_15305,N_12284,N_14559);
or U15306 (N_15306,N_11164,N_12820);
xor U15307 (N_15307,N_14159,N_13177);
nand U15308 (N_15308,N_12330,N_12638);
nand U15309 (N_15309,N_14513,N_13667);
nand U15310 (N_15310,N_13054,N_11764);
nand U15311 (N_15311,N_10806,N_10686);
and U15312 (N_15312,N_10269,N_13831);
xnor U15313 (N_15313,N_13063,N_14252);
nand U15314 (N_15314,N_10337,N_14721);
and U15315 (N_15315,N_11384,N_11650);
nand U15316 (N_15316,N_11955,N_14338);
xnor U15317 (N_15317,N_14728,N_14584);
xor U15318 (N_15318,N_12584,N_11969);
and U15319 (N_15319,N_14860,N_12923);
or U15320 (N_15320,N_11503,N_12740);
nand U15321 (N_15321,N_10781,N_13569);
nand U15322 (N_15322,N_12309,N_10599);
nor U15323 (N_15323,N_14201,N_11048);
or U15324 (N_15324,N_10236,N_10037);
nand U15325 (N_15325,N_12713,N_10639);
nor U15326 (N_15326,N_10986,N_14546);
xnor U15327 (N_15327,N_10937,N_10154);
or U15328 (N_15328,N_11656,N_11390);
and U15329 (N_15329,N_13523,N_12057);
xnor U15330 (N_15330,N_14512,N_13943);
or U15331 (N_15331,N_10809,N_13051);
nand U15332 (N_15332,N_10350,N_14759);
and U15333 (N_15333,N_10250,N_11023);
nor U15334 (N_15334,N_10585,N_14270);
nand U15335 (N_15335,N_13289,N_11345);
nor U15336 (N_15336,N_10976,N_13803);
or U15337 (N_15337,N_12494,N_13424);
xor U15338 (N_15338,N_13554,N_10066);
or U15339 (N_15339,N_10421,N_12268);
and U15340 (N_15340,N_14938,N_14430);
and U15341 (N_15341,N_10916,N_11507);
nand U15342 (N_15342,N_11024,N_11977);
or U15343 (N_15343,N_10080,N_11039);
nor U15344 (N_15344,N_12094,N_11891);
nand U15345 (N_15345,N_11347,N_11659);
nor U15346 (N_15346,N_12320,N_11794);
nand U15347 (N_15347,N_13703,N_13806);
nand U15348 (N_15348,N_12223,N_12017);
nor U15349 (N_15349,N_11922,N_13049);
and U15350 (N_15350,N_13680,N_14171);
or U15351 (N_15351,N_14745,N_11085);
or U15352 (N_15352,N_13771,N_14977);
nand U15353 (N_15353,N_14592,N_10238);
xnor U15354 (N_15354,N_10091,N_14629);
nor U15355 (N_15355,N_11736,N_11151);
nand U15356 (N_15356,N_11915,N_10044);
or U15357 (N_15357,N_10352,N_11343);
and U15358 (N_15358,N_10258,N_13407);
and U15359 (N_15359,N_11492,N_14814);
nor U15360 (N_15360,N_14197,N_14754);
nor U15361 (N_15361,N_12813,N_10076);
nor U15362 (N_15362,N_14150,N_10408);
or U15363 (N_15363,N_11042,N_13718);
or U15364 (N_15364,N_14328,N_11527);
and U15365 (N_15365,N_13065,N_14333);
and U15366 (N_15366,N_10172,N_14859);
nand U15367 (N_15367,N_13763,N_12520);
and U15368 (N_15368,N_12151,N_13622);
and U15369 (N_15369,N_13053,N_14499);
nand U15370 (N_15370,N_10028,N_14608);
or U15371 (N_15371,N_11130,N_12911);
or U15372 (N_15372,N_10543,N_10381);
nand U15373 (N_15373,N_12234,N_11315);
nor U15374 (N_15374,N_11846,N_14589);
nand U15375 (N_15375,N_11775,N_11239);
or U15376 (N_15376,N_13616,N_12828);
xor U15377 (N_15377,N_10354,N_12277);
or U15378 (N_15378,N_14738,N_11686);
nor U15379 (N_15379,N_12743,N_12724);
and U15380 (N_15380,N_13068,N_12791);
nand U15381 (N_15381,N_14111,N_11063);
nor U15382 (N_15382,N_12827,N_13497);
xnor U15383 (N_15383,N_10598,N_10490);
and U15384 (N_15384,N_13565,N_13203);
and U15385 (N_15385,N_14796,N_12083);
and U15386 (N_15386,N_13183,N_10170);
or U15387 (N_15387,N_12831,N_12972);
and U15388 (N_15388,N_14342,N_11299);
or U15389 (N_15389,N_14952,N_13440);
nor U15390 (N_15390,N_12435,N_12948);
or U15391 (N_15391,N_11592,N_13524);
or U15392 (N_15392,N_11687,N_12766);
and U15393 (N_15393,N_11038,N_14683);
xor U15394 (N_15394,N_11311,N_14433);
xnor U15395 (N_15395,N_11823,N_14354);
nand U15396 (N_15396,N_10115,N_11020);
xnor U15397 (N_15397,N_11072,N_12376);
or U15398 (N_15398,N_10366,N_14135);
nor U15399 (N_15399,N_10484,N_14834);
nand U15400 (N_15400,N_13376,N_12221);
nor U15401 (N_15401,N_13340,N_13039);
nand U15402 (N_15402,N_10331,N_14165);
nand U15403 (N_15403,N_12075,N_12767);
nor U15404 (N_15404,N_11776,N_10147);
nand U15405 (N_15405,N_12301,N_10592);
and U15406 (N_15406,N_11228,N_12940);
nor U15407 (N_15407,N_14990,N_11055);
xnor U15408 (N_15408,N_13433,N_14478);
and U15409 (N_15409,N_13986,N_14060);
and U15410 (N_15410,N_11121,N_11425);
nor U15411 (N_15411,N_10482,N_10577);
xnor U15412 (N_15412,N_11052,N_13865);
nor U15413 (N_15413,N_14669,N_10194);
or U15414 (N_15414,N_11387,N_14772);
and U15415 (N_15415,N_12708,N_10517);
nand U15416 (N_15416,N_14612,N_14119);
nor U15417 (N_15417,N_11236,N_11950);
nor U15418 (N_15418,N_12787,N_11000);
nand U15419 (N_15419,N_11168,N_10620);
or U15420 (N_15420,N_14080,N_10710);
nor U15421 (N_15421,N_14875,N_10672);
nor U15422 (N_15422,N_14316,N_10023);
or U15423 (N_15423,N_10438,N_10960);
nand U15424 (N_15424,N_12244,N_14174);
nor U15425 (N_15425,N_11994,N_10053);
nor U15426 (N_15426,N_13745,N_12852);
nor U15427 (N_15427,N_10914,N_13252);
xnor U15428 (N_15428,N_12572,N_11342);
or U15429 (N_15429,N_11470,N_11692);
nor U15430 (N_15430,N_13259,N_11783);
and U15431 (N_15431,N_12981,N_11396);
xnor U15432 (N_15432,N_10266,N_11103);
or U15433 (N_15433,N_13003,N_12365);
or U15434 (N_15434,N_13607,N_11313);
or U15435 (N_15435,N_13814,N_10711);
nor U15436 (N_15436,N_13164,N_12915);
nor U15437 (N_15437,N_10363,N_10578);
nor U15438 (N_15438,N_14138,N_14423);
or U15439 (N_15439,N_10658,N_12375);
or U15440 (N_15440,N_13635,N_12647);
or U15441 (N_15441,N_12762,N_13522);
nor U15442 (N_15442,N_12414,N_14903);
and U15443 (N_15443,N_11559,N_13776);
nand U15444 (N_15444,N_11981,N_10099);
or U15445 (N_15445,N_12240,N_10648);
and U15446 (N_15446,N_14352,N_12907);
nand U15447 (N_15447,N_13734,N_11172);
or U15448 (N_15448,N_12832,N_10391);
and U15449 (N_15449,N_14698,N_11460);
or U15450 (N_15450,N_11214,N_12854);
nor U15451 (N_15451,N_10205,N_12956);
or U15452 (N_15452,N_13950,N_14189);
nor U15453 (N_15453,N_13166,N_11041);
nor U15454 (N_15454,N_12991,N_12817);
nor U15455 (N_15455,N_11163,N_14872);
and U15456 (N_15456,N_13954,N_10560);
nand U15457 (N_15457,N_10280,N_12082);
nor U15458 (N_15458,N_14901,N_12283);
nand U15459 (N_15459,N_10545,N_14274);
nor U15460 (N_15460,N_12974,N_12067);
or U15461 (N_15461,N_14750,N_11127);
nor U15462 (N_15462,N_12860,N_10792);
nand U15463 (N_15463,N_10384,N_13562);
xnor U15464 (N_15464,N_14432,N_12855);
nand U15465 (N_15465,N_13979,N_12906);
xor U15466 (N_15466,N_10741,N_11141);
or U15467 (N_15467,N_11837,N_11801);
nor U15468 (N_15468,N_13791,N_12238);
xor U15469 (N_15469,N_10234,N_14636);
nand U15470 (N_15470,N_11361,N_11717);
and U15471 (N_15471,N_12355,N_14102);
or U15472 (N_15472,N_14692,N_14605);
or U15473 (N_15473,N_12977,N_13529);
nand U15474 (N_15474,N_10451,N_10525);
nor U15475 (N_15475,N_12348,N_14018);
nand U15476 (N_15476,N_12916,N_11542);
nor U15477 (N_15477,N_14881,N_10553);
xnor U15478 (N_15478,N_10325,N_13617);
nand U15479 (N_15479,N_14783,N_10059);
or U15480 (N_15480,N_10436,N_13794);
nor U15481 (N_15481,N_13017,N_10021);
nor U15482 (N_15482,N_10567,N_11802);
and U15483 (N_15483,N_11830,N_10036);
and U15484 (N_15484,N_11383,N_11282);
nand U15485 (N_15485,N_10597,N_14285);
and U15486 (N_15486,N_10471,N_12932);
xor U15487 (N_15487,N_11262,N_10073);
nor U15488 (N_15488,N_11497,N_12010);
and U15489 (N_15489,N_10182,N_10410);
or U15490 (N_15490,N_12390,N_12115);
nor U15491 (N_15491,N_10725,N_13301);
or U15492 (N_15492,N_12278,N_12220);
nor U15493 (N_15493,N_13571,N_11923);
xor U15494 (N_15494,N_14661,N_14765);
or U15495 (N_15495,N_12798,N_13662);
or U15496 (N_15496,N_11192,N_14148);
or U15497 (N_15497,N_12312,N_12368);
nand U15498 (N_15498,N_11199,N_12102);
xor U15499 (N_15499,N_10973,N_13792);
nor U15500 (N_15500,N_14838,N_10285);
nand U15501 (N_15501,N_12830,N_10819);
or U15502 (N_15502,N_13543,N_13824);
xor U15503 (N_15503,N_14906,N_11335);
nand U15504 (N_15504,N_11144,N_14717);
nand U15505 (N_15505,N_10265,N_10727);
or U15506 (N_15506,N_13346,N_10290);
nand U15507 (N_15507,N_13921,N_14904);
xor U15508 (N_15508,N_13488,N_14703);
nand U15509 (N_15509,N_14438,N_11909);
and U15510 (N_15510,N_14400,N_13432);
and U15511 (N_15511,N_10836,N_13624);
xnor U15512 (N_15512,N_11450,N_13202);
and U15513 (N_15513,N_11326,N_14852);
or U15514 (N_15514,N_14204,N_12819);
nand U15515 (N_15515,N_12920,N_12568);
nor U15516 (N_15516,N_12634,N_14017);
nand U15517 (N_15517,N_10564,N_12961);
nor U15518 (N_15518,N_14310,N_12664);
nor U15519 (N_15519,N_10975,N_14064);
and U15520 (N_15520,N_10343,N_11137);
nor U15521 (N_15521,N_10019,N_14287);
nand U15522 (N_15522,N_13674,N_11627);
nand U15523 (N_15523,N_14309,N_14585);
and U15524 (N_15524,N_14567,N_10169);
or U15525 (N_15525,N_12107,N_10126);
nor U15526 (N_15526,N_10649,N_14193);
nor U15527 (N_15527,N_10983,N_12280);
nand U15528 (N_15528,N_13122,N_10535);
or U15529 (N_15529,N_10892,N_14542);
and U15530 (N_15530,N_10752,N_11095);
nor U15531 (N_15531,N_11919,N_13071);
and U15532 (N_15532,N_12438,N_13422);
nand U15533 (N_15533,N_13169,N_12938);
nor U15534 (N_15534,N_12219,N_11803);
nor U15535 (N_15535,N_13176,N_10397);
or U15536 (N_15536,N_10197,N_11813);
nand U15537 (N_15537,N_14848,N_13572);
nor U15538 (N_15538,N_12926,N_14632);
or U15539 (N_15539,N_10958,N_13427);
nor U15540 (N_15540,N_10498,N_13881);
or U15541 (N_15541,N_11835,N_11789);
nand U15542 (N_15542,N_13325,N_12945);
nand U15543 (N_15543,N_12500,N_11793);
and U15544 (N_15544,N_12676,N_13391);
nor U15545 (N_15545,N_10129,N_14790);
or U15546 (N_15546,N_10621,N_12880);
and U15547 (N_15547,N_10622,N_13928);
nand U15548 (N_15548,N_11845,N_12371);
nor U15549 (N_15549,N_12835,N_11537);
nand U15550 (N_15550,N_11748,N_10463);
or U15551 (N_15551,N_13319,N_14829);
nand U15552 (N_15552,N_14957,N_11376);
xor U15553 (N_15553,N_12731,N_13078);
xor U15554 (N_15554,N_12587,N_10882);
nor U15555 (N_15555,N_11713,N_10309);
and U15556 (N_15556,N_10472,N_10608);
xnor U15557 (N_15557,N_12755,N_13330);
xor U15558 (N_15558,N_11979,N_12717);
nand U15559 (N_15559,N_14682,N_14458);
nand U15560 (N_15560,N_10870,N_12066);
nor U15561 (N_15561,N_11859,N_13728);
or U15562 (N_15562,N_13485,N_13251);
nand U15563 (N_15563,N_10681,N_14973);
xor U15564 (N_15564,N_12196,N_13908);
xor U15565 (N_15565,N_10510,N_11428);
nor U15566 (N_15566,N_13691,N_12544);
xnor U15567 (N_15567,N_13213,N_10824);
and U15568 (N_15568,N_14659,N_12398);
nor U15569 (N_15569,N_12499,N_10859);
nor U15570 (N_15570,N_12446,N_13438);
or U15571 (N_15571,N_10720,N_10796);
or U15572 (N_15572,N_13292,N_11125);
and U15573 (N_15573,N_11487,N_10749);
xnor U15574 (N_15574,N_14690,N_11987);
or U15575 (N_15575,N_11796,N_12537);
nand U15576 (N_15576,N_14096,N_14792);
and U15577 (N_15577,N_12271,N_14263);
nand U15578 (N_15578,N_12143,N_14773);
nand U15579 (N_15579,N_10972,N_10358);
and U15580 (N_15580,N_10619,N_11157);
nor U15581 (N_15581,N_11563,N_12122);
nor U15582 (N_15582,N_12085,N_10420);
xnor U15583 (N_15583,N_11220,N_12208);
nand U15584 (N_15584,N_10561,N_13219);
and U15585 (N_15585,N_14651,N_12228);
and U15586 (N_15586,N_12593,N_11516);
and U15587 (N_15587,N_14606,N_14112);
or U15588 (N_15588,N_13395,N_10175);
xor U15589 (N_15589,N_11218,N_14637);
xor U15590 (N_15590,N_13089,N_12670);
and U15591 (N_15591,N_14249,N_13742);
nand U15592 (N_15592,N_11572,N_10645);
nor U15593 (N_15593,N_13841,N_14262);
nand U15594 (N_15594,N_14920,N_10344);
and U15595 (N_15595,N_12073,N_11673);
nor U15596 (N_15596,N_10118,N_11581);
and U15597 (N_15597,N_13415,N_13857);
or U15598 (N_15598,N_13156,N_14855);
and U15599 (N_15599,N_10762,N_10237);
and U15600 (N_15600,N_14621,N_10540);
xor U15601 (N_15601,N_11855,N_13953);
xor U15602 (N_15602,N_14878,N_13073);
nand U15603 (N_15603,N_12856,N_13898);
nand U15604 (N_15604,N_12399,N_14428);
and U15605 (N_15605,N_14897,N_10295);
or U15606 (N_15606,N_12400,N_10057);
or U15607 (N_15607,N_10038,N_11643);
xor U15608 (N_15608,N_13494,N_14246);
and U15609 (N_15609,N_12296,N_14994);
and U15610 (N_15610,N_14645,N_12718);
and U15611 (N_15611,N_13915,N_13113);
xnor U15612 (N_15612,N_13548,N_11745);
nand U15613 (N_15613,N_10936,N_11876);
nand U15614 (N_15614,N_14281,N_14843);
nand U15615 (N_15615,N_12627,N_10627);
nor U15616 (N_15616,N_10283,N_11323);
xor U15617 (N_15617,N_10365,N_12513);
nor U15618 (N_15618,N_13779,N_14898);
and U15619 (N_15619,N_11740,N_10893);
xnor U15620 (N_15620,N_13653,N_14313);
and U15621 (N_15621,N_12667,N_13220);
or U15622 (N_15622,N_10128,N_10709);
xnor U15623 (N_15623,N_11509,N_12857);
xor U15624 (N_15624,N_12954,N_13557);
or U15625 (N_15625,N_11320,N_13595);
or U15626 (N_15626,N_11523,N_13525);
xnor U15627 (N_15627,N_11658,N_10163);
nand U15628 (N_15628,N_13590,N_11393);
xnor U15629 (N_15629,N_11426,N_14515);
xnor U15630 (N_15630,N_10167,N_13328);
nor U15631 (N_15631,N_10783,N_14439);
xor U15632 (N_15632,N_11216,N_12715);
and U15633 (N_15633,N_10114,N_10594);
nand U15634 (N_15634,N_12357,N_14345);
nor U15635 (N_15635,N_11732,N_12582);
nand U15636 (N_15636,N_14200,N_13347);
or U15637 (N_15637,N_12931,N_12205);
nor U15638 (N_15638,N_11062,N_12019);
or U15639 (N_15639,N_10558,N_13938);
or U15640 (N_15640,N_10908,N_10150);
and U15641 (N_15641,N_12826,N_10767);
nor U15642 (N_15642,N_13309,N_14633);
nor U15643 (N_15643,N_10616,N_11544);
xor U15644 (N_15644,N_13082,N_10079);
xor U15645 (N_15645,N_12668,N_11068);
xor U15646 (N_15646,N_12029,N_11797);
xnor U15647 (N_15647,N_14959,N_14794);
nor U15648 (N_15648,N_12255,N_14187);
nand U15649 (N_15649,N_12100,N_11392);
nand U15650 (N_15650,N_14614,N_10307);
nor U15651 (N_15651,N_11193,N_14290);
nor U15652 (N_15652,N_14217,N_14051);
xor U15653 (N_15653,N_11406,N_10953);
nand U15654 (N_15654,N_13945,N_13947);
nor U15655 (N_15655,N_12616,N_14654);
xor U15656 (N_15656,N_11791,N_13993);
nand U15657 (N_15657,N_13275,N_12628);
nand U15658 (N_15658,N_11074,N_13660);
xor U15659 (N_15659,N_12927,N_11580);
xnor U15660 (N_15660,N_12525,N_14550);
nand U15661 (N_15661,N_12741,N_10232);
xnor U15662 (N_15662,N_11107,N_12144);
and U15663 (N_15663,N_10158,N_10010);
nand U15664 (N_15664,N_13631,N_10298);
xnor U15665 (N_15665,N_10159,N_11248);
and U15666 (N_15666,N_14895,N_12729);
or U15667 (N_15667,N_13837,N_11625);
nor U15668 (N_15668,N_14541,N_10708);
or U15669 (N_15669,N_14876,N_14243);
xnor U15670 (N_15670,N_12349,N_10348);
xor U15671 (N_15671,N_12359,N_12132);
and U15672 (N_15672,N_10361,N_11571);
and U15673 (N_15673,N_13926,N_10810);
or U15674 (N_15674,N_11720,N_10222);
and U15675 (N_15675,N_13714,N_12150);
or U15676 (N_15676,N_14381,N_11598);
and U15677 (N_15677,N_11447,N_10766);
nor U15678 (N_15678,N_12055,N_10769);
xnor U15679 (N_15679,N_13705,N_11990);
xor U15680 (N_15680,N_10514,N_12846);
and U15681 (N_15681,N_10486,N_11456);
xnor U15682 (N_15682,N_11462,N_12074);
or U15683 (N_15683,N_10587,N_12410);
nand U15684 (N_15684,N_10475,N_11324);
xor U15685 (N_15685,N_12570,N_11778);
nand U15686 (N_15686,N_12261,N_13470);
nor U15687 (N_15687,N_12674,N_14232);
nor U15688 (N_15688,N_13855,N_13828);
or U15689 (N_15689,N_14213,N_11645);
nor U15690 (N_15690,N_11493,N_12432);
or U15691 (N_15691,N_10541,N_12710);
nand U15692 (N_15692,N_14315,N_10586);
nand U15693 (N_15693,N_11269,N_13658);
nand U15694 (N_15694,N_14770,N_11329);
nand U15695 (N_15695,N_10330,N_10656);
nor U15696 (N_15696,N_13040,N_14179);
nand U15697 (N_15697,N_11305,N_14302);
and U15698 (N_15698,N_11303,N_11132);
nand U15699 (N_15699,N_10511,N_10689);
nor U15700 (N_15700,N_12580,N_12901);
xnor U15701 (N_15701,N_14344,N_13620);
xor U15702 (N_15702,N_12209,N_14390);
and U15703 (N_15703,N_12407,N_10524);
and U15704 (N_15704,N_13699,N_14469);
xor U15705 (N_15705,N_14145,N_12988);
nand U15706 (N_15706,N_10626,N_11622);
and U15707 (N_15707,N_12428,N_13772);
or U15708 (N_15708,N_14454,N_11246);
nand U15709 (N_15709,N_14334,N_13573);
xnor U15710 (N_15710,N_10349,N_12893);
and U15711 (N_15711,N_13002,N_10926);
and U15712 (N_15712,N_14788,N_12697);
nand U15713 (N_15713,N_11540,N_14523);
nor U15714 (N_15714,N_12166,N_10174);
xor U15715 (N_15715,N_14514,N_12025);
or U15716 (N_15716,N_11946,N_14760);
xor U15717 (N_15717,N_11751,N_14784);
nand U15718 (N_15718,N_14486,N_14549);
xnor U15719 (N_15719,N_12851,N_10215);
nor U15720 (N_15720,N_11350,N_14413);
and U15721 (N_15721,N_14114,N_14247);
nor U15722 (N_15722,N_13312,N_10967);
xor U15723 (N_15723,N_14987,N_10125);
nand U15724 (N_15724,N_14644,N_11152);
nand U15725 (N_15725,N_11539,N_11495);
nand U15726 (N_15726,N_12793,N_13314);
and U15727 (N_15727,N_10923,N_11787);
xor U15728 (N_15728,N_10390,N_13104);
and U15729 (N_15729,N_14077,N_10117);
and U15730 (N_15730,N_10563,N_11870);
or U15731 (N_15731,N_14983,N_10437);
xor U15732 (N_15732,N_10719,N_11116);
nor U15733 (N_15733,N_13466,N_14564);
nor U15734 (N_15734,N_12894,N_13129);
and U15735 (N_15735,N_14055,N_10326);
and U15736 (N_15736,N_10803,N_12935);
and U15737 (N_15737,N_12521,N_13570);
nand U15738 (N_15738,N_13886,N_12356);
nand U15739 (N_15739,N_12236,N_11304);
nand U15740 (N_15740,N_14884,N_11225);
xor U15741 (N_15741,N_14052,N_12600);
and U15742 (N_15742,N_10464,N_10135);
nand U15743 (N_15743,N_14029,N_12987);
nor U15744 (N_15744,N_14874,N_13364);
xnor U15745 (N_15745,N_10666,N_12450);
and U15746 (N_15746,N_13553,N_12958);
nand U15747 (N_15747,N_11591,N_10758);
nor U15748 (N_15748,N_12046,N_11584);
and U15749 (N_15749,N_14599,N_11739);
or U15750 (N_15750,N_10652,N_13520);
and U15751 (N_15751,N_14968,N_12566);
nand U15752 (N_15752,N_10679,N_11298);
nand U15753 (N_15753,N_10509,N_11959);
nand U15754 (N_15754,N_14705,N_10576);
or U15755 (N_15755,N_13378,N_10879);
nor U15756 (N_15756,N_11785,N_13836);
and U15757 (N_15757,N_12040,N_12045);
xnor U15758 (N_15758,N_14936,N_14091);
nand U15759 (N_15759,N_13103,N_14468);
nand U15760 (N_15760,N_12101,N_14953);
or U15761 (N_15761,N_12789,N_11850);
xor U15762 (N_15762,N_11934,N_14912);
xnor U15763 (N_15763,N_12898,N_12061);
nand U15764 (N_15764,N_10083,N_10024);
or U15765 (N_15765,N_12796,N_13910);
or U15766 (N_15766,N_14407,N_13542);
nor U15767 (N_15767,N_14037,N_11341);
and U15768 (N_15768,N_12863,N_14978);
nor U15769 (N_15769,N_12892,N_11097);
nor U15770 (N_15770,N_13830,N_10119);
nor U15771 (N_15771,N_14825,N_11118);
and U15772 (N_15772,N_12821,N_11368);
and U15773 (N_15773,N_10006,N_11207);
or U15774 (N_15774,N_12555,N_11177);
nand U15775 (N_15775,N_12189,N_10522);
nand U15776 (N_15776,N_11485,N_14529);
and U15777 (N_15777,N_11819,N_14173);
xnor U15778 (N_15778,N_11918,N_11561);
xnor U15779 (N_15779,N_13004,N_13858);
nand U15780 (N_15780,N_13124,N_11769);
or U15781 (N_15781,N_13746,N_11570);
nand U15782 (N_15782,N_10881,N_11414);
or U15783 (N_15783,N_11174,N_14868);
nand U15784 (N_15784,N_12198,N_10837);
nor U15785 (N_15785,N_10866,N_13250);
nand U15786 (N_15786,N_10423,N_11264);
xor U15787 (N_15787,N_13454,N_11255);
nand U15788 (N_15788,N_10607,N_12753);
and U15789 (N_15789,N_14911,N_11661);
nor U15790 (N_15790,N_10685,N_10768);
and U15791 (N_15791,N_14446,N_12412);
xnor U15792 (N_15792,N_12161,N_13362);
or U15793 (N_15793,N_10306,N_12978);
nand U15794 (N_15794,N_10523,N_13833);
xor U15795 (N_15795,N_10318,N_10698);
nand U15796 (N_15796,N_11632,N_11353);
nand U15797 (N_15797,N_12809,N_11654);
or U15798 (N_15798,N_12178,N_12095);
nor U15799 (N_15799,N_14693,N_10777);
or U15800 (N_15800,N_14917,N_11811);
nand U15801 (N_15801,N_14151,N_14231);
xor U15802 (N_15802,N_11756,N_11010);
xnor U15803 (N_15803,N_11583,N_12966);
and U15804 (N_15804,N_11231,N_13244);
or U15805 (N_15805,N_11411,N_12560);
nor U15806 (N_15806,N_12392,N_10966);
xor U15807 (N_15807,N_13720,N_10750);
or U15808 (N_15808,N_11008,N_13411);
xor U15809 (N_15809,N_14078,N_13367);
or U15810 (N_15810,N_12881,N_14045);
nand U15811 (N_15811,N_13649,N_13329);
nand U15812 (N_15812,N_11672,N_14615);
nor U15813 (N_15813,N_10127,N_12995);
and U15814 (N_15814,N_14610,N_14300);
xnor U15815 (N_15815,N_11973,N_11634);
and U15816 (N_15816,N_14049,N_10581);
and U15817 (N_15817,N_10546,N_10200);
xnor U15818 (N_15818,N_12452,N_12601);
and U15819 (N_15819,N_11378,N_11101);
nor U15820 (N_15820,N_13994,N_13141);
and U15821 (N_15821,N_10605,N_11839);
nand U15822 (N_15822,N_14395,N_12318);
nand U15823 (N_15823,N_13802,N_12165);
or U15824 (N_15824,N_11865,N_10865);
or U15825 (N_15825,N_14239,N_11901);
xnor U15826 (N_15826,N_12337,N_12313);
or U15827 (N_15827,N_11014,N_13396);
xor U15828 (N_15828,N_13629,N_14704);
and U15829 (N_15829,N_13223,N_12603);
nor U15830 (N_15830,N_11173,N_13665);
or U15831 (N_15831,N_14989,N_14176);
and U15832 (N_15832,N_14396,N_13371);
xor U15833 (N_15833,N_10845,N_11957);
nand U15834 (N_15834,N_12325,N_13544);
nand U15835 (N_15835,N_13228,N_13604);
and U15836 (N_15836,N_13034,N_14427);
and U15837 (N_15837,N_14828,N_12653);
nor U15838 (N_15838,N_11325,N_10293);
nand U15839 (N_15839,N_13021,N_11452);
nand U15840 (N_15840,N_13740,N_12758);
xnor U15841 (N_15841,N_12050,N_10812);
or U15842 (N_15842,N_12563,N_14269);
nand U15843 (N_15843,N_10467,N_12692);
and U15844 (N_15844,N_10674,N_11394);
and U15845 (N_15845,N_11938,N_12769);
or U15846 (N_15846,N_11648,N_10075);
nand U15847 (N_15847,N_14972,N_13295);
nor U15848 (N_15848,N_14408,N_10297);
nand U15849 (N_15849,N_13736,N_11183);
nor U15850 (N_15850,N_13963,N_10479);
or U15851 (N_15851,N_12141,N_13756);
nand U15852 (N_15852,N_14308,N_14391);
and U15853 (N_15853,N_11524,N_12913);
nand U15854 (N_15854,N_13310,N_10143);
nand U15855 (N_15855,N_10797,N_13587);
or U15856 (N_15856,N_11562,N_11649);
and U15857 (N_15857,N_11422,N_12651);
xnor U15858 (N_15858,N_11980,N_13348);
nand U15859 (N_15859,N_13882,N_13108);
xor U15860 (N_15860,N_13760,N_14215);
nand U15861 (N_15861,N_12006,N_11670);
or U15862 (N_15862,N_11761,N_10505);
and U15863 (N_15863,N_14593,N_14752);
or U15864 (N_15864,N_14211,N_14639);
xor U15865 (N_15865,N_12685,N_10590);
or U15866 (N_15866,N_11257,N_12181);
nor U15867 (N_15867,N_11610,N_11178);
and U15868 (N_15868,N_13477,N_12535);
or U15869 (N_15869,N_13316,N_13001);
or U15870 (N_15870,N_11884,N_13972);
xor U15871 (N_15871,N_10104,N_10395);
xor U15872 (N_15872,N_10394,N_11241);
and U15873 (N_15873,N_11624,N_14995);
or U15874 (N_15874,N_13894,N_11856);
nor U15875 (N_15875,N_14404,N_12641);
xnor U15876 (N_15876,N_11129,N_14008);
nor U15877 (N_15877,N_14707,N_12682);
or U15878 (N_15878,N_13808,N_14195);
xnor U15879 (N_15879,N_12138,N_14240);
nor U15880 (N_15880,N_14470,N_10961);
and U15881 (N_15881,N_13187,N_12437);
nand U15882 (N_15882,N_11480,N_14434);
and U15883 (N_15883,N_10304,N_13648);
nor U15884 (N_15884,N_13765,N_13011);
and U15885 (N_15885,N_13998,N_11389);
or U15886 (N_15886,N_14130,N_14378);
nand U15887 (N_15887,N_13540,N_11995);
xnor U15888 (N_15888,N_14260,N_12976);
xor U15889 (N_15889,N_14706,N_11431);
or U15890 (N_15890,N_11338,N_13191);
xnor U15891 (N_15891,N_11028,N_14600);
and U15892 (N_15892,N_14540,N_10483);
nand U15893 (N_15893,N_11439,N_12807);
nor U15894 (N_15894,N_11498,N_10868);
or U15895 (N_15895,N_12140,N_12738);
or U15896 (N_15896,N_14357,N_11889);
xor U15897 (N_15897,N_12216,N_10638);
xnor U15898 (N_15898,N_13029,N_12970);
and U15899 (N_15899,N_11734,N_10992);
nor U15900 (N_15900,N_11712,N_10572);
nor U15901 (N_15901,N_12891,N_14914);
nor U15902 (N_15902,N_13727,N_13966);
or U15903 (N_15903,N_13133,N_12902);
xor U15904 (N_15904,N_13877,N_11375);
nand U15905 (N_15905,N_14420,N_13903);
or U15906 (N_15906,N_11604,N_10612);
nand U15907 (N_15907,N_13530,N_11729);
and U15908 (N_15908,N_11252,N_12556);
nand U15909 (N_15909,N_11538,N_10229);
and U15910 (N_15910,N_14634,N_12064);
nand U15911 (N_15911,N_14518,N_13227);
nand U15912 (N_15912,N_12658,N_13632);
nand U15913 (N_15913,N_11453,N_11469);
nand U15914 (N_15914,N_11804,N_13974);
xor U15915 (N_15915,N_12757,N_14865);
nand U15916 (N_15916,N_14880,N_12023);
or U15917 (N_15917,N_12879,N_11963);
or U15918 (N_15918,N_13127,N_13638);
nor U15919 (N_15919,N_13932,N_14525);
nand U15920 (N_15920,N_13146,N_12875);
or U15921 (N_15921,N_10334,N_11532);
xnor U15922 (N_15922,N_12293,N_14853);
or U15923 (N_15923,N_10573,N_14072);
nand U15924 (N_15924,N_10405,N_14387);
xor U15925 (N_15925,N_10957,N_14129);
or U15926 (N_15926,N_12815,N_14057);
or U15927 (N_15927,N_10226,N_13009);
xnor U15928 (N_15928,N_14555,N_13761);
xor U15929 (N_15929,N_13256,N_10434);
nand U15930 (N_15930,N_14244,N_10268);
xnor U15931 (N_15931,N_12308,N_14935);
nand U15932 (N_15932,N_13770,N_13956);
xor U15933 (N_15933,N_12777,N_13303);
xor U15934 (N_15934,N_12096,N_14998);
nand U15935 (N_15935,N_13165,N_11336);
or U15936 (N_15936,N_14816,N_10551);
nand U15937 (N_15937,N_10544,N_13692);
nor U15938 (N_15938,N_10415,N_14283);
or U15939 (N_15939,N_14474,N_14531);
and U15940 (N_15940,N_14444,N_14185);
nor U15941 (N_15941,N_14801,N_10849);
xnor U15942 (N_15942,N_11111,N_10520);
nor U15943 (N_15943,N_10927,N_13816);
nor U15944 (N_15944,N_12333,N_11723);
nand U15945 (N_15945,N_10896,N_12583);
nand U15946 (N_15946,N_14821,N_13492);
and U15947 (N_15947,N_10941,N_13484);
or U15948 (N_15948,N_10156,N_13610);
xor U15949 (N_15949,N_13175,N_10494);
nand U15950 (N_15950,N_11373,N_10690);
or U15951 (N_15951,N_14259,N_10855);
nor U15952 (N_15952,N_14565,N_13677);
nand U15953 (N_15953,N_10722,N_12380);
and U15954 (N_15954,N_10029,N_13056);
or U15955 (N_15955,N_14538,N_12868);
and U15956 (N_15956,N_14974,N_12273);
or U15957 (N_15957,N_12955,N_14753);
nand U15958 (N_15958,N_11646,N_12433);
or U15959 (N_15959,N_11685,N_13390);
and U15960 (N_15960,N_12712,N_14826);
xnor U15961 (N_15961,N_10173,N_10921);
nor U15962 (N_15962,N_14042,N_13257);
xor U15963 (N_15963,N_14136,N_11307);
and U15964 (N_15964,N_11879,N_12052);
nand U15965 (N_15965,N_11468,N_10507);
nand U15966 (N_15966,N_13405,N_12571);
nand U15967 (N_15967,N_13927,N_11349);
nand U15968 (N_15968,N_12080,N_13482);
and U15969 (N_15969,N_14152,N_10909);
nand U15970 (N_15970,N_10497,N_10360);
nor U15971 (N_15971,N_12162,N_10963);
and U15972 (N_15972,N_10374,N_12594);
or U15973 (N_15973,N_14646,N_12512);
xnor U15974 (N_15974,N_13006,N_13357);
nor U15975 (N_15975,N_12686,N_11821);
xnor U15976 (N_15976,N_12695,N_12173);
nand U15977 (N_15977,N_12020,N_13225);
or U15978 (N_15978,N_11534,N_10069);
nor U15979 (N_15979,N_12154,N_11210);
nand U15980 (N_15980,N_10116,N_12850);
and U15981 (N_15981,N_11337,N_14581);
xor U15982 (N_15982,N_12451,N_10131);
nand U15983 (N_15983,N_11718,N_12888);
nor U15984 (N_15984,N_12548,N_13121);
or U15985 (N_15985,N_13271,N_10907);
and U15986 (N_15986,N_11759,N_12177);
xor U15987 (N_15987,N_14519,N_11528);
nand U15988 (N_15988,N_14534,N_10902);
and U15989 (N_15989,N_14517,N_14004);
and U15990 (N_15990,N_10628,N_14330);
nand U15991 (N_15991,N_12950,N_14346);
nor U15992 (N_15992,N_11869,N_11122);
nor U15993 (N_15993,N_14554,N_10106);
or U15994 (N_15994,N_11021,N_10072);
nand U15995 (N_15995,N_14950,N_10313);
nand U15996 (N_15996,N_13914,N_10580);
nor U15997 (N_15997,N_11436,N_12586);
and U15998 (N_15998,N_12031,N_11605);
and U15999 (N_15999,N_11110,N_13441);
nand U16000 (N_16000,N_14284,N_10241);
and U16001 (N_16001,N_12252,N_14086);
or U16002 (N_16002,N_12951,N_12665);
or U16003 (N_16003,N_13241,N_14766);
nor U16004 (N_16004,N_13786,N_13890);
nor U16005 (N_16005,N_14163,N_13093);
and U16006 (N_16006,N_13719,N_13423);
or U16007 (N_16007,N_10864,N_11288);
xnor U16008 (N_16008,N_12790,N_13152);
and U16009 (N_16009,N_11822,N_12314);
nor U16010 (N_16010,N_13839,N_12136);
and U16011 (N_16011,N_10380,N_12391);
and U16012 (N_16012,N_13826,N_14622);
or U16013 (N_16013,N_13868,N_12367);
and U16014 (N_16014,N_13399,N_13904);
xor U16015 (N_16015,N_14297,N_12761);
and U16016 (N_16016,N_12156,N_10670);
xnor U16017 (N_16017,N_14168,N_11025);
nand U16018 (N_16018,N_10962,N_12015);
nor U16019 (N_16019,N_13472,N_11022);
or U16020 (N_16020,N_14806,N_11784);
nand U16021 (N_16021,N_11051,N_10195);
and U16022 (N_16022,N_10669,N_11607);
nand U16023 (N_16023,N_13160,N_13819);
or U16024 (N_16024,N_10138,N_12331);
and U16025 (N_16025,N_12805,N_14450);
nand U16026 (N_16026,N_12783,N_11574);
xor U16027 (N_16027,N_10211,N_12183);
nand U16028 (N_16028,N_10964,N_14804);
or U16029 (N_16029,N_11511,N_14896);
nor U16030 (N_16030,N_13153,N_11601);
nand U16031 (N_16031,N_14460,N_11233);
or U16032 (N_16032,N_13020,N_13627);
nor U16033 (N_16033,N_14643,N_13729);
or U16034 (N_16034,N_11044,N_10678);
nor U16035 (N_16035,N_10164,N_12012);
nand U16036 (N_16036,N_10492,N_10683);
or U16037 (N_16037,N_13086,N_13712);
xor U16038 (N_16038,N_10684,N_14623);
or U16039 (N_16039,N_13965,N_10166);
and U16040 (N_16040,N_10826,N_14141);
nand U16041 (N_16041,N_12448,N_12076);
xor U16042 (N_16042,N_14723,N_12985);
nor U16043 (N_16043,N_11514,N_11501);
xor U16044 (N_16044,N_10643,N_13249);
nor U16045 (N_16045,N_14472,N_10256);
nand U16046 (N_16046,N_10271,N_10460);
nand U16047 (N_16047,N_12069,N_13694);
xnor U16048 (N_16048,N_10602,N_12814);
and U16049 (N_16049,N_10291,N_11372);
xor U16050 (N_16050,N_14062,N_14126);
xnor U16051 (N_16051,N_10124,N_14190);
xnor U16052 (N_16052,N_12035,N_12617);
xor U16053 (N_16053,N_11209,N_14757);
xnor U16054 (N_16054,N_12360,N_12303);
nand U16055 (N_16055,N_10955,N_12129);
xor U16056 (N_16056,N_13290,N_10455);
nor U16057 (N_16057,N_14056,N_10160);
xor U16058 (N_16058,N_14591,N_14222);
and U16059 (N_16059,N_14588,N_13439);
or U16060 (N_16060,N_13777,N_11287);
xnor U16061 (N_16061,N_12688,N_13062);
nor U16062 (N_16062,N_14099,N_11221);
xnor U16063 (N_16063,N_10823,N_14482);
or U16064 (N_16064,N_11551,N_13871);
nand U16065 (N_16065,N_13911,N_10682);
or U16066 (N_16066,N_11727,N_10027);
xor U16067 (N_16067,N_14786,N_11319);
and U16068 (N_16068,N_12730,N_11590);
or U16069 (N_16069,N_13013,N_10518);
nand U16070 (N_16070,N_12933,N_11027);
nand U16071 (N_16071,N_13495,N_10852);
xor U16072 (N_16072,N_12873,N_11747);
and U16073 (N_16073,N_11181,N_10093);
nor U16074 (N_16074,N_10755,N_11330);
and U16075 (N_16075,N_10858,N_13050);
xor U16076 (N_16076,N_10090,N_10454);
nor U16077 (N_16077,N_12752,N_10485);
and U16078 (N_16078,N_12631,N_13107);
and U16079 (N_16079,N_12379,N_13342);
and U16080 (N_16080,N_13354,N_10706);
or U16081 (N_16081,N_14720,N_10856);
nand U16082 (N_16082,N_12152,N_14573);
and U16083 (N_16083,N_14504,N_13318);
nand U16084 (N_16084,N_11838,N_11318);
nor U16085 (N_16085,N_11613,N_14709);
nand U16086 (N_16086,N_11618,N_11006);
and U16087 (N_16087,N_12864,N_13280);
or U16088 (N_16088,N_12733,N_13064);
xor U16089 (N_16089,N_14835,N_10228);
xnor U16090 (N_16090,N_10245,N_13238);
xnor U16091 (N_16091,N_12889,N_11653);
or U16092 (N_16092,N_10888,N_13022);
nand U16093 (N_16093,N_13375,N_12147);
nor U16094 (N_16094,N_13502,N_13327);
nor U16095 (N_16095,N_13676,N_12347);
or U16096 (N_16096,N_12735,N_12256);
xnor U16097 (N_16097,N_14466,N_12302);
xnor U16098 (N_16098,N_14713,N_12049);
nor U16099 (N_16099,N_12874,N_10320);
xor U16100 (N_16100,N_12953,N_11159);
or U16101 (N_16101,N_11138,N_10419);
nor U16102 (N_16102,N_10784,N_14954);
nand U16103 (N_16103,N_12345,N_12417);
and U16104 (N_16104,N_13801,N_13916);
or U16105 (N_16105,N_11652,N_12746);
or U16106 (N_16106,N_11824,N_14586);
nor U16107 (N_16107,N_13246,N_14298);
and U16108 (N_16108,N_12469,N_14627);
nand U16109 (N_16109,N_13549,N_11285);
nor U16110 (N_16110,N_11873,N_12171);
xor U16111 (N_16111,N_10233,N_12316);
nand U16112 (N_16112,N_10820,N_12053);
and U16113 (N_16113,N_10191,N_12430);
and U16114 (N_16114,N_14793,N_11266);
nand U16115 (N_16115,N_13748,N_11366);
and U16116 (N_16116,N_13098,N_14477);
or U16117 (N_16117,N_10257,N_10335);
and U16118 (N_16118,N_12039,N_13591);
or U16119 (N_16119,N_11689,N_10058);
and U16120 (N_16120,N_13870,N_10183);
xnor U16121 (N_16121,N_14425,N_13320);
nor U16122 (N_16122,N_10542,N_13759);
xor U16123 (N_16123,N_10554,N_10244);
nor U16124 (N_16124,N_11888,N_12811);
and U16125 (N_16125,N_10281,N_10433);
or U16126 (N_16126,N_14317,N_10993);
or U16127 (N_16127,N_10070,N_12353);
and U16128 (N_16128,N_12327,N_10593);
and U16129 (N_16129,N_11695,N_10398);
or U16130 (N_16130,N_10878,N_11996);
or U16131 (N_16131,N_10736,N_11599);
and U16132 (N_16132,N_12257,N_13007);
or U16133 (N_16133,N_13035,N_13475);
nand U16134 (N_16134,N_14780,N_10407);
nand U16135 (N_16135,N_14336,N_14734);
or U16136 (N_16136,N_10008,N_13811);
xnor U16137 (N_16137,N_11237,N_12550);
and U16138 (N_16138,N_11092,N_14877);
nor U16139 (N_16139,N_11752,N_10251);
nor U16140 (N_16140,N_13895,N_14219);
or U16141 (N_16141,N_11641,N_11270);
nand U16142 (N_16142,N_10915,N_12103);
and U16143 (N_16143,N_11863,N_11308);
nand U16144 (N_16144,N_14089,N_13242);
xor U16145 (N_16145,N_12589,N_13155);
or U16146 (N_16146,N_10998,N_11834);
or U16147 (N_16147,N_14242,N_14265);
nand U16148 (N_16148,N_11924,N_13687);
xor U16149 (N_16149,N_13409,N_12335);
or U16150 (N_16150,N_10861,N_12557);
or U16151 (N_16151,N_14137,N_14133);
nand U16152 (N_16152,N_13417,N_14686);
nand U16153 (N_16153,N_11999,N_12607);
nand U16154 (N_16154,N_11683,N_10002);
and U16155 (N_16155,N_12833,N_11482);
or U16156 (N_16156,N_12689,N_11626);
nor U16157 (N_16157,N_14447,N_12344);
or U16158 (N_16158,N_12523,N_10120);
nor U16159 (N_16159,N_14002,N_13234);
and U16160 (N_16160,N_11015,N_14787);
xor U16161 (N_16161,N_10588,N_14492);
or U16162 (N_16162,N_10466,N_11681);
or U16163 (N_16163,N_10321,N_11954);
xnor U16164 (N_16164,N_14798,N_12120);
nor U16165 (N_16165,N_10165,N_14653);
or U16166 (N_16166,N_14558,N_11525);
or U16167 (N_16167,N_12310,N_14678);
or U16168 (N_16168,N_13935,N_12155);
and U16169 (N_16169,N_11007,N_12168);
nor U16170 (N_16170,N_11535,N_14142);
and U16171 (N_16171,N_14429,N_12869);
nor U16172 (N_16172,N_14410,N_13487);
nand U16173 (N_16173,N_11917,N_11942);
and U16174 (N_16174,N_13598,N_12285);
or U16175 (N_16175,N_13751,N_10949);
and U16176 (N_16176,N_10778,N_12397);
nand U16177 (N_16177,N_10025,N_12895);
or U16178 (N_16178,N_12663,N_10089);
nor U16179 (N_16179,N_12133,N_12439);
nand U16180 (N_16180,N_14380,N_12760);
or U16181 (N_16181,N_12997,N_10095);
or U16182 (N_16182,N_10456,N_11933);
nor U16183 (N_16183,N_11847,N_14041);
nand U16184 (N_16184,N_10213,N_11549);
or U16185 (N_16185,N_14324,N_10629);
xnor U16186 (N_16186,N_14095,N_12326);
nand U16187 (N_16187,N_12800,N_13783);
nor U16188 (N_16188,N_11808,N_13452);
or U16189 (N_16189,N_10278,N_11402);
or U16190 (N_16190,N_11292,N_12022);
nor U16191 (N_16191,N_11697,N_14023);
or U16192 (N_16192,N_11065,N_12613);
or U16193 (N_16193,N_13909,N_14294);
nor U16194 (N_16194,N_11230,N_10782);
nand U16195 (N_16195,N_14220,N_14708);
nor U16196 (N_16196,N_11688,N_11657);
or U16197 (N_16197,N_13528,N_12434);
nand U16198 (N_16198,N_11424,N_13812);
xnor U16199 (N_16199,N_13888,N_13730);
and U16200 (N_16200,N_14348,N_14749);
or U16201 (N_16201,N_11877,N_13429);
and U16202 (N_16202,N_12106,N_14696);
and U16203 (N_16203,N_13755,N_14451);
and U16204 (N_16204,N_13917,N_10440);
nor U16205 (N_16205,N_14115,N_13784);
or U16206 (N_16206,N_12546,N_11500);
nor U16207 (N_16207,N_10208,N_13744);
and U16208 (N_16208,N_13551,N_12661);
nand U16209 (N_16209,N_12597,N_11908);
xor U16210 (N_16210,N_10040,N_10827);
nor U16211 (N_16211,N_14490,N_14164);
nand U16212 (N_16212,N_14392,N_11259);
or U16213 (N_16213,N_14722,N_11896);
nor U16214 (N_16214,N_12960,N_12859);
nor U16215 (N_16215,N_12870,N_14288);
nand U16216 (N_16216,N_13757,N_12785);
xnor U16217 (N_16217,N_10074,N_11442);
nand U16218 (N_16218,N_10239,N_12957);
nor U16219 (N_16219,N_11242,N_11272);
nor U16220 (N_16220,N_13515,N_14882);
or U16221 (N_16221,N_13655,N_14850);
xnor U16222 (N_16222,N_14813,N_14457);
and U16223 (N_16223,N_13332,N_12726);
and U16224 (N_16224,N_14672,N_11573);
nor U16225 (N_16225,N_12226,N_14355);
and U16226 (N_16226,N_13924,N_13159);
xor U16227 (N_16227,N_13401,N_10137);
or U16228 (N_16228,N_14456,N_11247);
and U16229 (N_16229,N_14022,N_11356);
nor U16230 (N_16230,N_11443,N_13283);
or U16231 (N_16231,N_11429,N_12952);
xor U16232 (N_16232,N_14006,N_12030);
and U16233 (N_16233,N_10387,N_10033);
xnor U16234 (N_16234,N_12463,N_11403);
nor U16235 (N_16235,N_11810,N_10449);
nor U16236 (N_16236,N_12206,N_10733);
nand U16237 (N_16237,N_11161,N_10726);
xor U16238 (N_16238,N_13135,N_13725);
and U16239 (N_16239,N_12032,N_12319);
or U16240 (N_16240,N_10231,N_12944);
or U16241 (N_16241,N_13016,N_13434);
nor U16242 (N_16242,N_13991,N_11631);
xnor U16243 (N_16243,N_12799,N_14582);
or U16244 (N_16244,N_14894,N_13527);
xor U16245 (N_16245,N_11489,N_12562);
xor U16246 (N_16246,N_12113,N_12964);
or U16247 (N_16247,N_13095,N_12939);
and U16248 (N_16248,N_10417,N_12998);
nor U16249 (N_16249,N_12395,N_13893);
or U16250 (N_16250,N_14363,N_12358);
or U16251 (N_16251,N_10632,N_13370);
nand U16252 (N_16252,N_14485,N_14230);
nor U16253 (N_16253,N_11608,N_10301);
nand U16254 (N_16254,N_11096,N_11108);
nand U16255 (N_16255,N_11617,N_13218);
nor U16256 (N_16256,N_10373,N_10877);
xnor U16257 (N_16257,N_13931,N_13659);
or U16258 (N_16258,N_10991,N_11515);
nand U16259 (N_16259,N_14385,N_13393);
xnor U16260 (N_16260,N_13014,N_11932);
or U16261 (N_16261,N_10981,N_14040);
nor U16262 (N_16262,N_11250,N_11968);
nor U16263 (N_16263,N_10842,N_11045);
or U16264 (N_16264,N_11945,N_10883);
nand U16265 (N_16265,N_14375,N_10015);
nor U16266 (N_16266,N_13092,N_14981);
nor U16267 (N_16267,N_13780,N_11380);
nor U16268 (N_16268,N_11910,N_13537);
xor U16269 (N_16269,N_13560,N_13726);
and U16270 (N_16270,N_11704,N_11907);
and U16271 (N_16271,N_12501,N_10816);
or U16272 (N_16272,N_13929,N_14098);
and U16273 (N_16273,N_14397,N_14266);
and U16274 (N_16274,N_14268,N_11091);
and U16275 (N_16275,N_13120,N_10480);
xor U16276 (N_16276,N_13069,N_14347);
nand U16277 (N_16277,N_14496,N_13224);
or U16278 (N_16278,N_11983,N_14909);
xor U16279 (N_16279,N_11009,N_13443);
and U16280 (N_16280,N_14094,N_12495);
nor U16281 (N_16281,N_10378,N_12077);
or U16282 (N_16282,N_13070,N_12405);
xnor U16283 (N_16283,N_12245,N_10547);
nor U16284 (N_16284,N_14059,N_10371);
nand U16285 (N_16285,N_13717,N_13671);
and U16286 (N_16286,N_10003,N_12222);
xor U16287 (N_16287,N_11529,N_10818);
or U16288 (N_16288,N_10693,N_13374);
xor U16289 (N_16289,N_10985,N_12654);
nand U16290 (N_16290,N_13800,N_13365);
and U16291 (N_16291,N_11053,N_10566);
nor U16292 (N_16292,N_10193,N_10276);
nor U16293 (N_16293,N_10051,N_12163);
nor U16294 (N_16294,N_11208,N_14807);
xnor U16295 (N_16295,N_10591,N_13724);
or U16296 (N_16296,N_10207,N_13516);
nor U16297 (N_16297,N_14858,N_11722);
xnor U16298 (N_16298,N_12839,N_11635);
or U16299 (N_16299,N_13990,N_10500);
xor U16300 (N_16300,N_14402,N_11034);
and U16301 (N_16301,N_12378,N_14893);
nand U16302 (N_16302,N_10470,N_11944);
xor U16303 (N_16303,N_14663,N_10779);
and U16304 (N_16304,N_12574,N_10296);
xor U16305 (N_16305,N_13296,N_11364);
or U16306 (N_16306,N_12801,N_14631);
xnor U16307 (N_16307,N_11911,N_14000);
xnor U16308 (N_16308,N_14019,N_11682);
xnor U16309 (N_16309,N_13512,N_13158);
nor U16310 (N_16310,N_11893,N_12176);
nand U16311 (N_16311,N_10212,N_11467);
nor U16312 (N_16312,N_13650,N_12669);
and U16313 (N_16313,N_11700,N_12505);
or U16314 (N_16314,N_14740,N_13080);
nor U16315 (N_16315,N_10644,N_11788);
xnor U16316 (N_16316,N_14494,N_14351);
nand U16317 (N_16317,N_12727,N_13785);
and U16318 (N_16318,N_12211,N_12389);
xnor U16319 (N_16319,N_13618,N_13199);
nand U16320 (N_16320,N_10375,N_11076);
xnor U16321 (N_16321,N_12287,N_10203);
or U16322 (N_16322,N_13372,N_12186);
nand U16323 (N_16323,N_11781,N_10336);
nand U16324 (N_16324,N_11148,N_10799);
and U16325 (N_16325,N_14776,N_14003);
nor U16326 (N_16326,N_11352,N_13675);
nor U16327 (N_16327,N_12112,N_12458);
and U16328 (N_16328,N_12595,N_12445);
xor U16329 (N_16329,N_12253,N_12260);
or U16330 (N_16330,N_10432,N_11369);
and U16331 (N_16331,N_10452,N_12487);
nor U16332 (N_16332,N_14716,N_10399);
nor U16333 (N_16333,N_13198,N_11474);
nand U16334 (N_16334,N_10465,N_14399);
or U16335 (N_16335,N_10139,N_10931);
xor U16336 (N_16336,N_13430,N_10920);
or U16337 (N_16337,N_14823,N_13182);
and U16338 (N_16338,N_11106,N_11754);
nor U16339 (N_16339,N_14172,N_12473);
xor U16340 (N_16340,N_13823,N_11223);
nand U16341 (N_16341,N_12897,N_12079);
nor U16342 (N_16342,N_12065,N_10640);
or U16343 (N_16343,N_11512,N_11731);
xor U16344 (N_16344,N_14578,N_11112);
nand U16345 (N_16345,N_13905,N_11506);
nor U16346 (N_16346,N_11057,N_10801);
nor U16347 (N_16347,N_10771,N_13324);
xor U16348 (N_16348,N_12919,N_11708);
nand U16349 (N_16349,N_11935,N_13645);
nand U16350 (N_16350,N_10324,N_11567);
nor U16351 (N_16351,N_13406,N_10676);
xnor U16352 (N_16352,N_11832,N_14949);
nand U16353 (N_16353,N_11900,N_10954);
or U16354 (N_16354,N_10898,N_14368);
or U16355 (N_16355,N_11728,N_13368);
and U16356 (N_16356,N_13517,N_13852);
and U16357 (N_16357,N_14563,N_10108);
nand U16358 (N_16358,N_10260,N_14948);
xor U16359 (N_16359,N_12797,N_12779);
or U16360 (N_16360,N_11585,N_10959);
xor U16361 (N_16361,N_13605,N_13031);
nand U16362 (N_16362,N_10005,N_10789);
nor U16363 (N_16363,N_10811,N_14170);
nor U16364 (N_16364,N_12788,N_12299);
xnor U16365 (N_16365,N_12215,N_14715);
nand U16366 (N_16366,N_13041,N_14503);
or U16367 (N_16367,N_12818,N_13518);
or U16368 (N_16368,N_12058,N_11690);
nor U16369 (N_16369,N_13363,N_12016);
or U16370 (N_16370,N_10060,N_13207);
or U16371 (N_16371,N_14795,N_11067);
xor U16372 (N_16372,N_14360,N_13701);
or U16373 (N_16373,N_13245,N_14092);
nor U16374 (N_16374,N_14748,N_13023);
xor U16375 (N_16375,N_12506,N_10721);
or U16376 (N_16376,N_14979,N_13358);
xor U16377 (N_16377,N_13589,N_13101);
and U16378 (N_16378,N_14109,N_10052);
xnor U16379 (N_16379,N_12288,N_10579);
xor U16380 (N_16380,N_13984,N_13849);
nand U16381 (N_16381,N_12475,N_12698);
xor U16382 (N_16382,N_13414,N_13500);
and U16383 (N_16383,N_13232,N_11663);
or U16384 (N_16384,N_14840,N_13208);
or U16385 (N_16385,N_11357,N_13696);
xnor U16386 (N_16386,N_10333,N_10240);
nor U16387 (N_16387,N_12362,N_10948);
nor U16388 (N_16388,N_13181,N_10549);
and U16389 (N_16389,N_10930,N_14463);
nand U16390 (N_16390,N_11548,N_11416);
nand U16391 (N_16391,N_11816,N_12021);
or U16392 (N_16392,N_12164,N_11926);
xnor U16393 (N_16393,N_11033,N_11638);
and U16394 (N_16394,N_11966,N_13840);
or U16395 (N_16395,N_11651,N_10020);
nor U16396 (N_16396,N_11851,N_10940);
xor U16397 (N_16397,N_14830,N_13311);
nand U16398 (N_16398,N_13444,N_10704);
nor U16399 (N_16399,N_12286,N_11636);
or U16400 (N_16400,N_11245,N_12640);
nand U16401 (N_16401,N_12993,N_12237);
nand U16402 (N_16402,N_11943,N_11321);
xor U16403 (N_16403,N_12068,N_10196);
or U16404 (N_16404,N_13163,N_14924);
and U16405 (N_16405,N_13827,N_14650);
xor U16406 (N_16406,N_10042,N_14509);
nand U16407 (N_16407,N_11958,N_10952);
and U16408 (N_16408,N_10700,N_12401);
nand U16409 (N_16409,N_12201,N_14475);
xor U16410 (N_16410,N_12728,N_10687);
nand U16411 (N_16411,N_11263,N_11807);
and U16412 (N_16412,N_13576,N_10011);
or U16413 (N_16413,N_11662,N_14026);
xnor U16414 (N_16414,N_13483,N_11185);
nand U16415 (N_16415,N_12545,N_11279);
xnor U16416 (N_16416,N_11260,N_12218);
and U16417 (N_16417,N_12081,N_10255);
and U16418 (N_16418,N_12018,N_13602);
xnor U16419 (N_16419,N_13385,N_10102);
nor U16420 (N_16420,N_13541,N_14341);
nor U16421 (N_16421,N_12224,N_10548);
nor U16422 (N_16422,N_11772,N_12736);
nor U16423 (N_16423,N_13750,N_11434);
xor U16424 (N_16424,N_13268,N_11381);
or U16425 (N_16425,N_10235,N_14236);
nand U16426 (N_16426,N_13448,N_14657);
nand U16427 (N_16427,N_12108,N_10491);
nor U16428 (N_16428,N_12071,N_11843);
and U16429 (N_16429,N_11360,N_12486);
or U16430 (N_16430,N_13178,N_13313);
or U16431 (N_16431,N_11664,N_11188);
nand U16432 (N_16432,N_12605,N_13970);
nand U16433 (N_16433,N_13294,N_12748);
nand U16434 (N_16434,N_13951,N_10662);
and U16435 (N_16435,N_14202,N_12000);
or U16436 (N_16436,N_13630,N_11758);
and U16437 (N_16437,N_11575,N_11930);
xnor U16438 (N_16438,N_10737,N_14087);
xor U16439 (N_16439,N_13722,N_12497);
nor U16440 (N_16440,N_11069,N_10201);
and U16441 (N_16441,N_11432,N_13162);
and U16442 (N_16442,N_11753,N_13197);
xor U16443 (N_16443,N_14763,N_14350);
nand U16444 (N_16444,N_14038,N_12532);
and U16445 (N_16445,N_12373,N_11301);
nand U16446 (N_16446,N_13934,N_11774);
nor U16447 (N_16447,N_13651,N_14824);
and U16448 (N_16448,N_10978,N_11860);
xor U16449 (N_16449,N_14191,N_11293);
nor U16450 (N_16450,N_10288,N_10934);
xnor U16451 (N_16451,N_13835,N_12041);
or U16452 (N_16452,N_14984,N_14505);
nor U16453 (N_16453,N_10798,N_11577);
nor U16454 (N_16454,N_13856,N_13733);
and U16455 (N_16455,N_14831,N_10623);
nor U16456 (N_16456,N_14443,N_10181);
nor U16457 (N_16457,N_10026,N_11328);
nor U16458 (N_16458,N_12294,N_13221);
or U16459 (N_16459,N_10521,N_11741);
nand U16460 (N_16460,N_12836,N_10840);
xor U16461 (N_16461,N_13555,N_13942);
or U16462 (N_16462,N_13333,N_13539);
nand U16463 (N_16463,N_13884,N_10364);
xnor U16464 (N_16464,N_14508,N_10202);
nand U16465 (N_16465,N_12459,N_13531);
and U16466 (N_16466,N_11768,N_12038);
nand U16467 (N_16467,N_11398,N_11410);
nand U16468 (N_16468,N_12604,N_13106);
and U16469 (N_16469,N_13255,N_12078);
nor U16470 (N_16470,N_11284,N_13000);
and U16471 (N_16471,N_12169,N_13173);
nand U16472 (N_16472,N_12090,N_10123);
and U16473 (N_16473,N_10356,N_13273);
and U16474 (N_16474,N_11941,N_12871);
or U16475 (N_16475,N_12415,N_10383);
xnor U16476 (N_16476,N_10209,N_10739);
xnor U16477 (N_16477,N_10368,N_14411);
xor U16478 (N_16478,N_12470,N_11993);
and U16479 (N_16479,N_10900,N_13142);
and U16480 (N_16480,N_14188,N_11465);
or U16481 (N_16481,N_11105,N_12212);
nor U16482 (N_16482,N_12488,N_14118);
xor U16483 (N_16483,N_12072,N_10012);
or U16484 (N_16484,N_13983,N_12723);
and U16485 (N_16485,N_12004,N_11099);
xnor U16486 (N_16486,N_10552,N_12028);
xor U16487 (N_16487,N_13975,N_10041);
nor U16488 (N_16488,N_14743,N_11031);
xnor U16489 (N_16489,N_11377,N_13102);
and U16490 (N_16490,N_14562,N_10199);
nor U16491 (N_16491,N_11371,N_13510);
and U16492 (N_16492,N_11149,N_10872);
or U16493 (N_16493,N_12175,N_11359);
or U16494 (N_16494,N_14076,N_14837);
xnor U16495 (N_16495,N_10701,N_13930);
or U16496 (N_16496,N_12411,N_14366);
or U16497 (N_16497,N_10168,N_12291);
nand U16498 (N_16498,N_12547,N_12425);
xor U16499 (N_16499,N_11615,N_10667);
or U16500 (N_16500,N_10717,N_14603);
nor U16501 (N_16501,N_12217,N_12812);
nand U16502 (N_16502,N_13383,N_13229);
nor U16503 (N_16503,N_11224,N_10595);
nor U16504 (N_16504,N_14147,N_10067);
xor U16505 (N_16505,N_14014,N_14349);
nor U16506 (N_16506,N_14913,N_11639);
xnor U16507 (N_16507,N_10787,N_14647);
nor U16508 (N_16508,N_11435,N_12639);
or U16509 (N_16509,N_12922,N_14946);
nor U16510 (N_16510,N_10039,N_13798);
and U16511 (N_16511,N_14845,N_11314);
nor U16512 (N_16512,N_12569,N_12696);
nor U16513 (N_16513,N_14970,N_12756);
or U16514 (N_16514,N_11331,N_14303);
nor U16515 (N_16515,N_10425,N_10611);
nand U16516 (N_16516,N_13813,N_14177);
xor U16517 (N_16517,N_14932,N_12982);
or U16518 (N_16518,N_12579,N_12258);
nand U16519 (N_16519,N_11448,N_14815);
nand U16520 (N_16520,N_14082,N_10702);
and U16521 (N_16521,N_13210,N_10178);
xnor U16522 (N_16522,N_10259,N_13626);
or U16523 (N_16523,N_11871,N_10047);
nand U16524 (N_16524,N_11998,N_10345);
xnor U16525 (N_16525,N_11612,N_13478);
or U16526 (N_16526,N_12914,N_13493);
or U16527 (N_16527,N_11158,N_12248);
and U16528 (N_16528,N_14483,N_12502);
or U16529 (N_16529,N_14596,N_10817);
nand U16530 (N_16530,N_10068,N_13545);
nand U16531 (N_16531,N_12621,N_10136);
nor U16532 (N_16532,N_14453,N_11186);
xnor U16533 (N_16533,N_11295,N_13611);
nor U16534 (N_16534,N_10342,N_11477);
nor U16535 (N_16535,N_11836,N_12111);
or U16536 (N_16536,N_12249,N_13307);
nand U16537 (N_16537,N_11703,N_11564);
nor U16538 (N_16538,N_11374,N_11457);
nand U16539 (N_16539,N_10833,N_13274);
nor U16540 (N_16540,N_13795,N_14856);
nor U16541 (N_16541,N_11005,N_12507);
xnor U16542 (N_16542,N_14849,N_10748);
xnor U16543 (N_16543,N_14455,N_12194);
xnor U16544 (N_16544,N_13912,N_13033);
and U16545 (N_16545,N_14181,N_13386);
and U16546 (N_16546,N_11552,N_13656);
nand U16547 (N_16547,N_14607,N_10770);
xnor U16548 (N_16548,N_11437,N_13615);
or U16549 (N_16549,N_10869,N_12918);
nor U16550 (N_16550,N_13586,N_14569);
xnor U16551 (N_16551,N_14963,N_10262);
xor U16552 (N_16552,N_11451,N_13024);
or U16553 (N_16553,N_10110,N_12672);
or U16554 (N_16554,N_11113,N_14417);
nor U16555 (N_16555,N_10447,N_14522);
or U16556 (N_16556,N_14976,N_13848);
xor U16557 (N_16557,N_14746,N_13845);
nand U16558 (N_16558,N_14192,N_12862);
and U16559 (N_16559,N_14462,N_12269);
and U16560 (N_16560,N_12384,N_14020);
xnor U16561 (N_16561,N_12145,N_14031);
or U16562 (N_16562,N_12160,N_10946);
and U16563 (N_16563,N_10876,N_14070);
nor U16564 (N_16564,N_12195,N_13499);
and U16565 (N_16565,N_11861,N_12848);
nor U16566 (N_16566,N_10765,N_11724);
xor U16567 (N_16567,N_13212,N_11749);
and U16568 (N_16568,N_14340,N_13519);
nand U16569 (N_16569,N_13737,N_12946);
nor U16570 (N_16570,N_10641,N_11086);
nand U16571 (N_16571,N_11421,N_12251);
xnor U16572 (N_16572,N_11852,N_14376);
xnor U16573 (N_16573,N_11853,N_11903);
xor U16574 (N_16574,N_11709,N_14947);
nand U16575 (N_16575,N_11351,N_12388);
and U16576 (N_16576,N_11054,N_11011);
nand U16577 (N_16577,N_14292,N_14762);
xnor U16578 (N_16578,N_13693,N_14081);
nand U16579 (N_16579,N_10519,N_12994);
xnor U16580 (N_16580,N_14719,N_14253);
nand U16581 (N_16581,N_10157,N_12343);
xnor U16582 (N_16582,N_13214,N_12117);
and U16583 (N_16583,N_13172,N_14465);
xnor U16584 (N_16584,N_14590,N_11089);
and U16585 (N_16585,N_10122,N_14210);
xor U16586 (N_16586,N_13185,N_12971);
or U16587 (N_16587,N_12943,N_10831);
and U16588 (N_16588,N_11344,N_10970);
and U16589 (N_16589,N_10705,N_13253);
or U16590 (N_16590,N_12564,N_14833);
nand U16591 (N_16591,N_12259,N_11222);
xor U16592 (N_16592,N_14797,N_11951);
xnor U16593 (N_16593,N_14857,N_12056);
and U16594 (N_16594,N_13641,N_13474);
xnor U16595 (N_16595,N_13713,N_14476);
nand U16596 (N_16596,N_10430,N_12754);
xor U16597 (N_16597,N_13096,N_14526);
and U16598 (N_16598,N_13076,N_14011);
or U16599 (N_16599,N_10112,N_12949);
xor U16600 (N_16600,N_11253,N_13087);
nand U16601 (N_16601,N_12878,N_14574);
nor U16602 (N_16602,N_11058,N_10273);
xor U16603 (N_16603,N_12227,N_12182);
and U16604 (N_16604,N_12193,N_12387);
xor U16605 (N_16605,N_13222,N_11518);
and U16606 (N_16606,N_11674,N_10738);
and U16607 (N_16607,N_12576,N_13937);
and U16608 (N_16608,N_12573,N_14167);
and U16609 (N_16609,N_13437,N_14535);
nor U16610 (N_16610,N_12980,N_13838);
or U16611 (N_16611,N_14842,N_12126);
and U16612 (N_16612,N_10272,N_12590);
and U16613 (N_16613,N_11098,N_11276);
nor U16614 (N_16614,N_12214,N_12496);
nor U16615 (N_16615,N_12009,N_11508);
and U16616 (N_16616,N_11201,N_10562);
and U16617 (N_16617,N_12272,N_11792);
and U16618 (N_16618,N_11976,N_14889);
or U16619 (N_16619,N_12243,N_10176);
and U16620 (N_16620,N_11629,N_11560);
and U16621 (N_16621,N_12385,N_10773);
xnor U16622 (N_16622,N_12383,N_11050);
and U16623 (N_16623,N_10300,N_12427);
or U16624 (N_16624,N_14384,N_10488);
and U16625 (N_16625,N_13887,N_14616);
nand U16626 (N_16626,N_10571,N_10341);
or U16627 (N_16627,N_12884,N_14817);
nor U16628 (N_16628,N_14993,N_11885);
xnor U16629 (N_16629,N_12382,N_12300);
xnor U16630 (N_16630,N_14079,N_10223);
or U16631 (N_16631,N_13842,N_12242);
or U16632 (N_16632,N_10688,N_11547);
nand U16633 (N_16633,N_12858,N_13277);
nand U16634 (N_16634,N_10757,N_14104);
nor U16635 (N_16635,N_14071,N_14510);
xor U16636 (N_16636,N_13496,N_13578);
or U16637 (N_16637,N_14320,N_12498);
or U16638 (N_16638,N_11928,N_14493);
nor U16639 (N_16639,N_11800,N_13584);
and U16640 (N_16640,N_11986,N_10506);
and U16641 (N_16641,N_10943,N_12315);
xor U16642 (N_16642,N_13996,N_11219);
nor U16643 (N_16643,N_12900,N_14053);
or U16644 (N_16644,N_11833,N_13302);
xor U16645 (N_16645,N_13345,N_11317);
nand U16646 (N_16646,N_12693,N_10813);
nor U16647 (N_16647,N_11902,N_12386);
nor U16648 (N_16648,N_10617,N_13300);
or U16649 (N_16649,N_13684,N_11554);
nand U16650 (N_16650,N_10400,N_13509);
xor U16651 (N_16651,N_12822,N_14068);
or U16652 (N_16652,N_11866,N_12865);
and U16653 (N_16653,N_10242,N_10077);
or U16654 (N_16654,N_12847,N_12159);
and U16655 (N_16655,N_13297,N_11886);
or U16656 (N_16656,N_11449,N_14207);
nand U16657 (N_16657,N_11265,N_12060);
nor U16658 (N_16658,N_11569,N_12700);
nand U16659 (N_16659,N_11499,N_12872);
xnor U16660 (N_16660,N_13982,N_11971);
nand U16661 (N_16661,N_11536,N_11412);
or U16662 (N_16662,N_13955,N_12526);
and U16663 (N_16663,N_12424,N_11254);
and U16664 (N_16664,N_12003,N_11476);
nand U16665 (N_16665,N_12886,N_14710);
nand U16666 (N_16666,N_14131,N_14323);
or U16667 (N_16667,N_14638,N_13511);
or U16668 (N_16668,N_11760,N_14110);
nor U16669 (N_16669,N_13875,N_13613);
and U16670 (N_16670,N_12491,N_10468);
nand U16671 (N_16671,N_10261,N_13788);
or U16672 (N_16672,N_11669,N_10665);
nor U16673 (N_16673,N_11939,N_12008);
nor U16674 (N_16674,N_11167,N_13043);
or U16675 (N_16675,N_14677,N_13976);
xnor U16676 (N_16676,N_13045,N_13233);
or U16677 (N_16677,N_14128,N_10279);
and U16678 (N_16678,N_14103,N_13188);
nor U16679 (N_16679,N_13778,N_12305);
nand U16680 (N_16680,N_13536,N_10388);
and U16681 (N_16681,N_12908,N_11868);
and U16682 (N_16682,N_12324,N_11491);
nor U16683 (N_16683,N_11244,N_10162);
xnor U16684 (N_16684,N_10065,N_10109);
and U16685 (N_16685,N_14431,N_10282);
nor U16686 (N_16686,N_13025,N_10550);
or U16687 (N_16687,N_11194,N_12652);
or U16688 (N_16688,N_12051,N_14926);
or U16689 (N_16689,N_12768,N_10401);
or U16690 (N_16690,N_11628,N_10031);
nand U16691 (N_16691,N_12130,N_12795);
or U16692 (N_16692,N_14680,N_14771);
xor U16693 (N_16693,N_12037,N_13304);
and U16694 (N_16694,N_13394,N_11056);
or U16695 (N_16695,N_12876,N_14999);
nand U16696 (N_16696,N_14039,N_11948);
nand U16697 (N_16697,N_10516,N_14386);
nor U16698 (N_16698,N_12737,N_14808);
nand U16699 (N_16699,N_14149,N_12633);
nand U16700 (N_16700,N_14601,N_14524);
nor U16701 (N_16701,N_14295,N_13337);
nor U16702 (N_16702,N_14732,N_13105);
or U16703 (N_16703,N_11898,N_13344);
and U16704 (N_16704,N_13453,N_14846);
and U16705 (N_16705,N_13666,N_10322);
and U16706 (N_16706,N_13205,N_14506);
or U16707 (N_16707,N_11890,N_11757);
nor U16708 (N_16708,N_12591,N_13585);
nor U16709 (N_16709,N_12146,N_11281);
nand U16710 (N_16710,N_11073,N_10035);
nor U16711 (N_16711,N_12679,N_14228);
nand U16712 (N_16712,N_11309,N_11565);
nor U16713 (N_16713,N_10642,N_10637);
nand U16714 (N_16714,N_12007,N_14861);
or U16715 (N_16715,N_12536,N_12478);
or U16716 (N_16716,N_11644,N_14916);
xnor U16717 (N_16717,N_11798,N_14074);
nor U16718 (N_16718,N_12645,N_11215);
xor U16719 (N_16719,N_12702,N_11486);
xor U16720 (N_16720,N_13634,N_12377);
nor U16721 (N_16721,N_10589,N_10901);
xnor U16722 (N_16722,N_11715,N_14113);
or U16723 (N_16723,N_10828,N_11066);
and U16724 (N_16724,N_14134,N_12867);
nand U16725 (N_16725,N_12363,N_12110);
xnor U16726 (N_16726,N_13239,N_11586);
nor U16727 (N_16727,N_12471,N_12298);
or U16728 (N_16728,N_14261,N_10132);
or U16729 (N_16729,N_14630,N_13338);
nand U16730 (N_16730,N_10493,N_11277);
nor U16731 (N_16731,N_14121,N_12763);
or U16732 (N_16732,N_13873,N_14934);
and U16733 (N_16733,N_11226,N_11473);
or U16734 (N_16734,N_12099,N_12402);
nand U16735 (N_16735,N_12660,N_10328);
and U16736 (N_16736,N_11019,N_12413);
and U16737 (N_16737,N_13090,N_13769);
and U16738 (N_16738,N_14774,N_12334);
nor U16739 (N_16739,N_10764,N_11766);
nand U16740 (N_16740,N_10905,N_11229);
nor U16741 (N_16741,N_12127,N_11721);
nand U16742 (N_16742,N_13216,N_11240);
nand U16743 (N_16743,N_10730,N_10530);
nor U16744 (N_16744,N_10707,N_12877);
and U16745 (N_16745,N_10302,N_10527);
nand U16746 (N_16746,N_14652,N_14241);
nor U16747 (N_16747,N_11892,N_13192);
xnor U16748 (N_16748,N_10189,N_12440);
and U16749 (N_16749,N_10534,N_13913);
or U16750 (N_16750,N_12903,N_10716);
nor U16751 (N_16751,N_14671,N_10891);
or U16752 (N_16752,N_10890,N_14061);
nor U16753 (N_16753,N_11136,N_13614);
or U16754 (N_16754,N_14223,N_10984);
and U16755 (N_16755,N_14587,N_11036);
and U16756 (N_16756,N_12643,N_12366);
nor U16757 (N_16757,N_14702,N_10969);
and U16758 (N_16758,N_14484,N_14871);
nor U16759 (N_16759,N_13606,N_11595);
xnor U16760 (N_16760,N_14276,N_11733);
or U16761 (N_16761,N_11872,N_13138);
or U16762 (N_16762,N_13458,N_10851);
or U16763 (N_16763,N_13117,N_11602);
or U16764 (N_16764,N_11867,N_13985);
xnor U16765 (N_16765,N_13625,N_14180);
or U16766 (N_16766,N_13352,N_11213);
and U16767 (N_16767,N_14844,N_14184);
xnor U16768 (N_16768,N_11730,N_11367);
nand U16769 (N_16769,N_11521,N_14521);
or U16770 (N_16770,N_13732,N_12709);
nor U16771 (N_16771,N_10694,N_12711);
and U16772 (N_16772,N_11623,N_12508);
nand U16773 (N_16773,N_11212,N_12142);
or U16774 (N_16774,N_12436,N_14033);
nor U16775 (N_16775,N_14221,N_10919);
nand U16776 (N_16776,N_12322,N_14272);
xnor U16777 (N_16777,N_12675,N_12703);
and U16778 (N_16778,N_13010,N_11947);
xor U16779 (N_16779,N_14157,N_13978);
nand U16780 (N_16780,N_11707,N_11075);
or U16781 (N_16781,N_11755,N_13285);
and U16782 (N_16782,N_10054,N_13026);
xnor U16783 (N_16783,N_14755,N_12941);
and U16784 (N_16784,N_12823,N_14318);
xor U16785 (N_16785,N_11013,N_13944);
and U16786 (N_16786,N_12329,N_10582);
and U16787 (N_16787,N_12477,N_10793);
xnor U16788 (N_16788,N_12460,N_13291);
and U16789 (N_16789,N_13145,N_10635);
and U16790 (N_16790,N_12504,N_11738);
or U16791 (N_16791,N_11206,N_14902);
or U16792 (N_16792,N_11992,N_14156);
nand U16793 (N_16793,N_13379,N_13533);
or U16794 (N_16794,N_11333,N_12328);
or U16795 (N_16795,N_13467,N_13949);
nand U16796 (N_16796,N_11370,N_13940);
nor U16797 (N_16797,N_13211,N_12625);
xor U16798 (N_16798,N_12517,N_10653);
nor U16799 (N_16799,N_10538,N_14024);
xor U16800 (N_16800,N_11258,N_13005);
xnor U16801 (N_16801,N_14967,N_12364);
nand U16802 (N_16802,N_11029,N_10142);
or U16803 (N_16803,N_14097,N_11283);
xor U16804 (N_16804,N_10539,N_11799);
nand U16805 (N_16805,N_14047,N_13455);
xor U16806 (N_16806,N_12792,N_11484);
or U16807 (N_16807,N_12825,N_12374);
nand U16808 (N_16808,N_10763,N_11124);
xnor U16809 (N_16809,N_12930,N_10825);
and U16810 (N_16810,N_11256,N_12468);
and U16811 (N_16811,N_14327,N_11780);
and U16812 (N_16812,N_14101,N_12989);
xor U16813 (N_16813,N_11815,N_11300);
xor U16814 (N_16814,N_10990,N_14293);
or U16815 (N_16815,N_11198,N_12844);
and U16816 (N_16816,N_12602,N_10246);
nor U16817 (N_16817,N_11698,N_13706);
nand U16818 (N_16818,N_10134,N_11310);
xor U16819 (N_16819,N_11594,N_13404);
nor U16820 (N_16820,N_14335,N_12121);
or U16821 (N_16821,N_12925,N_13305);
nor U16822 (N_16822,N_11763,N_12027);
nand U16823 (N_16823,N_14892,N_12705);
and U16824 (N_16824,N_10918,N_10277);
xnor U16825 (N_16825,N_11109,N_11227);
and U16826 (N_16826,N_10353,N_12304);
and U16827 (N_16827,N_12464,N_14025);
and U16828 (N_16828,N_13151,N_10082);
or U16829 (N_16829,N_12853,N_12541);
nor U16830 (N_16830,N_14836,N_12070);
nor U16831 (N_16831,N_14779,N_14382);
nand U16832 (N_16832,N_13038,N_14888);
or U16833 (N_16833,N_11190,N_11180);
nor U16834 (N_16834,N_14169,N_10668);
xor U16835 (N_16835,N_14175,N_11267);
and U16836 (N_16836,N_13643,N_12816);
or U16837 (N_16837,N_14566,N_10061);
and U16838 (N_16838,N_13633,N_11433);
or U16839 (N_16839,N_10473,N_10088);
or U16840 (N_16840,N_12444,N_13880);
nor U16841 (N_16841,N_11795,N_12109);
nand U16842 (N_16842,N_14883,N_10501);
xor U16843 (N_16843,N_12599,N_12474);
or U16844 (N_16844,N_12241,N_13369);
or U16845 (N_16845,N_13583,N_11203);
nor U16846 (N_16846,N_13503,N_11666);
nor U16847 (N_16847,N_10995,N_12250);
and U16848 (N_16848,N_12983,N_10367);
and U16849 (N_16849,N_10575,N_11854);
and U16850 (N_16850,N_12481,N_14418);
nand U16851 (N_16851,N_13967,N_14034);
or U16852 (N_16852,N_13876,N_14543);
and U16853 (N_16853,N_12845,N_10098);
xor U16854 (N_16854,N_12699,N_12274);
or U16855 (N_16855,N_14879,N_10897);
and U16856 (N_16856,N_10329,N_10096);
nor U16857 (N_16857,N_12005,N_14016);
nand U16858 (N_16858,N_11881,N_13047);
nand U16859 (N_16859,N_10802,N_12942);
nor U16860 (N_16860,N_11104,N_11146);
nor U16861 (N_16861,N_12231,N_10867);
xor U16862 (N_16862,N_12225,N_12457);
nand U16863 (N_16863,N_11087,N_10319);
xnor U16864 (N_16864,N_11502,N_11046);
xnor U16865 (N_16865,N_10221,N_10584);
and U16866 (N_16866,N_12187,N_10651);
xor U16867 (N_16867,N_13136,N_12203);
xor U16868 (N_16868,N_14822,N_14730);
or U16869 (N_16869,N_10429,N_10839);
and U16870 (N_16870,N_14487,N_14088);
nor U16871 (N_16871,N_10724,N_13697);
nor U16872 (N_16872,N_14863,N_11671);
or U16873 (N_16873,N_11982,N_12167);
nand U16874 (N_16874,N_13834,N_14473);
or U16875 (N_16875,N_10655,N_14673);
nor U16876 (N_16876,N_14437,N_12098);
or U16877 (N_16877,N_10932,N_14685);
xnor U16878 (N_16878,N_14735,N_12611);
nor U16879 (N_16879,N_11997,N_14700);
nand U16880 (N_16880,N_12990,N_11696);
and U16881 (N_16881,N_10944,N_12204);
nor U16882 (N_16882,N_13579,N_13679);
and U16883 (N_16883,N_14552,N_13420);
and U16884 (N_16884,N_13782,N_13695);
xnor U16885 (N_16885,N_11916,N_12882);
xnor U16886 (N_16886,N_14768,N_10453);
or U16887 (N_16887,N_12493,N_13989);
and U16888 (N_16888,N_12745,N_11844);
and U16889 (N_16889,N_14422,N_13879);
and U16890 (N_16890,N_13654,N_12636);
or U16891 (N_16891,N_10503,N_14641);
nor U16892 (N_16892,N_14495,N_12311);
nor U16893 (N_16893,N_11899,N_12135);
or U16894 (N_16894,N_13652,N_10537);
nand U16895 (N_16895,N_10340,N_11078);
or U16896 (N_16896,N_14291,N_11940);
or U16897 (N_16897,N_13284,N_13504);
nand U16898 (N_16898,N_13140,N_13150);
and U16899 (N_16899,N_14501,N_12188);
nand U16900 (N_16900,N_11385,N_13754);
nand U16901 (N_16901,N_14548,N_11286);
xor U16902 (N_16902,N_13961,N_10103);
nor U16903 (N_16903,N_14699,N_11970);
and U16904 (N_16904,N_14084,N_13459);
nor U16905 (N_16905,N_10933,N_11912);
nor U16906 (N_16906,N_11123,N_13647);
and U16907 (N_16907,N_10210,N_11609);
nor U16908 (N_16908,N_14124,N_13075);
xnor U16909 (N_16909,N_11059,N_12899);
nand U16910 (N_16910,N_11831,N_12803);
nand U16911 (N_16911,N_11490,N_10703);
nand U16912 (N_16912,N_14572,N_12765);
or U16913 (N_16913,N_13902,N_11306);
nand U16914 (N_16914,N_10895,N_12742);
and U16915 (N_16915,N_14120,N_13670);
xor U16916 (N_16916,N_13987,N_10838);
nand U16917 (N_16917,N_11914,N_13247);
and U16918 (N_16918,N_14628,N_14620);
and U16919 (N_16919,N_13392,N_14282);
nor U16920 (N_16920,N_14069,N_11120);
nor U16921 (N_16921,N_14471,N_14370);
or U16922 (N_16922,N_12973,N_12704);
nand U16923 (N_16923,N_12936,N_13506);
xnor U16924 (N_16924,N_12528,N_13388);
or U16925 (N_16925,N_10422,N_10929);
xor U16926 (N_16926,N_14267,N_14406);
or U16927 (N_16927,N_13204,N_14985);
or U16928 (N_16928,N_13264,N_12609);
or U16929 (N_16929,N_12503,N_14958);
nand U16930 (N_16930,N_11826,N_14132);
xor U16931 (N_16931,N_14556,N_13977);
nand U16932 (N_16932,N_12527,N_10699);
xnor U16933 (N_16933,N_10692,N_10045);
and U16934 (N_16934,N_10996,N_13609);
and U16935 (N_16935,N_11936,N_14248);
nand U16936 (N_16936,N_11114,N_13161);
nand U16937 (N_16937,N_11365,N_13818);
xnor U16938 (N_16938,N_12370,N_13180);
nand U16939 (N_16939,N_14570,N_13700);
nand U16940 (N_16940,N_13469,N_14325);
or U16941 (N_16941,N_10832,N_11897);
and U16942 (N_16942,N_12553,N_14154);
and U16943 (N_16943,N_10854,N_10956);
nand U16944 (N_16944,N_10312,N_14921);
or U16945 (N_16945,N_12088,N_14545);
and U16946 (N_16946,N_13066,N_12905);
nor U16947 (N_16947,N_12552,N_10680);
nand U16948 (N_16948,N_10062,N_11840);
xnor U16949 (N_16949,N_11438,N_12969);
or U16950 (N_16950,N_14067,N_13171);
xor U16951 (N_16951,N_13425,N_10017);
xnor U16952 (N_16952,N_11102,N_10477);
nand U16953 (N_16953,N_13450,N_11399);
or U16954 (N_16954,N_14851,N_11217);
and U16955 (N_16955,N_11905,N_11083);
nor U16956 (N_16956,N_14726,N_11290);
nand U16957 (N_16957,N_10822,N_11975);
or U16958 (N_16958,N_14441,N_10152);
nand U16959 (N_16959,N_10732,N_13243);
xor U16960 (N_16960,N_14751,N_11550);
xor U16961 (N_16961,N_10529,N_13817);
and U16962 (N_16962,N_13690,N_12431);
xnor U16963 (N_16963,N_11017,N_14226);
nor U16964 (N_16964,N_10947,N_13526);
xnor U16965 (N_16965,N_13217,N_13461);
nor U16966 (N_16966,N_12649,N_14964);
xor U16967 (N_16967,N_13559,N_12773);
or U16968 (N_16968,N_10253,N_14123);
xor U16969 (N_16969,N_12422,N_12721);
and U16970 (N_16970,N_13099,N_10050);
xnor U16971 (N_16971,N_10230,N_10526);
nor U16972 (N_16972,N_10220,N_12321);
nor U16973 (N_16973,N_13298,N_12197);
nand U16974 (N_16974,N_13698,N_11849);
xor U16975 (N_16975,N_12323,N_12749);
nor U16976 (N_16976,N_10504,N_10691);
nand U16977 (N_16977,N_13883,N_10659);
nor U16978 (N_16978,N_13864,N_12921);
xnor U16979 (N_16979,N_12408,N_12342);
xor U16980 (N_16980,N_14971,N_10830);
xor U16981 (N_16981,N_13822,N_14679);
and U16982 (N_16982,N_13381,N_14597);
nor U16983 (N_16983,N_14887,N_12759);
xor U16984 (N_16984,N_14951,N_12683);
xor U16985 (N_16985,N_11558,N_13272);
or U16986 (N_16986,N_11679,N_13664);
xnor U16987 (N_16987,N_11710,N_12054);
and U16988 (N_16988,N_13008,N_14695);
nor U16989 (N_16989,N_12578,N_12279);
or U16990 (N_16990,N_11588,N_10631);
and U16991 (N_16991,N_10016,N_10013);
nor U16992 (N_16992,N_14085,N_13128);
and U16993 (N_16993,N_11363,N_12202);
nand U16994 (N_16994,N_10740,N_11504);
xnor U16995 (N_16995,N_14982,N_11030);
xor U16996 (N_16996,N_14312,N_14664);
nor U16997 (N_16997,N_14364,N_11170);
or U16998 (N_16998,N_14922,N_10085);
xnor U16999 (N_16999,N_14537,N_13753);
or U17000 (N_17000,N_14279,N_11705);
xor U17001 (N_17001,N_13787,N_11566);
and U17002 (N_17002,N_11827,N_14613);
nand U17003 (N_17003,N_12890,N_10382);
xnor U17004 (N_17004,N_11667,N_11496);
xor U17005 (N_17005,N_14737,N_10185);
nand U17006 (N_17006,N_12802,N_13768);
xnor U17007 (N_17007,N_10786,N_13621);
or U17008 (N_17008,N_14869,N_11171);
and U17009 (N_17009,N_10499,N_12394);
nand U17010 (N_17010,N_13380,N_12608);
and U17011 (N_17011,N_11200,N_10046);
xor U17012 (N_17012,N_14307,N_10657);
nor U17013 (N_17013,N_12624,N_11128);
xor U17014 (N_17014,N_10141,N_10939);
and U17015 (N_17015,N_11088,N_12629);
xor U17016 (N_17016,N_13490,N_10746);
nand U17017 (N_17017,N_13326,N_13112);
or U17018 (N_17018,N_10032,N_13286);
and U17019 (N_17019,N_10925,N_10713);
or U17020 (N_17020,N_10146,N_12317);
and U17021 (N_17021,N_13418,N_11488);
xnor U17022 (N_17022,N_12170,N_14146);
nand U17023 (N_17023,N_13446,N_11526);
nand U17024 (N_17024,N_14144,N_12534);
and U17025 (N_17025,N_13036,N_14286);
nand U17026 (N_17026,N_10729,N_13335);
nand U17027 (N_17027,N_13373,N_14662);
and U17028 (N_17028,N_12404,N_13323);
nor U17029 (N_17029,N_13421,N_10742);
nor U17030 (N_17030,N_11322,N_12680);
and U17031 (N_17031,N_11494,N_13184);
or U17032 (N_17032,N_14684,N_12292);
or U17033 (N_17033,N_13057,N_14640);
xor U17034 (N_17034,N_14127,N_14479);
nand U17035 (N_17035,N_14393,N_14575);
or U17036 (N_17036,N_12615,N_10673);
xor U17037 (N_17037,N_10780,N_14697);
or U17038 (N_17038,N_14229,N_14500);
or U17039 (N_17039,N_11505,N_11445);
nor U17040 (N_17040,N_13642,N_14233);
xnor U17041 (N_17041,N_12456,N_12447);
or U17042 (N_17042,N_11714,N_13872);
or U17043 (N_17043,N_13435,N_13397);
nand U17044 (N_17044,N_13804,N_10416);
nor U17045 (N_17045,N_13206,N_10788);
xor U17046 (N_17046,N_14930,N_14075);
or U17047 (N_17047,N_10745,N_14667);
nor U17048 (N_17048,N_11593,N_11546);
or U17049 (N_17049,N_14642,N_13174);
or U17050 (N_17050,N_10177,N_12834);
and U17051 (N_17051,N_11143,N_14264);
and U17052 (N_17052,N_14289,N_13847);
or U17053 (N_17053,N_12722,N_12131);
nand U17054 (N_17054,N_14319,N_12774);
xnor U17055 (N_17055,N_12567,N_13361);
nand U17056 (N_17056,N_10386,N_11401);
nand U17057 (N_17057,N_12354,N_14331);
nor U17058 (N_17058,N_12332,N_13168);
or U17059 (N_17059,N_14488,N_13416);
xor U17060 (N_17060,N_11191,N_12565);
nor U17061 (N_17061,N_12093,N_12912);
and U17062 (N_17062,N_14785,N_11032);
and U17063 (N_17063,N_14015,N_10795);
nand U17064 (N_17064,N_12263,N_13083);
xnor U17065 (N_17065,N_14314,N_12105);
nand U17066 (N_17066,N_14273,N_13636);
or U17067 (N_17067,N_10677,N_11358);
nor U17068 (N_17068,N_11155,N_12824);
nor U17069 (N_17069,N_12986,N_11814);
or U17070 (N_17070,N_11711,N_12409);
nor U17071 (N_17071,N_14832,N_11875);
and U17072 (N_17072,N_10751,N_11906);
nand U17073 (N_17073,N_11061,N_11016);
xor U17074 (N_17074,N_10445,N_10775);
xor U17075 (N_17075,N_14369,N_12026);
xnor U17076 (N_17076,N_13552,N_11419);
xor U17077 (N_17077,N_14238,N_10459);
or U17078 (N_17078,N_11533,N_12059);
nand U17079 (N_17079,N_12011,N_12352);
nor U17080 (N_17080,N_11079,N_10457);
nand U17081 (N_17081,N_10559,N_14812);
or U17082 (N_17082,N_11603,N_13721);
nand U17083 (N_17083,N_11779,N_12657);
nand U17084 (N_17084,N_14374,N_14942);
nand U17085 (N_17085,N_11777,N_10204);
nand U17086 (N_17086,N_14598,N_13738);
nand U17087 (N_17087,N_11169,N_11974);
or U17088 (N_17088,N_11828,N_10443);
and U17089 (N_17089,N_13825,N_13052);
and U17090 (N_17090,N_14899,N_14161);
and U17091 (N_17091,N_14955,N_11479);
xnor U17092 (N_17092,N_13534,N_14571);
and U17093 (N_17093,N_11145,N_11726);
xnor U17094 (N_17094,N_10372,N_12396);
xnor U17095 (N_17095,N_11458,N_13349);
xnor U17096 (N_17096,N_13960,N_14205);
nor U17097 (N_17097,N_12036,N_10761);
nor U17098 (N_17098,N_13688,N_10515);
xnor U17099 (N_17099,N_12128,N_14560);
nand U17100 (N_17100,N_10776,N_10248);
xnor U17101 (N_17101,N_10469,N_13389);
nand U17102 (N_17102,N_12810,N_10476);
nand U17103 (N_17103,N_12975,N_12467);
nor U17104 (N_17104,N_12013,N_10001);
or U17105 (N_17105,N_11647,N_14481);
and U17106 (N_17106,N_12842,N_11275);
or U17107 (N_17107,N_11765,N_10362);
xor U17108 (N_17108,N_12610,N_14125);
xnor U17109 (N_17109,N_12104,N_11135);
or U17110 (N_17110,N_11719,N_13260);
and U17111 (N_17111,N_13331,N_14681);
nor U17112 (N_17112,N_10743,N_11461);
or U17113 (N_17113,N_10735,N_11841);
xor U17114 (N_17114,N_11440,N_12648);
and U17115 (N_17115,N_10887,N_13293);
nor U17116 (N_17116,N_10850,N_13946);
or U17117 (N_17117,N_10913,N_11340);
or U17118 (N_17118,N_12509,N_13131);
xor U17119 (N_17119,N_12529,N_12158);
xnor U17120 (N_17120,N_14819,N_10198);
or U17121 (N_17121,N_12116,N_13215);
nor U17122 (N_17122,N_12184,N_12963);
nor U17123 (N_17123,N_12623,N_14036);
nor U17124 (N_17124,N_13962,N_13137);
or U17125 (N_17125,N_11596,N_11589);
nand U17126 (N_17126,N_12420,N_10275);
nand U17127 (N_17127,N_11417,N_14371);
nor U17128 (N_17128,N_13546,N_10971);
or U17129 (N_17129,N_11455,N_10536);
or U17130 (N_17130,N_14001,N_11878);
nor U17131 (N_17131,N_10604,N_12559);
nand U17132 (N_17132,N_13789,N_12577);
nor U17133 (N_17133,N_11404,N_12719);
nor U17134 (N_17134,N_14966,N_10610);
xnor U17135 (N_17135,N_14139,N_10048);
nand U17136 (N_17136,N_14945,N_13580);
xor U17137 (N_17137,N_13287,N_10646);
xnor U17138 (N_17138,N_10664,N_13189);
or U17139 (N_17139,N_13426,N_12996);
nor U17140 (N_17140,N_13410,N_13028);
xor U17141 (N_17141,N_14398,N_14580);
nand U17142 (N_17142,N_14873,N_13431);
or U17143 (N_17143,N_14739,N_13027);
nand U17144 (N_17144,N_10186,N_13683);
nor U17145 (N_17145,N_13413,N_11545);
or U17146 (N_17146,N_11557,N_11291);
nor U17147 (N_17147,N_13236,N_10487);
and U17148 (N_17148,N_14459,N_11964);
nor U17149 (N_17149,N_12042,N_12909);
or U17150 (N_17150,N_14907,N_13992);
nor U17151 (N_17151,N_13678,N_14414);
nand U17152 (N_17152,N_12297,N_13767);
or U17153 (N_17153,N_14960,N_10327);
and U17154 (N_17154,N_10426,N_12979);
nor U17155 (N_17155,N_11179,N_13094);
nor U17156 (N_17156,N_10249,N_12014);
and U17157 (N_17157,N_14066,N_12694);
nor U17158 (N_17158,N_14761,N_12598);
nor U17159 (N_17159,N_14712,N_10910);
or U17160 (N_17160,N_10723,N_10495);
or U17161 (N_17161,N_13566,N_13918);
nand U17162 (N_17162,N_12416,N_11984);
nor U17163 (N_17163,N_13084,N_10404);
and U17164 (N_17164,N_12372,N_11678);
nand U17165 (N_17165,N_14908,N_10846);
xnor U17166 (N_17166,N_13384,N_14449);
nand U17167 (N_17167,N_10294,N_13925);
xnor U17168 (N_17168,N_14256,N_10636);
nor U17169 (N_17169,N_14356,N_10151);
nor U17170 (N_17170,N_14992,N_13797);
xnor U17171 (N_17171,N_10323,N_10043);
or U17172 (N_17172,N_11620,N_12465);
or U17173 (N_17173,N_13936,N_11904);
xor U17174 (N_17174,N_13322,N_11081);
nand U17175 (N_17175,N_14711,N_13412);
or U17176 (N_17176,N_11616,N_11060);
nand U17177 (N_17177,N_11614,N_11927);
xnor U17178 (N_17178,N_14007,N_14742);
nand U17179 (N_17179,N_10843,N_10574);
nand U17180 (N_17180,N_13964,N_10263);
xor U17181 (N_17181,N_14359,N_13574);
and U17182 (N_17182,N_13891,N_11805);
nand U17183 (N_17183,N_13278,N_13669);
xor U17184 (N_17184,N_13508,N_12449);
or U17185 (N_17185,N_11702,N_14520);
nand U17186 (N_17186,N_10634,N_10299);
or U17187 (N_17187,N_14943,N_14436);
or U17188 (N_17188,N_11576,N_14326);
xor U17189 (N_17189,N_12780,N_14224);
or U17190 (N_17190,N_10489,N_10180);
xor U17191 (N_17191,N_13567,N_14379);
nand U17192 (N_17192,N_10807,N_12232);
nor U17193 (N_17193,N_10359,N_14383);
nor U17194 (N_17194,N_12999,N_11273);
nand U17195 (N_17195,N_10004,N_11790);
nand U17196 (N_17196,N_13781,N_14547);
nor U17197 (N_17197,N_14725,N_11202);
nand U17198 (N_17198,N_13514,N_11531);
nand U17199 (N_17199,N_13471,N_14373);
and U17200 (N_17200,N_12910,N_11459);
xnor U17201 (N_17201,N_11660,N_13959);
nor U17202 (N_17202,N_14108,N_13353);
nand U17203 (N_17203,N_12747,N_14162);
and U17204 (N_17204,N_11767,N_13851);
or U17205 (N_17205,N_13343,N_13265);
xnor U17206 (N_17206,N_12419,N_13317);
nor U17207 (N_17207,N_13582,N_10179);
nand U17208 (N_17208,N_14388,N_13764);
nor U17209 (N_17209,N_14933,N_14885);
nor U17210 (N_17210,N_14688,N_13170);
and U17211 (N_17211,N_12561,N_14054);
or U17212 (N_17212,N_14626,N_14691);
and U17213 (N_17213,N_14305,N_12340);
nor U17214 (N_17214,N_14214,N_14733);
nor U17215 (N_17215,N_12044,N_14532);
and U17216 (N_17216,N_11354,N_12666);
or U17217 (N_17217,N_10084,N_11189);
nor U17218 (N_17218,N_13263,N_11929);
xor U17219 (N_17219,N_14782,N_13334);
xnor U17220 (N_17220,N_12230,N_13100);
or U17221 (N_17221,N_13619,N_13144);
nor U17222 (N_17222,N_13308,N_14576);
or U17223 (N_17223,N_11409,N_11701);
xnor U17224 (N_17224,N_13315,N_13134);
nand U17225 (N_17225,N_13015,N_10022);
or U17226 (N_17226,N_14965,N_11725);
xor U17227 (N_17227,N_11953,N_10435);
xnor U17228 (N_17228,N_11420,N_14727);
nor U17229 (N_17229,N_12806,N_13115);
and U17230 (N_17230,N_10663,N_13190);
nand U17231 (N_17231,N_10731,N_12962);
and U17232 (N_17232,N_12965,N_13398);
xor U17233 (N_17233,N_10078,N_14905);
or U17234 (N_17234,N_14009,N_14301);
or U17235 (N_17235,N_12678,N_10377);
xnor U17236 (N_17236,N_10759,N_11582);
nand U17237 (N_17237,N_14969,N_10094);
nand U17238 (N_17238,N_12124,N_10951);
or U17239 (N_17239,N_14440,N_10171);
nand U17240 (N_17240,N_12612,N_12849);
nor U17241 (N_17241,N_13723,N_14442);
nand U17242 (N_17242,N_14032,N_13116);
and U17243 (N_17243,N_13844,N_13356);
nand U17244 (N_17244,N_10225,N_11234);
xnor U17245 (N_17245,N_11517,N_10772);
xor U17246 (N_17246,N_13018,N_12393);
or U17247 (N_17247,N_12091,N_13279);
nand U17248 (N_17248,N_10815,N_10431);
nand U17249 (N_17249,N_14343,N_13254);
and U17250 (N_17250,N_11522,N_13661);
and U17251 (N_17251,N_14841,N_14891);
and U17252 (N_17252,N_13154,N_11962);
or U17253 (N_17253,N_11355,N_10974);
and U17254 (N_17254,N_11471,N_11742);
nor U17255 (N_17255,N_14258,N_10695);
nand U17256 (N_17256,N_11196,N_10513);
xor U17257 (N_17257,N_11346,N_11894);
and U17258 (N_17258,N_11386,N_11895);
and U17259 (N_17259,N_10414,N_14714);
and U17260 (N_17260,N_10583,N_12684);
xnor U17261 (N_17261,N_12677,N_11035);
xnor U17262 (N_17262,N_14196,N_14046);
xnor U17263 (N_17263,N_13999,N_11466);
xor U17264 (N_17264,N_12551,N_10863);
nor U17265 (N_17265,N_13072,N_12454);
nor U17266 (N_17266,N_10081,N_12887);
and U17267 (N_17267,N_13861,N_12157);
nand U17268 (N_17268,N_12681,N_10614);
xor U17269 (N_17269,N_11579,N_12406);
nand U17270 (N_17270,N_10284,N_11510);
nand U17271 (N_17271,N_13952,N_10402);
xor U17272 (N_17272,N_10945,N_13892);
nand U17273 (N_17273,N_14277,N_10847);
or U17274 (N_17274,N_12883,N_10446);
nand U17275 (N_17275,N_14731,N_11680);
nand U17276 (N_17276,N_12266,N_14452);
or U17277 (N_17277,N_14665,N_13149);
and U17278 (N_17278,N_10379,N_10714);
nor U17279 (N_17279,N_12429,N_13810);
nor U17280 (N_17280,N_11655,N_14257);
and U17281 (N_17281,N_13762,N_13809);
xnor U17282 (N_17282,N_13132,N_13167);
nand U17283 (N_17283,N_13739,N_14227);
and U17284 (N_17284,N_14160,N_12089);
nand U17285 (N_17285,N_11988,N_12744);
nor U17286 (N_17286,N_11441,N_13906);
nor U17287 (N_17287,N_10339,N_10886);
or U17288 (N_17288,N_10502,N_13408);
nand U17289 (N_17289,N_10097,N_12786);
xnor U17290 (N_17290,N_13558,N_14799);
xnor U17291 (N_17291,N_14767,N_13449);
xnor U17292 (N_17292,N_13749,N_11049);
nand U17293 (N_17293,N_13126,N_11280);
or U17294 (N_17294,N_12606,N_12630);
nand U17295 (N_17295,N_14245,N_11043);
xnor U17296 (N_17296,N_11026,N_12490);
and U17297 (N_17297,N_11002,N_14862);
xor U17298 (N_17298,N_13704,N_12233);
nor U17299 (N_17299,N_11080,N_13628);
or U17300 (N_17300,N_11464,N_10149);
and U17301 (N_17301,N_10101,N_14489);
nor U17302 (N_17302,N_12776,N_12592);
and U17303 (N_17303,N_13451,N_13240);
and U17304 (N_17304,N_10332,N_11520);
nor U17305 (N_17305,N_12596,N_12538);
nand U17306 (N_17306,N_12706,N_13130);
xnor U17307 (N_17307,N_14005,N_12200);
or U17308 (N_17308,N_10924,N_10950);
nor U17309 (N_17309,N_14358,N_13139);
nand U17310 (N_17310,N_10315,N_10155);
nor U17311 (N_17311,N_13061,N_12904);
xor U17312 (N_17312,N_13850,N_13209);
xor U17313 (N_17313,N_10357,N_11444);
and U17314 (N_17314,N_11693,N_11587);
or U17315 (N_17315,N_14218,N_14035);
xnor U17316 (N_17316,N_14656,N_12917);
and U17317 (N_17317,N_12482,N_14527);
and U17318 (N_17318,N_12086,N_12659);
and U17319 (N_17319,N_14403,N_11913);
xnor U17320 (N_17320,N_13473,N_11478);
xnor U17321 (N_17321,N_10661,N_11205);
nand U17322 (N_17322,N_12192,N_13200);
and U17323 (N_17323,N_14611,N_13360);
nand U17324 (N_17324,N_10603,N_12524);
nand U17325 (N_17325,N_11187,N_11920);
or U17326 (N_17326,N_14666,N_12179);
and U17327 (N_17327,N_13639,N_14820);
xnor U17328 (N_17328,N_12207,N_12671);
xnor U17329 (N_17329,N_10409,N_10396);
or U17330 (N_17330,N_11882,N_12530);
nor U17331 (N_17331,N_14048,N_12764);
and U17332 (N_17332,N_13261,N_10977);
nand U17333 (N_17333,N_14073,N_12662);
or U17334 (N_17334,N_14299,N_11956);
nor U17335 (N_17335,N_13863,N_14083);
or U17336 (N_17336,N_12492,N_13350);
nand U17337 (N_17337,N_12190,N_14986);
nand U17338 (N_17338,N_10316,N_10411);
nor U17339 (N_17339,N_14777,N_14918);
nand U17340 (N_17340,N_10161,N_11668);
nor U17341 (N_17341,N_12229,N_14929);
nor U17342 (N_17342,N_14800,N_10774);
and U17343 (N_17343,N_11684,N_13521);
nand U17344 (N_17344,N_12338,N_13807);
nor U17345 (N_17345,N_13445,N_12725);
or U17346 (N_17346,N_10821,N_13501);
nor U17347 (N_17347,N_12701,N_10999);
xor U17348 (N_17348,N_12476,N_14867);
and U17349 (N_17349,N_14579,N_13118);
nand U17350 (N_17350,N_11556,N_10814);
and U17351 (N_17351,N_11773,N_14251);
and U17352 (N_17352,N_10140,N_14997);
xor U17353 (N_17353,N_12929,N_13194);
nor U17354 (N_17354,N_11142,N_13758);
nand U17355 (N_17355,N_12655,N_14093);
nand U17356 (N_17356,N_11446,N_14480);
xnor U17357 (N_17357,N_10369,N_11925);
nand U17358 (N_17358,N_13468,N_12984);
xnor U17359 (N_17359,N_13366,N_10968);
nor U17360 (N_17360,N_13907,N_14194);
nor U17361 (N_17361,N_10444,N_14928);
nor U17362 (N_17362,N_10873,N_12282);
and U17363 (N_17363,N_10481,N_11012);
or U17364 (N_17364,N_14927,N_13109);
or U17365 (N_17365,N_10671,N_12084);
nand U17366 (N_17366,N_13042,N_10808);
or U17367 (N_17367,N_14365,N_10227);
nand U17368 (N_17368,N_14140,N_14619);
nand U17369 (N_17369,N_12213,N_11825);
xor U17370 (N_17370,N_14758,N_10994);
nor U17371 (N_17371,N_14594,N_10618);
nand U17372 (N_17372,N_11991,N_10917);
nor U17373 (N_17373,N_10034,N_12087);
and U17374 (N_17374,N_13981,N_10860);
xor U17375 (N_17375,N_10987,N_10064);
or U17376 (N_17376,N_10712,N_13481);
xnor U17377 (N_17377,N_12781,N_12480);
nand U17378 (N_17378,N_13248,N_13505);
and U17379 (N_17379,N_10427,N_11809);
nor U17380 (N_17380,N_10596,N_11302);
nand U17381 (N_17381,N_11786,N_10403);
nor U17382 (N_17382,N_12554,N_11848);
nor U17383 (N_17383,N_13059,N_11812);
nor U17384 (N_17384,N_10461,N_14649);
nor U17385 (N_17385,N_12418,N_10413);
or U17386 (N_17386,N_11961,N_11675);
nand U17387 (N_17387,N_13919,N_11949);
nand U17388 (N_17388,N_13402,N_13111);
and U17389 (N_17389,N_13799,N_12782);
and U17390 (N_17390,N_11960,N_14012);
xor U17391 (N_17391,N_10346,N_14027);
and U17392 (N_17392,N_14811,N_12620);
xnor U17393 (N_17393,N_14931,N_12239);
nand U17394 (N_17394,N_11665,N_13447);
nor U17395 (N_17395,N_14183,N_14789);
nor U17396 (N_17396,N_13400,N_10338);
nand U17397 (N_17397,N_10609,N_14854);
xor U17398 (N_17398,N_12770,N_11568);
nand U17399 (N_17399,N_11937,N_11633);
xnor U17400 (N_17400,N_12307,N_13339);
nand U17401 (N_17401,N_11818,N_13476);
nand U17402 (N_17402,N_11195,N_14415);
xnor U17403 (N_17403,N_12148,N_10696);
and U17404 (N_17404,N_13359,N_10862);
or U17405 (N_17405,N_13498,N_12619);
and U17406 (N_17406,N_10718,N_10942);
nand U17407 (N_17407,N_10092,N_13077);
and U17408 (N_17408,N_12751,N_13973);
xor U17409 (N_17409,N_12281,N_14511);
nand U17410 (N_17410,N_11887,N_13897);
and U17411 (N_17411,N_10570,N_12575);
nor U17412 (N_17412,N_13867,N_11243);
nor U17413 (N_17413,N_10314,N_13997);
and U17414 (N_17414,N_13267,N_13299);
nand U17415 (N_17415,N_10274,N_12350);
nand U17416 (N_17416,N_11621,N_14530);
nor U17417 (N_17417,N_10308,N_13351);
nor U17418 (N_17418,N_14198,N_10834);
nor U17419 (N_17419,N_11694,N_13262);
xor U17420 (N_17420,N_13058,N_14445);
xor U17421 (N_17421,N_10804,N_11415);
xnor U17422 (N_17422,N_13226,N_10252);
nor U17423 (N_17423,N_10071,N_10496);
or U17424 (N_17424,N_10216,N_10565);
nand U17425 (N_17425,N_12306,N_13923);
nor U17426 (N_17426,N_13859,N_13600);
xor U17427 (N_17427,N_11294,N_10217);
xor U17428 (N_17428,N_10965,N_13707);
or U17429 (N_17429,N_14421,N_14604);
nor U17430 (N_17430,N_14116,N_11165);
nor U17431 (N_17431,N_11829,N_11348);
or U17432 (N_17432,N_10121,N_14122);
nor U17433 (N_17433,N_14010,N_11600);
and U17434 (N_17434,N_11154,N_10105);
or U17435 (N_17435,N_10697,N_11543);
nand U17436 (N_17436,N_13464,N_11541);
nand U17437 (N_17437,N_12114,N_14539);
and U17438 (N_17438,N_14595,N_14208);
xnor U17439 (N_17439,N_11238,N_11430);
nand U17440 (N_17440,N_10018,N_10289);
and U17441 (N_17441,N_10286,N_10532);
or U17442 (N_17442,N_11379,N_12515);
nand U17443 (N_17443,N_13594,N_11332);
nand U17444 (N_17444,N_11156,N_11606);
and U17445 (N_17445,N_10556,N_13556);
and U17446 (N_17446,N_12341,N_11806);
and U17447 (N_17447,N_11274,N_12656);
nor U17448 (N_17448,N_14296,N_11278);
xor U17449 (N_17449,N_13074,N_14311);
and U17450 (N_17450,N_14271,N_11117);
nor U17451 (N_17451,N_10894,N_13980);
and U17452 (N_17452,N_13889,N_11985);
and U17453 (N_17453,N_14827,N_13148);
nor U17454 (N_17454,N_10848,N_12519);
or U17455 (N_17455,N_11175,N_12191);
and U17456 (N_17456,N_11418,N_12720);
or U17457 (N_17457,N_12276,N_11842);
or U17458 (N_17458,N_11408,N_12137);
and U17459 (N_17459,N_11716,N_12461);
nor U17460 (N_17460,N_11597,N_14498);
nor U17461 (N_17461,N_10744,N_10790);
or U17462 (N_17462,N_10512,N_12968);
nand U17463 (N_17463,N_10982,N_13123);
xor U17464 (N_17464,N_14910,N_14724);
xnor U17465 (N_17465,N_12339,N_13269);
nand U17466 (N_17466,N_12270,N_10243);
nor U17467 (N_17467,N_13716,N_12540);
nor U17468 (N_17468,N_14203,N_10857);
nor U17469 (N_17469,N_10938,N_13428);
or U17470 (N_17470,N_14013,N_14805);
and U17471 (N_17471,N_14658,N_12466);
or U17472 (N_17472,N_14988,N_10441);
or U17473 (N_17473,N_14186,N_12804);
xnor U17474 (N_17474,N_13547,N_14337);
nand U17475 (N_17475,N_11553,N_11064);
nand U17476 (N_17476,N_13821,N_12346);
xor U17477 (N_17477,N_12794,N_13341);
xnor U17478 (N_17478,N_11454,N_12443);
and U17479 (N_17479,N_14839,N_14609);
and U17480 (N_17480,N_13237,N_11271);
xor U17481 (N_17481,N_11312,N_13479);
nor U17482 (N_17482,N_13563,N_14744);
and U17483 (N_17483,N_14178,N_10303);
and U17484 (N_17484,N_10660,N_14209);
nand U17485 (N_17485,N_12235,N_12489);
or U17486 (N_17486,N_12772,N_10056);
or U17487 (N_17487,N_12837,N_12843);
or U17488 (N_17488,N_12289,N_12262);
and U17489 (N_17489,N_13067,N_12928);
and U17490 (N_17490,N_12808,N_13306);
nor U17491 (N_17491,N_11115,N_12381);
nor U17492 (N_17492,N_13201,N_10928);
nor U17493 (N_17493,N_14155,N_14568);
and U17494 (N_17494,N_13282,N_13743);
and U17495 (N_17495,N_12048,N_13195);
xnor U17496 (N_17496,N_12642,N_12967);
nor U17497 (N_17497,N_12775,N_11232);
or U17498 (N_17498,N_14106,N_10997);
or U17499 (N_17499,N_11197,N_13193);
nor U17500 (N_17500,N_11529,N_13484);
xor U17501 (N_17501,N_10280,N_14726);
or U17502 (N_17502,N_14670,N_11313);
nor U17503 (N_17503,N_13615,N_13744);
xor U17504 (N_17504,N_14806,N_13529);
nand U17505 (N_17505,N_10265,N_12153);
nor U17506 (N_17506,N_11017,N_13306);
and U17507 (N_17507,N_14828,N_10479);
nor U17508 (N_17508,N_12750,N_11609);
and U17509 (N_17509,N_13978,N_12695);
nor U17510 (N_17510,N_14668,N_14427);
nand U17511 (N_17511,N_11536,N_14269);
nor U17512 (N_17512,N_13146,N_12833);
or U17513 (N_17513,N_12059,N_10937);
or U17514 (N_17514,N_12914,N_12566);
xnor U17515 (N_17515,N_11817,N_10410);
and U17516 (N_17516,N_12883,N_14286);
or U17517 (N_17517,N_11296,N_11462);
or U17518 (N_17518,N_11089,N_12489);
or U17519 (N_17519,N_11026,N_13269);
nor U17520 (N_17520,N_11012,N_14324);
and U17521 (N_17521,N_12371,N_13360);
nand U17522 (N_17522,N_13589,N_12276);
xnor U17523 (N_17523,N_10397,N_14061);
or U17524 (N_17524,N_14400,N_12724);
nor U17525 (N_17525,N_10118,N_12513);
nor U17526 (N_17526,N_11215,N_10425);
or U17527 (N_17527,N_11571,N_12036);
or U17528 (N_17528,N_11519,N_12730);
nand U17529 (N_17529,N_11868,N_14630);
or U17530 (N_17530,N_12003,N_11047);
xnor U17531 (N_17531,N_13013,N_12613);
nor U17532 (N_17532,N_13197,N_12464);
nor U17533 (N_17533,N_10744,N_14085);
nand U17534 (N_17534,N_12996,N_10570);
or U17535 (N_17535,N_10664,N_11131);
nand U17536 (N_17536,N_12519,N_14330);
or U17537 (N_17537,N_14400,N_14980);
or U17538 (N_17538,N_13952,N_10575);
xnor U17539 (N_17539,N_11571,N_13339);
or U17540 (N_17540,N_11491,N_12181);
and U17541 (N_17541,N_10678,N_11755);
and U17542 (N_17542,N_12645,N_12907);
xor U17543 (N_17543,N_13968,N_13328);
or U17544 (N_17544,N_13699,N_13302);
or U17545 (N_17545,N_13789,N_13674);
or U17546 (N_17546,N_12807,N_14976);
nand U17547 (N_17547,N_12711,N_13047);
or U17548 (N_17548,N_13255,N_13099);
nor U17549 (N_17549,N_12146,N_14563);
or U17550 (N_17550,N_13420,N_11439);
and U17551 (N_17551,N_13190,N_12452);
or U17552 (N_17552,N_13534,N_13016);
xor U17553 (N_17553,N_13814,N_10855);
xnor U17554 (N_17554,N_13204,N_11867);
and U17555 (N_17555,N_14076,N_11949);
and U17556 (N_17556,N_11394,N_12851);
xor U17557 (N_17557,N_14281,N_14252);
nand U17558 (N_17558,N_10704,N_14816);
and U17559 (N_17559,N_12429,N_12785);
nor U17560 (N_17560,N_14057,N_11193);
nor U17561 (N_17561,N_12606,N_10699);
or U17562 (N_17562,N_14857,N_14664);
or U17563 (N_17563,N_14821,N_14191);
xor U17564 (N_17564,N_12669,N_14936);
or U17565 (N_17565,N_12872,N_11767);
xnor U17566 (N_17566,N_12884,N_12349);
xor U17567 (N_17567,N_12357,N_12521);
or U17568 (N_17568,N_12786,N_12938);
or U17569 (N_17569,N_14507,N_10334);
or U17570 (N_17570,N_14883,N_10609);
nor U17571 (N_17571,N_10235,N_11978);
nand U17572 (N_17572,N_13897,N_11463);
nand U17573 (N_17573,N_13087,N_11763);
nor U17574 (N_17574,N_13869,N_13403);
xor U17575 (N_17575,N_12029,N_12166);
or U17576 (N_17576,N_14737,N_13196);
xor U17577 (N_17577,N_10961,N_14713);
and U17578 (N_17578,N_14452,N_13287);
nand U17579 (N_17579,N_14343,N_11360);
and U17580 (N_17580,N_14408,N_13544);
nand U17581 (N_17581,N_13738,N_12268);
nand U17582 (N_17582,N_14283,N_14222);
or U17583 (N_17583,N_11478,N_10027);
xnor U17584 (N_17584,N_13718,N_14997);
nor U17585 (N_17585,N_12220,N_12954);
and U17586 (N_17586,N_10171,N_12868);
or U17587 (N_17587,N_10904,N_12399);
nand U17588 (N_17588,N_13522,N_10086);
and U17589 (N_17589,N_12704,N_11865);
xnor U17590 (N_17590,N_14344,N_13599);
nand U17591 (N_17591,N_14795,N_12754);
or U17592 (N_17592,N_10265,N_10974);
or U17593 (N_17593,N_13592,N_12116);
nor U17594 (N_17594,N_14716,N_10432);
or U17595 (N_17595,N_14249,N_13604);
nor U17596 (N_17596,N_10998,N_13833);
xor U17597 (N_17597,N_10900,N_14515);
nor U17598 (N_17598,N_10033,N_14196);
and U17599 (N_17599,N_10104,N_10286);
nand U17600 (N_17600,N_10155,N_10766);
or U17601 (N_17601,N_10614,N_13554);
xnor U17602 (N_17602,N_13400,N_12924);
or U17603 (N_17603,N_12616,N_12285);
or U17604 (N_17604,N_10933,N_14600);
or U17605 (N_17605,N_10595,N_11922);
and U17606 (N_17606,N_14003,N_10075);
or U17607 (N_17607,N_14568,N_10420);
and U17608 (N_17608,N_12425,N_12237);
or U17609 (N_17609,N_10179,N_12883);
xnor U17610 (N_17610,N_11190,N_14001);
nand U17611 (N_17611,N_11968,N_12334);
xor U17612 (N_17612,N_12891,N_13769);
nand U17613 (N_17613,N_10957,N_10460);
nor U17614 (N_17614,N_13013,N_12618);
nand U17615 (N_17615,N_14014,N_11252);
nor U17616 (N_17616,N_10074,N_11089);
nand U17617 (N_17617,N_11820,N_13519);
and U17618 (N_17618,N_14879,N_10537);
xor U17619 (N_17619,N_13461,N_12752);
or U17620 (N_17620,N_13652,N_11863);
nor U17621 (N_17621,N_11396,N_14521);
nand U17622 (N_17622,N_13183,N_10207);
xor U17623 (N_17623,N_11074,N_10143);
and U17624 (N_17624,N_11856,N_14851);
nor U17625 (N_17625,N_11389,N_13185);
and U17626 (N_17626,N_11883,N_13179);
nor U17627 (N_17627,N_13518,N_14925);
nor U17628 (N_17628,N_12030,N_13892);
and U17629 (N_17629,N_11497,N_10432);
xnor U17630 (N_17630,N_12935,N_11829);
nand U17631 (N_17631,N_11645,N_13787);
xor U17632 (N_17632,N_12808,N_10700);
or U17633 (N_17633,N_11254,N_11482);
nor U17634 (N_17634,N_11544,N_11243);
or U17635 (N_17635,N_14029,N_11437);
or U17636 (N_17636,N_14670,N_10173);
nor U17637 (N_17637,N_12657,N_11289);
or U17638 (N_17638,N_12351,N_10960);
nor U17639 (N_17639,N_12809,N_13388);
or U17640 (N_17640,N_13991,N_10799);
or U17641 (N_17641,N_12685,N_14869);
and U17642 (N_17642,N_11865,N_12665);
nor U17643 (N_17643,N_11120,N_12891);
and U17644 (N_17644,N_10811,N_10943);
or U17645 (N_17645,N_14050,N_14947);
or U17646 (N_17646,N_10740,N_14796);
xor U17647 (N_17647,N_11012,N_14845);
xor U17648 (N_17648,N_12765,N_14842);
xor U17649 (N_17649,N_13006,N_10560);
or U17650 (N_17650,N_13325,N_12080);
xnor U17651 (N_17651,N_11587,N_11139);
nand U17652 (N_17652,N_12136,N_14560);
or U17653 (N_17653,N_11369,N_11480);
nand U17654 (N_17654,N_14629,N_14221);
nand U17655 (N_17655,N_13529,N_11105);
or U17656 (N_17656,N_11946,N_12919);
nand U17657 (N_17657,N_12337,N_13386);
xnor U17658 (N_17658,N_12180,N_14558);
or U17659 (N_17659,N_10566,N_10841);
and U17660 (N_17660,N_12576,N_13759);
or U17661 (N_17661,N_10114,N_10189);
nand U17662 (N_17662,N_14901,N_14295);
nand U17663 (N_17663,N_14490,N_11574);
nor U17664 (N_17664,N_13162,N_12962);
nand U17665 (N_17665,N_11240,N_12320);
nor U17666 (N_17666,N_12116,N_10640);
nand U17667 (N_17667,N_14901,N_11964);
xor U17668 (N_17668,N_11515,N_13044);
nand U17669 (N_17669,N_10457,N_14291);
nand U17670 (N_17670,N_14395,N_14384);
or U17671 (N_17671,N_14779,N_10570);
xor U17672 (N_17672,N_10582,N_10993);
or U17673 (N_17673,N_12049,N_14768);
nor U17674 (N_17674,N_10495,N_10687);
or U17675 (N_17675,N_14580,N_14923);
xnor U17676 (N_17676,N_14162,N_13245);
nand U17677 (N_17677,N_11267,N_14251);
xor U17678 (N_17678,N_13258,N_13828);
xnor U17679 (N_17679,N_12967,N_11894);
nand U17680 (N_17680,N_11742,N_14448);
and U17681 (N_17681,N_14689,N_14052);
nor U17682 (N_17682,N_12607,N_13841);
or U17683 (N_17683,N_11074,N_10691);
nor U17684 (N_17684,N_13094,N_10561);
nand U17685 (N_17685,N_13492,N_12863);
nand U17686 (N_17686,N_13970,N_14651);
nand U17687 (N_17687,N_14461,N_12605);
nor U17688 (N_17688,N_10429,N_10638);
or U17689 (N_17689,N_13049,N_14560);
nand U17690 (N_17690,N_10382,N_13844);
or U17691 (N_17691,N_11618,N_11682);
xor U17692 (N_17692,N_14605,N_13755);
or U17693 (N_17693,N_12856,N_10629);
xor U17694 (N_17694,N_13597,N_13135);
and U17695 (N_17695,N_10196,N_12112);
and U17696 (N_17696,N_10598,N_10074);
xor U17697 (N_17697,N_14494,N_13569);
or U17698 (N_17698,N_14045,N_13909);
nand U17699 (N_17699,N_13607,N_13828);
and U17700 (N_17700,N_13964,N_12093);
nand U17701 (N_17701,N_14953,N_13797);
xnor U17702 (N_17702,N_10190,N_11824);
nor U17703 (N_17703,N_12104,N_13350);
and U17704 (N_17704,N_11340,N_10367);
and U17705 (N_17705,N_11300,N_10724);
nor U17706 (N_17706,N_14512,N_13634);
nor U17707 (N_17707,N_14681,N_12212);
or U17708 (N_17708,N_12732,N_14595);
xnor U17709 (N_17709,N_10966,N_12187);
and U17710 (N_17710,N_14031,N_10574);
or U17711 (N_17711,N_12023,N_13567);
or U17712 (N_17712,N_13107,N_12652);
or U17713 (N_17713,N_10319,N_14889);
nor U17714 (N_17714,N_13848,N_12804);
xnor U17715 (N_17715,N_11576,N_13796);
nor U17716 (N_17716,N_10814,N_12908);
nand U17717 (N_17717,N_14236,N_13085);
xor U17718 (N_17718,N_11515,N_14171);
or U17719 (N_17719,N_10408,N_11912);
or U17720 (N_17720,N_12213,N_10793);
nor U17721 (N_17721,N_12911,N_10517);
or U17722 (N_17722,N_13994,N_12245);
and U17723 (N_17723,N_14136,N_12631);
or U17724 (N_17724,N_10985,N_13632);
nand U17725 (N_17725,N_11500,N_11373);
xor U17726 (N_17726,N_14581,N_12525);
and U17727 (N_17727,N_13994,N_10036);
and U17728 (N_17728,N_13535,N_14442);
nor U17729 (N_17729,N_11541,N_11281);
or U17730 (N_17730,N_13082,N_14521);
nand U17731 (N_17731,N_11995,N_13839);
and U17732 (N_17732,N_12071,N_14924);
nand U17733 (N_17733,N_12401,N_12032);
nand U17734 (N_17734,N_14810,N_10026);
nor U17735 (N_17735,N_14512,N_10344);
nand U17736 (N_17736,N_10898,N_13832);
xor U17737 (N_17737,N_12296,N_13825);
nor U17738 (N_17738,N_12237,N_13140);
nor U17739 (N_17739,N_13317,N_11257);
nand U17740 (N_17740,N_12672,N_11233);
and U17741 (N_17741,N_14788,N_11957);
or U17742 (N_17742,N_13455,N_14709);
and U17743 (N_17743,N_10284,N_11774);
or U17744 (N_17744,N_11530,N_12623);
xnor U17745 (N_17745,N_11083,N_12828);
or U17746 (N_17746,N_10700,N_10582);
xor U17747 (N_17747,N_11509,N_12492);
and U17748 (N_17748,N_14900,N_12416);
nand U17749 (N_17749,N_11684,N_13829);
or U17750 (N_17750,N_13375,N_12705);
or U17751 (N_17751,N_12299,N_10646);
nor U17752 (N_17752,N_10225,N_13221);
nor U17753 (N_17753,N_12459,N_14608);
nor U17754 (N_17754,N_14343,N_11686);
or U17755 (N_17755,N_11833,N_10318);
or U17756 (N_17756,N_12315,N_13933);
nand U17757 (N_17757,N_11981,N_13851);
and U17758 (N_17758,N_14577,N_12565);
nand U17759 (N_17759,N_13175,N_14467);
nand U17760 (N_17760,N_12097,N_10771);
or U17761 (N_17761,N_13957,N_13264);
nor U17762 (N_17762,N_12700,N_14189);
or U17763 (N_17763,N_14246,N_11741);
xnor U17764 (N_17764,N_11650,N_10464);
xor U17765 (N_17765,N_11618,N_10435);
nor U17766 (N_17766,N_12708,N_12933);
nand U17767 (N_17767,N_10315,N_12760);
and U17768 (N_17768,N_11154,N_11308);
xnor U17769 (N_17769,N_13393,N_10423);
and U17770 (N_17770,N_11468,N_10447);
and U17771 (N_17771,N_11405,N_12529);
and U17772 (N_17772,N_14887,N_12589);
and U17773 (N_17773,N_10756,N_10196);
and U17774 (N_17774,N_10411,N_11189);
and U17775 (N_17775,N_13165,N_11916);
or U17776 (N_17776,N_10984,N_12312);
or U17777 (N_17777,N_11674,N_12196);
nor U17778 (N_17778,N_13229,N_14585);
and U17779 (N_17779,N_12822,N_14057);
nand U17780 (N_17780,N_13930,N_13417);
and U17781 (N_17781,N_12814,N_12516);
nor U17782 (N_17782,N_12530,N_12894);
xor U17783 (N_17783,N_10924,N_14674);
and U17784 (N_17784,N_10252,N_14458);
nor U17785 (N_17785,N_11625,N_10273);
xor U17786 (N_17786,N_11441,N_12703);
xnor U17787 (N_17787,N_12507,N_11889);
and U17788 (N_17788,N_14989,N_11388);
and U17789 (N_17789,N_11047,N_13116);
xnor U17790 (N_17790,N_10978,N_14190);
xnor U17791 (N_17791,N_12561,N_12224);
and U17792 (N_17792,N_10068,N_12399);
nor U17793 (N_17793,N_11883,N_12629);
and U17794 (N_17794,N_10032,N_13273);
or U17795 (N_17795,N_14100,N_13707);
xor U17796 (N_17796,N_14086,N_12915);
and U17797 (N_17797,N_10156,N_10945);
nor U17798 (N_17798,N_11150,N_14408);
or U17799 (N_17799,N_14490,N_13697);
xor U17800 (N_17800,N_14734,N_11203);
nor U17801 (N_17801,N_14067,N_12592);
xor U17802 (N_17802,N_13752,N_14790);
nor U17803 (N_17803,N_13039,N_10552);
xnor U17804 (N_17804,N_14529,N_10637);
or U17805 (N_17805,N_14024,N_13699);
and U17806 (N_17806,N_12813,N_10572);
or U17807 (N_17807,N_14473,N_14228);
xor U17808 (N_17808,N_14177,N_10656);
xor U17809 (N_17809,N_10131,N_13461);
xor U17810 (N_17810,N_14947,N_10606);
nor U17811 (N_17811,N_13555,N_13352);
nor U17812 (N_17812,N_14422,N_12085);
nor U17813 (N_17813,N_11317,N_12589);
nor U17814 (N_17814,N_14596,N_10526);
and U17815 (N_17815,N_14194,N_10059);
and U17816 (N_17816,N_13814,N_13076);
nand U17817 (N_17817,N_10633,N_11593);
nor U17818 (N_17818,N_13243,N_11754);
and U17819 (N_17819,N_11724,N_10587);
xnor U17820 (N_17820,N_13964,N_13765);
and U17821 (N_17821,N_12799,N_10782);
and U17822 (N_17822,N_12065,N_14643);
and U17823 (N_17823,N_14565,N_13848);
nand U17824 (N_17824,N_10407,N_10299);
nor U17825 (N_17825,N_13827,N_10438);
nand U17826 (N_17826,N_13157,N_11903);
or U17827 (N_17827,N_11333,N_14736);
nand U17828 (N_17828,N_13646,N_11908);
or U17829 (N_17829,N_14344,N_11576);
nand U17830 (N_17830,N_14421,N_13216);
and U17831 (N_17831,N_10038,N_11516);
and U17832 (N_17832,N_12664,N_14093);
nand U17833 (N_17833,N_11091,N_10674);
nor U17834 (N_17834,N_10191,N_11290);
xor U17835 (N_17835,N_14898,N_11249);
and U17836 (N_17836,N_14703,N_14645);
or U17837 (N_17837,N_11443,N_14424);
nor U17838 (N_17838,N_12646,N_10219);
and U17839 (N_17839,N_12966,N_12392);
or U17840 (N_17840,N_11573,N_10426);
or U17841 (N_17841,N_14825,N_11458);
nand U17842 (N_17842,N_13586,N_12995);
xor U17843 (N_17843,N_14018,N_10949);
nand U17844 (N_17844,N_14632,N_12940);
nor U17845 (N_17845,N_12004,N_12253);
xor U17846 (N_17846,N_12028,N_14706);
or U17847 (N_17847,N_13563,N_14102);
or U17848 (N_17848,N_10636,N_14944);
nand U17849 (N_17849,N_10900,N_10037);
and U17850 (N_17850,N_13074,N_11831);
and U17851 (N_17851,N_13711,N_14338);
xnor U17852 (N_17852,N_14701,N_10614);
nand U17853 (N_17853,N_11844,N_14647);
and U17854 (N_17854,N_12038,N_12945);
xnor U17855 (N_17855,N_12033,N_12850);
nand U17856 (N_17856,N_14668,N_14986);
or U17857 (N_17857,N_13454,N_13670);
and U17858 (N_17858,N_12311,N_13982);
nor U17859 (N_17859,N_11187,N_13572);
xnor U17860 (N_17860,N_14326,N_14662);
nor U17861 (N_17861,N_12694,N_12455);
nand U17862 (N_17862,N_10519,N_14359);
and U17863 (N_17863,N_10832,N_11738);
xnor U17864 (N_17864,N_12779,N_10327);
nor U17865 (N_17865,N_13087,N_11978);
and U17866 (N_17866,N_14781,N_11933);
nand U17867 (N_17867,N_13367,N_10026);
and U17868 (N_17868,N_11566,N_14082);
and U17869 (N_17869,N_10037,N_11283);
nand U17870 (N_17870,N_11449,N_10753);
nor U17871 (N_17871,N_13255,N_13681);
nor U17872 (N_17872,N_11980,N_11492);
nor U17873 (N_17873,N_10428,N_12934);
nor U17874 (N_17874,N_12784,N_14419);
xor U17875 (N_17875,N_11986,N_14164);
or U17876 (N_17876,N_11926,N_10338);
and U17877 (N_17877,N_10986,N_11143);
nand U17878 (N_17878,N_14486,N_12860);
nand U17879 (N_17879,N_10787,N_14174);
nand U17880 (N_17880,N_12208,N_14732);
and U17881 (N_17881,N_14948,N_11293);
xnor U17882 (N_17882,N_14417,N_12427);
xnor U17883 (N_17883,N_10751,N_14554);
or U17884 (N_17884,N_12425,N_13797);
nor U17885 (N_17885,N_13645,N_14965);
nand U17886 (N_17886,N_13118,N_11931);
xnor U17887 (N_17887,N_14020,N_10827);
nand U17888 (N_17888,N_10265,N_11176);
or U17889 (N_17889,N_10148,N_12673);
and U17890 (N_17890,N_14479,N_14231);
and U17891 (N_17891,N_11031,N_14679);
xnor U17892 (N_17892,N_10167,N_13843);
xor U17893 (N_17893,N_11342,N_10322);
nand U17894 (N_17894,N_12095,N_13428);
xnor U17895 (N_17895,N_11888,N_12659);
or U17896 (N_17896,N_10269,N_13388);
nor U17897 (N_17897,N_10086,N_10818);
and U17898 (N_17898,N_14700,N_12440);
nor U17899 (N_17899,N_11163,N_12239);
and U17900 (N_17900,N_14070,N_14657);
xor U17901 (N_17901,N_11929,N_14729);
xor U17902 (N_17902,N_13432,N_13558);
and U17903 (N_17903,N_14279,N_13837);
nand U17904 (N_17904,N_10490,N_11090);
xor U17905 (N_17905,N_14489,N_10890);
nand U17906 (N_17906,N_14120,N_14475);
and U17907 (N_17907,N_11493,N_13150);
and U17908 (N_17908,N_14125,N_14241);
xnor U17909 (N_17909,N_14198,N_14217);
nor U17910 (N_17910,N_10103,N_12143);
nand U17911 (N_17911,N_10129,N_14709);
nor U17912 (N_17912,N_14286,N_14300);
xnor U17913 (N_17913,N_12085,N_10636);
xnor U17914 (N_17914,N_10553,N_13024);
nand U17915 (N_17915,N_11006,N_12244);
nor U17916 (N_17916,N_11169,N_14956);
or U17917 (N_17917,N_11365,N_13717);
or U17918 (N_17918,N_12114,N_11763);
and U17919 (N_17919,N_14244,N_12112);
xnor U17920 (N_17920,N_13986,N_14989);
and U17921 (N_17921,N_14830,N_13261);
nand U17922 (N_17922,N_11412,N_10024);
nor U17923 (N_17923,N_14290,N_14305);
and U17924 (N_17924,N_14295,N_10233);
and U17925 (N_17925,N_12335,N_10344);
nor U17926 (N_17926,N_14990,N_12686);
and U17927 (N_17927,N_12398,N_11890);
nor U17928 (N_17928,N_14663,N_11850);
or U17929 (N_17929,N_14388,N_10207);
and U17930 (N_17930,N_12623,N_11870);
nand U17931 (N_17931,N_12798,N_14379);
nand U17932 (N_17932,N_13484,N_14730);
or U17933 (N_17933,N_11155,N_13362);
nor U17934 (N_17934,N_10785,N_14539);
and U17935 (N_17935,N_12695,N_11082);
and U17936 (N_17936,N_10619,N_11024);
or U17937 (N_17937,N_10356,N_10119);
or U17938 (N_17938,N_11334,N_13215);
nor U17939 (N_17939,N_13805,N_14918);
xor U17940 (N_17940,N_10845,N_12009);
or U17941 (N_17941,N_12619,N_11294);
and U17942 (N_17942,N_14149,N_12885);
nand U17943 (N_17943,N_13694,N_10197);
nor U17944 (N_17944,N_11967,N_13631);
or U17945 (N_17945,N_11041,N_12275);
nand U17946 (N_17946,N_12425,N_13661);
nand U17947 (N_17947,N_10703,N_12602);
and U17948 (N_17948,N_10096,N_12913);
or U17949 (N_17949,N_11427,N_10434);
and U17950 (N_17950,N_10358,N_14786);
or U17951 (N_17951,N_12823,N_10572);
nor U17952 (N_17952,N_13522,N_12440);
and U17953 (N_17953,N_12235,N_10076);
nor U17954 (N_17954,N_14544,N_10387);
xnor U17955 (N_17955,N_10610,N_12276);
nor U17956 (N_17956,N_13942,N_11160);
nor U17957 (N_17957,N_12322,N_11500);
and U17958 (N_17958,N_10477,N_14958);
nand U17959 (N_17959,N_14107,N_10556);
nand U17960 (N_17960,N_12546,N_10615);
nand U17961 (N_17961,N_14886,N_12612);
and U17962 (N_17962,N_11370,N_12720);
and U17963 (N_17963,N_13084,N_10214);
nor U17964 (N_17964,N_11175,N_13826);
xor U17965 (N_17965,N_14479,N_10866);
nand U17966 (N_17966,N_10467,N_13264);
nand U17967 (N_17967,N_11889,N_14240);
nand U17968 (N_17968,N_12884,N_10629);
nor U17969 (N_17969,N_14256,N_12341);
nand U17970 (N_17970,N_13957,N_10176);
nand U17971 (N_17971,N_11031,N_14221);
and U17972 (N_17972,N_14575,N_12742);
nor U17973 (N_17973,N_13371,N_13269);
nor U17974 (N_17974,N_11070,N_10939);
and U17975 (N_17975,N_13940,N_13061);
and U17976 (N_17976,N_11304,N_13621);
nor U17977 (N_17977,N_10743,N_13218);
or U17978 (N_17978,N_11206,N_11421);
and U17979 (N_17979,N_11760,N_12750);
nand U17980 (N_17980,N_14190,N_12558);
nor U17981 (N_17981,N_10118,N_11936);
nand U17982 (N_17982,N_14339,N_12901);
nor U17983 (N_17983,N_11388,N_11898);
nor U17984 (N_17984,N_11771,N_11098);
nor U17985 (N_17985,N_12063,N_11336);
xnor U17986 (N_17986,N_13228,N_11849);
nor U17987 (N_17987,N_12209,N_14421);
nand U17988 (N_17988,N_14444,N_13570);
or U17989 (N_17989,N_10666,N_14936);
or U17990 (N_17990,N_12408,N_13803);
and U17991 (N_17991,N_12742,N_12865);
nor U17992 (N_17992,N_14948,N_12699);
nor U17993 (N_17993,N_14108,N_12051);
xnor U17994 (N_17994,N_11780,N_10581);
xnor U17995 (N_17995,N_14401,N_11411);
nor U17996 (N_17996,N_11906,N_14061);
xnor U17997 (N_17997,N_13468,N_11692);
nand U17998 (N_17998,N_13995,N_14911);
xnor U17999 (N_17999,N_14817,N_11602);
nor U18000 (N_18000,N_12931,N_12818);
nor U18001 (N_18001,N_10428,N_13563);
or U18002 (N_18002,N_13102,N_14895);
or U18003 (N_18003,N_14295,N_12784);
nor U18004 (N_18004,N_11891,N_10251);
and U18005 (N_18005,N_10661,N_10576);
nor U18006 (N_18006,N_14207,N_12993);
or U18007 (N_18007,N_12642,N_11592);
and U18008 (N_18008,N_12245,N_12916);
xor U18009 (N_18009,N_10129,N_13269);
xnor U18010 (N_18010,N_14841,N_11231);
nor U18011 (N_18011,N_13960,N_13104);
nor U18012 (N_18012,N_13468,N_13842);
xor U18013 (N_18013,N_12074,N_12804);
nor U18014 (N_18014,N_12319,N_11182);
and U18015 (N_18015,N_14300,N_10905);
and U18016 (N_18016,N_10234,N_11589);
and U18017 (N_18017,N_10262,N_10557);
nor U18018 (N_18018,N_10495,N_14034);
nand U18019 (N_18019,N_12834,N_12198);
nor U18020 (N_18020,N_11383,N_13935);
nor U18021 (N_18021,N_12327,N_14833);
or U18022 (N_18022,N_14088,N_14967);
and U18023 (N_18023,N_14372,N_11997);
nor U18024 (N_18024,N_11661,N_13852);
or U18025 (N_18025,N_10127,N_11825);
nand U18026 (N_18026,N_12726,N_13766);
and U18027 (N_18027,N_14370,N_10733);
or U18028 (N_18028,N_14687,N_13574);
or U18029 (N_18029,N_11350,N_13386);
nand U18030 (N_18030,N_10587,N_12620);
or U18031 (N_18031,N_13864,N_12685);
and U18032 (N_18032,N_13149,N_12449);
xor U18033 (N_18033,N_12006,N_10520);
nor U18034 (N_18034,N_12496,N_14696);
nor U18035 (N_18035,N_12514,N_14781);
or U18036 (N_18036,N_13400,N_13681);
xnor U18037 (N_18037,N_10127,N_13205);
nor U18038 (N_18038,N_11995,N_14013);
or U18039 (N_18039,N_14938,N_12945);
xor U18040 (N_18040,N_11144,N_12616);
and U18041 (N_18041,N_13358,N_12585);
xor U18042 (N_18042,N_12907,N_10545);
and U18043 (N_18043,N_10620,N_14041);
nand U18044 (N_18044,N_11493,N_12860);
xor U18045 (N_18045,N_12738,N_10453);
xnor U18046 (N_18046,N_13669,N_14824);
or U18047 (N_18047,N_13500,N_11093);
or U18048 (N_18048,N_14036,N_13387);
nand U18049 (N_18049,N_14960,N_11039);
and U18050 (N_18050,N_11034,N_14717);
nand U18051 (N_18051,N_14623,N_10331);
nor U18052 (N_18052,N_14580,N_14598);
nor U18053 (N_18053,N_14303,N_10018);
xnor U18054 (N_18054,N_12413,N_13392);
or U18055 (N_18055,N_10279,N_13578);
nand U18056 (N_18056,N_11945,N_11124);
and U18057 (N_18057,N_12900,N_10518);
nand U18058 (N_18058,N_13136,N_12171);
or U18059 (N_18059,N_10117,N_11989);
or U18060 (N_18060,N_11900,N_10337);
or U18061 (N_18061,N_11059,N_11656);
xnor U18062 (N_18062,N_10860,N_12046);
nand U18063 (N_18063,N_11555,N_10540);
or U18064 (N_18064,N_10265,N_10505);
xnor U18065 (N_18065,N_11172,N_12996);
or U18066 (N_18066,N_14722,N_10835);
nor U18067 (N_18067,N_11572,N_13100);
and U18068 (N_18068,N_14718,N_13675);
and U18069 (N_18069,N_13724,N_10904);
and U18070 (N_18070,N_14823,N_11973);
or U18071 (N_18071,N_10225,N_10256);
and U18072 (N_18072,N_14246,N_11489);
or U18073 (N_18073,N_11828,N_10265);
xnor U18074 (N_18074,N_13854,N_12494);
and U18075 (N_18075,N_13715,N_12118);
and U18076 (N_18076,N_12185,N_11349);
or U18077 (N_18077,N_14776,N_12505);
and U18078 (N_18078,N_13543,N_14076);
and U18079 (N_18079,N_14647,N_11211);
nand U18080 (N_18080,N_13591,N_10556);
xor U18081 (N_18081,N_10588,N_12647);
xor U18082 (N_18082,N_14937,N_12438);
and U18083 (N_18083,N_14165,N_12607);
and U18084 (N_18084,N_11310,N_10884);
or U18085 (N_18085,N_13263,N_12168);
or U18086 (N_18086,N_10926,N_10828);
or U18087 (N_18087,N_11039,N_10964);
or U18088 (N_18088,N_13799,N_11616);
and U18089 (N_18089,N_11429,N_13246);
xor U18090 (N_18090,N_10558,N_14369);
and U18091 (N_18091,N_13686,N_13892);
and U18092 (N_18092,N_13247,N_14543);
nand U18093 (N_18093,N_14017,N_11120);
xnor U18094 (N_18094,N_11886,N_10482);
nor U18095 (N_18095,N_12958,N_11571);
xor U18096 (N_18096,N_12615,N_14029);
xor U18097 (N_18097,N_10907,N_12135);
xnor U18098 (N_18098,N_11849,N_10803);
nor U18099 (N_18099,N_11441,N_11545);
nand U18100 (N_18100,N_12081,N_12101);
or U18101 (N_18101,N_10772,N_13139);
nand U18102 (N_18102,N_13294,N_12756);
nor U18103 (N_18103,N_11699,N_13200);
and U18104 (N_18104,N_11978,N_10123);
nand U18105 (N_18105,N_10310,N_12859);
or U18106 (N_18106,N_14211,N_13785);
nand U18107 (N_18107,N_14746,N_11480);
xor U18108 (N_18108,N_12018,N_14874);
xor U18109 (N_18109,N_13447,N_13435);
or U18110 (N_18110,N_12545,N_13932);
nand U18111 (N_18111,N_12225,N_13878);
nand U18112 (N_18112,N_11358,N_11461);
nor U18113 (N_18113,N_10852,N_11661);
and U18114 (N_18114,N_12648,N_10679);
nor U18115 (N_18115,N_11003,N_10544);
nor U18116 (N_18116,N_13789,N_11174);
xnor U18117 (N_18117,N_14656,N_14073);
xor U18118 (N_18118,N_13340,N_14283);
nand U18119 (N_18119,N_14541,N_12969);
nor U18120 (N_18120,N_13850,N_10100);
xnor U18121 (N_18121,N_12289,N_11324);
nand U18122 (N_18122,N_10967,N_13362);
xnor U18123 (N_18123,N_10237,N_13361);
xnor U18124 (N_18124,N_10942,N_12240);
and U18125 (N_18125,N_12942,N_12632);
nand U18126 (N_18126,N_10906,N_10056);
xnor U18127 (N_18127,N_12261,N_14089);
or U18128 (N_18128,N_14174,N_13183);
nand U18129 (N_18129,N_13405,N_10945);
xor U18130 (N_18130,N_14135,N_13252);
xnor U18131 (N_18131,N_11441,N_13644);
xor U18132 (N_18132,N_13550,N_12105);
nand U18133 (N_18133,N_11776,N_13152);
nand U18134 (N_18134,N_14829,N_10646);
nand U18135 (N_18135,N_10673,N_14228);
nand U18136 (N_18136,N_12187,N_14894);
or U18137 (N_18137,N_10776,N_10315);
nor U18138 (N_18138,N_11647,N_14349);
and U18139 (N_18139,N_14794,N_14930);
and U18140 (N_18140,N_11417,N_13941);
and U18141 (N_18141,N_14998,N_14786);
xor U18142 (N_18142,N_12044,N_10048);
or U18143 (N_18143,N_10141,N_14787);
nor U18144 (N_18144,N_12065,N_11236);
nand U18145 (N_18145,N_11537,N_11365);
nor U18146 (N_18146,N_10063,N_10439);
and U18147 (N_18147,N_13670,N_12728);
nand U18148 (N_18148,N_12602,N_12865);
nor U18149 (N_18149,N_14425,N_14866);
xor U18150 (N_18150,N_11287,N_10651);
or U18151 (N_18151,N_11756,N_14468);
and U18152 (N_18152,N_11499,N_12454);
xnor U18153 (N_18153,N_12370,N_11115);
nand U18154 (N_18154,N_14573,N_14467);
or U18155 (N_18155,N_14724,N_14827);
xnor U18156 (N_18156,N_11648,N_14446);
nand U18157 (N_18157,N_11637,N_12892);
nand U18158 (N_18158,N_13793,N_14257);
nand U18159 (N_18159,N_13160,N_10873);
xnor U18160 (N_18160,N_11114,N_12121);
nor U18161 (N_18161,N_13133,N_13403);
nor U18162 (N_18162,N_10057,N_10166);
or U18163 (N_18163,N_11613,N_13688);
and U18164 (N_18164,N_14512,N_10597);
nand U18165 (N_18165,N_12111,N_10248);
xnor U18166 (N_18166,N_13395,N_13289);
xor U18167 (N_18167,N_10202,N_14385);
or U18168 (N_18168,N_11206,N_13633);
or U18169 (N_18169,N_14232,N_13164);
xor U18170 (N_18170,N_13489,N_13363);
and U18171 (N_18171,N_10528,N_12031);
and U18172 (N_18172,N_13613,N_11402);
nor U18173 (N_18173,N_14315,N_12463);
nor U18174 (N_18174,N_11192,N_12148);
nand U18175 (N_18175,N_10102,N_10693);
nor U18176 (N_18176,N_10904,N_14122);
and U18177 (N_18177,N_12620,N_14736);
xor U18178 (N_18178,N_10489,N_14507);
or U18179 (N_18179,N_11032,N_13586);
nand U18180 (N_18180,N_10334,N_14814);
and U18181 (N_18181,N_11250,N_14495);
xor U18182 (N_18182,N_13372,N_12578);
nor U18183 (N_18183,N_14433,N_12172);
nor U18184 (N_18184,N_12276,N_11331);
nor U18185 (N_18185,N_10632,N_13354);
or U18186 (N_18186,N_10793,N_12515);
nor U18187 (N_18187,N_12641,N_11689);
xor U18188 (N_18188,N_14628,N_14961);
nand U18189 (N_18189,N_10768,N_13039);
or U18190 (N_18190,N_13817,N_10128);
nand U18191 (N_18191,N_11459,N_13159);
nand U18192 (N_18192,N_13135,N_13357);
xnor U18193 (N_18193,N_10976,N_13806);
or U18194 (N_18194,N_12221,N_13018);
nor U18195 (N_18195,N_14260,N_13203);
and U18196 (N_18196,N_13629,N_10791);
or U18197 (N_18197,N_13489,N_14986);
or U18198 (N_18198,N_13526,N_11962);
nand U18199 (N_18199,N_11502,N_11252);
nor U18200 (N_18200,N_14969,N_11238);
nor U18201 (N_18201,N_10457,N_10079);
xor U18202 (N_18202,N_10504,N_14425);
and U18203 (N_18203,N_10158,N_13415);
xnor U18204 (N_18204,N_13083,N_11745);
xor U18205 (N_18205,N_12509,N_12418);
xor U18206 (N_18206,N_11076,N_10721);
nand U18207 (N_18207,N_10600,N_10135);
or U18208 (N_18208,N_14803,N_13006);
and U18209 (N_18209,N_13314,N_14435);
and U18210 (N_18210,N_14618,N_10209);
or U18211 (N_18211,N_13025,N_12564);
nor U18212 (N_18212,N_12002,N_10999);
nor U18213 (N_18213,N_11505,N_14152);
and U18214 (N_18214,N_13495,N_14478);
xor U18215 (N_18215,N_13093,N_10433);
and U18216 (N_18216,N_11682,N_13012);
and U18217 (N_18217,N_12220,N_10942);
nor U18218 (N_18218,N_12242,N_10102);
xnor U18219 (N_18219,N_12228,N_14600);
nor U18220 (N_18220,N_10082,N_12602);
and U18221 (N_18221,N_11588,N_14002);
and U18222 (N_18222,N_12673,N_14822);
or U18223 (N_18223,N_12084,N_10166);
or U18224 (N_18224,N_13877,N_13730);
nand U18225 (N_18225,N_10459,N_10848);
nand U18226 (N_18226,N_10843,N_12026);
nor U18227 (N_18227,N_11035,N_10643);
xor U18228 (N_18228,N_14228,N_13930);
nand U18229 (N_18229,N_10732,N_11550);
xor U18230 (N_18230,N_13827,N_10070);
or U18231 (N_18231,N_12225,N_12740);
or U18232 (N_18232,N_13050,N_12295);
or U18233 (N_18233,N_11159,N_14766);
nand U18234 (N_18234,N_12034,N_12914);
xnor U18235 (N_18235,N_10516,N_14872);
and U18236 (N_18236,N_13859,N_11401);
nand U18237 (N_18237,N_11924,N_10370);
and U18238 (N_18238,N_10528,N_14031);
xor U18239 (N_18239,N_14009,N_10440);
nand U18240 (N_18240,N_14812,N_13709);
nor U18241 (N_18241,N_13782,N_14764);
and U18242 (N_18242,N_14715,N_13775);
and U18243 (N_18243,N_11157,N_14216);
nand U18244 (N_18244,N_11218,N_12244);
nand U18245 (N_18245,N_12906,N_13842);
and U18246 (N_18246,N_14254,N_14768);
nor U18247 (N_18247,N_10483,N_12142);
or U18248 (N_18248,N_14702,N_10399);
and U18249 (N_18249,N_11821,N_14248);
xor U18250 (N_18250,N_11012,N_11493);
or U18251 (N_18251,N_13805,N_14837);
nand U18252 (N_18252,N_14063,N_12830);
xor U18253 (N_18253,N_10643,N_10783);
or U18254 (N_18254,N_13631,N_13634);
or U18255 (N_18255,N_10483,N_14385);
nor U18256 (N_18256,N_11998,N_11880);
and U18257 (N_18257,N_13358,N_10460);
xor U18258 (N_18258,N_14528,N_13631);
or U18259 (N_18259,N_11869,N_14612);
xor U18260 (N_18260,N_12505,N_13669);
xnor U18261 (N_18261,N_10595,N_10160);
and U18262 (N_18262,N_10134,N_14942);
xnor U18263 (N_18263,N_13246,N_14668);
or U18264 (N_18264,N_14765,N_13481);
nand U18265 (N_18265,N_13595,N_10531);
and U18266 (N_18266,N_11553,N_12512);
or U18267 (N_18267,N_10676,N_13035);
or U18268 (N_18268,N_12165,N_12831);
and U18269 (N_18269,N_13710,N_13380);
or U18270 (N_18270,N_13718,N_13721);
nor U18271 (N_18271,N_12894,N_14821);
or U18272 (N_18272,N_13758,N_10062);
nor U18273 (N_18273,N_14635,N_14534);
nand U18274 (N_18274,N_11043,N_10645);
xor U18275 (N_18275,N_12568,N_13257);
nor U18276 (N_18276,N_10626,N_12040);
or U18277 (N_18277,N_13012,N_12583);
nor U18278 (N_18278,N_10451,N_14612);
xor U18279 (N_18279,N_12795,N_10049);
or U18280 (N_18280,N_14269,N_13142);
or U18281 (N_18281,N_11613,N_11300);
nor U18282 (N_18282,N_10646,N_13406);
nor U18283 (N_18283,N_10177,N_13303);
xor U18284 (N_18284,N_11995,N_10087);
and U18285 (N_18285,N_10226,N_14680);
xor U18286 (N_18286,N_14846,N_10007);
nand U18287 (N_18287,N_10075,N_10860);
and U18288 (N_18288,N_10812,N_12928);
xnor U18289 (N_18289,N_14590,N_13174);
nor U18290 (N_18290,N_12747,N_11212);
nor U18291 (N_18291,N_13862,N_14044);
nand U18292 (N_18292,N_12347,N_13527);
xnor U18293 (N_18293,N_10201,N_12204);
and U18294 (N_18294,N_13087,N_14604);
xnor U18295 (N_18295,N_14687,N_10349);
and U18296 (N_18296,N_12757,N_11391);
nor U18297 (N_18297,N_10223,N_11117);
or U18298 (N_18298,N_10494,N_13063);
nand U18299 (N_18299,N_12387,N_13513);
nor U18300 (N_18300,N_12450,N_12338);
nor U18301 (N_18301,N_13171,N_14221);
and U18302 (N_18302,N_13155,N_10108);
and U18303 (N_18303,N_12113,N_13407);
nor U18304 (N_18304,N_10733,N_11225);
nor U18305 (N_18305,N_11142,N_13673);
and U18306 (N_18306,N_12823,N_10660);
xor U18307 (N_18307,N_13079,N_13975);
or U18308 (N_18308,N_13280,N_10989);
nand U18309 (N_18309,N_13542,N_10754);
or U18310 (N_18310,N_13077,N_14740);
xnor U18311 (N_18311,N_13783,N_14655);
and U18312 (N_18312,N_11184,N_12089);
nor U18313 (N_18313,N_11873,N_10679);
xnor U18314 (N_18314,N_10263,N_10980);
nor U18315 (N_18315,N_14341,N_13359);
or U18316 (N_18316,N_10114,N_14767);
xnor U18317 (N_18317,N_13652,N_14880);
and U18318 (N_18318,N_12905,N_10111);
and U18319 (N_18319,N_10975,N_10006);
nor U18320 (N_18320,N_10061,N_13227);
nand U18321 (N_18321,N_11888,N_13644);
xor U18322 (N_18322,N_11645,N_12184);
and U18323 (N_18323,N_11121,N_13301);
and U18324 (N_18324,N_12189,N_12290);
nor U18325 (N_18325,N_11510,N_14681);
xor U18326 (N_18326,N_11851,N_10347);
or U18327 (N_18327,N_11251,N_14615);
nand U18328 (N_18328,N_12271,N_14438);
xor U18329 (N_18329,N_14701,N_14283);
xor U18330 (N_18330,N_13774,N_14409);
and U18331 (N_18331,N_13163,N_14134);
or U18332 (N_18332,N_12521,N_10856);
or U18333 (N_18333,N_13901,N_11581);
nand U18334 (N_18334,N_12991,N_12164);
nand U18335 (N_18335,N_11479,N_10035);
nand U18336 (N_18336,N_12425,N_13293);
nor U18337 (N_18337,N_10233,N_11835);
nand U18338 (N_18338,N_12564,N_14960);
nand U18339 (N_18339,N_14175,N_11717);
or U18340 (N_18340,N_11093,N_13875);
nand U18341 (N_18341,N_13406,N_13703);
nor U18342 (N_18342,N_14931,N_14652);
nor U18343 (N_18343,N_10496,N_11498);
and U18344 (N_18344,N_14406,N_10416);
or U18345 (N_18345,N_11804,N_12123);
xor U18346 (N_18346,N_11291,N_14940);
xnor U18347 (N_18347,N_13396,N_11923);
nor U18348 (N_18348,N_12303,N_14100);
xnor U18349 (N_18349,N_14511,N_10457);
nand U18350 (N_18350,N_10940,N_12798);
and U18351 (N_18351,N_10573,N_10888);
nand U18352 (N_18352,N_10453,N_11319);
or U18353 (N_18353,N_11143,N_13748);
nor U18354 (N_18354,N_10290,N_11980);
xnor U18355 (N_18355,N_11268,N_10556);
or U18356 (N_18356,N_12198,N_11794);
nand U18357 (N_18357,N_11743,N_14904);
xnor U18358 (N_18358,N_11502,N_12406);
nor U18359 (N_18359,N_11818,N_10199);
xor U18360 (N_18360,N_11078,N_11149);
and U18361 (N_18361,N_10045,N_11586);
nor U18362 (N_18362,N_10634,N_10635);
nand U18363 (N_18363,N_14249,N_10750);
and U18364 (N_18364,N_10043,N_13616);
nor U18365 (N_18365,N_12699,N_13048);
xor U18366 (N_18366,N_12551,N_14856);
nor U18367 (N_18367,N_11686,N_11317);
nor U18368 (N_18368,N_11421,N_13898);
and U18369 (N_18369,N_14303,N_12162);
or U18370 (N_18370,N_12093,N_12145);
nor U18371 (N_18371,N_11749,N_10929);
or U18372 (N_18372,N_10926,N_13106);
and U18373 (N_18373,N_11252,N_11230);
xor U18374 (N_18374,N_10741,N_11358);
xor U18375 (N_18375,N_10790,N_10073);
nand U18376 (N_18376,N_13515,N_11562);
nor U18377 (N_18377,N_12107,N_14773);
or U18378 (N_18378,N_13085,N_10831);
xnor U18379 (N_18379,N_14349,N_13060);
or U18380 (N_18380,N_14771,N_12149);
xor U18381 (N_18381,N_12620,N_12694);
xnor U18382 (N_18382,N_12089,N_11968);
nor U18383 (N_18383,N_10219,N_12831);
and U18384 (N_18384,N_13212,N_14481);
and U18385 (N_18385,N_10908,N_13464);
or U18386 (N_18386,N_11477,N_12090);
and U18387 (N_18387,N_14150,N_12958);
xnor U18388 (N_18388,N_11841,N_13393);
or U18389 (N_18389,N_11712,N_11963);
nand U18390 (N_18390,N_14032,N_11464);
nor U18391 (N_18391,N_12051,N_14267);
or U18392 (N_18392,N_13077,N_12508);
nand U18393 (N_18393,N_11961,N_11812);
nand U18394 (N_18394,N_13958,N_14730);
and U18395 (N_18395,N_10753,N_14258);
xor U18396 (N_18396,N_12660,N_12185);
xor U18397 (N_18397,N_14527,N_11625);
and U18398 (N_18398,N_11056,N_10468);
or U18399 (N_18399,N_12214,N_10336);
and U18400 (N_18400,N_14183,N_10424);
or U18401 (N_18401,N_14622,N_14785);
xnor U18402 (N_18402,N_10372,N_11895);
nor U18403 (N_18403,N_14943,N_14434);
nand U18404 (N_18404,N_10476,N_13273);
nand U18405 (N_18405,N_11175,N_14660);
xor U18406 (N_18406,N_10518,N_10928);
or U18407 (N_18407,N_11710,N_12443);
xor U18408 (N_18408,N_12830,N_13202);
nand U18409 (N_18409,N_11050,N_13890);
xnor U18410 (N_18410,N_10090,N_12460);
and U18411 (N_18411,N_12775,N_12453);
nand U18412 (N_18412,N_13175,N_14847);
xor U18413 (N_18413,N_14608,N_13018);
nor U18414 (N_18414,N_10498,N_11629);
nand U18415 (N_18415,N_13383,N_10994);
nand U18416 (N_18416,N_11518,N_11643);
or U18417 (N_18417,N_11773,N_11903);
xor U18418 (N_18418,N_12322,N_10177);
nor U18419 (N_18419,N_12092,N_13503);
or U18420 (N_18420,N_14227,N_11186);
nand U18421 (N_18421,N_13052,N_10615);
xnor U18422 (N_18422,N_11082,N_10974);
or U18423 (N_18423,N_10788,N_10052);
nor U18424 (N_18424,N_10978,N_14579);
nand U18425 (N_18425,N_14710,N_13735);
nand U18426 (N_18426,N_14568,N_10820);
nand U18427 (N_18427,N_12785,N_11341);
or U18428 (N_18428,N_14437,N_10838);
nand U18429 (N_18429,N_12109,N_11733);
and U18430 (N_18430,N_10162,N_14685);
nor U18431 (N_18431,N_12004,N_12130);
nand U18432 (N_18432,N_10689,N_13218);
and U18433 (N_18433,N_13929,N_12658);
or U18434 (N_18434,N_13979,N_13521);
nor U18435 (N_18435,N_13490,N_13876);
and U18436 (N_18436,N_13694,N_12771);
xnor U18437 (N_18437,N_11443,N_14584);
or U18438 (N_18438,N_12118,N_12316);
and U18439 (N_18439,N_14619,N_12493);
nand U18440 (N_18440,N_14823,N_10166);
xor U18441 (N_18441,N_13637,N_11195);
xor U18442 (N_18442,N_14083,N_10634);
xor U18443 (N_18443,N_10392,N_13211);
nand U18444 (N_18444,N_10085,N_14590);
and U18445 (N_18445,N_14886,N_12726);
or U18446 (N_18446,N_14866,N_13490);
or U18447 (N_18447,N_12958,N_12829);
nor U18448 (N_18448,N_13710,N_10960);
or U18449 (N_18449,N_14980,N_14661);
and U18450 (N_18450,N_12801,N_14911);
xor U18451 (N_18451,N_13340,N_10922);
and U18452 (N_18452,N_13848,N_10970);
or U18453 (N_18453,N_12205,N_13804);
and U18454 (N_18454,N_11536,N_12323);
nor U18455 (N_18455,N_12799,N_14372);
nand U18456 (N_18456,N_12462,N_13277);
nand U18457 (N_18457,N_14906,N_10577);
nand U18458 (N_18458,N_10473,N_11805);
nor U18459 (N_18459,N_14114,N_11844);
xnor U18460 (N_18460,N_11491,N_14187);
nor U18461 (N_18461,N_10406,N_13523);
nand U18462 (N_18462,N_11314,N_12658);
nor U18463 (N_18463,N_11170,N_10330);
and U18464 (N_18464,N_10356,N_10039);
or U18465 (N_18465,N_10077,N_14182);
nor U18466 (N_18466,N_10392,N_13393);
and U18467 (N_18467,N_12774,N_10128);
and U18468 (N_18468,N_13873,N_13936);
and U18469 (N_18469,N_12615,N_13927);
nand U18470 (N_18470,N_14147,N_13206);
nand U18471 (N_18471,N_13483,N_12283);
nand U18472 (N_18472,N_13310,N_13677);
or U18473 (N_18473,N_11414,N_12835);
nand U18474 (N_18474,N_13031,N_11339);
nor U18475 (N_18475,N_12630,N_12680);
or U18476 (N_18476,N_14450,N_10205);
or U18477 (N_18477,N_12787,N_10069);
nor U18478 (N_18478,N_12309,N_13896);
xor U18479 (N_18479,N_13817,N_12304);
xnor U18480 (N_18480,N_13198,N_10147);
nand U18481 (N_18481,N_12656,N_14484);
nor U18482 (N_18482,N_14679,N_10585);
xor U18483 (N_18483,N_12783,N_13744);
xor U18484 (N_18484,N_13589,N_11297);
xnor U18485 (N_18485,N_13890,N_11924);
or U18486 (N_18486,N_13760,N_12141);
or U18487 (N_18487,N_10832,N_14338);
nor U18488 (N_18488,N_13230,N_10385);
xnor U18489 (N_18489,N_12638,N_11703);
xnor U18490 (N_18490,N_11499,N_10270);
and U18491 (N_18491,N_11979,N_11282);
and U18492 (N_18492,N_12306,N_14015);
nand U18493 (N_18493,N_13028,N_12811);
and U18494 (N_18494,N_11724,N_10045);
or U18495 (N_18495,N_13626,N_11660);
or U18496 (N_18496,N_11993,N_10183);
nor U18497 (N_18497,N_10710,N_14587);
or U18498 (N_18498,N_11315,N_12652);
or U18499 (N_18499,N_12236,N_13230);
and U18500 (N_18500,N_14524,N_10842);
nand U18501 (N_18501,N_12458,N_10855);
nor U18502 (N_18502,N_11559,N_13082);
nand U18503 (N_18503,N_13923,N_14334);
and U18504 (N_18504,N_13020,N_12352);
nor U18505 (N_18505,N_11732,N_10560);
or U18506 (N_18506,N_10599,N_12928);
xor U18507 (N_18507,N_12111,N_10524);
nand U18508 (N_18508,N_11737,N_10100);
nor U18509 (N_18509,N_10180,N_14730);
nand U18510 (N_18510,N_12118,N_11838);
nor U18511 (N_18511,N_11032,N_14429);
and U18512 (N_18512,N_13925,N_10773);
nand U18513 (N_18513,N_14302,N_14265);
nor U18514 (N_18514,N_12066,N_11580);
nor U18515 (N_18515,N_11097,N_10455);
xor U18516 (N_18516,N_12429,N_10059);
or U18517 (N_18517,N_14733,N_11750);
or U18518 (N_18518,N_11960,N_14138);
or U18519 (N_18519,N_13040,N_11728);
xor U18520 (N_18520,N_12471,N_13891);
or U18521 (N_18521,N_14055,N_14231);
nand U18522 (N_18522,N_10606,N_12215);
xor U18523 (N_18523,N_14398,N_12065);
nand U18524 (N_18524,N_13588,N_12830);
nor U18525 (N_18525,N_14560,N_12261);
and U18526 (N_18526,N_10667,N_12390);
or U18527 (N_18527,N_11807,N_13713);
nor U18528 (N_18528,N_14777,N_13978);
or U18529 (N_18529,N_11942,N_10142);
or U18530 (N_18530,N_12492,N_11760);
nand U18531 (N_18531,N_13475,N_11110);
and U18532 (N_18532,N_11827,N_13580);
or U18533 (N_18533,N_14729,N_13261);
and U18534 (N_18534,N_12003,N_14930);
and U18535 (N_18535,N_14725,N_11751);
and U18536 (N_18536,N_12174,N_13196);
or U18537 (N_18537,N_11707,N_10309);
xnor U18538 (N_18538,N_11553,N_13071);
nand U18539 (N_18539,N_12086,N_14629);
and U18540 (N_18540,N_11907,N_10220);
or U18541 (N_18541,N_10774,N_10507);
xor U18542 (N_18542,N_13558,N_13925);
nor U18543 (N_18543,N_11493,N_13072);
nor U18544 (N_18544,N_12905,N_11253);
xnor U18545 (N_18545,N_12912,N_11907);
nand U18546 (N_18546,N_12019,N_14976);
nor U18547 (N_18547,N_13468,N_12843);
nor U18548 (N_18548,N_12076,N_10384);
or U18549 (N_18549,N_14043,N_10554);
nand U18550 (N_18550,N_14413,N_14079);
xor U18551 (N_18551,N_13843,N_14493);
nor U18552 (N_18552,N_10396,N_13581);
nand U18553 (N_18553,N_13678,N_12596);
nand U18554 (N_18554,N_14560,N_11751);
nor U18555 (N_18555,N_10794,N_14298);
or U18556 (N_18556,N_11341,N_12044);
nor U18557 (N_18557,N_13105,N_11313);
nand U18558 (N_18558,N_12583,N_11532);
nor U18559 (N_18559,N_14055,N_13533);
xor U18560 (N_18560,N_13416,N_13628);
or U18561 (N_18561,N_11132,N_14437);
nand U18562 (N_18562,N_10222,N_12013);
xnor U18563 (N_18563,N_11092,N_13700);
and U18564 (N_18564,N_14063,N_14851);
or U18565 (N_18565,N_14816,N_12752);
nor U18566 (N_18566,N_14145,N_10487);
xor U18567 (N_18567,N_10966,N_13829);
xor U18568 (N_18568,N_11811,N_14289);
or U18569 (N_18569,N_13308,N_14249);
nand U18570 (N_18570,N_12724,N_11440);
nand U18571 (N_18571,N_13375,N_14305);
and U18572 (N_18572,N_14428,N_12820);
and U18573 (N_18573,N_13079,N_11212);
nor U18574 (N_18574,N_14038,N_11952);
and U18575 (N_18575,N_11573,N_14997);
nand U18576 (N_18576,N_10743,N_11875);
and U18577 (N_18577,N_14036,N_11575);
and U18578 (N_18578,N_12955,N_14979);
and U18579 (N_18579,N_14565,N_13686);
nand U18580 (N_18580,N_13871,N_13191);
and U18581 (N_18581,N_14859,N_14511);
nor U18582 (N_18582,N_12452,N_11985);
nor U18583 (N_18583,N_14629,N_11457);
xnor U18584 (N_18584,N_14291,N_13159);
or U18585 (N_18585,N_12434,N_14708);
nor U18586 (N_18586,N_13658,N_14595);
or U18587 (N_18587,N_12781,N_12590);
or U18588 (N_18588,N_10671,N_13203);
nor U18589 (N_18589,N_13475,N_14864);
nor U18590 (N_18590,N_10231,N_12888);
nand U18591 (N_18591,N_14738,N_11451);
nand U18592 (N_18592,N_12272,N_13488);
nand U18593 (N_18593,N_10810,N_12340);
and U18594 (N_18594,N_14945,N_12056);
nor U18595 (N_18595,N_13643,N_13408);
nor U18596 (N_18596,N_11609,N_13111);
or U18597 (N_18597,N_13160,N_12783);
and U18598 (N_18598,N_13075,N_14765);
nor U18599 (N_18599,N_14076,N_12965);
nor U18600 (N_18600,N_10522,N_13258);
nand U18601 (N_18601,N_13895,N_12133);
xnor U18602 (N_18602,N_12503,N_10232);
xor U18603 (N_18603,N_12838,N_11241);
nand U18604 (N_18604,N_11247,N_10875);
or U18605 (N_18605,N_11268,N_10520);
nand U18606 (N_18606,N_11398,N_14237);
and U18607 (N_18607,N_12312,N_10003);
nor U18608 (N_18608,N_11090,N_10738);
nand U18609 (N_18609,N_12341,N_11309);
nand U18610 (N_18610,N_13551,N_13202);
nor U18611 (N_18611,N_11197,N_11899);
xor U18612 (N_18612,N_13371,N_10540);
or U18613 (N_18613,N_13770,N_12088);
and U18614 (N_18614,N_12592,N_12967);
nand U18615 (N_18615,N_12035,N_14503);
nand U18616 (N_18616,N_14460,N_10856);
and U18617 (N_18617,N_13523,N_14487);
or U18618 (N_18618,N_12957,N_13651);
and U18619 (N_18619,N_10085,N_14634);
and U18620 (N_18620,N_11470,N_10778);
and U18621 (N_18621,N_12198,N_10587);
and U18622 (N_18622,N_14293,N_10516);
xor U18623 (N_18623,N_10710,N_11671);
xor U18624 (N_18624,N_12086,N_12749);
nand U18625 (N_18625,N_10163,N_12125);
and U18626 (N_18626,N_12375,N_10028);
nor U18627 (N_18627,N_14448,N_11631);
xor U18628 (N_18628,N_12736,N_11364);
xnor U18629 (N_18629,N_10974,N_14436);
or U18630 (N_18630,N_13496,N_12827);
or U18631 (N_18631,N_13508,N_12355);
or U18632 (N_18632,N_10138,N_11287);
xnor U18633 (N_18633,N_10562,N_11724);
nor U18634 (N_18634,N_11352,N_10696);
and U18635 (N_18635,N_14300,N_10829);
nor U18636 (N_18636,N_14115,N_10750);
nand U18637 (N_18637,N_13464,N_10681);
and U18638 (N_18638,N_12162,N_14327);
or U18639 (N_18639,N_14893,N_14198);
or U18640 (N_18640,N_10049,N_11990);
and U18641 (N_18641,N_12099,N_13689);
nand U18642 (N_18642,N_14547,N_11714);
or U18643 (N_18643,N_10260,N_10318);
nor U18644 (N_18644,N_13678,N_11694);
or U18645 (N_18645,N_12707,N_13899);
xnor U18646 (N_18646,N_13711,N_12423);
xnor U18647 (N_18647,N_12542,N_12207);
nand U18648 (N_18648,N_11817,N_10436);
and U18649 (N_18649,N_11963,N_13215);
nand U18650 (N_18650,N_11679,N_12951);
and U18651 (N_18651,N_11716,N_11318);
nor U18652 (N_18652,N_13519,N_10060);
nand U18653 (N_18653,N_12014,N_10738);
or U18654 (N_18654,N_12928,N_11333);
nor U18655 (N_18655,N_14327,N_14703);
nand U18656 (N_18656,N_12339,N_10851);
and U18657 (N_18657,N_10196,N_11200);
nand U18658 (N_18658,N_10917,N_10093);
nor U18659 (N_18659,N_12933,N_11661);
or U18660 (N_18660,N_14159,N_11378);
xnor U18661 (N_18661,N_13323,N_10590);
and U18662 (N_18662,N_11114,N_12488);
xor U18663 (N_18663,N_11372,N_10850);
and U18664 (N_18664,N_13084,N_13665);
or U18665 (N_18665,N_12480,N_10035);
and U18666 (N_18666,N_11520,N_12079);
nand U18667 (N_18667,N_10292,N_14478);
xor U18668 (N_18668,N_12301,N_12437);
and U18669 (N_18669,N_11578,N_11190);
xor U18670 (N_18670,N_14729,N_13011);
xnor U18671 (N_18671,N_11787,N_10717);
or U18672 (N_18672,N_11386,N_10769);
or U18673 (N_18673,N_10536,N_14815);
nor U18674 (N_18674,N_14321,N_10545);
and U18675 (N_18675,N_13174,N_11620);
or U18676 (N_18676,N_13314,N_10913);
nor U18677 (N_18677,N_13488,N_14901);
and U18678 (N_18678,N_10700,N_10166);
and U18679 (N_18679,N_10389,N_12484);
nand U18680 (N_18680,N_13887,N_10129);
xnor U18681 (N_18681,N_14521,N_11167);
and U18682 (N_18682,N_13516,N_13028);
nor U18683 (N_18683,N_12422,N_13559);
xor U18684 (N_18684,N_13253,N_11500);
nor U18685 (N_18685,N_13312,N_10824);
nor U18686 (N_18686,N_14601,N_13875);
nand U18687 (N_18687,N_12329,N_14264);
nor U18688 (N_18688,N_12072,N_14372);
nor U18689 (N_18689,N_14213,N_13481);
or U18690 (N_18690,N_13468,N_14977);
and U18691 (N_18691,N_12321,N_12678);
nor U18692 (N_18692,N_10640,N_14529);
and U18693 (N_18693,N_14100,N_11205);
xor U18694 (N_18694,N_13563,N_13786);
or U18695 (N_18695,N_10522,N_14046);
and U18696 (N_18696,N_10259,N_10713);
nand U18697 (N_18697,N_13419,N_13073);
nand U18698 (N_18698,N_14881,N_14135);
and U18699 (N_18699,N_11978,N_10100);
or U18700 (N_18700,N_14834,N_11427);
nand U18701 (N_18701,N_13353,N_11498);
nand U18702 (N_18702,N_12074,N_13758);
or U18703 (N_18703,N_10120,N_12243);
xnor U18704 (N_18704,N_11264,N_13497);
nand U18705 (N_18705,N_12101,N_12354);
and U18706 (N_18706,N_12413,N_11825);
xnor U18707 (N_18707,N_13127,N_13591);
or U18708 (N_18708,N_14736,N_10770);
and U18709 (N_18709,N_14396,N_12466);
and U18710 (N_18710,N_13451,N_10329);
or U18711 (N_18711,N_13580,N_10295);
nand U18712 (N_18712,N_14384,N_13780);
or U18713 (N_18713,N_12680,N_10968);
xnor U18714 (N_18714,N_10284,N_12603);
nor U18715 (N_18715,N_13689,N_10414);
nor U18716 (N_18716,N_13033,N_13457);
or U18717 (N_18717,N_12471,N_10896);
xnor U18718 (N_18718,N_13565,N_14954);
and U18719 (N_18719,N_11983,N_13158);
nand U18720 (N_18720,N_10725,N_12481);
nand U18721 (N_18721,N_12596,N_13539);
nand U18722 (N_18722,N_10417,N_13971);
nor U18723 (N_18723,N_14023,N_14480);
nand U18724 (N_18724,N_14369,N_12224);
xor U18725 (N_18725,N_11572,N_14051);
xor U18726 (N_18726,N_13358,N_12485);
and U18727 (N_18727,N_12443,N_10087);
xor U18728 (N_18728,N_12014,N_14720);
xnor U18729 (N_18729,N_14326,N_10093);
nor U18730 (N_18730,N_11087,N_10166);
nor U18731 (N_18731,N_10128,N_11443);
nand U18732 (N_18732,N_14786,N_11498);
or U18733 (N_18733,N_11327,N_14579);
xnor U18734 (N_18734,N_11454,N_12160);
xnor U18735 (N_18735,N_12431,N_14519);
and U18736 (N_18736,N_13692,N_14430);
nand U18737 (N_18737,N_14194,N_13474);
nand U18738 (N_18738,N_10856,N_14631);
nand U18739 (N_18739,N_11648,N_12377);
and U18740 (N_18740,N_10929,N_14871);
or U18741 (N_18741,N_13592,N_14665);
nand U18742 (N_18742,N_13864,N_13112);
or U18743 (N_18743,N_14251,N_13375);
xor U18744 (N_18744,N_14827,N_10869);
nor U18745 (N_18745,N_14332,N_13677);
xnor U18746 (N_18746,N_12476,N_12283);
xor U18747 (N_18747,N_13377,N_11503);
nor U18748 (N_18748,N_14550,N_14649);
nor U18749 (N_18749,N_14488,N_12367);
and U18750 (N_18750,N_13567,N_10886);
nor U18751 (N_18751,N_14094,N_13713);
xor U18752 (N_18752,N_12713,N_11006);
or U18753 (N_18753,N_10248,N_14390);
xor U18754 (N_18754,N_14914,N_14483);
nor U18755 (N_18755,N_12075,N_14555);
nor U18756 (N_18756,N_14345,N_13837);
or U18757 (N_18757,N_11289,N_14797);
nor U18758 (N_18758,N_11492,N_12760);
xor U18759 (N_18759,N_10014,N_11563);
and U18760 (N_18760,N_13020,N_10117);
and U18761 (N_18761,N_13066,N_12370);
nand U18762 (N_18762,N_13779,N_10571);
nand U18763 (N_18763,N_11996,N_13526);
xnor U18764 (N_18764,N_13277,N_10530);
and U18765 (N_18765,N_14529,N_11667);
or U18766 (N_18766,N_10701,N_13486);
and U18767 (N_18767,N_14484,N_14878);
nand U18768 (N_18768,N_14499,N_11211);
or U18769 (N_18769,N_14525,N_12067);
xnor U18770 (N_18770,N_12071,N_10640);
or U18771 (N_18771,N_10597,N_14933);
or U18772 (N_18772,N_13705,N_14704);
xnor U18773 (N_18773,N_10712,N_10749);
or U18774 (N_18774,N_10704,N_12355);
nand U18775 (N_18775,N_11860,N_12757);
and U18776 (N_18776,N_10402,N_11301);
xor U18777 (N_18777,N_13608,N_14396);
and U18778 (N_18778,N_13920,N_14894);
and U18779 (N_18779,N_12746,N_14953);
xnor U18780 (N_18780,N_14970,N_13612);
and U18781 (N_18781,N_14943,N_13691);
and U18782 (N_18782,N_12896,N_10492);
nand U18783 (N_18783,N_10864,N_13631);
and U18784 (N_18784,N_12288,N_14344);
nor U18785 (N_18785,N_11700,N_13881);
or U18786 (N_18786,N_10869,N_10635);
or U18787 (N_18787,N_12452,N_10196);
xnor U18788 (N_18788,N_12591,N_10732);
nor U18789 (N_18789,N_12439,N_12737);
nand U18790 (N_18790,N_12223,N_12010);
nor U18791 (N_18791,N_10899,N_13858);
or U18792 (N_18792,N_12568,N_11031);
and U18793 (N_18793,N_10281,N_13918);
and U18794 (N_18794,N_12058,N_11397);
xnor U18795 (N_18795,N_10260,N_12887);
or U18796 (N_18796,N_13255,N_11121);
xnor U18797 (N_18797,N_12937,N_10738);
or U18798 (N_18798,N_13329,N_14764);
nand U18799 (N_18799,N_12399,N_10150);
nand U18800 (N_18800,N_11156,N_13730);
nor U18801 (N_18801,N_13269,N_12112);
xnor U18802 (N_18802,N_14834,N_13947);
and U18803 (N_18803,N_12987,N_12242);
nor U18804 (N_18804,N_10480,N_12994);
or U18805 (N_18805,N_14648,N_12139);
and U18806 (N_18806,N_12135,N_10399);
and U18807 (N_18807,N_10071,N_12692);
xor U18808 (N_18808,N_10934,N_13713);
xor U18809 (N_18809,N_13009,N_13919);
nor U18810 (N_18810,N_14163,N_13819);
or U18811 (N_18811,N_14421,N_13781);
xnor U18812 (N_18812,N_14170,N_13226);
or U18813 (N_18813,N_13660,N_10083);
nor U18814 (N_18814,N_13464,N_10597);
nor U18815 (N_18815,N_14643,N_11852);
and U18816 (N_18816,N_12194,N_12750);
and U18817 (N_18817,N_12580,N_10701);
or U18818 (N_18818,N_11834,N_13795);
nand U18819 (N_18819,N_11775,N_14335);
nor U18820 (N_18820,N_11100,N_12363);
nor U18821 (N_18821,N_11657,N_11633);
or U18822 (N_18822,N_13287,N_13021);
or U18823 (N_18823,N_12440,N_13127);
and U18824 (N_18824,N_14491,N_14910);
xor U18825 (N_18825,N_11107,N_14277);
xnor U18826 (N_18826,N_11892,N_13610);
nand U18827 (N_18827,N_13289,N_13520);
nor U18828 (N_18828,N_13055,N_10792);
and U18829 (N_18829,N_11297,N_10731);
nor U18830 (N_18830,N_13272,N_13313);
nor U18831 (N_18831,N_14241,N_11799);
xor U18832 (N_18832,N_14284,N_12726);
and U18833 (N_18833,N_14258,N_13909);
or U18834 (N_18834,N_13230,N_10600);
or U18835 (N_18835,N_14313,N_12080);
nor U18836 (N_18836,N_11089,N_10674);
or U18837 (N_18837,N_11172,N_14250);
or U18838 (N_18838,N_13578,N_14006);
nand U18839 (N_18839,N_14919,N_12468);
or U18840 (N_18840,N_10404,N_14344);
nand U18841 (N_18841,N_13859,N_11477);
nor U18842 (N_18842,N_13235,N_14571);
nor U18843 (N_18843,N_14825,N_13000);
and U18844 (N_18844,N_12566,N_13430);
or U18845 (N_18845,N_14540,N_13581);
or U18846 (N_18846,N_13497,N_10538);
and U18847 (N_18847,N_12499,N_11915);
or U18848 (N_18848,N_12584,N_12024);
nor U18849 (N_18849,N_13993,N_10346);
or U18850 (N_18850,N_11293,N_10892);
nand U18851 (N_18851,N_10146,N_13611);
nor U18852 (N_18852,N_10510,N_13042);
or U18853 (N_18853,N_14857,N_10133);
xnor U18854 (N_18854,N_12281,N_14168);
and U18855 (N_18855,N_14589,N_12119);
nor U18856 (N_18856,N_12442,N_14757);
or U18857 (N_18857,N_13725,N_12490);
or U18858 (N_18858,N_10482,N_10023);
nand U18859 (N_18859,N_10559,N_12176);
and U18860 (N_18860,N_14383,N_10273);
xnor U18861 (N_18861,N_10363,N_11925);
and U18862 (N_18862,N_13796,N_12718);
xor U18863 (N_18863,N_10218,N_14901);
nand U18864 (N_18864,N_14129,N_14648);
nor U18865 (N_18865,N_10166,N_12347);
or U18866 (N_18866,N_10772,N_13731);
nor U18867 (N_18867,N_11626,N_13776);
and U18868 (N_18868,N_11242,N_12329);
nor U18869 (N_18869,N_14912,N_14709);
nor U18870 (N_18870,N_10629,N_14334);
nand U18871 (N_18871,N_11079,N_14613);
nor U18872 (N_18872,N_12231,N_11418);
nor U18873 (N_18873,N_13901,N_11833);
nor U18874 (N_18874,N_11395,N_13576);
and U18875 (N_18875,N_10802,N_11732);
or U18876 (N_18876,N_10582,N_14094);
and U18877 (N_18877,N_13551,N_13925);
nand U18878 (N_18878,N_12422,N_13200);
xnor U18879 (N_18879,N_10119,N_12352);
nor U18880 (N_18880,N_10340,N_10905);
nand U18881 (N_18881,N_12935,N_11578);
nand U18882 (N_18882,N_14556,N_12014);
nand U18883 (N_18883,N_11791,N_14753);
and U18884 (N_18884,N_14749,N_14303);
or U18885 (N_18885,N_13643,N_11645);
or U18886 (N_18886,N_10705,N_14598);
nor U18887 (N_18887,N_10526,N_11341);
nand U18888 (N_18888,N_14998,N_11243);
nand U18889 (N_18889,N_10003,N_13362);
nand U18890 (N_18890,N_10456,N_11190);
xor U18891 (N_18891,N_11774,N_13555);
nor U18892 (N_18892,N_14188,N_13027);
nor U18893 (N_18893,N_12745,N_12656);
xnor U18894 (N_18894,N_13113,N_11159);
xor U18895 (N_18895,N_11111,N_13928);
nor U18896 (N_18896,N_11528,N_13516);
nand U18897 (N_18897,N_14879,N_14098);
and U18898 (N_18898,N_13831,N_14021);
nor U18899 (N_18899,N_10048,N_13937);
xor U18900 (N_18900,N_10011,N_10341);
nand U18901 (N_18901,N_10180,N_12785);
nand U18902 (N_18902,N_10834,N_12851);
xor U18903 (N_18903,N_11256,N_11665);
nand U18904 (N_18904,N_13246,N_12856);
nand U18905 (N_18905,N_13945,N_11377);
and U18906 (N_18906,N_10561,N_14824);
nor U18907 (N_18907,N_11907,N_14634);
nor U18908 (N_18908,N_10531,N_13025);
xnor U18909 (N_18909,N_10956,N_11118);
nand U18910 (N_18910,N_12487,N_12780);
nand U18911 (N_18911,N_10753,N_11877);
nor U18912 (N_18912,N_10929,N_13259);
xor U18913 (N_18913,N_12357,N_14719);
nor U18914 (N_18914,N_12195,N_13933);
xor U18915 (N_18915,N_13587,N_10818);
xnor U18916 (N_18916,N_12564,N_14187);
xnor U18917 (N_18917,N_11491,N_11985);
nor U18918 (N_18918,N_11717,N_12756);
or U18919 (N_18919,N_12897,N_12507);
or U18920 (N_18920,N_10456,N_14025);
nor U18921 (N_18921,N_10815,N_10412);
xor U18922 (N_18922,N_10177,N_14108);
or U18923 (N_18923,N_12142,N_11698);
and U18924 (N_18924,N_10448,N_14964);
and U18925 (N_18925,N_11758,N_14800);
or U18926 (N_18926,N_13163,N_11289);
nand U18927 (N_18927,N_14878,N_14801);
nand U18928 (N_18928,N_12347,N_10365);
or U18929 (N_18929,N_12168,N_13512);
and U18930 (N_18930,N_10077,N_14662);
nand U18931 (N_18931,N_10920,N_13527);
nor U18932 (N_18932,N_13729,N_10073);
or U18933 (N_18933,N_11131,N_11060);
or U18934 (N_18934,N_10608,N_10563);
and U18935 (N_18935,N_11911,N_11775);
and U18936 (N_18936,N_13144,N_10921);
and U18937 (N_18937,N_12971,N_10470);
or U18938 (N_18938,N_14203,N_13326);
nor U18939 (N_18939,N_12118,N_13998);
or U18940 (N_18940,N_11094,N_10444);
or U18941 (N_18941,N_10767,N_12891);
nand U18942 (N_18942,N_14318,N_11269);
or U18943 (N_18943,N_14262,N_14589);
nand U18944 (N_18944,N_11231,N_12220);
and U18945 (N_18945,N_12333,N_12750);
or U18946 (N_18946,N_14843,N_13293);
and U18947 (N_18947,N_14550,N_12748);
or U18948 (N_18948,N_13662,N_10313);
nor U18949 (N_18949,N_10024,N_14784);
and U18950 (N_18950,N_12271,N_13612);
xnor U18951 (N_18951,N_11585,N_14543);
and U18952 (N_18952,N_13076,N_14976);
nor U18953 (N_18953,N_10543,N_14207);
nor U18954 (N_18954,N_11030,N_12818);
nor U18955 (N_18955,N_12722,N_14031);
or U18956 (N_18956,N_14075,N_10232);
and U18957 (N_18957,N_11333,N_12710);
and U18958 (N_18958,N_10127,N_14104);
nand U18959 (N_18959,N_11698,N_12824);
or U18960 (N_18960,N_12236,N_11957);
or U18961 (N_18961,N_13840,N_14093);
nor U18962 (N_18962,N_10287,N_14426);
or U18963 (N_18963,N_10215,N_10439);
xor U18964 (N_18964,N_11974,N_13437);
nor U18965 (N_18965,N_14134,N_10106);
nor U18966 (N_18966,N_13017,N_10088);
nand U18967 (N_18967,N_10153,N_11758);
nor U18968 (N_18968,N_14231,N_12491);
nand U18969 (N_18969,N_14970,N_12081);
or U18970 (N_18970,N_13044,N_14669);
or U18971 (N_18971,N_13336,N_14811);
nor U18972 (N_18972,N_10810,N_11943);
and U18973 (N_18973,N_10489,N_12294);
and U18974 (N_18974,N_10151,N_10972);
and U18975 (N_18975,N_14850,N_14409);
nor U18976 (N_18976,N_10651,N_14503);
or U18977 (N_18977,N_10147,N_14281);
and U18978 (N_18978,N_13235,N_11774);
xnor U18979 (N_18979,N_10216,N_11193);
nor U18980 (N_18980,N_14095,N_14429);
or U18981 (N_18981,N_10858,N_13352);
nand U18982 (N_18982,N_11959,N_12462);
nand U18983 (N_18983,N_10197,N_11655);
or U18984 (N_18984,N_11760,N_13157);
nand U18985 (N_18985,N_14506,N_12267);
nor U18986 (N_18986,N_12081,N_12155);
or U18987 (N_18987,N_12164,N_13600);
or U18988 (N_18988,N_12557,N_13323);
nor U18989 (N_18989,N_10070,N_11719);
and U18990 (N_18990,N_11905,N_11196);
and U18991 (N_18991,N_10820,N_11245);
nor U18992 (N_18992,N_14898,N_11702);
xor U18993 (N_18993,N_11400,N_13333);
nand U18994 (N_18994,N_11272,N_14780);
nor U18995 (N_18995,N_10779,N_11813);
nor U18996 (N_18996,N_12689,N_14191);
nand U18997 (N_18997,N_11390,N_10720);
xnor U18998 (N_18998,N_13186,N_14829);
and U18999 (N_18999,N_12339,N_12608);
and U19000 (N_19000,N_10732,N_13080);
nor U19001 (N_19001,N_13172,N_13750);
xnor U19002 (N_19002,N_10382,N_12318);
or U19003 (N_19003,N_10350,N_11808);
and U19004 (N_19004,N_14937,N_11882);
or U19005 (N_19005,N_10729,N_10342);
nor U19006 (N_19006,N_11964,N_13422);
or U19007 (N_19007,N_13454,N_14655);
nor U19008 (N_19008,N_11980,N_10461);
nor U19009 (N_19009,N_12776,N_10309);
and U19010 (N_19010,N_14788,N_12488);
or U19011 (N_19011,N_10722,N_10933);
and U19012 (N_19012,N_12816,N_12036);
nand U19013 (N_19013,N_12350,N_10718);
xnor U19014 (N_19014,N_10675,N_13715);
xor U19015 (N_19015,N_14818,N_14720);
xnor U19016 (N_19016,N_14179,N_14910);
xnor U19017 (N_19017,N_14833,N_12140);
nor U19018 (N_19018,N_14382,N_12060);
xor U19019 (N_19019,N_14869,N_13328);
and U19020 (N_19020,N_10196,N_12333);
nor U19021 (N_19021,N_10118,N_13212);
nor U19022 (N_19022,N_12028,N_10517);
and U19023 (N_19023,N_14312,N_12337);
or U19024 (N_19024,N_13152,N_12518);
xor U19025 (N_19025,N_11669,N_10776);
nand U19026 (N_19026,N_11355,N_13284);
nor U19027 (N_19027,N_14915,N_11860);
nor U19028 (N_19028,N_10373,N_10557);
and U19029 (N_19029,N_13206,N_13087);
nand U19030 (N_19030,N_13864,N_11576);
xor U19031 (N_19031,N_10554,N_10739);
nor U19032 (N_19032,N_12415,N_14481);
xor U19033 (N_19033,N_13250,N_11171);
and U19034 (N_19034,N_11544,N_13986);
nor U19035 (N_19035,N_10739,N_10378);
and U19036 (N_19036,N_11461,N_12871);
or U19037 (N_19037,N_10331,N_10337);
xnor U19038 (N_19038,N_14819,N_14879);
nand U19039 (N_19039,N_12540,N_10924);
nand U19040 (N_19040,N_11581,N_12553);
nand U19041 (N_19041,N_10051,N_10334);
or U19042 (N_19042,N_13106,N_14376);
and U19043 (N_19043,N_10968,N_12797);
nor U19044 (N_19044,N_14054,N_11495);
or U19045 (N_19045,N_14899,N_12499);
nor U19046 (N_19046,N_10528,N_13220);
or U19047 (N_19047,N_13197,N_12940);
nor U19048 (N_19048,N_12948,N_11375);
xor U19049 (N_19049,N_12499,N_11291);
nor U19050 (N_19050,N_10512,N_13998);
and U19051 (N_19051,N_11835,N_10524);
nand U19052 (N_19052,N_13176,N_11448);
xor U19053 (N_19053,N_12267,N_14806);
xor U19054 (N_19054,N_13395,N_11028);
or U19055 (N_19055,N_12280,N_12201);
and U19056 (N_19056,N_14043,N_14025);
nor U19057 (N_19057,N_14034,N_14109);
xor U19058 (N_19058,N_12379,N_10997);
nor U19059 (N_19059,N_11839,N_14286);
xnor U19060 (N_19060,N_11292,N_14956);
xor U19061 (N_19061,N_11047,N_13935);
and U19062 (N_19062,N_14199,N_12176);
and U19063 (N_19063,N_13511,N_12241);
or U19064 (N_19064,N_11172,N_14026);
xnor U19065 (N_19065,N_14112,N_13589);
xor U19066 (N_19066,N_12791,N_14215);
or U19067 (N_19067,N_12199,N_13878);
and U19068 (N_19068,N_10131,N_11792);
xnor U19069 (N_19069,N_14872,N_14738);
nor U19070 (N_19070,N_14600,N_10435);
nand U19071 (N_19071,N_10498,N_14478);
nand U19072 (N_19072,N_10962,N_14873);
nand U19073 (N_19073,N_14842,N_10950);
or U19074 (N_19074,N_14139,N_10148);
or U19075 (N_19075,N_13414,N_12296);
or U19076 (N_19076,N_13819,N_13954);
or U19077 (N_19077,N_11169,N_12827);
nand U19078 (N_19078,N_10486,N_12100);
xnor U19079 (N_19079,N_10282,N_13167);
and U19080 (N_19080,N_11135,N_12701);
nor U19081 (N_19081,N_14051,N_14532);
and U19082 (N_19082,N_14361,N_13075);
or U19083 (N_19083,N_14287,N_12207);
xnor U19084 (N_19084,N_10491,N_10156);
nor U19085 (N_19085,N_11670,N_11610);
or U19086 (N_19086,N_12977,N_13147);
and U19087 (N_19087,N_13108,N_10250);
and U19088 (N_19088,N_14557,N_10409);
or U19089 (N_19089,N_10322,N_10755);
xnor U19090 (N_19090,N_10813,N_12276);
and U19091 (N_19091,N_13204,N_14563);
and U19092 (N_19092,N_13892,N_11581);
and U19093 (N_19093,N_13739,N_13750);
or U19094 (N_19094,N_13314,N_12801);
or U19095 (N_19095,N_11786,N_14573);
xnor U19096 (N_19096,N_11464,N_11967);
or U19097 (N_19097,N_11971,N_12721);
nand U19098 (N_19098,N_12714,N_11559);
or U19099 (N_19099,N_11757,N_12938);
xnor U19100 (N_19100,N_10377,N_13770);
nor U19101 (N_19101,N_11539,N_12647);
nand U19102 (N_19102,N_11986,N_14967);
nor U19103 (N_19103,N_10731,N_13781);
xor U19104 (N_19104,N_11105,N_10179);
nand U19105 (N_19105,N_11366,N_12338);
or U19106 (N_19106,N_14855,N_10717);
nand U19107 (N_19107,N_11908,N_14328);
and U19108 (N_19108,N_10116,N_11171);
nor U19109 (N_19109,N_14348,N_12218);
nand U19110 (N_19110,N_12675,N_12304);
and U19111 (N_19111,N_13515,N_12340);
xnor U19112 (N_19112,N_11393,N_10109);
xnor U19113 (N_19113,N_13414,N_13810);
nor U19114 (N_19114,N_11884,N_14826);
nand U19115 (N_19115,N_12308,N_10625);
nand U19116 (N_19116,N_11179,N_10807);
or U19117 (N_19117,N_12564,N_10470);
and U19118 (N_19118,N_14397,N_11068);
and U19119 (N_19119,N_13920,N_11544);
and U19120 (N_19120,N_11420,N_13345);
and U19121 (N_19121,N_11490,N_12527);
and U19122 (N_19122,N_13363,N_12935);
or U19123 (N_19123,N_11146,N_10317);
xnor U19124 (N_19124,N_14269,N_13227);
or U19125 (N_19125,N_11438,N_13443);
nand U19126 (N_19126,N_13537,N_11473);
nor U19127 (N_19127,N_14599,N_12849);
nor U19128 (N_19128,N_10824,N_14530);
xnor U19129 (N_19129,N_12698,N_12110);
nand U19130 (N_19130,N_10022,N_12974);
and U19131 (N_19131,N_12306,N_10921);
nor U19132 (N_19132,N_12275,N_11117);
nand U19133 (N_19133,N_11379,N_11002);
and U19134 (N_19134,N_13908,N_13174);
or U19135 (N_19135,N_11049,N_10750);
and U19136 (N_19136,N_11938,N_14132);
nand U19137 (N_19137,N_11632,N_10737);
or U19138 (N_19138,N_13458,N_13421);
nand U19139 (N_19139,N_12743,N_11653);
nor U19140 (N_19140,N_11729,N_13462);
nand U19141 (N_19141,N_13314,N_10664);
or U19142 (N_19142,N_12593,N_11906);
nor U19143 (N_19143,N_13938,N_14531);
and U19144 (N_19144,N_14239,N_11927);
xor U19145 (N_19145,N_14878,N_14330);
or U19146 (N_19146,N_11982,N_10993);
or U19147 (N_19147,N_13103,N_11162);
nor U19148 (N_19148,N_11122,N_13596);
and U19149 (N_19149,N_12711,N_12959);
or U19150 (N_19150,N_10463,N_11186);
and U19151 (N_19151,N_14812,N_14860);
nand U19152 (N_19152,N_13570,N_12157);
nor U19153 (N_19153,N_13868,N_12004);
nor U19154 (N_19154,N_12435,N_12335);
or U19155 (N_19155,N_13550,N_10117);
nor U19156 (N_19156,N_10970,N_14542);
xor U19157 (N_19157,N_10159,N_14511);
nand U19158 (N_19158,N_13078,N_11322);
nor U19159 (N_19159,N_11655,N_13674);
nor U19160 (N_19160,N_13533,N_10256);
xnor U19161 (N_19161,N_14665,N_12188);
nand U19162 (N_19162,N_12967,N_12666);
nor U19163 (N_19163,N_14003,N_11921);
xor U19164 (N_19164,N_13474,N_12189);
nand U19165 (N_19165,N_14907,N_14497);
or U19166 (N_19166,N_12844,N_12353);
and U19167 (N_19167,N_13492,N_10077);
nand U19168 (N_19168,N_12997,N_12540);
xnor U19169 (N_19169,N_10875,N_11194);
xnor U19170 (N_19170,N_12220,N_10388);
and U19171 (N_19171,N_13687,N_10525);
nor U19172 (N_19172,N_13227,N_12894);
nor U19173 (N_19173,N_12487,N_12270);
and U19174 (N_19174,N_14605,N_11950);
nor U19175 (N_19175,N_11686,N_13135);
and U19176 (N_19176,N_10443,N_11948);
nor U19177 (N_19177,N_11512,N_11264);
or U19178 (N_19178,N_11433,N_12246);
nand U19179 (N_19179,N_14458,N_11508);
nand U19180 (N_19180,N_12004,N_12544);
xor U19181 (N_19181,N_14931,N_10327);
xor U19182 (N_19182,N_12542,N_13980);
nor U19183 (N_19183,N_13482,N_11288);
nor U19184 (N_19184,N_14129,N_13092);
nor U19185 (N_19185,N_10196,N_10156);
and U19186 (N_19186,N_12874,N_13980);
xor U19187 (N_19187,N_11074,N_12039);
xnor U19188 (N_19188,N_12269,N_10200);
and U19189 (N_19189,N_14936,N_12409);
nand U19190 (N_19190,N_14452,N_13583);
or U19191 (N_19191,N_13099,N_12522);
or U19192 (N_19192,N_10152,N_12367);
and U19193 (N_19193,N_13884,N_11212);
and U19194 (N_19194,N_12301,N_11675);
xor U19195 (N_19195,N_13230,N_13100);
or U19196 (N_19196,N_12815,N_10039);
nor U19197 (N_19197,N_14768,N_10224);
nor U19198 (N_19198,N_11709,N_10506);
nor U19199 (N_19199,N_12083,N_11601);
or U19200 (N_19200,N_12003,N_13243);
xor U19201 (N_19201,N_12717,N_14124);
and U19202 (N_19202,N_14496,N_14173);
or U19203 (N_19203,N_10475,N_12100);
nand U19204 (N_19204,N_10094,N_12903);
nor U19205 (N_19205,N_12174,N_11923);
and U19206 (N_19206,N_14065,N_10715);
nor U19207 (N_19207,N_14488,N_14459);
xor U19208 (N_19208,N_14250,N_14468);
xor U19209 (N_19209,N_14323,N_10651);
xor U19210 (N_19210,N_11723,N_13040);
xor U19211 (N_19211,N_13417,N_12199);
nand U19212 (N_19212,N_10781,N_12398);
nand U19213 (N_19213,N_12537,N_13962);
nor U19214 (N_19214,N_13734,N_13180);
and U19215 (N_19215,N_12658,N_11701);
xnor U19216 (N_19216,N_10893,N_10789);
or U19217 (N_19217,N_11583,N_10337);
and U19218 (N_19218,N_12279,N_13320);
or U19219 (N_19219,N_11661,N_12842);
nand U19220 (N_19220,N_11163,N_11572);
or U19221 (N_19221,N_11439,N_11442);
xor U19222 (N_19222,N_14526,N_12861);
and U19223 (N_19223,N_13984,N_12615);
xor U19224 (N_19224,N_12464,N_14453);
and U19225 (N_19225,N_14617,N_13100);
nand U19226 (N_19226,N_14243,N_11646);
xnor U19227 (N_19227,N_10587,N_10572);
nand U19228 (N_19228,N_14721,N_13594);
xor U19229 (N_19229,N_14039,N_11049);
or U19230 (N_19230,N_11350,N_13641);
nor U19231 (N_19231,N_13788,N_11535);
or U19232 (N_19232,N_14603,N_14829);
xor U19233 (N_19233,N_14036,N_10815);
nand U19234 (N_19234,N_14652,N_10234);
nand U19235 (N_19235,N_11972,N_12280);
nand U19236 (N_19236,N_11172,N_10067);
nand U19237 (N_19237,N_10017,N_14337);
xor U19238 (N_19238,N_10244,N_10358);
or U19239 (N_19239,N_10655,N_10244);
nand U19240 (N_19240,N_12570,N_10049);
xnor U19241 (N_19241,N_10306,N_11471);
xnor U19242 (N_19242,N_14497,N_12031);
nand U19243 (N_19243,N_13676,N_14297);
or U19244 (N_19244,N_13417,N_10411);
nand U19245 (N_19245,N_13195,N_10256);
nor U19246 (N_19246,N_14185,N_14972);
and U19247 (N_19247,N_11829,N_12121);
and U19248 (N_19248,N_10683,N_11031);
nor U19249 (N_19249,N_12446,N_11956);
and U19250 (N_19250,N_13246,N_10585);
xnor U19251 (N_19251,N_13327,N_12251);
or U19252 (N_19252,N_10354,N_12164);
nor U19253 (N_19253,N_11513,N_10161);
or U19254 (N_19254,N_12722,N_10599);
or U19255 (N_19255,N_13045,N_12165);
or U19256 (N_19256,N_12434,N_12154);
nor U19257 (N_19257,N_14953,N_12977);
nand U19258 (N_19258,N_11839,N_11370);
nand U19259 (N_19259,N_12402,N_11603);
nor U19260 (N_19260,N_10356,N_13440);
and U19261 (N_19261,N_14544,N_10912);
nor U19262 (N_19262,N_12285,N_14643);
and U19263 (N_19263,N_13848,N_12248);
nor U19264 (N_19264,N_10797,N_11937);
nor U19265 (N_19265,N_10004,N_11855);
or U19266 (N_19266,N_14700,N_13359);
xor U19267 (N_19267,N_14509,N_10470);
or U19268 (N_19268,N_10805,N_11168);
and U19269 (N_19269,N_13780,N_10739);
or U19270 (N_19270,N_10112,N_13186);
xnor U19271 (N_19271,N_11212,N_10798);
and U19272 (N_19272,N_10550,N_14131);
xor U19273 (N_19273,N_12947,N_14279);
and U19274 (N_19274,N_11012,N_14348);
xor U19275 (N_19275,N_11198,N_11523);
and U19276 (N_19276,N_14560,N_13584);
and U19277 (N_19277,N_10127,N_12081);
nand U19278 (N_19278,N_14632,N_13413);
nor U19279 (N_19279,N_10338,N_12468);
xor U19280 (N_19280,N_10007,N_13895);
nor U19281 (N_19281,N_12532,N_14268);
nand U19282 (N_19282,N_14994,N_10840);
nand U19283 (N_19283,N_12748,N_14602);
or U19284 (N_19284,N_13332,N_11687);
nor U19285 (N_19285,N_14394,N_14719);
nor U19286 (N_19286,N_13313,N_14347);
or U19287 (N_19287,N_12834,N_12518);
or U19288 (N_19288,N_12128,N_14136);
nand U19289 (N_19289,N_10485,N_10646);
xnor U19290 (N_19290,N_11281,N_11141);
or U19291 (N_19291,N_10478,N_11891);
and U19292 (N_19292,N_14181,N_12846);
or U19293 (N_19293,N_10300,N_10073);
or U19294 (N_19294,N_13540,N_13352);
xnor U19295 (N_19295,N_10616,N_13025);
and U19296 (N_19296,N_11167,N_10345);
xor U19297 (N_19297,N_12160,N_14108);
and U19298 (N_19298,N_10469,N_11481);
and U19299 (N_19299,N_11789,N_14102);
or U19300 (N_19300,N_13025,N_12192);
or U19301 (N_19301,N_12426,N_12357);
or U19302 (N_19302,N_14758,N_11222);
nor U19303 (N_19303,N_14848,N_12485);
nand U19304 (N_19304,N_13000,N_10664);
nor U19305 (N_19305,N_14607,N_11398);
xnor U19306 (N_19306,N_12576,N_13734);
or U19307 (N_19307,N_14163,N_14919);
nor U19308 (N_19308,N_11979,N_14957);
nand U19309 (N_19309,N_14181,N_13914);
and U19310 (N_19310,N_10384,N_14924);
and U19311 (N_19311,N_13976,N_12584);
or U19312 (N_19312,N_14463,N_14475);
or U19313 (N_19313,N_11545,N_11865);
or U19314 (N_19314,N_13503,N_12194);
nand U19315 (N_19315,N_13014,N_14702);
or U19316 (N_19316,N_13482,N_14966);
and U19317 (N_19317,N_13078,N_14463);
and U19318 (N_19318,N_14184,N_13515);
and U19319 (N_19319,N_12030,N_12522);
or U19320 (N_19320,N_10029,N_10267);
or U19321 (N_19321,N_11089,N_14558);
nor U19322 (N_19322,N_13227,N_11255);
nand U19323 (N_19323,N_12028,N_13987);
xnor U19324 (N_19324,N_13432,N_10547);
or U19325 (N_19325,N_10196,N_10289);
or U19326 (N_19326,N_14026,N_10483);
and U19327 (N_19327,N_14610,N_13846);
and U19328 (N_19328,N_11539,N_14377);
and U19329 (N_19329,N_11256,N_12013);
nand U19330 (N_19330,N_13571,N_13548);
nor U19331 (N_19331,N_10150,N_10348);
and U19332 (N_19332,N_11403,N_11766);
nand U19333 (N_19333,N_11142,N_12160);
or U19334 (N_19334,N_12730,N_10266);
or U19335 (N_19335,N_12209,N_10059);
or U19336 (N_19336,N_12248,N_10861);
or U19337 (N_19337,N_11116,N_10003);
xnor U19338 (N_19338,N_13991,N_12764);
or U19339 (N_19339,N_10328,N_14438);
or U19340 (N_19340,N_11220,N_13492);
or U19341 (N_19341,N_10513,N_11950);
nor U19342 (N_19342,N_12938,N_12116);
or U19343 (N_19343,N_12283,N_11766);
nor U19344 (N_19344,N_10288,N_13559);
xor U19345 (N_19345,N_11029,N_12132);
or U19346 (N_19346,N_12032,N_12683);
xor U19347 (N_19347,N_11496,N_13610);
nand U19348 (N_19348,N_11466,N_11798);
xor U19349 (N_19349,N_13591,N_11870);
nor U19350 (N_19350,N_11609,N_14567);
or U19351 (N_19351,N_13743,N_11248);
nor U19352 (N_19352,N_13900,N_14914);
and U19353 (N_19353,N_14743,N_13729);
xnor U19354 (N_19354,N_10290,N_13472);
nand U19355 (N_19355,N_10903,N_12048);
nor U19356 (N_19356,N_10287,N_11085);
nand U19357 (N_19357,N_14620,N_10479);
and U19358 (N_19358,N_10498,N_13631);
nand U19359 (N_19359,N_11877,N_10831);
xor U19360 (N_19360,N_11764,N_11980);
nand U19361 (N_19361,N_13327,N_13746);
nand U19362 (N_19362,N_14682,N_14350);
nand U19363 (N_19363,N_10858,N_11037);
and U19364 (N_19364,N_10622,N_11485);
or U19365 (N_19365,N_13185,N_12676);
and U19366 (N_19366,N_10290,N_14062);
or U19367 (N_19367,N_11797,N_11393);
nor U19368 (N_19368,N_10370,N_14131);
xnor U19369 (N_19369,N_12915,N_10426);
nor U19370 (N_19370,N_10335,N_12347);
or U19371 (N_19371,N_12018,N_11693);
or U19372 (N_19372,N_10461,N_10363);
nor U19373 (N_19373,N_10187,N_11830);
and U19374 (N_19374,N_11288,N_12796);
xnor U19375 (N_19375,N_11021,N_13792);
nor U19376 (N_19376,N_11509,N_12226);
and U19377 (N_19377,N_13608,N_10026);
and U19378 (N_19378,N_10520,N_11807);
nor U19379 (N_19379,N_13445,N_14715);
xnor U19380 (N_19380,N_14226,N_14411);
nand U19381 (N_19381,N_10899,N_11335);
nand U19382 (N_19382,N_12713,N_13878);
nor U19383 (N_19383,N_14698,N_10885);
and U19384 (N_19384,N_11800,N_11760);
xor U19385 (N_19385,N_12606,N_10447);
or U19386 (N_19386,N_10438,N_11885);
nand U19387 (N_19387,N_14819,N_11417);
xor U19388 (N_19388,N_13037,N_14813);
xnor U19389 (N_19389,N_11030,N_14014);
and U19390 (N_19390,N_11877,N_11768);
nor U19391 (N_19391,N_13615,N_11574);
or U19392 (N_19392,N_12487,N_14565);
nand U19393 (N_19393,N_10794,N_10335);
or U19394 (N_19394,N_12453,N_13649);
nor U19395 (N_19395,N_11337,N_11808);
nor U19396 (N_19396,N_10801,N_10100);
or U19397 (N_19397,N_12689,N_14730);
or U19398 (N_19398,N_11805,N_13206);
xor U19399 (N_19399,N_10017,N_14774);
and U19400 (N_19400,N_12696,N_14460);
xnor U19401 (N_19401,N_14194,N_10463);
xnor U19402 (N_19402,N_11202,N_10369);
or U19403 (N_19403,N_14782,N_12342);
nand U19404 (N_19404,N_13228,N_10986);
or U19405 (N_19405,N_12265,N_10348);
or U19406 (N_19406,N_11783,N_10617);
xor U19407 (N_19407,N_14275,N_13426);
xor U19408 (N_19408,N_10843,N_14862);
nor U19409 (N_19409,N_12104,N_13553);
or U19410 (N_19410,N_11632,N_14482);
nand U19411 (N_19411,N_13747,N_12521);
nand U19412 (N_19412,N_10886,N_12134);
nand U19413 (N_19413,N_13817,N_11253);
xor U19414 (N_19414,N_10122,N_11160);
nand U19415 (N_19415,N_10049,N_11562);
nand U19416 (N_19416,N_11216,N_10114);
xor U19417 (N_19417,N_10073,N_12592);
xor U19418 (N_19418,N_11265,N_14988);
and U19419 (N_19419,N_13277,N_12373);
and U19420 (N_19420,N_13420,N_11893);
and U19421 (N_19421,N_12447,N_10657);
xor U19422 (N_19422,N_11535,N_10884);
or U19423 (N_19423,N_13153,N_10584);
xnor U19424 (N_19424,N_11349,N_10690);
nor U19425 (N_19425,N_13112,N_11317);
nand U19426 (N_19426,N_14599,N_11928);
xor U19427 (N_19427,N_11047,N_14810);
xor U19428 (N_19428,N_11434,N_10232);
and U19429 (N_19429,N_14361,N_14551);
or U19430 (N_19430,N_14191,N_12747);
xor U19431 (N_19431,N_10901,N_10091);
and U19432 (N_19432,N_14258,N_12458);
nor U19433 (N_19433,N_11454,N_14016);
xnor U19434 (N_19434,N_14533,N_13455);
and U19435 (N_19435,N_10191,N_12003);
and U19436 (N_19436,N_10677,N_11063);
and U19437 (N_19437,N_10874,N_13291);
and U19438 (N_19438,N_14423,N_11038);
nand U19439 (N_19439,N_12030,N_12989);
nand U19440 (N_19440,N_14888,N_12328);
nand U19441 (N_19441,N_10946,N_14781);
nand U19442 (N_19442,N_13200,N_13961);
xor U19443 (N_19443,N_12115,N_11131);
nor U19444 (N_19444,N_12220,N_13970);
xnor U19445 (N_19445,N_11867,N_11558);
and U19446 (N_19446,N_11291,N_11655);
nor U19447 (N_19447,N_13730,N_13462);
or U19448 (N_19448,N_13845,N_10839);
and U19449 (N_19449,N_13769,N_11300);
or U19450 (N_19450,N_10923,N_14575);
nand U19451 (N_19451,N_11557,N_14113);
xnor U19452 (N_19452,N_10999,N_12489);
nand U19453 (N_19453,N_14689,N_10849);
and U19454 (N_19454,N_10130,N_14614);
nand U19455 (N_19455,N_12309,N_13427);
xor U19456 (N_19456,N_12157,N_10159);
nand U19457 (N_19457,N_10232,N_10651);
nand U19458 (N_19458,N_10296,N_13337);
nor U19459 (N_19459,N_14603,N_14221);
and U19460 (N_19460,N_11353,N_10090);
xor U19461 (N_19461,N_12716,N_12458);
nand U19462 (N_19462,N_13672,N_11345);
or U19463 (N_19463,N_14411,N_10605);
nor U19464 (N_19464,N_10385,N_14354);
and U19465 (N_19465,N_11464,N_13720);
or U19466 (N_19466,N_13255,N_10884);
and U19467 (N_19467,N_10687,N_13178);
and U19468 (N_19468,N_13094,N_11914);
nand U19469 (N_19469,N_13116,N_12428);
and U19470 (N_19470,N_11022,N_13046);
and U19471 (N_19471,N_12768,N_13385);
nand U19472 (N_19472,N_11148,N_10084);
or U19473 (N_19473,N_10209,N_13087);
or U19474 (N_19474,N_12678,N_10745);
nor U19475 (N_19475,N_14464,N_12534);
or U19476 (N_19476,N_14805,N_14749);
nand U19477 (N_19477,N_12794,N_14354);
nor U19478 (N_19478,N_14925,N_13901);
and U19479 (N_19479,N_11681,N_10816);
and U19480 (N_19480,N_11771,N_10030);
nor U19481 (N_19481,N_11689,N_12049);
nor U19482 (N_19482,N_10497,N_14118);
nand U19483 (N_19483,N_10092,N_11545);
nor U19484 (N_19484,N_11872,N_14470);
nand U19485 (N_19485,N_14209,N_14927);
nor U19486 (N_19486,N_11221,N_10735);
or U19487 (N_19487,N_12983,N_10218);
and U19488 (N_19488,N_13477,N_14974);
or U19489 (N_19489,N_14742,N_10200);
and U19490 (N_19490,N_10199,N_13739);
nor U19491 (N_19491,N_12005,N_10769);
and U19492 (N_19492,N_14158,N_12824);
or U19493 (N_19493,N_12364,N_13083);
xnor U19494 (N_19494,N_10599,N_12897);
nor U19495 (N_19495,N_11278,N_14651);
nand U19496 (N_19496,N_14853,N_13014);
xnor U19497 (N_19497,N_13569,N_11716);
or U19498 (N_19498,N_14283,N_14562);
and U19499 (N_19499,N_12603,N_10013);
nand U19500 (N_19500,N_11129,N_10488);
xor U19501 (N_19501,N_14939,N_13988);
or U19502 (N_19502,N_12704,N_14215);
nor U19503 (N_19503,N_14241,N_10380);
and U19504 (N_19504,N_14049,N_10197);
or U19505 (N_19505,N_10163,N_11152);
nand U19506 (N_19506,N_10939,N_13612);
xor U19507 (N_19507,N_14754,N_12803);
or U19508 (N_19508,N_14199,N_14999);
xor U19509 (N_19509,N_14717,N_13648);
nor U19510 (N_19510,N_11882,N_11501);
nor U19511 (N_19511,N_10947,N_11324);
and U19512 (N_19512,N_10325,N_14036);
xnor U19513 (N_19513,N_12127,N_11081);
xnor U19514 (N_19514,N_12691,N_12787);
nand U19515 (N_19515,N_14764,N_10373);
nand U19516 (N_19516,N_13010,N_14126);
or U19517 (N_19517,N_12781,N_12357);
nand U19518 (N_19518,N_12320,N_13405);
nor U19519 (N_19519,N_11709,N_14000);
or U19520 (N_19520,N_12813,N_11886);
xnor U19521 (N_19521,N_10496,N_10601);
nand U19522 (N_19522,N_10151,N_13915);
nand U19523 (N_19523,N_13262,N_12935);
or U19524 (N_19524,N_14228,N_11541);
nand U19525 (N_19525,N_11819,N_12869);
nand U19526 (N_19526,N_14037,N_10234);
nor U19527 (N_19527,N_14119,N_12967);
or U19528 (N_19528,N_12446,N_14739);
xnor U19529 (N_19529,N_11702,N_10531);
nand U19530 (N_19530,N_14566,N_13378);
nand U19531 (N_19531,N_11148,N_14489);
xnor U19532 (N_19532,N_11891,N_14739);
xnor U19533 (N_19533,N_12047,N_10708);
and U19534 (N_19534,N_13444,N_13104);
or U19535 (N_19535,N_14232,N_12796);
and U19536 (N_19536,N_11451,N_14390);
nand U19537 (N_19537,N_13689,N_12730);
and U19538 (N_19538,N_13221,N_10329);
nor U19539 (N_19539,N_12983,N_14195);
or U19540 (N_19540,N_11553,N_13945);
xnor U19541 (N_19541,N_12326,N_10468);
nand U19542 (N_19542,N_10211,N_12695);
nand U19543 (N_19543,N_12705,N_12736);
or U19544 (N_19544,N_12071,N_10746);
or U19545 (N_19545,N_11360,N_13041);
and U19546 (N_19546,N_12830,N_10079);
nand U19547 (N_19547,N_13741,N_11461);
nand U19548 (N_19548,N_14325,N_13820);
nand U19549 (N_19549,N_13079,N_12185);
nor U19550 (N_19550,N_14749,N_14763);
or U19551 (N_19551,N_14973,N_14103);
or U19552 (N_19552,N_12483,N_12252);
xnor U19553 (N_19553,N_10041,N_11295);
xor U19554 (N_19554,N_10947,N_13443);
or U19555 (N_19555,N_13602,N_11897);
and U19556 (N_19556,N_14888,N_10535);
nand U19557 (N_19557,N_10223,N_10198);
or U19558 (N_19558,N_10743,N_11445);
xor U19559 (N_19559,N_14433,N_14153);
nor U19560 (N_19560,N_11672,N_12445);
xnor U19561 (N_19561,N_12343,N_10774);
or U19562 (N_19562,N_10342,N_14635);
xnor U19563 (N_19563,N_10231,N_14460);
and U19564 (N_19564,N_13737,N_11512);
or U19565 (N_19565,N_10022,N_13785);
nor U19566 (N_19566,N_12799,N_12324);
xor U19567 (N_19567,N_12131,N_13397);
nand U19568 (N_19568,N_11493,N_14980);
xor U19569 (N_19569,N_13372,N_14764);
xor U19570 (N_19570,N_11849,N_10260);
or U19571 (N_19571,N_13375,N_10551);
nand U19572 (N_19572,N_13589,N_11253);
or U19573 (N_19573,N_14798,N_12557);
nand U19574 (N_19574,N_14683,N_11013);
and U19575 (N_19575,N_14963,N_10570);
nor U19576 (N_19576,N_14880,N_13404);
or U19577 (N_19577,N_13714,N_13297);
nor U19578 (N_19578,N_11976,N_11630);
xnor U19579 (N_19579,N_12003,N_14503);
and U19580 (N_19580,N_14969,N_14872);
nand U19581 (N_19581,N_10420,N_11511);
nor U19582 (N_19582,N_10123,N_13278);
nand U19583 (N_19583,N_10780,N_13936);
or U19584 (N_19584,N_11459,N_10197);
nor U19585 (N_19585,N_11929,N_10405);
xor U19586 (N_19586,N_14290,N_14713);
or U19587 (N_19587,N_12699,N_13642);
and U19588 (N_19588,N_14248,N_13652);
nor U19589 (N_19589,N_10874,N_14864);
or U19590 (N_19590,N_13506,N_11787);
xnor U19591 (N_19591,N_13974,N_10173);
and U19592 (N_19592,N_10312,N_11613);
and U19593 (N_19593,N_10694,N_14946);
and U19594 (N_19594,N_13020,N_14672);
nand U19595 (N_19595,N_10302,N_12863);
and U19596 (N_19596,N_12010,N_13493);
xnor U19597 (N_19597,N_12804,N_14852);
or U19598 (N_19598,N_12133,N_11599);
xor U19599 (N_19599,N_12974,N_10788);
nor U19600 (N_19600,N_13177,N_13962);
xnor U19601 (N_19601,N_10315,N_13714);
or U19602 (N_19602,N_11385,N_13890);
nand U19603 (N_19603,N_14654,N_14374);
and U19604 (N_19604,N_10243,N_14176);
or U19605 (N_19605,N_11517,N_14528);
nor U19606 (N_19606,N_14684,N_12802);
and U19607 (N_19607,N_13442,N_13990);
or U19608 (N_19608,N_10793,N_13661);
and U19609 (N_19609,N_13997,N_12538);
nor U19610 (N_19610,N_10081,N_11680);
and U19611 (N_19611,N_14006,N_13913);
xor U19612 (N_19612,N_14388,N_13952);
and U19613 (N_19613,N_12526,N_14981);
nand U19614 (N_19614,N_10924,N_13959);
or U19615 (N_19615,N_14560,N_12357);
nor U19616 (N_19616,N_12047,N_14967);
nor U19617 (N_19617,N_13980,N_12256);
and U19618 (N_19618,N_10026,N_13531);
nand U19619 (N_19619,N_14779,N_12190);
nand U19620 (N_19620,N_14137,N_13353);
or U19621 (N_19621,N_13872,N_11911);
or U19622 (N_19622,N_10118,N_14569);
and U19623 (N_19623,N_14815,N_13201);
and U19624 (N_19624,N_13102,N_14041);
xor U19625 (N_19625,N_10476,N_13008);
xor U19626 (N_19626,N_14258,N_12656);
xor U19627 (N_19627,N_12668,N_11244);
nand U19628 (N_19628,N_12648,N_12169);
xnor U19629 (N_19629,N_10929,N_10207);
and U19630 (N_19630,N_13893,N_12510);
xnor U19631 (N_19631,N_10689,N_10402);
xnor U19632 (N_19632,N_13898,N_11233);
and U19633 (N_19633,N_13704,N_12364);
nand U19634 (N_19634,N_13597,N_10577);
nor U19635 (N_19635,N_14704,N_10906);
or U19636 (N_19636,N_10410,N_13177);
nand U19637 (N_19637,N_10638,N_14735);
nor U19638 (N_19638,N_14500,N_14769);
xnor U19639 (N_19639,N_11155,N_13622);
and U19640 (N_19640,N_11363,N_13848);
nor U19641 (N_19641,N_14075,N_10348);
or U19642 (N_19642,N_14139,N_13434);
xor U19643 (N_19643,N_13457,N_13952);
nor U19644 (N_19644,N_13610,N_12396);
and U19645 (N_19645,N_13680,N_13326);
nand U19646 (N_19646,N_10940,N_10232);
xnor U19647 (N_19647,N_11941,N_13738);
xnor U19648 (N_19648,N_14532,N_14340);
or U19649 (N_19649,N_14208,N_12883);
xnor U19650 (N_19650,N_11619,N_10911);
nor U19651 (N_19651,N_13746,N_12326);
xnor U19652 (N_19652,N_12323,N_10286);
nor U19653 (N_19653,N_11064,N_13279);
and U19654 (N_19654,N_11068,N_13567);
xnor U19655 (N_19655,N_12518,N_14916);
nor U19656 (N_19656,N_12050,N_14595);
nor U19657 (N_19657,N_13478,N_13644);
nand U19658 (N_19658,N_14846,N_10434);
and U19659 (N_19659,N_10574,N_13635);
nor U19660 (N_19660,N_14743,N_10826);
xor U19661 (N_19661,N_11277,N_12455);
and U19662 (N_19662,N_14197,N_10444);
and U19663 (N_19663,N_10260,N_10311);
nand U19664 (N_19664,N_13103,N_13506);
xnor U19665 (N_19665,N_13162,N_11359);
xor U19666 (N_19666,N_14662,N_11539);
or U19667 (N_19667,N_14963,N_10708);
nand U19668 (N_19668,N_10572,N_10445);
nor U19669 (N_19669,N_13920,N_10692);
and U19670 (N_19670,N_14468,N_11949);
xor U19671 (N_19671,N_14102,N_14552);
nor U19672 (N_19672,N_12446,N_13032);
or U19673 (N_19673,N_13667,N_14449);
or U19674 (N_19674,N_13717,N_11286);
and U19675 (N_19675,N_11635,N_13443);
nor U19676 (N_19676,N_12985,N_14004);
and U19677 (N_19677,N_11671,N_11049);
or U19678 (N_19678,N_13743,N_11282);
or U19679 (N_19679,N_13880,N_12541);
nand U19680 (N_19680,N_14111,N_12519);
nor U19681 (N_19681,N_14517,N_10841);
nand U19682 (N_19682,N_13720,N_11480);
xor U19683 (N_19683,N_14483,N_13153);
nor U19684 (N_19684,N_10182,N_13750);
and U19685 (N_19685,N_10290,N_14593);
nor U19686 (N_19686,N_12609,N_14401);
nor U19687 (N_19687,N_13783,N_12974);
xnor U19688 (N_19688,N_13113,N_12457);
or U19689 (N_19689,N_13558,N_11357);
nand U19690 (N_19690,N_10199,N_11463);
nand U19691 (N_19691,N_10768,N_11879);
nor U19692 (N_19692,N_11999,N_11083);
and U19693 (N_19693,N_11986,N_14778);
xor U19694 (N_19694,N_11929,N_14610);
and U19695 (N_19695,N_13760,N_12469);
and U19696 (N_19696,N_13073,N_13713);
nor U19697 (N_19697,N_12508,N_14025);
nor U19698 (N_19698,N_11453,N_14233);
or U19699 (N_19699,N_14238,N_12158);
xor U19700 (N_19700,N_14490,N_14454);
xnor U19701 (N_19701,N_10164,N_10927);
and U19702 (N_19702,N_12340,N_11031);
xor U19703 (N_19703,N_13956,N_11113);
nor U19704 (N_19704,N_11730,N_13655);
nand U19705 (N_19705,N_12908,N_13143);
and U19706 (N_19706,N_10599,N_12555);
nor U19707 (N_19707,N_12664,N_13874);
xnor U19708 (N_19708,N_14482,N_11049);
and U19709 (N_19709,N_11535,N_13538);
nor U19710 (N_19710,N_13846,N_11668);
or U19711 (N_19711,N_12038,N_12452);
xor U19712 (N_19712,N_12603,N_13757);
and U19713 (N_19713,N_10507,N_14860);
nand U19714 (N_19714,N_10288,N_12973);
or U19715 (N_19715,N_11220,N_12111);
or U19716 (N_19716,N_13077,N_14208);
nand U19717 (N_19717,N_10253,N_11709);
xnor U19718 (N_19718,N_10496,N_13884);
or U19719 (N_19719,N_14404,N_10205);
nand U19720 (N_19720,N_10459,N_11646);
xor U19721 (N_19721,N_14208,N_14956);
nor U19722 (N_19722,N_13505,N_14653);
xnor U19723 (N_19723,N_14868,N_12114);
or U19724 (N_19724,N_10220,N_12026);
xnor U19725 (N_19725,N_11329,N_10993);
or U19726 (N_19726,N_12407,N_10537);
nand U19727 (N_19727,N_11344,N_11706);
xnor U19728 (N_19728,N_14200,N_11157);
and U19729 (N_19729,N_10292,N_13259);
nand U19730 (N_19730,N_11290,N_14099);
or U19731 (N_19731,N_12502,N_13533);
nand U19732 (N_19732,N_14853,N_13042);
or U19733 (N_19733,N_11056,N_10508);
or U19734 (N_19734,N_13924,N_14728);
nand U19735 (N_19735,N_12060,N_14060);
nor U19736 (N_19736,N_10808,N_11553);
nand U19737 (N_19737,N_10507,N_12486);
nor U19738 (N_19738,N_10683,N_10098);
nand U19739 (N_19739,N_14649,N_14585);
nor U19740 (N_19740,N_13335,N_10141);
and U19741 (N_19741,N_13398,N_10388);
or U19742 (N_19742,N_13358,N_14811);
nor U19743 (N_19743,N_14695,N_14885);
and U19744 (N_19744,N_10750,N_14470);
nor U19745 (N_19745,N_10818,N_10319);
nand U19746 (N_19746,N_10989,N_11557);
and U19747 (N_19747,N_14199,N_14013);
xor U19748 (N_19748,N_10730,N_14177);
nor U19749 (N_19749,N_12923,N_14275);
and U19750 (N_19750,N_13367,N_12281);
and U19751 (N_19751,N_10031,N_12020);
and U19752 (N_19752,N_13938,N_12157);
nand U19753 (N_19753,N_11123,N_12600);
or U19754 (N_19754,N_11346,N_13217);
nor U19755 (N_19755,N_10919,N_10384);
and U19756 (N_19756,N_11665,N_11525);
xnor U19757 (N_19757,N_12956,N_12029);
xor U19758 (N_19758,N_11006,N_13497);
nor U19759 (N_19759,N_14010,N_14613);
or U19760 (N_19760,N_12347,N_10108);
nor U19761 (N_19761,N_13337,N_13366);
and U19762 (N_19762,N_12140,N_11964);
nor U19763 (N_19763,N_10738,N_13606);
or U19764 (N_19764,N_12130,N_11037);
or U19765 (N_19765,N_13554,N_10830);
and U19766 (N_19766,N_14468,N_11478);
nand U19767 (N_19767,N_11770,N_10715);
or U19768 (N_19768,N_12056,N_14321);
xnor U19769 (N_19769,N_13151,N_12758);
or U19770 (N_19770,N_12599,N_14630);
nand U19771 (N_19771,N_10684,N_14670);
or U19772 (N_19772,N_14605,N_14016);
or U19773 (N_19773,N_13626,N_12942);
nand U19774 (N_19774,N_14427,N_11302);
nor U19775 (N_19775,N_14092,N_10931);
nand U19776 (N_19776,N_13427,N_13908);
xor U19777 (N_19777,N_11188,N_11995);
and U19778 (N_19778,N_11630,N_13627);
nand U19779 (N_19779,N_14185,N_14909);
or U19780 (N_19780,N_11888,N_14372);
xor U19781 (N_19781,N_12678,N_13695);
or U19782 (N_19782,N_13756,N_12467);
xnor U19783 (N_19783,N_10615,N_14745);
xnor U19784 (N_19784,N_13781,N_14969);
nor U19785 (N_19785,N_11801,N_12321);
and U19786 (N_19786,N_10170,N_13736);
and U19787 (N_19787,N_12425,N_11373);
nor U19788 (N_19788,N_13583,N_13769);
xor U19789 (N_19789,N_13966,N_11388);
xor U19790 (N_19790,N_12766,N_10658);
or U19791 (N_19791,N_14331,N_10593);
xnor U19792 (N_19792,N_11806,N_13375);
nand U19793 (N_19793,N_13214,N_12322);
and U19794 (N_19794,N_14213,N_13270);
or U19795 (N_19795,N_13607,N_10002);
xor U19796 (N_19796,N_12975,N_10058);
xor U19797 (N_19797,N_12045,N_10355);
nor U19798 (N_19798,N_11468,N_10650);
nor U19799 (N_19799,N_14620,N_11989);
nor U19800 (N_19800,N_13690,N_11290);
xnor U19801 (N_19801,N_10112,N_12352);
xor U19802 (N_19802,N_14014,N_10383);
nor U19803 (N_19803,N_12595,N_11816);
nor U19804 (N_19804,N_10772,N_13267);
nor U19805 (N_19805,N_12754,N_10783);
or U19806 (N_19806,N_11086,N_13250);
or U19807 (N_19807,N_14577,N_13823);
and U19808 (N_19808,N_14058,N_13575);
xor U19809 (N_19809,N_14779,N_12889);
or U19810 (N_19810,N_13215,N_11635);
nand U19811 (N_19811,N_13970,N_14068);
and U19812 (N_19812,N_12412,N_14644);
or U19813 (N_19813,N_10358,N_14535);
nand U19814 (N_19814,N_13187,N_13820);
xnor U19815 (N_19815,N_12871,N_12228);
or U19816 (N_19816,N_12372,N_14616);
nor U19817 (N_19817,N_14512,N_14681);
or U19818 (N_19818,N_11612,N_14233);
and U19819 (N_19819,N_12623,N_12317);
nand U19820 (N_19820,N_14153,N_10549);
or U19821 (N_19821,N_10714,N_13037);
xnor U19822 (N_19822,N_11891,N_10374);
nand U19823 (N_19823,N_10099,N_11758);
nor U19824 (N_19824,N_11866,N_13933);
or U19825 (N_19825,N_14026,N_12371);
nand U19826 (N_19826,N_10956,N_12449);
xnor U19827 (N_19827,N_12604,N_10661);
nand U19828 (N_19828,N_14873,N_13278);
or U19829 (N_19829,N_11347,N_12927);
xnor U19830 (N_19830,N_14514,N_11248);
or U19831 (N_19831,N_11112,N_13516);
and U19832 (N_19832,N_13806,N_14567);
or U19833 (N_19833,N_12807,N_12157);
and U19834 (N_19834,N_12037,N_12905);
nor U19835 (N_19835,N_14661,N_12032);
nand U19836 (N_19836,N_11928,N_10751);
nor U19837 (N_19837,N_12361,N_10960);
xor U19838 (N_19838,N_11228,N_13152);
xor U19839 (N_19839,N_13747,N_12231);
xnor U19840 (N_19840,N_11857,N_12437);
or U19841 (N_19841,N_13973,N_11259);
and U19842 (N_19842,N_11946,N_14224);
and U19843 (N_19843,N_10463,N_12243);
nor U19844 (N_19844,N_12680,N_13939);
or U19845 (N_19845,N_14840,N_10064);
or U19846 (N_19846,N_14570,N_14686);
xor U19847 (N_19847,N_10060,N_14927);
nor U19848 (N_19848,N_12374,N_13414);
or U19849 (N_19849,N_11868,N_14975);
nor U19850 (N_19850,N_10574,N_12003);
and U19851 (N_19851,N_14940,N_11010);
or U19852 (N_19852,N_12994,N_10946);
nand U19853 (N_19853,N_12001,N_11325);
nor U19854 (N_19854,N_14426,N_10601);
or U19855 (N_19855,N_14931,N_12361);
nand U19856 (N_19856,N_11267,N_12195);
nand U19857 (N_19857,N_12082,N_12250);
or U19858 (N_19858,N_14141,N_10858);
or U19859 (N_19859,N_13825,N_13896);
nand U19860 (N_19860,N_13660,N_14915);
xnor U19861 (N_19861,N_11093,N_11278);
and U19862 (N_19862,N_13795,N_11812);
nand U19863 (N_19863,N_11779,N_10449);
nor U19864 (N_19864,N_12037,N_14608);
nor U19865 (N_19865,N_14269,N_10821);
or U19866 (N_19866,N_10377,N_10401);
and U19867 (N_19867,N_11018,N_14663);
and U19868 (N_19868,N_13345,N_14251);
nor U19869 (N_19869,N_14182,N_14177);
and U19870 (N_19870,N_14318,N_12138);
nand U19871 (N_19871,N_11983,N_10554);
nor U19872 (N_19872,N_14847,N_11414);
xnor U19873 (N_19873,N_11085,N_11803);
and U19874 (N_19874,N_10429,N_10613);
or U19875 (N_19875,N_14629,N_13175);
or U19876 (N_19876,N_12776,N_12254);
nor U19877 (N_19877,N_14572,N_11070);
nor U19878 (N_19878,N_11412,N_13843);
xor U19879 (N_19879,N_11771,N_13188);
or U19880 (N_19880,N_13464,N_13661);
or U19881 (N_19881,N_14503,N_11308);
or U19882 (N_19882,N_11020,N_10614);
nand U19883 (N_19883,N_12197,N_14869);
and U19884 (N_19884,N_14989,N_13704);
nand U19885 (N_19885,N_11487,N_14811);
nand U19886 (N_19886,N_13019,N_11508);
xor U19887 (N_19887,N_14158,N_14114);
or U19888 (N_19888,N_13749,N_10072);
nor U19889 (N_19889,N_10109,N_10932);
and U19890 (N_19890,N_13006,N_12006);
nor U19891 (N_19891,N_10367,N_10413);
nand U19892 (N_19892,N_14699,N_14690);
nor U19893 (N_19893,N_10240,N_10599);
nand U19894 (N_19894,N_11249,N_10915);
or U19895 (N_19895,N_13625,N_10485);
or U19896 (N_19896,N_14693,N_11230);
xnor U19897 (N_19897,N_14811,N_14720);
nor U19898 (N_19898,N_12094,N_10429);
xor U19899 (N_19899,N_11387,N_10074);
or U19900 (N_19900,N_14226,N_13830);
xor U19901 (N_19901,N_10495,N_14220);
or U19902 (N_19902,N_14809,N_13390);
nor U19903 (N_19903,N_11667,N_13283);
or U19904 (N_19904,N_11774,N_12813);
nand U19905 (N_19905,N_11434,N_10405);
nand U19906 (N_19906,N_13713,N_14341);
and U19907 (N_19907,N_11638,N_13014);
nand U19908 (N_19908,N_10689,N_13055);
and U19909 (N_19909,N_14847,N_13061);
nor U19910 (N_19910,N_11404,N_13015);
or U19911 (N_19911,N_14598,N_10940);
and U19912 (N_19912,N_11839,N_13181);
and U19913 (N_19913,N_11603,N_14003);
xnor U19914 (N_19914,N_14490,N_13947);
or U19915 (N_19915,N_11886,N_11409);
xor U19916 (N_19916,N_11465,N_12391);
xor U19917 (N_19917,N_10118,N_13414);
or U19918 (N_19918,N_11547,N_12861);
and U19919 (N_19919,N_13894,N_10219);
xor U19920 (N_19920,N_11277,N_11555);
and U19921 (N_19921,N_11482,N_12880);
xnor U19922 (N_19922,N_14438,N_14445);
and U19923 (N_19923,N_12860,N_11121);
or U19924 (N_19924,N_10579,N_13102);
or U19925 (N_19925,N_12415,N_11265);
nand U19926 (N_19926,N_12068,N_14114);
and U19927 (N_19927,N_14066,N_13665);
nor U19928 (N_19928,N_14419,N_13341);
nand U19929 (N_19929,N_14230,N_14877);
nor U19930 (N_19930,N_10394,N_11898);
nand U19931 (N_19931,N_12893,N_14825);
or U19932 (N_19932,N_10873,N_14311);
xor U19933 (N_19933,N_10626,N_11808);
nand U19934 (N_19934,N_12041,N_10760);
or U19935 (N_19935,N_11131,N_12843);
nand U19936 (N_19936,N_10095,N_13224);
or U19937 (N_19937,N_14039,N_13618);
nand U19938 (N_19938,N_14351,N_10820);
nor U19939 (N_19939,N_13969,N_11785);
xor U19940 (N_19940,N_14487,N_12576);
or U19941 (N_19941,N_11883,N_12664);
nor U19942 (N_19942,N_12383,N_12695);
and U19943 (N_19943,N_10445,N_12618);
xor U19944 (N_19944,N_14924,N_14122);
nand U19945 (N_19945,N_12881,N_13466);
or U19946 (N_19946,N_14889,N_11874);
xnor U19947 (N_19947,N_12667,N_11437);
or U19948 (N_19948,N_11635,N_10593);
or U19949 (N_19949,N_12807,N_11337);
nand U19950 (N_19950,N_14274,N_12217);
nand U19951 (N_19951,N_10175,N_10002);
or U19952 (N_19952,N_10965,N_12388);
nor U19953 (N_19953,N_12260,N_11653);
or U19954 (N_19954,N_14662,N_12775);
nor U19955 (N_19955,N_14925,N_12983);
nand U19956 (N_19956,N_14202,N_13290);
and U19957 (N_19957,N_13300,N_11744);
xnor U19958 (N_19958,N_14557,N_11045);
and U19959 (N_19959,N_12431,N_10543);
nor U19960 (N_19960,N_13854,N_13194);
nand U19961 (N_19961,N_14523,N_12753);
xnor U19962 (N_19962,N_11663,N_13553);
nand U19963 (N_19963,N_11335,N_12844);
nand U19964 (N_19964,N_14925,N_12397);
and U19965 (N_19965,N_11430,N_10390);
and U19966 (N_19966,N_10030,N_14198);
or U19967 (N_19967,N_11714,N_10096);
nor U19968 (N_19968,N_12739,N_10694);
xnor U19969 (N_19969,N_12591,N_11281);
and U19970 (N_19970,N_14805,N_13527);
or U19971 (N_19971,N_14264,N_10810);
xor U19972 (N_19972,N_13531,N_10001);
xor U19973 (N_19973,N_11613,N_13212);
nand U19974 (N_19974,N_14008,N_13345);
nand U19975 (N_19975,N_10433,N_13844);
or U19976 (N_19976,N_14477,N_13729);
nand U19977 (N_19977,N_10731,N_12993);
nand U19978 (N_19978,N_14307,N_10225);
nand U19979 (N_19979,N_13978,N_11934);
nand U19980 (N_19980,N_12830,N_14046);
xor U19981 (N_19981,N_10703,N_13787);
or U19982 (N_19982,N_13721,N_13326);
nor U19983 (N_19983,N_13469,N_12046);
xnor U19984 (N_19984,N_12041,N_13438);
and U19985 (N_19985,N_11703,N_12824);
nand U19986 (N_19986,N_14724,N_11586);
or U19987 (N_19987,N_10925,N_14427);
or U19988 (N_19988,N_11521,N_10118);
and U19989 (N_19989,N_13257,N_11329);
xnor U19990 (N_19990,N_10149,N_10136);
nand U19991 (N_19991,N_13450,N_14896);
and U19992 (N_19992,N_12782,N_14229);
xnor U19993 (N_19993,N_10588,N_10026);
nand U19994 (N_19994,N_14230,N_12629);
nand U19995 (N_19995,N_14924,N_13792);
and U19996 (N_19996,N_12174,N_12497);
and U19997 (N_19997,N_12426,N_11934);
nor U19998 (N_19998,N_13167,N_10813);
nand U19999 (N_19999,N_12668,N_10432);
nand U20000 (N_20000,N_18376,N_16826);
nor U20001 (N_20001,N_18068,N_15770);
or U20002 (N_20002,N_18796,N_17626);
and U20003 (N_20003,N_17365,N_19004);
nand U20004 (N_20004,N_19679,N_19391);
nand U20005 (N_20005,N_17456,N_17855);
or U20006 (N_20006,N_18942,N_16140);
and U20007 (N_20007,N_16263,N_16170);
xor U20008 (N_20008,N_19827,N_15386);
nor U20009 (N_20009,N_18529,N_15750);
and U20010 (N_20010,N_17722,N_16278);
nand U20011 (N_20011,N_18270,N_17991);
and U20012 (N_20012,N_16935,N_18253);
xnor U20013 (N_20013,N_19543,N_19330);
nand U20014 (N_20014,N_19488,N_15331);
nor U20015 (N_20015,N_19582,N_16754);
nand U20016 (N_20016,N_16657,N_19451);
nor U20017 (N_20017,N_19584,N_15080);
nand U20018 (N_20018,N_18455,N_19599);
xnor U20019 (N_20019,N_15335,N_19625);
or U20020 (N_20020,N_15121,N_15940);
and U20021 (N_20021,N_16542,N_15767);
nand U20022 (N_20022,N_19471,N_18204);
or U20023 (N_20023,N_16078,N_19510);
nand U20024 (N_20024,N_16898,N_19424);
nand U20025 (N_20025,N_17426,N_18478);
nor U20026 (N_20026,N_17845,N_18386);
and U20027 (N_20027,N_19672,N_16001);
nand U20028 (N_20028,N_16839,N_16763);
or U20029 (N_20029,N_16403,N_17778);
nor U20030 (N_20030,N_15971,N_19895);
or U20031 (N_20031,N_18557,N_18312);
or U20032 (N_20032,N_19955,N_19900);
nor U20033 (N_20033,N_18626,N_19881);
xor U20034 (N_20034,N_17966,N_19917);
or U20035 (N_20035,N_15402,N_19892);
nand U20036 (N_20036,N_19311,N_15865);
xnor U20037 (N_20037,N_19089,N_17749);
nand U20038 (N_20038,N_17977,N_17262);
nor U20039 (N_20039,N_17844,N_19341);
nor U20040 (N_20040,N_18090,N_15455);
and U20041 (N_20041,N_19415,N_16332);
nor U20042 (N_20042,N_19213,N_16107);
xor U20043 (N_20043,N_19052,N_19739);
and U20044 (N_20044,N_18224,N_18170);
xor U20045 (N_20045,N_18385,N_16479);
nand U20046 (N_20046,N_15195,N_18742);
nor U20047 (N_20047,N_17980,N_17022);
nand U20048 (N_20048,N_18433,N_18681);
nor U20049 (N_20049,N_18842,N_15276);
nor U20050 (N_20050,N_17942,N_16847);
nor U20051 (N_20051,N_17227,N_15790);
or U20052 (N_20052,N_19244,N_15274);
nor U20053 (N_20053,N_18106,N_15120);
and U20054 (N_20054,N_19877,N_17318);
or U20055 (N_20055,N_18486,N_15248);
nor U20056 (N_20056,N_15685,N_18899);
nand U20057 (N_20057,N_15107,N_15293);
and U20058 (N_20058,N_16094,N_16882);
and U20059 (N_20059,N_15078,N_18728);
nor U20060 (N_20060,N_17806,N_16300);
or U20061 (N_20061,N_17092,N_17981);
nor U20062 (N_20062,N_15132,N_15892);
or U20063 (N_20063,N_15809,N_18944);
xor U20064 (N_20064,N_19318,N_15821);
or U20065 (N_20065,N_15098,N_18867);
and U20066 (N_20066,N_19541,N_17536);
nor U20067 (N_20067,N_15600,N_15085);
or U20068 (N_20068,N_19194,N_19624);
or U20069 (N_20069,N_15145,N_16943);
xnor U20070 (N_20070,N_16761,N_15167);
or U20071 (N_20071,N_18780,N_17978);
and U20072 (N_20072,N_19355,N_18804);
and U20073 (N_20073,N_16036,N_16640);
xor U20074 (N_20074,N_18731,N_17382);
nand U20075 (N_20075,N_16687,N_16212);
nor U20076 (N_20076,N_17246,N_16370);
xnor U20077 (N_20077,N_19487,N_16553);
xnor U20078 (N_20078,N_17742,N_18398);
xnor U20079 (N_20079,N_19644,N_18847);
or U20080 (N_20080,N_15029,N_16123);
nand U20081 (N_20081,N_16106,N_17415);
nand U20082 (N_20082,N_19239,N_16686);
or U20083 (N_20083,N_16684,N_19162);
nor U20084 (N_20084,N_17355,N_16905);
nor U20085 (N_20085,N_15568,N_15820);
or U20086 (N_20086,N_15933,N_19240);
nor U20087 (N_20087,N_19883,N_15642);
nand U20088 (N_20088,N_17903,N_18801);
or U20089 (N_20089,N_15227,N_16270);
nand U20090 (N_20090,N_16373,N_17555);
nand U20091 (N_20091,N_18313,N_19389);
nand U20092 (N_20092,N_16115,N_17795);
or U20093 (N_20093,N_16303,N_15044);
and U20094 (N_20094,N_16196,N_18508);
nor U20095 (N_20095,N_16872,N_19496);
xnor U20096 (N_20096,N_18881,N_17771);
xnor U20097 (N_20097,N_17691,N_19158);
or U20098 (N_20098,N_18908,N_16246);
or U20099 (N_20099,N_16353,N_16803);
or U20100 (N_20100,N_17234,N_18069);
and U20101 (N_20101,N_18636,N_15288);
nand U20102 (N_20102,N_19852,N_17420);
or U20103 (N_20103,N_18029,N_15793);
or U20104 (N_20104,N_16151,N_17604);
xnor U20105 (N_20105,N_19022,N_19091);
nand U20106 (N_20106,N_17427,N_19690);
nand U20107 (N_20107,N_18672,N_19208);
or U20108 (N_20108,N_17994,N_15887);
or U20109 (N_20109,N_18448,N_16772);
nand U20110 (N_20110,N_15840,N_15135);
or U20111 (N_20111,N_17501,N_18549);
and U20112 (N_20112,N_15058,N_18920);
nor U20113 (N_20113,N_18164,N_18097);
or U20114 (N_20114,N_17949,N_19726);
nand U20115 (N_20115,N_15799,N_19112);
or U20116 (N_20116,N_17702,N_17263);
or U20117 (N_20117,N_15075,N_16306);
and U20118 (N_20118,N_15670,N_15502);
and U20119 (N_20119,N_19676,N_19361);
and U20120 (N_20120,N_15748,N_16105);
nor U20121 (N_20121,N_18434,N_16846);
nand U20122 (N_20122,N_16389,N_15077);
xor U20123 (N_20123,N_16626,N_18992);
nand U20124 (N_20124,N_18355,N_19390);
nand U20125 (N_20125,N_16878,N_15571);
or U20126 (N_20126,N_16526,N_18275);
and U20127 (N_20127,N_19594,N_19097);
or U20128 (N_20128,N_15728,N_17134);
xor U20129 (N_20129,N_17886,N_15932);
and U20130 (N_20130,N_17574,N_18473);
or U20131 (N_20131,N_16157,N_19869);
and U20132 (N_20132,N_15751,N_19713);
xnor U20133 (N_20133,N_18160,N_18382);
or U20134 (N_20134,N_17049,N_17221);
and U20135 (N_20135,N_18790,N_19765);
xnor U20136 (N_20136,N_16964,N_18991);
xor U20137 (N_20137,N_19916,N_15005);
nor U20138 (N_20138,N_19971,N_15904);
or U20139 (N_20139,N_17010,N_19670);
xor U20140 (N_20140,N_18218,N_18730);
and U20141 (N_20141,N_17218,N_15146);
or U20142 (N_20142,N_19267,N_16215);
and U20143 (N_20143,N_15023,N_15119);
nor U20144 (N_20144,N_16746,N_16741);
or U20145 (N_20145,N_18807,N_17087);
or U20146 (N_20146,N_19100,N_18083);
and U20147 (N_20147,N_17492,N_19150);
xor U20148 (N_20148,N_19121,N_15757);
and U20149 (N_20149,N_17310,N_17960);
nand U20150 (N_20150,N_17736,N_18359);
and U20151 (N_20151,N_16587,N_18406);
and U20152 (N_20152,N_18271,N_19538);
nand U20153 (N_20153,N_18716,N_18241);
xor U20154 (N_20154,N_18436,N_19693);
nand U20155 (N_20155,N_18460,N_15429);
nor U20156 (N_20156,N_16261,N_15312);
nor U20157 (N_20157,N_19411,N_18775);
or U20158 (N_20158,N_18323,N_19157);
xor U20159 (N_20159,N_17001,N_18366);
nor U20160 (N_20160,N_16226,N_18247);
or U20161 (N_20161,N_15835,N_17392);
or U20162 (N_20162,N_17755,N_15562);
xor U20163 (N_20163,N_18357,N_17147);
xnor U20164 (N_20164,N_18843,N_15516);
or U20165 (N_20165,N_19296,N_17723);
xor U20166 (N_20166,N_17098,N_18717);
nand U20167 (N_20167,N_15059,N_15396);
nor U20168 (N_20168,N_16701,N_16920);
nand U20169 (N_20169,N_19226,N_17096);
and U20170 (N_20170,N_16320,N_16220);
nand U20171 (N_20171,N_18134,N_19122);
and U20172 (N_20172,N_19042,N_16810);
xor U20173 (N_20173,N_19377,N_15254);
or U20174 (N_20174,N_16216,N_16432);
nand U20175 (N_20175,N_16792,N_18765);
nor U20176 (N_20176,N_18354,N_16331);
nand U20177 (N_20177,N_17648,N_16769);
nor U20178 (N_20178,N_18608,N_15661);
or U20179 (N_20179,N_16429,N_19119);
or U20180 (N_20180,N_16022,N_19165);
or U20181 (N_20181,N_16985,N_18751);
xnor U20182 (N_20182,N_15390,N_18598);
nor U20183 (N_20183,N_17792,N_17832);
nand U20184 (N_20184,N_16632,N_16809);
nand U20185 (N_20185,N_16255,N_19408);
or U20186 (N_20186,N_17085,N_15106);
nand U20187 (N_20187,N_17607,N_17592);
xor U20188 (N_20188,N_18380,N_18683);
nand U20189 (N_20189,N_18130,N_19830);
or U20190 (N_20190,N_16834,N_17156);
or U20191 (N_20191,N_15497,N_16516);
nor U20192 (N_20192,N_15539,N_15854);
nand U20193 (N_20193,N_16280,N_16869);
nor U20194 (N_20194,N_18425,N_17658);
nor U20195 (N_20195,N_18747,N_18479);
nor U20196 (N_20196,N_19853,N_15879);
nor U20197 (N_20197,N_15710,N_17895);
or U20198 (N_20198,N_19569,N_15399);
nor U20199 (N_20199,N_17395,N_19927);
nor U20200 (N_20200,N_16464,N_19474);
or U20201 (N_20201,N_18395,N_19257);
and U20202 (N_20202,N_17959,N_19247);
or U20203 (N_20203,N_18456,N_19107);
nand U20204 (N_20204,N_17322,N_19283);
nand U20205 (N_20205,N_16498,N_19346);
nor U20206 (N_20206,N_15141,N_15627);
nand U20207 (N_20207,N_16352,N_19254);
or U20208 (N_20208,N_18795,N_19778);
xnor U20209 (N_20209,N_18553,N_17018);
nand U20210 (N_20210,N_15307,N_18840);
and U20211 (N_20211,N_18752,N_17768);
xnor U20212 (N_20212,N_18703,N_15918);
and U20213 (N_20213,N_18267,N_19490);
or U20214 (N_20214,N_15957,N_16065);
nand U20215 (N_20215,N_18773,N_16340);
xnor U20216 (N_20216,N_18037,N_18470);
or U20217 (N_20217,N_19313,N_17651);
nand U20218 (N_20218,N_17242,N_15921);
nand U20219 (N_20219,N_18581,N_15963);
xnor U20220 (N_20220,N_18670,N_16521);
and U20221 (N_20221,N_18040,N_16031);
and U20222 (N_20222,N_15693,N_17834);
nor U20223 (N_20223,N_16122,N_18923);
nor U20224 (N_20224,N_16930,N_15880);
nand U20225 (N_20225,N_19896,N_17911);
and U20226 (N_20226,N_19295,N_16650);
or U20227 (N_20227,N_19609,N_18101);
or U20228 (N_20228,N_19170,N_15352);
nand U20229 (N_20229,N_19735,N_15191);
or U20230 (N_20230,N_18171,N_16674);
nor U20231 (N_20231,N_18396,N_18278);
nand U20232 (N_20232,N_18988,N_19727);
and U20233 (N_20233,N_16194,N_16435);
or U20234 (N_20234,N_18285,N_18310);
nand U20235 (N_20235,N_15127,N_18558);
nand U20236 (N_20236,N_16709,N_17717);
and U20237 (N_20237,N_19535,N_16490);
nand U20238 (N_20238,N_16544,N_19745);
nand U20239 (N_20239,N_18405,N_17454);
or U20240 (N_20240,N_16906,N_17204);
nand U20241 (N_20241,N_17562,N_18835);
and U20242 (N_20242,N_18692,N_15925);
or U20243 (N_20243,N_15717,N_16713);
or U20244 (N_20244,N_19706,N_16776);
xor U20245 (N_20245,N_17449,N_19858);
nand U20246 (N_20246,N_19358,N_18336);
xor U20247 (N_20247,N_17037,N_17111);
xor U20248 (N_20248,N_18732,N_19807);
or U20249 (N_20249,N_15542,N_16604);
nor U20250 (N_20250,N_18199,N_16975);
xor U20251 (N_20251,N_18032,N_16092);
or U20252 (N_20252,N_18146,N_16887);
nand U20253 (N_20253,N_15772,N_15950);
or U20254 (N_20254,N_19251,N_15013);
nor U20255 (N_20255,N_19552,N_18978);
or U20256 (N_20256,N_15047,N_16893);
or U20257 (N_20257,N_16046,N_15482);
nand U20258 (N_20258,N_19140,N_18712);
or U20259 (N_20259,N_18065,N_19482);
xor U20260 (N_20260,N_15764,N_18067);
or U20261 (N_20261,N_17578,N_18886);
and U20262 (N_20262,N_19159,N_18221);
and U20263 (N_20263,N_16736,N_16510);
and U20264 (N_20264,N_16272,N_16478);
xnor U20265 (N_20265,N_16148,N_19872);
nor U20266 (N_20266,N_18754,N_15472);
xnor U20267 (N_20267,N_19785,N_15545);
nor U20268 (N_20268,N_18868,N_18294);
or U20269 (N_20269,N_17284,N_16925);
or U20270 (N_20270,N_16924,N_19792);
xor U20271 (N_20271,N_18587,N_17625);
xor U20272 (N_20272,N_19419,N_17835);
or U20273 (N_20273,N_19930,N_15235);
xor U20274 (N_20274,N_15201,N_16731);
nor U20275 (N_20275,N_19749,N_17861);
nor U20276 (N_20276,N_18126,N_19902);
nor U20277 (N_20277,N_17672,N_15682);
or U20278 (N_20278,N_17142,N_17992);
or U20279 (N_20279,N_16366,N_19874);
and U20280 (N_20280,N_15558,N_16957);
and U20281 (N_20281,N_18488,N_18105);
or U20282 (N_20282,N_15373,N_15526);
nor U20283 (N_20283,N_18372,N_16168);
nor U20284 (N_20284,N_18196,N_17414);
and U20285 (N_20285,N_16383,N_15566);
nand U20286 (N_20286,N_18656,N_19120);
nand U20287 (N_20287,N_16328,N_15103);
nor U20288 (N_20288,N_17095,N_16646);
xor U20289 (N_20289,N_15485,N_16474);
or U20290 (N_20290,N_19442,N_17593);
xnor U20291 (N_20291,N_15941,N_18337);
nand U20292 (N_20292,N_18924,N_16322);
nand U20293 (N_20293,N_17388,N_18518);
nand U20294 (N_20294,N_16384,N_17097);
xnor U20295 (N_20295,N_17850,N_19542);
and U20296 (N_20296,N_19685,N_16454);
nor U20297 (N_20297,N_18628,N_17348);
or U20298 (N_20298,N_19175,N_16462);
or U20299 (N_20299,N_15376,N_15742);
or U20300 (N_20300,N_18953,N_16381);
nand U20301 (N_20301,N_18458,N_15233);
and U20302 (N_20302,N_19714,N_15505);
and U20303 (N_20303,N_15438,N_15045);
xnor U20304 (N_20304,N_15786,N_19844);
nand U20305 (N_20305,N_19559,N_17505);
nor U20306 (N_20306,N_19991,N_18848);
xor U20307 (N_20307,N_17528,N_15048);
or U20308 (N_20308,N_16997,N_17802);
xor U20309 (N_20309,N_18137,N_17436);
nand U20310 (N_20310,N_15150,N_17174);
or U20311 (N_20311,N_17565,N_18157);
or U20312 (N_20312,N_15645,N_19768);
nand U20313 (N_20313,N_19933,N_18047);
and U20314 (N_20314,N_19264,N_15382);
xor U20315 (N_20315,N_18031,N_15099);
and U20316 (N_20316,N_18237,N_16199);
and U20317 (N_20317,N_18482,N_19999);
xnor U20318 (N_20318,N_16477,N_19832);
and U20319 (N_20319,N_15454,N_19036);
or U20320 (N_20320,N_16696,N_19232);
nand U20321 (N_20321,N_16368,N_15237);
xor U20322 (N_20322,N_17453,N_15931);
nand U20323 (N_20323,N_18659,N_17356);
nand U20324 (N_20324,N_19104,N_16266);
nand U20325 (N_20325,N_19190,N_17165);
nor U20326 (N_20326,N_18548,N_15624);
nor U20327 (N_20327,N_18321,N_18234);
nand U20328 (N_20328,N_17888,N_15697);
nand U20329 (N_20329,N_15997,N_17965);
nand U20330 (N_20330,N_17402,N_18616);
xnor U20331 (N_20331,N_16683,N_18227);
and U20332 (N_20332,N_16350,N_19741);
nand U20333 (N_20333,N_18539,N_19154);
and U20334 (N_20334,N_17586,N_19101);
and U20335 (N_20335,N_16780,N_18609);
or U20336 (N_20336,N_19789,N_16377);
nor U20337 (N_20337,N_18111,N_15729);
and U20338 (N_20338,N_16806,N_17239);
nand U20339 (N_20339,N_19695,N_18643);
nand U20340 (N_20340,N_17086,N_19299);
nand U20341 (N_20341,N_18483,N_18454);
or U20342 (N_20342,N_15952,N_16862);
nor U20343 (N_20343,N_18882,N_16880);
nand U20344 (N_20344,N_16532,N_17937);
nor U20345 (N_20345,N_19585,N_17024);
and U20346 (N_20346,N_16223,N_16149);
or U20347 (N_20347,N_17143,N_17192);
nand U20348 (N_20348,N_15839,N_18825);
nand U20349 (N_20349,N_19805,N_17982);
nor U20350 (N_20350,N_17953,N_19234);
nand U20351 (N_20351,N_19098,N_18726);
or U20352 (N_20352,N_18411,N_19623);
xor U20353 (N_20353,N_18110,N_19824);
and U20354 (N_20354,N_15247,N_19646);
or U20355 (N_20355,N_19448,N_18602);
nand U20356 (N_20356,N_17248,N_16811);
and U20357 (N_20357,N_18573,N_15342);
and U20358 (N_20358,N_16505,N_16312);
nor U20359 (N_20359,N_16970,N_18949);
nand U20360 (N_20360,N_16257,N_19836);
or U20361 (N_20361,N_17237,N_17660);
xnor U20362 (N_20362,N_19353,N_18063);
xor U20363 (N_20363,N_18390,N_15303);
nand U20364 (N_20364,N_19435,N_16718);
nor U20365 (N_20365,N_18315,N_16018);
and U20366 (N_20366,N_15513,N_15129);
xnor U20367 (N_20367,N_15464,N_16129);
xor U20368 (N_20368,N_19109,N_15547);
xor U20369 (N_20369,N_19055,N_15988);
or U20370 (N_20370,N_17915,N_17194);
or U20371 (N_20371,N_19828,N_15859);
nor U20372 (N_20372,N_17532,N_19956);
and U20373 (N_20373,N_15978,N_16936);
nand U20374 (N_20374,N_15453,N_18829);
or U20375 (N_20375,N_16304,N_16918);
and U20376 (N_20376,N_16917,N_19506);
nor U20377 (N_20377,N_19040,N_16064);
nor U20378 (N_20378,N_15423,N_18710);
nor U20379 (N_20379,N_15291,N_17063);
or U20380 (N_20380,N_19043,N_17551);
nand U20381 (N_20381,N_17438,N_15692);
and U20382 (N_20382,N_17474,N_17351);
xnor U20383 (N_20383,N_17278,N_15158);
and U20384 (N_20384,N_19041,N_18145);
nor U20385 (N_20385,N_19534,N_15659);
nand U20386 (N_20386,N_15720,N_15965);
nor U20387 (N_20387,N_17659,N_18967);
and U20388 (N_20388,N_19889,N_16556);
xor U20389 (N_20389,N_17898,N_16325);
or U20390 (N_20390,N_17635,N_15828);
and U20391 (N_20391,N_16428,N_15056);
nand U20392 (N_20392,N_16494,N_16147);
or U20393 (N_20393,N_19751,N_19823);
or U20394 (N_20394,N_15392,N_18084);
nor U20395 (N_20395,N_17842,N_18777);
or U20396 (N_20396,N_17502,N_16002);
xnor U20397 (N_20397,N_15553,N_15620);
nand U20398 (N_20398,N_17434,N_15236);
xor U20399 (N_20399,N_17784,N_17685);
or U20400 (N_20400,N_18869,N_18296);
nor U20401 (N_20401,N_17885,N_17601);
nand U20402 (N_20402,N_16663,N_15725);
or U20403 (N_20403,N_17056,N_18753);
xnor U20404 (N_20404,N_17917,N_17788);
nor U20405 (N_20405,N_17347,N_18964);
nor U20406 (N_20406,N_19182,N_19343);
or U20407 (N_20407,N_15827,N_16823);
nand U20408 (N_20408,N_17196,N_16380);
xor U20409 (N_20409,N_16773,N_15510);
nand U20410 (N_20410,N_19406,N_16956);
nand U20411 (N_20411,N_17827,N_19861);
or U20412 (N_20412,N_19650,N_16507);
nor U20413 (N_20413,N_16849,N_18158);
or U20414 (N_20414,N_15959,N_17952);
or U20415 (N_20415,N_19266,N_16421);
nand U20416 (N_20416,N_19317,N_16671);
nand U20417 (N_20417,N_18734,N_17558);
nor U20418 (N_20418,N_15061,N_16870);
or U20419 (N_20419,N_15524,N_19284);
nand U20420 (N_20420,N_18652,N_18414);
xor U20421 (N_20421,N_15721,N_18055);
or U20422 (N_20422,N_18528,N_19253);
xor U20423 (N_20423,N_18788,N_15649);
xnor U20424 (N_20424,N_19648,N_18073);
or U20425 (N_20425,N_16475,N_18220);
nand U20426 (N_20426,N_16613,N_18798);
nor U20427 (N_20427,N_16682,N_17759);
nand U20428 (N_20428,N_16060,N_15888);
xnor U20429 (N_20429,N_17972,N_17516);
and U20430 (N_20430,N_18416,N_15460);
and U20431 (N_20431,N_17865,N_19596);
xnor U20432 (N_20432,N_17777,N_18412);
nand U20433 (N_20433,N_19303,N_15758);
nor U20434 (N_20434,N_17709,N_15518);
and U20435 (N_20435,N_15700,N_19405);
xnor U20436 (N_20436,N_18800,N_19309);
and U20437 (N_20437,N_18420,N_19574);
or U20438 (N_20438,N_15610,N_15522);
nand U20439 (N_20439,N_17294,N_15109);
xnor U20440 (N_20440,N_15646,N_17031);
nand U20441 (N_20441,N_19855,N_17897);
nand U20442 (N_20442,N_15481,N_15890);
nor U20443 (N_20443,N_17882,N_18085);
xor U20444 (N_20444,N_15671,N_18962);
xor U20445 (N_20445,N_19978,N_17059);
or U20446 (N_20446,N_17857,N_18346);
or U20447 (N_20447,N_17153,N_15084);
xnor U20448 (N_20448,N_19659,N_18516);
or U20449 (N_20449,N_15492,N_17210);
xnor U20450 (N_20450,N_17164,N_15014);
nor U20451 (N_20451,N_19907,N_15051);
nand U20452 (N_20452,N_17618,N_15180);
xor U20453 (N_20453,N_17317,N_19694);
nand U20454 (N_20454,N_15445,N_18045);
or U20455 (N_20455,N_15234,N_18012);
xnor U20456 (N_20456,N_16425,N_18613);
nor U20457 (N_20457,N_18184,N_18173);
and U20458 (N_20458,N_18524,N_18919);
nand U20459 (N_20459,N_15205,N_17631);
xor U20460 (N_20460,N_19241,N_19252);
xnor U20461 (N_20461,N_19617,N_15134);
xnor U20462 (N_20462,N_15424,N_15681);
or U20463 (N_20463,N_17397,N_17557);
nor U20464 (N_20464,N_17418,N_16753);
or U20465 (N_20465,N_15055,N_18383);
nor U20466 (N_20466,N_19180,N_19293);
xnor U20467 (N_20467,N_17363,N_15552);
xor U20468 (N_20468,N_18254,N_16364);
nand U20469 (N_20469,N_18048,N_19787);
xnor U20470 (N_20470,N_15713,N_15092);
or U20471 (N_20471,N_17491,N_15930);
and U20472 (N_20472,N_19595,N_17496);
or U20473 (N_20473,N_18087,N_18678);
xnor U20474 (N_20474,N_17511,N_15707);
nand U20475 (N_20475,N_16117,N_17091);
xor U20476 (N_20476,N_16119,N_18737);
or U20477 (N_20477,N_15258,N_19530);
nand U20478 (N_20478,N_15733,N_17805);
nor U20479 (N_20479,N_19417,N_18371);
and U20480 (N_20480,N_16641,N_15576);
or U20481 (N_20481,N_18606,N_16787);
and U20482 (N_20482,N_16737,N_16241);
nor U20483 (N_20483,N_19513,N_18654);
nand U20484 (N_20484,N_16111,N_19547);
and U20485 (N_20485,N_18298,N_19786);
or U20486 (N_20486,N_18578,N_18530);
nor U20487 (N_20487,N_15806,N_15804);
and U20488 (N_20488,N_15724,N_16555);
nand U20489 (N_20489,N_16347,N_17787);
and U20490 (N_20490,N_17123,N_16557);
nand U20491 (N_20491,N_19953,N_17376);
nor U20492 (N_20492,N_18117,N_15118);
nor U20493 (N_20493,N_15252,N_18627);
and U20494 (N_20494,N_19636,N_18050);
and U20495 (N_20495,N_16181,N_19654);
nand U20496 (N_20496,N_16706,N_18286);
nand U20497 (N_20497,N_17288,N_16450);
nor U20498 (N_20498,N_15567,N_18116);
nand U20499 (N_20499,N_16601,N_16690);
or U20500 (N_20500,N_19776,N_17761);
and U20501 (N_20501,N_19833,N_18580);
and U20502 (N_20502,N_17180,N_17325);
nor U20503 (N_20503,N_15228,N_19375);
and U20504 (N_20504,N_17679,N_19891);
xor U20505 (N_20505,N_18256,N_15861);
or U20506 (N_20506,N_17140,N_15320);
nand U20507 (N_20507,N_19038,N_16135);
or U20508 (N_20508,N_16230,N_18612);
and U20509 (N_20509,N_17178,N_19176);
nand U20510 (N_20510,N_19527,N_15884);
nand U20511 (N_20511,N_15613,N_16865);
or U20512 (N_20512,N_18600,N_19740);
nand U20513 (N_20513,N_18466,N_17042);
nor U20514 (N_20514,N_16467,N_15208);
and U20515 (N_20515,N_17490,N_16339);
nand U20516 (N_20516,N_19952,N_16351);
or U20517 (N_20517,N_15469,N_19431);
xor U20518 (N_20518,N_15560,N_17330);
or U20519 (N_20519,N_16459,N_18056);
nor U20520 (N_20520,N_17328,N_16013);
or U20521 (N_20521,N_16842,N_15546);
nand U20522 (N_20522,N_18295,N_16296);
nand U20523 (N_20523,N_18242,N_19583);
xor U20524 (N_20524,N_16791,N_16609);
and U20525 (N_20525,N_18291,N_16444);
and U20526 (N_20526,N_17688,N_16099);
nand U20527 (N_20527,N_19230,N_18431);
and U20528 (N_20528,N_16540,N_18714);
xor U20529 (N_20529,N_19439,N_17615);
and U20530 (N_20530,N_16897,N_17863);
nand U20531 (N_20531,N_16982,N_17231);
or U20532 (N_20532,N_16726,N_16044);
and U20533 (N_20533,N_19308,N_19279);
and U20534 (N_20534,N_17657,N_19643);
and U20535 (N_20535,N_16003,N_19132);
nand U20536 (N_20536,N_19656,N_16393);
nand U20537 (N_20537,N_18075,N_19763);
xnor U20538 (N_20538,N_15290,N_17515);
and U20539 (N_20539,N_15203,N_17051);
or U20540 (N_20540,N_15372,N_15273);
and U20541 (N_20541,N_18292,N_18903);
and U20542 (N_20542,N_19666,N_17112);
and U20543 (N_20543,N_19328,N_19380);
or U20544 (N_20544,N_17694,N_16785);
xor U20545 (N_20545,N_19362,N_18208);
xor U20546 (N_20546,N_18341,N_17486);
xor U20547 (N_20547,N_17267,N_15073);
or U20548 (N_20548,N_18144,N_17896);
xnor U20549 (N_20549,N_15763,N_17577);
nand U20550 (N_20550,N_19015,N_15537);
and U20551 (N_20551,N_15732,N_18972);
and U20552 (N_20552,N_15444,N_15934);
and U20553 (N_20553,N_16578,N_19393);
or U20554 (N_20554,N_16538,N_15130);
or U20555 (N_20555,N_18914,N_17971);
xnor U20556 (N_20556,N_18845,N_15583);
nor U20557 (N_20557,N_17706,N_19188);
or U20558 (N_20558,N_17398,N_19321);
nor U20559 (N_20559,N_15142,N_19359);
and U20560 (N_20560,N_15410,N_19704);
nor U20561 (N_20561,N_19944,N_16375);
nand U20562 (N_20562,N_16725,N_19007);
and U20563 (N_20563,N_15421,N_19750);
xor U20564 (N_20564,N_17384,N_18092);
nand U20565 (N_20565,N_17352,N_18941);
nor U20566 (N_20566,N_17945,N_17671);
xor U20567 (N_20567,N_18408,N_15500);
nand U20568 (N_20568,N_15466,N_18533);
and U20569 (N_20569,N_19555,N_15090);
nand U20570 (N_20570,N_17853,N_16323);
nand U20571 (N_20571,N_16088,N_15128);
xnor U20572 (N_20572,N_16728,N_16314);
xnor U20573 (N_20573,N_19385,N_16911);
nand U20574 (N_20574,N_15315,N_17250);
and U20575 (N_20575,N_19151,N_19001);
nor U20576 (N_20576,N_17057,N_19387);
or U20577 (N_20577,N_15436,N_17197);
nor U20578 (N_20578,N_15967,N_16193);
nand U20579 (N_20579,N_18900,N_18956);
nand U20580 (N_20580,N_16665,N_19192);
or U20581 (N_20581,N_18968,N_16771);
and U20582 (N_20582,N_16275,N_17910);
xnor U20583 (N_20583,N_15531,N_15032);
and U20584 (N_20584,N_15885,N_15490);
or U20585 (N_20585,N_19235,N_16829);
nand U20586 (N_20586,N_16136,N_19430);
nor U20587 (N_20587,N_15304,N_19322);
nor U20588 (N_20588,N_18507,N_15789);
nor U20589 (N_20589,N_16011,N_15829);
nor U20590 (N_20590,N_16967,N_17193);
or U20591 (N_20591,N_18397,N_19647);
xnor U20592 (N_20592,N_17054,N_15960);
nand U20593 (N_20593,N_16611,N_16007);
nor U20594 (N_20594,N_15657,N_15036);
or U20595 (N_20595,N_17306,N_19286);
nand U20596 (N_20596,N_19110,N_15782);
nor U20597 (N_20597,N_17877,N_15428);
nor U20598 (N_20598,N_17137,N_19456);
or U20599 (N_20599,N_16622,N_17387);
and U20600 (N_20600,N_19081,N_19551);
or U20601 (N_20601,N_16824,N_18025);
xor U20602 (N_20602,N_16868,N_16009);
nand U20603 (N_20603,N_15544,N_15812);
nor U20604 (N_20604,N_15690,N_18435);
nand U20605 (N_20605,N_16150,N_19621);
and U20606 (N_20606,N_19124,N_16672);
nand U20607 (N_20607,N_18307,N_18922);
nor U20608 (N_20608,N_17594,N_17364);
xnor U20609 (N_20609,N_19412,N_16596);
xor U20610 (N_20610,N_15337,N_15901);
nand U20611 (N_20611,N_15394,N_17393);
nand U20612 (N_20612,N_19118,N_16667);
and U20613 (N_20613,N_18595,N_19762);
xor U20614 (N_20614,N_18030,N_18407);
nor U20615 (N_20615,N_19281,N_16670);
and U20616 (N_20616,N_16681,N_17650);
xor U20617 (N_20617,N_18546,N_15149);
or U20618 (N_20618,N_17168,N_18662);
nor U20619 (N_20619,N_16126,N_16644);
xor U20620 (N_20620,N_17763,N_19423);
or U20621 (N_20621,N_19843,N_16160);
nor U20622 (N_20622,N_15439,N_16248);
nor U20623 (N_20623,N_19139,N_19237);
nand U20624 (N_20624,N_18485,N_15271);
and U20625 (N_20625,N_18094,N_16919);
nor U20626 (N_20626,N_16828,N_16413);
nand U20627 (N_20627,N_19711,N_18238);
nor U20628 (N_20628,N_18880,N_19425);
nand U20629 (N_20629,N_19628,N_18430);
nor U20630 (N_20630,N_16045,N_17148);
nor U20631 (N_20631,N_17526,N_16590);
or U20632 (N_20632,N_18190,N_18660);
nor U20633 (N_20633,N_19518,N_18839);
or U20634 (N_20634,N_17697,N_15289);
and U20635 (N_20635,N_15222,N_17421);
nor U20636 (N_20636,N_17233,N_15617);
xnor U20637 (N_20637,N_17003,N_16837);
or U20638 (N_20638,N_15629,N_16026);
and U20639 (N_20639,N_18687,N_16372);
nand U20640 (N_20640,N_15604,N_18679);
nand U20641 (N_20641,N_16027,N_15683);
and U20642 (N_20642,N_16568,N_15961);
nand U20643 (N_20643,N_15338,N_16677);
or U20644 (N_20644,N_18082,N_19006);
nor U20645 (N_20645,N_15412,N_18861);
or U20646 (N_20646,N_18020,N_18876);
nand U20647 (N_20647,N_16748,N_15223);
nand U20648 (N_20648,N_18452,N_19642);
and U20649 (N_20649,N_15066,N_19705);
nand U20650 (N_20650,N_16299,N_18774);
and U20651 (N_20651,N_15361,N_16237);
xnor U20652 (N_20652,N_15634,N_18973);
or U20653 (N_20653,N_16500,N_15768);
xor U20654 (N_20654,N_19893,N_17214);
or U20655 (N_20655,N_17859,N_17595);
nand U20656 (N_20656,N_15603,N_16624);
or U20657 (N_20657,N_18695,N_18179);
nor U20658 (N_20658,N_17206,N_17349);
or U20659 (N_20659,N_15696,N_17485);
and U20660 (N_20660,N_16177,N_19980);
nand U20661 (N_20661,N_18148,N_15496);
xor U20662 (N_20662,N_19878,N_15487);
nor U20663 (N_20663,N_15691,N_17312);
and U20664 (N_20664,N_16190,N_16120);
nand U20665 (N_20665,N_16852,N_17727);
xor U20666 (N_20666,N_17762,N_18230);
nor U20667 (N_20667,N_16503,N_19127);
or U20668 (N_20668,N_19102,N_17724);
and U20669 (N_20669,N_17542,N_19985);
nand U20670 (N_20670,N_15299,N_17666);
nand U20671 (N_20671,N_16415,N_16131);
or U20672 (N_20672,N_19616,N_17841);
xor U20673 (N_20673,N_17831,N_15097);
or U20674 (N_20674,N_16520,N_18477);
nor U20675 (N_20675,N_19185,N_16914);
or U20676 (N_20676,N_19152,N_15367);
xor U20677 (N_20677,N_19717,N_18965);
nand U20678 (N_20678,N_19783,N_17998);
nor U20679 (N_20679,N_16605,N_16756);
xor U20680 (N_20680,N_19056,N_18667);
xnor U20681 (N_20681,N_17446,N_19093);
nor U20682 (N_20682,N_16227,N_17425);
and U20683 (N_20683,N_19868,N_18021);
nor U20684 (N_20684,N_19444,N_15877);
or U20685 (N_20685,N_16493,N_19564);
and U20686 (N_20686,N_17020,N_16030);
nand U20687 (N_20687,N_15152,N_16749);
nand U20688 (N_20688,N_17396,N_15136);
nor U20689 (N_20689,N_19184,N_18358);
nand U20690 (N_20690,N_16835,N_16260);
xor U20691 (N_20691,N_18240,N_19106);
nand U20692 (N_20692,N_17276,N_16714);
and U20693 (N_20693,N_18691,N_15962);
or U20694 (N_20694,N_15062,N_15385);
nor U20695 (N_20695,N_16819,N_19722);
and U20696 (N_20696,N_19243,N_16042);
nor U20697 (N_20697,N_16016,N_19661);
nand U20698 (N_20698,N_17235,N_17498);
and U20699 (N_20699,N_18006,N_18772);
or U20700 (N_20700,N_18114,N_19379);
and U20701 (N_20701,N_18233,N_17000);
xnor U20702 (N_20702,N_16205,N_17493);
xor U20703 (N_20703,N_17407,N_18480);
xor U20704 (N_20704,N_19683,N_17251);
and U20705 (N_20705,N_15639,N_18155);
xnor U20706 (N_20706,N_15656,N_19629);
and U20707 (N_20707,N_15011,N_19094);
and U20708 (N_20708,N_18827,N_17993);
nor U20709 (N_20709,N_17646,N_19850);
or U20710 (N_20710,N_15830,N_15841);
nand U20711 (N_20711,N_15587,N_17600);
xor U20712 (N_20712,N_19914,N_19949);
nor U20713 (N_20713,N_16420,N_16903);
xor U20714 (N_20714,N_17588,N_17136);
or U20715 (N_20715,N_16987,N_19873);
xnor U20716 (N_20716,N_19202,N_15549);
xor U20717 (N_20717,N_16253,N_18631);
or U20718 (N_20718,N_17879,N_17731);
or U20719 (N_20719,N_17662,N_15095);
xor U20720 (N_20720,N_15411,N_19876);
or U20721 (N_20721,N_18623,N_19024);
nor U20722 (N_20722,N_16569,N_15582);
xnor U20723 (N_20723,N_17932,N_15040);
and U20724 (N_20724,N_19462,N_17464);
nor U20725 (N_20725,N_15667,N_16574);
xnor U20726 (N_20726,N_19682,N_16816);
and U20727 (N_20727,N_15631,N_15817);
xor U20728 (N_20728,N_16922,N_15565);
nand U20729 (N_20729,N_18159,N_15096);
or U20730 (N_20730,N_19492,N_16699);
nand U20731 (N_20731,N_19626,N_19062);
nand U20732 (N_20732,N_18532,N_15573);
nor U20733 (N_20733,N_16745,N_17734);
or U20734 (N_20734,N_17072,N_19333);
xnor U20735 (N_20735,N_17240,N_17026);
and U20736 (N_20736,N_16760,N_15781);
and U20737 (N_20737,N_17359,N_17941);
nand U20738 (N_20738,N_18232,N_16360);
or U20739 (N_20739,N_18072,N_17944);
nor U20740 (N_20740,N_16451,N_17487);
and U20741 (N_20741,N_16221,N_16301);
nand U20742 (N_20742,N_17326,N_19607);
nor U20743 (N_20743,N_15407,N_18402);
and U20744 (N_20744,N_19206,N_16946);
and U20745 (N_20745,N_19080,N_16993);
xor U20746 (N_20746,N_17745,N_17570);
xor U20747 (N_20747,N_15473,N_17852);
or U20748 (N_20748,N_17340,N_19712);
and U20749 (N_20749,N_15270,N_19452);
or U20750 (N_20750,N_19085,N_16537);
nor U20751 (N_20751,N_18326,N_18637);
nand U20752 (N_20752,N_17120,N_19515);
and U20753 (N_20753,N_17228,N_15194);
xnor U20754 (N_20754,N_16598,N_19466);
and U20755 (N_20755,N_15694,N_16759);
and U20756 (N_20756,N_15938,N_18935);
or U20757 (N_20757,N_15022,N_17126);
xnor U20758 (N_20758,N_19501,N_16200);
xor U20759 (N_20759,N_19048,N_17344);
xor U20760 (N_20760,N_17583,N_17247);
or U20761 (N_20761,N_17177,N_15818);
and U20762 (N_20762,N_19147,N_16784);
nand U20763 (N_20763,N_17411,N_16326);
xor U20764 (N_20764,N_15752,N_19516);
or U20765 (N_20765,N_17299,N_15046);
xor U20766 (N_20766,N_15592,N_17121);
nand U20767 (N_20767,N_15297,N_17188);
or U20768 (N_20768,N_17378,N_17224);
nor U20769 (N_20769,N_18635,N_19812);
and U20770 (N_20770,N_17070,N_15192);
xnor U20771 (N_20771,N_16015,N_16790);
xor U20772 (N_20772,N_15265,N_15322);
nor U20773 (N_20773,N_17799,N_18127);
nand U20774 (N_20774,N_18163,N_18214);
nand U20775 (N_20775,N_15256,N_16043);
nand U20776 (N_20776,N_18484,N_16496);
nand U20777 (N_20777,N_19223,N_16620);
nor U20778 (N_20778,N_16021,N_16702);
or U20779 (N_20779,N_19113,N_17524);
xnor U20780 (N_20780,N_18644,N_19529);
or U20781 (N_20781,N_17171,N_18819);
or U20782 (N_20782,N_16234,N_15155);
and U20783 (N_20783,N_16591,N_18981);
nand U20784 (N_20784,N_19536,N_18887);
nand U20785 (N_20785,N_18519,N_15086);
nand U20786 (N_20786,N_19619,N_16912);
xor U20787 (N_20787,N_16645,N_16827);
and U20788 (N_20788,N_17107,N_17447);
nor U20789 (N_20789,N_17357,N_18474);
xnor U20790 (N_20790,N_19499,N_17441);
nand U20791 (N_20791,N_19128,N_15173);
and U20792 (N_20792,N_18989,N_17881);
xnor U20793 (N_20793,N_16083,N_16511);
or U20794 (N_20794,N_17064,N_18394);
xor U20795 (N_20795,N_19149,N_16302);
and U20796 (N_20796,N_19769,N_18552);
and U20797 (N_20797,N_15899,N_16004);
or U20798 (N_20798,N_18120,N_15590);
nor U20799 (N_20799,N_15172,N_15079);
xor U20800 (N_20800,N_16483,N_17909);
xnor U20801 (N_20801,N_16074,N_18713);
or U20802 (N_20802,N_19875,N_17628);
and U20803 (N_20803,N_17404,N_18102);
xnor U20804 (N_20804,N_18915,N_17668);
or U20805 (N_20805,N_18209,N_19066);
and U20806 (N_20806,N_15916,N_17617);
nor U20807 (N_20807,N_17368,N_17919);
or U20808 (N_20808,N_16536,N_18760);
xnor U20809 (N_20809,N_18585,N_17290);
xnor U20810 (N_20810,N_19665,N_15251);
nand U20811 (N_20811,N_17684,N_17336);
nor U20812 (N_20812,N_17078,N_19565);
or U20813 (N_20813,N_19278,N_19177);
nand U20814 (N_20814,N_17517,N_17100);
nand U20815 (N_20815,N_18818,N_19773);
nand U20816 (N_20816,N_18250,N_15499);
nand U20817 (N_20817,N_19637,N_16891);
or U20818 (N_20818,N_18682,N_19511);
or U20819 (N_20819,N_15614,N_15114);
xnor U20820 (N_20820,N_16529,N_18725);
and U20821 (N_20821,N_18000,N_16877);
xor U20822 (N_20822,N_16767,N_15282);
or U20823 (N_20823,N_17687,N_18008);
and U20824 (N_20824,N_18178,N_19716);
and U20825 (N_20825,N_16307,N_16209);
and U20826 (N_20826,N_19378,N_17225);
and U20827 (N_20827,N_15908,N_15184);
nor U20828 (N_20828,N_17608,N_16802);
nand U20829 (N_20829,N_17305,N_15801);
and U20830 (N_20830,N_17538,N_19033);
nor U20831 (N_20831,N_15112,N_19854);
and U20832 (N_20832,N_17812,N_16694);
nand U20833 (N_20833,N_19720,N_19684);
or U20834 (N_20834,N_19988,N_17988);
nor U20835 (N_20835,N_18288,N_19968);
nand U20836 (N_20836,N_19926,N_19514);
or U20837 (N_20837,N_18853,N_19220);
and U20838 (N_20838,N_17207,N_18010);
nor U20839 (N_20839,N_16426,N_17243);
and U20840 (N_20840,N_16546,N_15787);
nor U20841 (N_20841,N_15329,N_15360);
nor U20842 (N_20842,N_16999,N_19732);
nor U20843 (N_20843,N_15648,N_17775);
or U20844 (N_20844,N_17254,N_16589);
nand U20845 (N_20845,N_18305,N_19986);
xnor U20846 (N_20846,N_19897,N_16482);
nor U20847 (N_20847,N_18700,N_18838);
nor U20848 (N_20848,N_19172,N_16093);
nor U20849 (N_20849,N_16349,N_17629);
nor U20850 (N_20850,N_18834,N_15334);
nor U20851 (N_20851,N_17793,N_17475);
and U20852 (N_20852,N_18970,N_18808);
or U20853 (N_20853,N_19691,N_16958);
xnor U20854 (N_20854,N_15895,N_19938);
xor U20855 (N_20855,N_17400,N_19434);
nand U20856 (N_20856,N_19087,N_18428);
nor U20857 (N_20857,N_16162,N_19924);
nand U20858 (N_20858,N_15714,N_19357);
or U20859 (N_20859,N_15712,N_16281);
and U20860 (N_20860,N_15495,N_17465);
xor U20861 (N_20861,N_19179,N_19138);
nor U20862 (N_20862,N_18770,N_19934);
nand U20863 (N_20863,N_17539,N_15832);
nand U20864 (N_20864,N_18098,N_19143);
and U20865 (N_20865,N_15672,N_17431);
and U20866 (N_20866,N_16192,N_18640);
and U20867 (N_20867,N_17315,N_15246);
nand U20868 (N_20868,N_16916,N_15384);
nor U20869 (N_20869,N_15309,N_17190);
xnor U20870 (N_20870,N_16186,N_15622);
and U20871 (N_20871,N_16305,N_16928);
and U20872 (N_20872,N_19407,N_18872);
or U20873 (N_20873,N_18338,N_17955);
xnor U20874 (N_20874,N_18723,N_17280);
or U20875 (N_20875,N_18863,N_18610);
xor U20876 (N_20876,N_18750,N_17105);
or U20877 (N_20877,N_19025,N_19486);
and U20878 (N_20878,N_16469,N_16739);
xor U20879 (N_20879,N_16715,N_15991);
or U20880 (N_20880,N_17027,N_17321);
xor U20881 (N_20881,N_17236,N_18064);
or U20882 (N_20882,N_17634,N_19131);
nand U20883 (N_20883,N_17925,N_18205);
nor U20884 (N_20884,N_15577,N_16324);
nor U20885 (N_20885,N_17912,N_15012);
and U20886 (N_20886,N_18515,N_19508);
and U20887 (N_20887,N_16337,N_16139);
or U20888 (N_20888,N_18034,N_16434);
and U20889 (N_20889,N_15595,N_16535);
and U20890 (N_20890,N_19560,N_18038);
or U20891 (N_20891,N_15475,N_19340);
and U20892 (N_20892,N_15715,N_16900);
nand U20893 (N_20893,N_18534,N_16402);
and U20894 (N_20894,N_15431,N_15224);
xor U20895 (N_20895,N_17437,N_16388);
or U20896 (N_20896,N_16386,N_16379);
or U20897 (N_20897,N_18653,N_17350);
or U20898 (N_20898,N_16412,N_16669);
xor U20899 (N_20899,N_19590,N_18511);
nor U20900 (N_20900,N_15442,N_17935);
nand U20901 (N_20901,N_18393,N_16560);
nand U20902 (N_20902,N_17202,N_17710);
nor U20903 (N_20903,N_17726,N_19825);
nand U20904 (N_20904,N_15579,N_19929);
nor U20905 (N_20905,N_16284,N_19020);
or U20906 (N_20906,N_18864,N_19903);
xnor U20907 (N_20907,N_17122,N_16075);
and U20908 (N_20908,N_16218,N_16243);
nor U20909 (N_20909,N_18186,N_15860);
and U20910 (N_20910,N_16416,N_17360);
nor U20911 (N_20911,N_17567,N_17302);
nand U20912 (N_20912,N_17011,N_17596);
and U20913 (N_20913,N_17733,N_19573);
nor U20914 (N_20914,N_16025,N_17323);
nor U20915 (N_20915,N_16566,N_18169);
xor U20916 (N_20916,N_16330,N_19418);
and U20917 (N_20917,N_17052,N_16907);
nor U20918 (N_20918,N_16962,N_15678);
nand U20919 (N_20919,N_18846,N_15776);
xor U20920 (N_20920,N_17334,N_15628);
or U20921 (N_20921,N_16539,N_15984);
nor U20922 (N_20922,N_19627,N_17813);
and U20923 (N_20923,N_18715,N_18841);
and U20924 (N_20924,N_18215,N_16169);
xor U20925 (N_20925,N_17119,N_16053);
nand U20926 (N_20926,N_15087,N_18248);
or U20927 (N_20927,N_16858,N_15953);
nor U20928 (N_20928,N_15777,N_15457);
nand U20929 (N_20929,N_15006,N_17975);
xnor U20930 (N_20930,N_15311,N_15550);
and U20931 (N_20931,N_16315,N_17752);
and U20932 (N_20932,N_15476,N_18614);
nor U20933 (N_20933,N_18364,N_18496);
nand U20934 (N_20934,N_19306,N_17118);
nor U20935 (N_20935,N_15243,N_16676);
or U20936 (N_20936,N_19925,N_18343);
nand U20937 (N_20937,N_19593,N_19859);
nand U20938 (N_20938,N_16680,N_15593);
and U20939 (N_20939,N_18370,N_15640);
or U20940 (N_20940,N_15973,N_16603);
or U20941 (N_20941,N_17152,N_16822);
nor U20942 (N_20942,N_19285,N_19483);
nand U20943 (N_20943,N_16176,N_17716);
nor U20944 (N_20944,N_19133,N_17353);
nand U20945 (N_20945,N_18079,N_19817);
nand U20946 (N_20946,N_16259,N_17815);
or U20947 (N_20947,N_17967,N_15515);
nand U20948 (N_20948,N_17531,N_17090);
and U20949 (N_20949,N_17630,N_17826);
nand U20950 (N_20950,N_16250,N_15755);
nand U20951 (N_20951,N_19302,N_15214);
xnor U20952 (N_20952,N_17016,N_17403);
nand U20953 (N_20953,N_17568,N_17132);
xnor U20954 (N_20954,N_15796,N_17699);
nor U20955 (N_20955,N_16528,N_17048);
xnor U20956 (N_20956,N_19497,N_16817);
and U20957 (N_20957,N_18074,N_16664);
or U20958 (N_20958,N_17848,N_18004);
nor U20959 (N_20959,N_19915,N_15745);
and U20960 (N_20960,N_17253,N_15824);
or U20961 (N_20961,N_19238,N_17683);
nand U20962 (N_20962,N_18057,N_16652);
nor U20963 (N_20963,N_17104,N_16481);
and U20964 (N_20964,N_17598,N_17891);
and U20965 (N_20965,N_16417,N_17905);
xnor U20966 (N_20966,N_17375,N_15943);
xnor U20967 (N_20967,N_19972,N_18175);
or U20968 (N_20968,N_17451,N_15433);
nand U20969 (N_20969,N_17808,N_16992);
and U20970 (N_20970,N_18832,N_15060);
or U20971 (N_20971,N_17543,N_15819);
xor U20972 (N_20972,N_17468,N_18429);
xnor U20973 (N_20973,N_17737,N_18810);
nor U20974 (N_20974,N_19021,N_16866);
or U20975 (N_20975,N_16955,N_18513);
or U20976 (N_20976,N_18361,N_16821);
xor U20977 (N_20977,N_19935,N_19524);
nand U20978 (N_20978,N_19838,N_19123);
xnor U20979 (N_20979,N_18290,N_18918);
nor U20980 (N_20980,N_19401,N_16143);
nand U20981 (N_20981,N_15417,N_17015);
and U20982 (N_20982,N_17219,N_15813);
and U20983 (N_20983,N_19641,N_17663);
xnor U20984 (N_20984,N_17461,N_15067);
nor U20985 (N_20985,N_16639,N_19307);
nand U20986 (N_20986,N_15528,N_17677);
nor U20987 (N_20987,N_19342,N_15494);
nand U20988 (N_20988,N_17007,N_18883);
nor U20989 (N_20989,N_15655,N_16523);
and U20990 (N_20990,N_18870,N_18289);
and U20991 (N_20991,N_15520,N_18453);
nor U20992 (N_20992,N_16121,N_16146);
and U20993 (N_20993,N_17869,N_15939);
nor U20994 (N_20994,N_19702,N_19354);
or U20995 (N_20995,N_19707,N_18815);
nand U20996 (N_20996,N_18333,N_16774);
xnor U20997 (N_20997,N_15321,N_16145);
nor U20998 (N_20998,N_16424,N_18542);
xor U20999 (N_20999,N_15186,N_19886);
nor U21000 (N_21000,N_17405,N_19550);
nor U21001 (N_21001,N_18658,N_16588);
nor U21002 (N_21002,N_19806,N_16175);
or U21003 (N_21003,N_17374,N_15596);
or U21004 (N_21004,N_18878,N_19409);
or U21005 (N_21005,N_17872,N_17066);
xnor U21006 (N_21006,N_15883,N_19111);
and U21007 (N_21007,N_15913,N_19075);
xor U21008 (N_21008,N_18349,N_18514);
or U21009 (N_21009,N_17452,N_15705);
and U21010 (N_21010,N_18650,N_18391);
nor U21011 (N_21011,N_17970,N_15589);
or U21012 (N_21012,N_19117,N_16319);
and U21013 (N_21013,N_17361,N_19586);
nor U21014 (N_21014,N_18044,N_18156);
xnor U21015 (N_21015,N_17301,N_18521);
nor U21016 (N_21016,N_18257,N_16265);
xnor U21017 (N_21017,N_17222,N_17563);
xnor U21018 (N_21018,N_17753,N_18243);
nor U21019 (N_21019,N_15695,N_16134);
or U21020 (N_21020,N_17220,N_17983);
nor U21021 (N_21021,N_15189,N_19888);
and U21022 (N_21022,N_16293,N_16952);
xnor U21023 (N_21023,N_19031,N_18124);
or U21024 (N_21024,N_18709,N_15024);
and U21025 (N_21025,N_16519,N_16549);
and U21026 (N_21026,N_17610,N_15000);
xnor U21027 (N_21027,N_17319,N_19099);
or U21028 (N_21028,N_17483,N_17282);
or U21029 (N_21029,N_19197,N_18450);
nor U21030 (N_21030,N_15730,N_19316);
xor U21031 (N_21031,N_16172,N_16480);
xor U21032 (N_21032,N_16051,N_15292);
and U21033 (N_21033,N_18168,N_16857);
or U21034 (N_21034,N_18392,N_17423);
or U21035 (N_21035,N_18141,N_17829);
nor U21036 (N_21036,N_17466,N_19181);
nor U21037 (N_21037,N_19947,N_15115);
nor U21038 (N_21038,N_19561,N_17013);
or U21039 (N_21039,N_19049,N_16489);
nand U21040 (N_21040,N_15598,N_15569);
or U21041 (N_21041,N_16990,N_18554);
and U21042 (N_21042,N_15615,N_19829);
or U21043 (N_21043,N_17139,N_19034);
or U21044 (N_21044,N_15199,N_18119);
and U21045 (N_21045,N_19849,N_19939);
and U21046 (N_21046,N_18472,N_15740);
and U21047 (N_21047,N_17892,N_15775);
nand U21048 (N_21048,N_17481,N_19957);
nor U21049 (N_21049,N_16630,N_17951);
or U21050 (N_21050,N_17450,N_17170);
xor U21051 (N_21051,N_15076,N_17367);
xor U21052 (N_21052,N_18109,N_18347);
nor U21053 (N_21053,N_17783,N_19277);
xor U21054 (N_21054,N_18059,N_16072);
and U21055 (N_21055,N_17612,N_16843);
xor U21056 (N_21056,N_17605,N_19023);
or U21057 (N_21057,N_15535,N_17145);
or U21058 (N_21058,N_19310,N_16562);
and U21059 (N_21059,N_17033,N_15213);
xor U21060 (N_21060,N_15182,N_18125);
or U21061 (N_21061,N_16224,N_17069);
nor U21062 (N_21062,N_16581,N_18745);
or U21063 (N_21063,N_15365,N_17435);
and U21064 (N_21064,N_17509,N_16994);
or U21065 (N_21065,N_15268,N_17408);
and U21066 (N_21066,N_18579,N_15702);
nor U21067 (N_21067,N_16066,N_18211);
and U21068 (N_21068,N_16636,N_17017);
xnor U21069 (N_21069,N_18550,N_18824);
xnor U21070 (N_21070,N_19557,N_15317);
nand U21071 (N_21071,N_16222,N_18113);
or U21072 (N_21072,N_19579,N_15635);
and U21073 (N_21073,N_17469,N_15906);
or U21074 (N_21074,N_17179,N_15391);
and U21075 (N_21075,N_18415,N_18301);
xor U21076 (N_21076,N_18857,N_19958);
or U21077 (N_21077,N_15071,N_18035);
or U21078 (N_21078,N_16673,N_16487);
and U21079 (N_21079,N_17973,N_15644);
and U21080 (N_21080,N_16801,N_15842);
or U21081 (N_21081,N_16017,N_17094);
nand U21082 (N_21082,N_18561,N_18786);
nor U21083 (N_21083,N_15232,N_15788);
and U21084 (N_21084,N_17544,N_18497);
nor U21085 (N_21085,N_17703,N_17157);
or U21086 (N_21086,N_15478,N_16762);
nand U21087 (N_21087,N_17252,N_19979);
xor U21088 (N_21088,N_19070,N_16976);
nor U21089 (N_21089,N_17135,N_16274);
nor U21090 (N_21090,N_18517,N_17715);
xnor U21091 (N_21091,N_17867,N_17457);
nor U21092 (N_21092,N_17948,N_18260);
nor U21093 (N_21093,N_19005,N_15666);
nand U21094 (N_21094,N_15975,N_19729);
nor U21095 (N_21095,N_17390,N_18368);
and U21096 (N_21096,N_18822,N_18619);
nor U21097 (N_21097,N_15463,N_16138);
and U21098 (N_21098,N_15137,N_16988);
nand U21099 (N_21099,N_15443,N_17673);
nor U21100 (N_21100,N_17488,N_17738);
and U21101 (N_21101,N_18096,N_15441);
nor U21102 (N_21102,N_17124,N_16693);
and U21103 (N_21103,N_19604,N_15353);
nand U21104 (N_21104,N_18365,N_16874);
and U21105 (N_21105,N_15452,N_18642);
nor U21106 (N_21106,N_17921,N_18374);
xor U21107 (N_21107,N_15379,N_16940);
or U21108 (N_21108,N_17036,N_18225);
and U21109 (N_21109,N_19697,N_15295);
xnor U21110 (N_21110,N_17748,N_15856);
xor U21111 (N_21111,N_18107,N_16163);
xor U21112 (N_21112,N_19819,N_19772);
and U21113 (N_21113,N_16734,N_15853);
nor U21114 (N_21114,N_16161,N_16298);
xor U21115 (N_21115,N_18564,N_16385);
and U21116 (N_21116,N_18566,N_17223);
and U21117 (N_21117,N_16392,N_15570);
nor U21118 (N_21118,N_17548,N_18671);
and U21119 (N_21119,N_18487,N_15404);
or U21120 (N_21120,N_19245,N_18625);
and U21121 (N_21121,N_15922,N_17409);
nand U21122 (N_21122,N_19961,N_17127);
nor U21123 (N_21123,N_15909,N_17985);
nor U21124 (N_21124,N_17433,N_18711);
and U21125 (N_21125,N_18066,N_19084);
and U21126 (N_21126,N_15318,N_19082);
and U21127 (N_21127,N_19289,N_18837);
nand U21128 (N_21128,N_17669,N_17261);
nor U21129 (N_21129,N_18702,N_15766);
and U21130 (N_21130,N_16485,N_18593);
nor U21131 (N_21131,N_15995,N_17429);
xnor U21132 (N_21132,N_16779,N_16142);
and U21133 (N_21133,N_18620,N_16398);
and U21134 (N_21134,N_18297,N_15958);
xor U21135 (N_21135,N_15039,N_17274);
nand U21136 (N_21136,N_19187,N_17856);
nand U21137 (N_21137,N_17824,N_17088);
and U21138 (N_21138,N_18499,N_16056);
or U21139 (N_21139,N_16798,N_19718);
and U21140 (N_21140,N_15171,N_19906);
nor U21141 (N_21141,N_19205,N_19919);
nand U21142 (N_21142,N_19416,N_18467);
and U21143 (N_21143,N_17244,N_17144);
nand U21144 (N_21144,N_19791,N_15255);
nor U21145 (N_21145,N_19608,N_15294);
nand U21146 (N_21146,N_15179,N_19793);
xnor U21147 (N_21147,N_18300,N_17028);
or U21148 (N_21148,N_16850,N_19090);
xor U21149 (N_21149,N_19164,N_16104);
xor U21150 (N_21150,N_16593,N_16808);
nand U21151 (N_21151,N_19198,N_15753);
or U21152 (N_21152,N_17782,N_15253);
xnor U21153 (N_21153,N_19760,N_16619);
nor U21154 (N_21154,N_16969,N_16730);
xor U21155 (N_21155,N_16573,N_17899);
and U21156 (N_21156,N_19890,N_15533);
or U21157 (N_21157,N_18821,N_15873);
or U21158 (N_21158,N_19324,N_15489);
xnor U21159 (N_21159,N_17499,N_16267);
nand U21160 (N_21160,N_18443,N_17080);
or U21161 (N_21161,N_18410,N_15305);
and U21162 (N_21162,N_18570,N_19523);
xor U21163 (N_21163,N_17614,N_18226);
and U21164 (N_21164,N_15301,N_19461);
or U21165 (N_21165,N_19166,N_17732);
nor U21166 (N_21166,N_16440,N_17692);
xor U21167 (N_21167,N_15028,N_15994);
or U21168 (N_21168,N_17590,N_18180);
and U21169 (N_21169,N_15874,N_19847);
xnor U21170 (N_21170,N_16476,N_18684);
nand U21171 (N_21171,N_17969,N_17729);
or U21172 (N_21172,N_16054,N_19348);
xor U21173 (N_21173,N_17295,N_18939);
xnor U21174 (N_21174,N_16465,N_17798);
nand U21175 (N_21175,N_19191,N_15637);
and U21176 (N_21176,N_16873,N_19460);
or U21177 (N_21177,N_15534,N_19808);
or U21178 (N_21178,N_15990,N_18136);
nand U21179 (N_21179,N_16534,N_15870);
nor U21180 (N_21180,N_19774,N_19314);
nand U21181 (N_21181,N_18172,N_15437);
nand U21182 (N_21182,N_18803,N_15982);
nor U21183 (N_21183,N_18306,N_19970);
and U21184 (N_21184,N_19334,N_15354);
nor U21185 (N_21185,N_19429,N_16171);
xnor U21186 (N_21186,N_16453,N_15327);
xor U21187 (N_21187,N_19936,N_19580);
and U21188 (N_21188,N_16055,N_19937);
or U21189 (N_21189,N_17076,N_18940);
or U21190 (N_21190,N_17711,N_18081);
nand U21191 (N_21191,N_15698,N_16095);
xor U21192 (N_21192,N_19657,N_19671);
nor U21193 (N_21193,N_18904,N_15529);
or U21194 (N_21194,N_18228,N_17772);
nand U21195 (N_21195,N_19413,N_19820);
nand U21196 (N_21196,N_16518,N_19631);
and U21197 (N_21197,N_17656,N_17936);
nand U21198 (N_21198,N_16113,N_19136);
nor U21199 (N_21199,N_18469,N_16344);
xor U21200 (N_21200,N_18632,N_15362);
or U21201 (N_21201,N_16841,N_19545);
nor U21202 (N_21202,N_19941,N_17974);
nand U21203 (N_21203,N_19531,N_15669);
or U21204 (N_21204,N_17259,N_18762);
or U21205 (N_21205,N_17009,N_18437);
xor U21206 (N_21206,N_15989,N_19973);
and U21207 (N_21207,N_18182,N_19525);
nor U21208 (N_21208,N_15749,N_17708);
nor U21209 (N_21209,N_19592,N_17265);
or U21210 (N_21210,N_16517,N_18054);
and U21211 (N_21211,N_19800,N_18498);
or U21212 (N_21212,N_16968,N_16742);
nor U21213 (N_21213,N_16933,N_16355);
or U21214 (N_21214,N_16688,N_18771);
or U21215 (N_21215,N_18975,N_16195);
and U21216 (N_21216,N_19743,N_16886);
xnor U21217 (N_21217,N_18009,N_18262);
nand U21218 (N_21218,N_16998,N_17103);
nand U21219 (N_21219,N_16781,N_17701);
and U21220 (N_21220,N_16855,N_16085);
nand U21221 (N_21221,N_18462,N_17455);
or U21222 (N_21222,N_17162,N_18969);
or U21223 (N_21223,N_16721,N_18118);
or U21224 (N_21224,N_19549,N_15356);
xnor U21225 (N_21225,N_17264,N_15881);
nor U21226 (N_21226,N_15783,N_15117);
nand U21227 (N_21227,N_16382,N_16932);
nand U21228 (N_21228,N_17159,N_18255);
xnor U21229 (N_21229,N_19225,N_15559);
nor U21230 (N_21230,N_15389,N_19747);
xnor U21231 (N_21231,N_17060,N_16287);
or U21232 (N_21232,N_19035,N_16100);
nor U21233 (N_21233,N_17109,N_18806);
or U21234 (N_21234,N_16229,N_17307);
xor U21235 (N_21235,N_17211,N_18476);
or U21236 (N_21236,N_18540,N_15347);
and U21237 (N_21237,N_19554,N_15083);
or U21238 (N_21238,N_18093,N_18112);
nand U21239 (N_21239,N_15229,N_18510);
nand U21240 (N_21240,N_19203,N_18417);
and U21241 (N_21241,N_19207,N_16439);
and U21242 (N_21242,N_19047,N_15876);
xnor U21243 (N_21243,N_15088,N_16249);
and U21244 (N_21244,N_19994,N_19480);
xor U21245 (N_21245,N_19367,N_16471);
or U21246 (N_21246,N_19376,N_19032);
xnor U21247 (N_21247,N_16245,N_19153);
xnor U21248 (N_21248,N_18576,N_18003);
or U21249 (N_21249,N_18802,N_19686);
xnor U21250 (N_21250,N_15110,N_18022);
or U21251 (N_21251,N_19567,N_17479);
and U21252 (N_21252,N_16941,N_18638);
and U21253 (N_21253,N_16080,N_17704);
nor U21254 (N_21254,N_17527,N_19703);
xor U21255 (N_21255,N_16931,N_16996);
and U21256 (N_21256,N_19029,N_17846);
xnor U21257 (N_21257,N_15217,N_15016);
xnor U21258 (N_21258,N_15643,N_18945);
nor U21259 (N_21259,N_15064,N_19802);
xor U21260 (N_21260,N_16468,N_17275);
or U21261 (N_21261,N_17963,N_17163);
nor U21262 (N_21262,N_15422,N_16010);
or U21263 (N_21263,N_16971,N_15686);
nor U21264 (N_21264,N_18018,N_15979);
and U21265 (N_21265,N_15833,N_19601);
nor U21266 (N_21266,N_18844,N_19145);
xnor U21267 (N_21267,N_16211,N_16079);
or U21268 (N_21268,N_16853,N_16883);
nand U21269 (N_21269,N_16840,N_17758);
xor U21270 (N_21270,N_18909,N_18925);
nor U21271 (N_21271,N_18859,N_15951);
nand U21272 (N_21272,N_18356,N_18198);
nor U21273 (N_21273,N_15001,N_15937);
nor U21274 (N_21274,N_16551,N_18946);
nor U21275 (N_21275,N_19719,N_17249);
or U21276 (N_21276,N_18565,N_18502);
nor U21277 (N_21277,N_16288,N_19003);
and U21278 (N_21278,N_16354,N_17627);
nand U21279 (N_21279,N_19236,N_18727);
and U21280 (N_21280,N_18335,N_19016);
and U21281 (N_21281,N_18266,N_18805);
and U21282 (N_21282,N_16789,N_15609);
or U21283 (N_21283,N_17581,N_19692);
or U21284 (N_21284,N_15584,N_17285);
nand U21285 (N_21285,N_18559,N_18633);
or U21286 (N_21286,N_16219,N_17665);
xor U21287 (N_21287,N_19851,N_15405);
xnor U21288 (N_21288,N_19570,N_19509);
nor U21289 (N_21289,N_17838,N_19857);
and U21290 (N_21290,N_17216,N_18329);
or U21291 (N_21291,N_15459,N_15514);
or U21292 (N_21292,N_15015,N_19227);
nand U21293 (N_21293,N_19011,N_17341);
or U21294 (N_21294,N_18555,N_16618);
xor U21295 (N_21295,N_15284,N_19532);
xnor U21296 (N_21296,N_19459,N_17954);
or U21297 (N_21297,N_16710,N_16597);
nand U21298 (N_21298,N_16369,N_18388);
nor U21299 (N_21299,N_15654,N_15484);
xor U21300 (N_21300,N_16727,N_16127);
nor U21301 (N_21301,N_17597,N_16418);
nor U21302 (N_21302,N_18833,N_16408);
xnor U21303 (N_21303,N_17843,N_15398);
nand U21304 (N_21304,N_16399,N_19764);
nor U21305 (N_21305,N_19211,N_17484);
and U21306 (N_21306,N_18693,N_17916);
and U21307 (N_21307,N_15508,N_16563);
nor U21308 (N_21308,N_19489,N_17083);
or U21309 (N_21309,N_16879,N_19105);
and U21310 (N_21310,N_16908,N_19782);
nor U21311 (N_21311,N_16101,N_16210);
or U21312 (N_21312,N_15743,N_15035);
or U21313 (N_21313,N_15281,N_18027);
nor U21314 (N_21314,N_18907,N_17268);
and U21315 (N_21315,N_16513,N_17928);
nand U21316 (N_21316,N_18562,N_17149);
nand U21317 (N_21317,N_19300,N_16856);
nor U21318 (N_21318,N_19575,N_15111);
or U21319 (N_21319,N_16580,N_17154);
nand U21320 (N_21320,N_18663,N_17854);
nand U21321 (N_21321,N_17893,N_18569);
xnor U21322 (N_21322,N_17819,N_16679);
nand U21323 (N_21323,N_15872,N_16419);
nand U21324 (N_21324,N_15574,N_16795);
xnor U21325 (N_21325,N_15031,N_18509);
nand U21326 (N_21326,N_15653,N_15709);
or U21327 (N_21327,N_18123,N_15053);
nor U21328 (N_21328,N_15731,N_17519);
nor U21329 (N_21329,N_15564,N_15122);
nor U21330 (N_21330,N_15359,N_17389);
nand U21331 (N_21331,N_18706,N_17766);
nor U21332 (N_21332,N_18974,N_16600);
nor U21333 (N_21333,N_16697,N_16980);
or U21334 (N_21334,N_16348,N_16724);
xor U21335 (N_21335,N_17720,N_18665);
and U21336 (N_21336,N_16165,N_17331);
xor U21337 (N_21337,N_15942,N_17811);
xnor U21338 (N_21338,N_19517,N_19271);
xor U21339 (N_21339,N_15741,N_18122);
nand U21340 (N_21340,N_17394,N_16653);
nor U21341 (N_21341,N_17642,N_16238);
or U21342 (N_21342,N_18645,N_18293);
or U21343 (N_21343,N_16814,N_19141);
nor U21344 (N_21344,N_17012,N_18139);
nand U21345 (N_21345,N_19210,N_19397);
and U21346 (N_21346,N_18895,N_16006);
and U21347 (N_21347,N_18885,N_19992);
and U21348 (N_21348,N_18767,N_15196);
nand U21349 (N_21349,N_15688,N_15374);
nor U21350 (N_21350,N_16572,N_17467);
nand U21351 (N_21351,N_19012,N_15848);
or U21352 (N_21352,N_18142,N_15800);
xnor U21353 (N_21353,N_16024,N_19521);
nor U21354 (N_21354,N_15340,N_15727);
and U21355 (N_21355,N_19519,N_16926);
and U21356 (N_21356,N_17575,N_19775);
nor U21357 (N_21357,N_15471,N_17238);
and U21358 (N_21358,N_16048,N_18177);
nor U21359 (N_21359,N_19349,N_19974);
or U21360 (N_21360,N_19984,N_19837);
or U21361 (N_21361,N_16005,N_19894);
nand U21362 (N_21362,N_19598,N_19485);
and U21363 (N_21363,N_16860,N_15900);
nor U21364 (N_21364,N_17797,N_16945);
nand U21365 (N_21365,N_15807,N_15283);
and U21366 (N_21366,N_15004,N_18769);
and U21367 (N_21367,N_18015,N_15949);
or U21368 (N_21368,N_15754,N_16712);
nand U21369 (N_21369,N_15057,N_18937);
nand U21370 (N_21370,N_17497,N_16583);
nor U21371 (N_21371,N_15869,N_18379);
nor U21372 (N_21372,N_17093,N_19263);
nor U21373 (N_21373,N_17113,N_16273);
or U21374 (N_21374,N_16090,N_17507);
nand U21375 (N_21375,N_17346,N_17199);
nor U21376 (N_21376,N_19632,N_19400);
or U21377 (N_21377,N_15034,N_15889);
xnor U21378 (N_21378,N_17308,N_17613);
and U21379 (N_21379,N_15216,N_15187);
and U21380 (N_21380,N_18584,N_19942);
nor U21381 (N_21381,N_19484,N_15886);
nand U21382 (N_21382,N_19290,N_18778);
and U21383 (N_21383,N_16167,N_15650);
xnor U21384 (N_21384,N_18865,N_15704);
xor U21385 (N_21385,N_17637,N_16570);
nand U21386 (N_21386,N_15735,N_16554);
nand U21387 (N_21387,N_15027,N_15538);
nand U21388 (N_21388,N_17986,N_16567);
xor U21389 (N_21389,N_18877,N_18244);
nor U21390 (N_21390,N_18689,N_15948);
or U21391 (N_21391,N_19305,N_15719);
or U21392 (N_21392,N_16110,N_17473);
or U21393 (N_21393,N_18782,N_16838);
and U21394 (N_21394,N_16691,N_19350);
nand U21395 (N_21395,N_15070,N_16201);
nand U21396 (N_21396,N_18866,N_15357);
or U21397 (N_21397,N_15792,N_15333);
xnor U21398 (N_21398,N_15928,N_16390);
xnor U21399 (N_21399,N_17289,N_19148);
xor U21400 (N_21400,N_18950,N_18784);
nand U21401 (N_21401,N_17632,N_19095);
or U21402 (N_21402,N_16738,N_19721);
and U21403 (N_21403,N_15175,N_19975);
nor U21404 (N_21404,N_16023,N_19079);
and U21405 (N_21405,N_17458,N_17874);
xnor U21406 (N_21406,N_15190,N_17924);
xnor U21407 (N_21407,N_17482,N_16543);
and U21408 (N_21408,N_17533,N_15176);
nor U21409 (N_21409,N_17023,N_15221);
nand U21410 (N_21410,N_18611,N_18605);
and U21411 (N_21411,N_19553,N_19137);
nand U21412 (N_21412,N_19183,N_19500);
nor U21413 (N_21413,N_18830,N_15151);
nor U21414 (N_21414,N_19288,N_17904);
xnor U21415 (N_21415,N_19498,N_16057);
xnor U21416 (N_21416,N_19074,N_16735);
nor U21417 (N_21417,N_18758,N_18669);
nor U21418 (N_21418,N_18983,N_16889);
or U21419 (N_21419,N_18026,N_19338);
nor U21420 (N_21420,N_17930,N_19144);
nor U21421 (N_21421,N_19229,N_17226);
or U21422 (N_21422,N_18320,N_19761);
and U21423 (N_21423,N_17213,N_15636);
xor U21424 (N_21424,N_15093,N_18894);
or U21425 (N_21425,N_15286,N_16431);
and U21426 (N_21426,N_16457,N_18115);
or U21427 (N_21427,N_18987,N_17198);
xor U21428 (N_21428,N_19998,N_19731);
nand U21429 (N_21429,N_19057,N_15483);
and U21430 (N_21430,N_15449,N_17914);
nor U21431 (N_21431,N_16228,N_18071);
and U21432 (N_21432,N_17939,N_15619);
or U21433 (N_21433,N_17311,N_15351);
or U21434 (N_21434,N_16938,N_15905);
nor U21435 (N_21435,N_19770,N_17038);
and U21436 (N_21436,N_17560,N_18503);
nor U21437 (N_21437,N_19045,N_15240);
nor U21438 (N_21438,N_15003,N_15677);
or U21439 (N_21439,N_17585,N_17030);
nor U21440 (N_21440,N_18892,N_19212);
nor U21441 (N_21441,N_18647,N_18489);
and U21442 (N_21442,N_19835,N_19472);
nor U21443 (N_21443,N_19620,N_17823);
nand U21444 (N_21444,N_18685,N_17101);
xor U21445 (N_21445,N_15857,N_18089);
or U21446 (N_21446,N_15955,N_15414);
nor U21447 (N_21447,N_18258,N_17366);
nor U21448 (N_21448,N_15585,N_19381);
nand U21449 (N_21449,N_18902,N_19261);
and U21450 (N_21450,N_15279,N_19142);
nand U21451 (N_21451,N_15597,N_17686);
and U21452 (N_21452,N_19969,N_17741);
nor U21453 (N_21453,N_16052,N_18422);
xnor U21454 (N_21454,N_16232,N_16062);
nor U21455 (N_21455,N_17297,N_19155);
nor U21456 (N_21456,N_19458,N_17114);
nor U21457 (N_21457,N_17480,N_18705);
or U21458 (N_21458,N_16396,N_19454);
or U21459 (N_21459,N_16719,N_15488);
nand U21460 (N_21460,N_18912,N_16901);
or U21461 (N_21461,N_16108,N_16659);
nand U21462 (N_21462,N_17693,N_16156);
and U21463 (N_21463,N_15259,N_18399);
xnor U21464 (N_21464,N_16269,N_18591);
and U21465 (N_21465,N_18722,N_15561);
nand U21466 (N_21466,N_15773,N_17166);
nand U21467 (N_21467,N_16942,N_17645);
xor U21468 (N_21468,N_17459,N_17298);
and U21469 (N_21469,N_18108,N_16185);
and U21470 (N_21470,N_16239,N_16356);
nand U21471 (N_21471,N_18200,N_19384);
xor U21472 (N_21472,N_18577,N_19809);
or U21473 (N_21473,N_16376,N_19678);
xnor U21474 (N_21474,N_17901,N_15113);
and U21475 (N_21475,N_18328,N_15795);
and U21476 (N_21476,N_17894,N_15316);
and U21477 (N_21477,N_19063,N_17478);
or U21478 (N_21478,N_15927,N_16125);
xnor U21479 (N_21479,N_15660,N_16217);
or U21480 (N_21480,N_16722,N_16595);
and U21481 (N_21481,N_19064,N_19540);
and U21482 (N_21482,N_16815,N_19951);
and U21483 (N_21483,N_19558,N_17471);
xor U21484 (N_21484,N_18929,N_18149);
and U21485 (N_21485,N_16130,N_18543);
nor U21486 (N_21486,N_17495,N_17958);
or U21487 (N_21487,N_16244,N_18677);
nor U21488 (N_21488,N_15007,N_18639);
or U21489 (N_21489,N_15041,N_15911);
and U21490 (N_21490,N_19347,N_15375);
or U21491 (N_21491,N_16775,N_18739);
nand U21492 (N_21492,N_17195,N_16698);
nand U21493 (N_21493,N_19655,N_15737);
or U21494 (N_21494,N_17169,N_15467);
nand U21495 (N_21495,N_17906,N_18451);
nor U21496 (N_21496,N_15212,N_17128);
xnor U21497 (N_21497,N_18229,N_15388);
nor U21498 (N_21498,N_18261,N_18194);
nor U21499 (N_21499,N_18024,N_18423);
nand U21500 (N_21500,N_18525,N_16695);
and U21501 (N_21501,N_17369,N_18091);
or U21502 (N_21502,N_17200,N_17756);
nor U21503 (N_21503,N_16365,N_15893);
nor U21504 (N_21504,N_18203,N_19948);
xor U21505 (N_21505,N_17889,N_15010);
nor U21506 (N_21506,N_15393,N_17934);
nand U21507 (N_21507,N_17181,N_15348);
nor U21508 (N_21508,N_17599,N_16617);
and U21509 (N_21509,N_16047,N_19258);
and U21510 (N_21510,N_15736,N_16073);
xnor U21511 (N_21511,N_16502,N_19613);
nor U21512 (N_21512,N_17439,N_16041);
nor U21513 (N_21513,N_16430,N_18187);
and U21514 (N_21514,N_19335,N_15231);
or U21515 (N_21515,N_19399,N_17337);
nor U21516 (N_21516,N_17639,N_18947);
xnor U21517 (N_21517,N_19345,N_15275);
nor U21518 (N_21518,N_16397,N_17997);
or U21519 (N_21519,N_19742,N_15765);
and U21520 (N_21520,N_16978,N_16951);
nand U21521 (N_21521,N_15746,N_19344);
nand U21522 (N_21522,N_15380,N_16778);
or U21523 (N_21523,N_17556,N_15703);
xnor U21524 (N_21524,N_15555,N_17883);
xnor U21525 (N_21525,N_17940,N_18001);
nand U21526 (N_21526,N_19028,N_17554);
xnor U21527 (N_21527,N_17653,N_17858);
or U21528 (N_21528,N_17638,N_15519);
nor U21529 (N_21529,N_15896,N_16133);
xor U21530 (N_21530,N_15138,N_16144);
xnor U21531 (N_21531,N_19315,N_19753);
xnor U21532 (N_21532,N_15033,N_16443);
nor U21533 (N_21533,N_15554,N_17700);
nand U21534 (N_21534,N_17796,N_15981);
and U21535 (N_21535,N_17292,N_19233);
xnor U21536 (N_21536,N_15448,N_19699);
nand U21537 (N_21537,N_15894,N_17296);
nor U21538 (N_21538,N_16077,N_15843);
and U21539 (N_21539,N_17545,N_19186);
or U21540 (N_21540,N_16564,N_16297);
nand U21541 (N_21541,N_17412,N_15269);
xor U21542 (N_21542,N_15652,N_16864);
nor U21543 (N_21543,N_19537,N_17643);
nor U21544 (N_21544,N_17184,N_18099);
nor U21545 (N_21545,N_18490,N_18438);
nor U21546 (N_21546,N_19909,N_15206);
nor U21547 (N_21547,N_18792,N_16910);
xor U21548 (N_21548,N_16086,N_15968);
and U21549 (N_21549,N_18345,N_18181);
nand U21550 (N_21550,N_17816,N_18604);
or U21551 (N_21551,N_16091,N_19959);
xor U21552 (N_21552,N_17014,N_15837);
or U21553 (N_21553,N_19242,N_17146);
nand U21554 (N_21554,N_15866,N_17371);
nand U21555 (N_21555,N_15599,N_15543);
nand U21556 (N_21556,N_15521,N_18277);
nor U21557 (N_21557,N_17902,N_18527);
nor U21558 (N_21558,N_15986,N_15249);
or U21559 (N_21559,N_17358,N_17068);
nor U21560 (N_21560,N_17106,N_15723);
and U21561 (N_21561,N_15462,N_19814);
or U21562 (N_21562,N_17667,N_17800);
nand U21563 (N_21563,N_18287,N_15594);
and U21564 (N_21564,N_15133,N_15684);
or U21565 (N_21565,N_19422,N_18738);
and U21566 (N_21566,N_18891,N_18958);
nand U21567 (N_21567,N_16154,N_16116);
or U21568 (N_21568,N_19976,N_16818);
xor U21569 (N_21569,N_19053,N_17040);
xnor U21570 (N_21570,N_17537,N_15108);
or U21571 (N_21571,N_18471,N_15674);
nand U21572 (N_21572,N_17757,N_17277);
nor U21573 (N_21573,N_18133,N_17138);
nor U21574 (N_21574,N_18649,N_16638);
nor U21575 (N_21575,N_15017,N_15588);
xnor U21576 (N_21576,N_16561,N_17725);
or U21577 (N_21577,N_18274,N_19675);
and U21578 (N_21578,N_19394,N_16394);
nor U21579 (N_21579,N_19493,N_16294);
nand U21580 (N_21580,N_17343,N_15477);
nor U21581 (N_21581,N_19589,N_16191);
or U21582 (N_21582,N_16506,N_16321);
or U21583 (N_21583,N_17707,N_19221);
xnor U21584 (N_21584,N_17534,N_19262);
xor U21585 (N_21585,N_17345,N_15068);
and U21586 (N_21586,N_18426,N_16032);
or U21587 (N_21587,N_16514,N_18166);
xor U21588 (N_21588,N_15350,N_16308);
and U21589 (N_21589,N_17316,N_16973);
or U21590 (N_21590,N_16395,N_19269);
or U21591 (N_21591,N_19320,N_17230);
nand U21592 (N_21592,N_16634,N_16628);
xor U21593 (N_21593,N_18193,N_18246);
and U21594 (N_21594,N_17807,N_19605);
nor U21595 (N_21595,N_16888,N_15983);
nor U21596 (N_21596,N_18571,N_19766);
or U21597 (N_21597,N_18781,N_16658);
xor U21598 (N_21598,N_19905,N_18588);
nand U21599 (N_21599,N_15446,N_19860);
nand U21600 (N_21600,N_19804,N_18816);
xnor U21601 (N_21601,N_18216,N_19982);
nand U21602 (N_21602,N_19096,N_17522);
or U21603 (N_21603,N_19388,N_15002);
nand U21604 (N_21604,N_18748,N_18272);
and U21605 (N_21605,N_18360,N_16173);
nand U21606 (N_21606,N_19673,N_18607);
nor U21607 (N_21607,N_18916,N_15370);
nor U21608 (N_21608,N_17115,N_18720);
xnor U21609 (N_21609,N_19539,N_16777);
nor U21610 (N_21610,N_19790,N_19563);
or U21611 (N_21611,N_18794,N_19848);
nor U21612 (N_21612,N_15756,N_15504);
or U21613 (N_21613,N_17791,N_18701);
or U21614 (N_21614,N_18252,N_15260);
or U21615 (N_21615,N_17445,N_18629);
or U21616 (N_21616,N_19200,N_15779);
nand U21617 (N_21617,N_15037,N_16081);
nor U21618 (N_21618,N_16606,N_15054);
xnor U21619 (N_21619,N_18151,N_16794);
nor U21620 (N_21620,N_15708,N_16575);
nand U21621 (N_21621,N_16258,N_18724);
or U21622 (N_21622,N_16966,N_17546);
nor U21623 (N_21623,N_15823,N_19634);
nor U21624 (N_21624,N_15626,N_17770);
nor U21625 (N_21625,N_16703,N_16019);
nor U21626 (N_21626,N_19755,N_19960);
and U21627 (N_21627,N_16008,N_16977);
or U21628 (N_21628,N_17313,N_19989);
nand U21629 (N_21629,N_16179,N_18707);
xnor U21630 (N_21630,N_19781,N_19779);
nor U21631 (N_21631,N_19436,N_16183);
and U21632 (N_21632,N_15468,N_15345);
or U21633 (N_21633,N_16608,N_16076);
or U21634 (N_21634,N_18060,N_15836);
xnor U21635 (N_21635,N_18442,N_16770);
or U21636 (N_21636,N_18615,N_18995);
nor U21637 (N_21637,N_18330,N_17920);
nand U21638 (N_21638,N_15174,N_18934);
and U21639 (N_21639,N_19463,N_17619);
and U21640 (N_21640,N_16407,N_18704);
and U21641 (N_21641,N_16410,N_19688);
nand U21642 (N_21642,N_18282,N_18464);
nor U21643 (N_21643,N_18135,N_18348);
and U21644 (N_21644,N_18002,N_15815);
and U21645 (N_21645,N_18729,N_18624);
xor U21646 (N_21646,N_19587,N_17754);
nor U21647 (N_21647,N_17764,N_16153);
nand U21648 (N_21648,N_18501,N_15680);
and U21649 (N_21649,N_18041,N_19445);
xnor U21650 (N_21650,N_16188,N_18817);
nand U21651 (N_21651,N_18121,N_19282);
or U21652 (N_21652,N_16470,N_18304);
xnor U21653 (N_21653,N_18400,N_18641);
nand U21654 (N_21654,N_19372,N_17789);
xor U21655 (N_21655,N_17339,N_15852);
nand U21656 (N_21656,N_19161,N_18375);
nand U21657 (N_21657,N_19059,N_18813);
or U21658 (N_21658,N_19928,N_19556);
xnor U21659 (N_21659,N_15116,N_15451);
xnor U21660 (N_21660,N_18926,N_16438);
nand U21661 (N_21661,N_17256,N_16602);
and U21662 (N_21662,N_16069,N_17270);
or U21663 (N_21663,N_18381,N_19453);
or U21664 (N_21664,N_16648,N_16565);
or U21665 (N_21665,N_16000,N_16820);
xnor U21666 (N_21666,N_18505,N_18369);
nor U21667 (N_21667,N_18219,N_15936);
or U21668 (N_21668,N_18873,N_15687);
nor U21669 (N_21669,N_16371,N_19746);
nor U21670 (N_21670,N_19494,N_19816);
and U21671 (N_21671,N_18927,N_19169);
xnor U21672 (N_21672,N_19871,N_18522);
nor U21673 (N_21673,N_17820,N_19912);
xnor U21674 (N_21674,N_18592,N_16182);
or U21675 (N_21675,N_18646,N_17690);
nor U21676 (N_21676,N_17931,N_17416);
xnor U21677 (N_21677,N_17847,N_18387);
nor U21678 (N_21678,N_18007,N_18049);
nor U21679 (N_21679,N_15977,N_18538);
xor U21680 (N_21680,N_16484,N_16251);
or U21681 (N_21681,N_18823,N_18921);
xnor U21682 (N_21682,N_16592,N_18911);
nand U21683 (N_21683,N_17286,N_18362);
nor U21684 (N_21684,N_18189,N_18938);
nor U21685 (N_21685,N_17004,N_17335);
nor U21686 (N_21686,N_17406,N_19696);
nor U21687 (N_21687,N_17155,N_15302);
and U21688 (N_21688,N_19365,N_16449);
nand U21689 (N_21689,N_16717,N_16446);
nor U21690 (N_21690,N_18468,N_19856);
xor U21691 (N_21691,N_18062,N_17035);
xnor U21692 (N_21692,N_15408,N_17947);
nand U21693 (N_21693,N_16068,N_19173);
and U21694 (N_21694,N_17561,N_16899);
or U21695 (N_21695,N_19966,N_18269);
or U21696 (N_21696,N_19867,N_17383);
or U21697 (N_21697,N_15419,N_15811);
and U21698 (N_21698,N_15089,N_16292);
and U21699 (N_21699,N_15094,N_19503);
or U21700 (N_21700,N_16637,N_19013);
nor U21701 (N_21701,N_17825,N_16114);
or U21702 (N_21702,N_16367,N_19428);
nor U21703 (N_21703,N_17257,N_18996);
nand U21704 (N_21704,N_16805,N_16892);
nor U21705 (N_21705,N_16959,N_17212);
or U21706 (N_21706,N_15139,N_15917);
or U21707 (N_21707,N_17822,N_15601);
or U21708 (N_21708,N_19071,N_19997);
and U21709 (N_21709,N_16038,N_18898);
xnor U21710 (N_21710,N_18694,N_16254);
and U21711 (N_21711,N_15025,N_18879);
nand U21712 (N_21712,N_19759,N_16929);
or U21713 (N_21713,N_17518,N_15998);
or U21714 (N_21714,N_15914,N_15278);
nor U21715 (N_21715,N_15633,N_19943);
nor U21716 (N_21716,N_16178,N_18618);
and U21717 (N_21717,N_16831,N_15219);
xnor U21718 (N_21718,N_19918,N_17391);
nand U21719 (N_21719,N_15082,N_17175);
nor U21720 (N_21720,N_18236,N_17587);
nand U21721 (N_21721,N_19522,N_18327);
nor U21722 (N_21722,N_19963,N_15244);
xnor U21723 (N_21723,N_19339,N_17380);
and U21724 (N_21724,N_18673,N_15557);
and U21725 (N_21725,N_18560,N_17167);
nor U21726 (N_21726,N_18061,N_17833);
nor U21727 (N_21727,N_18997,N_19215);
xor U21728 (N_21728,N_17676,N_18799);
xnor U21729 (N_21729,N_16995,N_15810);
xor U21730 (N_21730,N_15298,N_16207);
nand U21731 (N_21731,N_17125,N_17862);
and U21732 (N_21732,N_16289,N_19002);
or U21733 (N_21733,N_16463,N_19922);
nand U21734 (N_21734,N_17081,N_16247);
nand U21735 (N_21735,N_17622,N_16983);
or U21736 (N_21736,N_15426,N_19327);
nand U21737 (N_21737,N_19115,N_16904);
and U21738 (N_21738,N_19795,N_18523);
or U21739 (N_21739,N_16651,N_18980);
nand U21740 (N_21740,N_18764,N_17354);
and U21741 (N_21741,N_17571,N_19108);
and U21742 (N_21742,N_16084,N_15280);
or U21743 (N_21743,N_18787,N_18331);
nor U21744 (N_21744,N_19134,N_15902);
and U21745 (N_21745,N_15314,N_18005);
nand U21746 (N_21746,N_19754,N_19255);
nand U21747 (N_21747,N_17209,N_16747);
and U21748 (N_21748,N_17075,N_16550);
nand U21749 (N_21749,N_19505,N_19373);
and U21750 (N_21750,N_17043,N_17381);
nor U21751 (N_21751,N_16189,N_19272);
and U21752 (N_21752,N_16813,N_15250);
and U21753 (N_21753,N_15330,N_19810);
xor U21754 (N_21754,N_16863,N_17654);
or U21755 (N_21755,N_18506,N_18162);
xor U21756 (N_21756,N_16558,N_18756);
or U21757 (N_21757,N_17293,N_17880);
and U21758 (N_21758,N_18826,N_18039);
nand U21759 (N_21759,N_18076,N_18299);
xor U21760 (N_21760,N_15474,N_19639);
or U21761 (N_21761,N_15159,N_19332);
and U21762 (N_21762,N_17141,N_18575);
xor U21763 (N_21763,N_17714,N_18621);
and U21764 (N_21764,N_19414,N_18023);
nor U21765 (N_21765,N_19911,N_19821);
nor U21766 (N_21766,N_17271,N_15100);
xor U21767 (N_21767,N_18265,N_19222);
nand U21768 (N_21768,N_17780,N_17837);
nor U21769 (N_21769,N_16334,N_16799);
and U21770 (N_21770,N_17172,N_15845);
or U21771 (N_21771,N_16159,N_16584);
and U21772 (N_21772,N_16271,N_17327);
xor U21773 (N_21773,N_19420,N_19009);
xnor U21774 (N_21774,N_17640,N_16213);
xor U21775 (N_21775,N_15734,N_15381);
nand U21776 (N_21776,N_17386,N_19822);
nand U21777 (N_21777,N_16033,N_18152);
nor U21778 (N_21778,N_18699,N_15406);
or U21779 (N_21779,N_18721,N_16034);
nand U21780 (N_21780,N_16495,N_18334);
or U21781 (N_21781,N_19008,N_15944);
nand U21782 (N_21782,N_19700,N_15915);
nand U21783 (N_21783,N_17047,N_17602);
xnor U21784 (N_21784,N_16545,N_15215);
xnor U21785 (N_21785,N_19259,N_17508);
xnor U21786 (N_21786,N_18404,N_15328);
xor U21787 (N_21787,N_16063,N_16552);
and U21788 (N_21788,N_16452,N_16902);
xor U21789 (N_21789,N_16362,N_19798);
nor U21790 (N_21790,N_15160,N_18583);
or U21791 (N_21791,N_18648,N_15479);
nor U21792 (N_21792,N_18013,N_19366);
nand U21793 (N_21793,N_15416,N_18249);
or U21794 (N_21794,N_17045,N_19910);
xnor U21795 (N_21795,N_19432,N_18931);
xor U21796 (N_21796,N_16283,N_17245);
or U21797 (N_21797,N_16832,N_17513);
or U21798 (N_21798,N_16466,N_19864);
and U21799 (N_21799,N_17370,N_18077);
nor U21800 (N_21800,N_15143,N_16414);
nand U21801 (N_21801,N_17821,N_19796);
nand U21802 (N_21802,N_17183,N_15226);
nand U21803 (N_21803,N_19054,N_18541);
nor U21804 (N_21804,N_16037,N_17215);
and U21805 (N_21805,N_19908,N_18344);
and U21806 (N_21806,N_18202,N_15947);
and U21807 (N_21807,N_17440,N_18128);
nor U21808 (N_21808,N_16204,N_15262);
nor U21809 (N_21809,N_15784,N_17258);
or U21810 (N_21810,N_15868,N_16458);
and U21811 (N_21811,N_19195,N_17689);
and U21812 (N_21812,N_18100,N_15964);
nand U21813 (N_21813,N_16264,N_19291);
and U21814 (N_21814,N_15689,N_15104);
or U21815 (N_21815,N_17419,N_19325);
xor U21816 (N_21816,N_19351,N_19612);
and U21817 (N_21817,N_18928,N_19086);
and U21818 (N_21818,N_15456,N_16400);
nand U21819 (N_21819,N_18378,N_19356);
xnor U21820 (N_21820,N_17442,N_18019);
nor U21821 (N_21821,N_18536,N_16087);
nand U21822 (N_21822,N_19879,N_19752);
and U21823 (N_21823,N_18622,N_16401);
and U21824 (N_21824,N_18791,N_18210);
and U21825 (N_21825,N_15987,N_16757);
xnor U21826 (N_21826,N_15401,N_19983);
nand U21827 (N_21827,N_17589,N_18545);
or U21828 (N_21828,N_15091,N_19658);
xnor U21829 (N_21829,N_19280,N_18666);
and U21830 (N_21830,N_18051,N_15272);
nand U21831 (N_21831,N_17002,N_16286);
nor U21832 (N_21832,N_15863,N_16733);
xnor U21833 (N_21833,N_19709,N_17830);
and U21834 (N_21834,N_15140,N_19421);
nand U21835 (N_21835,N_17773,N_17413);
or U21836 (N_21836,N_18708,N_19426);
and U21837 (N_21837,N_18377,N_16515);
nand U21838 (N_21838,N_18617,N_19733);
xor U21839 (N_21839,N_18913,N_17606);
or U21840 (N_21840,N_18836,N_19304);
or U21841 (N_21841,N_19962,N_19163);
nand U21842 (N_21842,N_18740,N_16960);
nor U21843 (N_21843,N_16896,N_16720);
nor U21844 (N_21844,N_18563,N_18537);
nor U21845 (N_21845,N_16660,N_17870);
nand U21846 (N_21846,N_18657,N_19687);
nor U21847 (N_21847,N_16965,N_15378);
or U21848 (N_21848,N_16522,N_16097);
and U21849 (N_21849,N_16242,N_16309);
nor U21850 (N_21850,N_18789,N_18551);
nand U21851 (N_21851,N_16233,N_19019);
nand U21852 (N_21852,N_15923,N_17034);
nand U21853 (N_21853,N_18132,N_17287);
xnor U21854 (N_21854,N_17779,N_19777);
nand U21855 (N_21855,N_15760,N_17900);
xor U21856 (N_21856,N_16082,N_18688);
or U21857 (N_21857,N_17283,N_17705);
xnor U21858 (N_21858,N_15572,N_18053);
nor U21859 (N_21859,N_18655,N_16909);
xor U21860 (N_21860,N_19689,N_18948);
nor U21861 (N_21861,N_17814,N_18933);
xnor U21862 (N_21862,N_15325,N_15397);
xor U21863 (N_21863,N_18279,N_15864);
nor U21864 (N_21864,N_15910,N_17923);
nand U21865 (N_21865,N_19044,N_19546);
xor U21866 (N_21866,N_19865,N_19398);
nand U21867 (N_21867,N_17025,N_16206);
nor U21868 (N_21868,N_16961,N_15166);
and U21869 (N_21869,N_15946,N_19710);
xor U21870 (N_21870,N_16268,N_15008);
nand U21871 (N_21871,N_19728,N_19651);
nor U21872 (N_21872,N_15625,N_17926);
and U21873 (N_21873,N_16501,N_17890);
and U21874 (N_21874,N_18309,N_16954);
or U21875 (N_21875,N_18757,N_17055);
nor U21876 (N_21876,N_17549,N_18284);
or U21877 (N_21877,N_18698,N_18070);
or U21878 (N_21878,N_18603,N_15197);
xnor U21879 (N_21879,N_16750,N_17039);
and U21880 (N_21880,N_15101,N_15850);
or U21881 (N_21881,N_15178,N_16028);
xor U21882 (N_21882,N_17817,N_16921);
or U21883 (N_21883,N_17470,N_18675);
nor U21884 (N_21884,N_19797,N_18932);
or U21885 (N_21885,N_15346,N_15632);
nor U21886 (N_21886,N_16508,N_19507);
and U21887 (N_21887,N_15069,N_16881);
xor U21888 (N_21888,N_17876,N_17786);
nor U21889 (N_21889,N_17102,N_18535);
or U21890 (N_21890,N_15540,N_18943);
and U21891 (N_21891,N_15493,N_17695);
nand U21892 (N_21892,N_16668,N_19946);
or U21893 (N_21893,N_16631,N_18849);
and U21894 (N_21894,N_15400,N_16844);
nor U21895 (N_21895,N_16472,N_18674);
and U21896 (N_21896,N_15336,N_15602);
and U21897 (N_21897,N_18890,N_17005);
nor U21898 (N_21898,N_16944,N_18033);
or U21899 (N_21899,N_17655,N_18418);
nand U21900 (N_21900,N_19945,N_19274);
xor U21901 (N_21901,N_16012,N_19653);
or U21902 (N_21902,N_16884,N_17281);
xnor U21903 (N_21903,N_19010,N_16623);
nand U21904 (N_21904,N_19635,N_17129);
and U21905 (N_21905,N_15630,N_17550);
and U21906 (N_21906,N_16282,N_15447);
and U21907 (N_21907,N_19885,N_17675);
nor U21908 (N_21908,N_19818,N_17611);
or U21909 (N_21909,N_15844,N_16231);
nand U21910 (N_21910,N_16423,N_16363);
xor U21911 (N_21911,N_19219,N_19887);
nand U21912 (N_21912,N_18755,N_16768);
and U21913 (N_21913,N_15154,N_15501);
and U21914 (N_21914,N_17943,N_18961);
nor U21915 (N_21915,N_17652,N_19146);
and U21916 (N_21916,N_19940,N_15285);
and U21917 (N_21917,N_16621,N_15355);
nor U21918 (N_21918,N_19904,N_18951);
or U21919 (N_21919,N_18893,N_19292);
nand U21920 (N_21920,N_18809,N_17424);
or U21921 (N_21921,N_17520,N_16290);
or U21922 (N_21922,N_19475,N_16504);
nand U21923 (N_21923,N_15074,N_19780);
and U21924 (N_21924,N_15929,N_19427);
and U21925 (N_21925,N_15816,N_19135);
xnor U21926 (N_21926,N_16812,N_19901);
nand U21927 (N_21927,N_15148,N_19884);
and U21928 (N_21928,N_18766,N_16643);
and U21929 (N_21929,N_19723,N_19771);
and U21930 (N_21930,N_19329,N_18432);
or U21931 (N_21931,N_18028,N_19130);
or U21932 (N_21932,N_19065,N_16655);
nand U21933 (N_21933,N_19736,N_15976);
and U21934 (N_21934,N_16707,N_15551);
or U21935 (N_21935,N_16050,N_19866);
nor U21936 (N_21936,N_16705,N_17514);
and U21937 (N_21937,N_17750,N_19588);
and U21938 (N_21938,N_18352,N_15161);
or U21939 (N_21939,N_16527,N_15364);
and U21940 (N_21940,N_15156,N_17875);
or U21941 (N_21941,N_17968,N_16491);
and U21942 (N_21942,N_17747,N_17260);
or U21943 (N_21943,N_19178,N_16387);
nor U21944 (N_21944,N_19680,N_17873);
nand U21945 (N_21945,N_16627,N_17448);
xor U21946 (N_21946,N_16509,N_16685);
nand U21947 (N_21947,N_19630,N_16174);
nor U21948 (N_21948,N_18147,N_15440);
nor U21949 (N_21949,N_17525,N_19479);
and U21950 (N_21950,N_16765,N_15344);
xnor U21951 (N_21951,N_15102,N_19231);
xnor U21952 (N_21952,N_19652,N_17160);
nand U21953 (N_21953,N_17131,N_17332);
nand U21954 (N_21954,N_18596,N_16202);
and U21955 (N_21955,N_15105,N_17373);
and U21956 (N_21956,N_17329,N_18212);
or U21957 (N_21957,N_19337,N_15676);
nor U21958 (N_21958,N_17765,N_15465);
xor U21959 (N_21959,N_16460,N_19571);
xor U21960 (N_21960,N_17907,N_18744);
nor U21961 (N_21961,N_18901,N_15805);
xor U21962 (N_21962,N_19473,N_17918);
xnor U21963 (N_21963,N_19312,N_17379);
nor U21964 (N_21964,N_19576,N_17681);
nor U21965 (N_21965,N_18512,N_18814);
nor U21966 (N_21966,N_15470,N_15527);
nand U21967 (N_21967,N_19708,N_16124);
nand U21968 (N_21968,N_15532,N_19640);
nor U21969 (N_21969,N_15498,N_16096);
nor U21970 (N_21970,N_15701,N_16067);
and U21971 (N_21971,N_19987,N_17661);
nor U21972 (N_21972,N_18820,N_19520);
xnor U21973 (N_21973,N_18495,N_15230);
and U21974 (N_21974,N_15332,N_16049);
xor U21975 (N_21975,N_16317,N_18042);
xnor U21976 (N_21976,N_19799,N_18986);
xor U21977 (N_21977,N_18862,N_17116);
or U21978 (N_21978,N_17584,N_17739);
or U21979 (N_21979,N_17500,N_16152);
or U21980 (N_21980,N_19478,N_17205);
and U21981 (N_21981,N_17089,N_15662);
xnor U21982 (N_21982,N_18314,N_15181);
and U21983 (N_21983,N_15738,N_19077);
nor U21984 (N_21984,N_16409,N_19014);
or U21985 (N_21985,N_19602,N_19533);
nand U21986 (N_21986,N_16934,N_15618);
nor U21987 (N_21987,N_19464,N_16740);
or U21988 (N_21988,N_17839,N_16533);
or U21989 (N_21989,N_18735,N_16039);
or U21990 (N_21990,N_19502,N_17670);
xor U21991 (N_21991,N_17062,N_18167);
and U21992 (N_21992,N_16014,N_15525);
and U21993 (N_21993,N_16357,N_16436);
xnor U21994 (N_21994,N_19352,N_18197);
xnor U21995 (N_21995,N_18316,N_17073);
nand U21996 (N_21996,N_19039,N_19067);
xnor U21997 (N_21997,N_16374,N_19270);
or U21998 (N_21998,N_17029,N_15263);
and U21999 (N_21999,N_16986,N_18351);
and U22000 (N_22000,N_15339,N_17309);
or U22001 (N_22001,N_18439,N_18461);
or U22002 (N_22002,N_16981,N_17878);
or U22003 (N_22003,N_15970,N_15791);
or U22004 (N_22004,N_19610,N_17187);
and U22005 (N_22005,N_15009,N_16214);
xor U22006 (N_22006,N_19060,N_16437);
nand U22007 (N_22007,N_18129,N_15287);
and U22008 (N_22008,N_19512,N_18409);
xnor U22009 (N_22009,N_15049,N_18960);
nand U22010 (N_22010,N_18874,N_16723);
nand U22011 (N_22011,N_16716,N_17718);
nand U22012 (N_22012,N_19395,N_17566);
xor U22013 (N_22013,N_15413,N_19217);
or U22014 (N_22014,N_15605,N_18680);
or U22015 (N_22015,N_18776,N_16615);
or U22016 (N_22016,N_19331,N_17540);
xnor U22017 (N_22017,N_16456,N_18206);
nor U22018 (N_22018,N_16972,N_16497);
nand U22019 (N_22019,N_18222,N_17176);
nand U22020 (N_22020,N_19990,N_16391);
or U22021 (N_22021,N_15207,N_19756);
xnor U22022 (N_22022,N_15785,N_18500);
nand U22023 (N_22023,N_15606,N_16295);
or U22024 (N_22024,N_15326,N_18403);
nor U22025 (N_22025,N_17621,N_18544);
or U22026 (N_22026,N_19441,N_15586);
or U22027 (N_22027,N_16579,N_17021);
or U22028 (N_22028,N_19068,N_18743);
and U22029 (N_22029,N_18174,N_15030);
and U22030 (N_22030,N_19591,N_18143);
xnor U22031 (N_22031,N_19526,N_19996);
and U22032 (N_22032,N_16225,N_18140);
nand U22033 (N_22033,N_16531,N_17460);
xor U22034 (N_22034,N_18531,N_17333);
or U22035 (N_22035,N_17868,N_19477);
xor U22036 (N_22036,N_18273,N_18259);
and U22037 (N_22037,N_15430,N_17860);
or U22038 (N_22038,N_19050,N_17828);
nor U22039 (N_22039,N_16599,N_15898);
or U22040 (N_22040,N_16346,N_16335);
nand U22041 (N_22041,N_15507,N_15308);
nor U22042 (N_22042,N_17624,N_18858);
nand U22043 (N_22043,N_18875,N_16455);
xor U22044 (N_22044,N_16279,N_18191);
nor U22045 (N_22045,N_16704,N_17633);
or U22046 (N_22046,N_19196,N_18888);
and U22047 (N_22047,N_17591,N_16758);
xor U22048 (N_22048,N_18384,N_19268);
or U22049 (N_22049,N_15699,N_16895);
or U22050 (N_22050,N_18325,N_19882);
nand U22051 (N_22051,N_15163,N_18339);
nand U22052 (N_22052,N_17428,N_16336);
or U22053 (N_22053,N_17399,N_18910);
xnor U22054 (N_22054,N_18401,N_19663);
or U22055 (N_22055,N_15124,N_16830);
nor U22056 (N_22056,N_19301,N_15168);
and U22057 (N_22057,N_15349,N_17541);
and U22058 (N_22058,N_15123,N_16404);
nor U22059 (N_22059,N_19156,N_16166);
xor U22060 (N_22060,N_16894,N_16118);
nor U22061 (N_22061,N_17836,N_15956);
and U22062 (N_22062,N_15616,N_16848);
nand U22063 (N_22063,N_19977,N_17110);
nor U22064 (N_22064,N_18447,N_16610);
nand U22065 (N_22065,N_18150,N_18779);
nand U22066 (N_22066,N_16875,N_18058);
xor U22067 (N_22067,N_17576,N_15722);
nand U22068 (N_22068,N_15177,N_17999);
nand U22069 (N_22069,N_16291,N_18954);
xnor U22070 (N_22070,N_18930,N_16913);
and U22071 (N_22071,N_16927,N_17494);
nor U22072 (N_22072,N_18572,N_16576);
nor U22073 (N_22073,N_15461,N_17573);
nor U22074 (N_22074,N_19297,N_15668);
nor U22075 (N_22075,N_18192,N_18917);
and U22076 (N_22076,N_16871,N_16642);
and U22077 (N_22077,N_18188,N_18668);
or U22078 (N_22078,N_19457,N_16164);
xor U22079 (N_22079,N_15261,N_15257);
xnor U22080 (N_22080,N_19528,N_18283);
nor U22081 (N_22081,N_19298,N_17241);
and U22082 (N_22082,N_16979,N_15855);
and U22083 (N_22083,N_19396,N_15838);
nand U22084 (N_22084,N_19078,N_15019);
xnor U22085 (N_22085,N_17979,N_19465);
nor U22086 (N_22086,N_15871,N_19954);
or U22087 (N_22087,N_17804,N_15245);
nor U22088 (N_22088,N_15623,N_19438);
and U22089 (N_22089,N_17079,N_15387);
or U22090 (N_22090,N_17887,N_15907);
and U22091 (N_22091,N_19058,N_15144);
or U22092 (N_22092,N_15266,N_15972);
nand U22093 (N_22093,N_18213,N_16313);
or U22094 (N_22094,N_16488,N_19404);
or U22095 (N_22095,N_19030,N_19737);
nand U22096 (N_22096,N_17477,N_15306);
xnor U22097 (N_22097,N_19730,N_16422);
and U22098 (N_22098,N_19826,N_17444);
nand U22099 (N_22099,N_15198,N_17984);
and U22100 (N_22100,N_19544,N_19701);
nand U22101 (N_22101,N_19758,N_15021);
or U22102 (N_22102,N_19246,N_15371);
xnor U22103 (N_22103,N_15026,N_19392);
and U22104 (N_22104,N_19360,N_18207);
nor U22105 (N_22105,N_16020,N_17579);
xor U22106 (N_22106,N_17746,N_18785);
or U22107 (N_22107,N_18982,N_18311);
nand U22108 (N_22108,N_19116,N_15403);
xnor U22109 (N_22109,N_15267,N_17422);
nor U22110 (N_22110,N_17186,N_17950);
and U22111 (N_22111,N_17084,N_15711);
xnor U22112 (N_22112,N_18161,N_16661);
and U22113 (N_22113,N_16345,N_19862);
nor U22114 (N_22114,N_16793,N_16059);
or U22115 (N_22115,N_15300,N_19249);
nor U22116 (N_22116,N_18812,N_18318);
xor U22117 (N_22117,N_16525,N_16711);
or U22118 (N_22118,N_18263,N_17767);
xnor U22119 (N_22119,N_16198,N_15778);
and U22120 (N_22120,N_18424,N_19898);
xor U22121 (N_22121,N_15242,N_18860);
or U22122 (N_22122,N_15218,N_19467);
or U22123 (N_22123,N_17680,N_15563);
xnor U22124 (N_22124,N_15450,N_16647);
nor U22125 (N_22125,N_18797,N_16333);
or U22126 (N_22126,N_17866,N_16358);
nor U22127 (N_22127,N_17074,N_18884);
or U22128 (N_22128,N_16441,N_17964);
or U22129 (N_22129,N_19674,N_19899);
xor U22130 (N_22130,N_16571,N_18078);
nor U22131 (N_22131,N_15999,N_16678);
or U22132 (N_22132,N_19788,N_15912);
nor U22133 (N_22133,N_18046,N_17044);
xnor U22134 (N_22134,N_18686,N_15050);
or U22135 (N_22135,N_18223,N_18183);
xnor U22136 (N_22136,N_18828,N_19088);
and U22137 (N_22137,N_15343,N_15204);
and U22138 (N_22138,N_16915,N_17272);
nand U22139 (N_22139,N_18104,N_18856);
nor U22140 (N_22140,N_18303,N_18195);
and U22141 (N_22141,N_16825,N_17266);
nand U22142 (N_22142,N_18696,N_16708);
and U22143 (N_22143,N_18746,N_18741);
and U22144 (N_22144,N_16800,N_15210);
or U22145 (N_22145,N_15162,N_16329);
and U22146 (N_22146,N_17712,N_16796);
nand U22147 (N_22147,N_17229,N_16256);
xor U22148 (N_22148,N_16923,N_16547);
nand U22149 (N_22149,N_16128,N_18317);
or U22150 (N_22150,N_17050,N_19114);
xnor U22151 (N_22151,N_17189,N_17161);
nand U22152 (N_22152,N_19276,N_15607);
nor U22153 (N_22153,N_19577,N_15851);
xor U22154 (N_22154,N_15774,N_17849);
nor U22155 (N_22155,N_19913,N_15825);
xor U22156 (N_22156,N_17809,N_15369);
and U22157 (N_22157,N_18998,N_16700);
and U22158 (N_22158,N_15486,N_19193);
nor U22159 (N_22159,N_17053,N_16461);
xnor U22160 (N_22160,N_15523,N_16851);
nor U22161 (N_22161,N_16098,N_17760);
nor U22162 (N_22162,N_17636,N_19189);
or U22163 (N_22163,N_19840,N_16607);
or U22164 (N_22164,N_19449,N_18088);
or U22165 (N_22165,N_19103,N_15826);
xnor U22166 (N_22166,N_16310,N_16486);
and U22167 (N_22167,N_15310,N_17781);
or U22168 (N_22168,N_15065,N_18446);
or U22169 (N_22169,N_15706,N_19174);
or U22170 (N_22170,N_19265,N_15992);
nor U22171 (N_22171,N_15814,N_16752);
or U22172 (N_22172,N_18831,N_15954);
nand U22173 (N_22173,N_17864,N_19846);
xnor U22174 (N_22174,N_15726,N_17996);
nand U22175 (N_22175,N_16180,N_17790);
xor U22176 (N_22176,N_15211,N_18759);
nand U22177 (N_22177,N_18586,N_15503);
or U22178 (N_22178,N_18768,N_15020);
nand U22179 (N_22179,N_17884,N_16949);
or U22180 (N_22180,N_18052,N_16654);
and U22181 (N_22181,N_15935,N_16499);
xor U22182 (N_22182,N_19757,N_15980);
and U22183 (N_22183,N_18854,N_18957);
xor U22184 (N_22184,N_16155,N_18494);
nor U22185 (N_22185,N_18990,N_17058);
nor U22186 (N_22186,N_15802,N_17664);
and U22187 (N_22187,N_17957,N_15621);
nand U22188 (N_22188,N_16885,N_18324);
nor U22189 (N_22189,N_16585,N_19603);
or U22190 (N_22190,N_16692,N_15663);
or U22191 (N_22191,N_19256,N_16666);
and U22192 (N_22192,N_16836,N_18661);
and U22193 (N_22193,N_17314,N_15769);
nor U22194 (N_22194,N_18016,N_19443);
nand U22195 (N_22195,N_15875,N_15803);
xor U22196 (N_22196,N_19410,N_19964);
nor U22197 (N_22197,N_15153,N_16035);
nand U22198 (N_22198,N_17173,N_19446);
or U22199 (N_22199,N_19725,N_19813);
nor U22200 (N_22200,N_19845,N_19294);
and U22201 (N_22201,N_15323,N_15548);
and U22202 (N_22202,N_17871,N_18697);
nand U22203 (N_22203,N_18651,N_15638);
xor U22204 (N_22204,N_18719,N_19784);
nor U22205 (N_22205,N_17529,N_16689);
nor U22206 (N_22206,N_19815,N_18763);
nand U22207 (N_22207,N_18011,N_18855);
xor U22208 (N_22208,N_18567,N_18389);
nor U22209 (N_22209,N_19965,N_17082);
and U22210 (N_22210,N_19228,N_15849);
and U22211 (N_22211,N_16341,N_19834);
nand U22212 (N_22212,N_16861,N_16492);
or U22213 (N_22213,N_19386,N_15862);
nor U22214 (N_22214,N_15277,N_16586);
xnor U22215 (N_22215,N_15052,N_17117);
or U22216 (N_22216,N_18095,N_15427);
xor U22217 (N_22217,N_16040,N_19017);
xnor U22218 (N_22218,N_15926,N_17721);
and U22219 (N_22219,N_19027,N_18457);
xnor U22220 (N_22220,N_19993,N_15383);
and U22221 (N_22221,N_19681,N_15822);
or U22222 (N_22222,N_15608,N_18165);
and U22223 (N_22223,N_19581,N_19369);
and U22224 (N_22224,N_15759,N_17338);
and U22225 (N_22225,N_19069,N_15363);
or U22226 (N_22226,N_16577,N_16786);
and U22227 (N_22227,N_16411,N_18985);
xor U22228 (N_22228,N_15185,N_17913);
nand U22229 (N_22229,N_17443,N_16656);
xnor U22230 (N_22230,N_15993,N_17041);
xor U22231 (N_22231,N_16327,N_19046);
or U22232 (N_22232,N_17995,N_19214);
and U22233 (N_22233,N_19018,N_19618);
nand U22234 (N_22234,N_18664,N_16729);
and U22235 (N_22235,N_18590,N_15183);
nor U22236 (N_22236,N_18851,N_15858);
xor U22237 (N_22237,N_16594,N_17108);
nand U22238 (N_22238,N_18280,N_19051);
or U22239 (N_22239,N_17641,N_19037);
nand U22240 (N_22240,N_19455,N_17158);
or U22241 (N_22241,N_17150,N_19633);
nor U22242 (N_22242,N_19364,N_17232);
or U22243 (N_22243,N_16984,N_19481);
nand U22244 (N_22244,N_16783,N_15985);
nor U22245 (N_22245,N_17061,N_17929);
or U22246 (N_22246,N_17649,N_17273);
or U22247 (N_22247,N_18427,N_15506);
and U22248 (N_22248,N_17510,N_19000);
xor U22249 (N_22249,N_17938,N_16236);
or U22250 (N_22250,N_16766,N_16316);
xor U22251 (N_22251,N_16512,N_19491);
nand U22252 (N_22252,N_19495,N_17506);
nor U22253 (N_22253,N_17735,N_17751);
nor U22254 (N_22254,N_19677,N_17303);
nand U22255 (N_22255,N_17430,N_17008);
nor U22256 (N_22256,N_17476,N_17818);
nor U22257 (N_22257,N_16953,N_17840);
xor U22258 (N_22258,N_19841,N_19842);
nand U22259 (N_22259,N_19383,N_16342);
or U22260 (N_22260,N_16854,N_17291);
nor U22261 (N_22261,N_18905,N_19450);
nor U22262 (N_22262,N_19611,N_17922);
and U22263 (N_22263,N_17908,N_17462);
nor U22264 (N_22264,N_18504,N_15996);
nor U22265 (N_22265,N_15739,N_15409);
or U22266 (N_22266,N_18984,N_19767);
xor U22267 (N_22267,N_19578,N_15063);
nand U22268 (N_22268,N_17324,N_17201);
nor U22269 (N_22269,N_19923,N_18014);
or U22270 (N_22270,N_19368,N_19323);
nor U22271 (N_22271,N_16732,N_19469);
nand U22272 (N_22272,N_19950,N_18491);
or U22273 (N_22273,N_17472,N_16109);
nor U22274 (N_22274,N_17032,N_18264);
and U22275 (N_22275,N_15131,N_19734);
xor U22276 (N_22276,N_15530,N_19083);
nor U22277 (N_22277,N_19981,N_16991);
nor U22278 (N_22278,N_18492,N_19382);
xnor U22279 (N_22279,N_15718,N_18245);
or U22280 (N_22280,N_15920,N_19669);
nand U22281 (N_22281,N_16187,N_17744);
nor U22282 (N_22282,N_18103,N_15794);
nand U22283 (N_22283,N_16311,N_18235);
nand U22284 (N_22284,N_17564,N_18589);
xnor U22285 (N_22285,N_19748,N_18017);
and U22286 (N_22286,N_16530,N_17523);
nand U22287 (N_22287,N_15209,N_19363);
and U22288 (N_22288,N_15395,N_16112);
xnor U22289 (N_22289,N_15797,N_18319);
or U22290 (N_22290,N_17644,N_15651);
nand U22291 (N_22291,N_17719,N_16876);
xor U22292 (N_22292,N_15664,N_19076);
and U22293 (N_22293,N_17133,N_16445);
or U22294 (N_22294,N_18963,N_19504);
or U22295 (N_22295,N_18955,N_16318);
and U22296 (N_22296,N_16089,N_18268);
and U22297 (N_22297,N_16262,N_19476);
xnor U22298 (N_22298,N_17740,N_15165);
nor U22299 (N_22299,N_18080,N_15480);
nand U22300 (N_22300,N_19794,N_19801);
or U22301 (N_22301,N_19698,N_17530);
and U22302 (N_22302,N_17603,N_17946);
xor U22303 (N_22303,N_15324,N_19371);
xnor U22304 (N_22304,N_17743,N_17803);
and U22305 (N_22305,N_18481,N_19668);
or U22306 (N_22306,N_19660,N_15157);
or U22307 (N_22307,N_18526,N_15358);
xnor U22308 (N_22308,N_16963,N_16744);
xor U22309 (N_22309,N_19126,N_19562);
or U22310 (N_22310,N_17774,N_15081);
nand U22311 (N_22311,N_19614,N_16447);
nor U22312 (N_22312,N_17559,N_18976);
nor U22313 (N_22313,N_18154,N_16277);
or U22314 (N_22314,N_15580,N_17417);
and U22315 (N_22315,N_17217,N_16633);
xnor U22316 (N_22316,N_15834,N_19803);
and U22317 (N_22317,N_15882,N_19026);
nor U22318 (N_22318,N_18966,N_18332);
nor U22319 (N_22319,N_15541,N_18475);
nor U22320 (N_22320,N_15434,N_16285);
nand U22321 (N_22321,N_15313,N_18749);
or U22322 (N_22322,N_15193,N_17255);
nor U22323 (N_22323,N_18153,N_18276);
and U22324 (N_22324,N_15238,N_18733);
or U22325 (N_22325,N_16950,N_16184);
or U22326 (N_22326,N_19209,N_15612);
nand U22327 (N_22327,N_17077,N_18449);
xnor U22328 (N_22328,N_15264,N_15038);
or U22329 (N_22329,N_15747,N_17769);
nand U22330 (N_22330,N_15891,N_15536);
nor U22331 (N_22331,N_18185,N_17401);
nand U22332 (N_22332,N_18363,N_15126);
nor U22333 (N_22333,N_18952,N_15170);
nand U22334 (N_22334,N_18556,N_19468);
nand U22335 (N_22335,N_16675,N_18761);
and U22336 (N_22336,N_18993,N_19967);
nor U22337 (N_22337,N_19863,N_18459);
xor U22338 (N_22338,N_15341,N_18350);
and U22339 (N_22339,N_16833,N_18440);
nor U22340 (N_22340,N_19171,N_15432);
nor U22341 (N_22341,N_18871,N_16764);
and U22342 (N_22342,N_17512,N_15969);
xor U22343 (N_22343,N_17372,N_19870);
nand U22344 (N_22344,N_16406,N_17552);
xor U22345 (N_22345,N_19319,N_15647);
and U22346 (N_22346,N_15296,N_18176);
nor U22347 (N_22347,N_19649,N_16541);
or U22348 (N_22348,N_15611,N_17728);
nor U22349 (N_22349,N_16058,N_17385);
xnor U22350 (N_22350,N_16442,N_15974);
or U22351 (N_22351,N_16070,N_16235);
nand U22352 (N_22352,N_19167,N_18367);
nand U22353 (N_22353,N_19218,N_16559);
xor U22354 (N_22354,N_17342,N_16867);
and U22355 (N_22355,N_19600,N_15415);
and U22356 (N_22356,N_19568,N_18445);
and U22357 (N_22357,N_19645,N_17851);
or U22358 (N_22358,N_17410,N_19811);
nand U22359 (N_22359,N_15966,N_15771);
nand U22360 (N_22360,N_16625,N_19072);
nor U22361 (N_22361,N_15169,N_18582);
nor U22362 (N_22362,N_15239,N_15761);
or U22363 (N_22363,N_17503,N_15847);
xor U22364 (N_22364,N_17320,N_15945);
xnor U22365 (N_22365,N_17130,N_16548);
nand U22366 (N_22366,N_15744,N_18896);
nor U22367 (N_22367,N_18568,N_15578);
nand U22368 (N_22368,N_16029,N_18850);
and U22369 (N_22369,N_18444,N_15125);
xnor U22370 (N_22370,N_18634,N_18793);
xnor U22371 (N_22371,N_15420,N_16859);
or U22372 (N_22372,N_17006,N_18251);
nor U22373 (N_22373,N_17976,N_17580);
and U22374 (N_22374,N_17269,N_16132);
xnor U22375 (N_22375,N_19336,N_15425);
or U22376 (N_22376,N_19248,N_19440);
or U22377 (N_22377,N_18811,N_18465);
or U22378 (N_22378,N_17616,N_18036);
nor U22379 (N_22379,N_19931,N_17609);
nand U22380 (N_22380,N_15716,N_15556);
nand U22381 (N_22381,N_19615,N_19061);
nor U22382 (N_22382,N_19921,N_16782);
nand U22383 (N_22383,N_19662,N_15366);
xor U22384 (N_22384,N_16629,N_19597);
or U22385 (N_22385,N_19168,N_17304);
nor U22386 (N_22386,N_16197,N_19572);
nor U22387 (N_22387,N_18308,N_18594);
or U22388 (N_22388,N_19995,N_19566);
xnor U22389 (N_22389,N_18353,N_18340);
or U22390 (N_22390,N_18441,N_15511);
and U22391 (N_22391,N_17674,N_15042);
and U22392 (N_22392,N_18676,N_18977);
nor U22393 (N_22393,N_15846,N_19437);
and U22394 (N_22394,N_17208,N_15780);
and U22395 (N_22395,N_18736,N_15509);
nor U22396 (N_22396,N_19548,N_19447);
or U22397 (N_22397,N_16751,N_18373);
nor U22398 (N_22398,N_15018,N_16473);
and U22399 (N_22399,N_18959,N_18852);
nor U22400 (N_22400,N_19260,N_16448);
nor U22401 (N_22401,N_15878,N_15202);
or U22402 (N_22402,N_18936,N_17810);
xor U22403 (N_22403,N_18043,N_17962);
or U22404 (N_22404,N_19326,N_15641);
and U22405 (N_22405,N_16948,N_15435);
xnor U22406 (N_22406,N_18322,N_17300);
nand U22407 (N_22407,N_16662,N_17933);
or U22408 (N_22408,N_16807,N_17071);
nand U22409 (N_22409,N_16102,N_15164);
nor U22410 (N_22410,N_16614,N_19664);
nor U22411 (N_22411,N_17801,N_16158);
xnor U22412 (N_22412,N_16103,N_18520);
nand U22413 (N_22413,N_18138,N_19403);
xnor U22414 (N_22414,N_16378,N_15798);
or U22415 (N_22415,N_17067,N_18971);
xor U22416 (N_22416,N_17678,N_18906);
or U22417 (N_22417,N_15903,N_19125);
xor U22418 (N_22418,N_16061,N_18413);
nor U22419 (N_22419,N_17989,N_17489);
or U22420 (N_22420,N_17569,N_16405);
nor U22421 (N_22421,N_16343,N_19724);
xor U22422 (N_22422,N_15072,N_19275);
nand U22423 (N_22423,N_15220,N_18889);
xor U22424 (N_22424,N_15147,N_16616);
and U22425 (N_22425,N_17682,N_17432);
nand U22426 (N_22426,N_19374,N_19667);
nor U22427 (N_22427,N_19287,N_17582);
and U22428 (N_22428,N_15658,N_17956);
or U22429 (N_22429,N_18979,N_16612);
nor U22430 (N_22430,N_17961,N_16755);
nor U22431 (N_22431,N_17990,N_18281);
and U22432 (N_22432,N_18601,N_17463);
or U22433 (N_22433,N_15673,N_19638);
nor U22434 (N_22434,N_17776,N_18419);
nor U22435 (N_22435,N_17553,N_18239);
nor U22436 (N_22436,N_18086,N_15377);
nand U22437 (N_22437,N_17185,N_17203);
nand U22438 (N_22438,N_18630,N_17794);
or U22439 (N_22439,N_18231,N_16788);
nor U22440 (N_22440,N_15188,N_17521);
and U22441 (N_22441,N_17698,N_18994);
nor U22442 (N_22442,N_16989,N_15575);
nor U22443 (N_22443,N_19204,N_15591);
or U22444 (N_22444,N_18342,N_17019);
nand U22445 (N_22445,N_16137,N_17046);
xnor U22446 (N_22446,N_17547,N_18783);
and U22447 (N_22447,N_19160,N_16974);
nor U22448 (N_22448,N_15491,N_17572);
or U22449 (N_22449,N_18302,N_17182);
and U22450 (N_22450,N_19606,N_19224);
and U22451 (N_22451,N_16203,N_16338);
nand U22452 (N_22452,N_16071,N_15418);
nor U22453 (N_22453,N_19250,N_16939);
nand U22454 (N_22454,N_17191,N_18493);
or U22455 (N_22455,N_16635,N_18599);
nand U22456 (N_22456,N_19744,N_19370);
or U22457 (N_22457,N_16649,N_15043);
xor U22458 (N_22458,N_19622,N_15867);
xor U22459 (N_22459,N_16240,N_16433);
xnor U22460 (N_22460,N_19932,N_17377);
or U22461 (N_22461,N_15581,N_19199);
nand U22462 (N_22462,N_15831,N_17362);
or U22463 (N_22463,N_19715,N_15919);
nor U22464 (N_22464,N_17504,N_18718);
or U22465 (N_22465,N_19920,N_17535);
xor U22466 (N_22466,N_17927,N_16890);
nand U22467 (N_22467,N_19273,N_17065);
and U22468 (N_22468,N_16276,N_15762);
xor U22469 (N_22469,N_17987,N_16359);
or U22470 (N_22470,N_15512,N_17713);
nor U22471 (N_22471,N_16208,N_15458);
or U22472 (N_22472,N_18421,N_15665);
nand U22473 (N_22473,N_17730,N_17279);
and U22474 (N_22474,N_18690,N_19073);
nand U22475 (N_22475,N_16141,N_15319);
nor U22476 (N_22476,N_16797,N_16845);
xor U22477 (N_22477,N_19738,N_17647);
nor U22478 (N_22478,N_16524,N_18217);
xnor U22479 (N_22479,N_19092,N_15225);
nor U22480 (N_22480,N_16427,N_18131);
and U22481 (N_22481,N_18597,N_18897);
nand U22482 (N_22482,N_16804,N_17623);
nand U22483 (N_22483,N_17696,N_15675);
xnor U22484 (N_22484,N_15897,N_15517);
or U22485 (N_22485,N_15200,N_19402);
nand U22486 (N_22486,N_19129,N_15679);
and U22487 (N_22487,N_17785,N_18574);
xor U22488 (N_22488,N_16582,N_17151);
and U22489 (N_22489,N_15924,N_18201);
or U22490 (N_22490,N_15368,N_18463);
nand U22491 (N_22491,N_17099,N_18999);
and U22492 (N_22492,N_15808,N_18547);
nor U22493 (N_22493,N_15241,N_19470);
nor U22494 (N_22494,N_16252,N_19831);
nor U22495 (N_22495,N_19201,N_16947);
or U22496 (N_22496,N_19880,N_17620);
xor U22497 (N_22497,N_19216,N_19433);
or U22498 (N_22498,N_19839,N_16937);
or U22499 (N_22499,N_16361,N_16743);
or U22500 (N_22500,N_16330,N_18597);
and U22501 (N_22501,N_19577,N_16011);
or U22502 (N_22502,N_15447,N_15190);
xnor U22503 (N_22503,N_19168,N_19716);
nand U22504 (N_22504,N_15774,N_16942);
nor U22505 (N_22505,N_18956,N_19180);
xnor U22506 (N_22506,N_19828,N_17443);
xor U22507 (N_22507,N_19973,N_18441);
nor U22508 (N_22508,N_17238,N_15541);
nand U22509 (N_22509,N_17519,N_17693);
nor U22510 (N_22510,N_19719,N_16207);
or U22511 (N_22511,N_15927,N_18693);
nand U22512 (N_22512,N_15109,N_16391);
xor U22513 (N_22513,N_16905,N_15715);
nand U22514 (N_22514,N_16502,N_15057);
nand U22515 (N_22515,N_15658,N_18535);
and U22516 (N_22516,N_15411,N_17211);
and U22517 (N_22517,N_15236,N_16921);
xnor U22518 (N_22518,N_16673,N_16529);
xnor U22519 (N_22519,N_15861,N_18940);
nand U22520 (N_22520,N_18354,N_18793);
and U22521 (N_22521,N_19741,N_16661);
nand U22522 (N_22522,N_18016,N_19880);
and U22523 (N_22523,N_18141,N_17863);
nand U22524 (N_22524,N_19500,N_15322);
nor U22525 (N_22525,N_16639,N_19070);
or U22526 (N_22526,N_18495,N_17160);
or U22527 (N_22527,N_16093,N_15464);
and U22528 (N_22528,N_17496,N_18197);
and U22529 (N_22529,N_15816,N_19444);
xnor U22530 (N_22530,N_16645,N_18203);
and U22531 (N_22531,N_19624,N_17508);
and U22532 (N_22532,N_18203,N_15661);
or U22533 (N_22533,N_16379,N_19299);
or U22534 (N_22534,N_19655,N_18763);
or U22535 (N_22535,N_15565,N_19938);
or U22536 (N_22536,N_16242,N_17642);
or U22537 (N_22537,N_18944,N_18973);
or U22538 (N_22538,N_19084,N_18081);
nand U22539 (N_22539,N_18335,N_15735);
nand U22540 (N_22540,N_18641,N_18483);
nand U22541 (N_22541,N_17915,N_19986);
or U22542 (N_22542,N_16267,N_17028);
nor U22543 (N_22543,N_17340,N_18067);
nand U22544 (N_22544,N_18966,N_17377);
xor U22545 (N_22545,N_18834,N_15770);
or U22546 (N_22546,N_19379,N_17172);
xor U22547 (N_22547,N_17925,N_17445);
nand U22548 (N_22548,N_18002,N_18538);
nand U22549 (N_22549,N_16910,N_19743);
xor U22550 (N_22550,N_16935,N_18964);
and U22551 (N_22551,N_18236,N_15027);
or U22552 (N_22552,N_19997,N_18981);
or U22553 (N_22553,N_18703,N_16798);
and U22554 (N_22554,N_15558,N_19511);
and U22555 (N_22555,N_15045,N_19086);
xor U22556 (N_22556,N_18931,N_15395);
xnor U22557 (N_22557,N_16443,N_16171);
or U22558 (N_22558,N_16503,N_19704);
or U22559 (N_22559,N_19422,N_19238);
nor U22560 (N_22560,N_15720,N_15813);
xor U22561 (N_22561,N_19749,N_17505);
nand U22562 (N_22562,N_16876,N_15094);
xnor U22563 (N_22563,N_15245,N_18026);
xor U22564 (N_22564,N_17918,N_15812);
or U22565 (N_22565,N_19539,N_16188);
nand U22566 (N_22566,N_15141,N_19963);
xnor U22567 (N_22567,N_19770,N_19125);
or U22568 (N_22568,N_15684,N_17898);
and U22569 (N_22569,N_17233,N_16723);
and U22570 (N_22570,N_16788,N_16413);
nor U22571 (N_22571,N_18091,N_18771);
and U22572 (N_22572,N_17500,N_16616);
nor U22573 (N_22573,N_17322,N_18787);
nor U22574 (N_22574,N_18126,N_19136);
nor U22575 (N_22575,N_15777,N_18983);
xor U22576 (N_22576,N_18992,N_18893);
nor U22577 (N_22577,N_19653,N_17965);
nand U22578 (N_22578,N_16716,N_15569);
nor U22579 (N_22579,N_16246,N_18431);
nand U22580 (N_22580,N_15989,N_16696);
xnor U22581 (N_22581,N_15345,N_16490);
nor U22582 (N_22582,N_19566,N_18276);
nor U22583 (N_22583,N_18274,N_15197);
nor U22584 (N_22584,N_18388,N_15092);
nand U22585 (N_22585,N_17394,N_18081);
nand U22586 (N_22586,N_17086,N_16710);
nor U22587 (N_22587,N_15393,N_18870);
nand U22588 (N_22588,N_15541,N_15320);
nand U22589 (N_22589,N_15043,N_19616);
nor U22590 (N_22590,N_16381,N_17141);
and U22591 (N_22591,N_15499,N_16247);
nor U22592 (N_22592,N_15042,N_19003);
nand U22593 (N_22593,N_19991,N_19489);
nor U22594 (N_22594,N_15079,N_16547);
nor U22595 (N_22595,N_16565,N_17937);
and U22596 (N_22596,N_19460,N_17372);
nor U22597 (N_22597,N_19198,N_18781);
and U22598 (N_22598,N_16809,N_19819);
nand U22599 (N_22599,N_18623,N_15903);
nor U22600 (N_22600,N_19881,N_18593);
or U22601 (N_22601,N_17501,N_18103);
or U22602 (N_22602,N_19445,N_16581);
nand U22603 (N_22603,N_15112,N_15400);
and U22604 (N_22604,N_16095,N_18753);
nor U22605 (N_22605,N_15211,N_17389);
nor U22606 (N_22606,N_19751,N_19975);
nor U22607 (N_22607,N_17038,N_18260);
nand U22608 (N_22608,N_16238,N_17828);
nor U22609 (N_22609,N_15193,N_18374);
nand U22610 (N_22610,N_17348,N_15701);
xnor U22611 (N_22611,N_16325,N_16744);
or U22612 (N_22612,N_16596,N_16431);
nor U22613 (N_22613,N_18423,N_17671);
xnor U22614 (N_22614,N_16892,N_17835);
and U22615 (N_22615,N_18571,N_16077);
nor U22616 (N_22616,N_17835,N_17850);
nand U22617 (N_22617,N_18516,N_16152);
nand U22618 (N_22618,N_18726,N_19576);
nand U22619 (N_22619,N_18873,N_16889);
xor U22620 (N_22620,N_18524,N_15885);
nand U22621 (N_22621,N_19615,N_15334);
and U22622 (N_22622,N_18951,N_15091);
nand U22623 (N_22623,N_16608,N_15675);
xor U22624 (N_22624,N_15811,N_19930);
nor U22625 (N_22625,N_16763,N_17879);
and U22626 (N_22626,N_16559,N_18752);
and U22627 (N_22627,N_18633,N_16155);
or U22628 (N_22628,N_15082,N_18173);
nor U22629 (N_22629,N_17745,N_16028);
xor U22630 (N_22630,N_18210,N_16419);
and U22631 (N_22631,N_18440,N_15217);
xnor U22632 (N_22632,N_16854,N_19172);
nor U22633 (N_22633,N_17816,N_16726);
and U22634 (N_22634,N_19908,N_18044);
nor U22635 (N_22635,N_18185,N_18071);
nor U22636 (N_22636,N_15083,N_15366);
or U22637 (N_22637,N_18572,N_15657);
and U22638 (N_22638,N_19126,N_17774);
or U22639 (N_22639,N_17702,N_18262);
and U22640 (N_22640,N_18584,N_18523);
or U22641 (N_22641,N_19226,N_16782);
or U22642 (N_22642,N_18225,N_18100);
nand U22643 (N_22643,N_16082,N_16323);
or U22644 (N_22644,N_19046,N_19250);
nand U22645 (N_22645,N_16205,N_18716);
nand U22646 (N_22646,N_16891,N_18850);
nor U22647 (N_22647,N_18365,N_17093);
nor U22648 (N_22648,N_15369,N_18125);
or U22649 (N_22649,N_16518,N_18496);
xor U22650 (N_22650,N_17187,N_15089);
nand U22651 (N_22651,N_16049,N_17771);
and U22652 (N_22652,N_17586,N_18179);
nand U22653 (N_22653,N_18377,N_18292);
xnor U22654 (N_22654,N_15272,N_17409);
xor U22655 (N_22655,N_19390,N_16331);
nand U22656 (N_22656,N_19209,N_16932);
or U22657 (N_22657,N_17680,N_17467);
or U22658 (N_22658,N_17843,N_17680);
nand U22659 (N_22659,N_17174,N_16843);
nand U22660 (N_22660,N_16724,N_18058);
nand U22661 (N_22661,N_15717,N_19265);
and U22662 (N_22662,N_18505,N_16594);
nor U22663 (N_22663,N_19444,N_15302);
and U22664 (N_22664,N_17399,N_19167);
xnor U22665 (N_22665,N_18974,N_17570);
or U22666 (N_22666,N_16156,N_15000);
xor U22667 (N_22667,N_19061,N_19845);
and U22668 (N_22668,N_19860,N_15675);
or U22669 (N_22669,N_19988,N_19176);
xnor U22670 (N_22670,N_18330,N_19421);
nand U22671 (N_22671,N_15144,N_18408);
or U22672 (N_22672,N_18460,N_15325);
nor U22673 (N_22673,N_17891,N_16839);
xnor U22674 (N_22674,N_19008,N_16784);
and U22675 (N_22675,N_17072,N_16751);
and U22676 (N_22676,N_17329,N_16319);
xnor U22677 (N_22677,N_15657,N_17236);
and U22678 (N_22678,N_15629,N_15856);
and U22679 (N_22679,N_19028,N_15183);
xor U22680 (N_22680,N_17204,N_17130);
xnor U22681 (N_22681,N_17866,N_15154);
nand U22682 (N_22682,N_19182,N_19348);
nor U22683 (N_22683,N_16901,N_17063);
and U22684 (N_22684,N_19769,N_19541);
nor U22685 (N_22685,N_16495,N_18805);
or U22686 (N_22686,N_19894,N_18788);
nor U22687 (N_22687,N_19784,N_19336);
or U22688 (N_22688,N_18165,N_16119);
or U22689 (N_22689,N_16730,N_15500);
or U22690 (N_22690,N_15966,N_15640);
nor U22691 (N_22691,N_16397,N_18559);
nand U22692 (N_22692,N_18573,N_19700);
or U22693 (N_22693,N_19352,N_16030);
and U22694 (N_22694,N_16997,N_18234);
nand U22695 (N_22695,N_17421,N_18444);
and U22696 (N_22696,N_15511,N_18866);
nor U22697 (N_22697,N_17333,N_18645);
xor U22698 (N_22698,N_15932,N_16316);
or U22699 (N_22699,N_15404,N_15319);
nand U22700 (N_22700,N_18455,N_19336);
or U22701 (N_22701,N_17549,N_16318);
xnor U22702 (N_22702,N_15123,N_16043);
or U22703 (N_22703,N_18120,N_17779);
xnor U22704 (N_22704,N_18537,N_18261);
nand U22705 (N_22705,N_17225,N_19972);
nand U22706 (N_22706,N_17426,N_19328);
xor U22707 (N_22707,N_15939,N_15483);
or U22708 (N_22708,N_15544,N_18387);
or U22709 (N_22709,N_17559,N_15216);
nor U22710 (N_22710,N_15972,N_19926);
nand U22711 (N_22711,N_18806,N_18023);
and U22712 (N_22712,N_15037,N_19995);
and U22713 (N_22713,N_17489,N_18925);
xnor U22714 (N_22714,N_19797,N_18875);
nor U22715 (N_22715,N_18496,N_16348);
or U22716 (N_22716,N_15620,N_18471);
or U22717 (N_22717,N_17653,N_18425);
and U22718 (N_22718,N_19225,N_19322);
and U22719 (N_22719,N_18063,N_19834);
nor U22720 (N_22720,N_19401,N_17663);
nor U22721 (N_22721,N_15101,N_15416);
nand U22722 (N_22722,N_19498,N_18710);
xor U22723 (N_22723,N_16269,N_15558);
nand U22724 (N_22724,N_17392,N_16676);
nand U22725 (N_22725,N_18791,N_18494);
nor U22726 (N_22726,N_17593,N_15000);
or U22727 (N_22727,N_15477,N_17057);
nor U22728 (N_22728,N_17972,N_18782);
or U22729 (N_22729,N_19867,N_18180);
and U22730 (N_22730,N_16703,N_16704);
and U22731 (N_22731,N_15148,N_16888);
and U22732 (N_22732,N_17192,N_18232);
nor U22733 (N_22733,N_18239,N_16470);
and U22734 (N_22734,N_17451,N_16057);
and U22735 (N_22735,N_16638,N_17475);
nor U22736 (N_22736,N_18200,N_19043);
nand U22737 (N_22737,N_18720,N_16453);
nor U22738 (N_22738,N_18014,N_15600);
and U22739 (N_22739,N_16494,N_15876);
nand U22740 (N_22740,N_17395,N_17462);
nor U22741 (N_22741,N_18527,N_17537);
or U22742 (N_22742,N_19479,N_19289);
nand U22743 (N_22743,N_15365,N_15462);
nor U22744 (N_22744,N_16818,N_18109);
nand U22745 (N_22745,N_19775,N_19233);
nor U22746 (N_22746,N_18271,N_16375);
and U22747 (N_22747,N_15696,N_16741);
xor U22748 (N_22748,N_16988,N_16462);
xor U22749 (N_22749,N_19776,N_19912);
nand U22750 (N_22750,N_17060,N_19396);
nand U22751 (N_22751,N_18034,N_19527);
or U22752 (N_22752,N_15659,N_17688);
xor U22753 (N_22753,N_17417,N_15925);
nand U22754 (N_22754,N_18671,N_17949);
nor U22755 (N_22755,N_18793,N_15117);
nand U22756 (N_22756,N_15730,N_15771);
or U22757 (N_22757,N_19389,N_18299);
or U22758 (N_22758,N_16394,N_16695);
and U22759 (N_22759,N_18313,N_16382);
xor U22760 (N_22760,N_19963,N_16117);
nor U22761 (N_22761,N_16065,N_17917);
nand U22762 (N_22762,N_17990,N_16235);
or U22763 (N_22763,N_18642,N_15074);
xnor U22764 (N_22764,N_16537,N_18230);
nor U22765 (N_22765,N_16940,N_17924);
xor U22766 (N_22766,N_18630,N_16823);
or U22767 (N_22767,N_15831,N_17835);
xor U22768 (N_22768,N_19173,N_18318);
or U22769 (N_22769,N_15980,N_16808);
xnor U22770 (N_22770,N_17983,N_17332);
xnor U22771 (N_22771,N_15778,N_17316);
nand U22772 (N_22772,N_16990,N_17724);
xnor U22773 (N_22773,N_18334,N_16308);
xnor U22774 (N_22774,N_16822,N_17407);
nand U22775 (N_22775,N_18323,N_15658);
and U22776 (N_22776,N_19896,N_18789);
or U22777 (N_22777,N_15699,N_17631);
nand U22778 (N_22778,N_15217,N_17287);
or U22779 (N_22779,N_17056,N_19751);
nor U22780 (N_22780,N_16219,N_17782);
and U22781 (N_22781,N_18621,N_17085);
and U22782 (N_22782,N_18967,N_16224);
nand U22783 (N_22783,N_18736,N_15937);
or U22784 (N_22784,N_18791,N_18015);
nand U22785 (N_22785,N_16694,N_18714);
xor U22786 (N_22786,N_15497,N_17698);
or U22787 (N_22787,N_16796,N_16016);
nand U22788 (N_22788,N_19132,N_19868);
and U22789 (N_22789,N_18335,N_16805);
and U22790 (N_22790,N_19969,N_18188);
nand U22791 (N_22791,N_15670,N_17746);
and U22792 (N_22792,N_19374,N_17551);
or U22793 (N_22793,N_18043,N_19288);
and U22794 (N_22794,N_18164,N_18709);
nor U22795 (N_22795,N_18785,N_17152);
nand U22796 (N_22796,N_19993,N_15420);
xnor U22797 (N_22797,N_16253,N_18179);
xnor U22798 (N_22798,N_18249,N_15285);
or U22799 (N_22799,N_15560,N_17117);
xor U22800 (N_22800,N_16481,N_18993);
xor U22801 (N_22801,N_18164,N_16281);
nand U22802 (N_22802,N_16193,N_19520);
nand U22803 (N_22803,N_16799,N_19732);
and U22804 (N_22804,N_15261,N_19121);
nor U22805 (N_22805,N_19754,N_18786);
and U22806 (N_22806,N_18206,N_19086);
or U22807 (N_22807,N_19417,N_16603);
nor U22808 (N_22808,N_19177,N_16827);
nor U22809 (N_22809,N_19398,N_17862);
or U22810 (N_22810,N_19655,N_16019);
or U22811 (N_22811,N_19962,N_19972);
or U22812 (N_22812,N_19179,N_18126);
nor U22813 (N_22813,N_15676,N_16739);
or U22814 (N_22814,N_15193,N_16638);
nand U22815 (N_22815,N_19228,N_17313);
nor U22816 (N_22816,N_19031,N_15656);
nor U22817 (N_22817,N_15821,N_15878);
and U22818 (N_22818,N_17244,N_17600);
nor U22819 (N_22819,N_17267,N_19449);
or U22820 (N_22820,N_19916,N_17939);
nand U22821 (N_22821,N_16355,N_16872);
or U22822 (N_22822,N_18752,N_17046);
xnor U22823 (N_22823,N_17931,N_15873);
xnor U22824 (N_22824,N_18891,N_18972);
and U22825 (N_22825,N_19893,N_18634);
nand U22826 (N_22826,N_18436,N_16395);
nor U22827 (N_22827,N_19356,N_17345);
and U22828 (N_22828,N_16145,N_18417);
xnor U22829 (N_22829,N_16695,N_17597);
xor U22830 (N_22830,N_15247,N_19853);
nand U22831 (N_22831,N_15770,N_16327);
and U22832 (N_22832,N_16030,N_15011);
and U22833 (N_22833,N_18605,N_18362);
or U22834 (N_22834,N_18319,N_16514);
nor U22835 (N_22835,N_15394,N_16991);
or U22836 (N_22836,N_17760,N_15899);
and U22837 (N_22837,N_19492,N_15156);
nor U22838 (N_22838,N_19726,N_15965);
xor U22839 (N_22839,N_18818,N_19358);
and U22840 (N_22840,N_16276,N_18955);
nand U22841 (N_22841,N_15266,N_15774);
and U22842 (N_22842,N_19240,N_16977);
xor U22843 (N_22843,N_17530,N_18174);
or U22844 (N_22844,N_19408,N_17851);
or U22845 (N_22845,N_15637,N_18132);
nor U22846 (N_22846,N_18907,N_15847);
nor U22847 (N_22847,N_18474,N_19525);
nand U22848 (N_22848,N_15531,N_18331);
nand U22849 (N_22849,N_19654,N_15236);
xnor U22850 (N_22850,N_19988,N_15938);
nand U22851 (N_22851,N_16061,N_16373);
nand U22852 (N_22852,N_19024,N_17608);
or U22853 (N_22853,N_19548,N_18410);
xnor U22854 (N_22854,N_17251,N_15225);
nand U22855 (N_22855,N_17615,N_19587);
nor U22856 (N_22856,N_15734,N_15041);
nor U22857 (N_22857,N_18985,N_16407);
and U22858 (N_22858,N_17764,N_15384);
nor U22859 (N_22859,N_16136,N_17105);
and U22860 (N_22860,N_15799,N_19076);
and U22861 (N_22861,N_15819,N_15050);
and U22862 (N_22862,N_19738,N_15422);
nand U22863 (N_22863,N_19632,N_17242);
nand U22864 (N_22864,N_16138,N_18327);
nand U22865 (N_22865,N_17188,N_19708);
nor U22866 (N_22866,N_19564,N_15605);
nand U22867 (N_22867,N_17301,N_17283);
nor U22868 (N_22868,N_19603,N_15064);
and U22869 (N_22869,N_16312,N_15014);
xor U22870 (N_22870,N_18958,N_15701);
nor U22871 (N_22871,N_17339,N_19260);
nor U22872 (N_22872,N_19645,N_18088);
or U22873 (N_22873,N_19904,N_15542);
nor U22874 (N_22874,N_17512,N_15003);
and U22875 (N_22875,N_16530,N_16687);
xnor U22876 (N_22876,N_18768,N_15289);
nand U22877 (N_22877,N_19020,N_17073);
xor U22878 (N_22878,N_15496,N_19994);
nor U22879 (N_22879,N_15355,N_16425);
or U22880 (N_22880,N_15088,N_19286);
and U22881 (N_22881,N_15614,N_17650);
nor U22882 (N_22882,N_17240,N_15212);
nand U22883 (N_22883,N_17040,N_16564);
nand U22884 (N_22884,N_16367,N_15510);
nor U22885 (N_22885,N_18580,N_17895);
or U22886 (N_22886,N_16035,N_19309);
or U22887 (N_22887,N_18683,N_16717);
nand U22888 (N_22888,N_15506,N_15677);
and U22889 (N_22889,N_16729,N_16582);
nor U22890 (N_22890,N_16949,N_19302);
nand U22891 (N_22891,N_16927,N_16097);
xnor U22892 (N_22892,N_16679,N_18723);
and U22893 (N_22893,N_16525,N_15900);
or U22894 (N_22894,N_17457,N_16577);
or U22895 (N_22895,N_15582,N_17516);
and U22896 (N_22896,N_17935,N_15805);
and U22897 (N_22897,N_19490,N_17978);
nor U22898 (N_22898,N_15152,N_19512);
or U22899 (N_22899,N_15176,N_19943);
xnor U22900 (N_22900,N_17793,N_16389);
nor U22901 (N_22901,N_19604,N_17368);
nor U22902 (N_22902,N_17450,N_17730);
and U22903 (N_22903,N_19647,N_19513);
nand U22904 (N_22904,N_15874,N_18988);
nand U22905 (N_22905,N_17997,N_18746);
nor U22906 (N_22906,N_15548,N_16813);
and U22907 (N_22907,N_17134,N_18985);
xor U22908 (N_22908,N_19862,N_19600);
and U22909 (N_22909,N_18707,N_18426);
nand U22910 (N_22910,N_18835,N_16503);
xor U22911 (N_22911,N_17719,N_18861);
or U22912 (N_22912,N_15446,N_17329);
nor U22913 (N_22913,N_19139,N_19396);
xor U22914 (N_22914,N_16987,N_16696);
nor U22915 (N_22915,N_15524,N_16295);
xnor U22916 (N_22916,N_17646,N_19396);
or U22917 (N_22917,N_18767,N_18879);
nand U22918 (N_22918,N_16069,N_18485);
xor U22919 (N_22919,N_17822,N_15370);
and U22920 (N_22920,N_16329,N_19520);
or U22921 (N_22921,N_18537,N_15015);
and U22922 (N_22922,N_18879,N_19217);
and U22923 (N_22923,N_16993,N_18917);
nand U22924 (N_22924,N_18033,N_19048);
nand U22925 (N_22925,N_19625,N_16515);
nand U22926 (N_22926,N_18629,N_15413);
nor U22927 (N_22927,N_19418,N_17984);
nand U22928 (N_22928,N_17293,N_16520);
nor U22929 (N_22929,N_15254,N_15949);
nor U22930 (N_22930,N_17203,N_17414);
xnor U22931 (N_22931,N_15488,N_15644);
nor U22932 (N_22932,N_19438,N_18467);
and U22933 (N_22933,N_19217,N_15280);
nand U22934 (N_22934,N_17173,N_16791);
nand U22935 (N_22935,N_18154,N_16024);
xor U22936 (N_22936,N_15571,N_19198);
and U22937 (N_22937,N_18857,N_15499);
or U22938 (N_22938,N_18347,N_18835);
nor U22939 (N_22939,N_18975,N_18170);
nand U22940 (N_22940,N_19509,N_18339);
and U22941 (N_22941,N_15172,N_18537);
or U22942 (N_22942,N_16619,N_17556);
and U22943 (N_22943,N_19784,N_18021);
and U22944 (N_22944,N_18564,N_17509);
xor U22945 (N_22945,N_15121,N_19323);
xnor U22946 (N_22946,N_17378,N_16395);
and U22947 (N_22947,N_15714,N_15167);
nor U22948 (N_22948,N_19219,N_17281);
and U22949 (N_22949,N_19519,N_15727);
and U22950 (N_22950,N_18049,N_17818);
nor U22951 (N_22951,N_17574,N_18468);
nand U22952 (N_22952,N_16962,N_18351);
or U22953 (N_22953,N_16569,N_18218);
nand U22954 (N_22954,N_15281,N_17463);
or U22955 (N_22955,N_15144,N_18388);
nor U22956 (N_22956,N_16468,N_18487);
nand U22957 (N_22957,N_19415,N_19490);
xnor U22958 (N_22958,N_16598,N_16148);
and U22959 (N_22959,N_15294,N_19103);
and U22960 (N_22960,N_15400,N_19657);
and U22961 (N_22961,N_18208,N_18120);
nor U22962 (N_22962,N_18569,N_17227);
or U22963 (N_22963,N_18724,N_18888);
or U22964 (N_22964,N_17207,N_18625);
nor U22965 (N_22965,N_15477,N_15656);
and U22966 (N_22966,N_16995,N_19077);
nor U22967 (N_22967,N_16082,N_19727);
nor U22968 (N_22968,N_15741,N_17155);
xor U22969 (N_22969,N_16021,N_18195);
or U22970 (N_22970,N_18176,N_17222);
xnor U22971 (N_22971,N_16344,N_17420);
or U22972 (N_22972,N_17916,N_18075);
nand U22973 (N_22973,N_16507,N_16483);
or U22974 (N_22974,N_18891,N_17287);
xnor U22975 (N_22975,N_18912,N_16092);
and U22976 (N_22976,N_17830,N_16248);
or U22977 (N_22977,N_18543,N_19867);
and U22978 (N_22978,N_16930,N_19167);
nor U22979 (N_22979,N_17987,N_15753);
or U22980 (N_22980,N_15488,N_19303);
and U22981 (N_22981,N_15406,N_18006);
nor U22982 (N_22982,N_18142,N_17833);
nand U22983 (N_22983,N_15043,N_18747);
and U22984 (N_22984,N_16069,N_17310);
and U22985 (N_22985,N_15019,N_15713);
or U22986 (N_22986,N_16252,N_18914);
nand U22987 (N_22987,N_17255,N_19704);
nor U22988 (N_22988,N_17995,N_15918);
nand U22989 (N_22989,N_19959,N_15012);
nor U22990 (N_22990,N_15605,N_18138);
nand U22991 (N_22991,N_18555,N_17190);
and U22992 (N_22992,N_19941,N_18677);
xor U22993 (N_22993,N_17323,N_16256);
nor U22994 (N_22994,N_15172,N_15331);
nand U22995 (N_22995,N_16783,N_17087);
nor U22996 (N_22996,N_19628,N_17040);
xor U22997 (N_22997,N_15954,N_15276);
nand U22998 (N_22998,N_16300,N_18804);
nand U22999 (N_22999,N_19011,N_17233);
nand U23000 (N_23000,N_15263,N_15362);
and U23001 (N_23001,N_16056,N_16791);
nor U23002 (N_23002,N_18161,N_18284);
nand U23003 (N_23003,N_18320,N_15269);
nand U23004 (N_23004,N_19077,N_19544);
or U23005 (N_23005,N_19031,N_17411);
and U23006 (N_23006,N_18085,N_17216);
and U23007 (N_23007,N_18559,N_15055);
nor U23008 (N_23008,N_15361,N_17839);
nand U23009 (N_23009,N_17595,N_16891);
and U23010 (N_23010,N_16350,N_18646);
xor U23011 (N_23011,N_19828,N_15167);
nor U23012 (N_23012,N_16308,N_19581);
xor U23013 (N_23013,N_15342,N_19910);
nor U23014 (N_23014,N_17604,N_19278);
xnor U23015 (N_23015,N_19120,N_18425);
and U23016 (N_23016,N_15834,N_18920);
nor U23017 (N_23017,N_15282,N_18240);
nand U23018 (N_23018,N_17145,N_15608);
nand U23019 (N_23019,N_19313,N_19600);
nor U23020 (N_23020,N_17776,N_16543);
and U23021 (N_23021,N_16583,N_17197);
and U23022 (N_23022,N_16653,N_15900);
nand U23023 (N_23023,N_17082,N_15703);
and U23024 (N_23024,N_16625,N_19460);
nand U23025 (N_23025,N_15808,N_16752);
nand U23026 (N_23026,N_18975,N_16087);
nand U23027 (N_23027,N_19213,N_18753);
nor U23028 (N_23028,N_16075,N_15558);
xor U23029 (N_23029,N_17743,N_18129);
xor U23030 (N_23030,N_19440,N_17949);
and U23031 (N_23031,N_18754,N_17367);
nor U23032 (N_23032,N_16177,N_15320);
nand U23033 (N_23033,N_17742,N_15858);
xnor U23034 (N_23034,N_18785,N_18523);
nor U23035 (N_23035,N_19512,N_15969);
and U23036 (N_23036,N_18136,N_17252);
nand U23037 (N_23037,N_19736,N_17289);
nand U23038 (N_23038,N_15298,N_15287);
and U23039 (N_23039,N_15112,N_18060);
or U23040 (N_23040,N_17678,N_19717);
and U23041 (N_23041,N_16864,N_19611);
nand U23042 (N_23042,N_15728,N_17993);
xnor U23043 (N_23043,N_18477,N_16661);
and U23044 (N_23044,N_16592,N_19032);
nor U23045 (N_23045,N_19737,N_18452);
nor U23046 (N_23046,N_15418,N_15649);
nand U23047 (N_23047,N_19447,N_16774);
nor U23048 (N_23048,N_18894,N_18326);
and U23049 (N_23049,N_18160,N_18208);
nor U23050 (N_23050,N_18220,N_19063);
or U23051 (N_23051,N_17934,N_16321);
nand U23052 (N_23052,N_18397,N_18034);
nand U23053 (N_23053,N_18621,N_16991);
or U23054 (N_23054,N_19174,N_19279);
and U23055 (N_23055,N_18360,N_19406);
xor U23056 (N_23056,N_15430,N_19350);
and U23057 (N_23057,N_19208,N_17391);
xor U23058 (N_23058,N_17540,N_19172);
and U23059 (N_23059,N_17716,N_18641);
or U23060 (N_23060,N_16763,N_17176);
xnor U23061 (N_23061,N_18365,N_17605);
or U23062 (N_23062,N_17952,N_16585);
and U23063 (N_23063,N_17790,N_16897);
nand U23064 (N_23064,N_17482,N_16160);
or U23065 (N_23065,N_17675,N_18993);
xnor U23066 (N_23066,N_16001,N_16251);
or U23067 (N_23067,N_16023,N_18836);
xor U23068 (N_23068,N_18973,N_18194);
xor U23069 (N_23069,N_18718,N_19127);
xor U23070 (N_23070,N_18024,N_18254);
nand U23071 (N_23071,N_16267,N_18620);
xor U23072 (N_23072,N_19870,N_15719);
nand U23073 (N_23073,N_16863,N_17883);
xor U23074 (N_23074,N_19944,N_19132);
nand U23075 (N_23075,N_16419,N_16666);
nand U23076 (N_23076,N_15264,N_15700);
nor U23077 (N_23077,N_18131,N_17982);
and U23078 (N_23078,N_15834,N_17846);
or U23079 (N_23079,N_16189,N_18130);
nand U23080 (N_23080,N_16856,N_17644);
nand U23081 (N_23081,N_15631,N_19914);
nand U23082 (N_23082,N_18482,N_17594);
and U23083 (N_23083,N_19269,N_16839);
nand U23084 (N_23084,N_15158,N_17170);
xnor U23085 (N_23085,N_15633,N_16498);
xor U23086 (N_23086,N_17604,N_17306);
nor U23087 (N_23087,N_16749,N_16737);
or U23088 (N_23088,N_16254,N_18760);
nand U23089 (N_23089,N_19594,N_18741);
nand U23090 (N_23090,N_17711,N_18170);
or U23091 (N_23091,N_17698,N_18395);
or U23092 (N_23092,N_16793,N_16551);
and U23093 (N_23093,N_18555,N_17804);
nor U23094 (N_23094,N_15705,N_16106);
xor U23095 (N_23095,N_17128,N_17607);
nor U23096 (N_23096,N_19481,N_18781);
xnor U23097 (N_23097,N_19228,N_18565);
or U23098 (N_23098,N_15666,N_17642);
and U23099 (N_23099,N_17124,N_16962);
xor U23100 (N_23100,N_15716,N_16592);
nand U23101 (N_23101,N_17092,N_19379);
xor U23102 (N_23102,N_19330,N_16110);
and U23103 (N_23103,N_18253,N_15763);
or U23104 (N_23104,N_16599,N_19359);
and U23105 (N_23105,N_16739,N_15548);
xor U23106 (N_23106,N_15640,N_17618);
xnor U23107 (N_23107,N_19083,N_18037);
nand U23108 (N_23108,N_18433,N_15117);
xnor U23109 (N_23109,N_19218,N_17988);
nand U23110 (N_23110,N_15949,N_17800);
xor U23111 (N_23111,N_17898,N_19661);
or U23112 (N_23112,N_19943,N_19761);
nand U23113 (N_23113,N_17521,N_19583);
nand U23114 (N_23114,N_15308,N_15067);
nor U23115 (N_23115,N_18391,N_19297);
xor U23116 (N_23116,N_19689,N_18978);
nand U23117 (N_23117,N_19580,N_17201);
and U23118 (N_23118,N_17359,N_15915);
and U23119 (N_23119,N_17893,N_15139);
nor U23120 (N_23120,N_15663,N_17086);
nor U23121 (N_23121,N_18596,N_15709);
nand U23122 (N_23122,N_16948,N_19826);
nor U23123 (N_23123,N_15511,N_16699);
nand U23124 (N_23124,N_15052,N_19301);
and U23125 (N_23125,N_15516,N_16258);
xor U23126 (N_23126,N_15281,N_18305);
nor U23127 (N_23127,N_19601,N_18803);
nand U23128 (N_23128,N_17684,N_16849);
nor U23129 (N_23129,N_15012,N_17520);
and U23130 (N_23130,N_18021,N_19335);
xor U23131 (N_23131,N_18165,N_18098);
xnor U23132 (N_23132,N_15579,N_19119);
nor U23133 (N_23133,N_17283,N_19863);
and U23134 (N_23134,N_17615,N_15057);
nor U23135 (N_23135,N_17928,N_17300);
nand U23136 (N_23136,N_18734,N_19848);
nand U23137 (N_23137,N_16745,N_16761);
nor U23138 (N_23138,N_16631,N_16002);
nor U23139 (N_23139,N_15317,N_17434);
nand U23140 (N_23140,N_19964,N_17776);
and U23141 (N_23141,N_17519,N_16107);
xnor U23142 (N_23142,N_15252,N_17198);
or U23143 (N_23143,N_16561,N_19802);
nor U23144 (N_23144,N_19065,N_19272);
and U23145 (N_23145,N_17963,N_18355);
nand U23146 (N_23146,N_19106,N_17436);
and U23147 (N_23147,N_17648,N_16989);
or U23148 (N_23148,N_16303,N_15985);
xnor U23149 (N_23149,N_18649,N_19712);
xnor U23150 (N_23150,N_15103,N_17912);
xnor U23151 (N_23151,N_16940,N_17944);
nor U23152 (N_23152,N_16689,N_18911);
nor U23153 (N_23153,N_17885,N_19752);
nand U23154 (N_23154,N_18646,N_16252);
nor U23155 (N_23155,N_15998,N_17664);
nand U23156 (N_23156,N_17728,N_15390);
xnor U23157 (N_23157,N_15654,N_18702);
xnor U23158 (N_23158,N_18628,N_16587);
nand U23159 (N_23159,N_18830,N_16283);
nor U23160 (N_23160,N_17389,N_18329);
nor U23161 (N_23161,N_16766,N_18601);
and U23162 (N_23162,N_15715,N_17280);
or U23163 (N_23163,N_15457,N_16422);
xor U23164 (N_23164,N_16284,N_15870);
xor U23165 (N_23165,N_16564,N_16143);
or U23166 (N_23166,N_19916,N_17415);
xor U23167 (N_23167,N_18208,N_18547);
xnor U23168 (N_23168,N_17161,N_17702);
and U23169 (N_23169,N_16503,N_15390);
nor U23170 (N_23170,N_17806,N_15457);
nor U23171 (N_23171,N_19075,N_15666);
nand U23172 (N_23172,N_17534,N_19762);
nor U23173 (N_23173,N_17719,N_15450);
nand U23174 (N_23174,N_16144,N_15417);
and U23175 (N_23175,N_18062,N_16482);
and U23176 (N_23176,N_19814,N_16452);
nand U23177 (N_23177,N_17788,N_19981);
and U23178 (N_23178,N_19324,N_15300);
nand U23179 (N_23179,N_16937,N_16548);
and U23180 (N_23180,N_17020,N_15684);
nand U23181 (N_23181,N_17160,N_19528);
xnor U23182 (N_23182,N_18097,N_15784);
nand U23183 (N_23183,N_16657,N_18987);
nor U23184 (N_23184,N_18897,N_19774);
nand U23185 (N_23185,N_17491,N_18915);
and U23186 (N_23186,N_15286,N_19426);
nor U23187 (N_23187,N_17320,N_18214);
nor U23188 (N_23188,N_18599,N_15483);
nand U23189 (N_23189,N_18546,N_15883);
xor U23190 (N_23190,N_16505,N_15482);
nor U23191 (N_23191,N_17063,N_15112);
and U23192 (N_23192,N_18431,N_19975);
or U23193 (N_23193,N_19369,N_17084);
xor U23194 (N_23194,N_17512,N_15267);
or U23195 (N_23195,N_15404,N_19004);
xnor U23196 (N_23196,N_17355,N_18188);
nor U23197 (N_23197,N_17637,N_16797);
nor U23198 (N_23198,N_17857,N_17983);
nor U23199 (N_23199,N_15607,N_16718);
xnor U23200 (N_23200,N_19157,N_17185);
xnor U23201 (N_23201,N_17874,N_15135);
or U23202 (N_23202,N_19663,N_16395);
nand U23203 (N_23203,N_16281,N_18210);
and U23204 (N_23204,N_18021,N_16485);
xor U23205 (N_23205,N_16172,N_16679);
and U23206 (N_23206,N_15675,N_16097);
xnor U23207 (N_23207,N_15492,N_15872);
xor U23208 (N_23208,N_15179,N_19260);
xnor U23209 (N_23209,N_15937,N_18580);
nand U23210 (N_23210,N_17116,N_16805);
nand U23211 (N_23211,N_16724,N_16643);
and U23212 (N_23212,N_15145,N_18525);
and U23213 (N_23213,N_16684,N_19358);
nor U23214 (N_23214,N_18023,N_16316);
and U23215 (N_23215,N_19850,N_15185);
nor U23216 (N_23216,N_15005,N_19057);
and U23217 (N_23217,N_16794,N_15548);
and U23218 (N_23218,N_18944,N_19573);
and U23219 (N_23219,N_15307,N_16778);
or U23220 (N_23220,N_16917,N_15265);
nor U23221 (N_23221,N_15590,N_18439);
nor U23222 (N_23222,N_19899,N_17519);
and U23223 (N_23223,N_19838,N_18128);
nor U23224 (N_23224,N_18414,N_15762);
xor U23225 (N_23225,N_17672,N_18008);
nor U23226 (N_23226,N_16104,N_15952);
nor U23227 (N_23227,N_17053,N_15343);
nor U23228 (N_23228,N_15674,N_18396);
nor U23229 (N_23229,N_16381,N_19204);
xnor U23230 (N_23230,N_19009,N_17969);
nor U23231 (N_23231,N_17028,N_17126);
or U23232 (N_23232,N_19437,N_19651);
or U23233 (N_23233,N_19729,N_15627);
and U23234 (N_23234,N_18416,N_19042);
xnor U23235 (N_23235,N_18134,N_15623);
xor U23236 (N_23236,N_19571,N_15879);
xor U23237 (N_23237,N_19785,N_16835);
nor U23238 (N_23238,N_18459,N_16146);
xor U23239 (N_23239,N_15841,N_15373);
nor U23240 (N_23240,N_15514,N_19013);
nand U23241 (N_23241,N_18378,N_15052);
xnor U23242 (N_23242,N_17739,N_19300);
nand U23243 (N_23243,N_17775,N_15395);
and U23244 (N_23244,N_16272,N_15781);
xnor U23245 (N_23245,N_19498,N_15132);
nand U23246 (N_23246,N_19550,N_17025);
and U23247 (N_23247,N_17115,N_17345);
and U23248 (N_23248,N_18399,N_18801);
nand U23249 (N_23249,N_19977,N_17917);
nand U23250 (N_23250,N_16168,N_19979);
and U23251 (N_23251,N_19830,N_18187);
and U23252 (N_23252,N_17440,N_19818);
and U23253 (N_23253,N_17709,N_15566);
and U23254 (N_23254,N_16357,N_18190);
xor U23255 (N_23255,N_17832,N_18569);
or U23256 (N_23256,N_15951,N_19112);
nand U23257 (N_23257,N_19867,N_15151);
nor U23258 (N_23258,N_18910,N_15417);
or U23259 (N_23259,N_18809,N_15106);
or U23260 (N_23260,N_17748,N_16561);
and U23261 (N_23261,N_17590,N_18205);
nor U23262 (N_23262,N_17371,N_19904);
nand U23263 (N_23263,N_17094,N_18869);
xnor U23264 (N_23264,N_17494,N_19420);
nand U23265 (N_23265,N_19719,N_19237);
xnor U23266 (N_23266,N_18637,N_19071);
nor U23267 (N_23267,N_15823,N_19953);
xor U23268 (N_23268,N_17538,N_17635);
xor U23269 (N_23269,N_16912,N_19888);
nor U23270 (N_23270,N_18290,N_19225);
and U23271 (N_23271,N_18951,N_16935);
nand U23272 (N_23272,N_15422,N_16627);
and U23273 (N_23273,N_19060,N_17545);
nand U23274 (N_23274,N_17650,N_16829);
and U23275 (N_23275,N_18709,N_19767);
and U23276 (N_23276,N_17066,N_17484);
xnor U23277 (N_23277,N_17617,N_19527);
and U23278 (N_23278,N_16793,N_17795);
and U23279 (N_23279,N_16523,N_17679);
nand U23280 (N_23280,N_16990,N_18783);
xnor U23281 (N_23281,N_15850,N_15012);
or U23282 (N_23282,N_18546,N_15139);
xnor U23283 (N_23283,N_19401,N_15172);
nor U23284 (N_23284,N_15647,N_15549);
and U23285 (N_23285,N_17401,N_18503);
or U23286 (N_23286,N_17979,N_16508);
xor U23287 (N_23287,N_19333,N_16297);
xnor U23288 (N_23288,N_16266,N_15125);
xnor U23289 (N_23289,N_18341,N_18072);
or U23290 (N_23290,N_18348,N_15118);
and U23291 (N_23291,N_15987,N_15222);
or U23292 (N_23292,N_16501,N_17740);
or U23293 (N_23293,N_19670,N_15531);
and U23294 (N_23294,N_15554,N_15228);
nand U23295 (N_23295,N_15105,N_15564);
nand U23296 (N_23296,N_18269,N_17558);
xor U23297 (N_23297,N_15570,N_19050);
nor U23298 (N_23298,N_15756,N_19483);
and U23299 (N_23299,N_17786,N_15946);
nor U23300 (N_23300,N_17699,N_16066);
nand U23301 (N_23301,N_18256,N_15332);
nand U23302 (N_23302,N_15187,N_18285);
nand U23303 (N_23303,N_18447,N_15923);
xor U23304 (N_23304,N_19729,N_18106);
nor U23305 (N_23305,N_19197,N_17209);
and U23306 (N_23306,N_19036,N_19352);
or U23307 (N_23307,N_15421,N_15823);
nand U23308 (N_23308,N_16452,N_15279);
nand U23309 (N_23309,N_15366,N_15477);
nor U23310 (N_23310,N_19300,N_15110);
nand U23311 (N_23311,N_17755,N_17374);
or U23312 (N_23312,N_15445,N_18997);
xnor U23313 (N_23313,N_16916,N_19678);
or U23314 (N_23314,N_17593,N_18280);
nand U23315 (N_23315,N_16810,N_17994);
nand U23316 (N_23316,N_17854,N_17829);
or U23317 (N_23317,N_16780,N_15974);
nand U23318 (N_23318,N_15165,N_17358);
or U23319 (N_23319,N_16793,N_17652);
and U23320 (N_23320,N_19782,N_16186);
and U23321 (N_23321,N_19645,N_16003);
xnor U23322 (N_23322,N_18021,N_18384);
or U23323 (N_23323,N_17941,N_18144);
xor U23324 (N_23324,N_18794,N_18488);
nand U23325 (N_23325,N_19619,N_18367);
xnor U23326 (N_23326,N_18398,N_16691);
or U23327 (N_23327,N_19382,N_19738);
nand U23328 (N_23328,N_15238,N_15459);
or U23329 (N_23329,N_17959,N_18544);
nor U23330 (N_23330,N_16853,N_15713);
or U23331 (N_23331,N_17073,N_18574);
nand U23332 (N_23332,N_18549,N_19593);
or U23333 (N_23333,N_18164,N_18290);
or U23334 (N_23334,N_19038,N_19987);
and U23335 (N_23335,N_15202,N_17706);
and U23336 (N_23336,N_15927,N_17801);
nand U23337 (N_23337,N_17921,N_16143);
and U23338 (N_23338,N_16860,N_18140);
nand U23339 (N_23339,N_17872,N_17562);
or U23340 (N_23340,N_16603,N_15069);
and U23341 (N_23341,N_15890,N_18138);
nand U23342 (N_23342,N_17761,N_17793);
nor U23343 (N_23343,N_15719,N_17612);
xnor U23344 (N_23344,N_17104,N_17069);
xor U23345 (N_23345,N_15842,N_16737);
nor U23346 (N_23346,N_16880,N_17994);
and U23347 (N_23347,N_17247,N_19238);
xnor U23348 (N_23348,N_19222,N_19965);
and U23349 (N_23349,N_17236,N_19388);
nand U23350 (N_23350,N_15445,N_15277);
or U23351 (N_23351,N_15831,N_18422);
xnor U23352 (N_23352,N_17648,N_17194);
and U23353 (N_23353,N_17808,N_17294);
xor U23354 (N_23354,N_18705,N_18585);
or U23355 (N_23355,N_18298,N_15065);
xnor U23356 (N_23356,N_18956,N_19813);
xnor U23357 (N_23357,N_19975,N_15216);
and U23358 (N_23358,N_15278,N_19609);
and U23359 (N_23359,N_17048,N_16241);
nand U23360 (N_23360,N_16415,N_15271);
and U23361 (N_23361,N_17870,N_17864);
and U23362 (N_23362,N_19468,N_15645);
and U23363 (N_23363,N_17547,N_17373);
nor U23364 (N_23364,N_18154,N_16790);
nor U23365 (N_23365,N_18572,N_15329);
nor U23366 (N_23366,N_15769,N_18074);
xnor U23367 (N_23367,N_18656,N_19072);
xor U23368 (N_23368,N_18633,N_15427);
nor U23369 (N_23369,N_17911,N_19266);
xnor U23370 (N_23370,N_19727,N_16579);
nor U23371 (N_23371,N_17941,N_15172);
or U23372 (N_23372,N_16251,N_17870);
nor U23373 (N_23373,N_17299,N_19434);
nand U23374 (N_23374,N_16815,N_15430);
nand U23375 (N_23375,N_15250,N_18678);
xnor U23376 (N_23376,N_15993,N_19847);
nand U23377 (N_23377,N_19147,N_19637);
xor U23378 (N_23378,N_17436,N_18670);
nor U23379 (N_23379,N_15258,N_19375);
and U23380 (N_23380,N_17210,N_18744);
nor U23381 (N_23381,N_18713,N_19498);
or U23382 (N_23382,N_18980,N_17165);
or U23383 (N_23383,N_15041,N_15040);
nor U23384 (N_23384,N_17998,N_16215);
nor U23385 (N_23385,N_18146,N_16692);
nand U23386 (N_23386,N_17525,N_18632);
nand U23387 (N_23387,N_19548,N_17237);
xnor U23388 (N_23388,N_15950,N_17709);
nand U23389 (N_23389,N_19876,N_16412);
nor U23390 (N_23390,N_16255,N_16898);
nand U23391 (N_23391,N_19335,N_19424);
nor U23392 (N_23392,N_19151,N_18883);
nor U23393 (N_23393,N_18956,N_19762);
or U23394 (N_23394,N_19501,N_17280);
nand U23395 (N_23395,N_19507,N_18468);
nand U23396 (N_23396,N_16090,N_15473);
nor U23397 (N_23397,N_19007,N_15925);
and U23398 (N_23398,N_17408,N_16795);
and U23399 (N_23399,N_19010,N_15698);
nand U23400 (N_23400,N_17159,N_19355);
nor U23401 (N_23401,N_18013,N_16135);
nor U23402 (N_23402,N_16313,N_17227);
xnor U23403 (N_23403,N_18260,N_18484);
and U23404 (N_23404,N_16366,N_15837);
and U23405 (N_23405,N_16744,N_18644);
nor U23406 (N_23406,N_19746,N_19538);
nor U23407 (N_23407,N_15371,N_17698);
or U23408 (N_23408,N_15442,N_17389);
xnor U23409 (N_23409,N_15274,N_18990);
nor U23410 (N_23410,N_17198,N_17681);
nor U23411 (N_23411,N_19346,N_17665);
or U23412 (N_23412,N_18008,N_19692);
xor U23413 (N_23413,N_16076,N_16921);
and U23414 (N_23414,N_18629,N_15211);
nand U23415 (N_23415,N_17489,N_15999);
and U23416 (N_23416,N_15454,N_17850);
or U23417 (N_23417,N_16066,N_15601);
nand U23418 (N_23418,N_16387,N_17332);
nor U23419 (N_23419,N_16996,N_15258);
and U23420 (N_23420,N_17747,N_19219);
and U23421 (N_23421,N_19661,N_15133);
or U23422 (N_23422,N_18128,N_16822);
or U23423 (N_23423,N_16195,N_15435);
nand U23424 (N_23424,N_15148,N_16523);
xor U23425 (N_23425,N_18418,N_15363);
xnor U23426 (N_23426,N_17329,N_17224);
nand U23427 (N_23427,N_19731,N_17132);
nor U23428 (N_23428,N_19344,N_16529);
and U23429 (N_23429,N_17117,N_19036);
nor U23430 (N_23430,N_19533,N_15702);
or U23431 (N_23431,N_18491,N_19336);
xnor U23432 (N_23432,N_17708,N_17999);
or U23433 (N_23433,N_17930,N_19875);
nor U23434 (N_23434,N_16291,N_18582);
or U23435 (N_23435,N_15496,N_18285);
nor U23436 (N_23436,N_15988,N_17930);
or U23437 (N_23437,N_15549,N_17157);
nor U23438 (N_23438,N_17155,N_19196);
xor U23439 (N_23439,N_16374,N_19621);
and U23440 (N_23440,N_19564,N_16095);
nor U23441 (N_23441,N_17139,N_15841);
xnor U23442 (N_23442,N_17314,N_19526);
nor U23443 (N_23443,N_16870,N_18376);
nand U23444 (N_23444,N_16473,N_15890);
and U23445 (N_23445,N_19891,N_18330);
and U23446 (N_23446,N_18729,N_17467);
xor U23447 (N_23447,N_17396,N_16672);
or U23448 (N_23448,N_18252,N_18194);
and U23449 (N_23449,N_15585,N_19726);
nor U23450 (N_23450,N_19181,N_18155);
or U23451 (N_23451,N_15157,N_18995);
and U23452 (N_23452,N_16566,N_18834);
and U23453 (N_23453,N_18858,N_18935);
and U23454 (N_23454,N_18363,N_16262);
and U23455 (N_23455,N_18066,N_18183);
xor U23456 (N_23456,N_18685,N_19058);
nor U23457 (N_23457,N_16739,N_17542);
or U23458 (N_23458,N_17212,N_15902);
nand U23459 (N_23459,N_17620,N_17450);
nand U23460 (N_23460,N_17100,N_15146);
xnor U23461 (N_23461,N_15464,N_15567);
and U23462 (N_23462,N_17467,N_16177);
xor U23463 (N_23463,N_17173,N_19713);
xnor U23464 (N_23464,N_18929,N_16905);
nor U23465 (N_23465,N_18399,N_16401);
and U23466 (N_23466,N_19650,N_17360);
and U23467 (N_23467,N_19508,N_17525);
or U23468 (N_23468,N_15159,N_15617);
nor U23469 (N_23469,N_18337,N_15210);
xnor U23470 (N_23470,N_16455,N_16260);
xnor U23471 (N_23471,N_19744,N_19598);
nor U23472 (N_23472,N_16797,N_15634);
and U23473 (N_23473,N_17294,N_16046);
and U23474 (N_23474,N_16875,N_15208);
nand U23475 (N_23475,N_19256,N_17797);
nor U23476 (N_23476,N_19641,N_19816);
nand U23477 (N_23477,N_15498,N_17301);
and U23478 (N_23478,N_16213,N_18275);
nand U23479 (N_23479,N_18943,N_15442);
or U23480 (N_23480,N_17270,N_15074);
xnor U23481 (N_23481,N_19309,N_19208);
nand U23482 (N_23482,N_16427,N_19758);
nor U23483 (N_23483,N_16917,N_16372);
or U23484 (N_23484,N_16340,N_16413);
and U23485 (N_23485,N_19667,N_19894);
xor U23486 (N_23486,N_16402,N_15829);
xnor U23487 (N_23487,N_18934,N_15958);
or U23488 (N_23488,N_19537,N_16914);
nor U23489 (N_23489,N_17773,N_15310);
xnor U23490 (N_23490,N_18773,N_18642);
xor U23491 (N_23491,N_15547,N_18579);
or U23492 (N_23492,N_19625,N_19520);
nor U23493 (N_23493,N_17521,N_17477);
nor U23494 (N_23494,N_15200,N_17126);
nand U23495 (N_23495,N_19428,N_19987);
nand U23496 (N_23496,N_16529,N_15537);
or U23497 (N_23497,N_18534,N_16632);
and U23498 (N_23498,N_18931,N_19131);
nand U23499 (N_23499,N_15213,N_17127);
nor U23500 (N_23500,N_16060,N_19841);
nand U23501 (N_23501,N_18285,N_18639);
or U23502 (N_23502,N_18951,N_18750);
xnor U23503 (N_23503,N_18907,N_18383);
nand U23504 (N_23504,N_18889,N_19100);
or U23505 (N_23505,N_19486,N_15142);
and U23506 (N_23506,N_18444,N_16195);
nor U23507 (N_23507,N_17196,N_15497);
nor U23508 (N_23508,N_16356,N_15585);
nor U23509 (N_23509,N_18187,N_18352);
xnor U23510 (N_23510,N_17040,N_16316);
and U23511 (N_23511,N_17685,N_18263);
or U23512 (N_23512,N_18365,N_18951);
xor U23513 (N_23513,N_17799,N_16991);
or U23514 (N_23514,N_17024,N_18664);
xor U23515 (N_23515,N_19542,N_16436);
xnor U23516 (N_23516,N_15560,N_16981);
and U23517 (N_23517,N_19583,N_16702);
xor U23518 (N_23518,N_17239,N_15406);
and U23519 (N_23519,N_19681,N_18989);
xnor U23520 (N_23520,N_19052,N_19720);
nor U23521 (N_23521,N_16953,N_15728);
nand U23522 (N_23522,N_16825,N_18125);
or U23523 (N_23523,N_16172,N_15843);
or U23524 (N_23524,N_19020,N_16699);
nor U23525 (N_23525,N_18806,N_18423);
and U23526 (N_23526,N_16219,N_18928);
xnor U23527 (N_23527,N_15599,N_17258);
nand U23528 (N_23528,N_19956,N_15250);
nand U23529 (N_23529,N_16367,N_19521);
or U23530 (N_23530,N_16188,N_16393);
or U23531 (N_23531,N_18936,N_15697);
nand U23532 (N_23532,N_15774,N_16043);
xor U23533 (N_23533,N_18578,N_19534);
xnor U23534 (N_23534,N_18677,N_19136);
nor U23535 (N_23535,N_15969,N_19820);
xor U23536 (N_23536,N_18230,N_15320);
nor U23537 (N_23537,N_16088,N_15385);
nand U23538 (N_23538,N_18308,N_15073);
or U23539 (N_23539,N_17275,N_15339);
xor U23540 (N_23540,N_19537,N_19568);
nand U23541 (N_23541,N_18515,N_18318);
and U23542 (N_23542,N_15838,N_16735);
nand U23543 (N_23543,N_15567,N_15171);
xor U23544 (N_23544,N_17625,N_19890);
nand U23545 (N_23545,N_15578,N_18602);
nor U23546 (N_23546,N_16738,N_15456);
or U23547 (N_23547,N_15331,N_18875);
nand U23548 (N_23548,N_16424,N_19471);
nor U23549 (N_23549,N_19540,N_16597);
and U23550 (N_23550,N_16171,N_18659);
or U23551 (N_23551,N_15223,N_19223);
nor U23552 (N_23552,N_19652,N_17689);
nor U23553 (N_23553,N_15512,N_16164);
and U23554 (N_23554,N_17515,N_19523);
or U23555 (N_23555,N_15381,N_17717);
xnor U23556 (N_23556,N_17290,N_15558);
nor U23557 (N_23557,N_19530,N_16187);
or U23558 (N_23558,N_18635,N_17767);
or U23559 (N_23559,N_19793,N_17616);
nand U23560 (N_23560,N_16286,N_16255);
nor U23561 (N_23561,N_19135,N_15217);
and U23562 (N_23562,N_19218,N_16005);
and U23563 (N_23563,N_19913,N_16042);
nand U23564 (N_23564,N_15965,N_17798);
and U23565 (N_23565,N_16089,N_19054);
and U23566 (N_23566,N_15132,N_15742);
and U23567 (N_23567,N_18309,N_18847);
nor U23568 (N_23568,N_17922,N_16199);
or U23569 (N_23569,N_19076,N_17643);
xnor U23570 (N_23570,N_16756,N_19543);
nor U23571 (N_23571,N_19107,N_19202);
nor U23572 (N_23572,N_17667,N_17615);
nor U23573 (N_23573,N_19752,N_19537);
nor U23574 (N_23574,N_18688,N_16473);
xnor U23575 (N_23575,N_17366,N_18091);
nand U23576 (N_23576,N_16019,N_16476);
xor U23577 (N_23577,N_19231,N_18403);
xnor U23578 (N_23578,N_19204,N_17610);
or U23579 (N_23579,N_18181,N_19114);
nor U23580 (N_23580,N_17312,N_17479);
nor U23581 (N_23581,N_15920,N_17891);
nor U23582 (N_23582,N_18722,N_19687);
nand U23583 (N_23583,N_16855,N_17543);
or U23584 (N_23584,N_19320,N_19163);
and U23585 (N_23585,N_17444,N_15465);
xnor U23586 (N_23586,N_16545,N_19083);
or U23587 (N_23587,N_15540,N_15879);
xnor U23588 (N_23588,N_15487,N_19148);
and U23589 (N_23589,N_17143,N_16022);
or U23590 (N_23590,N_16996,N_19698);
or U23591 (N_23591,N_15611,N_19588);
nand U23592 (N_23592,N_19745,N_19921);
or U23593 (N_23593,N_16617,N_16902);
nor U23594 (N_23594,N_19437,N_18945);
and U23595 (N_23595,N_18587,N_18820);
nand U23596 (N_23596,N_18781,N_17199);
xnor U23597 (N_23597,N_19438,N_19086);
xnor U23598 (N_23598,N_17994,N_15907);
and U23599 (N_23599,N_19827,N_16838);
or U23600 (N_23600,N_18988,N_16642);
and U23601 (N_23601,N_18859,N_17557);
xor U23602 (N_23602,N_16153,N_16054);
or U23603 (N_23603,N_18349,N_17037);
or U23604 (N_23604,N_18942,N_17288);
or U23605 (N_23605,N_15027,N_17573);
nand U23606 (N_23606,N_19326,N_18339);
or U23607 (N_23607,N_19769,N_15115);
nand U23608 (N_23608,N_15982,N_17531);
and U23609 (N_23609,N_15050,N_16663);
nor U23610 (N_23610,N_16185,N_16271);
and U23611 (N_23611,N_17350,N_15545);
or U23612 (N_23612,N_18640,N_19642);
and U23613 (N_23613,N_17703,N_17916);
xnor U23614 (N_23614,N_15649,N_16690);
and U23615 (N_23615,N_19665,N_17238);
nor U23616 (N_23616,N_16982,N_19230);
nand U23617 (N_23617,N_17162,N_17194);
and U23618 (N_23618,N_19785,N_16954);
nand U23619 (N_23619,N_18554,N_16027);
nor U23620 (N_23620,N_16976,N_19102);
nor U23621 (N_23621,N_19027,N_15425);
nand U23622 (N_23622,N_15526,N_15432);
or U23623 (N_23623,N_18021,N_17622);
nor U23624 (N_23624,N_17649,N_17461);
nor U23625 (N_23625,N_18415,N_15333);
nor U23626 (N_23626,N_15417,N_19569);
or U23627 (N_23627,N_18647,N_16263);
nor U23628 (N_23628,N_18953,N_18595);
or U23629 (N_23629,N_17192,N_17209);
xnor U23630 (N_23630,N_15710,N_16524);
xor U23631 (N_23631,N_15483,N_15590);
nor U23632 (N_23632,N_16629,N_18850);
and U23633 (N_23633,N_15099,N_15688);
and U23634 (N_23634,N_17475,N_19199);
nand U23635 (N_23635,N_16661,N_15932);
or U23636 (N_23636,N_19318,N_18267);
and U23637 (N_23637,N_17997,N_15138);
and U23638 (N_23638,N_19673,N_15765);
nand U23639 (N_23639,N_16971,N_19719);
nand U23640 (N_23640,N_18987,N_18483);
nand U23641 (N_23641,N_19920,N_18543);
and U23642 (N_23642,N_19714,N_18930);
and U23643 (N_23643,N_15914,N_18684);
xnor U23644 (N_23644,N_15902,N_19039);
xor U23645 (N_23645,N_19650,N_15543);
or U23646 (N_23646,N_19185,N_16656);
nor U23647 (N_23647,N_17954,N_18610);
xor U23648 (N_23648,N_16316,N_19473);
nor U23649 (N_23649,N_17924,N_19044);
nor U23650 (N_23650,N_18559,N_18685);
nand U23651 (N_23651,N_18252,N_18586);
and U23652 (N_23652,N_16958,N_18188);
and U23653 (N_23653,N_15365,N_15065);
nor U23654 (N_23654,N_18672,N_17517);
and U23655 (N_23655,N_17679,N_18819);
nor U23656 (N_23656,N_15033,N_15256);
and U23657 (N_23657,N_18081,N_19821);
and U23658 (N_23658,N_16403,N_17835);
or U23659 (N_23659,N_18877,N_18405);
nand U23660 (N_23660,N_15031,N_17767);
or U23661 (N_23661,N_16214,N_15569);
xnor U23662 (N_23662,N_18177,N_18978);
nand U23663 (N_23663,N_15789,N_15909);
xnor U23664 (N_23664,N_16602,N_18814);
nand U23665 (N_23665,N_19173,N_15235);
or U23666 (N_23666,N_18052,N_16868);
or U23667 (N_23667,N_18994,N_19085);
xor U23668 (N_23668,N_18290,N_17816);
or U23669 (N_23669,N_16619,N_16477);
and U23670 (N_23670,N_19019,N_17774);
or U23671 (N_23671,N_17554,N_15806);
xor U23672 (N_23672,N_16404,N_17694);
xor U23673 (N_23673,N_19841,N_15468);
or U23674 (N_23674,N_15135,N_15578);
or U23675 (N_23675,N_16636,N_15356);
and U23676 (N_23676,N_16838,N_15778);
nor U23677 (N_23677,N_19000,N_18290);
and U23678 (N_23678,N_19004,N_16916);
or U23679 (N_23679,N_17377,N_16676);
and U23680 (N_23680,N_17639,N_18959);
xor U23681 (N_23681,N_19233,N_15705);
and U23682 (N_23682,N_19823,N_17707);
or U23683 (N_23683,N_17635,N_18960);
nand U23684 (N_23684,N_16049,N_16246);
or U23685 (N_23685,N_18699,N_15519);
xnor U23686 (N_23686,N_17396,N_17385);
nand U23687 (N_23687,N_17551,N_16175);
xor U23688 (N_23688,N_17930,N_18583);
nand U23689 (N_23689,N_16682,N_16763);
and U23690 (N_23690,N_15781,N_15210);
nor U23691 (N_23691,N_16919,N_18923);
or U23692 (N_23692,N_17996,N_18136);
nor U23693 (N_23693,N_15608,N_16892);
xor U23694 (N_23694,N_18286,N_18625);
nand U23695 (N_23695,N_17379,N_18344);
nor U23696 (N_23696,N_17655,N_18859);
nor U23697 (N_23697,N_18215,N_18600);
or U23698 (N_23698,N_19611,N_16833);
and U23699 (N_23699,N_16549,N_18025);
nand U23700 (N_23700,N_16498,N_19765);
xnor U23701 (N_23701,N_18504,N_17152);
xor U23702 (N_23702,N_18604,N_16378);
and U23703 (N_23703,N_18774,N_17958);
and U23704 (N_23704,N_17142,N_17276);
nand U23705 (N_23705,N_17953,N_19494);
or U23706 (N_23706,N_17030,N_19090);
nand U23707 (N_23707,N_18323,N_16329);
nand U23708 (N_23708,N_19936,N_15450);
xnor U23709 (N_23709,N_16688,N_15437);
nand U23710 (N_23710,N_17696,N_15920);
nor U23711 (N_23711,N_15395,N_19956);
nor U23712 (N_23712,N_16474,N_19150);
nand U23713 (N_23713,N_19378,N_17271);
nand U23714 (N_23714,N_17128,N_16840);
or U23715 (N_23715,N_18608,N_17804);
nor U23716 (N_23716,N_17508,N_16581);
xor U23717 (N_23717,N_17694,N_19556);
nor U23718 (N_23718,N_15290,N_19301);
nor U23719 (N_23719,N_15730,N_18451);
or U23720 (N_23720,N_16554,N_15277);
xnor U23721 (N_23721,N_17388,N_19112);
and U23722 (N_23722,N_16304,N_16960);
or U23723 (N_23723,N_19180,N_17942);
xnor U23724 (N_23724,N_18449,N_15222);
and U23725 (N_23725,N_18809,N_17182);
or U23726 (N_23726,N_18206,N_19239);
and U23727 (N_23727,N_18540,N_18785);
nand U23728 (N_23728,N_17798,N_16901);
nand U23729 (N_23729,N_18215,N_16025);
nand U23730 (N_23730,N_16359,N_16030);
nor U23731 (N_23731,N_17886,N_16195);
or U23732 (N_23732,N_18758,N_17397);
and U23733 (N_23733,N_16005,N_15021);
or U23734 (N_23734,N_19488,N_18212);
nor U23735 (N_23735,N_18327,N_19426);
nor U23736 (N_23736,N_17005,N_19644);
xor U23737 (N_23737,N_17374,N_19498);
nor U23738 (N_23738,N_17145,N_16162);
and U23739 (N_23739,N_18412,N_19427);
and U23740 (N_23740,N_18724,N_15984);
or U23741 (N_23741,N_19056,N_16422);
or U23742 (N_23742,N_17258,N_16143);
nand U23743 (N_23743,N_19865,N_17219);
or U23744 (N_23744,N_19216,N_16963);
and U23745 (N_23745,N_19274,N_18739);
nor U23746 (N_23746,N_17325,N_16440);
xor U23747 (N_23747,N_17102,N_18810);
nor U23748 (N_23748,N_16919,N_16191);
nand U23749 (N_23749,N_18520,N_19232);
nor U23750 (N_23750,N_16195,N_17148);
and U23751 (N_23751,N_17111,N_16062);
nand U23752 (N_23752,N_18172,N_15428);
or U23753 (N_23753,N_16824,N_17899);
nor U23754 (N_23754,N_16920,N_19002);
nor U23755 (N_23755,N_16044,N_19621);
nand U23756 (N_23756,N_16136,N_16999);
nor U23757 (N_23757,N_18004,N_16645);
or U23758 (N_23758,N_19058,N_17127);
xnor U23759 (N_23759,N_18009,N_18505);
or U23760 (N_23760,N_17079,N_17325);
nand U23761 (N_23761,N_17860,N_15208);
xnor U23762 (N_23762,N_17259,N_19581);
nand U23763 (N_23763,N_19110,N_19939);
xnor U23764 (N_23764,N_16914,N_18317);
xnor U23765 (N_23765,N_19990,N_15148);
or U23766 (N_23766,N_19587,N_18384);
or U23767 (N_23767,N_16367,N_15371);
xnor U23768 (N_23768,N_18363,N_17008);
xor U23769 (N_23769,N_17052,N_17945);
or U23770 (N_23770,N_15963,N_16073);
nand U23771 (N_23771,N_17630,N_18033);
and U23772 (N_23772,N_18761,N_17881);
or U23773 (N_23773,N_19007,N_17579);
nand U23774 (N_23774,N_17907,N_15223);
and U23775 (N_23775,N_19498,N_16053);
nand U23776 (N_23776,N_19368,N_19729);
nor U23777 (N_23777,N_16567,N_16954);
or U23778 (N_23778,N_16082,N_16478);
xnor U23779 (N_23779,N_18110,N_18817);
and U23780 (N_23780,N_15368,N_15824);
or U23781 (N_23781,N_17967,N_17884);
nand U23782 (N_23782,N_18158,N_18580);
xnor U23783 (N_23783,N_17806,N_16078);
nor U23784 (N_23784,N_16901,N_15426);
nor U23785 (N_23785,N_16481,N_18096);
nor U23786 (N_23786,N_18245,N_19706);
nand U23787 (N_23787,N_19216,N_18359);
xnor U23788 (N_23788,N_18386,N_17696);
nor U23789 (N_23789,N_18389,N_17177);
nor U23790 (N_23790,N_15569,N_17428);
and U23791 (N_23791,N_18545,N_18011);
and U23792 (N_23792,N_19767,N_19904);
xnor U23793 (N_23793,N_18890,N_16484);
nand U23794 (N_23794,N_19653,N_19608);
xnor U23795 (N_23795,N_17949,N_18421);
nand U23796 (N_23796,N_18079,N_15607);
and U23797 (N_23797,N_18646,N_17525);
nand U23798 (N_23798,N_19571,N_18609);
and U23799 (N_23799,N_18515,N_16094);
nor U23800 (N_23800,N_16210,N_19955);
and U23801 (N_23801,N_18846,N_16941);
nand U23802 (N_23802,N_15839,N_18609);
xnor U23803 (N_23803,N_15369,N_15914);
xnor U23804 (N_23804,N_17822,N_16431);
and U23805 (N_23805,N_19175,N_19851);
nand U23806 (N_23806,N_16771,N_16348);
nor U23807 (N_23807,N_16560,N_17183);
and U23808 (N_23808,N_16386,N_16826);
xnor U23809 (N_23809,N_15034,N_16238);
or U23810 (N_23810,N_17817,N_16391);
xnor U23811 (N_23811,N_15023,N_17908);
and U23812 (N_23812,N_18817,N_19442);
and U23813 (N_23813,N_19042,N_19475);
nor U23814 (N_23814,N_16216,N_17543);
or U23815 (N_23815,N_18168,N_17884);
xnor U23816 (N_23816,N_15716,N_19091);
nor U23817 (N_23817,N_16492,N_16005);
xnor U23818 (N_23818,N_19296,N_16557);
or U23819 (N_23819,N_18899,N_19846);
xnor U23820 (N_23820,N_15562,N_17088);
nand U23821 (N_23821,N_17539,N_15300);
or U23822 (N_23822,N_16502,N_19640);
xor U23823 (N_23823,N_15539,N_18176);
and U23824 (N_23824,N_17770,N_19141);
xnor U23825 (N_23825,N_18009,N_15072);
xnor U23826 (N_23826,N_16810,N_16417);
or U23827 (N_23827,N_15475,N_18085);
nor U23828 (N_23828,N_16341,N_15513);
and U23829 (N_23829,N_17348,N_19139);
and U23830 (N_23830,N_19891,N_17796);
and U23831 (N_23831,N_19612,N_19100);
nand U23832 (N_23832,N_17159,N_15697);
xnor U23833 (N_23833,N_17590,N_15333);
or U23834 (N_23834,N_17361,N_19477);
xnor U23835 (N_23835,N_16511,N_16899);
nand U23836 (N_23836,N_16085,N_16895);
and U23837 (N_23837,N_18313,N_17413);
nand U23838 (N_23838,N_15557,N_16462);
and U23839 (N_23839,N_16003,N_19164);
xor U23840 (N_23840,N_18847,N_19202);
xnor U23841 (N_23841,N_16643,N_16740);
nand U23842 (N_23842,N_17424,N_19101);
nand U23843 (N_23843,N_16150,N_16260);
and U23844 (N_23844,N_15516,N_15146);
nor U23845 (N_23845,N_15253,N_17494);
and U23846 (N_23846,N_15576,N_18122);
and U23847 (N_23847,N_18885,N_19714);
xor U23848 (N_23848,N_16962,N_19031);
nor U23849 (N_23849,N_19412,N_19094);
and U23850 (N_23850,N_15810,N_17163);
and U23851 (N_23851,N_16335,N_19636);
and U23852 (N_23852,N_15263,N_18128);
nand U23853 (N_23853,N_18980,N_17747);
nand U23854 (N_23854,N_19303,N_19847);
xor U23855 (N_23855,N_15239,N_16285);
nand U23856 (N_23856,N_15509,N_17765);
or U23857 (N_23857,N_17699,N_18041);
nor U23858 (N_23858,N_15589,N_15538);
or U23859 (N_23859,N_15705,N_19320);
nand U23860 (N_23860,N_15066,N_17518);
nor U23861 (N_23861,N_16279,N_15928);
nor U23862 (N_23862,N_15249,N_19294);
nor U23863 (N_23863,N_19862,N_17533);
and U23864 (N_23864,N_19400,N_19087);
xor U23865 (N_23865,N_16528,N_18775);
xor U23866 (N_23866,N_16716,N_17914);
or U23867 (N_23867,N_16454,N_15955);
xnor U23868 (N_23868,N_18103,N_15989);
nand U23869 (N_23869,N_17735,N_18449);
and U23870 (N_23870,N_17140,N_16053);
nand U23871 (N_23871,N_19566,N_17609);
and U23872 (N_23872,N_19864,N_18506);
and U23873 (N_23873,N_16176,N_17695);
or U23874 (N_23874,N_15142,N_16834);
nand U23875 (N_23875,N_19859,N_18152);
nand U23876 (N_23876,N_17195,N_15283);
nand U23877 (N_23877,N_16470,N_16762);
nand U23878 (N_23878,N_15461,N_18100);
nand U23879 (N_23879,N_18675,N_19287);
or U23880 (N_23880,N_18856,N_17687);
nand U23881 (N_23881,N_15445,N_16670);
or U23882 (N_23882,N_17285,N_17598);
nor U23883 (N_23883,N_17384,N_15676);
and U23884 (N_23884,N_19718,N_18707);
nor U23885 (N_23885,N_15140,N_19855);
nor U23886 (N_23886,N_19242,N_15780);
nand U23887 (N_23887,N_18096,N_19271);
and U23888 (N_23888,N_16439,N_18360);
or U23889 (N_23889,N_19916,N_16590);
or U23890 (N_23890,N_16345,N_15002);
and U23891 (N_23891,N_19759,N_16675);
xor U23892 (N_23892,N_16579,N_19121);
nor U23893 (N_23893,N_18315,N_15473);
nand U23894 (N_23894,N_19646,N_18843);
and U23895 (N_23895,N_19520,N_19096);
and U23896 (N_23896,N_17628,N_16365);
and U23897 (N_23897,N_18498,N_16649);
xnor U23898 (N_23898,N_17323,N_19679);
nand U23899 (N_23899,N_17069,N_16474);
or U23900 (N_23900,N_18473,N_16244);
xor U23901 (N_23901,N_17124,N_17002);
nor U23902 (N_23902,N_15986,N_19406);
xor U23903 (N_23903,N_18240,N_16990);
nor U23904 (N_23904,N_19897,N_18852);
and U23905 (N_23905,N_18017,N_15495);
or U23906 (N_23906,N_16803,N_15507);
and U23907 (N_23907,N_19611,N_18505);
nand U23908 (N_23908,N_18712,N_19030);
nor U23909 (N_23909,N_18077,N_18714);
or U23910 (N_23910,N_17122,N_19354);
xor U23911 (N_23911,N_16935,N_16409);
nor U23912 (N_23912,N_19653,N_17737);
xnor U23913 (N_23913,N_15048,N_19661);
and U23914 (N_23914,N_15689,N_18565);
and U23915 (N_23915,N_16729,N_19650);
and U23916 (N_23916,N_18472,N_16874);
and U23917 (N_23917,N_19264,N_17874);
or U23918 (N_23918,N_16254,N_16528);
xor U23919 (N_23919,N_18495,N_17606);
xor U23920 (N_23920,N_17629,N_16390);
nand U23921 (N_23921,N_15905,N_16798);
nor U23922 (N_23922,N_18482,N_16143);
and U23923 (N_23923,N_17616,N_18138);
and U23924 (N_23924,N_18724,N_15852);
xor U23925 (N_23925,N_15113,N_15947);
and U23926 (N_23926,N_18623,N_17201);
or U23927 (N_23927,N_17267,N_16887);
xnor U23928 (N_23928,N_18248,N_17593);
and U23929 (N_23929,N_16270,N_16143);
xor U23930 (N_23930,N_15678,N_15984);
xor U23931 (N_23931,N_19544,N_16179);
and U23932 (N_23932,N_17482,N_16570);
xor U23933 (N_23933,N_18000,N_16932);
nor U23934 (N_23934,N_18523,N_16978);
or U23935 (N_23935,N_15193,N_19268);
xnor U23936 (N_23936,N_19745,N_19352);
or U23937 (N_23937,N_17448,N_19301);
or U23938 (N_23938,N_18819,N_19169);
nor U23939 (N_23939,N_17648,N_15736);
and U23940 (N_23940,N_18937,N_18205);
nor U23941 (N_23941,N_15129,N_17685);
and U23942 (N_23942,N_18034,N_19574);
nor U23943 (N_23943,N_15110,N_19923);
and U23944 (N_23944,N_18583,N_19503);
or U23945 (N_23945,N_18454,N_18908);
xnor U23946 (N_23946,N_17085,N_16537);
nand U23947 (N_23947,N_15712,N_18994);
or U23948 (N_23948,N_17458,N_18502);
nand U23949 (N_23949,N_18582,N_19719);
nand U23950 (N_23950,N_16651,N_15308);
nand U23951 (N_23951,N_18287,N_19881);
nor U23952 (N_23952,N_17630,N_17738);
and U23953 (N_23953,N_16990,N_19649);
xor U23954 (N_23954,N_16779,N_19331);
and U23955 (N_23955,N_15707,N_15639);
and U23956 (N_23956,N_15903,N_16149);
or U23957 (N_23957,N_16745,N_16223);
or U23958 (N_23958,N_17953,N_18263);
nor U23959 (N_23959,N_15705,N_15204);
nand U23960 (N_23960,N_16608,N_18409);
and U23961 (N_23961,N_15952,N_19025);
or U23962 (N_23962,N_16784,N_18202);
and U23963 (N_23963,N_18136,N_17339);
and U23964 (N_23964,N_16084,N_15908);
and U23965 (N_23965,N_18953,N_15653);
xnor U23966 (N_23966,N_18320,N_17089);
nor U23967 (N_23967,N_17849,N_16900);
or U23968 (N_23968,N_19892,N_15081);
or U23969 (N_23969,N_19552,N_15975);
and U23970 (N_23970,N_17707,N_16737);
or U23971 (N_23971,N_15797,N_17561);
and U23972 (N_23972,N_18085,N_16833);
and U23973 (N_23973,N_15407,N_18428);
or U23974 (N_23974,N_17593,N_17927);
and U23975 (N_23975,N_16887,N_17555);
or U23976 (N_23976,N_18120,N_16355);
nand U23977 (N_23977,N_18546,N_18845);
xnor U23978 (N_23978,N_17091,N_16812);
nor U23979 (N_23979,N_18344,N_16406);
nand U23980 (N_23980,N_15551,N_19020);
or U23981 (N_23981,N_17721,N_16266);
or U23982 (N_23982,N_19072,N_15975);
or U23983 (N_23983,N_17414,N_18383);
nand U23984 (N_23984,N_19196,N_15027);
and U23985 (N_23985,N_15197,N_16588);
and U23986 (N_23986,N_15007,N_17700);
xnor U23987 (N_23987,N_16667,N_19906);
and U23988 (N_23988,N_16378,N_16240);
and U23989 (N_23989,N_15003,N_17123);
xor U23990 (N_23990,N_15118,N_18760);
or U23991 (N_23991,N_18220,N_16330);
or U23992 (N_23992,N_19522,N_18810);
or U23993 (N_23993,N_18698,N_16540);
nand U23994 (N_23994,N_16742,N_18925);
and U23995 (N_23995,N_19397,N_17796);
xor U23996 (N_23996,N_16401,N_15944);
xor U23997 (N_23997,N_19698,N_16092);
xor U23998 (N_23998,N_16540,N_16722);
and U23999 (N_23999,N_15220,N_18813);
xnor U24000 (N_24000,N_15605,N_17439);
and U24001 (N_24001,N_16953,N_16763);
nor U24002 (N_24002,N_15708,N_18306);
and U24003 (N_24003,N_19061,N_17128);
xor U24004 (N_24004,N_19970,N_19675);
nor U24005 (N_24005,N_18232,N_17436);
nor U24006 (N_24006,N_15111,N_17389);
nand U24007 (N_24007,N_18921,N_18657);
nand U24008 (N_24008,N_16402,N_16261);
or U24009 (N_24009,N_19635,N_19211);
nand U24010 (N_24010,N_16609,N_16182);
and U24011 (N_24011,N_18316,N_18578);
nand U24012 (N_24012,N_15518,N_16470);
xnor U24013 (N_24013,N_19088,N_18910);
or U24014 (N_24014,N_18830,N_19331);
nor U24015 (N_24015,N_18624,N_15861);
nor U24016 (N_24016,N_19635,N_17626);
nand U24017 (N_24017,N_15821,N_18402);
and U24018 (N_24018,N_17752,N_17804);
and U24019 (N_24019,N_15494,N_15724);
xor U24020 (N_24020,N_17849,N_15652);
nor U24021 (N_24021,N_19041,N_17703);
or U24022 (N_24022,N_19043,N_18905);
or U24023 (N_24023,N_16990,N_19658);
or U24024 (N_24024,N_19108,N_16286);
nand U24025 (N_24025,N_15078,N_19824);
and U24026 (N_24026,N_15484,N_17845);
nor U24027 (N_24027,N_18232,N_19651);
and U24028 (N_24028,N_18346,N_18903);
nor U24029 (N_24029,N_15719,N_15303);
or U24030 (N_24030,N_15059,N_15183);
nand U24031 (N_24031,N_17402,N_19784);
or U24032 (N_24032,N_18172,N_19576);
nor U24033 (N_24033,N_16743,N_16154);
or U24034 (N_24034,N_17362,N_19215);
nor U24035 (N_24035,N_17304,N_19194);
nor U24036 (N_24036,N_18067,N_17883);
or U24037 (N_24037,N_19810,N_15426);
or U24038 (N_24038,N_18064,N_17320);
nand U24039 (N_24039,N_15388,N_15975);
nand U24040 (N_24040,N_18889,N_16011);
nor U24041 (N_24041,N_19435,N_16330);
and U24042 (N_24042,N_19332,N_16372);
or U24043 (N_24043,N_19445,N_19392);
and U24044 (N_24044,N_17584,N_15283);
xnor U24045 (N_24045,N_18183,N_19186);
nand U24046 (N_24046,N_16536,N_16725);
nor U24047 (N_24047,N_15667,N_17750);
and U24048 (N_24048,N_19106,N_18981);
nand U24049 (N_24049,N_15485,N_15008);
or U24050 (N_24050,N_18692,N_15680);
nand U24051 (N_24051,N_18940,N_18838);
xor U24052 (N_24052,N_15810,N_15738);
xor U24053 (N_24053,N_15537,N_18815);
and U24054 (N_24054,N_17000,N_16457);
and U24055 (N_24055,N_19267,N_19634);
nand U24056 (N_24056,N_18791,N_15568);
nor U24057 (N_24057,N_18562,N_18757);
or U24058 (N_24058,N_16172,N_15431);
nand U24059 (N_24059,N_17954,N_16358);
xor U24060 (N_24060,N_17271,N_17096);
and U24061 (N_24061,N_18554,N_17555);
nand U24062 (N_24062,N_16202,N_16920);
xor U24063 (N_24063,N_17926,N_16554);
nand U24064 (N_24064,N_18099,N_16422);
nand U24065 (N_24065,N_16529,N_18001);
xor U24066 (N_24066,N_19994,N_18975);
nor U24067 (N_24067,N_15202,N_15756);
nor U24068 (N_24068,N_15982,N_19831);
or U24069 (N_24069,N_18187,N_16263);
and U24070 (N_24070,N_16475,N_17822);
and U24071 (N_24071,N_18209,N_15058);
xor U24072 (N_24072,N_17283,N_15598);
xor U24073 (N_24073,N_15902,N_15540);
nand U24074 (N_24074,N_15746,N_17515);
xnor U24075 (N_24075,N_17861,N_17125);
or U24076 (N_24076,N_17502,N_19400);
and U24077 (N_24077,N_15967,N_17708);
nand U24078 (N_24078,N_17076,N_17941);
and U24079 (N_24079,N_15899,N_16651);
nand U24080 (N_24080,N_18248,N_16523);
xor U24081 (N_24081,N_16011,N_17311);
and U24082 (N_24082,N_18088,N_17692);
xor U24083 (N_24083,N_19948,N_19424);
nor U24084 (N_24084,N_17900,N_16632);
nand U24085 (N_24085,N_17881,N_18624);
nand U24086 (N_24086,N_18185,N_16457);
xor U24087 (N_24087,N_17484,N_17438);
nor U24088 (N_24088,N_17385,N_18285);
xor U24089 (N_24089,N_19979,N_16241);
and U24090 (N_24090,N_17353,N_19656);
nand U24091 (N_24091,N_15461,N_16226);
xnor U24092 (N_24092,N_19175,N_16105);
and U24093 (N_24093,N_18674,N_16058);
and U24094 (N_24094,N_15596,N_19852);
xnor U24095 (N_24095,N_17905,N_18757);
and U24096 (N_24096,N_19330,N_17195);
nor U24097 (N_24097,N_16405,N_18666);
and U24098 (N_24098,N_18706,N_17846);
or U24099 (N_24099,N_18088,N_18261);
xor U24100 (N_24100,N_18371,N_19801);
xnor U24101 (N_24101,N_19391,N_17506);
and U24102 (N_24102,N_16456,N_15228);
and U24103 (N_24103,N_15977,N_19619);
nor U24104 (N_24104,N_19786,N_19240);
or U24105 (N_24105,N_19876,N_15303);
xnor U24106 (N_24106,N_16675,N_16924);
nor U24107 (N_24107,N_16629,N_15952);
xor U24108 (N_24108,N_17830,N_19265);
or U24109 (N_24109,N_17685,N_18968);
xnor U24110 (N_24110,N_19739,N_18972);
or U24111 (N_24111,N_16915,N_16474);
nor U24112 (N_24112,N_17283,N_18829);
xnor U24113 (N_24113,N_18608,N_18784);
nor U24114 (N_24114,N_16137,N_17982);
nand U24115 (N_24115,N_19002,N_15998);
and U24116 (N_24116,N_16140,N_17027);
or U24117 (N_24117,N_19287,N_18802);
or U24118 (N_24118,N_15168,N_16637);
or U24119 (N_24119,N_16143,N_19503);
and U24120 (N_24120,N_17559,N_15746);
and U24121 (N_24121,N_19441,N_17987);
or U24122 (N_24122,N_17619,N_18427);
or U24123 (N_24123,N_17845,N_15868);
xor U24124 (N_24124,N_18412,N_15594);
xnor U24125 (N_24125,N_16885,N_16242);
or U24126 (N_24126,N_18561,N_19952);
and U24127 (N_24127,N_18080,N_17206);
xnor U24128 (N_24128,N_16393,N_18440);
xnor U24129 (N_24129,N_19300,N_18017);
nand U24130 (N_24130,N_17301,N_18832);
or U24131 (N_24131,N_19307,N_18457);
nand U24132 (N_24132,N_16733,N_18532);
or U24133 (N_24133,N_16794,N_15274);
and U24134 (N_24134,N_16868,N_19949);
or U24135 (N_24135,N_17424,N_15946);
xnor U24136 (N_24136,N_15610,N_18467);
xor U24137 (N_24137,N_17439,N_17344);
nor U24138 (N_24138,N_15696,N_16055);
nand U24139 (N_24139,N_16003,N_16930);
xnor U24140 (N_24140,N_17913,N_15868);
nor U24141 (N_24141,N_16823,N_18726);
nand U24142 (N_24142,N_18165,N_15988);
nor U24143 (N_24143,N_16991,N_18180);
nor U24144 (N_24144,N_16983,N_15370);
nand U24145 (N_24145,N_15559,N_15184);
xnor U24146 (N_24146,N_16955,N_18281);
xor U24147 (N_24147,N_18227,N_15450);
nor U24148 (N_24148,N_19212,N_17918);
or U24149 (N_24149,N_16804,N_16561);
or U24150 (N_24150,N_19434,N_16608);
nor U24151 (N_24151,N_18017,N_19222);
or U24152 (N_24152,N_15743,N_17901);
and U24153 (N_24153,N_19544,N_19371);
and U24154 (N_24154,N_16264,N_15168);
nor U24155 (N_24155,N_18345,N_17277);
xnor U24156 (N_24156,N_19606,N_16354);
nand U24157 (N_24157,N_18539,N_18360);
xor U24158 (N_24158,N_17338,N_15843);
nand U24159 (N_24159,N_19780,N_18361);
and U24160 (N_24160,N_15454,N_19883);
nor U24161 (N_24161,N_17452,N_19709);
nor U24162 (N_24162,N_15050,N_19412);
or U24163 (N_24163,N_19591,N_17151);
nor U24164 (N_24164,N_16714,N_17461);
and U24165 (N_24165,N_15856,N_18562);
nor U24166 (N_24166,N_19919,N_19137);
nand U24167 (N_24167,N_19064,N_19940);
and U24168 (N_24168,N_17480,N_19786);
nor U24169 (N_24169,N_19816,N_19711);
or U24170 (N_24170,N_19964,N_15042);
and U24171 (N_24171,N_19468,N_17142);
and U24172 (N_24172,N_15560,N_18250);
nor U24173 (N_24173,N_19426,N_16015);
and U24174 (N_24174,N_16670,N_19829);
nor U24175 (N_24175,N_16637,N_19707);
nand U24176 (N_24176,N_18816,N_18773);
nor U24177 (N_24177,N_17353,N_18598);
nand U24178 (N_24178,N_17705,N_15370);
nand U24179 (N_24179,N_16671,N_15405);
and U24180 (N_24180,N_17305,N_18365);
nand U24181 (N_24181,N_15137,N_18115);
xnor U24182 (N_24182,N_16808,N_16100);
xor U24183 (N_24183,N_15772,N_18894);
nand U24184 (N_24184,N_18703,N_18339);
or U24185 (N_24185,N_16461,N_15025);
nand U24186 (N_24186,N_17828,N_17607);
or U24187 (N_24187,N_15314,N_15802);
nor U24188 (N_24188,N_16980,N_15276);
nor U24189 (N_24189,N_19311,N_17544);
xnor U24190 (N_24190,N_19896,N_18508);
xnor U24191 (N_24191,N_18405,N_16565);
nand U24192 (N_24192,N_17758,N_18687);
and U24193 (N_24193,N_17990,N_19274);
nand U24194 (N_24194,N_16333,N_19043);
nor U24195 (N_24195,N_17479,N_15912);
and U24196 (N_24196,N_15908,N_18867);
nand U24197 (N_24197,N_18730,N_15713);
nor U24198 (N_24198,N_15208,N_16294);
nor U24199 (N_24199,N_19429,N_18352);
nand U24200 (N_24200,N_17655,N_18187);
nor U24201 (N_24201,N_18407,N_18672);
xnor U24202 (N_24202,N_17045,N_18670);
or U24203 (N_24203,N_19810,N_17787);
nand U24204 (N_24204,N_17785,N_19764);
nor U24205 (N_24205,N_17096,N_18468);
xor U24206 (N_24206,N_15381,N_15405);
nor U24207 (N_24207,N_17937,N_19571);
nand U24208 (N_24208,N_17733,N_18585);
nor U24209 (N_24209,N_19720,N_17422);
nor U24210 (N_24210,N_15673,N_19203);
xnor U24211 (N_24211,N_18646,N_19790);
nor U24212 (N_24212,N_18142,N_15518);
xor U24213 (N_24213,N_17612,N_18956);
or U24214 (N_24214,N_19778,N_15245);
and U24215 (N_24215,N_16934,N_15875);
nand U24216 (N_24216,N_16926,N_16502);
or U24217 (N_24217,N_19467,N_18885);
and U24218 (N_24218,N_15965,N_18685);
nor U24219 (N_24219,N_17219,N_19154);
nand U24220 (N_24220,N_19704,N_19545);
xnor U24221 (N_24221,N_15251,N_19488);
nor U24222 (N_24222,N_17596,N_16181);
or U24223 (N_24223,N_18915,N_16160);
xnor U24224 (N_24224,N_16603,N_19408);
nor U24225 (N_24225,N_18700,N_17129);
nor U24226 (N_24226,N_15110,N_16177);
nor U24227 (N_24227,N_15235,N_15818);
and U24228 (N_24228,N_16379,N_17109);
nand U24229 (N_24229,N_18155,N_19995);
and U24230 (N_24230,N_18327,N_18322);
and U24231 (N_24231,N_15929,N_18807);
nor U24232 (N_24232,N_18818,N_19303);
or U24233 (N_24233,N_17762,N_15731);
and U24234 (N_24234,N_16764,N_15173);
and U24235 (N_24235,N_16041,N_18910);
nand U24236 (N_24236,N_16105,N_16567);
nand U24237 (N_24237,N_18551,N_15389);
nand U24238 (N_24238,N_19926,N_19710);
nor U24239 (N_24239,N_18374,N_19942);
nor U24240 (N_24240,N_16079,N_18569);
nand U24241 (N_24241,N_15484,N_17086);
and U24242 (N_24242,N_18822,N_15300);
nand U24243 (N_24243,N_15267,N_15270);
nand U24244 (N_24244,N_15111,N_19447);
xnor U24245 (N_24245,N_18473,N_18855);
nand U24246 (N_24246,N_16259,N_18909);
nand U24247 (N_24247,N_17307,N_15134);
nand U24248 (N_24248,N_19704,N_19021);
or U24249 (N_24249,N_17535,N_16148);
or U24250 (N_24250,N_16953,N_18728);
nand U24251 (N_24251,N_18592,N_15425);
xnor U24252 (N_24252,N_19272,N_16098);
nand U24253 (N_24253,N_18340,N_17702);
and U24254 (N_24254,N_15490,N_15894);
nor U24255 (N_24255,N_17797,N_16427);
xor U24256 (N_24256,N_19345,N_15996);
nor U24257 (N_24257,N_17417,N_18962);
or U24258 (N_24258,N_19415,N_17512);
xnor U24259 (N_24259,N_16912,N_16779);
xor U24260 (N_24260,N_17571,N_17450);
nor U24261 (N_24261,N_15405,N_17750);
nor U24262 (N_24262,N_16143,N_17832);
and U24263 (N_24263,N_19642,N_18187);
nand U24264 (N_24264,N_19269,N_18942);
nor U24265 (N_24265,N_19686,N_17526);
nand U24266 (N_24266,N_15754,N_16570);
and U24267 (N_24267,N_17145,N_16519);
xnor U24268 (N_24268,N_16361,N_17111);
or U24269 (N_24269,N_18407,N_17482);
xor U24270 (N_24270,N_17261,N_18957);
nand U24271 (N_24271,N_18778,N_19952);
xor U24272 (N_24272,N_17093,N_17149);
nand U24273 (N_24273,N_19394,N_17182);
nand U24274 (N_24274,N_17082,N_18363);
nor U24275 (N_24275,N_15077,N_16630);
xnor U24276 (N_24276,N_15699,N_19504);
or U24277 (N_24277,N_18896,N_17720);
or U24278 (N_24278,N_18912,N_17421);
or U24279 (N_24279,N_17895,N_17481);
and U24280 (N_24280,N_16591,N_15726);
nor U24281 (N_24281,N_17432,N_16929);
nor U24282 (N_24282,N_19582,N_17418);
and U24283 (N_24283,N_19767,N_19409);
or U24284 (N_24284,N_18613,N_16137);
or U24285 (N_24285,N_16103,N_15261);
nor U24286 (N_24286,N_15546,N_17447);
nor U24287 (N_24287,N_17909,N_16427);
nor U24288 (N_24288,N_19793,N_19089);
nand U24289 (N_24289,N_17170,N_15968);
or U24290 (N_24290,N_15074,N_18010);
xnor U24291 (N_24291,N_16820,N_18569);
or U24292 (N_24292,N_15300,N_16153);
nand U24293 (N_24293,N_16417,N_15059);
nand U24294 (N_24294,N_18958,N_19055);
or U24295 (N_24295,N_17484,N_17264);
nand U24296 (N_24296,N_16255,N_16772);
nand U24297 (N_24297,N_17499,N_19691);
nand U24298 (N_24298,N_16074,N_15969);
nand U24299 (N_24299,N_17090,N_18076);
xnor U24300 (N_24300,N_19754,N_16199);
nand U24301 (N_24301,N_15491,N_16537);
nand U24302 (N_24302,N_17567,N_15417);
and U24303 (N_24303,N_17898,N_19328);
and U24304 (N_24304,N_18942,N_15967);
nand U24305 (N_24305,N_19623,N_17572);
and U24306 (N_24306,N_19868,N_18620);
or U24307 (N_24307,N_15435,N_15125);
nor U24308 (N_24308,N_15446,N_16470);
nand U24309 (N_24309,N_17989,N_16618);
and U24310 (N_24310,N_19529,N_15805);
nor U24311 (N_24311,N_19845,N_16402);
or U24312 (N_24312,N_18413,N_17171);
and U24313 (N_24313,N_15574,N_15710);
or U24314 (N_24314,N_19650,N_17380);
nand U24315 (N_24315,N_15577,N_17803);
or U24316 (N_24316,N_16781,N_16411);
xor U24317 (N_24317,N_17134,N_18977);
nand U24318 (N_24318,N_17908,N_17214);
and U24319 (N_24319,N_15418,N_18705);
xor U24320 (N_24320,N_18442,N_19156);
nor U24321 (N_24321,N_17653,N_19965);
or U24322 (N_24322,N_16318,N_18865);
xnor U24323 (N_24323,N_18078,N_16550);
or U24324 (N_24324,N_19235,N_19059);
nor U24325 (N_24325,N_16091,N_18156);
or U24326 (N_24326,N_17697,N_15891);
nor U24327 (N_24327,N_16674,N_19881);
nor U24328 (N_24328,N_16709,N_18653);
and U24329 (N_24329,N_17372,N_17790);
xnor U24330 (N_24330,N_18484,N_19268);
xor U24331 (N_24331,N_17559,N_19044);
xnor U24332 (N_24332,N_17717,N_17947);
xor U24333 (N_24333,N_15424,N_18171);
nor U24334 (N_24334,N_19672,N_17959);
nor U24335 (N_24335,N_19485,N_19843);
or U24336 (N_24336,N_15734,N_18039);
nand U24337 (N_24337,N_15146,N_19249);
or U24338 (N_24338,N_15746,N_19830);
xor U24339 (N_24339,N_18110,N_17176);
nor U24340 (N_24340,N_18032,N_16477);
and U24341 (N_24341,N_18943,N_17957);
xor U24342 (N_24342,N_17842,N_16335);
or U24343 (N_24343,N_15413,N_19786);
and U24344 (N_24344,N_16528,N_17928);
or U24345 (N_24345,N_17409,N_18130);
or U24346 (N_24346,N_18036,N_16660);
xor U24347 (N_24347,N_15746,N_15950);
or U24348 (N_24348,N_15619,N_17455);
nand U24349 (N_24349,N_19712,N_17473);
nor U24350 (N_24350,N_16151,N_18263);
or U24351 (N_24351,N_19684,N_15500);
and U24352 (N_24352,N_19018,N_17308);
xnor U24353 (N_24353,N_15366,N_18257);
xnor U24354 (N_24354,N_16579,N_19859);
or U24355 (N_24355,N_19336,N_15637);
xnor U24356 (N_24356,N_19504,N_18722);
nand U24357 (N_24357,N_15035,N_15579);
and U24358 (N_24358,N_17526,N_15078);
nor U24359 (N_24359,N_19416,N_18270);
and U24360 (N_24360,N_19859,N_17484);
or U24361 (N_24361,N_16749,N_17937);
xor U24362 (N_24362,N_17721,N_19757);
nand U24363 (N_24363,N_15990,N_15801);
or U24364 (N_24364,N_19756,N_17820);
and U24365 (N_24365,N_19643,N_17403);
nor U24366 (N_24366,N_16830,N_15694);
or U24367 (N_24367,N_15639,N_19228);
or U24368 (N_24368,N_18505,N_17691);
nor U24369 (N_24369,N_15517,N_19831);
xnor U24370 (N_24370,N_16986,N_17907);
xnor U24371 (N_24371,N_19074,N_19645);
and U24372 (N_24372,N_15239,N_18741);
or U24373 (N_24373,N_15428,N_19272);
and U24374 (N_24374,N_18643,N_18201);
or U24375 (N_24375,N_19901,N_15832);
and U24376 (N_24376,N_19741,N_15885);
and U24377 (N_24377,N_18296,N_16407);
nand U24378 (N_24378,N_16471,N_16520);
nand U24379 (N_24379,N_17232,N_15113);
nor U24380 (N_24380,N_17444,N_17648);
xor U24381 (N_24381,N_17989,N_16071);
or U24382 (N_24382,N_16472,N_19079);
xor U24383 (N_24383,N_18782,N_17536);
and U24384 (N_24384,N_18690,N_17787);
nor U24385 (N_24385,N_16233,N_16824);
nand U24386 (N_24386,N_15835,N_16205);
or U24387 (N_24387,N_18900,N_19380);
or U24388 (N_24388,N_19071,N_17325);
nor U24389 (N_24389,N_15878,N_19456);
nand U24390 (N_24390,N_19878,N_16637);
and U24391 (N_24391,N_15576,N_15080);
or U24392 (N_24392,N_16600,N_16737);
nor U24393 (N_24393,N_17270,N_18185);
or U24394 (N_24394,N_15979,N_16062);
xor U24395 (N_24395,N_16174,N_17480);
nor U24396 (N_24396,N_15066,N_18740);
and U24397 (N_24397,N_17582,N_16072);
xnor U24398 (N_24398,N_16510,N_17530);
and U24399 (N_24399,N_17205,N_17817);
or U24400 (N_24400,N_16576,N_15999);
and U24401 (N_24401,N_18713,N_17655);
xor U24402 (N_24402,N_17116,N_19765);
nor U24403 (N_24403,N_16707,N_15163);
nand U24404 (N_24404,N_18484,N_19001);
xor U24405 (N_24405,N_16794,N_18630);
xnor U24406 (N_24406,N_16425,N_17687);
and U24407 (N_24407,N_18487,N_15328);
xnor U24408 (N_24408,N_19049,N_16675);
nor U24409 (N_24409,N_17289,N_15113);
nand U24410 (N_24410,N_16974,N_19923);
or U24411 (N_24411,N_19702,N_19978);
xnor U24412 (N_24412,N_19530,N_17182);
and U24413 (N_24413,N_15099,N_19189);
or U24414 (N_24414,N_18946,N_18526);
nand U24415 (N_24415,N_19910,N_15125);
or U24416 (N_24416,N_18455,N_17664);
nand U24417 (N_24417,N_19006,N_16198);
nor U24418 (N_24418,N_16335,N_18415);
or U24419 (N_24419,N_17362,N_15823);
nand U24420 (N_24420,N_17548,N_17278);
xor U24421 (N_24421,N_19112,N_18251);
xor U24422 (N_24422,N_16807,N_17797);
nand U24423 (N_24423,N_17829,N_18594);
nand U24424 (N_24424,N_15796,N_18134);
xnor U24425 (N_24425,N_18174,N_17849);
or U24426 (N_24426,N_17250,N_18684);
xor U24427 (N_24427,N_18721,N_17196);
nor U24428 (N_24428,N_18830,N_17254);
or U24429 (N_24429,N_16197,N_15340);
and U24430 (N_24430,N_15388,N_17569);
or U24431 (N_24431,N_15974,N_16788);
and U24432 (N_24432,N_16223,N_16002);
and U24433 (N_24433,N_17784,N_19387);
nor U24434 (N_24434,N_16585,N_18759);
nand U24435 (N_24435,N_15225,N_18551);
nor U24436 (N_24436,N_16325,N_16856);
or U24437 (N_24437,N_17738,N_15447);
and U24438 (N_24438,N_19776,N_16771);
nand U24439 (N_24439,N_15366,N_18934);
nor U24440 (N_24440,N_16616,N_18266);
and U24441 (N_24441,N_15269,N_19701);
xnor U24442 (N_24442,N_15013,N_19679);
nand U24443 (N_24443,N_15389,N_18420);
nand U24444 (N_24444,N_15798,N_19778);
xnor U24445 (N_24445,N_18978,N_19086);
xor U24446 (N_24446,N_15200,N_18631);
nor U24447 (N_24447,N_16436,N_18683);
nor U24448 (N_24448,N_15351,N_17931);
nand U24449 (N_24449,N_17961,N_17427);
and U24450 (N_24450,N_15168,N_18854);
xnor U24451 (N_24451,N_19768,N_18691);
or U24452 (N_24452,N_19299,N_15342);
and U24453 (N_24453,N_18828,N_19771);
nand U24454 (N_24454,N_19848,N_17743);
nor U24455 (N_24455,N_19866,N_18724);
nand U24456 (N_24456,N_15977,N_17305);
xnor U24457 (N_24457,N_19710,N_16735);
nor U24458 (N_24458,N_15180,N_17491);
nand U24459 (N_24459,N_18557,N_17890);
nand U24460 (N_24460,N_15144,N_15499);
or U24461 (N_24461,N_18503,N_15099);
nor U24462 (N_24462,N_15843,N_19230);
nand U24463 (N_24463,N_19477,N_19409);
xnor U24464 (N_24464,N_18326,N_17147);
xnor U24465 (N_24465,N_15737,N_18597);
nor U24466 (N_24466,N_18213,N_16374);
nand U24467 (N_24467,N_15956,N_15547);
xor U24468 (N_24468,N_16462,N_19119);
or U24469 (N_24469,N_15790,N_16148);
nand U24470 (N_24470,N_18592,N_19145);
or U24471 (N_24471,N_17303,N_18076);
nor U24472 (N_24472,N_15094,N_19338);
nor U24473 (N_24473,N_18360,N_17587);
or U24474 (N_24474,N_19115,N_18541);
nor U24475 (N_24475,N_17560,N_16102);
or U24476 (N_24476,N_16134,N_16055);
and U24477 (N_24477,N_16053,N_15131);
xor U24478 (N_24478,N_18150,N_19421);
nor U24479 (N_24479,N_16524,N_16181);
nor U24480 (N_24480,N_17935,N_19652);
nand U24481 (N_24481,N_18156,N_19504);
nor U24482 (N_24482,N_18308,N_15133);
xor U24483 (N_24483,N_16943,N_15110);
nand U24484 (N_24484,N_18220,N_16716);
nor U24485 (N_24485,N_15744,N_16977);
nand U24486 (N_24486,N_19783,N_18181);
nor U24487 (N_24487,N_18830,N_15062);
and U24488 (N_24488,N_17322,N_16234);
nand U24489 (N_24489,N_18432,N_16530);
nor U24490 (N_24490,N_15160,N_19825);
nand U24491 (N_24491,N_18830,N_17751);
or U24492 (N_24492,N_19984,N_16694);
and U24493 (N_24493,N_19250,N_19166);
nor U24494 (N_24494,N_18610,N_15504);
and U24495 (N_24495,N_18193,N_19422);
and U24496 (N_24496,N_18996,N_17362);
nand U24497 (N_24497,N_19893,N_18083);
and U24498 (N_24498,N_15344,N_18023);
nor U24499 (N_24499,N_19707,N_16709);
and U24500 (N_24500,N_18548,N_16804);
nand U24501 (N_24501,N_15735,N_15807);
xnor U24502 (N_24502,N_17534,N_15995);
nand U24503 (N_24503,N_15851,N_16090);
nor U24504 (N_24504,N_18772,N_17456);
and U24505 (N_24505,N_16110,N_16921);
or U24506 (N_24506,N_16532,N_15006);
xnor U24507 (N_24507,N_16084,N_18410);
or U24508 (N_24508,N_19478,N_17679);
or U24509 (N_24509,N_15910,N_15516);
nand U24510 (N_24510,N_18398,N_16762);
nand U24511 (N_24511,N_15520,N_17458);
and U24512 (N_24512,N_16008,N_15383);
nor U24513 (N_24513,N_19259,N_19494);
nand U24514 (N_24514,N_16380,N_15977);
nand U24515 (N_24515,N_15058,N_18795);
or U24516 (N_24516,N_16523,N_19517);
or U24517 (N_24517,N_17592,N_15120);
and U24518 (N_24518,N_17410,N_18280);
and U24519 (N_24519,N_17566,N_19567);
nor U24520 (N_24520,N_15065,N_18736);
xnor U24521 (N_24521,N_15504,N_15416);
xnor U24522 (N_24522,N_18760,N_18381);
or U24523 (N_24523,N_15425,N_19199);
and U24524 (N_24524,N_18484,N_15052);
nand U24525 (N_24525,N_15472,N_18257);
and U24526 (N_24526,N_16109,N_15541);
xnor U24527 (N_24527,N_18001,N_19540);
or U24528 (N_24528,N_17242,N_15577);
nor U24529 (N_24529,N_16381,N_16713);
nand U24530 (N_24530,N_18339,N_16454);
nand U24531 (N_24531,N_15215,N_18772);
and U24532 (N_24532,N_18940,N_17970);
or U24533 (N_24533,N_19079,N_16632);
nor U24534 (N_24534,N_19396,N_19504);
nand U24535 (N_24535,N_19616,N_17579);
and U24536 (N_24536,N_17361,N_15267);
nor U24537 (N_24537,N_18610,N_17756);
xor U24538 (N_24538,N_17266,N_17965);
nor U24539 (N_24539,N_19621,N_18871);
or U24540 (N_24540,N_19301,N_18133);
and U24541 (N_24541,N_19300,N_18569);
xor U24542 (N_24542,N_17318,N_16343);
nor U24543 (N_24543,N_17747,N_16070);
nor U24544 (N_24544,N_16987,N_19603);
and U24545 (N_24545,N_18408,N_19925);
xnor U24546 (N_24546,N_16430,N_19678);
xnor U24547 (N_24547,N_19989,N_19348);
xnor U24548 (N_24548,N_17836,N_17957);
or U24549 (N_24549,N_17036,N_16184);
and U24550 (N_24550,N_19579,N_17984);
nand U24551 (N_24551,N_17823,N_19677);
or U24552 (N_24552,N_16766,N_17541);
or U24553 (N_24553,N_15051,N_18661);
xor U24554 (N_24554,N_18795,N_16164);
nor U24555 (N_24555,N_18322,N_17046);
or U24556 (N_24556,N_16930,N_18288);
nand U24557 (N_24557,N_15545,N_15113);
nand U24558 (N_24558,N_17797,N_17596);
and U24559 (N_24559,N_16883,N_17992);
and U24560 (N_24560,N_17837,N_18234);
or U24561 (N_24561,N_16414,N_18228);
nor U24562 (N_24562,N_15005,N_17204);
nand U24563 (N_24563,N_19534,N_19641);
nor U24564 (N_24564,N_18852,N_18062);
xor U24565 (N_24565,N_17712,N_19904);
nand U24566 (N_24566,N_19169,N_19756);
xnor U24567 (N_24567,N_16105,N_15339);
or U24568 (N_24568,N_15367,N_16057);
and U24569 (N_24569,N_19273,N_19841);
nor U24570 (N_24570,N_18288,N_18784);
and U24571 (N_24571,N_19542,N_15930);
and U24572 (N_24572,N_17854,N_18017);
nor U24573 (N_24573,N_19770,N_17203);
nor U24574 (N_24574,N_18947,N_17422);
nand U24575 (N_24575,N_19082,N_17140);
and U24576 (N_24576,N_15928,N_16067);
or U24577 (N_24577,N_16004,N_17896);
or U24578 (N_24578,N_15954,N_17991);
xnor U24579 (N_24579,N_16245,N_19832);
nor U24580 (N_24580,N_15241,N_18727);
xnor U24581 (N_24581,N_15403,N_19829);
xnor U24582 (N_24582,N_19022,N_19289);
and U24583 (N_24583,N_19817,N_18432);
xnor U24584 (N_24584,N_15267,N_18909);
and U24585 (N_24585,N_18525,N_19204);
nand U24586 (N_24586,N_16807,N_19239);
nand U24587 (N_24587,N_17592,N_16534);
xor U24588 (N_24588,N_19109,N_18593);
nand U24589 (N_24589,N_18863,N_15526);
nand U24590 (N_24590,N_19578,N_16518);
nand U24591 (N_24591,N_19288,N_15113);
nor U24592 (N_24592,N_16479,N_19089);
nand U24593 (N_24593,N_15667,N_19280);
or U24594 (N_24594,N_17646,N_17320);
or U24595 (N_24595,N_15082,N_15059);
nor U24596 (N_24596,N_17022,N_15081);
xnor U24597 (N_24597,N_17889,N_15401);
xnor U24598 (N_24598,N_15853,N_17570);
or U24599 (N_24599,N_19343,N_16145);
and U24600 (N_24600,N_18205,N_16103);
or U24601 (N_24601,N_18577,N_18048);
and U24602 (N_24602,N_19858,N_15614);
nor U24603 (N_24603,N_16940,N_19815);
nor U24604 (N_24604,N_19233,N_17164);
nand U24605 (N_24605,N_18896,N_19248);
xnor U24606 (N_24606,N_17192,N_17076);
nand U24607 (N_24607,N_16321,N_18963);
nor U24608 (N_24608,N_19494,N_19107);
and U24609 (N_24609,N_19169,N_17361);
and U24610 (N_24610,N_19210,N_17687);
nand U24611 (N_24611,N_15255,N_15609);
xor U24612 (N_24612,N_18683,N_18056);
nor U24613 (N_24613,N_19212,N_19649);
or U24614 (N_24614,N_18305,N_18991);
xor U24615 (N_24615,N_16540,N_18716);
and U24616 (N_24616,N_16658,N_18132);
nor U24617 (N_24617,N_19388,N_17486);
nor U24618 (N_24618,N_19351,N_18719);
xor U24619 (N_24619,N_19020,N_15284);
nand U24620 (N_24620,N_16213,N_15824);
or U24621 (N_24621,N_19506,N_18946);
nand U24622 (N_24622,N_16048,N_18646);
and U24623 (N_24623,N_16057,N_19463);
and U24624 (N_24624,N_17803,N_15206);
nor U24625 (N_24625,N_18827,N_16780);
nor U24626 (N_24626,N_18099,N_16084);
xor U24627 (N_24627,N_15209,N_16638);
or U24628 (N_24628,N_18125,N_17452);
nand U24629 (N_24629,N_17018,N_16692);
and U24630 (N_24630,N_18142,N_17975);
or U24631 (N_24631,N_15185,N_16137);
nand U24632 (N_24632,N_17302,N_18320);
and U24633 (N_24633,N_19505,N_19295);
xnor U24634 (N_24634,N_18111,N_18506);
xor U24635 (N_24635,N_15644,N_16522);
nor U24636 (N_24636,N_18641,N_16228);
and U24637 (N_24637,N_19147,N_15466);
or U24638 (N_24638,N_18265,N_18790);
xnor U24639 (N_24639,N_19058,N_15073);
nor U24640 (N_24640,N_16681,N_16970);
xor U24641 (N_24641,N_17654,N_17453);
nand U24642 (N_24642,N_16038,N_19919);
nor U24643 (N_24643,N_16269,N_15022);
nand U24644 (N_24644,N_19431,N_17688);
nor U24645 (N_24645,N_18795,N_17384);
or U24646 (N_24646,N_16874,N_17696);
or U24647 (N_24647,N_18509,N_19352);
nor U24648 (N_24648,N_17561,N_18385);
nand U24649 (N_24649,N_15101,N_19306);
nand U24650 (N_24650,N_17865,N_18169);
nand U24651 (N_24651,N_17231,N_18075);
and U24652 (N_24652,N_16895,N_15013);
xnor U24653 (N_24653,N_16509,N_19709);
xnor U24654 (N_24654,N_19532,N_17617);
nor U24655 (N_24655,N_19019,N_18810);
xor U24656 (N_24656,N_17905,N_19244);
nand U24657 (N_24657,N_18932,N_15369);
xor U24658 (N_24658,N_18092,N_19488);
nor U24659 (N_24659,N_16999,N_17661);
xnor U24660 (N_24660,N_19350,N_18783);
nand U24661 (N_24661,N_15267,N_19022);
nor U24662 (N_24662,N_18047,N_17227);
and U24663 (N_24663,N_19116,N_18403);
nor U24664 (N_24664,N_17029,N_15240);
nor U24665 (N_24665,N_15474,N_17703);
nor U24666 (N_24666,N_18255,N_19209);
nand U24667 (N_24667,N_15176,N_15703);
or U24668 (N_24668,N_17913,N_17301);
nand U24669 (N_24669,N_15254,N_17272);
nor U24670 (N_24670,N_15120,N_15918);
or U24671 (N_24671,N_17686,N_16930);
nor U24672 (N_24672,N_19293,N_17555);
or U24673 (N_24673,N_15301,N_19172);
or U24674 (N_24674,N_18867,N_16648);
xor U24675 (N_24675,N_19740,N_18406);
or U24676 (N_24676,N_16076,N_15388);
xnor U24677 (N_24677,N_16746,N_16911);
or U24678 (N_24678,N_17222,N_19674);
nand U24679 (N_24679,N_19802,N_18560);
or U24680 (N_24680,N_19618,N_16495);
and U24681 (N_24681,N_19083,N_18117);
nand U24682 (N_24682,N_15548,N_17535);
and U24683 (N_24683,N_18342,N_19084);
nand U24684 (N_24684,N_18989,N_17612);
xor U24685 (N_24685,N_18852,N_17022);
and U24686 (N_24686,N_15068,N_19312);
or U24687 (N_24687,N_16185,N_16031);
xnor U24688 (N_24688,N_18072,N_16628);
or U24689 (N_24689,N_17499,N_15002);
xor U24690 (N_24690,N_18538,N_19750);
nand U24691 (N_24691,N_15376,N_17632);
and U24692 (N_24692,N_16302,N_15630);
or U24693 (N_24693,N_16030,N_17094);
nor U24694 (N_24694,N_17647,N_15794);
and U24695 (N_24695,N_19148,N_18478);
nor U24696 (N_24696,N_17544,N_19430);
xor U24697 (N_24697,N_19876,N_17784);
nand U24698 (N_24698,N_15495,N_18024);
and U24699 (N_24699,N_15628,N_19958);
nand U24700 (N_24700,N_16125,N_18022);
nand U24701 (N_24701,N_15328,N_15341);
or U24702 (N_24702,N_16169,N_18542);
and U24703 (N_24703,N_16616,N_15045);
xor U24704 (N_24704,N_18235,N_18327);
or U24705 (N_24705,N_15992,N_16688);
and U24706 (N_24706,N_18817,N_17289);
xnor U24707 (N_24707,N_18454,N_17648);
xor U24708 (N_24708,N_16877,N_17850);
nand U24709 (N_24709,N_15153,N_16471);
or U24710 (N_24710,N_19630,N_17395);
or U24711 (N_24711,N_18062,N_16499);
nor U24712 (N_24712,N_16582,N_16004);
nor U24713 (N_24713,N_19642,N_15290);
and U24714 (N_24714,N_16706,N_15709);
and U24715 (N_24715,N_17552,N_16129);
nand U24716 (N_24716,N_18629,N_18621);
nor U24717 (N_24717,N_15494,N_15423);
or U24718 (N_24718,N_19713,N_19795);
xnor U24719 (N_24719,N_18745,N_16948);
nand U24720 (N_24720,N_18124,N_16024);
nor U24721 (N_24721,N_17777,N_16782);
nor U24722 (N_24722,N_19779,N_19352);
and U24723 (N_24723,N_17397,N_18915);
nor U24724 (N_24724,N_16087,N_15607);
xnor U24725 (N_24725,N_15073,N_17982);
xnor U24726 (N_24726,N_15461,N_16700);
or U24727 (N_24727,N_16429,N_19490);
or U24728 (N_24728,N_15146,N_15439);
or U24729 (N_24729,N_16591,N_19175);
or U24730 (N_24730,N_15253,N_16486);
or U24731 (N_24731,N_16021,N_18411);
nor U24732 (N_24732,N_18090,N_17220);
nand U24733 (N_24733,N_19900,N_16899);
nor U24734 (N_24734,N_15020,N_17075);
nand U24735 (N_24735,N_19352,N_16234);
or U24736 (N_24736,N_16430,N_17449);
or U24737 (N_24737,N_17389,N_16539);
xor U24738 (N_24738,N_19195,N_17382);
nand U24739 (N_24739,N_16622,N_16386);
and U24740 (N_24740,N_19716,N_18570);
or U24741 (N_24741,N_18154,N_16468);
and U24742 (N_24742,N_18346,N_17150);
nor U24743 (N_24743,N_19138,N_17254);
and U24744 (N_24744,N_16569,N_15695);
xor U24745 (N_24745,N_15247,N_19711);
nor U24746 (N_24746,N_19724,N_19189);
nor U24747 (N_24747,N_19934,N_16514);
and U24748 (N_24748,N_16621,N_17518);
or U24749 (N_24749,N_16905,N_18500);
nand U24750 (N_24750,N_16788,N_18931);
nand U24751 (N_24751,N_16108,N_16106);
or U24752 (N_24752,N_15881,N_19497);
xnor U24753 (N_24753,N_17581,N_17504);
and U24754 (N_24754,N_15314,N_16961);
nand U24755 (N_24755,N_16236,N_17319);
and U24756 (N_24756,N_15456,N_17373);
nor U24757 (N_24757,N_18353,N_19773);
nor U24758 (N_24758,N_16565,N_15402);
nor U24759 (N_24759,N_16923,N_19775);
nor U24760 (N_24760,N_19921,N_18346);
xnor U24761 (N_24761,N_18057,N_16240);
nand U24762 (N_24762,N_19286,N_19932);
nor U24763 (N_24763,N_18008,N_16066);
and U24764 (N_24764,N_17286,N_17287);
xor U24765 (N_24765,N_17686,N_16347);
nor U24766 (N_24766,N_17158,N_15989);
xnor U24767 (N_24767,N_16540,N_19951);
nand U24768 (N_24768,N_17269,N_19459);
and U24769 (N_24769,N_15731,N_17213);
nor U24770 (N_24770,N_17857,N_16738);
nand U24771 (N_24771,N_18726,N_19017);
or U24772 (N_24772,N_15790,N_17695);
xor U24773 (N_24773,N_17638,N_19919);
and U24774 (N_24774,N_16245,N_15751);
nand U24775 (N_24775,N_19064,N_16102);
or U24776 (N_24776,N_17170,N_19877);
nor U24777 (N_24777,N_16960,N_18306);
and U24778 (N_24778,N_19762,N_17687);
xnor U24779 (N_24779,N_19226,N_15490);
or U24780 (N_24780,N_18225,N_17099);
xor U24781 (N_24781,N_16204,N_18202);
nand U24782 (N_24782,N_19430,N_18952);
xnor U24783 (N_24783,N_18313,N_18334);
and U24784 (N_24784,N_15525,N_18448);
and U24785 (N_24785,N_18905,N_18520);
xor U24786 (N_24786,N_19559,N_17470);
or U24787 (N_24787,N_15358,N_19112);
nand U24788 (N_24788,N_17191,N_16139);
or U24789 (N_24789,N_18787,N_17040);
or U24790 (N_24790,N_18116,N_15332);
nand U24791 (N_24791,N_15399,N_16045);
nor U24792 (N_24792,N_15217,N_18973);
nand U24793 (N_24793,N_16198,N_19821);
and U24794 (N_24794,N_16902,N_16932);
or U24795 (N_24795,N_19567,N_16121);
nor U24796 (N_24796,N_15596,N_16559);
xor U24797 (N_24797,N_18903,N_15580);
nor U24798 (N_24798,N_19149,N_17144);
or U24799 (N_24799,N_15926,N_16158);
nand U24800 (N_24800,N_16505,N_17032);
xor U24801 (N_24801,N_15292,N_19046);
nand U24802 (N_24802,N_15943,N_17469);
or U24803 (N_24803,N_16563,N_17388);
nand U24804 (N_24804,N_17291,N_19202);
nor U24805 (N_24805,N_17961,N_18336);
or U24806 (N_24806,N_17520,N_18678);
xor U24807 (N_24807,N_17133,N_18416);
nor U24808 (N_24808,N_16695,N_18606);
or U24809 (N_24809,N_17607,N_19520);
nor U24810 (N_24810,N_15840,N_18488);
nand U24811 (N_24811,N_15983,N_17061);
xnor U24812 (N_24812,N_18966,N_17956);
nor U24813 (N_24813,N_19346,N_17245);
nor U24814 (N_24814,N_17063,N_15320);
and U24815 (N_24815,N_19504,N_15348);
and U24816 (N_24816,N_19575,N_19083);
and U24817 (N_24817,N_16459,N_16161);
or U24818 (N_24818,N_15211,N_19057);
or U24819 (N_24819,N_16024,N_17596);
nand U24820 (N_24820,N_16197,N_19956);
or U24821 (N_24821,N_19770,N_17376);
nor U24822 (N_24822,N_17656,N_15150);
nor U24823 (N_24823,N_18554,N_17172);
xnor U24824 (N_24824,N_16893,N_19781);
or U24825 (N_24825,N_16241,N_18179);
nor U24826 (N_24826,N_19432,N_15365);
and U24827 (N_24827,N_19919,N_15767);
and U24828 (N_24828,N_19568,N_16326);
nor U24829 (N_24829,N_18861,N_19974);
nor U24830 (N_24830,N_19855,N_19423);
xor U24831 (N_24831,N_18628,N_15289);
or U24832 (N_24832,N_19503,N_19779);
or U24833 (N_24833,N_18954,N_18910);
nand U24834 (N_24834,N_19170,N_17925);
xor U24835 (N_24835,N_17844,N_15788);
nand U24836 (N_24836,N_18217,N_17160);
and U24837 (N_24837,N_19353,N_18140);
and U24838 (N_24838,N_18107,N_16351);
or U24839 (N_24839,N_18712,N_16415);
nand U24840 (N_24840,N_18355,N_18929);
xnor U24841 (N_24841,N_16203,N_16881);
and U24842 (N_24842,N_18247,N_19397);
nor U24843 (N_24843,N_19359,N_18092);
xnor U24844 (N_24844,N_17918,N_19455);
or U24845 (N_24845,N_19989,N_15036);
xnor U24846 (N_24846,N_17282,N_16523);
nor U24847 (N_24847,N_16143,N_15914);
or U24848 (N_24848,N_19609,N_16054);
nor U24849 (N_24849,N_19274,N_19830);
or U24850 (N_24850,N_15939,N_16583);
and U24851 (N_24851,N_16597,N_16513);
xor U24852 (N_24852,N_18905,N_16931);
xnor U24853 (N_24853,N_19219,N_18794);
xnor U24854 (N_24854,N_18802,N_16605);
nor U24855 (N_24855,N_16799,N_19426);
or U24856 (N_24856,N_17144,N_18207);
xor U24857 (N_24857,N_18676,N_18585);
xor U24858 (N_24858,N_17970,N_16714);
or U24859 (N_24859,N_17105,N_18917);
xor U24860 (N_24860,N_19285,N_19760);
xor U24861 (N_24861,N_19719,N_15515);
nor U24862 (N_24862,N_16785,N_17551);
or U24863 (N_24863,N_15970,N_19518);
nand U24864 (N_24864,N_17306,N_15110);
and U24865 (N_24865,N_17579,N_18095);
or U24866 (N_24866,N_16793,N_17615);
nor U24867 (N_24867,N_18164,N_15492);
xor U24868 (N_24868,N_16685,N_17438);
xnor U24869 (N_24869,N_16841,N_15203);
nand U24870 (N_24870,N_16718,N_16543);
or U24871 (N_24871,N_15666,N_16760);
nand U24872 (N_24872,N_16161,N_19597);
or U24873 (N_24873,N_16371,N_19716);
xnor U24874 (N_24874,N_18045,N_17467);
xnor U24875 (N_24875,N_17183,N_17791);
or U24876 (N_24876,N_15034,N_15615);
and U24877 (N_24877,N_17406,N_19847);
or U24878 (N_24878,N_19880,N_15979);
xnor U24879 (N_24879,N_19211,N_15490);
nand U24880 (N_24880,N_16913,N_15897);
nor U24881 (N_24881,N_17525,N_16568);
or U24882 (N_24882,N_19597,N_16968);
or U24883 (N_24883,N_17211,N_17689);
or U24884 (N_24884,N_18650,N_19607);
and U24885 (N_24885,N_17977,N_16127);
xnor U24886 (N_24886,N_15858,N_15569);
or U24887 (N_24887,N_16072,N_18598);
xor U24888 (N_24888,N_17835,N_15904);
xnor U24889 (N_24889,N_18865,N_15982);
and U24890 (N_24890,N_16272,N_16461);
and U24891 (N_24891,N_18138,N_18113);
xnor U24892 (N_24892,N_19730,N_17781);
or U24893 (N_24893,N_15692,N_19461);
or U24894 (N_24894,N_16207,N_16468);
nand U24895 (N_24895,N_18436,N_15377);
and U24896 (N_24896,N_19855,N_19406);
nor U24897 (N_24897,N_16265,N_16576);
nor U24898 (N_24898,N_15684,N_18531);
nor U24899 (N_24899,N_16995,N_15507);
nand U24900 (N_24900,N_18143,N_16271);
xnor U24901 (N_24901,N_16669,N_18245);
xnor U24902 (N_24902,N_17987,N_16894);
nand U24903 (N_24903,N_15270,N_19023);
xor U24904 (N_24904,N_18112,N_15358);
nand U24905 (N_24905,N_19121,N_17784);
and U24906 (N_24906,N_17207,N_19246);
nor U24907 (N_24907,N_19638,N_15879);
nand U24908 (N_24908,N_18024,N_15270);
nand U24909 (N_24909,N_15903,N_16452);
xor U24910 (N_24910,N_16922,N_19365);
nand U24911 (N_24911,N_18411,N_17345);
xor U24912 (N_24912,N_16399,N_15437);
nor U24913 (N_24913,N_18678,N_16758);
or U24914 (N_24914,N_17247,N_17560);
nor U24915 (N_24915,N_18674,N_15388);
xnor U24916 (N_24916,N_17917,N_16975);
and U24917 (N_24917,N_15242,N_15814);
nand U24918 (N_24918,N_15755,N_18302);
xor U24919 (N_24919,N_17278,N_16903);
nand U24920 (N_24920,N_17379,N_15358);
and U24921 (N_24921,N_19936,N_18746);
xor U24922 (N_24922,N_15486,N_15137);
or U24923 (N_24923,N_19741,N_19148);
nand U24924 (N_24924,N_17870,N_16270);
and U24925 (N_24925,N_16147,N_15579);
or U24926 (N_24926,N_18750,N_18018);
and U24927 (N_24927,N_17192,N_18745);
nor U24928 (N_24928,N_16037,N_17013);
nor U24929 (N_24929,N_18304,N_19394);
nor U24930 (N_24930,N_17774,N_16053);
or U24931 (N_24931,N_16025,N_16646);
nor U24932 (N_24932,N_17454,N_17890);
or U24933 (N_24933,N_16924,N_19364);
xor U24934 (N_24934,N_19676,N_19431);
xnor U24935 (N_24935,N_18112,N_18239);
and U24936 (N_24936,N_18876,N_15588);
and U24937 (N_24937,N_15141,N_15031);
xor U24938 (N_24938,N_18306,N_16868);
or U24939 (N_24939,N_17922,N_19933);
and U24940 (N_24940,N_16048,N_16227);
nor U24941 (N_24941,N_18809,N_17357);
nor U24942 (N_24942,N_15320,N_19773);
and U24943 (N_24943,N_19167,N_16516);
xnor U24944 (N_24944,N_15200,N_16889);
and U24945 (N_24945,N_18822,N_15129);
xnor U24946 (N_24946,N_15187,N_17286);
nand U24947 (N_24947,N_15907,N_17257);
nor U24948 (N_24948,N_16608,N_18905);
or U24949 (N_24949,N_17491,N_15407);
nor U24950 (N_24950,N_16565,N_19290);
nand U24951 (N_24951,N_16219,N_15998);
xor U24952 (N_24952,N_19141,N_15508);
nand U24953 (N_24953,N_18716,N_19023);
or U24954 (N_24954,N_19198,N_19841);
nor U24955 (N_24955,N_16240,N_17884);
xor U24956 (N_24956,N_15656,N_16924);
nor U24957 (N_24957,N_17340,N_15318);
or U24958 (N_24958,N_17544,N_17017);
and U24959 (N_24959,N_19130,N_17506);
nor U24960 (N_24960,N_15254,N_15070);
and U24961 (N_24961,N_17371,N_18217);
or U24962 (N_24962,N_18937,N_18594);
and U24963 (N_24963,N_15348,N_17247);
xnor U24964 (N_24964,N_16128,N_19387);
nand U24965 (N_24965,N_15872,N_16771);
xnor U24966 (N_24966,N_15977,N_18778);
xor U24967 (N_24967,N_16602,N_15114);
xor U24968 (N_24968,N_19314,N_16566);
or U24969 (N_24969,N_15082,N_16903);
or U24970 (N_24970,N_17106,N_15598);
xnor U24971 (N_24971,N_17463,N_16782);
nand U24972 (N_24972,N_16009,N_18978);
nand U24973 (N_24973,N_19354,N_17085);
xnor U24974 (N_24974,N_16680,N_19409);
nand U24975 (N_24975,N_17187,N_17630);
and U24976 (N_24976,N_17121,N_19820);
xor U24977 (N_24977,N_15472,N_16470);
and U24978 (N_24978,N_17385,N_16735);
nor U24979 (N_24979,N_16231,N_16546);
and U24980 (N_24980,N_15410,N_16557);
and U24981 (N_24981,N_17712,N_15329);
xor U24982 (N_24982,N_16115,N_19969);
nor U24983 (N_24983,N_16210,N_17294);
nor U24984 (N_24984,N_18911,N_16862);
nand U24985 (N_24985,N_17532,N_19458);
or U24986 (N_24986,N_19899,N_19460);
xor U24987 (N_24987,N_15565,N_19072);
and U24988 (N_24988,N_19739,N_18210);
or U24989 (N_24989,N_17085,N_18158);
nor U24990 (N_24990,N_18372,N_17269);
or U24991 (N_24991,N_19398,N_19724);
and U24992 (N_24992,N_17387,N_16938);
nand U24993 (N_24993,N_19203,N_17196);
and U24994 (N_24994,N_15566,N_16058);
nor U24995 (N_24995,N_15917,N_19777);
or U24996 (N_24996,N_19574,N_17773);
xnor U24997 (N_24997,N_19789,N_17386);
xnor U24998 (N_24998,N_17063,N_15214);
or U24999 (N_24999,N_18362,N_15092);
and U25000 (N_25000,N_24128,N_21354);
xor U25001 (N_25001,N_20128,N_22646);
or U25002 (N_25002,N_21676,N_22173);
xor U25003 (N_25003,N_23530,N_23021);
nand U25004 (N_25004,N_22780,N_23627);
nand U25005 (N_25005,N_20309,N_22264);
and U25006 (N_25006,N_21132,N_22903);
nand U25007 (N_25007,N_22016,N_20894);
nor U25008 (N_25008,N_24400,N_20419);
and U25009 (N_25009,N_20876,N_22927);
nand U25010 (N_25010,N_22214,N_21342);
xor U25011 (N_25011,N_21957,N_21367);
and U25012 (N_25012,N_21781,N_21417);
and U25013 (N_25013,N_23697,N_21815);
nand U25014 (N_25014,N_24253,N_22490);
or U25015 (N_25015,N_21476,N_22141);
and U25016 (N_25016,N_22955,N_22128);
nor U25017 (N_25017,N_24319,N_22569);
nor U25018 (N_25018,N_23362,N_23531);
and U25019 (N_25019,N_24290,N_24043);
xor U25020 (N_25020,N_22262,N_24893);
nor U25021 (N_25021,N_24864,N_22279);
nor U25022 (N_25022,N_22288,N_20688);
nor U25023 (N_25023,N_22861,N_20553);
or U25024 (N_25024,N_24873,N_21489);
or U25025 (N_25025,N_23161,N_21110);
xnor U25026 (N_25026,N_24740,N_21929);
or U25027 (N_25027,N_22649,N_24477);
or U25028 (N_25028,N_20961,N_20262);
or U25029 (N_25029,N_21604,N_21718);
nor U25030 (N_25030,N_24183,N_23398);
nor U25031 (N_25031,N_24769,N_21337);
or U25032 (N_25032,N_22337,N_24537);
xor U25033 (N_25033,N_23248,N_20918);
and U25034 (N_25034,N_22851,N_21142);
nor U25035 (N_25035,N_23411,N_21714);
or U25036 (N_25036,N_22893,N_20330);
nor U25037 (N_25037,N_22554,N_23813);
and U25038 (N_25038,N_21124,N_23453);
nand U25039 (N_25039,N_23311,N_24854);
nor U25040 (N_25040,N_20805,N_22584);
or U25041 (N_25041,N_24387,N_22838);
or U25042 (N_25042,N_23785,N_23635);
xnor U25043 (N_25043,N_20463,N_22402);
xnor U25044 (N_25044,N_22842,N_21953);
xnor U25045 (N_25045,N_20239,N_21620);
and U25046 (N_25046,N_20441,N_24193);
and U25047 (N_25047,N_23672,N_20332);
nand U25048 (N_25048,N_24841,N_24073);
and U25049 (N_25049,N_22041,N_21192);
xnor U25050 (N_25050,N_24294,N_23526);
or U25051 (N_25051,N_20049,N_21126);
nor U25052 (N_25052,N_20323,N_23938);
and U25053 (N_25053,N_23669,N_24037);
xor U25054 (N_25054,N_21669,N_22166);
xor U25055 (N_25055,N_21698,N_24094);
xnor U25056 (N_25056,N_22715,N_24713);
and U25057 (N_25057,N_21673,N_22561);
or U25058 (N_25058,N_24863,N_22997);
nand U25059 (N_25059,N_20452,N_23005);
xnor U25060 (N_25060,N_21278,N_21801);
nand U25061 (N_25061,N_23843,N_21593);
and U25062 (N_25062,N_20637,N_21234);
nor U25063 (N_25063,N_20191,N_21980);
or U25064 (N_25064,N_24258,N_20968);
nand U25065 (N_25065,N_22527,N_23443);
nor U25066 (N_25066,N_20222,N_23979);
nor U25067 (N_25067,N_20376,N_23050);
xor U25068 (N_25068,N_20734,N_23111);
nand U25069 (N_25069,N_20901,N_23514);
nor U25070 (N_25070,N_22832,N_20792);
and U25071 (N_25071,N_24492,N_24778);
nand U25072 (N_25072,N_22974,N_20075);
nand U25073 (N_25073,N_22667,N_23873);
nor U25074 (N_25074,N_20118,N_21903);
xnor U25075 (N_25075,N_20598,N_23297);
or U25076 (N_25076,N_22548,N_21158);
and U25077 (N_25077,N_24923,N_21370);
nand U25078 (N_25078,N_24126,N_24816);
xor U25079 (N_25079,N_22776,N_22465);
nand U25080 (N_25080,N_24001,N_20400);
nand U25081 (N_25081,N_21761,N_21931);
xor U25082 (N_25082,N_23011,N_21486);
and U25083 (N_25083,N_24842,N_21825);
nand U25084 (N_25084,N_24158,N_21228);
and U25085 (N_25085,N_21360,N_22314);
and U25086 (N_25086,N_21112,N_21134);
nand U25087 (N_25087,N_21910,N_23388);
nand U25088 (N_25088,N_23188,N_21413);
nand U25089 (N_25089,N_24718,N_21275);
xor U25090 (N_25090,N_24962,N_23437);
and U25091 (N_25091,N_21883,N_22525);
nand U25092 (N_25092,N_22790,N_24056);
xor U25093 (N_25093,N_22217,N_22785);
or U25094 (N_25094,N_24658,N_22825);
or U25095 (N_25095,N_21920,N_22393);
nor U25096 (N_25096,N_23772,N_22310);
xnor U25097 (N_25097,N_21616,N_22845);
xnor U25098 (N_25098,N_21197,N_20728);
or U25099 (N_25099,N_24327,N_20035);
nor U25100 (N_25100,N_24997,N_24661);
xnor U25101 (N_25101,N_20385,N_24730);
nand U25102 (N_25102,N_22140,N_22232);
nand U25103 (N_25103,N_24760,N_21173);
nor U25104 (N_25104,N_24283,N_22432);
and U25105 (N_25105,N_20321,N_20011);
nand U25106 (N_25106,N_24803,N_24737);
xor U25107 (N_25107,N_21170,N_22835);
nand U25108 (N_25108,N_20313,N_20166);
nor U25109 (N_25109,N_21996,N_23625);
xor U25110 (N_25110,N_24699,N_23808);
and U25111 (N_25111,N_24144,N_20758);
or U25112 (N_25112,N_23083,N_20819);
and U25113 (N_25113,N_20856,N_21252);
or U25114 (N_25114,N_20572,N_24942);
and U25115 (N_25115,N_24596,N_23107);
nand U25116 (N_25116,N_22730,N_21947);
and U25117 (N_25117,N_24714,N_23752);
or U25118 (N_25118,N_24727,N_20829);
nor U25119 (N_25119,N_21856,N_23704);
nand U25120 (N_25120,N_21217,N_22874);
or U25121 (N_25121,N_20018,N_21611);
or U25122 (N_25122,N_20426,N_21432);
nand U25123 (N_25123,N_22856,N_20037);
and U25124 (N_25124,N_21597,N_23053);
or U25125 (N_25125,N_24885,N_21219);
or U25126 (N_25126,N_24301,N_21240);
nor U25127 (N_25127,N_21594,N_24905);
nor U25128 (N_25128,N_20512,N_20378);
nor U25129 (N_25129,N_22272,N_23482);
nor U25130 (N_25130,N_23686,N_24871);
and U25131 (N_25131,N_21932,N_21582);
or U25132 (N_25132,N_24826,N_21079);
and U25133 (N_25133,N_24366,N_21827);
or U25134 (N_25134,N_23851,N_23145);
or U25135 (N_25135,N_22341,N_20840);
nand U25136 (N_25136,N_21227,N_24916);
or U25137 (N_25137,N_23156,N_22003);
or U25138 (N_25138,N_22238,N_21960);
xnor U25139 (N_25139,N_24310,N_24855);
nor U25140 (N_25140,N_20556,N_22481);
xnor U25141 (N_25141,N_22726,N_21470);
nand U25142 (N_25142,N_21341,N_20971);
nand U25143 (N_25143,N_22579,N_22309);
or U25144 (N_25144,N_21114,N_22532);
nand U25145 (N_25145,N_22333,N_24894);
xnor U25146 (N_25146,N_24593,N_21685);
xor U25147 (N_25147,N_20520,N_20051);
nor U25148 (N_25148,N_21571,N_24805);
and U25149 (N_25149,N_21458,N_20267);
nor U25150 (N_25150,N_20163,N_23010);
xnor U25151 (N_25151,N_21231,N_24521);
or U25152 (N_25152,N_22981,N_22088);
xnor U25153 (N_25153,N_23324,N_20745);
or U25154 (N_25154,N_21697,N_20358);
nand U25155 (N_25155,N_23250,N_23995);
xor U25156 (N_25156,N_22446,N_24662);
nand U25157 (N_25157,N_21330,N_23992);
nor U25158 (N_25158,N_24512,N_23164);
nand U25159 (N_25159,N_22713,N_22261);
nand U25160 (N_25160,N_23774,N_22191);
nand U25161 (N_25161,N_24720,N_24022);
or U25162 (N_25162,N_23573,N_23764);
xor U25163 (N_25163,N_24218,N_23160);
xnor U25164 (N_25164,N_24407,N_20743);
or U25165 (N_25165,N_24861,N_21006);
or U25166 (N_25166,N_21215,N_22320);
or U25167 (N_25167,N_21291,N_22717);
or U25168 (N_25168,N_21959,N_21422);
nand U25169 (N_25169,N_24039,N_23396);
or U25170 (N_25170,N_22581,N_23999);
xor U25171 (N_25171,N_23756,N_22537);
nand U25172 (N_25172,N_21648,N_21999);
nand U25173 (N_25173,N_23750,N_24638);
xnor U25174 (N_25174,N_23049,N_20720);
and U25175 (N_25175,N_20697,N_22451);
or U25176 (N_25176,N_21468,N_21975);
nor U25177 (N_25177,N_24766,N_21970);
and U25178 (N_25178,N_23492,N_21510);
or U25179 (N_25179,N_24583,N_24089);
xnor U25180 (N_25180,N_20260,N_20081);
nor U25181 (N_25181,N_21816,N_22152);
nor U25182 (N_25182,N_24426,N_22043);
nand U25183 (N_25183,N_24656,N_23186);
or U25184 (N_25184,N_22211,N_22904);
or U25185 (N_25185,N_23494,N_20089);
xor U25186 (N_25186,N_21819,N_22163);
or U25187 (N_25187,N_23912,N_22850);
or U25188 (N_25188,N_23063,N_22652);
and U25189 (N_25189,N_24839,N_21366);
nor U25190 (N_25190,N_21490,N_22752);
or U25191 (N_25191,N_24579,N_22468);
nand U25192 (N_25192,N_22226,N_20458);
xnor U25193 (N_25193,N_21770,N_23178);
or U25194 (N_25194,N_22268,N_20233);
and U25195 (N_25195,N_22102,N_24024);
xnor U25196 (N_25196,N_21334,N_23462);
nand U25197 (N_25197,N_24082,N_22588);
nand U25198 (N_25198,N_22080,N_21508);
and U25199 (N_25199,N_21484,N_22171);
or U25200 (N_25200,N_22111,N_21075);
nor U25201 (N_25201,N_22883,N_20938);
nand U25202 (N_25202,N_24186,N_20314);
xor U25203 (N_25203,N_24858,N_22389);
nand U25204 (N_25204,N_22386,N_24907);
nand U25205 (N_25205,N_23582,N_20896);
and U25206 (N_25206,N_20232,N_23612);
nor U25207 (N_25207,N_24909,N_24988);
or U25208 (N_25208,N_20429,N_22249);
or U25209 (N_25209,N_21624,N_21105);
and U25210 (N_25210,N_22302,N_24626);
nor U25211 (N_25211,N_23835,N_23257);
and U25212 (N_25212,N_21711,N_21242);
or U25213 (N_25213,N_21729,N_23022);
xor U25214 (N_25214,N_24751,N_20006);
and U25215 (N_25215,N_22415,N_20167);
xnor U25216 (N_25216,N_23430,N_20401);
nand U25217 (N_25217,N_23440,N_23079);
nand U25218 (N_25218,N_22792,N_23058);
and U25219 (N_25219,N_21861,N_22925);
nand U25220 (N_25220,N_21579,N_21093);
or U25221 (N_25221,N_21289,N_23129);
or U25222 (N_25222,N_22696,N_22884);
nor U25223 (N_25223,N_22582,N_22810);
nor U25224 (N_25224,N_24881,N_24215);
nand U25225 (N_25225,N_21915,N_21137);
nand U25226 (N_25226,N_21054,N_21055);
or U25227 (N_25227,N_24653,N_20301);
nor U25228 (N_25228,N_24747,N_23412);
and U25229 (N_25229,N_22420,N_21260);
nand U25230 (N_25230,N_23140,N_23900);
xor U25231 (N_25231,N_23998,N_22467);
nor U25232 (N_25232,N_24787,N_22693);
nand U25233 (N_25233,N_22378,N_24978);
nand U25234 (N_25234,N_23486,N_24609);
nor U25235 (N_25235,N_22566,N_24783);
and U25236 (N_25236,N_21352,N_23823);
nor U25237 (N_25237,N_21397,N_21531);
and U25238 (N_25238,N_23465,N_23002);
nand U25239 (N_25239,N_21011,N_21704);
or U25240 (N_25240,N_24474,N_20142);
and U25241 (N_25241,N_24784,N_22134);
and U25242 (N_25242,N_20382,N_24305);
or U25243 (N_25243,N_22710,N_23378);
nor U25244 (N_25244,N_24996,N_21545);
xnor U25245 (N_25245,N_22517,N_20028);
nand U25246 (N_25246,N_20913,N_20927);
nand U25247 (N_25247,N_21057,N_20404);
xnor U25248 (N_25248,N_23424,N_23405);
nand U25249 (N_25249,N_20906,N_20564);
or U25250 (N_25250,N_20969,N_24865);
and U25251 (N_25251,N_20808,N_20015);
and U25252 (N_25252,N_20433,N_22784);
nand U25253 (N_25253,N_20182,N_21670);
nor U25254 (N_25254,N_23480,N_22245);
nand U25255 (N_25255,N_21693,N_21097);
nor U25256 (N_25256,N_23298,N_21628);
and U25257 (N_25257,N_22400,N_23825);
nor U25258 (N_25258,N_23986,N_23521);
and U25259 (N_25259,N_22511,N_22344);
or U25260 (N_25260,N_22256,N_20516);
nor U25261 (N_25261,N_24610,N_21991);
nand U25262 (N_25262,N_22225,N_22476);
nand U25263 (N_25263,N_22564,N_20496);
nor U25264 (N_25264,N_22599,N_22718);
nor U25265 (N_25265,N_24749,N_20671);
xnor U25266 (N_25266,N_21713,N_22198);
or U25267 (N_25267,N_20641,N_22266);
and U25268 (N_25268,N_21687,N_20278);
xor U25269 (N_25269,N_20818,N_22781);
xor U25270 (N_25270,N_23723,N_22546);
nand U25271 (N_25271,N_23426,N_22472);
or U25272 (N_25272,N_24723,N_22686);
or U25273 (N_25273,N_21286,N_21420);
and U25274 (N_25274,N_22677,N_21353);
and U25275 (N_25275,N_24745,N_22486);
xor U25276 (N_25276,N_23108,N_21518);
nor U25277 (N_25277,N_23077,N_22750);
xnor U25278 (N_25278,N_23122,N_21712);
and U25279 (N_25279,N_21956,N_21067);
nor U25280 (N_25280,N_21135,N_24932);
or U25281 (N_25281,N_22937,N_22755);
nand U25282 (N_25282,N_24199,N_20636);
nor U25283 (N_25283,N_20228,N_22875);
and U25284 (N_25284,N_23868,N_20681);
and U25285 (N_25285,N_20447,N_22159);
nor U25286 (N_25286,N_23935,N_23379);
nand U25287 (N_25287,N_20067,N_21482);
xnor U25288 (N_25288,N_22782,N_21835);
nand U25289 (N_25289,N_24330,N_24159);
or U25290 (N_25290,N_23862,N_21674);
nand U25291 (N_25291,N_24875,N_24313);
nand U25292 (N_25292,N_24143,N_22109);
nand U25293 (N_25293,N_22644,N_21277);
or U25294 (N_25294,N_23965,N_20281);
nand U25295 (N_25295,N_21782,N_21058);
or U25296 (N_25296,N_21877,N_24790);
nand U25297 (N_25297,N_22706,N_21283);
nor U25298 (N_25298,N_23566,N_22922);
xor U25299 (N_25299,N_23768,N_20711);
nor U25300 (N_25300,N_20384,N_23571);
and U25301 (N_25301,N_24761,N_21329);
and U25302 (N_25302,N_22192,N_21943);
nor U25303 (N_25303,N_24821,N_23202);
xor U25304 (N_25304,N_22948,N_21439);
nor U25305 (N_25305,N_23146,N_23280);
nor U25306 (N_25306,N_24684,N_21962);
xnor U25307 (N_25307,N_24237,N_23251);
nor U25308 (N_25308,N_20104,N_20687);
or U25309 (N_25309,N_22255,N_24493);
or U25310 (N_25310,N_23678,N_22126);
nand U25311 (N_25311,N_20470,N_23180);
nand U25312 (N_25312,N_21701,N_22658);
and U25313 (N_25313,N_24198,N_20653);
or U25314 (N_25314,N_20440,N_22805);
nor U25315 (N_25315,N_22243,N_21811);
nor U25316 (N_25316,N_20835,N_23515);
or U25317 (N_25317,N_24478,N_24897);
and U25318 (N_25318,N_21990,N_21441);
nor U25319 (N_25319,N_22612,N_22025);
xnor U25320 (N_25320,N_20910,N_24631);
and U25321 (N_25321,N_23767,N_23288);
nand U25322 (N_25322,N_23427,N_23074);
or U25323 (N_25323,N_20955,N_21014);
nand U25324 (N_25324,N_24166,N_21948);
xnor U25325 (N_25325,N_24121,N_20515);
xnor U25326 (N_25326,N_24637,N_20416);
and U25327 (N_25327,N_22469,N_22898);
xor U25328 (N_25328,N_21066,N_24984);
or U25329 (N_25329,N_24018,N_20246);
and U25330 (N_25330,N_23225,N_22777);
or U25331 (N_25331,N_20693,N_24872);
or U25332 (N_25332,N_20528,N_22031);
or U25333 (N_25333,N_22096,N_22870);
xnor U25334 (N_25334,N_22992,N_24464);
or U25335 (N_25335,N_20206,N_23247);
nand U25336 (N_25336,N_22452,N_24560);
xnor U25337 (N_25337,N_21878,N_24220);
nor U25338 (N_25338,N_22963,N_21113);
xor U25339 (N_25339,N_21279,N_22724);
xnor U25340 (N_25340,N_22355,N_23585);
nand U25341 (N_25341,N_24109,N_22229);
and U25342 (N_25342,N_20219,N_24027);
and U25343 (N_25343,N_20117,N_21400);
nand U25344 (N_25344,N_24389,N_22296);
nor U25345 (N_25345,N_21979,N_22675);
or U25346 (N_25346,N_21448,N_23335);
nand U25347 (N_25347,N_22058,N_22975);
nor U25348 (N_25348,N_21303,N_21740);
nand U25349 (N_25349,N_22801,N_20658);
nand U25350 (N_25350,N_20843,N_24476);
nand U25351 (N_25351,N_20058,N_20996);
or U25352 (N_25352,N_22627,N_20878);
nand U25353 (N_25353,N_20303,N_22095);
xnor U25354 (N_25354,N_22553,N_23149);
and U25355 (N_25355,N_23842,N_22104);
nand U25356 (N_25356,N_24038,N_20199);
and U25357 (N_25357,N_20611,N_20057);
and U25358 (N_25358,N_21069,N_21818);
xnor U25359 (N_25359,N_24910,N_20978);
or U25360 (N_25360,N_24321,N_24743);
xnor U25361 (N_25361,N_23836,N_22551);
and U25362 (N_25362,N_23957,N_21301);
and U25363 (N_25363,N_24976,N_24163);
nand U25364 (N_25364,N_20092,N_22999);
and U25365 (N_25365,N_20771,N_24295);
nand U25366 (N_25366,N_20541,N_22340);
nand U25367 (N_25367,N_21106,N_20097);
xor U25368 (N_25368,N_20582,N_22045);
nand U25369 (N_25369,N_24811,N_23501);
and U25370 (N_25370,N_22453,N_22086);
and U25371 (N_25371,N_20388,N_20511);
nor U25372 (N_25372,N_24710,N_24045);
xnor U25373 (N_25373,N_21843,N_23264);
xnor U25374 (N_25374,N_21407,N_23834);
or U25375 (N_25375,N_20225,N_24234);
or U25376 (N_25376,N_23624,N_24960);
and U25377 (N_25377,N_24598,N_24982);
and U25378 (N_25378,N_24167,N_23461);
nand U25379 (N_25379,N_22390,N_22924);
xnor U25380 (N_25380,N_24884,N_21882);
nand U25381 (N_25381,N_21070,N_22774);
nand U25382 (N_25382,N_20629,N_23743);
or U25383 (N_25383,N_21282,N_23605);
or U25384 (N_25384,N_20663,N_21913);
nor U25385 (N_25385,N_22939,N_21602);
and U25386 (N_25386,N_22769,N_20112);
or U25387 (N_25387,N_20634,N_22269);
nor U25388 (N_25388,N_22410,N_23824);
or U25389 (N_25389,N_20250,N_21427);
xor U25390 (N_25390,N_24519,N_20699);
nand U25391 (N_25391,N_22504,N_21188);
nand U25392 (N_25392,N_21424,N_23755);
or U25393 (N_25393,N_20234,N_20500);
and U25394 (N_25394,N_20529,N_21187);
or U25395 (N_25395,N_21176,N_23616);
nor U25396 (N_25396,N_20079,N_24418);
or U25397 (N_25397,N_23073,N_21829);
nor U25398 (N_25398,N_23702,N_24210);
nor U25399 (N_25399,N_23651,N_21037);
nor U25400 (N_25400,N_20831,N_24005);
xnor U25401 (N_25401,N_24336,N_22007);
and U25402 (N_25402,N_23629,N_20230);
nand U25403 (N_25403,N_22032,N_23062);
nand U25404 (N_25404,N_20914,N_20499);
or U25405 (N_25405,N_20369,N_24368);
or U25406 (N_25406,N_20976,N_22411);
xor U25407 (N_25407,N_20253,N_20148);
xor U25408 (N_25408,N_22280,N_24162);
or U25409 (N_25409,N_20434,N_22613);
or U25410 (N_25410,N_22023,N_20754);
xor U25411 (N_25411,N_20576,N_20543);
xnor U25412 (N_25412,N_20735,N_20152);
and U25413 (N_25413,N_20620,N_21378);
xnor U25414 (N_25414,N_21559,N_23713);
or U25415 (N_25415,N_21859,N_23738);
or U25416 (N_25416,N_23506,N_23961);
nand U25417 (N_25417,N_21733,N_21088);
and U25418 (N_25418,N_22170,N_20255);
and U25419 (N_25419,N_21453,N_20700);
xor U25420 (N_25420,N_22258,N_24232);
nor U25421 (N_25421,N_21024,N_20570);
xor U25422 (N_25422,N_22574,N_24097);
nor U25423 (N_25423,N_22608,N_23676);
or U25424 (N_25424,N_24028,N_21689);
nand U25425 (N_25425,N_24009,N_22972);
or U25426 (N_25426,N_24986,N_22220);
nor U25427 (N_25427,N_22908,N_22449);
and U25428 (N_25428,N_21230,N_21204);
or U25429 (N_25429,N_24472,N_22738);
nand U25430 (N_25430,N_22077,N_22580);
nor U25431 (N_25431,N_24507,N_22384);
xor U25432 (N_25432,N_23783,N_24475);
nand U25433 (N_25433,N_22811,N_21254);
nor U25434 (N_25434,N_23954,N_20909);
nor U25435 (N_25435,N_21042,N_23206);
or U25436 (N_25436,N_23761,N_22920);
and U25437 (N_25437,N_21321,N_21732);
nand U25438 (N_25438,N_21524,N_24180);
nor U25439 (N_25439,N_24957,N_23777);
nor U25440 (N_25440,N_21633,N_24345);
xnor U25441 (N_25441,N_22909,N_22763);
nor U25442 (N_25442,N_23204,N_21927);
xor U25443 (N_25443,N_23646,N_22442);
xnor U25444 (N_25444,N_20580,N_20612);
nor U25445 (N_25445,N_23942,N_23393);
xor U25446 (N_25446,N_21416,N_21389);
nand U25447 (N_25447,N_21431,N_23456);
nand U25448 (N_25448,N_24624,N_21068);
nor U25449 (N_25449,N_23137,N_24599);
nor U25450 (N_25450,N_23245,N_22707);
nand U25451 (N_25451,N_22815,N_21032);
nor U25452 (N_25452,N_22347,N_23828);
nand U25453 (N_25453,N_23897,N_22421);
nand U25454 (N_25454,N_22768,N_22751);
nor U25455 (N_25455,N_23775,N_23061);
nand U25456 (N_25456,N_24528,N_21863);
xnor U25457 (N_25457,N_21989,N_22153);
nor U25458 (N_25458,N_23508,N_23125);
xnor U25459 (N_25459,N_24411,N_22090);
xnor U25460 (N_25460,N_22005,N_21190);
and U25461 (N_25461,N_23326,N_23725);
xnor U25462 (N_25462,N_20038,N_20151);
and U25463 (N_25463,N_20351,N_22299);
and U25464 (N_25464,N_23425,N_22316);
and U25465 (N_25465,N_22114,N_21048);
nor U25466 (N_25466,N_21887,N_24654);
or U25467 (N_25467,N_22387,N_22146);
xnor U25468 (N_25468,N_20124,N_23159);
or U25469 (N_25469,N_21864,N_24194);
and U25470 (N_25470,N_23559,N_24573);
nand U25471 (N_25471,N_21534,N_22363);
and U25472 (N_25472,N_20443,N_20537);
nor U25473 (N_25473,N_20946,N_24269);
nand U25474 (N_25474,N_20951,N_21333);
nor U25475 (N_25475,N_23004,N_21671);
xnor U25476 (N_25476,N_21934,N_20348);
and U25477 (N_25477,N_20205,N_23788);
nor U25478 (N_25478,N_23679,N_24792);
and U25479 (N_25479,N_20875,N_21596);
nand U25480 (N_25480,N_23881,N_21734);
xnor U25481 (N_25481,N_23306,N_24522);
xnor U25482 (N_25482,N_23347,N_23940);
nand U25483 (N_25483,N_22455,N_20566);
nor U25484 (N_25484,N_21963,N_21474);
nand U25485 (N_25485,N_20651,N_24665);
nor U25486 (N_25486,N_24495,N_21942);
or U25487 (N_25487,N_21748,N_21937);
nor U25488 (N_25488,N_24852,N_22590);
nor U25489 (N_25489,N_21136,N_23352);
nor U25490 (N_25490,N_20956,N_24645);
xnor U25491 (N_25491,N_24035,N_21750);
xnor U25492 (N_25492,N_23476,N_20904);
nand U25493 (N_25493,N_21186,N_22770);
or U25494 (N_25494,N_20574,N_22246);
nand U25495 (N_25495,N_21884,N_23040);
nand U25496 (N_25496,N_24979,N_24025);
and U25497 (N_25497,N_23662,N_20784);
or U25498 (N_25498,N_21675,N_20394);
nor U25499 (N_25499,N_21769,N_20957);
xor U25500 (N_25500,N_20002,N_21590);
nor U25501 (N_25501,N_23996,N_21382);
xor U25502 (N_25502,N_23115,N_24990);
nor U25503 (N_25503,N_21386,N_24421);
nand U25504 (N_25504,N_21598,N_20939);
xnor U25505 (N_25505,N_22250,N_22403);
and U25506 (N_25506,N_21184,N_24732);
and U25507 (N_25507,N_21033,N_23663);
nor U25508 (N_25508,N_21259,N_21377);
and U25509 (N_25509,N_21774,N_20237);
nand U25510 (N_25510,N_22712,N_21065);
xnor U25511 (N_25511,N_23056,N_22300);
and U25512 (N_25512,N_23356,N_24482);
nor U25513 (N_25513,N_22408,N_22611);
or U25514 (N_25514,N_24931,N_23016);
and U25515 (N_25515,N_21257,N_24074);
nand U25516 (N_25516,N_23974,N_23595);
xnor U25517 (N_25517,N_21710,N_23766);
or U25518 (N_25518,N_22181,N_22459);
nor U25519 (N_25519,N_22965,N_23421);
and U25520 (N_25520,N_23402,N_21660);
or U25521 (N_25521,N_21383,N_23441);
xor U25522 (N_25522,N_23519,N_24033);
nand U25523 (N_25523,N_23574,N_20763);
nand U25524 (N_25524,N_22097,N_21573);
nor U25525 (N_25525,N_22259,N_22430);
nand U25526 (N_25526,N_21457,N_20273);
nand U25527 (N_25527,N_21690,N_21274);
nor U25528 (N_25528,N_24454,N_20928);
nor U25529 (N_25529,N_21166,N_22227);
and U25530 (N_25530,N_22149,N_24221);
nor U25531 (N_25531,N_23431,N_24547);
xor U25532 (N_25532,N_21185,N_22085);
nand U25533 (N_25533,N_22368,N_23760);
and U25534 (N_25534,N_20202,N_23317);
xnor U25535 (N_25535,N_24849,N_24349);
xor U25536 (N_25536,N_24998,N_23187);
xor U25537 (N_25537,N_21644,N_24533);
xnor U25538 (N_25538,N_22779,N_21865);
xor U25539 (N_25539,N_22961,N_24563);
nand U25540 (N_25540,N_21198,N_23964);
nor U25541 (N_25541,N_23294,N_24669);
nand U25542 (N_25542,N_23351,N_22711);
xor U25543 (N_25543,N_24453,N_23036);
or U25544 (N_25544,N_24217,N_21414);
nand U25545 (N_25545,N_22206,N_24552);
or U25546 (N_25546,N_23096,N_23232);
or U25547 (N_25547,N_24249,N_20254);
or U25548 (N_25548,N_23953,N_20519);
nor U25549 (N_25549,N_21575,N_24110);
and U25550 (N_25550,N_22332,N_22622);
xor U25551 (N_25551,N_24322,N_24452);
nor U25552 (N_25552,N_22480,N_24520);
and U25553 (N_25553,N_24002,N_23630);
xor U25554 (N_25554,N_23837,N_23404);
nor U25555 (N_25555,N_20153,N_23549);
or U25556 (N_25556,N_20768,N_21500);
nor U25557 (N_25557,N_21376,N_20765);
or U25558 (N_25558,N_22092,N_24758);
nand U25559 (N_25559,N_24264,N_21077);
xor U25560 (N_25560,N_24619,N_22860);
nand U25561 (N_25561,N_21401,N_21973);
or U25562 (N_25562,N_21694,N_24332);
or U25563 (N_25563,N_23523,N_23231);
xor U25564 (N_25564,N_21777,N_20999);
and U25565 (N_25565,N_21201,N_20773);
or U25566 (N_25566,N_23176,N_23390);
nor U25567 (N_25567,N_20274,N_21908);
nand U25568 (N_25568,N_21911,N_21563);
and U25569 (N_25569,N_20781,N_21415);
and U25570 (N_25570,N_20258,N_23367);
nand U25571 (N_25571,N_23887,N_21758);
or U25572 (N_25572,N_21300,N_20296);
nor U25573 (N_25573,N_23373,N_24735);
nand U25574 (N_25574,N_24613,N_23154);
nand U25575 (N_25575,N_22645,N_20544);
and U25576 (N_25576,N_23455,N_21869);
xnor U25577 (N_25577,N_22679,N_20517);
nand U25578 (N_25578,N_22518,N_24333);
nand U25579 (N_25579,N_21668,N_20606);
xnor U25580 (N_25580,N_23793,N_22803);
nand U25581 (N_25581,N_24196,N_22901);
or U25582 (N_25582,N_22643,N_23711);
nand U25583 (N_25583,N_24939,N_24611);
or U25584 (N_25584,N_22308,N_23028);
and U25585 (N_25585,N_20106,N_24632);
and U25586 (N_25586,N_22534,N_20422);
or U25587 (N_25587,N_22448,N_20837);
nand U25588 (N_25588,N_23401,N_21672);
and U25589 (N_25589,N_24244,N_23433);
nand U25590 (N_25590,N_21357,N_21349);
nand U25591 (N_25591,N_22562,N_21623);
xnor U25592 (N_25592,N_23721,N_20887);
xor U25593 (N_25593,N_23445,N_23174);
and U25594 (N_25594,N_22374,N_21700);
or U25595 (N_25595,N_20494,N_24235);
nand U25596 (N_25596,N_23089,N_23918);
xor U25597 (N_25597,N_23548,N_21211);
or U25598 (N_25598,N_21735,N_20802);
xnor U25599 (N_25599,N_23106,N_21543);
and U25600 (N_25600,N_23119,N_20832);
and U25601 (N_25601,N_23141,N_23608);
xnor U25602 (N_25602,N_21061,N_24207);
xnor U25603 (N_25603,N_22823,N_20959);
and U25604 (N_25604,N_20372,N_23578);
nand U25605 (N_25605,N_20746,N_24625);
or U25606 (N_25606,N_22385,N_23551);
nand U25607 (N_25607,N_24843,N_23849);
xor U25608 (N_25608,N_22284,N_24980);
nor U25609 (N_25609,N_22624,N_23806);
xor U25610 (N_25610,N_20310,N_23299);
or U25611 (N_25611,N_20855,N_24832);
nor U25612 (N_25612,N_24700,N_20925);
nand U25613 (N_25613,N_23195,N_24281);
nor U25614 (N_25614,N_24096,N_22951);
nor U25615 (N_25615,N_24768,N_22057);
nor U25616 (N_25616,N_24945,N_24947);
or U25617 (N_25617,N_21161,N_22075);
and U25618 (N_25618,N_22787,N_22900);
and U25619 (N_25619,N_21629,N_21122);
nor U25620 (N_25620,N_22491,N_24728);
and U25621 (N_25621,N_23165,N_20324);
and U25622 (N_25622,N_20346,N_23977);
xor U25623 (N_25623,N_23820,N_23092);
nor U25624 (N_25624,N_23261,N_21101);
and U25625 (N_25625,N_20170,N_20136);
xnor U25626 (N_25626,N_23220,N_23221);
xor U25627 (N_25627,N_21746,N_20677);
or U25628 (N_25628,N_20625,N_24602);
or U25629 (N_25629,N_20851,N_23109);
nor U25630 (N_25630,N_20169,N_24915);
nor U25631 (N_25631,N_22461,N_21521);
and U25632 (N_25632,N_24886,N_24209);
or U25633 (N_25633,N_21297,N_21359);
or U25634 (N_25634,N_21139,N_20102);
or U25635 (N_25635,N_21862,N_24185);
nand U25636 (N_25636,N_23592,N_24456);
and U25637 (N_25637,N_21647,N_21847);
or U25638 (N_25638,N_23510,N_24913);
xor U25639 (N_25639,N_23026,N_21040);
nand U25640 (N_25640,N_24856,N_21914);
or U25641 (N_25641,N_20391,N_20751);
and U25642 (N_25642,N_20005,N_22257);
and U25643 (N_25643,N_24558,N_22053);
or U25644 (N_25644,N_24657,N_23601);
nor U25645 (N_25645,N_20012,N_20727);
nand U25646 (N_25646,N_23325,N_24413);
xnor U25647 (N_25647,N_20269,N_23305);
nor U25648 (N_25648,N_24054,N_22484);
xnor U25649 (N_25649,N_21541,N_22274);
nand U25650 (N_25650,N_23504,N_20125);
nor U25651 (N_25651,N_20633,N_20180);
nand U25652 (N_25652,N_20617,N_24791);
nand U25653 (N_25653,N_24702,N_20270);
nor U25654 (N_25654,N_23917,N_24680);
xor U25655 (N_25655,N_24975,N_20750);
xor U25656 (N_25656,N_22573,N_21371);
and U25657 (N_25657,N_20645,N_20858);
or U25658 (N_25658,N_20066,N_22988);
nand U25659 (N_25659,N_21396,N_24238);
and U25660 (N_25660,N_21812,N_22688);
and U25661 (N_25661,N_23891,N_24090);
or U25662 (N_25662,N_21350,N_22589);
and U25663 (N_25663,N_22941,N_22709);
nand U25664 (N_25664,N_22583,N_20705);
and U25665 (N_25665,N_22354,N_24795);
nor U25666 (N_25666,N_23117,N_21762);
or U25667 (N_25667,N_23706,N_23179);
nor U25668 (N_25668,N_21464,N_22167);
xnor U25669 (N_25669,N_21591,N_24000);
nor U25670 (N_25670,N_21739,N_23271);
nor U25671 (N_25671,N_20584,N_23444);
xnor U25672 (N_25672,N_23555,N_23346);
xor U25673 (N_25673,N_21823,N_23331);
and U25674 (N_25674,N_21890,N_22074);
or U25675 (N_25675,N_22121,N_22783);
xor U25676 (N_25676,N_22840,N_20341);
xnor U25677 (N_25677,N_20108,N_22959);
and U25678 (N_25678,N_24880,N_22231);
nor U25679 (N_25679,N_20605,N_21085);
and U25680 (N_25680,N_21246,N_21398);
nand U25681 (N_25681,N_21243,N_22911);
and U25682 (N_25682,N_20526,N_21327);
and U25683 (N_25683,N_24906,N_21392);
nand U25684 (N_25684,N_23126,N_20929);
nor U25685 (N_25685,N_20173,N_20538);
and U25686 (N_25686,N_23959,N_20579);
nand U25687 (N_25687,N_21368,N_22021);
or U25688 (N_25688,N_23472,N_24892);
nor U25689 (N_25689,N_20053,N_23014);
nor U25690 (N_25690,N_20485,N_24652);
nor U25691 (N_25691,N_24388,N_22929);
nor U25692 (N_25692,N_21302,N_23268);
and U25693 (N_25693,N_20958,N_24717);
or U25694 (N_25694,N_20138,N_24851);
xnor U25695 (N_25695,N_22692,N_23491);
nor U25696 (N_25696,N_21630,N_20798);
and U25697 (N_25697,N_22575,N_24663);
nand U25698 (N_25698,N_24172,N_23169);
xnor U25699 (N_25699,N_20474,N_20383);
xor U25700 (N_25700,N_23720,N_23950);
nor U25701 (N_25701,N_20505,N_21844);
and U25702 (N_25702,N_23477,N_22366);
xnor U25703 (N_25703,N_21503,N_20312);
and U25704 (N_25704,N_23602,N_22775);
nor U25705 (N_25705,N_20337,N_22767);
nor U25706 (N_25706,N_22543,N_22184);
or U25707 (N_25707,N_20860,N_23330);
xor U25708 (N_25708,N_22670,N_21245);
xor U25709 (N_25709,N_21722,N_23841);
and U25710 (N_25710,N_24772,N_24689);
or U25711 (N_25711,N_22169,N_21893);
nand U25712 (N_25712,N_22002,N_24845);
nor U25713 (N_25713,N_20032,N_22772);
or U25714 (N_25714,N_21759,N_21410);
or U25715 (N_25715,N_23854,N_23173);
xor U25716 (N_25716,N_23255,N_21542);
or U25717 (N_25717,N_24788,N_22103);
nand U25718 (N_25718,N_22158,N_20221);
xnor U25719 (N_25719,N_24859,N_24174);
nor U25720 (N_25720,N_21403,N_23300);
or U25721 (N_25721,N_20898,N_23552);
nand U25722 (N_25722,N_24600,N_20662);
and U25723 (N_25723,N_24177,N_20774);
nand U25724 (N_25724,N_24759,N_20469);
xor U25725 (N_25725,N_23383,N_23816);
and U25726 (N_25726,N_22623,N_20670);
nor U25727 (N_25727,N_20578,N_22218);
nor U25728 (N_25728,N_22592,N_24691);
xnor U25729 (N_25729,N_20039,N_23034);
xor U25730 (N_25730,N_23355,N_22325);
nand U25731 (N_25731,N_24967,N_22321);
xor U25732 (N_25732,N_21226,N_24922);
nor U25733 (N_25733,N_21885,N_23745);
xor U25734 (N_25734,N_24918,N_24348);
nor U25735 (N_25735,N_20643,N_23447);
and U25736 (N_25736,N_21967,N_21520);
nor U25737 (N_25737,N_23417,N_24328);
and U25738 (N_25738,N_20395,N_24325);
nor U25739 (N_25739,N_23889,N_23481);
nand U25740 (N_25740,N_21880,N_23254);
xnor U25741 (N_25741,N_24398,N_23558);
xor U25742 (N_25742,N_23031,N_23201);
nor U25743 (N_25743,N_22843,N_21646);
nand U25744 (N_25744,N_21331,N_23442);
nand U25745 (N_25745,N_24707,N_23547);
nor U25746 (N_25746,N_24324,N_22203);
and U25747 (N_25747,N_21525,N_20189);
xnor U25748 (N_25748,N_24111,N_24155);
nand U25749 (N_25749,N_20007,N_22078);
xnor U25750 (N_25750,N_23037,N_21030);
xor U25751 (N_25751,N_23270,N_24291);
and U25752 (N_25752,N_21062,N_24424);
and U25753 (N_25753,N_24981,N_20019);
xor U25754 (N_25754,N_20982,N_21940);
nand U25755 (N_25755,N_23072,N_21567);
nand U25756 (N_25756,N_23018,N_22849);
xor U25757 (N_25757,N_24867,N_22721);
xor U25758 (N_25758,N_22604,N_21565);
and U25759 (N_25759,N_20095,N_22377);
and U25760 (N_25760,N_24357,N_23650);
or U25761 (N_25761,N_20420,N_23576);
or U25762 (N_25762,N_22819,N_22736);
and U25763 (N_25763,N_23588,N_23328);
or U25764 (N_25764,N_20917,N_24995);
nand U25765 (N_25765,N_24353,N_22425);
nor U25766 (N_25766,N_22514,N_23934);
and U25767 (N_25767,N_24935,N_23786);
nor U25768 (N_25768,N_24703,N_24289);
or U25769 (N_25769,N_20827,N_23933);
nor U25770 (N_25770,N_20060,N_23923);
xnor U25771 (N_25771,N_21540,N_20306);
nand U25772 (N_25772,N_21501,N_20954);
xnor U25773 (N_25773,N_21152,N_21318);
xnor U25774 (N_25774,N_20730,N_21547);
nor U25775 (N_25775,N_23333,N_21269);
or U25776 (N_25776,N_20162,N_20088);
and U25777 (N_25777,N_22329,N_23997);
xnor U25778 (N_25778,N_23970,N_21324);
or U25779 (N_25779,N_23069,N_23597);
nor U25780 (N_25780,N_23978,N_20527);
and U25781 (N_25781,N_20532,N_24574);
nor U25782 (N_25782,N_24127,N_21892);
or U25783 (N_25783,N_21183,N_22946);
and U25784 (N_25784,N_21255,N_23438);
nand U25785 (N_25785,N_21043,N_20672);
or U25786 (N_25786,N_20607,N_24550);
nor U25787 (N_25787,N_20806,N_23265);
nand U25788 (N_25788,N_24427,N_23914);
nor U25789 (N_25789,N_22567,N_23336);
nor U25790 (N_25790,N_24687,N_22671);
xor U25791 (N_25791,N_24734,N_23916);
xnor U25792 (N_25792,N_22488,N_20044);
nand U25793 (N_25793,N_24231,N_22757);
xor U25794 (N_25794,N_20050,N_22748);
nand U25795 (N_25795,N_23064,N_22866);
and U25796 (N_25796,N_20047,N_23172);
xnor U25797 (N_25797,N_23973,N_22863);
and U25798 (N_25798,N_22962,N_23683);
or U25799 (N_25799,N_20271,N_21745);
or U25800 (N_25800,N_22265,N_22099);
or U25801 (N_25801,N_20145,N_20839);
nor U25802 (N_25802,N_24314,N_21576);
nand U25803 (N_25803,N_23980,N_24262);
nor U25804 (N_25804,N_20673,N_22353);
nor U25805 (N_25805,N_21379,N_22331);
and U25806 (N_25806,N_23946,N_24084);
nand U25807 (N_25807,N_21619,N_20975);
or U25808 (N_25808,N_23386,N_24065);
and U25809 (N_25809,N_20087,N_21631);
or U25810 (N_25810,N_24259,N_24075);
and U25811 (N_25811,N_23643,N_21850);
or U25812 (N_25812,N_22905,N_22594);
or U25813 (N_25813,N_22471,N_22684);
xnor U25814 (N_25814,N_23493,N_23790);
xnor U25815 (N_25815,N_22600,N_23338);
nand U25816 (N_25816,N_24003,N_22230);
or U25817 (N_25817,N_22727,N_21522);
nor U25818 (N_25818,N_24770,N_23360);
nand U25819 (N_25819,N_22433,N_21116);
or U25820 (N_25820,N_22487,N_20504);
xnor U25821 (N_25821,N_20589,N_23628);
nor U25822 (N_25822,N_21881,N_24712);
or U25823 (N_25823,N_22116,N_24603);
xor U25824 (N_25824,N_23927,N_21587);
and U25825 (N_25825,N_24921,N_24773);
or U25826 (N_25826,N_22797,N_22298);
nand U25827 (N_25827,N_20698,N_24334);
xor U25828 (N_25828,N_24079,N_22113);
or U25829 (N_25829,N_24970,N_21328);
and U25830 (N_25830,N_20708,N_23925);
nand U25831 (N_25831,N_24704,N_22665);
nor U25832 (N_25832,N_22731,N_21493);
xnor U25833 (N_25833,N_24888,N_22263);
xor U25834 (N_25834,N_20565,N_22859);
or U25835 (N_25835,N_20863,N_23621);
xor U25836 (N_25836,N_23705,N_23698);
or U25837 (N_25837,N_24195,N_23323);
and U25838 (N_25838,N_21127,N_22424);
and U25839 (N_25839,N_22142,N_24165);
nand U25840 (N_25840,N_24042,N_20680);
or U25841 (N_25841,N_20801,N_20669);
or U25842 (N_25842,N_24070,N_24088);
xor U25843 (N_25843,N_22180,N_21047);
nand U25844 (N_25844,N_21663,N_20211);
and U25845 (N_25845,N_24125,N_23478);
nand U25846 (N_25846,N_20070,N_21237);
or U25847 (N_25847,N_20506,N_20503);
nor U25848 (N_25848,N_21015,N_22493);
xnor U25849 (N_25849,N_24137,N_22212);
nor U25850 (N_25850,N_24211,N_22470);
or U25851 (N_25851,N_20571,N_21073);
and U25852 (N_25852,N_20782,N_22969);
xor U25853 (N_25853,N_22680,N_24069);
xor U25854 (N_25854,N_22295,N_22894);
nand U25855 (N_25855,N_21150,N_21307);
and U25856 (N_25856,N_21191,N_21529);
and U25857 (N_25857,N_24987,N_23369);
or U25858 (N_25858,N_23522,N_23733);
and U25859 (N_25859,N_21857,N_21281);
or U25860 (N_25860,N_20461,N_20945);
nand U25861 (N_25861,N_23505,N_22915);
nand U25862 (N_25862,N_20297,N_24448);
or U25863 (N_25863,N_23693,N_20783);
nor U25864 (N_25864,N_24176,N_20176);
xnor U25865 (N_25865,N_24634,N_23048);
nor U25866 (N_25866,N_21820,N_24565);
nand U25867 (N_25867,N_23876,N_20283);
xnor U25868 (N_25868,N_22401,N_21051);
xnor U25869 (N_25869,N_21340,N_21517);
or U25870 (N_25870,N_24650,N_21200);
xnor U25871 (N_25871,N_21952,N_23839);
and U25872 (N_25872,N_21380,N_20872);
and U25873 (N_25873,N_22115,N_22931);
and U25874 (N_25874,N_24595,N_22022);
xor U25875 (N_25875,N_21322,N_23138);
xnor U25876 (N_25876,N_20885,N_24030);
nand U25877 (N_25877,N_23278,N_24809);
nand U25878 (N_25878,N_22858,N_23792);
nor U25879 (N_25879,N_20853,N_20729);
and U25880 (N_25880,N_20998,N_22394);
xor U25881 (N_25881,N_22084,N_22867);
or U25882 (N_25882,N_21430,N_23182);
nand U25883 (N_25883,N_24581,N_22327);
nor U25884 (N_25884,N_21175,N_20891);
or U25885 (N_25885,N_23253,N_24557);
nand U25886 (N_25886,N_24678,N_22737);
xnor U25887 (N_25887,N_24021,N_24399);
xor U25888 (N_25888,N_22489,N_20599);
xor U25889 (N_25889,N_22070,N_20456);
or U25890 (N_25890,N_22734,N_22044);
xor U25891 (N_25891,N_21221,N_21858);
and U25892 (N_25892,N_23874,N_24460);
and U25893 (N_25893,N_22285,N_24391);
xor U25894 (N_25894,N_20405,N_23878);
xnor U25895 (N_25895,N_22117,N_23293);
xor U25896 (N_25896,N_23006,N_21535);
nand U25897 (N_25897,N_24529,N_24819);
nor U25898 (N_25898,N_22055,N_20967);
xor U25899 (N_25899,N_23737,N_24635);
and U25900 (N_25900,N_23619,N_22479);
or U25901 (N_25901,N_23668,N_23671);
and U25902 (N_25902,N_21805,N_22541);
or U25903 (N_25903,N_23511,N_24455);
nand U25904 (N_25904,N_23060,N_22143);
and U25905 (N_25905,N_23029,N_21707);
xnor U25906 (N_25906,N_20777,N_24912);
nand U25907 (N_25907,N_20174,N_20327);
or U25908 (N_25908,N_22703,N_22978);
xnor U25909 (N_25909,N_22216,N_24868);
nor U25910 (N_25910,N_21171,N_22252);
xor U25911 (N_25911,N_22602,N_24504);
and U25912 (N_25912,N_23327,N_21404);
xor U25913 (N_25913,N_23802,N_23982);
or U25914 (N_25914,N_22607,N_20014);
xnor U25915 (N_25915,N_24490,N_20739);
nor U25916 (N_25916,N_23432,N_20640);
and U25917 (N_25917,N_20040,N_24430);
nand U25918 (N_25918,N_21635,N_20399);
xnor U25919 (N_25919,N_24359,N_22242);
and U25920 (N_25920,N_23316,N_24369);
nor U25921 (N_25921,N_22209,N_21691);
nor U25922 (N_25922,N_20023,N_24484);
nor U25923 (N_25923,N_20738,N_24469);
nand U25924 (N_25924,N_23665,N_23148);
xnor U25925 (N_25925,N_21572,N_22289);
and U25926 (N_25926,N_22947,N_21783);
xnor U25927 (N_25927,N_24060,N_22505);
or U25928 (N_25928,N_23068,N_23847);
and U25929 (N_25929,N_24640,N_23540);
nand U25930 (N_25930,N_20844,N_23649);
nor U25931 (N_25931,N_20847,N_21118);
or U25932 (N_25932,N_23237,N_23798);
xor U25933 (N_25933,N_21298,N_23675);
and U25934 (N_25934,N_20706,N_22391);
xnor U25935 (N_25935,N_24122,N_24887);
nand U25936 (N_25936,N_22854,N_23968);
nand U25937 (N_25937,N_22839,N_23210);
and U25938 (N_25938,N_21029,N_20650);
nand U25939 (N_25939,N_22530,N_21494);
and U25940 (N_25940,N_20175,N_22899);
nor U25941 (N_25941,N_21926,N_24317);
or U25942 (N_25942,N_24937,N_23276);
nor U25943 (N_25943,N_20741,N_21552);
or U25944 (N_25944,N_20409,N_24847);
or U25945 (N_25945,N_21028,N_22064);
and U25946 (N_25946,N_22598,N_24877);
and U25947 (N_25947,N_24245,N_21146);
nor U25948 (N_25948,N_22923,N_21898);
nand U25949 (N_25949,N_20350,N_24267);
nor U25950 (N_25950,N_20888,N_22427);
nor U25951 (N_25951,N_24390,N_22195);
nor U25952 (N_25952,N_24335,N_22637);
or U25953 (N_25953,N_24806,N_21326);
or U25954 (N_25954,N_24374,N_22609);
or U25955 (N_25955,N_24692,N_20583);
nand U25956 (N_25956,N_20766,N_21220);
and U25957 (N_25957,N_22254,N_23163);
nor U25958 (N_25958,N_22814,N_21316);
nor U25959 (N_25959,N_21408,N_21609);
xor U25960 (N_25960,N_21613,N_22926);
or U25961 (N_25961,N_20336,N_24246);
xnor U25962 (N_25962,N_24200,N_24955);
xnor U25963 (N_25963,N_23435,N_22593);
xor U25964 (N_25964,N_20791,N_24439);
and U25965 (N_25965,N_22788,N_23177);
or U25966 (N_25966,N_23136,N_22046);
nand U25967 (N_25967,N_21643,N_24973);
nor U25968 (N_25968,N_24733,N_20074);
or U25969 (N_25969,N_23735,N_22935);
nand U25970 (N_25970,N_21723,N_23805);
and U25971 (N_25971,N_22197,N_22990);
or U25972 (N_25972,N_24952,N_24874);
or U25973 (N_25973,N_24890,N_21738);
nor U25974 (N_25974,N_23027,N_22656);
xnor U25975 (N_25975,N_20361,N_24300);
nand U25976 (N_25976,N_20343,N_24901);
nor U25977 (N_25977,N_24487,N_21141);
nor U25978 (N_25978,N_23500,N_20282);
nand U25979 (N_25979,N_21945,N_24059);
xor U25980 (N_25980,N_22928,N_24248);
xor U25981 (N_25981,N_20974,N_20287);
nand U25982 (N_25982,N_24927,N_22910);
xor U25983 (N_25983,N_24446,N_24741);
and U25984 (N_25984,N_20119,N_20842);
xnor U25985 (N_25985,N_22024,N_20455);
nor U25986 (N_25986,N_20449,N_22610);
xor U25987 (N_25987,N_20613,N_23844);
and U25988 (N_25988,N_20638,N_22000);
nor U25989 (N_25989,N_23707,N_23641);
nand U25990 (N_25990,N_22367,N_21537);
nand U25991 (N_25991,N_21581,N_20227);
nand U25992 (N_25992,N_23238,N_24168);
nor U25993 (N_25993,N_22507,N_22560);
and U25994 (N_25994,N_22087,N_20562);
xor U25995 (N_25995,N_21921,N_20657);
or U25996 (N_25996,N_23888,N_21406);
and U25997 (N_25997,N_23568,N_22572);
and U25998 (N_25998,N_24471,N_21652);
or U25999 (N_25999,N_22542,N_21096);
or U26000 (N_26000,N_22793,N_20073);
xnor U26001 (N_26001,N_23944,N_21941);
xor U26002 (N_26002,N_22139,N_22303);
nand U26003 (N_26003,N_23587,N_24617);
and U26004 (N_26004,N_23971,N_22112);
xnor U26005 (N_26005,N_20085,N_20139);
and U26006 (N_26006,N_23262,N_24564);
nand U26007 (N_26007,N_21059,N_23945);
xnor U26008 (N_26008,N_21614,N_20857);
or U26009 (N_26009,N_21617,N_22155);
and U26010 (N_26010,N_21034,N_21627);
or U26011 (N_26011,N_22440,N_24659);
nor U26012 (N_26012,N_22210,N_21013);
nand U26013 (N_26013,N_20962,N_22676);
xnor U26014 (N_26014,N_21080,N_22290);
xor U26015 (N_26015,N_23086,N_22683);
xor U26016 (N_26016,N_21459,N_20816);
nand U26017 (N_26017,N_20980,N_23087);
nor U26018 (N_26018,N_20315,N_22287);
nand U26019 (N_26019,N_22701,N_20289);
and U26020 (N_26020,N_20703,N_24160);
or U26021 (N_26021,N_20375,N_23598);
and U26022 (N_26022,N_20359,N_20702);
xor U26023 (N_26023,N_24444,N_20772);
or U26024 (N_26024,N_20370,N_24814);
nand U26025 (N_26025,N_22740,N_22382);
nand U26026 (N_26026,N_23260,N_23610);
or U26027 (N_26027,N_20787,N_22651);
nand U26028 (N_26028,N_21249,N_24278);
nor U26029 (N_26029,N_20497,N_23217);
nor U26030 (N_26030,N_24748,N_22700);
nor U26031 (N_26031,N_24403,N_23189);
or U26032 (N_26032,N_20757,N_20726);
or U26033 (N_26033,N_22723,N_24530);
xor U26034 (N_26034,N_22405,N_24182);
nor U26035 (N_26035,N_24964,N_20964);
and U26036 (N_26036,N_21364,N_24306);
xor U26037 (N_26037,N_24179,N_20569);
xor U26038 (N_26038,N_23282,N_20435);
nor U26039 (N_26039,N_21776,N_22056);
and U26040 (N_26040,N_23371,N_20815);
xor U26041 (N_26041,N_24461,N_20534);
or U26042 (N_26042,N_22164,N_24311);
nor U26043 (N_26043,N_22539,N_24508);
nand U26044 (N_26044,N_22841,N_20308);
and U26045 (N_26045,N_23162,N_24457);
nor U26046 (N_26046,N_21848,N_20021);
or U26047 (N_26047,N_22964,N_23784);
or U26048 (N_26048,N_20457,N_23015);
and U26049 (N_26049,N_23133,N_21639);
xor U26050 (N_26050,N_20432,N_23422);
nor U26051 (N_26051,N_24739,N_21010);
nand U26052 (N_26052,N_23279,N_20603);
or U26053 (N_26053,N_21923,N_22986);
nor U26054 (N_26054,N_24799,N_20123);
nor U26055 (N_26055,N_22873,N_22906);
nand U26056 (N_26056,N_24954,N_22276);
nor U26057 (N_26057,N_20970,N_20713);
nand U26058 (N_26058,N_24974,N_22392);
and U26059 (N_26059,N_24683,N_23730);
and U26060 (N_26060,N_22501,N_23000);
and U26061 (N_26061,N_22027,N_22887);
or U26062 (N_26062,N_22156,N_20387);
or U26063 (N_26063,N_22343,N_20981);
xor U26064 (N_26064,N_21938,N_21605);
xor U26065 (N_26065,N_22862,N_24309);
nand U26066 (N_26066,N_24649,N_21451);
and U26067 (N_26067,N_22809,N_22271);
xnor U26068 (N_26068,N_24646,N_23458);
xor U26069 (N_26069,N_21875,N_23315);
nor U26070 (N_26070,N_20134,N_24420);
nor U26071 (N_26071,N_20036,N_24242);
and U26072 (N_26072,N_21483,N_22076);
xnor U26073 (N_26073,N_24148,N_24376);
and U26074 (N_26074,N_22513,N_21218);
nand U26075 (N_26075,N_24642,N_23076);
and U26076 (N_26076,N_24342,N_24969);
or U26077 (N_26077,N_20208,N_24340);
nor U26078 (N_26078,N_24812,N_21978);
and U26079 (N_26079,N_23969,N_20160);
nor U26080 (N_26080,N_21790,N_22147);
or U26081 (N_26081,N_20454,N_23171);
nor U26082 (N_26082,N_24343,N_23560);
xnor U26083 (N_26083,N_24365,N_22136);
nand U26084 (N_26084,N_23657,N_21256);
xnor U26085 (N_26085,N_20261,N_22091);
nand U26086 (N_26086,N_23600,N_24606);
and U26087 (N_26087,N_22338,N_24032);
xor U26088 (N_26088,N_24671,N_20172);
xor U26089 (N_26089,N_22399,N_22606);
and U26090 (N_26090,N_22960,N_22483);
nor U26091 (N_26091,N_23509,N_24549);
or U26092 (N_26092,N_24762,N_24586);
nand U26093 (N_26093,N_21555,N_23308);
xor U26094 (N_26094,N_23801,N_21958);
xnor U26095 (N_26095,N_24431,N_21270);
and U26096 (N_26096,N_23054,N_24026);
and U26097 (N_26097,N_22065,N_21082);
nor U26098 (N_26098,N_22145,N_24303);
and U26099 (N_26099,N_20356,N_22376);
xnor U26100 (N_26100,N_21253,N_24746);
xor U26101 (N_26101,N_20795,N_20291);
xor U26102 (N_26102,N_22342,N_20575);
and U26103 (N_26103,N_21130,N_24375);
nor U26104 (N_26104,N_20922,N_20238);
or U26105 (N_26105,N_21145,N_22640);
nand U26106 (N_26106,N_20100,N_20290);
and U26107 (N_26107,N_24417,N_23846);
nor U26108 (N_26108,N_23542,N_21180);
nor U26109 (N_26109,N_22423,N_21977);
or U26110 (N_26110,N_21463,N_24869);
or U26111 (N_26111,N_20193,N_23563);
nand U26112 (N_26112,N_20916,N_21405);
nand U26113 (N_26113,N_21901,N_22881);
or U26114 (N_26114,N_20732,N_23208);
and U26115 (N_26115,N_24006,N_24250);
or U26116 (N_26116,N_21677,N_24802);
xnor U26117 (N_26117,N_22702,N_24326);
and U26118 (N_26118,N_22621,N_23105);
or U26119 (N_26119,N_23128,N_20062);
nand U26120 (N_26120,N_22083,N_20338);
or U26121 (N_26121,N_22855,N_23561);
nor U26122 (N_26122,N_20817,N_20923);
nor U26123 (N_26123,N_23017,N_23170);
or U26124 (N_26124,N_24757,N_24071);
or U26125 (N_26125,N_22311,N_21214);
nor U26126 (N_26126,N_21479,N_23984);
nor U26127 (N_26127,N_20897,N_21466);
nor U26128 (N_26128,N_22100,N_23502);
nand U26129 (N_26129,N_21399,N_22011);
xor U26130 (N_26130,N_20328,N_24655);
xor U26131 (N_26131,N_24150,N_24972);
xnor U26132 (N_26132,N_21928,N_21595);
xor U26133 (N_26133,N_24266,N_24156);
and U26134 (N_26134,N_20477,N_22654);
nand U26135 (N_26135,N_22334,N_23949);
nor U26136 (N_26136,N_20299,N_23193);
nor U26137 (N_26137,N_21830,N_20304);
nor U26138 (N_26138,N_22460,N_21786);
nand U26139 (N_26139,N_22586,N_24286);
or U26140 (N_26140,N_23219,N_24046);
and U26141 (N_26141,N_22704,N_24824);
nor U26142 (N_26142,N_22557,N_20334);
and U26143 (N_26143,N_24985,N_22519);
xor U26144 (N_26144,N_20320,N_20275);
and U26145 (N_26145,N_23372,N_22932);
and U26146 (N_26146,N_24607,N_22208);
or U26147 (N_26147,N_23507,N_24837);
xor U26148 (N_26148,N_20090,N_20624);
xnor U26149 (N_26149,N_24187,N_20179);
nand U26150 (N_26150,N_21084,N_23032);
xor U26151 (N_26151,N_21640,N_24721);
or U26152 (N_26152,N_22373,N_21363);
xor U26153 (N_26153,N_24914,N_24672);
xor U26154 (N_26154,N_23084,N_20884);
or U26155 (N_26155,N_24977,N_24698);
xnor U26156 (N_26156,N_21976,N_24938);
nor U26157 (N_26157,N_21154,N_24225);
nand U26158 (N_26158,N_24542,N_23463);
and U26159 (N_26159,N_20667,N_24793);
nor U26160 (N_26160,N_24331,N_23932);
nor U26161 (N_26161,N_24107,N_23135);
nor U26162 (N_26162,N_23537,N_20307);
or U26163 (N_26163,N_23081,N_24948);
nand U26164 (N_26164,N_23580,N_24275);
nor U26165 (N_26165,N_20764,N_21104);
nor U26166 (N_26166,N_23899,N_24946);
xnor U26167 (N_26167,N_23203,N_23384);
nand U26168 (N_26168,N_22635,N_21310);
nor U26169 (N_26169,N_23606,N_23467);
or U26170 (N_26170,N_24800,N_22953);
xor U26171 (N_26171,N_24055,N_24068);
xnor U26172 (N_26172,N_20899,N_20821);
or U26173 (N_26173,N_23688,N_24276);
or U26174 (N_26174,N_20277,N_24197);
and U26175 (N_26175,N_21266,N_22500);
xnor U26176 (N_26176,N_21306,N_24515);
nand U26177 (N_26177,N_24020,N_23901);
or U26178 (N_26178,N_23239,N_23863);
xnor U26179 (N_26179,N_24372,N_22035);
xor U26180 (N_26180,N_21332,N_20948);
and U26181 (N_26181,N_22048,N_21339);
xor U26182 (N_26182,N_21196,N_20865);
nor U26183 (N_26183,N_20335,N_20411);
nand U26184 (N_26184,N_24505,N_22597);
or U26185 (N_26185,N_23155,N_22847);
nor U26186 (N_26186,N_21742,N_23332);
nand U26187 (N_26187,N_21796,N_24373);
nor U26188 (N_26188,N_23365,N_23468);
nor U26189 (N_26189,N_24813,N_22498);
nor U26190 (N_26190,N_21412,N_20679);
xnor U26191 (N_26191,N_23464,N_23252);
nor U26192 (N_26192,N_23313,N_20510);
or U26193 (N_26193,N_22089,N_20025);
nand U26194 (N_26194,N_20059,N_24796);
and U26195 (N_26195,N_24685,N_24358);
or U26196 (N_26196,N_22428,N_24526);
nand U26197 (N_26197,N_20588,N_20209);
nor U26198 (N_26198,N_21264,N_20616);
nor U26199 (N_26199,N_22985,N_20983);
or U26200 (N_26200,N_21870,N_24798);
nand U26201 (N_26201,N_24535,N_23055);
nor U26202 (N_26202,N_21346,N_20052);
nor U26203 (N_26203,N_20631,N_23303);
and U26204 (N_26204,N_20410,N_21969);
nand U26205 (N_26205,N_20495,N_22098);
or U26206 (N_26206,N_22697,N_20696);
and U26207 (N_26207,N_24623,N_23722);
and U26208 (N_26208,N_20168,N_20001);
nand U26209 (N_26209,N_22626,N_21288);
and U26210 (N_26210,N_21899,N_24140);
xor U26211 (N_26211,N_21261,N_23655);
nand U26212 (N_26212,N_23765,N_24102);
nand U26213 (N_26213,N_21800,N_20188);
nor U26214 (N_26214,N_23184,N_24081);
and U26215 (N_26215,N_20992,N_24113);
nor U26216 (N_26216,N_21528,N_24397);
nor U26217 (N_26217,N_22183,N_21836);
and U26218 (N_26218,N_20924,N_22012);
nand U26219 (N_26219,N_24618,N_24360);
and U26220 (N_26220,N_20280,N_21680);
nor U26221 (N_26221,N_24393,N_21872);
and U26222 (N_26222,N_20294,N_22754);
or U26223 (N_26223,N_22068,N_24428);
nand U26224 (N_26224,N_22417,N_24352);
or U26225 (N_26225,N_20484,N_21131);
nor U26226 (N_26226,N_23214,N_22892);
or U26227 (N_26227,N_22033,N_20183);
and U26228 (N_26228,N_20717,N_20471);
or U26229 (N_26229,N_24993,N_23659);
and U26230 (N_26230,N_23213,N_22535);
nand U26231 (N_26231,N_21111,N_23142);
nor U26232 (N_26232,N_20947,N_20709);
nor U26233 (N_26233,N_22416,N_23150);
and U26234 (N_26234,N_23937,N_21026);
xor U26235 (N_26235,N_20622,N_21299);
nand U26236 (N_26236,N_24468,N_20780);
nor U26237 (N_26237,N_20789,N_20311);
nor U26238 (N_26238,N_24775,N_21313);
xor U26239 (N_26239,N_23550,N_23632);
nor U26240 (N_26240,N_23770,N_24750);
or U26241 (N_26241,N_22178,N_20201);
or U26242 (N_26242,N_22037,N_23094);
or U26243 (N_26243,N_20597,N_23922);
nand U26244 (N_26244,N_21411,N_20776);
xor U26245 (N_26245,N_23867,N_24170);
nand U26246 (N_26246,N_20834,N_21157);
or U26247 (N_26247,N_24971,N_22496);
xnor U26248 (N_26248,N_23557,N_20488);
nor U26249 (N_26249,N_22729,N_24061);
xnor U26250 (N_26250,N_24620,N_21840);
xnor U26251 (N_26251,N_21107,N_20710);
xor U26252 (N_26252,N_23833,N_24480);
or U26253 (N_26253,N_24926,N_24010);
nand U26254 (N_26254,N_24674,N_23274);
nor U26255 (N_26255,N_21159,N_21744);
nand U26256 (N_26256,N_20266,N_23024);
xor U26257 (N_26257,N_24866,N_21645);
nor U26258 (N_26258,N_22069,N_23538);
and U26259 (N_26259,N_21514,N_21165);
and U26260 (N_26260,N_24355,N_21478);
or U26261 (N_26261,N_24367,N_24442);
xnor U26262 (N_26262,N_23848,N_21709);
or U26263 (N_26263,N_23095,N_23310);
and U26264 (N_26264,N_24363,N_22725);
xor U26265 (N_26265,N_22868,N_20744);
or U26266 (N_26266,N_24386,N_22834);
xnor U26267 (N_26267,N_22996,N_24499);
and U26268 (N_26268,N_23185,N_23196);
nor U26269 (N_26269,N_20316,N_22794);
nand U26270 (N_26270,N_24031,N_21891);
xor U26271 (N_26271,N_21174,N_22123);
xnor U26272 (N_26272,N_23044,N_24889);
or U26273 (N_26273,N_21505,N_23830);
nor U26274 (N_26274,N_22993,N_20345);
or U26275 (N_26275,N_20623,N_22239);
xnor U26276 (N_26276,N_21155,N_24251);
xor U26277 (N_26277,N_23284,N_20105);
xor U26278 (N_26278,N_20272,N_22942);
or U26279 (N_26279,N_22662,N_22716);
or U26280 (N_26280,N_24100,N_24736);
or U26281 (N_26281,N_22339,N_21568);
nand U26282 (N_26282,N_20991,N_20215);
and U26283 (N_26283,N_23318,N_20340);
and U26284 (N_26284,N_20468,N_22897);
nand U26285 (N_26285,N_21156,N_22943);
xnor U26286 (N_26286,N_20716,N_21515);
nand U26287 (N_26287,N_23827,N_22375);
and U26288 (N_26288,N_24763,N_20719);
and U26289 (N_26289,N_20759,N_23795);
or U26290 (N_26290,N_24882,N_20686);
or U26291 (N_26291,N_22081,N_20451);
nor U26292 (N_26292,N_21585,N_20055);
nor U26293 (N_26293,N_22827,N_22708);
nand U26294 (N_26294,N_22865,N_21536);
nor U26295 (N_26295,N_24173,N_24527);
or U26296 (N_26296,N_20753,N_22950);
nor U26297 (N_26297,N_22270,N_22013);
nor U26298 (N_26298,N_22615,N_20355);
or U26299 (N_26299,N_21981,N_20869);
and U26300 (N_26300,N_24941,N_20103);
nor U26301 (N_26301,N_20462,N_23205);
or U26302 (N_26302,N_20412,N_22429);
nand U26303 (N_26303,N_23536,N_23712);
and U26304 (N_26304,N_21115,N_22595);
nor U26305 (N_26305,N_20788,N_24483);
and U26306 (N_26306,N_23218,N_23246);
and U26307 (N_26307,N_20305,N_22396);
and U26308 (N_26308,N_21229,N_23009);
or U26309 (N_26309,N_23320,N_22808);
and U26310 (N_26310,N_22407,N_20704);
or U26311 (N_26311,N_23475,N_22426);
nand U26312 (N_26312,N_24119,N_22397);
or U26313 (N_26313,N_22336,N_23886);
xor U26314 (N_26314,N_22240,N_20442);
nor U26315 (N_26315,N_22668,N_22570);
nor U26316 (N_26316,N_23975,N_24288);
and U26317 (N_26317,N_22372,N_20943);
and U26318 (N_26318,N_20364,N_24722);
or U26319 (N_26319,N_20203,N_22766);
nor U26320 (N_26320,N_23637,N_24708);
and U26321 (N_26321,N_21438,N_20198);
or U26322 (N_26322,N_20020,N_20135);
nand U26323 (N_26323,N_21961,N_21148);
xnor U26324 (N_26324,N_20627,N_24087);
xor U26325 (N_26325,N_20800,N_24604);
xor U26326 (N_26326,N_23894,N_20033);
nor U26327 (N_26327,N_21049,N_23654);
and U26328 (N_26328,N_22512,N_24531);
nor U26329 (N_26329,N_22681,N_22361);
xor U26330 (N_26330,N_21083,N_20874);
and U26331 (N_26331,N_22743,N_20952);
or U26332 (N_26332,N_24742,N_20171);
nor U26333 (N_26333,N_20557,N_23545);
or U26334 (N_26334,N_24744,N_24963);
nand U26335 (N_26335,N_23696,N_23098);
and U26336 (N_26336,N_22526,N_24688);
nor U26337 (N_26337,N_24580,N_24019);
and U26338 (N_26338,N_22185,N_24966);
nand U26339 (N_26339,N_21338,N_22120);
nand U26340 (N_26340,N_20586,N_24902);
xor U26341 (N_26341,N_20056,N_20155);
nor U26342 (N_26342,N_20812,N_20559);
xor U26343 (N_26343,N_22533,N_23858);
xnor U26344 (N_26344,N_20121,N_23377);
and U26345 (N_26345,N_20116,N_23381);
nand U26346 (N_26346,N_24228,N_23198);
and U26347 (N_26347,N_21098,N_23479);
xor U26348 (N_26348,N_23459,N_23543);
nand U26349 (N_26349,N_24447,N_23235);
xor U26350 (N_26350,N_21661,N_24346);
and U26351 (N_26351,N_20086,N_21642);
xor U26352 (N_26352,N_21496,N_23939);
or U26353 (N_26353,N_21442,N_21716);
xnor U26354 (N_26354,N_22101,N_22162);
nor U26355 (N_26355,N_21721,N_21109);
and U26356 (N_26356,N_20132,N_23409);
or U26357 (N_26357,N_21755,N_20247);
xor U26358 (N_26358,N_22735,N_23674);
xor U26359 (N_26359,N_22168,N_23042);
nand U26360 (N_26360,N_23457,N_23121);
and U26361 (N_26361,N_20521,N_20010);
nand U26362 (N_26362,N_21793,N_21103);
nor U26363 (N_26363,N_20501,N_24142);
xnor U26364 (N_26364,N_24051,N_23617);
nand U26365 (N_26365,N_23046,N_24169);
and U26366 (N_26366,N_22746,N_23692);
or U26367 (N_26367,N_21428,N_21060);
nand U26368 (N_26368,N_24956,N_24154);
xnor U26369 (N_26369,N_20293,N_22018);
nor U26370 (N_26370,N_21888,N_21736);
nor U26371 (N_26371,N_23778,N_22648);
nand U26372 (N_26372,N_21036,N_20695);
or U26373 (N_26373,N_24463,N_22552);
nand U26374 (N_26374,N_24394,N_20094);
xor U26375 (N_26375,N_22015,N_24083);
xnor U26376 (N_26376,N_20192,N_22165);
xor U26377 (N_26377,N_21144,N_21785);
nor U26378 (N_26378,N_21005,N_22829);
xor U26379 (N_26379,N_20354,N_23731);
and U26380 (N_26380,N_20465,N_23586);
xnor U26381 (N_26381,N_22322,N_24414);
and U26382 (N_26382,N_24153,N_23872);
and U26383 (N_26383,N_20828,N_22059);
and U26384 (N_26384,N_21798,N_22984);
nand U26385 (N_26385,N_24765,N_21771);
and U26386 (N_26386,N_23256,N_23281);
or U26387 (N_26387,N_22362,N_23884);
and U26388 (N_26388,N_24724,N_24261);
nor U26389 (N_26389,N_20099,N_20549);
or U26390 (N_26390,N_24896,N_22445);
or U26391 (N_26391,N_20413,N_23423);
nor U26392 (N_26392,N_22315,N_24614);
nor U26393 (N_26393,N_23474,N_23882);
nand U26394 (N_26394,N_23337,N_23395);
and U26395 (N_26395,N_21570,N_24950);
nand U26396 (N_26396,N_22558,N_20114);
nand U26397 (N_26397,N_23123,N_21737);
nor U26398 (N_26398,N_24272,N_23910);
or U26399 (N_26399,N_22235,N_23499);
nand U26400 (N_26400,N_21809,N_22728);
and U26401 (N_26401,N_24440,N_21606);
or U26402 (N_26402,N_21436,N_21705);
xnor U26403 (N_26403,N_22879,N_24833);
nand U26404 (N_26404,N_22036,N_23039);
nand U26405 (N_26405,N_22828,N_24190);
xor U26406 (N_26406,N_23166,N_20450);
nand U26407 (N_26407,N_24664,N_21071);
or U26408 (N_26408,N_20406,N_23471);
nor U26409 (N_26409,N_21311,N_21467);
or U26410 (N_26410,N_23687,N_21684);
or U26411 (N_26411,N_24514,N_22857);
or U26412 (N_26412,N_21873,N_24298);
nand U26413 (N_26413,N_20886,N_20661);
or U26414 (N_26414,N_23358,N_23572);
xnor U26415 (N_26415,N_20785,N_24506);
or U26416 (N_26416,N_20694,N_23319);
nand U26417 (N_26417,N_24752,N_24134);
or U26418 (N_26418,N_21791,N_24621);
nand U26419 (N_26419,N_22968,N_23191);
and U26420 (N_26420,N_23236,N_21195);
xor U26421 (N_26421,N_21151,N_20259);
nand U26422 (N_26422,N_23483,N_22917);
nor U26423 (N_26423,N_21072,N_23789);
and U26424 (N_26424,N_23865,N_23920);
xnor U26425 (N_26425,N_20226,N_20041);
xor U26426 (N_26426,N_20937,N_20331);
xor U26427 (N_26427,N_20016,N_21168);
or U26428 (N_26428,N_21599,N_23645);
or U26429 (N_26429,N_23528,N_24208);
or U26430 (N_26430,N_23413,N_23418);
nor U26431 (N_26431,N_24379,N_24516);
nor U26432 (N_26432,N_24362,N_20748);
nor U26433 (N_26433,N_20072,N_20326);
nor U26434 (N_26434,N_24382,N_23546);
nand U26435 (N_26435,N_24511,N_22577);
nand U26436 (N_26436,N_20048,N_21760);
xor U26437 (N_26437,N_21095,N_24615);
xnor U26438 (N_26438,N_20533,N_22418);
nand U26439 (N_26439,N_20475,N_20165);
xnor U26440 (N_26440,N_22807,N_20554);
and U26441 (N_26441,N_21460,N_21485);
and U26442 (N_26442,N_22719,N_24395);
or U26443 (N_26443,N_24808,N_21419);
nor U26444 (N_26444,N_20034,N_20684);
and U26445 (N_26445,N_20487,N_24597);
or U26446 (N_26446,N_20592,N_22054);
xnor U26447 (N_26447,N_22916,N_24101);
xor U26448 (N_26448,N_24222,N_22190);
nand U26449 (N_26449,N_22765,N_21272);
xor U26450 (N_26450,N_20042,N_24050);
nand U26451 (N_26451,N_23963,N_23565);
xor U26452 (N_26452,N_24822,N_22323);
and U26453 (N_26453,N_23078,N_21375);
nand U26454 (N_26454,N_23831,N_21971);
or U26455 (N_26455,N_20083,N_21936);
xor U26456 (N_26456,N_20213,N_23211);
nor U26457 (N_26457,N_24928,N_22485);
and U26458 (N_26458,N_20082,N_21280);
nor U26459 (N_26459,N_21916,N_21817);
or U26460 (N_26460,N_21172,N_21550);
xnor U26461 (N_26461,N_22215,N_24497);
nand U26462 (N_26462,N_20063,N_20178);
nor U26463 (N_26463,N_20701,N_22370);
nor U26464 (N_26464,N_24587,N_21251);
nand U26465 (N_26465,N_20986,N_24630);
xnor U26466 (N_26466,N_22798,N_22520);
and U26467 (N_26467,N_23579,N_20749);
nand U26468 (N_26468,N_23670,N_23727);
or U26469 (N_26469,N_22638,N_24092);
or U26470 (N_26470,N_23071,N_21539);
nor U26471 (N_26471,N_23875,N_21584);
nand U26472 (N_26472,N_22186,N_24486);
nor U26473 (N_26473,N_24106,N_23989);
nand U26474 (N_26474,N_20423,N_23449);
or U26475 (N_26475,N_24999,N_23446);
nor U26476 (N_26476,N_21906,N_22933);
or U26477 (N_26477,N_24120,N_24577);
and U26478 (N_26478,N_23695,N_21651);
nand U26479 (N_26479,N_20127,N_24828);
and U26480 (N_26480,N_21855,N_21757);
or U26481 (N_26481,N_24840,N_22655);
or U26482 (N_26482,N_21193,N_23090);
and U26483 (N_26483,N_20249,N_24838);
nor U26484 (N_26484,N_24738,N_24458);
or U26485 (N_26485,N_20257,N_22778);
and U26486 (N_26486,N_21064,N_20445);
nand U26487 (N_26487,N_20467,N_23623);
nand U26488 (N_26488,N_24994,N_23639);
and U26489 (N_26489,N_20360,N_24135);
and U26490 (N_26490,N_24572,N_21538);
or U26491 (N_26491,N_20417,N_22179);
nor U26492 (N_26492,N_21471,N_22042);
xnor U26493 (N_26493,N_24961,N_23285);
nand U26494 (N_26494,N_23091,N_20596);
and U26495 (N_26495,N_21634,N_23972);
and U26496 (N_26496,N_20482,N_22538);
and U26497 (N_26497,N_24627,N_24271);
xor U26498 (N_26498,N_20109,N_22660);
and U26499 (N_26499,N_24681,N_22380);
nand U26500 (N_26500,N_21622,N_21833);
and U26501 (N_26501,N_22699,N_23724);
and U26502 (N_26502,N_20133,N_23956);
and U26503 (N_26503,N_23642,N_20009);
or U26504 (N_26504,N_22293,N_21641);
or U26505 (N_26505,N_20536,N_24568);
nand U26506 (N_26506,N_20514,N_24293);
and U26507 (N_26507,N_20220,N_20676);
nor U26508 (N_26508,N_23748,N_24498);
nor U26509 (N_26509,N_23342,N_24820);
nand U26510 (N_26510,N_24284,N_20767);
xnor U26511 (N_26511,N_23051,N_24494);
and U26512 (N_26512,N_22657,N_23594);
and U26513 (N_26513,N_23604,N_22105);
xor U26514 (N_26514,N_23631,N_21498);
and U26515 (N_26515,N_20235,N_20344);
or U26516 (N_26516,N_20386,N_23222);
and U26517 (N_26517,N_23908,N_22307);
nand U26518 (N_26518,N_24229,N_20866);
and U26519 (N_26519,N_23958,N_22565);
and U26520 (N_26520,N_20466,N_24541);
or U26521 (N_26521,N_23680,N_24481);
nand U26522 (N_26522,N_23314,N_21421);
or U26523 (N_26523,N_20003,N_20200);
or U26524 (N_26524,N_22176,N_23622);
nand U26525 (N_26525,N_24934,N_22934);
and U26526 (N_26526,N_21446,N_23277);
nand U26527 (N_26527,N_24409,N_20900);
nor U26528 (N_26528,N_21724,N_24145);
or U26529 (N_26529,N_24629,N_21335);
and U26530 (N_26530,N_24908,N_23618);
nor U26531 (N_26531,N_24898,N_21659);
nor U26532 (N_26532,N_24936,N_20689);
xor U26533 (N_26533,N_21087,N_24219);
nor U26534 (N_26534,N_22983,N_23012);
or U26535 (N_26535,N_24205,N_22995);
nor U26536 (N_26536,N_21876,N_24445);
nand U26537 (N_26537,N_22672,N_21499);
xnor U26538 (N_26538,N_20231,N_22956);
nand U26539 (N_26539,N_22871,N_22830);
xor U26540 (N_26540,N_20977,N_23810);
and U26541 (N_26541,N_24589,N_20833);
and U26542 (N_26542,N_23460,N_22973);
and U26543 (N_26543,N_22050,N_21232);
nor U26544 (N_26544,N_23153,N_23025);
nand U26545 (N_26545,N_24270,N_21469);
nand U26546 (N_26546,N_20715,N_24585);
xor U26547 (N_26547,N_24146,N_23286);
nor U26548 (N_26548,N_22691,N_21409);
nor U26549 (N_26549,N_24239,N_21021);
or U26550 (N_26550,N_23489,N_23233);
nor U26551 (N_26551,N_21806,N_23158);
or U26552 (N_26552,N_21741,N_23883);
nand U26553 (N_26553,N_24323,N_21182);
nand U26554 (N_26554,N_21607,N_23215);
or U26555 (N_26555,N_20595,N_24257);
nor U26556 (N_26556,N_20187,N_21385);
nand U26557 (N_26557,N_21250,N_24044);
nand U26558 (N_26558,N_23636,N_22029);
or U26559 (N_26559,N_20244,N_21362);
nand U26560 (N_26560,N_22764,N_24224);
nand U26561 (N_26561,N_23907,N_21149);
or U26562 (N_26562,N_22124,N_20476);
and U26563 (N_26563,N_23924,N_23591);
nor U26564 (N_26564,N_24178,N_21803);
nand U26565 (N_26565,N_20295,N_20357);
and U26566 (N_26566,N_23139,N_21358);
and U26567 (N_26567,N_21347,N_21450);
nand U26568 (N_26568,N_20979,N_20691);
xor U26569 (N_26569,N_21650,N_24233);
nor U26570 (N_26570,N_24416,N_23734);
nand U26571 (N_26571,N_23003,N_21993);
or U26572 (N_26572,N_22383,N_20154);
or U26573 (N_26573,N_22172,N_22559);
or U26574 (N_26574,N_21775,N_23392);
and U26575 (N_26575,N_21348,N_23451);
xnor U26576 (N_26576,N_21695,N_23498);
nand U26577 (N_26577,N_22351,N_21216);
and U26578 (N_26578,N_20993,N_22936);
nor U26579 (N_26579,N_21703,N_23866);
nand U26580 (N_26580,N_21834,N_21236);
or U26581 (N_26581,N_21889,N_20724);
or U26582 (N_26582,N_20893,N_22918);
and U26583 (N_26583,N_20390,N_22587);
nor U26584 (N_26584,N_24693,N_22877);
and U26585 (N_26585,N_21813,N_24227);
nor U26586 (N_26586,N_22348,N_22244);
xor U26587 (N_26587,N_21778,N_24149);
nand U26588 (N_26588,N_23667,N_20046);
and U26589 (N_26589,N_21189,N_21162);
xor U26590 (N_26590,N_23484,N_22444);
xnor U26591 (N_26591,N_23368,N_20248);
nand U26592 (N_26592,N_22357,N_22456);
nor U26593 (N_26593,N_23714,N_22641);
xnor U26594 (N_26594,N_24285,N_24879);
nand U26595 (N_26595,N_21625,N_22118);
and U26596 (N_26596,N_21203,N_21199);
nand U26597 (N_26597,N_21210,N_20161);
and U26598 (N_26598,N_20963,N_21852);
or U26599 (N_26599,N_21549,N_20848);
xor U26600 (N_26600,N_22073,N_22224);
xnor U26601 (N_26601,N_23354,N_21751);
or U26602 (N_26602,N_23080,N_22236);
xor U26603 (N_26603,N_20882,N_21907);
nand U26604 (N_26604,N_20600,N_21974);
and U26605 (N_26605,N_21102,N_21129);
nand U26606 (N_26606,N_24371,N_20392);
nor U26607 (N_26607,N_22356,N_22313);
nand U26608 (N_26608,N_22650,N_20649);
or U26609 (N_26609,N_21558,N_20850);
nand U26610 (N_26610,N_24786,N_22902);
nor U26611 (N_26611,N_20194,N_23817);
and U26612 (N_26612,N_24489,N_24103);
and U26613 (N_26613,N_22502,N_21121);
xor U26614 (N_26614,N_21133,N_23389);
nor U26615 (N_26615,N_23023,N_23240);
xnor U26616 (N_26616,N_24280,N_23812);
and U26617 (N_26617,N_24057,N_20427);
nand U26618 (N_26618,N_23541,N_21731);
xor U26619 (N_26619,N_20096,N_22324);
xnor U26620 (N_26620,N_22913,N_20242);
xnor U26621 (N_26621,N_24450,N_21965);
and U26622 (N_26622,N_21930,N_22747);
and U26623 (N_26623,N_24384,N_23045);
or U26624 (N_26624,N_22970,N_24304);
and U26625 (N_26625,N_21902,N_24862);
nand U26626 (N_26626,N_24252,N_21343);
or U26627 (N_26627,N_20459,N_24091);
or U26628 (N_26628,N_24562,N_20903);
and U26629 (N_26629,N_23302,N_23682);
nor U26630 (N_26630,N_21023,N_20143);
and U26631 (N_26631,N_20017,N_23194);
and U26632 (N_26632,N_24466,N_21086);
nor U26633 (N_26633,N_20648,N_21276);
and U26634 (N_26634,N_21295,N_23569);
xnor U26635 (N_26635,N_21637,N_24551);
xor U26636 (N_26636,N_22806,N_24406);
or U26637 (N_26637,N_22634,N_22079);
xnor U26638 (N_26638,N_20054,N_20013);
nor U26639 (N_26639,N_24052,N_21919);
nor U26640 (N_26640,N_23747,N_21997);
nor U26641 (N_26641,N_22720,N_22466);
xor U26642 (N_26642,N_24968,N_24341);
nand U26643 (N_26643,N_22853,N_20618);
or U26644 (N_26644,N_21512,N_20403);
nor U26645 (N_26645,N_20473,N_20742);
xnor U26646 (N_26646,N_23370,N_23797);
nand U26647 (N_26647,N_24297,N_20811);
and U26648 (N_26648,N_23590,N_24965);
nor U26649 (N_26649,N_21754,N_21372);
nor U26650 (N_26650,N_23131,N_23893);
or U26651 (N_26651,N_23520,N_20555);
and U26652 (N_26652,N_20396,N_21449);
xnor U26653 (N_26653,N_21344,N_21949);
and U26654 (N_26654,N_21764,N_20140);
nand U26655 (N_26655,N_23691,N_20184);
nand U26656 (N_26656,N_24086,N_22888);
nor U26657 (N_26657,N_20558,N_24354);
xor U26658 (N_26658,N_20944,N_24815);
or U26659 (N_26659,N_20864,N_21747);
xor U26660 (N_26660,N_23981,N_20276);
nand U26661 (N_26661,N_23321,N_20158);
nor U26662 (N_26662,N_20614,N_20675);
nand U26663 (N_26663,N_24639,N_24588);
nor U26664 (N_26664,N_23581,N_22154);
nor U26665 (N_26665,N_24566,N_21140);
and U26666 (N_26666,N_24777,N_20489);
or U26667 (N_26667,N_24953,N_20164);
or U26668 (N_26668,N_20481,N_22349);
nand U26669 (N_26669,N_20522,N_20478);
or U26670 (N_26670,N_21369,N_22435);
xnor U26671 (N_26671,N_22371,N_20824);
nor U26672 (N_26672,N_22038,N_22233);
and U26673 (N_26673,N_20402,N_23267);
nor U26674 (N_26674,N_24014,N_24451);
or U26675 (N_26675,N_21789,N_22204);
nor U26676 (N_26676,N_22817,N_20714);
and U26677 (N_26677,N_23941,N_20859);
nand U26678 (N_26678,N_21091,N_23334);
and U26679 (N_26679,N_21336,N_21656);
nand U26680 (N_26680,N_20393,N_20329);
xnor U26681 (N_26681,N_23815,N_23524);
nor U26682 (N_26682,N_20144,N_23226);
and U26683 (N_26683,N_23596,N_21050);
and U26684 (N_26684,N_21164,N_24433);
nand U26685 (N_26685,N_22182,N_23626);
xnor U26686 (N_26686,N_24012,N_24124);
nor U26687 (N_26687,N_20398,N_20585);
nor U26688 (N_26688,N_24449,N_20251);
nor U26689 (N_26689,N_24628,N_23832);
xor U26690 (N_26690,N_21749,N_22816);
and U26691 (N_26691,N_24903,N_23583);
nor U26692 (N_26692,N_22219,N_23266);
nor U26693 (N_26693,N_20985,N_24807);
or U26694 (N_26694,N_23809,N_21294);
nand U26695 (N_26695,N_21387,N_20581);
nor U26696 (N_26696,N_23729,N_22698);
and U26697 (N_26697,N_20577,N_23088);
nor U26698 (N_26698,N_24518,N_24308);
and U26699 (N_26699,N_24643,N_21031);
nand U26700 (N_26700,N_20268,N_22761);
xor U26701 (N_26701,N_20919,N_22207);
and U26702 (N_26702,N_23701,N_23577);
nand U26703 (N_26703,N_24047,N_21679);
nand U26704 (N_26704,N_24008,N_24133);
and U26705 (N_26705,N_24063,N_22297);
or U26706 (N_26706,N_23344,N_20285);
nand U26707 (N_26707,N_21608,N_20915);
nor U26708 (N_26708,N_21900,N_23681);
and U26709 (N_26709,N_20936,N_23988);
nand U26710 (N_26710,N_22438,N_23439);
and U26711 (N_26711,N_24265,N_23740);
nor U26712 (N_26712,N_23609,N_21839);
nand U26713 (N_26713,N_20797,N_23838);
xnor U26714 (N_26714,N_21225,N_22260);
nand U26715 (N_26715,N_20813,N_23718);
xnor U26716 (N_26716,N_23857,N_22072);
xnor U26717 (N_26717,N_23190,N_21763);
nor U26718 (N_26718,N_23800,N_22318);
nor U26719 (N_26719,N_20682,N_20177);
or U26720 (N_26720,N_21719,N_22998);
xnor U26721 (N_26721,N_22919,N_22944);
xnor U26722 (N_26722,N_23168,N_21233);
nand U26723 (N_26723,N_24236,N_22150);
and U26724 (N_26724,N_23690,N_22129);
nand U26725 (N_26725,N_22278,N_24835);
or U26726 (N_26726,N_20240,N_21886);
xnor U26727 (N_26727,N_20026,N_23726);
and U26728 (N_26728,N_20439,N_23387);
or U26729 (N_26729,N_20838,N_22516);
and U26730 (N_26730,N_21374,N_20377);
or U26731 (N_26731,N_20652,N_22633);
nor U26732 (N_26732,N_22813,N_24899);
and U26733 (N_26733,N_21726,N_20523);
nor U26734 (N_26734,N_23466,N_22196);
or U26735 (N_26735,N_21692,N_23366);
and U26736 (N_26736,N_23599,N_23207);
xor U26737 (N_26737,N_24536,N_24829);
nand U26738 (N_26738,N_21027,N_20539);
xor U26739 (N_26739,N_22742,N_23909);
and U26740 (N_26740,N_22540,N_21008);
nand U26741 (N_26741,N_22826,N_22799);
or U26742 (N_26742,N_24415,N_22521);
nand U26743 (N_26743,N_21108,N_21516);
or U26744 (N_26744,N_22267,N_22273);
xor U26745 (N_26745,N_24706,N_20630);
nand U26746 (N_26746,N_24544,N_22047);
nand U26747 (N_26747,N_23781,N_22462);
nor U26748 (N_26748,N_21860,N_24123);
nor U26749 (N_26749,N_21797,N_20064);
xor U26750 (N_26750,N_24925,N_24917);
and U26751 (N_26751,N_21461,N_24356);
and U26752 (N_26752,N_21653,N_23553);
and U26753 (N_26753,N_21799,N_23570);
nor U26754 (N_26754,N_22921,N_23269);
nand U26755 (N_26755,N_22020,N_24983);
xnor U26756 (N_26756,N_21954,N_21052);
xor U26757 (N_26757,N_21016,N_21832);
xor U26758 (N_26758,N_23947,N_21897);
xnor U26759 (N_26759,N_20093,N_20867);
and U26760 (N_26760,N_22175,N_24731);
nand U26761 (N_26761,N_21871,N_22802);
nor U26762 (N_26762,N_20960,N_21128);
nand U26763 (N_26763,N_22749,N_21896);
nand U26764 (N_26764,N_24780,N_22052);
nor U26765 (N_26765,N_20642,N_20830);
xnor U26766 (N_26766,N_24992,N_24015);
nand U26767 (N_26767,N_21998,N_20298);
xor U26768 (N_26768,N_24254,N_23814);
and U26769 (N_26769,N_21784,N_24690);
xor U26770 (N_26770,N_23911,N_20043);
nor U26771 (N_26771,N_24860,N_22492);
and U26772 (N_26772,N_20733,N_20861);
or U26773 (N_26773,N_20890,N_24540);
or U26774 (N_26774,N_21681,N_21905);
or U26775 (N_26775,N_20809,N_22642);
or U26776 (N_26776,N_22980,N_23955);
or U26777 (N_26777,N_23749,N_24115);
and U26778 (N_26778,N_22478,N_20550);
nand U26779 (N_26779,N_21018,N_24850);
and U26780 (N_26780,N_24919,N_21153);
and U26781 (N_26781,N_21053,N_20542);
or U26782 (N_26782,N_22189,N_20707);
or U26783 (N_26783,N_21209,N_20609);
nor U26784 (N_26784,N_21966,N_22741);
and U26785 (N_26785,N_20022,N_20498);
nor U26786 (N_26786,N_20513,N_21202);
or U26787 (N_26787,N_20907,N_22364);
and U26788 (N_26788,N_21235,N_20852);
and U26789 (N_26789,N_23929,N_23341);
and U26790 (N_26790,N_24118,N_23241);
xnor U26791 (N_26791,N_24755,N_24622);
xnor U26792 (N_26792,N_22890,N_20552);
or U26793 (N_26793,N_20935,N_21922);
nand U26794 (N_26794,N_21994,N_20480);
xnor U26795 (N_26795,N_24781,N_22967);
nor U26796 (N_26796,N_20065,N_21867);
and U26797 (N_26797,N_22199,N_23529);
or U26798 (N_26798,N_20362,N_22653);
nand U26799 (N_26799,N_20472,N_22093);
xnor U26800 (N_26800,N_21138,N_23290);
and U26801 (N_26801,N_24776,N_24116);
xor U26802 (N_26802,N_22689,N_20920);
and U26803 (N_26803,N_23132,N_23717);
xnor U26804 (N_26804,N_22536,N_21456);
xor U26805 (N_26805,N_24425,N_22125);
nor U26806 (N_26806,N_23716,N_21491);
and U26807 (N_26807,N_24924,N_20389);
nor U26808 (N_26808,N_20965,N_23008);
and U26809 (N_26809,N_20186,N_23532);
and U26810 (N_26810,N_23019,N_21814);
or U26811 (N_26811,N_22222,N_22614);
and U26812 (N_26812,N_21756,N_22639);
xor U26813 (N_26813,N_24230,N_21017);
and U26814 (N_26814,N_22110,N_24441);
xor U26815 (N_26815,N_23052,N_21117);
or U26816 (N_26816,N_22795,N_21497);
nand U26817 (N_26817,N_20342,N_21548);
xor U26818 (N_26818,N_22283,N_24462);
and U26819 (N_26819,N_24377,N_21169);
nor U26820 (N_26820,N_20731,N_21924);
nor U26821 (N_26821,N_23564,N_24085);
or U26822 (N_26822,N_23794,N_24076);
and U26823 (N_26823,N_24338,N_23556);
nand U26824 (N_26824,N_21523,N_24870);
or U26825 (N_26825,N_21000,N_21429);
or U26826 (N_26826,N_23903,N_23773);
or U26827 (N_26827,N_23470,N_21207);
xor U26828 (N_26828,N_24878,N_21546);
nor U26829 (N_26829,N_23242,N_20084);
nor U26830 (N_26830,N_23931,N_24151);
and U26831 (N_26831,N_23826,N_21772);
and U26832 (N_26832,N_21787,N_22019);
nor U26833 (N_26833,N_21879,N_24695);
nand U26834 (N_26834,N_21481,N_20871);
and U26835 (N_26835,N_22545,N_21794);
xnor U26836 (N_26836,N_24189,N_22524);
nor U26837 (N_26837,N_22522,N_22319);
and U26838 (N_26838,N_22200,N_23151);
nand U26839 (N_26839,N_22350,N_20181);
nand U26840 (N_26840,N_21715,N_23562);
and U26841 (N_26841,N_21682,N_24099);
or U26842 (N_26842,N_22406,N_24705);
nand U26843 (N_26843,N_20762,N_22632);
nor U26844 (N_26844,N_23415,N_20655);
nand U26845 (N_26845,N_24105,N_23684);
or U26846 (N_26846,N_21773,N_21530);
and U26847 (N_26847,N_20414,N_22122);
or U26848 (N_26848,N_23234,N_21356);
xnor U26849 (N_26849,N_23554,N_20666);
and U26850 (N_26850,N_23685,N_21753);
nor U26851 (N_26851,N_23322,N_21662);
and U26852 (N_26852,N_23380,N_21917);
xor U26853 (N_26853,N_24753,N_24412);
and U26854 (N_26854,N_23075,N_21802);
nand U26855 (N_26855,N_20548,N_20593);
nor U26856 (N_26856,N_23799,N_23496);
or U26857 (N_26857,N_21765,N_20892);
and U26858 (N_26858,N_20591,N_23007);
xnor U26859 (N_26859,N_20769,N_23348);
nand U26860 (N_26860,N_21477,N_23776);
nor U26861 (N_26861,N_23936,N_22976);
nand U26862 (N_26862,N_22454,N_23066);
nor U26863 (N_26863,N_21725,N_24212);
and U26864 (N_26864,N_20547,N_24876);
or U26865 (N_26865,N_21063,N_21720);
xnor U26866 (N_26866,N_20912,N_20540);
nor U26867 (N_26867,N_21317,N_23349);
and U26868 (N_26868,N_23791,N_22820);
and U26869 (N_26869,N_20810,N_22286);
xnor U26870 (N_26870,N_23065,N_24524);
xor U26871 (N_26871,N_22458,N_22335);
xor U26872 (N_26872,N_21090,N_20508);
nand U26873 (N_26873,N_24344,N_23450);
xor U26874 (N_26874,N_22547,N_22161);
nor U26875 (N_26875,N_23116,N_23708);
and U26876 (N_26876,N_21824,N_24904);
nor U26877 (N_26877,N_21502,N_23085);
or U26878 (N_26878,N_23821,N_24040);
nand U26879 (N_26879,N_22508,N_24129);
xor U26880 (N_26880,N_23420,N_22678);
xnor U26881 (N_26881,N_24350,N_24666);
nand U26882 (N_26882,N_24435,N_22151);
nand U26883 (N_26883,N_21904,N_22202);
nor U26884 (N_26884,N_24836,N_24378);
or U26885 (N_26885,N_23157,N_21632);
and U26886 (N_26886,N_24268,N_24567);
or U26887 (N_26887,N_21025,N_22248);
nand U26888 (N_26888,N_22494,N_20212);
nand U26889 (N_26889,N_21315,N_22422);
nor U26890 (N_26890,N_22982,N_21287);
nor U26891 (N_26891,N_22398,N_21178);
and U26892 (N_26892,N_22177,N_22409);
nand U26893 (N_26893,N_21727,N_21527);
or U26894 (N_26894,N_20632,N_22753);
nand U26895 (N_26895,N_24582,N_20849);
and U26896 (N_26896,N_22544,N_20725);
nor U26897 (N_26897,N_24823,N_20339);
or U26898 (N_26898,N_23410,N_24605);
and U26899 (N_26899,N_23197,N_23689);
xnor U26900 (N_26900,N_23101,N_21390);
or U26901 (N_26901,N_23406,N_23488);
xor U26902 (N_26902,N_24347,N_24754);
and U26903 (N_26903,N_24517,N_20621);
and U26904 (N_26904,N_20775,N_22831);
xnor U26905 (N_26905,N_23363,N_22066);
or U26906 (N_26906,N_22989,N_24818);
and U26907 (N_26907,N_23469,N_23634);
or U26908 (N_26908,N_23753,N_24141);
or U26909 (N_26909,N_22878,N_24940);
nor U26910 (N_26910,N_24036,N_20674);
xor U26911 (N_26911,N_21224,N_20263);
nor U26912 (N_26912,N_24594,N_20424);
or U26913 (N_26913,N_21987,N_23699);
or U26914 (N_26914,N_20889,N_21472);
and U26915 (N_26915,N_22563,N_21577);
nand U26916 (N_26916,N_21480,N_21434);
and U26917 (N_26917,N_24117,N_24900);
and U26918 (N_26918,N_23870,N_24774);
nor U26919 (N_26919,N_24570,N_24682);
nand U26920 (N_26920,N_21968,N_23782);
and U26921 (N_26921,N_22131,N_22949);
and U26922 (N_26922,N_23485,N_23224);
nor U26923 (N_26923,N_21267,N_22666);
nand U26924 (N_26924,N_23715,N_20881);
and U26925 (N_26925,N_20755,N_21125);
nand U26926 (N_26926,N_22281,N_24108);
nand U26927 (N_26927,N_20286,N_21081);
and U26928 (N_26928,N_24559,N_20483);
and U26929 (N_26929,N_22848,N_22360);
xnor U26930 (N_26930,N_24857,N_20646);
and U26931 (N_26931,N_22616,N_22659);
xor U26932 (N_26932,N_22796,N_22629);
or U26933 (N_26933,N_21683,N_21509);
and U26934 (N_26934,N_20008,N_24104);
xor U26935 (N_26935,N_21638,N_21418);
nor U26936 (N_26936,N_22006,N_21488);
xor U26937 (N_26937,N_24571,N_24500);
and U26938 (N_26938,N_24801,N_21985);
and U26939 (N_26939,N_21222,N_21325);
nand U26940 (N_26940,N_20490,N_20668);
xnor U26941 (N_26941,N_20425,N_21394);
nor U26942 (N_26942,N_21435,N_23200);
nor U26943 (N_26943,N_24636,N_20218);
xor U26944 (N_26944,N_22515,N_23130);
or U26945 (N_26945,N_23001,N_23864);
and U26946 (N_26946,N_22550,N_20573);
nor U26947 (N_26947,N_22412,N_23879);
and U26948 (N_26948,N_23860,N_20071);
nand U26949 (N_26949,N_20546,N_20129);
nand U26950 (N_26950,N_21285,N_20846);
nor U26951 (N_26951,N_22690,N_23852);
nand U26952 (N_26952,N_21918,N_21708);
and U26953 (N_26953,N_20656,N_20525);
nand U26954 (N_26954,N_20921,N_21454);
and U26955 (N_26955,N_21437,N_21319);
nand U26956 (N_26956,N_20243,N_22119);
or U26957 (N_26957,N_24676,N_22882);
and U26958 (N_26958,N_24510,N_22201);
or U26959 (N_26959,N_24785,N_24502);
and U26960 (N_26960,N_24320,N_23885);
and U26961 (N_26961,N_22247,N_24891);
and U26962 (N_26962,N_24711,N_23408);
nor U26963 (N_26963,N_21610,N_24385);
nand U26964 (N_26964,N_20594,N_22869);
nand U26965 (N_26965,N_22994,N_22529);
or U26966 (N_26966,N_22695,N_22301);
nand U26967 (N_26967,N_23223,N_22306);
nor U26968 (N_26968,N_22317,N_20587);
nand U26969 (N_26969,N_20790,N_24380);
nor U26970 (N_26970,N_22060,N_20770);
nand U26971 (N_26971,N_23227,N_24554);
and U26972 (N_26972,N_20654,N_24846);
and U26973 (N_26973,N_21636,N_20460);
and U26974 (N_26974,N_21147,N_20932);
and U26975 (N_26975,N_21667,N_20365);
or U26976 (N_26976,N_23340,N_24370);
or U26977 (N_26977,N_24064,N_24670);
nor U26978 (N_26978,N_23343,N_24578);
nor U26979 (N_26979,N_23856,N_20110);
and U26980 (N_26980,N_20563,N_24255);
and U26981 (N_26981,N_23244,N_24053);
and U26982 (N_26982,N_24633,N_23751);
nor U26983 (N_26983,N_22601,N_21445);
nand U26984 (N_26984,N_22523,N_22071);
or U26985 (N_26985,N_24192,N_21455);
and U26986 (N_26986,N_24243,N_22886);
and U26987 (N_26987,N_24556,N_24696);
nor U26988 (N_26988,N_21912,N_21717);
or U26989 (N_26989,N_21600,N_21580);
xnor U26990 (N_26990,N_21177,N_24181);
and U26991 (N_26991,N_23732,N_20264);
xor U26992 (N_26992,N_24213,N_22194);
and U26993 (N_26993,N_21944,N_23994);
xor U26994 (N_26994,N_20279,N_24072);
nor U26995 (N_26995,N_20107,N_20794);
xnor U26996 (N_26996,N_21988,N_23853);
xor U26997 (N_26997,N_21841,N_23880);
xnor U26998 (N_26998,N_21583,N_24789);
or U26999 (N_26999,N_23822,N_22193);
and U27000 (N_27000,N_20031,N_22758);
or U27001 (N_27001,N_22625,N_24171);
nand U27002 (N_27002,N_24729,N_21895);
nand U27003 (N_27003,N_21273,N_22132);
nor U27004 (N_27004,N_22620,N_22714);
and U27005 (N_27005,N_20130,N_24616);
nand U27006 (N_27006,N_21533,N_20841);
and U27007 (N_27007,N_22596,N_24034);
or U27008 (N_27008,N_24496,N_22762);
xor U27009 (N_27009,N_24895,N_22063);
nand U27010 (N_27010,N_24175,N_23416);
or U27011 (N_27011,N_23273,N_24402);
and U27012 (N_27012,N_20608,N_23407);
nand U27013 (N_27013,N_22051,N_21972);
or U27014 (N_27014,N_20933,N_21946);
and U27015 (N_27015,N_24644,N_20492);
and U27016 (N_27016,N_20418,N_24273);
xor U27017 (N_27017,N_24575,N_22001);
xor U27018 (N_27018,N_21304,N_21795);
xnor U27019 (N_27019,N_21001,N_20825);
xor U27020 (N_27020,N_24525,N_24188);
nor U27021 (N_27021,N_22130,N_24157);
nor U27022 (N_27022,N_24016,N_24098);
nand U27023 (N_27023,N_22914,N_21519);
and U27024 (N_27024,N_23694,N_20997);
nor U27025 (N_27025,N_21092,N_20101);
or U27026 (N_27026,N_21241,N_20804);
and U27027 (N_27027,N_21615,N_22509);
and U27028 (N_27028,N_20639,N_20665);
nand U27029 (N_27029,N_21035,N_21351);
nor U27030 (N_27030,N_20987,N_20080);
nor U27031 (N_27031,N_20862,N_24601);
or U27032 (N_27032,N_20966,N_22506);
nand U27033 (N_27033,N_21603,N_20615);
and U27034 (N_27034,N_22556,N_22358);
and U27035 (N_27035,N_22441,N_20229);
or U27036 (N_27036,N_22895,N_24951);
or U27037 (N_27037,N_21044,N_20190);
xor U27038 (N_27038,N_20453,N_23525);
and U27039 (N_27039,N_23454,N_21056);
nand U27040 (N_27040,N_24312,N_20941);
nand U27041 (N_27041,N_23746,N_22004);
nor U27042 (N_27042,N_23710,N_22234);
nand U27043 (N_27043,N_24651,N_20027);
xnor U27044 (N_27044,N_23869,N_22437);
and U27045 (N_27045,N_21495,N_21078);
xnor U27046 (N_27046,N_20146,N_23043);
and U27047 (N_27047,N_22578,N_22474);
nor U27048 (N_27048,N_21984,N_24958);
xor U27049 (N_27049,N_22292,N_23047);
xor U27050 (N_27050,N_23104,N_24066);
nand U27051 (N_27051,N_20374,N_22673);
or U27052 (N_27052,N_20352,N_22413);
nand U27053 (N_27053,N_20644,N_21846);
nand U27054 (N_27054,N_20325,N_23414);
and U27055 (N_27055,N_21557,N_20207);
nor U27056 (N_27056,N_23243,N_20988);
or U27057 (N_27057,N_22885,N_22062);
or U27058 (N_27058,N_24029,N_23987);
xor U27059 (N_27059,N_21074,N_22034);
xnor U27060 (N_27060,N_24405,N_21009);
nor U27061 (N_27061,N_23575,N_20628);
xnor U27062 (N_27062,N_21831,N_23099);
xnor U27063 (N_27063,N_21365,N_22661);
and U27064 (N_27064,N_24470,N_23181);
or U27065 (N_27065,N_20868,N_22253);
xor U27066 (N_27066,N_22991,N_24329);
xnor U27067 (N_27067,N_24488,N_24277);
nor U27068 (N_27068,N_24883,N_21381);
nand U27069 (N_27069,N_21462,N_20973);
nand U27070 (N_27070,N_21179,N_22127);
and U27071 (N_27071,N_22030,N_22663);
nor U27072 (N_27072,N_20149,N_23114);
nand U27073 (N_27073,N_22395,N_21247);
and U27074 (N_27074,N_20807,N_22277);
nand U27075 (N_27075,N_22473,N_22061);
xor U27076 (N_27076,N_24299,N_22722);
or U27077 (N_27077,N_20061,N_20115);
and U27078 (N_27078,N_23452,N_23301);
or U27079 (N_27079,N_24569,N_21995);
and U27080 (N_27080,N_20349,N_20363);
nand U27081 (N_27081,N_20024,N_24240);
nor U27082 (N_27082,N_24282,N_21526);
or U27083 (N_27083,N_20740,N_24204);
and U27084 (N_27084,N_24553,N_22436);
xor U27085 (N_27085,N_23518,N_23385);
xnor U27086 (N_27086,N_20091,N_23059);
xnor U27087 (N_27087,N_22499,N_23898);
and U27088 (N_27088,N_23742,N_21866);
nor U27089 (N_27089,N_23289,N_23589);
and U27090 (N_27090,N_22039,N_22312);
or U27091 (N_27091,N_23656,N_23905);
xnor U27092 (N_27092,N_21935,N_23948);
xnor U27093 (N_27093,N_22148,N_22791);
xnor U27094 (N_27094,N_22477,N_21041);
and U27095 (N_27095,N_20000,N_22872);
nand U27096 (N_27096,N_21618,N_20436);
nor U27097 (N_27097,N_24247,N_23307);
or U27098 (N_27098,N_20635,N_24114);
and U27099 (N_27099,N_23124,N_23375);
nand U27100 (N_27100,N_23329,N_23593);
xnor U27101 (N_27101,N_21780,N_21039);
and U27102 (N_27102,N_23394,N_20590);
nor U27103 (N_27103,N_24767,N_20926);
xor U27104 (N_27104,N_21423,N_24318);
or U27105 (N_27105,N_24911,N_21779);
and U27106 (N_27106,N_23112,N_24667);
xor U27107 (N_27107,N_23216,N_22987);
nand U27108 (N_27108,N_21696,N_24513);
or U27109 (N_27109,N_22822,N_20045);
nor U27110 (N_27110,N_23890,N_22864);
xor U27111 (N_27111,N_20972,N_21657);
nor U27112 (N_27112,N_23082,N_21426);
and U27113 (N_27113,N_23350,N_24719);
nor U27114 (N_27114,N_22760,N_22852);
nand U27115 (N_27115,N_22528,N_22213);
or U27116 (N_27116,N_23183,N_21909);
xnor U27117 (N_27117,N_24933,N_23757);
or U27118 (N_27118,N_20737,N_20214);
nor U27119 (N_27119,N_23097,N_22733);
or U27120 (N_27120,N_21808,N_24532);
and U27121 (N_27121,N_23397,N_23658);
xnor U27122 (N_27122,N_23304,N_20317);
xor U27123 (N_27123,N_20990,N_23175);
or U27124 (N_27124,N_22187,N_24726);
or U27125 (N_27125,N_23666,N_24491);
nor U27126 (N_27126,N_20156,N_20252);
nand U27127 (N_27127,N_20204,N_23895);
xor U27128 (N_27128,N_24989,N_20779);
xnor U27129 (N_27129,N_23361,N_22223);
nor U27130 (N_27130,N_23804,N_23620);
nor U27131 (N_27131,N_24827,N_20373);
or U27132 (N_27132,N_23769,N_24112);
nand U27133 (N_27133,N_22510,N_20626);
nand U27134 (N_27134,N_22786,N_20265);
nor U27135 (N_27135,N_23067,N_23345);
nand U27136 (N_27136,N_22800,N_21810);
nor U27137 (N_27137,N_23364,N_24339);
and U27138 (N_27138,N_24641,N_23030);
and U27139 (N_27139,N_20845,N_23309);
or U27140 (N_27140,N_24432,N_20491);
nor U27141 (N_27141,N_23400,N_24351);
and U27142 (N_27142,N_20551,N_21473);
nand U27143 (N_27143,N_23448,N_22759);
nand U27144 (N_27144,N_23640,N_20803);
nand U27145 (N_27145,N_20371,N_23357);
and U27146 (N_27146,N_22896,N_23811);
or U27147 (N_27147,N_21244,N_21258);
nor U27148 (N_27148,N_23661,N_20486);
and U27149 (N_27149,N_20822,N_22912);
or U27150 (N_27150,N_20464,N_20380);
and U27151 (N_27151,N_24263,N_24944);
nor U27152 (N_27152,N_21447,N_24256);
nand U27153 (N_27153,N_24392,N_24930);
nor U27154 (N_27154,N_24797,N_22628);
nor U27155 (N_27155,N_22463,N_21612);
nand U27156 (N_27156,N_22907,N_20902);
and U27157 (N_27157,N_24337,N_20479);
nor U27158 (N_27158,N_24147,N_23057);
nor U27159 (N_27159,N_23533,N_23845);
or U27160 (N_27160,N_24591,N_23020);
nor U27161 (N_27161,N_21305,N_24756);
and U27162 (N_27162,N_24576,N_23633);
and U27163 (N_27163,N_20989,N_21361);
nand U27164 (N_27164,N_24539,N_23199);
and U27165 (N_27165,N_23353,N_21586);
nor U27166 (N_27166,N_22294,N_22094);
and U27167 (N_27167,N_23652,N_20796);
nor U27168 (N_27168,N_20159,N_24501);
xnor U27169 (N_27169,N_21290,N_24677);
or U27170 (N_27170,N_24543,N_23647);
and U27171 (N_27171,N_20647,N_24408);
nand U27172 (N_27172,N_21308,N_20302);
xnor U27173 (N_27173,N_20535,N_20147);
or U27174 (N_27174,N_20678,N_21163);
xnor U27175 (N_27175,N_22419,N_21933);
nor U27176 (N_27176,N_23495,N_24438);
and U27177 (N_27177,N_22771,N_24410);
nand U27178 (N_27178,N_24138,N_22205);
nor U27179 (N_27179,N_21688,N_22404);
nand U27180 (N_27180,N_20905,N_21574);
nand U27181 (N_27181,N_22954,N_23754);
or U27182 (N_27182,N_21094,N_21004);
nor U27183 (N_27183,N_20333,N_21626);
and U27184 (N_27184,N_22138,N_22591);
nor U27185 (N_27185,N_22836,N_23382);
nor U27186 (N_27186,N_24260,N_20415);
xor U27187 (N_27187,N_22457,N_23209);
nor U27188 (N_27188,N_20531,N_23312);
xor U27189 (N_27189,N_22732,N_20367);
nor U27190 (N_27190,N_22221,N_22821);
and U27191 (N_27191,N_24779,N_24017);
or U27192 (N_27192,N_22009,N_20994);
nor U27193 (N_27193,N_22014,N_23913);
and U27194 (N_27194,N_21293,N_20195);
and U27195 (N_27195,N_22503,N_20799);
nor U27196 (N_27196,N_24459,N_23527);
nand U27197 (N_27197,N_22028,N_23906);
nor U27198 (N_27198,N_23503,N_20995);
nor U27199 (N_27199,N_23230,N_20431);
xnor U27200 (N_27200,N_22326,N_23673);
xor U27201 (N_27201,N_21743,N_21022);
and U27202 (N_27202,N_21487,N_23147);
xor U27203 (N_27203,N_21822,N_22251);
or U27204 (N_27204,N_20950,N_22345);
xor U27205 (N_27205,N_23607,N_23758);
nand U27206 (N_27206,N_23391,N_23990);
and U27207 (N_27207,N_24694,N_22977);
nand U27208 (N_27208,N_22952,N_21206);
and U27209 (N_27209,N_24548,N_23359);
and U27210 (N_27210,N_22664,N_21492);
nor U27211 (N_27211,N_21842,N_24590);
xnor U27212 (N_27212,N_22844,N_21678);
and U27213 (N_27213,N_21752,N_24485);
or U27214 (N_27214,N_20942,N_24296);
or U27215 (N_27215,N_21475,N_24381);
or U27216 (N_27216,N_23513,N_21561);
nand U27217 (N_27217,N_22889,N_22464);
or U27218 (N_27218,N_24023,N_23660);
nand U27219 (N_27219,N_23926,N_23967);
xnor U27220 (N_27220,N_20430,N_24058);
xor U27221 (N_27221,N_21654,N_24041);
nor U27222 (N_27222,N_21433,N_23952);
xor U27223 (N_27223,N_21849,N_22966);
nand U27224 (N_27224,N_24584,N_21045);
xnor U27225 (N_27225,N_23295,N_20664);
and U27226 (N_27226,N_21248,N_20908);
nor U27227 (N_27227,N_23840,N_20502);
nand U27228 (N_27228,N_23292,N_21239);
and U27229 (N_27229,N_20245,N_21589);
xnor U27230 (N_27230,N_20934,N_24202);
xnor U27231 (N_27231,N_21265,N_24503);
or U27232 (N_27232,N_23374,N_21556);
nand U27233 (N_27233,N_22352,N_20756);
nor U27234 (N_27234,N_24383,N_20760);
xor U27235 (N_27235,N_21444,N_23719);
nor U27236 (N_27236,N_20509,N_24830);
nand U27237 (N_27237,N_21296,N_22938);
xor U27238 (N_27238,N_24929,N_23436);
or U27239 (N_27239,N_22647,N_21223);
or U27240 (N_27240,N_20224,N_23892);
and U27241 (N_27241,N_24078,N_21532);
xor U27242 (N_27242,N_22745,N_24561);
nand U27243 (N_27243,N_24848,N_21730);
nand U27244 (N_27244,N_22824,N_22837);
and U27245 (N_27245,N_24592,N_22108);
or U27246 (N_27246,N_22241,N_24216);
xor U27247 (N_27247,N_21002,N_20880);
or U27248 (N_27248,N_21951,N_22833);
and U27249 (N_27249,N_20736,N_22282);
nor U27250 (N_27250,N_20446,N_21076);
nand U27251 (N_27251,N_21564,N_20381);
nand U27252 (N_27252,N_21964,N_21019);
nor U27253 (N_27253,N_23376,N_20718);
or U27254 (N_27254,N_22605,N_21578);
or U27255 (N_27255,N_23013,N_21792);
nand U27256 (N_27256,N_22495,N_23819);
or U27257 (N_27257,N_20318,N_20721);
xnor U27258 (N_27258,N_23993,N_23296);
nand U27259 (N_27259,N_21649,N_21388);
or U27260 (N_27260,N_21268,N_23249);
nor U27261 (N_27261,N_23534,N_23787);
nor U27262 (N_27262,N_21837,N_22106);
nand U27263 (N_27263,N_21553,N_20437);
or U27264 (N_27264,N_21003,N_23700);
nor U27265 (N_27265,N_24716,N_23771);
nor U27266 (N_27266,N_20078,N_21807);
nand U27267 (N_27267,N_24152,N_22133);
xnor U27268 (N_27268,N_23517,N_21089);
nand U27269 (N_27269,N_20076,N_22414);
xor U27270 (N_27270,N_20493,N_24226);
xor U27271 (N_27271,N_20660,N_21355);
nand U27272 (N_27272,N_21699,N_22475);
or U27273 (N_27273,N_24697,N_22359);
xnor U27274 (N_27274,N_24292,N_24361);
nor U27275 (N_27275,N_22228,N_21345);
nand U27276 (N_27276,N_21194,N_23648);
or U27277 (N_27277,N_22682,N_24007);
and U27278 (N_27278,N_23603,N_22017);
nor U27279 (N_27279,N_20428,N_20196);
and U27280 (N_27280,N_24302,N_20568);
or U27281 (N_27281,N_20911,N_20561);
and U27282 (N_27282,N_22107,N_23902);
xor U27283 (N_27283,N_20930,N_22328);
or U27284 (N_27284,N_21119,N_23709);
nor U27285 (N_27285,N_23614,N_21588);
xnor U27286 (N_27286,N_23102,N_20004);
nor U27287 (N_27287,N_23861,N_22305);
and U27288 (N_27288,N_21271,N_20408);
or U27289 (N_27289,N_22531,N_21544);
nor U27290 (N_27290,N_24810,N_21868);
or U27291 (N_27291,N_22049,N_22237);
nor U27292 (N_27292,N_24206,N_24274);
or U27293 (N_27293,N_20444,N_22549);
or U27294 (N_27294,N_23951,N_23100);
and U27295 (N_27295,N_24831,N_21292);
nand U27296 (N_27296,N_22971,N_24943);
xor U27297 (N_27297,N_20786,N_20131);
xor U27298 (N_27298,N_24555,N_23127);
and U27299 (N_27299,N_22026,N_24201);
nor U27300 (N_27300,N_20098,N_24817);
and U27301 (N_27301,N_23258,N_21986);
xor U27302 (N_27302,N_20368,N_22137);
and U27303 (N_27303,N_22756,N_20659);
xnor U27304 (N_27304,N_20141,N_23118);
nand U27305 (N_27305,N_23991,N_24725);
or U27306 (N_27306,N_21143,N_23490);
nor U27307 (N_27307,N_22876,N_21373);
xor U27308 (N_27308,N_24214,N_21323);
and U27309 (N_27309,N_23516,N_20236);
xnor U27310 (N_27310,N_20185,N_20879);
nand U27311 (N_27311,N_24132,N_23567);
and U27312 (N_27312,N_22846,N_23930);
nor U27313 (N_27313,N_24844,N_24764);
nand U27314 (N_27314,N_22618,N_21939);
or U27315 (N_27315,N_23291,N_24130);
xnor U27316 (N_27316,N_21181,N_23110);
nand U27317 (N_27317,N_24473,N_23744);
nor U27318 (N_27318,N_23035,N_23807);
or U27319 (N_27319,N_23928,N_22330);
xor U27320 (N_27320,N_23943,N_22930);
nand U27321 (N_27321,N_21621,N_20685);
and U27322 (N_27322,N_24396,N_22705);
or U27323 (N_27323,N_24184,N_22443);
xor U27324 (N_27324,N_24479,N_20747);
xnor U27325 (N_27325,N_21440,N_23167);
xnor U27326 (N_27326,N_23638,N_20397);
nor U27327 (N_27327,N_21686,N_24067);
or U27328 (N_27328,N_22636,N_22568);
or U27329 (N_27329,N_23275,N_24825);
or U27330 (N_27330,N_22940,N_22674);
nand U27331 (N_27331,N_21982,N_21702);
and U27332 (N_27332,N_22744,N_22630);
nor U27333 (N_27333,N_21983,N_24131);
nand U27334 (N_27334,N_23192,N_24443);
nand U27335 (N_27335,N_23739,N_21238);
nand U27336 (N_27336,N_20823,N_20137);
or U27337 (N_27337,N_20157,N_22010);
xnor U27338 (N_27338,N_23664,N_21012);
nor U27339 (N_27339,N_20069,N_20545);
or U27340 (N_27340,N_20610,N_22812);
nand U27341 (N_27341,N_23877,N_24136);
xor U27342 (N_27342,N_24546,N_22067);
and U27343 (N_27343,N_21212,N_24419);
and U27344 (N_27344,N_20984,N_23921);
or U27345 (N_27345,N_21845,N_21666);
xnor U27346 (N_27346,N_24048,N_24673);
nor U27347 (N_27347,N_20870,N_23728);
nor U27348 (N_27348,N_24701,N_24093);
nor U27349 (N_27349,N_24647,N_21309);
or U27350 (N_27350,N_21838,N_21821);
nor U27351 (N_27351,N_21569,N_20723);
or U27352 (N_27352,N_20940,N_20223);
and U27353 (N_27353,N_21665,N_20111);
nor U27354 (N_27354,N_24467,N_23144);
or U27355 (N_27355,N_24203,N_21955);
and U27356 (N_27356,N_24011,N_20604);
and U27357 (N_27357,N_20122,N_22291);
xor U27358 (N_27358,N_24715,N_23263);
or U27359 (N_27359,N_24095,N_20197);
xor U27360 (N_27360,N_24364,N_21804);
or U27361 (N_27361,N_20692,N_22379);
nand U27362 (N_27362,N_23212,N_20602);
xnor U27363 (N_27363,N_22135,N_22789);
nand U27364 (N_27364,N_23762,N_22773);
nor U27365 (N_27365,N_24434,N_23512);
xnor U27366 (N_27366,N_20029,N_20300);
and U27367 (N_27367,N_24401,N_20256);
nand U27368 (N_27368,N_24538,N_21020);
or U27369 (N_27369,N_21768,N_24949);
nand U27370 (N_27370,N_23780,N_21284);
nor U27371 (N_27371,N_21120,N_23741);
nor U27372 (N_27372,N_21425,N_24013);
or U27373 (N_27373,N_21205,N_23429);
and U27374 (N_27374,N_21664,N_20949);
and U27375 (N_27375,N_20288,N_21507);
or U27376 (N_27376,N_21391,N_23497);
nand U27377 (N_27377,N_22447,N_24049);
or U27378 (N_27378,N_20126,N_22304);
xor U27379 (N_27379,N_23960,N_22439);
and U27380 (N_27380,N_21925,N_21384);
or U27381 (N_27381,N_23228,N_20407);
and U27382 (N_27382,N_20619,N_21554);
nor U27383 (N_27383,N_21099,N_21504);
or U27384 (N_27384,N_24612,N_21513);
and U27385 (N_27385,N_24077,N_24920);
xnor U27386 (N_27386,N_23113,N_23871);
or U27387 (N_27387,N_23535,N_20530);
or U27388 (N_27388,N_23272,N_21766);
xor U27389 (N_27389,N_21854,N_23985);
and U27390 (N_27390,N_21100,N_20793);
or U27391 (N_27391,N_23103,N_21452);
nand U27392 (N_27392,N_24423,N_22157);
xnor U27393 (N_27393,N_20322,N_21562);
or U27394 (N_27394,N_20712,N_20030);
nand U27395 (N_27395,N_24668,N_20507);
and U27396 (N_27396,N_24709,N_20836);
xnor U27397 (N_27397,N_24794,N_21894);
nand U27398 (N_27398,N_22979,N_21853);
nor U27399 (N_27399,N_21167,N_21208);
nor U27400 (N_27400,N_24429,N_24660);
or U27401 (N_27401,N_24771,N_20722);
or U27402 (N_27402,N_22082,N_23759);
and U27403 (N_27403,N_21263,N_24509);
xor U27404 (N_27404,N_23904,N_22669);
or U27405 (N_27405,N_22434,N_20077);
or U27406 (N_27406,N_24404,N_22694);
or U27407 (N_27407,N_23644,N_20347);
or U27408 (N_27408,N_24062,N_23677);
and U27409 (N_27409,N_22275,N_22431);
nor U27410 (N_27410,N_20778,N_23428);
nand U27411 (N_27411,N_23976,N_24648);
or U27412 (N_27412,N_21314,N_21262);
and U27413 (N_27413,N_21160,N_22617);
nand U27414 (N_27414,N_23611,N_20068);
xor U27415 (N_27415,N_24139,N_23653);
or U27416 (N_27416,N_21992,N_22619);
or U27417 (N_27417,N_24679,N_21566);
or U27418 (N_27418,N_24422,N_23615);
xor U27419 (N_27419,N_21601,N_22388);
or U27420 (N_27420,N_23703,N_23473);
xor U27421 (N_27421,N_20953,N_21123);
or U27422 (N_27422,N_23829,N_22685);
xnor U27423 (N_27423,N_22346,N_24307);
nor U27424 (N_27424,N_20216,N_22958);
and U27425 (N_27425,N_23434,N_24991);
or U27426 (N_27426,N_21393,N_20820);
and U27427 (N_27427,N_22450,N_24279);
xnor U27428 (N_27428,N_24223,N_22008);
nor U27429 (N_27429,N_22482,N_20883);
nand U27430 (N_27430,N_22631,N_24804);
nand U27431 (N_27431,N_22571,N_20353);
or U27432 (N_27432,N_21465,N_23134);
and U27433 (N_27433,N_23818,N_24853);
xnor U27434 (N_27434,N_21443,N_21007);
and U27435 (N_27435,N_20931,N_21851);
and U27436 (N_27436,N_22687,N_20150);
and U27437 (N_27437,N_23539,N_20854);
nand U27438 (N_27438,N_20319,N_22945);
and U27439 (N_27439,N_23736,N_20560);
xor U27440 (N_27440,N_21706,N_24161);
nor U27441 (N_27441,N_21874,N_21046);
nor U27442 (N_27442,N_21658,N_24534);
xor U27443 (N_27443,N_20683,N_23070);
xor U27444 (N_27444,N_22174,N_20826);
nand U27445 (N_27445,N_22369,N_23259);
or U27446 (N_27446,N_21592,N_24608);
nand U27447 (N_27447,N_22381,N_23033);
or U27448 (N_27448,N_23283,N_20448);
or U27449 (N_27449,N_23584,N_23152);
nor U27450 (N_27450,N_23919,N_21038);
xnor U27451 (N_27451,N_20366,N_22497);
nand U27452 (N_27452,N_20217,N_22585);
nor U27453 (N_27453,N_24315,N_24080);
or U27454 (N_27454,N_21551,N_23850);
and U27455 (N_27455,N_20241,N_21511);
and U27456 (N_27456,N_22804,N_21395);
nand U27457 (N_27457,N_22739,N_24686);
xnor U27458 (N_27458,N_23763,N_23038);
or U27459 (N_27459,N_24465,N_20873);
nand U27460 (N_27460,N_23339,N_24287);
nor U27461 (N_27461,N_23403,N_20690);
and U27462 (N_27462,N_22040,N_24782);
xor U27463 (N_27463,N_23093,N_20877);
and U27464 (N_27464,N_23966,N_24959);
nor U27465 (N_27465,N_21788,N_20518);
nor U27466 (N_27466,N_20284,N_23803);
and U27467 (N_27467,N_24241,N_20567);
xor U27468 (N_27468,N_23859,N_21728);
xor U27469 (N_27469,N_20752,N_24316);
xor U27470 (N_27470,N_22555,N_21828);
and U27471 (N_27471,N_24675,N_24545);
xnor U27472 (N_27472,N_21506,N_23983);
and U27473 (N_27473,N_21320,N_21213);
nor U27474 (N_27474,N_23896,N_23120);
xor U27475 (N_27475,N_22957,N_20895);
xnor U27476 (N_27476,N_22880,N_20379);
and U27477 (N_27477,N_23796,N_21950);
nor U27478 (N_27478,N_22188,N_23041);
nor U27479 (N_27479,N_23143,N_23419);
nor U27480 (N_27480,N_22160,N_24834);
xnor U27481 (N_27481,N_21826,N_22891);
xor U27482 (N_27482,N_21402,N_20524);
nor U27483 (N_27483,N_23287,N_21767);
nor U27484 (N_27484,N_24436,N_23855);
xnor U27485 (N_27485,N_21560,N_21312);
nand U27486 (N_27486,N_20120,N_24191);
and U27487 (N_27487,N_22365,N_20421);
or U27488 (N_27488,N_21655,N_20814);
or U27489 (N_27489,N_20292,N_22144);
nand U27490 (N_27490,N_24004,N_23962);
nor U27491 (N_27491,N_24523,N_23613);
or U27492 (N_27492,N_24164,N_20438);
or U27493 (N_27493,N_22603,N_23779);
or U27494 (N_27494,N_23399,N_23229);
nor U27495 (N_27495,N_20761,N_20210);
nand U27496 (N_27496,N_24437,N_23915);
and U27497 (N_27497,N_20601,N_23544);
or U27498 (N_27498,N_23487,N_22818);
and U27499 (N_27499,N_22576,N_20113);
or U27500 (N_27500,N_23506,N_22709);
xnor U27501 (N_27501,N_21047,N_24224);
nand U27502 (N_27502,N_24063,N_23164);
and U27503 (N_27503,N_22000,N_21222);
nand U27504 (N_27504,N_20731,N_24472);
and U27505 (N_27505,N_23053,N_24544);
xnor U27506 (N_27506,N_22169,N_20523);
xnor U27507 (N_27507,N_24969,N_20749);
and U27508 (N_27508,N_20340,N_24561);
or U27509 (N_27509,N_24472,N_23961);
nor U27510 (N_27510,N_22619,N_23787);
nor U27511 (N_27511,N_21738,N_21621);
or U27512 (N_27512,N_21316,N_21858);
nand U27513 (N_27513,N_23538,N_21483);
or U27514 (N_27514,N_24451,N_20898);
nand U27515 (N_27515,N_22256,N_22023);
nor U27516 (N_27516,N_21816,N_20832);
or U27517 (N_27517,N_22400,N_20807);
nor U27518 (N_27518,N_23293,N_23512);
and U27519 (N_27519,N_23729,N_20206);
or U27520 (N_27520,N_22331,N_20032);
and U27521 (N_27521,N_23867,N_20183);
xnor U27522 (N_27522,N_21018,N_22476);
nand U27523 (N_27523,N_24189,N_24735);
nand U27524 (N_27524,N_20692,N_21407);
nor U27525 (N_27525,N_24477,N_23982);
nand U27526 (N_27526,N_24106,N_23793);
and U27527 (N_27527,N_21145,N_23003);
xnor U27528 (N_27528,N_24792,N_21877);
and U27529 (N_27529,N_22236,N_21282);
or U27530 (N_27530,N_22081,N_23207);
nor U27531 (N_27531,N_24270,N_22309);
nor U27532 (N_27532,N_22137,N_23966);
or U27533 (N_27533,N_20714,N_24589);
nand U27534 (N_27534,N_22686,N_20339);
nor U27535 (N_27535,N_23663,N_23579);
and U27536 (N_27536,N_21656,N_20346);
nand U27537 (N_27537,N_20569,N_22442);
nand U27538 (N_27538,N_20517,N_22433);
and U27539 (N_27539,N_21543,N_22351);
nand U27540 (N_27540,N_23891,N_23928);
and U27541 (N_27541,N_24681,N_21873);
nor U27542 (N_27542,N_24797,N_20701);
xor U27543 (N_27543,N_24996,N_21438);
or U27544 (N_27544,N_24210,N_23118);
and U27545 (N_27545,N_23425,N_20906);
and U27546 (N_27546,N_23790,N_22364);
or U27547 (N_27547,N_21848,N_24653);
or U27548 (N_27548,N_21096,N_20467);
or U27549 (N_27549,N_24569,N_22841);
or U27550 (N_27550,N_23247,N_20977);
or U27551 (N_27551,N_24351,N_22984);
nor U27552 (N_27552,N_21441,N_23283);
nand U27553 (N_27553,N_21425,N_24785);
or U27554 (N_27554,N_24988,N_22208);
xor U27555 (N_27555,N_20252,N_22181);
or U27556 (N_27556,N_23318,N_21114);
or U27557 (N_27557,N_23841,N_23901);
nor U27558 (N_27558,N_20698,N_20473);
or U27559 (N_27559,N_22526,N_23579);
or U27560 (N_27560,N_24907,N_24939);
xor U27561 (N_27561,N_20163,N_22323);
nor U27562 (N_27562,N_23299,N_22194);
and U27563 (N_27563,N_20604,N_20967);
nor U27564 (N_27564,N_23342,N_24111);
nor U27565 (N_27565,N_22920,N_21877);
nor U27566 (N_27566,N_21323,N_24450);
or U27567 (N_27567,N_22743,N_21954);
and U27568 (N_27568,N_24725,N_22587);
nor U27569 (N_27569,N_23688,N_22871);
and U27570 (N_27570,N_23645,N_21021);
or U27571 (N_27571,N_23762,N_20927);
nand U27572 (N_27572,N_23059,N_20149);
or U27573 (N_27573,N_21920,N_24522);
or U27574 (N_27574,N_20521,N_23501);
nor U27575 (N_27575,N_23559,N_20586);
xnor U27576 (N_27576,N_20451,N_21529);
nand U27577 (N_27577,N_21889,N_21593);
or U27578 (N_27578,N_20961,N_23360);
nand U27579 (N_27579,N_22102,N_24989);
and U27580 (N_27580,N_21595,N_22994);
and U27581 (N_27581,N_20394,N_23223);
nor U27582 (N_27582,N_22529,N_22699);
or U27583 (N_27583,N_22217,N_24865);
or U27584 (N_27584,N_23510,N_22171);
and U27585 (N_27585,N_22178,N_23687);
and U27586 (N_27586,N_22977,N_22062);
and U27587 (N_27587,N_22641,N_23451);
and U27588 (N_27588,N_21916,N_24056);
and U27589 (N_27589,N_23892,N_21747);
xnor U27590 (N_27590,N_21109,N_23105);
xor U27591 (N_27591,N_22470,N_22112);
and U27592 (N_27592,N_22182,N_22438);
nor U27593 (N_27593,N_20617,N_24346);
xnor U27594 (N_27594,N_22708,N_24634);
xor U27595 (N_27595,N_23871,N_23670);
nor U27596 (N_27596,N_23716,N_20892);
nand U27597 (N_27597,N_20110,N_21480);
nor U27598 (N_27598,N_23183,N_24845);
nand U27599 (N_27599,N_24426,N_24421);
nor U27600 (N_27600,N_21472,N_20931);
or U27601 (N_27601,N_21942,N_21551);
nand U27602 (N_27602,N_22868,N_21343);
or U27603 (N_27603,N_20456,N_22069);
or U27604 (N_27604,N_20471,N_23696);
nor U27605 (N_27605,N_21988,N_20101);
nor U27606 (N_27606,N_22656,N_21290);
nand U27607 (N_27607,N_22083,N_20500);
and U27608 (N_27608,N_22622,N_23384);
nor U27609 (N_27609,N_24889,N_24519);
xor U27610 (N_27610,N_20396,N_24425);
and U27611 (N_27611,N_24676,N_23356);
nor U27612 (N_27612,N_20426,N_23630);
or U27613 (N_27613,N_20199,N_23840);
nor U27614 (N_27614,N_20725,N_21222);
or U27615 (N_27615,N_24052,N_24823);
xor U27616 (N_27616,N_24815,N_20529);
and U27617 (N_27617,N_20884,N_21956);
nand U27618 (N_27618,N_20130,N_21452);
nand U27619 (N_27619,N_21079,N_24065);
or U27620 (N_27620,N_24519,N_22799);
xor U27621 (N_27621,N_20405,N_23671);
nand U27622 (N_27622,N_21779,N_22640);
nand U27623 (N_27623,N_22139,N_20133);
or U27624 (N_27624,N_24657,N_20036);
xnor U27625 (N_27625,N_23845,N_23996);
nor U27626 (N_27626,N_24404,N_23535);
nor U27627 (N_27627,N_21552,N_24772);
xor U27628 (N_27628,N_24395,N_22800);
or U27629 (N_27629,N_24552,N_20397);
or U27630 (N_27630,N_20764,N_24302);
or U27631 (N_27631,N_22932,N_20975);
and U27632 (N_27632,N_24721,N_21600);
xnor U27633 (N_27633,N_22776,N_22038);
or U27634 (N_27634,N_22466,N_24402);
or U27635 (N_27635,N_21066,N_24419);
nor U27636 (N_27636,N_21369,N_24817);
nor U27637 (N_27637,N_23921,N_22225);
nor U27638 (N_27638,N_20250,N_20016);
and U27639 (N_27639,N_20731,N_21573);
nand U27640 (N_27640,N_24944,N_21594);
nand U27641 (N_27641,N_22330,N_21908);
nand U27642 (N_27642,N_22383,N_23007);
xnor U27643 (N_27643,N_22656,N_20757);
xor U27644 (N_27644,N_20857,N_24947);
xnor U27645 (N_27645,N_24189,N_24978);
nor U27646 (N_27646,N_20150,N_22738);
nand U27647 (N_27647,N_20550,N_23601);
xor U27648 (N_27648,N_24981,N_21296);
xor U27649 (N_27649,N_23046,N_21832);
nor U27650 (N_27650,N_23733,N_21982);
xnor U27651 (N_27651,N_21450,N_24798);
nor U27652 (N_27652,N_23638,N_24565);
xnor U27653 (N_27653,N_22882,N_22336);
nand U27654 (N_27654,N_20561,N_21558);
and U27655 (N_27655,N_20855,N_20242);
xor U27656 (N_27656,N_23911,N_21674);
xnor U27657 (N_27657,N_20248,N_24773);
xnor U27658 (N_27658,N_21406,N_20746);
and U27659 (N_27659,N_21417,N_20078);
and U27660 (N_27660,N_20599,N_20601);
or U27661 (N_27661,N_20048,N_22800);
xnor U27662 (N_27662,N_23156,N_24354);
nor U27663 (N_27663,N_24675,N_20849);
or U27664 (N_27664,N_21190,N_22471);
or U27665 (N_27665,N_21847,N_21638);
nand U27666 (N_27666,N_24603,N_22515);
xnor U27667 (N_27667,N_24708,N_23224);
or U27668 (N_27668,N_22342,N_20232);
and U27669 (N_27669,N_22383,N_23805);
xor U27670 (N_27670,N_24203,N_24515);
or U27671 (N_27671,N_24013,N_21982);
and U27672 (N_27672,N_21560,N_24900);
and U27673 (N_27673,N_21419,N_20250);
xnor U27674 (N_27674,N_22043,N_23843);
or U27675 (N_27675,N_23920,N_22425);
nor U27676 (N_27676,N_24542,N_20281);
nand U27677 (N_27677,N_22105,N_21405);
nand U27678 (N_27678,N_23826,N_21881);
nand U27679 (N_27679,N_23328,N_22485);
nand U27680 (N_27680,N_24252,N_22511);
or U27681 (N_27681,N_24895,N_21903);
and U27682 (N_27682,N_21067,N_23121);
or U27683 (N_27683,N_22893,N_23047);
and U27684 (N_27684,N_20457,N_20721);
or U27685 (N_27685,N_21704,N_21291);
or U27686 (N_27686,N_22641,N_22701);
nand U27687 (N_27687,N_21237,N_24911);
and U27688 (N_27688,N_21219,N_21368);
nand U27689 (N_27689,N_20668,N_20892);
or U27690 (N_27690,N_22769,N_23815);
xor U27691 (N_27691,N_21648,N_21820);
or U27692 (N_27692,N_20260,N_24978);
or U27693 (N_27693,N_21006,N_24638);
and U27694 (N_27694,N_20467,N_22295);
or U27695 (N_27695,N_22580,N_21770);
or U27696 (N_27696,N_20809,N_23950);
and U27697 (N_27697,N_21733,N_23588);
nand U27698 (N_27698,N_23306,N_22729);
nand U27699 (N_27699,N_23483,N_24466);
nor U27700 (N_27700,N_20773,N_23392);
xor U27701 (N_27701,N_21757,N_20954);
and U27702 (N_27702,N_21055,N_24557);
and U27703 (N_27703,N_21615,N_20196);
or U27704 (N_27704,N_22979,N_21080);
and U27705 (N_27705,N_21315,N_21821);
or U27706 (N_27706,N_21546,N_23941);
xor U27707 (N_27707,N_24446,N_23585);
xor U27708 (N_27708,N_23448,N_23266);
xor U27709 (N_27709,N_23875,N_21333);
nand U27710 (N_27710,N_20514,N_24210);
xor U27711 (N_27711,N_22609,N_23474);
and U27712 (N_27712,N_20337,N_22614);
and U27713 (N_27713,N_20595,N_20028);
xnor U27714 (N_27714,N_24827,N_22308);
nor U27715 (N_27715,N_20434,N_21811);
nand U27716 (N_27716,N_20912,N_20485);
nor U27717 (N_27717,N_21035,N_22734);
nor U27718 (N_27718,N_21483,N_21619);
nand U27719 (N_27719,N_23343,N_20037);
nor U27720 (N_27720,N_22892,N_23145);
nor U27721 (N_27721,N_22351,N_20061);
and U27722 (N_27722,N_21578,N_24294);
xnor U27723 (N_27723,N_20477,N_24178);
or U27724 (N_27724,N_22983,N_21769);
xor U27725 (N_27725,N_23875,N_23103);
xnor U27726 (N_27726,N_23277,N_21651);
or U27727 (N_27727,N_24408,N_22513);
or U27728 (N_27728,N_24138,N_24133);
nand U27729 (N_27729,N_21757,N_24355);
nand U27730 (N_27730,N_23449,N_20867);
nor U27731 (N_27731,N_21985,N_20452);
nand U27732 (N_27732,N_23963,N_21667);
and U27733 (N_27733,N_23996,N_21031);
nand U27734 (N_27734,N_22160,N_24446);
nand U27735 (N_27735,N_23995,N_23889);
nand U27736 (N_27736,N_23410,N_20834);
xor U27737 (N_27737,N_22821,N_24449);
nor U27738 (N_27738,N_21779,N_21514);
and U27739 (N_27739,N_22728,N_21102);
and U27740 (N_27740,N_24596,N_24957);
nor U27741 (N_27741,N_21405,N_22345);
xor U27742 (N_27742,N_20618,N_24807);
and U27743 (N_27743,N_22638,N_21428);
or U27744 (N_27744,N_20940,N_20627);
or U27745 (N_27745,N_20972,N_22496);
xor U27746 (N_27746,N_21436,N_23279);
xor U27747 (N_27747,N_22353,N_23917);
nand U27748 (N_27748,N_22558,N_23966);
or U27749 (N_27749,N_20258,N_21084);
nand U27750 (N_27750,N_22641,N_23126);
nand U27751 (N_27751,N_20407,N_23727);
nor U27752 (N_27752,N_20845,N_24117);
and U27753 (N_27753,N_22554,N_23758);
nor U27754 (N_27754,N_20499,N_20836);
or U27755 (N_27755,N_21466,N_22988);
or U27756 (N_27756,N_23556,N_22215);
or U27757 (N_27757,N_23887,N_23188);
or U27758 (N_27758,N_21162,N_21021);
and U27759 (N_27759,N_21115,N_24699);
and U27760 (N_27760,N_21468,N_24835);
xor U27761 (N_27761,N_20364,N_22792);
or U27762 (N_27762,N_24432,N_21297);
and U27763 (N_27763,N_23589,N_23432);
nor U27764 (N_27764,N_22722,N_23286);
and U27765 (N_27765,N_23705,N_24970);
nor U27766 (N_27766,N_24291,N_21605);
nand U27767 (N_27767,N_20985,N_22054);
and U27768 (N_27768,N_20630,N_20748);
xnor U27769 (N_27769,N_21745,N_21308);
xor U27770 (N_27770,N_20855,N_21241);
nor U27771 (N_27771,N_24175,N_23029);
nand U27772 (N_27772,N_23627,N_24168);
xnor U27773 (N_27773,N_21249,N_23720);
xor U27774 (N_27774,N_22716,N_21335);
or U27775 (N_27775,N_21916,N_21170);
and U27776 (N_27776,N_22734,N_24462);
nor U27777 (N_27777,N_20293,N_22944);
xnor U27778 (N_27778,N_20146,N_23432);
xor U27779 (N_27779,N_23269,N_24802);
nor U27780 (N_27780,N_22869,N_24119);
and U27781 (N_27781,N_22645,N_23129);
or U27782 (N_27782,N_20975,N_21906);
nand U27783 (N_27783,N_22361,N_20885);
nor U27784 (N_27784,N_23291,N_21854);
nand U27785 (N_27785,N_22079,N_20487);
xor U27786 (N_27786,N_21595,N_24447);
or U27787 (N_27787,N_24762,N_23316);
nor U27788 (N_27788,N_24229,N_21965);
xor U27789 (N_27789,N_20913,N_23080);
or U27790 (N_27790,N_22919,N_22176);
or U27791 (N_27791,N_23886,N_20530);
nor U27792 (N_27792,N_20432,N_23144);
xor U27793 (N_27793,N_22554,N_21660);
or U27794 (N_27794,N_21544,N_22154);
and U27795 (N_27795,N_22787,N_23248);
and U27796 (N_27796,N_23807,N_20628);
and U27797 (N_27797,N_24939,N_22139);
or U27798 (N_27798,N_21466,N_23033);
nand U27799 (N_27799,N_23836,N_20370);
and U27800 (N_27800,N_24470,N_24873);
xnor U27801 (N_27801,N_20095,N_24499);
nor U27802 (N_27802,N_23516,N_21671);
nor U27803 (N_27803,N_23358,N_20369);
and U27804 (N_27804,N_24587,N_24896);
nand U27805 (N_27805,N_23183,N_21447);
xnor U27806 (N_27806,N_24801,N_20370);
nand U27807 (N_27807,N_20587,N_22118);
and U27808 (N_27808,N_24607,N_20454);
or U27809 (N_27809,N_21340,N_20761);
xor U27810 (N_27810,N_22816,N_21027);
and U27811 (N_27811,N_21395,N_22227);
nor U27812 (N_27812,N_23253,N_21380);
or U27813 (N_27813,N_20243,N_20471);
or U27814 (N_27814,N_21531,N_22700);
nand U27815 (N_27815,N_21506,N_24048);
and U27816 (N_27816,N_22785,N_21460);
or U27817 (N_27817,N_23819,N_22632);
and U27818 (N_27818,N_21549,N_24209);
xnor U27819 (N_27819,N_23648,N_21302);
and U27820 (N_27820,N_23874,N_24157);
nor U27821 (N_27821,N_23470,N_21051);
nor U27822 (N_27822,N_21942,N_24826);
nor U27823 (N_27823,N_24627,N_24945);
or U27824 (N_27824,N_24663,N_23769);
nand U27825 (N_27825,N_20323,N_21930);
and U27826 (N_27826,N_24739,N_23525);
nand U27827 (N_27827,N_21318,N_21980);
nor U27828 (N_27828,N_24746,N_22337);
xor U27829 (N_27829,N_24260,N_21218);
xnor U27830 (N_27830,N_23588,N_22066);
nor U27831 (N_27831,N_20448,N_23173);
or U27832 (N_27832,N_23439,N_20212);
nand U27833 (N_27833,N_20249,N_20610);
nand U27834 (N_27834,N_20607,N_22395);
nand U27835 (N_27835,N_24108,N_20843);
nor U27836 (N_27836,N_21875,N_21625);
xor U27837 (N_27837,N_24919,N_21992);
nor U27838 (N_27838,N_22138,N_22924);
or U27839 (N_27839,N_21526,N_24123);
or U27840 (N_27840,N_24504,N_22222);
and U27841 (N_27841,N_24864,N_23238);
xor U27842 (N_27842,N_22772,N_24350);
nand U27843 (N_27843,N_24736,N_22850);
or U27844 (N_27844,N_22020,N_21273);
or U27845 (N_27845,N_20557,N_24351);
nand U27846 (N_27846,N_22226,N_21506);
nand U27847 (N_27847,N_24293,N_22644);
nor U27848 (N_27848,N_21505,N_24000);
nor U27849 (N_27849,N_22899,N_22959);
and U27850 (N_27850,N_21929,N_24609);
or U27851 (N_27851,N_20007,N_23191);
nor U27852 (N_27852,N_21046,N_22698);
xor U27853 (N_27853,N_21088,N_20600);
xnor U27854 (N_27854,N_23883,N_21968);
and U27855 (N_27855,N_23825,N_20712);
and U27856 (N_27856,N_23182,N_21031);
nand U27857 (N_27857,N_22568,N_20280);
nand U27858 (N_27858,N_23313,N_20810);
nor U27859 (N_27859,N_21070,N_22801);
and U27860 (N_27860,N_20173,N_21639);
nand U27861 (N_27861,N_23976,N_23548);
or U27862 (N_27862,N_23180,N_20427);
nor U27863 (N_27863,N_22207,N_23220);
nand U27864 (N_27864,N_24502,N_24317);
or U27865 (N_27865,N_20803,N_24010);
nand U27866 (N_27866,N_24637,N_22928);
nor U27867 (N_27867,N_24520,N_23395);
nand U27868 (N_27868,N_21398,N_20989);
and U27869 (N_27869,N_21293,N_23414);
and U27870 (N_27870,N_22954,N_23448);
xnor U27871 (N_27871,N_24125,N_23591);
xnor U27872 (N_27872,N_23542,N_22456);
and U27873 (N_27873,N_21899,N_20256);
xor U27874 (N_27874,N_20702,N_22510);
nor U27875 (N_27875,N_21956,N_22202);
nor U27876 (N_27876,N_21503,N_22184);
nand U27877 (N_27877,N_24404,N_22434);
or U27878 (N_27878,N_24441,N_22634);
xnor U27879 (N_27879,N_21071,N_23633);
nor U27880 (N_27880,N_24345,N_22026);
nor U27881 (N_27881,N_23561,N_20631);
nand U27882 (N_27882,N_24878,N_22753);
xnor U27883 (N_27883,N_21562,N_20635);
nor U27884 (N_27884,N_20106,N_20617);
nand U27885 (N_27885,N_20518,N_22988);
and U27886 (N_27886,N_20903,N_22357);
nand U27887 (N_27887,N_24142,N_22617);
nor U27888 (N_27888,N_23710,N_21076);
xnor U27889 (N_27889,N_22795,N_21136);
xor U27890 (N_27890,N_22084,N_20556);
and U27891 (N_27891,N_22163,N_21573);
or U27892 (N_27892,N_21979,N_22859);
and U27893 (N_27893,N_23105,N_21377);
nand U27894 (N_27894,N_22511,N_22611);
nand U27895 (N_27895,N_21105,N_22184);
xor U27896 (N_27896,N_22986,N_23934);
nor U27897 (N_27897,N_24607,N_21593);
and U27898 (N_27898,N_22551,N_22782);
and U27899 (N_27899,N_23034,N_22669);
and U27900 (N_27900,N_22641,N_23389);
nand U27901 (N_27901,N_22905,N_20909);
nand U27902 (N_27902,N_23902,N_21997);
or U27903 (N_27903,N_22596,N_20519);
and U27904 (N_27904,N_20507,N_24572);
nor U27905 (N_27905,N_21245,N_24123);
or U27906 (N_27906,N_21737,N_20754);
and U27907 (N_27907,N_22066,N_21792);
nor U27908 (N_27908,N_22455,N_23830);
xnor U27909 (N_27909,N_20806,N_21094);
and U27910 (N_27910,N_24022,N_22987);
nand U27911 (N_27911,N_20228,N_23907);
nand U27912 (N_27912,N_22654,N_24594);
or U27913 (N_27913,N_24599,N_20464);
nand U27914 (N_27914,N_21346,N_21258);
nor U27915 (N_27915,N_21308,N_21234);
nand U27916 (N_27916,N_22482,N_24198);
nor U27917 (N_27917,N_21941,N_23559);
nand U27918 (N_27918,N_24632,N_23598);
nand U27919 (N_27919,N_24330,N_22994);
and U27920 (N_27920,N_22261,N_23864);
or U27921 (N_27921,N_20089,N_21206);
and U27922 (N_27922,N_21711,N_23116);
nand U27923 (N_27923,N_20012,N_22766);
or U27924 (N_27924,N_21796,N_24918);
and U27925 (N_27925,N_23513,N_24625);
or U27926 (N_27926,N_21637,N_21893);
nor U27927 (N_27927,N_23285,N_23607);
nand U27928 (N_27928,N_21448,N_22379);
or U27929 (N_27929,N_24175,N_22746);
xnor U27930 (N_27930,N_21354,N_20606);
and U27931 (N_27931,N_21575,N_22314);
xor U27932 (N_27932,N_24749,N_24270);
and U27933 (N_27933,N_20969,N_20453);
nand U27934 (N_27934,N_22911,N_22765);
xnor U27935 (N_27935,N_20252,N_21470);
nor U27936 (N_27936,N_22607,N_20645);
or U27937 (N_27937,N_21590,N_23978);
xor U27938 (N_27938,N_24892,N_21732);
nand U27939 (N_27939,N_20924,N_22264);
xor U27940 (N_27940,N_22291,N_21108);
and U27941 (N_27941,N_24630,N_22998);
or U27942 (N_27942,N_23463,N_21181);
nor U27943 (N_27943,N_24591,N_21990);
or U27944 (N_27944,N_20272,N_20971);
nand U27945 (N_27945,N_23528,N_22093);
xnor U27946 (N_27946,N_21720,N_20727);
nand U27947 (N_27947,N_20963,N_21745);
nand U27948 (N_27948,N_22256,N_23165);
nor U27949 (N_27949,N_23073,N_24875);
and U27950 (N_27950,N_24556,N_22107);
nand U27951 (N_27951,N_21636,N_23444);
nand U27952 (N_27952,N_21322,N_21562);
or U27953 (N_27953,N_22041,N_21043);
and U27954 (N_27954,N_20659,N_21093);
nand U27955 (N_27955,N_24436,N_23564);
or U27956 (N_27956,N_23655,N_22248);
nor U27957 (N_27957,N_24118,N_23060);
nand U27958 (N_27958,N_20867,N_23873);
nand U27959 (N_27959,N_24362,N_21288);
or U27960 (N_27960,N_20568,N_21370);
or U27961 (N_27961,N_20804,N_22050);
xor U27962 (N_27962,N_22726,N_22538);
xnor U27963 (N_27963,N_20201,N_21346);
nand U27964 (N_27964,N_23405,N_24430);
nand U27965 (N_27965,N_23556,N_22046);
or U27966 (N_27966,N_23620,N_24358);
nor U27967 (N_27967,N_22129,N_21170);
and U27968 (N_27968,N_21481,N_22184);
nand U27969 (N_27969,N_24996,N_24291);
nand U27970 (N_27970,N_24892,N_20457);
xnor U27971 (N_27971,N_24839,N_24007);
xor U27972 (N_27972,N_23179,N_21958);
xor U27973 (N_27973,N_21578,N_24811);
nor U27974 (N_27974,N_22213,N_23815);
xnor U27975 (N_27975,N_21426,N_24354);
nand U27976 (N_27976,N_23967,N_23798);
or U27977 (N_27977,N_23044,N_24233);
and U27978 (N_27978,N_24169,N_22692);
or U27979 (N_27979,N_24044,N_20759);
xnor U27980 (N_27980,N_20030,N_21752);
and U27981 (N_27981,N_21786,N_20954);
nor U27982 (N_27982,N_22732,N_20849);
or U27983 (N_27983,N_22485,N_24216);
nor U27984 (N_27984,N_22783,N_20481);
or U27985 (N_27985,N_21932,N_21212);
xor U27986 (N_27986,N_21366,N_20679);
or U27987 (N_27987,N_21082,N_24560);
xnor U27988 (N_27988,N_20236,N_22863);
nand U27989 (N_27989,N_24887,N_24155);
xor U27990 (N_27990,N_20227,N_24383);
xnor U27991 (N_27991,N_23915,N_20361);
nand U27992 (N_27992,N_24239,N_20379);
xnor U27993 (N_27993,N_23811,N_23125);
nand U27994 (N_27994,N_24804,N_24443);
or U27995 (N_27995,N_23067,N_21802);
xnor U27996 (N_27996,N_21938,N_23199);
xnor U27997 (N_27997,N_22370,N_22242);
nand U27998 (N_27998,N_22159,N_20073);
nor U27999 (N_27999,N_20341,N_20158);
xnor U28000 (N_28000,N_23706,N_24374);
or U28001 (N_28001,N_23968,N_23519);
or U28002 (N_28002,N_20692,N_22756);
nand U28003 (N_28003,N_22748,N_20394);
nand U28004 (N_28004,N_24140,N_23678);
and U28005 (N_28005,N_22253,N_24044);
nand U28006 (N_28006,N_24624,N_24970);
xnor U28007 (N_28007,N_24552,N_20686);
nor U28008 (N_28008,N_24253,N_24575);
nor U28009 (N_28009,N_24185,N_24242);
nand U28010 (N_28010,N_24042,N_22035);
nand U28011 (N_28011,N_23536,N_23827);
xnor U28012 (N_28012,N_24133,N_21953);
xor U28013 (N_28013,N_20533,N_22868);
and U28014 (N_28014,N_23101,N_24014);
and U28015 (N_28015,N_22825,N_20949);
xnor U28016 (N_28016,N_21106,N_22375);
and U28017 (N_28017,N_21095,N_22465);
nor U28018 (N_28018,N_23242,N_20344);
nand U28019 (N_28019,N_23863,N_24513);
and U28020 (N_28020,N_22923,N_24831);
and U28021 (N_28021,N_22107,N_23233);
and U28022 (N_28022,N_21545,N_23756);
or U28023 (N_28023,N_22636,N_20664);
nand U28024 (N_28024,N_23918,N_24129);
nand U28025 (N_28025,N_23124,N_22092);
and U28026 (N_28026,N_23675,N_22013);
and U28027 (N_28027,N_22651,N_20082);
nand U28028 (N_28028,N_23277,N_23355);
nor U28029 (N_28029,N_22517,N_21752);
and U28030 (N_28030,N_23463,N_21982);
nand U28031 (N_28031,N_21809,N_22717);
or U28032 (N_28032,N_20199,N_23982);
or U28033 (N_28033,N_21817,N_22910);
nand U28034 (N_28034,N_24283,N_21640);
xnor U28035 (N_28035,N_22088,N_24993);
nand U28036 (N_28036,N_23743,N_23009);
nor U28037 (N_28037,N_22889,N_24619);
or U28038 (N_28038,N_21500,N_24665);
or U28039 (N_28039,N_22605,N_24423);
and U28040 (N_28040,N_20998,N_23575);
or U28041 (N_28041,N_22396,N_23729);
nor U28042 (N_28042,N_21603,N_23527);
nor U28043 (N_28043,N_24898,N_21406);
or U28044 (N_28044,N_21965,N_20504);
or U28045 (N_28045,N_24275,N_24050);
nor U28046 (N_28046,N_22780,N_23003);
or U28047 (N_28047,N_24428,N_24177);
or U28048 (N_28048,N_20586,N_20958);
nor U28049 (N_28049,N_21643,N_21531);
nor U28050 (N_28050,N_20704,N_20878);
xor U28051 (N_28051,N_23200,N_20439);
xnor U28052 (N_28052,N_20394,N_23722);
nor U28053 (N_28053,N_21030,N_20925);
xnor U28054 (N_28054,N_24926,N_21079);
and U28055 (N_28055,N_22320,N_24669);
or U28056 (N_28056,N_23493,N_21096);
nand U28057 (N_28057,N_23411,N_24749);
or U28058 (N_28058,N_22130,N_24725);
nor U28059 (N_28059,N_21983,N_24881);
xnor U28060 (N_28060,N_21641,N_22631);
xor U28061 (N_28061,N_20528,N_22662);
and U28062 (N_28062,N_24884,N_24867);
nor U28063 (N_28063,N_24607,N_24431);
nand U28064 (N_28064,N_24873,N_20622);
nand U28065 (N_28065,N_22744,N_21523);
nand U28066 (N_28066,N_24270,N_20796);
nor U28067 (N_28067,N_21780,N_21440);
and U28068 (N_28068,N_22851,N_24761);
nor U28069 (N_28069,N_22800,N_23917);
nand U28070 (N_28070,N_22191,N_21904);
and U28071 (N_28071,N_21018,N_23498);
nand U28072 (N_28072,N_24313,N_22554);
nand U28073 (N_28073,N_24034,N_22862);
or U28074 (N_28074,N_22312,N_22609);
and U28075 (N_28075,N_24567,N_21897);
xor U28076 (N_28076,N_23041,N_24168);
xnor U28077 (N_28077,N_20398,N_22627);
xor U28078 (N_28078,N_23281,N_23205);
xnor U28079 (N_28079,N_20267,N_23557);
xnor U28080 (N_28080,N_20588,N_24900);
nand U28081 (N_28081,N_22645,N_20695);
and U28082 (N_28082,N_20951,N_23336);
nor U28083 (N_28083,N_23643,N_22462);
nand U28084 (N_28084,N_22515,N_22048);
nor U28085 (N_28085,N_22038,N_21963);
xor U28086 (N_28086,N_24894,N_22911);
nand U28087 (N_28087,N_20492,N_21566);
or U28088 (N_28088,N_22619,N_21349);
nand U28089 (N_28089,N_23038,N_23835);
or U28090 (N_28090,N_21477,N_23620);
nor U28091 (N_28091,N_23746,N_23771);
and U28092 (N_28092,N_23698,N_20301);
nor U28093 (N_28093,N_22676,N_24864);
or U28094 (N_28094,N_21216,N_21256);
and U28095 (N_28095,N_20517,N_23885);
xnor U28096 (N_28096,N_23253,N_23798);
xnor U28097 (N_28097,N_20149,N_20336);
nand U28098 (N_28098,N_24267,N_21495);
xnor U28099 (N_28099,N_23599,N_23564);
nand U28100 (N_28100,N_24692,N_20286);
and U28101 (N_28101,N_24434,N_24810);
nand U28102 (N_28102,N_24128,N_20037);
or U28103 (N_28103,N_22680,N_23030);
nand U28104 (N_28104,N_24898,N_20505);
nor U28105 (N_28105,N_22081,N_24116);
and U28106 (N_28106,N_21678,N_21702);
xnor U28107 (N_28107,N_24086,N_20701);
and U28108 (N_28108,N_24392,N_20300);
xor U28109 (N_28109,N_23402,N_22496);
xnor U28110 (N_28110,N_22815,N_21343);
nor U28111 (N_28111,N_20468,N_22701);
nand U28112 (N_28112,N_21944,N_22440);
and U28113 (N_28113,N_23593,N_23324);
xor U28114 (N_28114,N_23276,N_21453);
xor U28115 (N_28115,N_20576,N_24230);
nor U28116 (N_28116,N_23916,N_20775);
or U28117 (N_28117,N_22278,N_23660);
xor U28118 (N_28118,N_24815,N_24847);
xor U28119 (N_28119,N_22561,N_22542);
or U28120 (N_28120,N_24718,N_22901);
xnor U28121 (N_28121,N_21457,N_22705);
nor U28122 (N_28122,N_24513,N_21593);
nand U28123 (N_28123,N_21397,N_23347);
and U28124 (N_28124,N_22827,N_23290);
and U28125 (N_28125,N_23052,N_21142);
nand U28126 (N_28126,N_20261,N_22082);
or U28127 (N_28127,N_23031,N_20355);
xnor U28128 (N_28128,N_22807,N_20612);
nand U28129 (N_28129,N_20038,N_24430);
nand U28130 (N_28130,N_21751,N_23556);
nor U28131 (N_28131,N_23910,N_21528);
xnor U28132 (N_28132,N_21648,N_22541);
xor U28133 (N_28133,N_21227,N_22319);
nor U28134 (N_28134,N_21038,N_23385);
xnor U28135 (N_28135,N_21905,N_20512);
and U28136 (N_28136,N_21107,N_21309);
nand U28137 (N_28137,N_24666,N_24280);
nand U28138 (N_28138,N_21676,N_24571);
or U28139 (N_28139,N_20433,N_22720);
nand U28140 (N_28140,N_23305,N_20512);
and U28141 (N_28141,N_23872,N_22452);
nor U28142 (N_28142,N_23939,N_24928);
nor U28143 (N_28143,N_21097,N_21924);
xnor U28144 (N_28144,N_23778,N_21349);
or U28145 (N_28145,N_21834,N_21486);
nor U28146 (N_28146,N_24364,N_21313);
xnor U28147 (N_28147,N_24282,N_20863);
and U28148 (N_28148,N_22383,N_23915);
or U28149 (N_28149,N_24977,N_20107);
nor U28150 (N_28150,N_20292,N_23263);
and U28151 (N_28151,N_23176,N_21734);
nor U28152 (N_28152,N_21202,N_20798);
nor U28153 (N_28153,N_23405,N_22446);
nand U28154 (N_28154,N_24279,N_20736);
nand U28155 (N_28155,N_20103,N_24990);
nand U28156 (N_28156,N_24377,N_21211);
nand U28157 (N_28157,N_23601,N_20947);
xnor U28158 (N_28158,N_21040,N_20349);
nor U28159 (N_28159,N_21322,N_20354);
xor U28160 (N_28160,N_23446,N_21288);
nor U28161 (N_28161,N_20856,N_20174);
and U28162 (N_28162,N_23646,N_24925);
and U28163 (N_28163,N_24013,N_22020);
nor U28164 (N_28164,N_23830,N_20776);
or U28165 (N_28165,N_21028,N_21613);
nand U28166 (N_28166,N_22603,N_21870);
nand U28167 (N_28167,N_22542,N_22332);
nand U28168 (N_28168,N_21279,N_22929);
or U28169 (N_28169,N_22342,N_20999);
nor U28170 (N_28170,N_22910,N_23223);
or U28171 (N_28171,N_24791,N_21040);
xnor U28172 (N_28172,N_21356,N_22513);
or U28173 (N_28173,N_24051,N_22400);
xor U28174 (N_28174,N_23316,N_21921);
nor U28175 (N_28175,N_22800,N_21767);
xnor U28176 (N_28176,N_23582,N_23690);
xnor U28177 (N_28177,N_20957,N_23744);
and U28178 (N_28178,N_21095,N_24841);
nand U28179 (N_28179,N_23729,N_20018);
xor U28180 (N_28180,N_20403,N_21303);
nand U28181 (N_28181,N_23203,N_24271);
nand U28182 (N_28182,N_20610,N_23608);
or U28183 (N_28183,N_21976,N_23437);
nand U28184 (N_28184,N_22151,N_21162);
nor U28185 (N_28185,N_21068,N_24228);
nor U28186 (N_28186,N_22835,N_21539);
nand U28187 (N_28187,N_24206,N_21902);
and U28188 (N_28188,N_24702,N_23273);
nor U28189 (N_28189,N_24917,N_23185);
or U28190 (N_28190,N_20674,N_24125);
nand U28191 (N_28191,N_24854,N_21177);
nor U28192 (N_28192,N_22155,N_22319);
and U28193 (N_28193,N_20143,N_21231);
and U28194 (N_28194,N_22049,N_20422);
nand U28195 (N_28195,N_22950,N_23797);
or U28196 (N_28196,N_20859,N_22103);
or U28197 (N_28197,N_22648,N_24186);
nand U28198 (N_28198,N_22973,N_21464);
or U28199 (N_28199,N_22610,N_21489);
and U28200 (N_28200,N_20010,N_23489);
nor U28201 (N_28201,N_23169,N_22361);
xor U28202 (N_28202,N_23222,N_24319);
and U28203 (N_28203,N_24806,N_24545);
nor U28204 (N_28204,N_21684,N_24807);
or U28205 (N_28205,N_22385,N_21066);
and U28206 (N_28206,N_20821,N_20253);
nand U28207 (N_28207,N_20574,N_24226);
or U28208 (N_28208,N_20695,N_24331);
nand U28209 (N_28209,N_22190,N_21950);
or U28210 (N_28210,N_23860,N_24119);
or U28211 (N_28211,N_23435,N_23018);
or U28212 (N_28212,N_22985,N_21096);
or U28213 (N_28213,N_20013,N_22841);
or U28214 (N_28214,N_22436,N_23516);
or U28215 (N_28215,N_23039,N_22917);
xor U28216 (N_28216,N_22845,N_20190);
or U28217 (N_28217,N_24084,N_21492);
nand U28218 (N_28218,N_23990,N_22446);
or U28219 (N_28219,N_20368,N_21777);
nand U28220 (N_28220,N_22785,N_22525);
and U28221 (N_28221,N_22560,N_24921);
nand U28222 (N_28222,N_22627,N_24662);
and U28223 (N_28223,N_23301,N_21249);
nand U28224 (N_28224,N_22487,N_22734);
nand U28225 (N_28225,N_22742,N_22965);
nand U28226 (N_28226,N_21811,N_20011);
nand U28227 (N_28227,N_20891,N_23601);
and U28228 (N_28228,N_20459,N_21868);
and U28229 (N_28229,N_21618,N_23360);
nor U28230 (N_28230,N_24620,N_20260);
xnor U28231 (N_28231,N_23732,N_22063);
nor U28232 (N_28232,N_22046,N_24196);
and U28233 (N_28233,N_22853,N_22343);
or U28234 (N_28234,N_24653,N_20916);
xnor U28235 (N_28235,N_20978,N_21020);
nor U28236 (N_28236,N_23221,N_24109);
xor U28237 (N_28237,N_23412,N_24015);
xor U28238 (N_28238,N_23005,N_23799);
and U28239 (N_28239,N_24077,N_20842);
nor U28240 (N_28240,N_22961,N_23122);
xor U28241 (N_28241,N_22064,N_24856);
xor U28242 (N_28242,N_20742,N_20781);
or U28243 (N_28243,N_22174,N_22169);
or U28244 (N_28244,N_24731,N_22161);
or U28245 (N_28245,N_22797,N_21442);
nand U28246 (N_28246,N_23634,N_22418);
or U28247 (N_28247,N_22410,N_24029);
nand U28248 (N_28248,N_24036,N_24309);
nand U28249 (N_28249,N_21612,N_21639);
and U28250 (N_28250,N_22324,N_24183);
nand U28251 (N_28251,N_22888,N_20381);
nor U28252 (N_28252,N_21991,N_22518);
xnor U28253 (N_28253,N_20926,N_24449);
xnor U28254 (N_28254,N_24566,N_20949);
xor U28255 (N_28255,N_24330,N_22208);
or U28256 (N_28256,N_23225,N_24586);
nand U28257 (N_28257,N_22451,N_23364);
nor U28258 (N_28258,N_23145,N_24092);
or U28259 (N_28259,N_22465,N_24984);
or U28260 (N_28260,N_22584,N_21521);
nand U28261 (N_28261,N_23443,N_20120);
nor U28262 (N_28262,N_20141,N_21004);
xor U28263 (N_28263,N_21108,N_24783);
nand U28264 (N_28264,N_20756,N_20958);
xor U28265 (N_28265,N_20147,N_22931);
nor U28266 (N_28266,N_20611,N_23480);
or U28267 (N_28267,N_23905,N_20382);
and U28268 (N_28268,N_20745,N_24578);
nand U28269 (N_28269,N_22198,N_21801);
or U28270 (N_28270,N_20668,N_21243);
nand U28271 (N_28271,N_20048,N_24010);
xor U28272 (N_28272,N_21623,N_20467);
or U28273 (N_28273,N_22894,N_23106);
nand U28274 (N_28274,N_24676,N_21343);
xnor U28275 (N_28275,N_22677,N_21087);
nand U28276 (N_28276,N_20556,N_24485);
or U28277 (N_28277,N_20366,N_24120);
nor U28278 (N_28278,N_24051,N_24699);
xor U28279 (N_28279,N_23845,N_24391);
xor U28280 (N_28280,N_24076,N_20251);
or U28281 (N_28281,N_24579,N_23754);
nand U28282 (N_28282,N_24723,N_24382);
or U28283 (N_28283,N_22879,N_22885);
and U28284 (N_28284,N_21022,N_21858);
and U28285 (N_28285,N_20043,N_20511);
xor U28286 (N_28286,N_24810,N_24086);
and U28287 (N_28287,N_22910,N_24890);
or U28288 (N_28288,N_24194,N_22232);
xnor U28289 (N_28289,N_20867,N_24390);
or U28290 (N_28290,N_22172,N_23497);
and U28291 (N_28291,N_20806,N_20400);
or U28292 (N_28292,N_23952,N_24598);
nor U28293 (N_28293,N_21191,N_24102);
and U28294 (N_28294,N_22132,N_23128);
and U28295 (N_28295,N_20501,N_22201);
or U28296 (N_28296,N_23611,N_22697);
or U28297 (N_28297,N_20486,N_20402);
nand U28298 (N_28298,N_20483,N_23794);
nand U28299 (N_28299,N_24249,N_23021);
and U28300 (N_28300,N_23036,N_22804);
or U28301 (N_28301,N_21235,N_24104);
nor U28302 (N_28302,N_20708,N_22476);
or U28303 (N_28303,N_23810,N_22337);
and U28304 (N_28304,N_23691,N_20566);
nand U28305 (N_28305,N_20313,N_21244);
nor U28306 (N_28306,N_20674,N_24986);
nand U28307 (N_28307,N_20223,N_21626);
nor U28308 (N_28308,N_24485,N_24373);
nor U28309 (N_28309,N_20807,N_21591);
xor U28310 (N_28310,N_21315,N_21762);
xnor U28311 (N_28311,N_23505,N_21049);
nand U28312 (N_28312,N_21432,N_22032);
nand U28313 (N_28313,N_21016,N_24868);
nand U28314 (N_28314,N_23245,N_21972);
and U28315 (N_28315,N_22814,N_20055);
and U28316 (N_28316,N_23453,N_20172);
xnor U28317 (N_28317,N_20573,N_24854);
nor U28318 (N_28318,N_21061,N_24455);
nor U28319 (N_28319,N_21502,N_24939);
xor U28320 (N_28320,N_20627,N_20104);
nor U28321 (N_28321,N_23256,N_22262);
nand U28322 (N_28322,N_22554,N_22149);
nor U28323 (N_28323,N_20794,N_20485);
nand U28324 (N_28324,N_23309,N_20759);
nand U28325 (N_28325,N_24855,N_22510);
nor U28326 (N_28326,N_24496,N_23937);
nor U28327 (N_28327,N_21570,N_20853);
or U28328 (N_28328,N_21719,N_23677);
or U28329 (N_28329,N_24557,N_21355);
nand U28330 (N_28330,N_23200,N_21935);
or U28331 (N_28331,N_20456,N_23391);
nor U28332 (N_28332,N_22332,N_24139);
and U28333 (N_28333,N_21208,N_23837);
nor U28334 (N_28334,N_22942,N_20255);
and U28335 (N_28335,N_24090,N_23265);
xnor U28336 (N_28336,N_21084,N_20990);
xnor U28337 (N_28337,N_24083,N_21188);
nor U28338 (N_28338,N_21566,N_24271);
xor U28339 (N_28339,N_24811,N_22755);
nor U28340 (N_28340,N_21190,N_21634);
or U28341 (N_28341,N_21891,N_24258);
nand U28342 (N_28342,N_20621,N_22702);
nor U28343 (N_28343,N_20238,N_21813);
or U28344 (N_28344,N_23090,N_20400);
xor U28345 (N_28345,N_20143,N_20862);
xor U28346 (N_28346,N_23240,N_20846);
and U28347 (N_28347,N_20607,N_24956);
xor U28348 (N_28348,N_23968,N_20879);
xnor U28349 (N_28349,N_24018,N_20907);
nor U28350 (N_28350,N_22752,N_21072);
nand U28351 (N_28351,N_24332,N_22035);
xor U28352 (N_28352,N_24108,N_24110);
nor U28353 (N_28353,N_24782,N_24507);
and U28354 (N_28354,N_23905,N_23362);
nor U28355 (N_28355,N_21446,N_22193);
and U28356 (N_28356,N_20329,N_23037);
nor U28357 (N_28357,N_23894,N_20002);
xnor U28358 (N_28358,N_21039,N_22134);
nand U28359 (N_28359,N_24845,N_24153);
and U28360 (N_28360,N_20273,N_20448);
nand U28361 (N_28361,N_24681,N_20703);
nand U28362 (N_28362,N_20090,N_24062);
nor U28363 (N_28363,N_23692,N_24261);
or U28364 (N_28364,N_23881,N_24368);
and U28365 (N_28365,N_23677,N_21062);
xor U28366 (N_28366,N_22544,N_21564);
nand U28367 (N_28367,N_21737,N_21402);
xor U28368 (N_28368,N_22380,N_21400);
nor U28369 (N_28369,N_23382,N_20374);
and U28370 (N_28370,N_24213,N_20792);
and U28371 (N_28371,N_21480,N_23213);
and U28372 (N_28372,N_20122,N_22889);
nand U28373 (N_28373,N_21133,N_20668);
nand U28374 (N_28374,N_20689,N_21621);
nor U28375 (N_28375,N_22070,N_22535);
xnor U28376 (N_28376,N_24947,N_23441);
and U28377 (N_28377,N_22782,N_20695);
nor U28378 (N_28378,N_20783,N_24972);
nand U28379 (N_28379,N_22149,N_22960);
xor U28380 (N_28380,N_23956,N_24224);
and U28381 (N_28381,N_23229,N_20222);
nor U28382 (N_28382,N_24586,N_21684);
nor U28383 (N_28383,N_21078,N_20498);
nand U28384 (N_28384,N_22288,N_21943);
or U28385 (N_28385,N_24805,N_24284);
or U28386 (N_28386,N_21413,N_21987);
nor U28387 (N_28387,N_21095,N_22641);
nand U28388 (N_28388,N_21617,N_23402);
nand U28389 (N_28389,N_21418,N_21117);
nand U28390 (N_28390,N_24685,N_23390);
nand U28391 (N_28391,N_21880,N_23341);
xor U28392 (N_28392,N_21524,N_21086);
or U28393 (N_28393,N_21720,N_22103);
nor U28394 (N_28394,N_24468,N_23241);
nand U28395 (N_28395,N_21726,N_21218);
nand U28396 (N_28396,N_21762,N_21482);
or U28397 (N_28397,N_23732,N_22091);
xor U28398 (N_28398,N_24777,N_24440);
nor U28399 (N_28399,N_20373,N_21943);
and U28400 (N_28400,N_23359,N_21585);
nor U28401 (N_28401,N_20610,N_24204);
and U28402 (N_28402,N_21869,N_23607);
or U28403 (N_28403,N_23282,N_22274);
or U28404 (N_28404,N_20578,N_21901);
or U28405 (N_28405,N_20977,N_20112);
nand U28406 (N_28406,N_24893,N_20154);
nand U28407 (N_28407,N_23230,N_20651);
and U28408 (N_28408,N_20763,N_20199);
nand U28409 (N_28409,N_23476,N_21274);
nor U28410 (N_28410,N_21751,N_21612);
xnor U28411 (N_28411,N_23629,N_21666);
nand U28412 (N_28412,N_20376,N_20438);
or U28413 (N_28413,N_22493,N_24207);
xor U28414 (N_28414,N_21084,N_23203);
and U28415 (N_28415,N_23370,N_20203);
nor U28416 (N_28416,N_22895,N_23002);
xor U28417 (N_28417,N_24381,N_23131);
xnor U28418 (N_28418,N_24708,N_24792);
or U28419 (N_28419,N_23587,N_22018);
and U28420 (N_28420,N_23948,N_22208);
or U28421 (N_28421,N_22357,N_20379);
and U28422 (N_28422,N_23391,N_22327);
or U28423 (N_28423,N_20837,N_20378);
nor U28424 (N_28424,N_24723,N_23125);
and U28425 (N_28425,N_22386,N_22732);
nand U28426 (N_28426,N_20684,N_22954);
nand U28427 (N_28427,N_21519,N_24672);
xnor U28428 (N_28428,N_21099,N_23034);
nor U28429 (N_28429,N_24547,N_21318);
xor U28430 (N_28430,N_23990,N_20522);
and U28431 (N_28431,N_22163,N_22385);
nand U28432 (N_28432,N_20563,N_22220);
or U28433 (N_28433,N_21078,N_24121);
xor U28434 (N_28434,N_23081,N_21795);
and U28435 (N_28435,N_24478,N_24241);
xnor U28436 (N_28436,N_23257,N_21564);
nand U28437 (N_28437,N_20869,N_24129);
nand U28438 (N_28438,N_24003,N_22721);
nor U28439 (N_28439,N_24153,N_24920);
nor U28440 (N_28440,N_20054,N_22007);
xor U28441 (N_28441,N_23661,N_23003);
or U28442 (N_28442,N_21217,N_23230);
nor U28443 (N_28443,N_21353,N_20242);
nor U28444 (N_28444,N_24378,N_21298);
xor U28445 (N_28445,N_20619,N_23536);
and U28446 (N_28446,N_24545,N_21854);
nand U28447 (N_28447,N_21151,N_23591);
and U28448 (N_28448,N_21090,N_22600);
nand U28449 (N_28449,N_24808,N_23080);
or U28450 (N_28450,N_21754,N_23835);
nand U28451 (N_28451,N_21968,N_22908);
or U28452 (N_28452,N_21985,N_24931);
and U28453 (N_28453,N_22211,N_20095);
nand U28454 (N_28454,N_20977,N_24177);
and U28455 (N_28455,N_21020,N_23865);
nand U28456 (N_28456,N_22338,N_20443);
nand U28457 (N_28457,N_22140,N_24987);
or U28458 (N_28458,N_20519,N_21898);
nand U28459 (N_28459,N_20890,N_21041);
nor U28460 (N_28460,N_23838,N_22700);
nand U28461 (N_28461,N_21289,N_23714);
nand U28462 (N_28462,N_23196,N_24927);
and U28463 (N_28463,N_22038,N_23305);
xor U28464 (N_28464,N_22008,N_21391);
xnor U28465 (N_28465,N_20971,N_21645);
xor U28466 (N_28466,N_23142,N_20255);
nor U28467 (N_28467,N_23015,N_23295);
nor U28468 (N_28468,N_20583,N_24017);
nand U28469 (N_28469,N_21471,N_20344);
and U28470 (N_28470,N_20807,N_23152);
and U28471 (N_28471,N_21545,N_20226);
xnor U28472 (N_28472,N_23141,N_24721);
xnor U28473 (N_28473,N_20005,N_20278);
xor U28474 (N_28474,N_23508,N_20100);
and U28475 (N_28475,N_22199,N_21063);
and U28476 (N_28476,N_20721,N_21942);
and U28477 (N_28477,N_21538,N_21528);
nor U28478 (N_28478,N_21235,N_24023);
nand U28479 (N_28479,N_23030,N_20809);
xnor U28480 (N_28480,N_22835,N_24351);
or U28481 (N_28481,N_20329,N_22982);
nand U28482 (N_28482,N_24885,N_23880);
nor U28483 (N_28483,N_22846,N_21113);
nor U28484 (N_28484,N_23957,N_24714);
or U28485 (N_28485,N_23934,N_22060);
nor U28486 (N_28486,N_20040,N_23805);
nor U28487 (N_28487,N_22618,N_21669);
xor U28488 (N_28488,N_21834,N_21250);
and U28489 (N_28489,N_21689,N_21271);
and U28490 (N_28490,N_22440,N_24964);
and U28491 (N_28491,N_20702,N_24332);
or U28492 (N_28492,N_23349,N_23671);
and U28493 (N_28493,N_20494,N_23675);
nor U28494 (N_28494,N_21057,N_22197);
and U28495 (N_28495,N_24414,N_23499);
xor U28496 (N_28496,N_20698,N_22220);
or U28497 (N_28497,N_21595,N_24363);
nor U28498 (N_28498,N_22995,N_24559);
nor U28499 (N_28499,N_23514,N_20156);
and U28500 (N_28500,N_22936,N_21256);
nor U28501 (N_28501,N_22630,N_21288);
nor U28502 (N_28502,N_23769,N_20720);
and U28503 (N_28503,N_23192,N_21115);
or U28504 (N_28504,N_23926,N_20647);
and U28505 (N_28505,N_21930,N_21010);
nor U28506 (N_28506,N_23095,N_22893);
xor U28507 (N_28507,N_22864,N_20211);
nand U28508 (N_28508,N_20285,N_21038);
and U28509 (N_28509,N_21148,N_21919);
and U28510 (N_28510,N_24891,N_21805);
xnor U28511 (N_28511,N_22767,N_21352);
or U28512 (N_28512,N_20527,N_24838);
and U28513 (N_28513,N_22639,N_21909);
and U28514 (N_28514,N_22851,N_21950);
xnor U28515 (N_28515,N_21039,N_23009);
xor U28516 (N_28516,N_24851,N_21596);
and U28517 (N_28517,N_20245,N_22082);
or U28518 (N_28518,N_23566,N_22240);
and U28519 (N_28519,N_22387,N_20188);
or U28520 (N_28520,N_21105,N_21245);
nand U28521 (N_28521,N_24247,N_20532);
xnor U28522 (N_28522,N_23618,N_20999);
nor U28523 (N_28523,N_20622,N_20292);
xor U28524 (N_28524,N_20059,N_22784);
or U28525 (N_28525,N_20733,N_20486);
and U28526 (N_28526,N_22360,N_20515);
or U28527 (N_28527,N_20745,N_20347);
nor U28528 (N_28528,N_23022,N_24921);
xor U28529 (N_28529,N_22122,N_24696);
xor U28530 (N_28530,N_20843,N_22008);
or U28531 (N_28531,N_23488,N_21359);
and U28532 (N_28532,N_21336,N_22956);
and U28533 (N_28533,N_23034,N_20483);
xor U28534 (N_28534,N_21216,N_22232);
xor U28535 (N_28535,N_24360,N_23940);
and U28536 (N_28536,N_23264,N_23566);
nand U28537 (N_28537,N_20953,N_22453);
xor U28538 (N_28538,N_24621,N_21395);
nor U28539 (N_28539,N_24364,N_23306);
and U28540 (N_28540,N_21791,N_24135);
and U28541 (N_28541,N_24789,N_20568);
nand U28542 (N_28542,N_21407,N_21171);
and U28543 (N_28543,N_22746,N_24768);
and U28544 (N_28544,N_21346,N_23299);
nand U28545 (N_28545,N_22589,N_24105);
nor U28546 (N_28546,N_22766,N_24916);
or U28547 (N_28547,N_22928,N_20221);
and U28548 (N_28548,N_20780,N_22541);
nor U28549 (N_28549,N_22322,N_23570);
nand U28550 (N_28550,N_21017,N_21959);
xor U28551 (N_28551,N_23908,N_20272);
xor U28552 (N_28552,N_24300,N_24991);
nand U28553 (N_28553,N_22868,N_20288);
and U28554 (N_28554,N_24905,N_24676);
nand U28555 (N_28555,N_21592,N_21111);
and U28556 (N_28556,N_21896,N_21781);
nand U28557 (N_28557,N_22250,N_23753);
or U28558 (N_28558,N_23642,N_22117);
xnor U28559 (N_28559,N_22808,N_20914);
nor U28560 (N_28560,N_20275,N_20135);
or U28561 (N_28561,N_24056,N_21934);
and U28562 (N_28562,N_24013,N_22645);
nand U28563 (N_28563,N_24118,N_21533);
and U28564 (N_28564,N_23456,N_20532);
and U28565 (N_28565,N_21908,N_21312);
and U28566 (N_28566,N_24445,N_20348);
and U28567 (N_28567,N_20401,N_22225);
and U28568 (N_28568,N_24593,N_23229);
and U28569 (N_28569,N_23672,N_21545);
and U28570 (N_28570,N_24765,N_20608);
xnor U28571 (N_28571,N_21428,N_22212);
nor U28572 (N_28572,N_22656,N_22488);
and U28573 (N_28573,N_23756,N_20217);
xor U28574 (N_28574,N_20221,N_23341);
xor U28575 (N_28575,N_24160,N_23726);
and U28576 (N_28576,N_24690,N_22503);
and U28577 (N_28577,N_24339,N_23719);
nor U28578 (N_28578,N_21812,N_24323);
and U28579 (N_28579,N_22154,N_24987);
xnor U28580 (N_28580,N_23566,N_21154);
nand U28581 (N_28581,N_21619,N_21180);
nor U28582 (N_28582,N_20616,N_20307);
nor U28583 (N_28583,N_21456,N_22873);
nor U28584 (N_28584,N_20120,N_22178);
nor U28585 (N_28585,N_23130,N_24911);
nor U28586 (N_28586,N_21662,N_20228);
and U28587 (N_28587,N_23497,N_23243);
nand U28588 (N_28588,N_20021,N_20234);
nor U28589 (N_28589,N_21336,N_21077);
xor U28590 (N_28590,N_21478,N_21114);
xor U28591 (N_28591,N_20328,N_20857);
xor U28592 (N_28592,N_22076,N_21763);
or U28593 (N_28593,N_24860,N_23310);
and U28594 (N_28594,N_20473,N_23659);
and U28595 (N_28595,N_24214,N_23743);
or U28596 (N_28596,N_24378,N_22073);
xnor U28597 (N_28597,N_22504,N_21479);
xnor U28598 (N_28598,N_21249,N_24469);
nand U28599 (N_28599,N_23460,N_24341);
nor U28600 (N_28600,N_24529,N_21759);
xnor U28601 (N_28601,N_24562,N_22132);
or U28602 (N_28602,N_24730,N_23744);
xor U28603 (N_28603,N_21457,N_24252);
nand U28604 (N_28604,N_24888,N_23727);
nor U28605 (N_28605,N_23255,N_23911);
xor U28606 (N_28606,N_20598,N_23236);
nor U28607 (N_28607,N_20797,N_24365);
or U28608 (N_28608,N_20320,N_20216);
xnor U28609 (N_28609,N_24100,N_22099);
nor U28610 (N_28610,N_21360,N_22762);
xor U28611 (N_28611,N_21093,N_24625);
or U28612 (N_28612,N_20452,N_21525);
nand U28613 (N_28613,N_20436,N_20730);
or U28614 (N_28614,N_24037,N_24872);
and U28615 (N_28615,N_23066,N_24496);
xor U28616 (N_28616,N_20876,N_20135);
and U28617 (N_28617,N_24718,N_24237);
and U28618 (N_28618,N_22346,N_20254);
or U28619 (N_28619,N_20751,N_21408);
and U28620 (N_28620,N_22717,N_24580);
nor U28621 (N_28621,N_22816,N_20495);
nor U28622 (N_28622,N_20406,N_21503);
xor U28623 (N_28623,N_24334,N_20112);
and U28624 (N_28624,N_23344,N_23844);
and U28625 (N_28625,N_23465,N_24233);
xnor U28626 (N_28626,N_22512,N_23374);
xnor U28627 (N_28627,N_23051,N_23358);
nor U28628 (N_28628,N_23419,N_22816);
nand U28629 (N_28629,N_23965,N_23944);
and U28630 (N_28630,N_20373,N_23899);
nand U28631 (N_28631,N_21306,N_22239);
nor U28632 (N_28632,N_23163,N_23629);
or U28633 (N_28633,N_20898,N_20938);
nand U28634 (N_28634,N_21788,N_23470);
and U28635 (N_28635,N_24771,N_20091);
xor U28636 (N_28636,N_22490,N_23855);
nand U28637 (N_28637,N_22160,N_22391);
and U28638 (N_28638,N_22620,N_23763);
and U28639 (N_28639,N_21250,N_21227);
and U28640 (N_28640,N_23307,N_22346);
nand U28641 (N_28641,N_21711,N_20901);
xnor U28642 (N_28642,N_24927,N_21467);
nand U28643 (N_28643,N_22148,N_20309);
or U28644 (N_28644,N_24933,N_20717);
or U28645 (N_28645,N_20276,N_20137);
and U28646 (N_28646,N_21339,N_23265);
xor U28647 (N_28647,N_24778,N_22755);
nor U28648 (N_28648,N_20930,N_24698);
xor U28649 (N_28649,N_22299,N_23836);
and U28650 (N_28650,N_23953,N_23740);
or U28651 (N_28651,N_21288,N_21947);
xor U28652 (N_28652,N_20300,N_20496);
xnor U28653 (N_28653,N_24133,N_21099);
and U28654 (N_28654,N_21187,N_20331);
nand U28655 (N_28655,N_20177,N_23392);
nor U28656 (N_28656,N_21140,N_20158);
nand U28657 (N_28657,N_22519,N_23621);
nor U28658 (N_28658,N_21941,N_21610);
nand U28659 (N_28659,N_21095,N_20848);
nand U28660 (N_28660,N_23134,N_24764);
xor U28661 (N_28661,N_24913,N_20227);
nand U28662 (N_28662,N_24630,N_22348);
and U28663 (N_28663,N_24614,N_20687);
and U28664 (N_28664,N_23859,N_24056);
and U28665 (N_28665,N_22026,N_21459);
and U28666 (N_28666,N_23457,N_23720);
nand U28667 (N_28667,N_20652,N_20632);
nor U28668 (N_28668,N_20821,N_21410);
nand U28669 (N_28669,N_24283,N_21142);
or U28670 (N_28670,N_23035,N_20723);
and U28671 (N_28671,N_20122,N_23797);
nor U28672 (N_28672,N_24799,N_24714);
nand U28673 (N_28673,N_24090,N_20059);
or U28674 (N_28674,N_22232,N_24278);
and U28675 (N_28675,N_23355,N_24049);
or U28676 (N_28676,N_23637,N_24546);
nand U28677 (N_28677,N_23481,N_20637);
nor U28678 (N_28678,N_24024,N_23195);
and U28679 (N_28679,N_21477,N_21496);
nor U28680 (N_28680,N_23985,N_24657);
nand U28681 (N_28681,N_24437,N_22570);
nand U28682 (N_28682,N_23636,N_22772);
or U28683 (N_28683,N_23433,N_24230);
nor U28684 (N_28684,N_23673,N_22324);
nand U28685 (N_28685,N_23372,N_20937);
nor U28686 (N_28686,N_22878,N_20666);
or U28687 (N_28687,N_23302,N_23733);
nor U28688 (N_28688,N_20326,N_22642);
xnor U28689 (N_28689,N_23303,N_24659);
nand U28690 (N_28690,N_22110,N_23575);
or U28691 (N_28691,N_23650,N_23820);
xor U28692 (N_28692,N_21585,N_24603);
nand U28693 (N_28693,N_21521,N_23580);
and U28694 (N_28694,N_21682,N_20472);
nor U28695 (N_28695,N_20001,N_24618);
or U28696 (N_28696,N_20825,N_22662);
or U28697 (N_28697,N_22827,N_23319);
or U28698 (N_28698,N_24090,N_24510);
nor U28699 (N_28699,N_21842,N_23522);
or U28700 (N_28700,N_23893,N_22528);
xnor U28701 (N_28701,N_22333,N_24884);
and U28702 (N_28702,N_21136,N_22717);
and U28703 (N_28703,N_20822,N_20757);
or U28704 (N_28704,N_20394,N_23256);
nand U28705 (N_28705,N_21396,N_22840);
or U28706 (N_28706,N_20244,N_23676);
or U28707 (N_28707,N_23025,N_23794);
nor U28708 (N_28708,N_24641,N_24336);
nor U28709 (N_28709,N_21590,N_20040);
and U28710 (N_28710,N_24941,N_20486);
nand U28711 (N_28711,N_22484,N_23044);
or U28712 (N_28712,N_23138,N_21572);
xor U28713 (N_28713,N_21126,N_24994);
and U28714 (N_28714,N_21093,N_20207);
and U28715 (N_28715,N_23906,N_22183);
xor U28716 (N_28716,N_21157,N_23462);
xnor U28717 (N_28717,N_24992,N_24681);
and U28718 (N_28718,N_20292,N_21979);
xor U28719 (N_28719,N_20587,N_24898);
or U28720 (N_28720,N_23100,N_20122);
nand U28721 (N_28721,N_23379,N_24239);
nand U28722 (N_28722,N_23807,N_22158);
nand U28723 (N_28723,N_24761,N_21333);
and U28724 (N_28724,N_23633,N_20536);
or U28725 (N_28725,N_21236,N_21663);
and U28726 (N_28726,N_21174,N_23133);
xor U28727 (N_28727,N_20718,N_21590);
nand U28728 (N_28728,N_20447,N_24541);
or U28729 (N_28729,N_22841,N_22550);
and U28730 (N_28730,N_21717,N_22045);
and U28731 (N_28731,N_21298,N_24482);
or U28732 (N_28732,N_22026,N_24628);
nand U28733 (N_28733,N_24328,N_21727);
nand U28734 (N_28734,N_21562,N_23083);
or U28735 (N_28735,N_20027,N_21237);
and U28736 (N_28736,N_22269,N_23466);
nor U28737 (N_28737,N_20998,N_24168);
xnor U28738 (N_28738,N_24366,N_22850);
nor U28739 (N_28739,N_21527,N_24260);
nand U28740 (N_28740,N_24229,N_24575);
and U28741 (N_28741,N_24377,N_20292);
nor U28742 (N_28742,N_23803,N_22811);
xor U28743 (N_28743,N_20094,N_20212);
and U28744 (N_28744,N_23795,N_21017);
xor U28745 (N_28745,N_21324,N_23287);
nor U28746 (N_28746,N_21942,N_21837);
nor U28747 (N_28747,N_22913,N_23837);
or U28748 (N_28748,N_21150,N_24291);
and U28749 (N_28749,N_22656,N_23967);
xor U28750 (N_28750,N_23696,N_23545);
nand U28751 (N_28751,N_21157,N_23595);
nor U28752 (N_28752,N_21738,N_21472);
xnor U28753 (N_28753,N_24367,N_20743);
nor U28754 (N_28754,N_23519,N_24169);
or U28755 (N_28755,N_23743,N_20604);
or U28756 (N_28756,N_22507,N_23072);
xnor U28757 (N_28757,N_20191,N_20055);
xnor U28758 (N_28758,N_22944,N_23290);
nand U28759 (N_28759,N_22306,N_23636);
nor U28760 (N_28760,N_23240,N_21411);
or U28761 (N_28761,N_24119,N_24173);
and U28762 (N_28762,N_22772,N_24123);
nand U28763 (N_28763,N_24013,N_21661);
and U28764 (N_28764,N_20848,N_23017);
nand U28765 (N_28765,N_22737,N_21353);
xor U28766 (N_28766,N_22446,N_22003);
and U28767 (N_28767,N_22261,N_23663);
xnor U28768 (N_28768,N_22508,N_21585);
xor U28769 (N_28769,N_20433,N_23609);
nor U28770 (N_28770,N_21767,N_22167);
or U28771 (N_28771,N_21893,N_20294);
and U28772 (N_28772,N_21165,N_22957);
nor U28773 (N_28773,N_22341,N_20920);
nand U28774 (N_28774,N_22937,N_21525);
nor U28775 (N_28775,N_24490,N_21405);
xor U28776 (N_28776,N_22052,N_23063);
xor U28777 (N_28777,N_20130,N_23114);
and U28778 (N_28778,N_20119,N_23207);
nand U28779 (N_28779,N_23282,N_23484);
nor U28780 (N_28780,N_23639,N_23402);
and U28781 (N_28781,N_21821,N_20851);
nand U28782 (N_28782,N_24373,N_21233);
and U28783 (N_28783,N_22161,N_22071);
nand U28784 (N_28784,N_20194,N_20994);
and U28785 (N_28785,N_21666,N_24214);
and U28786 (N_28786,N_20945,N_24136);
nor U28787 (N_28787,N_24859,N_22230);
xor U28788 (N_28788,N_22909,N_24448);
and U28789 (N_28789,N_22307,N_23810);
and U28790 (N_28790,N_22535,N_20280);
nand U28791 (N_28791,N_21650,N_20119);
and U28792 (N_28792,N_21288,N_23650);
or U28793 (N_28793,N_20793,N_24419);
or U28794 (N_28794,N_24508,N_20341);
and U28795 (N_28795,N_21671,N_22157);
nand U28796 (N_28796,N_23174,N_21978);
and U28797 (N_28797,N_20176,N_21131);
nor U28798 (N_28798,N_23135,N_24178);
and U28799 (N_28799,N_21144,N_23316);
or U28800 (N_28800,N_24364,N_23273);
nor U28801 (N_28801,N_24611,N_21757);
and U28802 (N_28802,N_24067,N_22581);
and U28803 (N_28803,N_24304,N_24123);
or U28804 (N_28804,N_23518,N_24792);
nor U28805 (N_28805,N_22064,N_23036);
or U28806 (N_28806,N_24053,N_23584);
xor U28807 (N_28807,N_24689,N_21005);
or U28808 (N_28808,N_24747,N_22785);
xor U28809 (N_28809,N_21869,N_21993);
or U28810 (N_28810,N_24397,N_20130);
and U28811 (N_28811,N_20834,N_24485);
or U28812 (N_28812,N_22803,N_23424);
and U28813 (N_28813,N_24991,N_23410);
nand U28814 (N_28814,N_22982,N_20010);
nor U28815 (N_28815,N_21792,N_24116);
nor U28816 (N_28816,N_20723,N_20426);
and U28817 (N_28817,N_20872,N_24167);
nand U28818 (N_28818,N_24131,N_20599);
and U28819 (N_28819,N_23683,N_21755);
and U28820 (N_28820,N_23010,N_21321);
nor U28821 (N_28821,N_23974,N_24730);
xor U28822 (N_28822,N_20508,N_24977);
nor U28823 (N_28823,N_20175,N_20688);
and U28824 (N_28824,N_20113,N_21402);
or U28825 (N_28825,N_20349,N_24971);
and U28826 (N_28826,N_20778,N_23203);
and U28827 (N_28827,N_22680,N_21828);
or U28828 (N_28828,N_21405,N_20336);
or U28829 (N_28829,N_20851,N_22752);
or U28830 (N_28830,N_23810,N_21649);
nor U28831 (N_28831,N_23161,N_21123);
nor U28832 (N_28832,N_21031,N_21557);
and U28833 (N_28833,N_20514,N_20333);
or U28834 (N_28834,N_22783,N_20905);
nor U28835 (N_28835,N_20405,N_20975);
xnor U28836 (N_28836,N_24654,N_22233);
nand U28837 (N_28837,N_23552,N_22436);
nand U28838 (N_28838,N_23026,N_24139);
nand U28839 (N_28839,N_23909,N_20971);
and U28840 (N_28840,N_20582,N_21853);
or U28841 (N_28841,N_21242,N_20550);
and U28842 (N_28842,N_24635,N_21238);
xnor U28843 (N_28843,N_21731,N_24985);
xnor U28844 (N_28844,N_22512,N_23682);
xnor U28845 (N_28845,N_21578,N_24491);
or U28846 (N_28846,N_21421,N_21850);
or U28847 (N_28847,N_21819,N_24173);
nor U28848 (N_28848,N_21996,N_21317);
or U28849 (N_28849,N_20710,N_22685);
or U28850 (N_28850,N_20519,N_23028);
or U28851 (N_28851,N_22233,N_24319);
xnor U28852 (N_28852,N_20056,N_24750);
nand U28853 (N_28853,N_24703,N_24208);
nand U28854 (N_28854,N_24543,N_23082);
and U28855 (N_28855,N_23160,N_20481);
and U28856 (N_28856,N_21440,N_20786);
or U28857 (N_28857,N_24557,N_23411);
nor U28858 (N_28858,N_21791,N_24889);
xor U28859 (N_28859,N_21998,N_23662);
nand U28860 (N_28860,N_22291,N_23803);
nand U28861 (N_28861,N_20357,N_22529);
or U28862 (N_28862,N_20153,N_23641);
nand U28863 (N_28863,N_23171,N_22424);
nand U28864 (N_28864,N_20692,N_20685);
or U28865 (N_28865,N_21032,N_21485);
or U28866 (N_28866,N_20189,N_23472);
nand U28867 (N_28867,N_20511,N_24144);
xor U28868 (N_28868,N_23945,N_20336);
and U28869 (N_28869,N_24282,N_23624);
or U28870 (N_28870,N_20319,N_23337);
and U28871 (N_28871,N_20713,N_22010);
nand U28872 (N_28872,N_23617,N_20605);
and U28873 (N_28873,N_24300,N_21914);
xor U28874 (N_28874,N_21891,N_23128);
nor U28875 (N_28875,N_24951,N_24027);
xnor U28876 (N_28876,N_23462,N_22976);
or U28877 (N_28877,N_21684,N_21295);
and U28878 (N_28878,N_23181,N_21904);
and U28879 (N_28879,N_24701,N_22231);
and U28880 (N_28880,N_24549,N_23192);
nor U28881 (N_28881,N_24155,N_24952);
nor U28882 (N_28882,N_21416,N_24067);
nor U28883 (N_28883,N_20871,N_24804);
or U28884 (N_28884,N_20001,N_21685);
and U28885 (N_28885,N_24936,N_21888);
nand U28886 (N_28886,N_22597,N_22754);
or U28887 (N_28887,N_24159,N_22014);
nand U28888 (N_28888,N_20566,N_20886);
and U28889 (N_28889,N_23942,N_22529);
nand U28890 (N_28890,N_23603,N_22027);
and U28891 (N_28891,N_23726,N_24872);
nand U28892 (N_28892,N_24834,N_24763);
or U28893 (N_28893,N_20039,N_22731);
and U28894 (N_28894,N_21532,N_21494);
or U28895 (N_28895,N_22479,N_22078);
nand U28896 (N_28896,N_20260,N_20854);
nor U28897 (N_28897,N_22986,N_23435);
nand U28898 (N_28898,N_22336,N_21388);
and U28899 (N_28899,N_24888,N_21570);
nor U28900 (N_28900,N_23098,N_23754);
nand U28901 (N_28901,N_24476,N_24706);
and U28902 (N_28902,N_22404,N_23932);
nor U28903 (N_28903,N_21985,N_22508);
and U28904 (N_28904,N_21520,N_23227);
nand U28905 (N_28905,N_24845,N_24844);
and U28906 (N_28906,N_20337,N_23531);
and U28907 (N_28907,N_23427,N_23591);
nand U28908 (N_28908,N_21762,N_24979);
or U28909 (N_28909,N_20950,N_20784);
nand U28910 (N_28910,N_22002,N_23065);
nand U28911 (N_28911,N_24971,N_21271);
and U28912 (N_28912,N_22708,N_23003);
nor U28913 (N_28913,N_24242,N_21406);
xor U28914 (N_28914,N_23719,N_21579);
and U28915 (N_28915,N_24199,N_23097);
or U28916 (N_28916,N_21484,N_24674);
and U28917 (N_28917,N_20017,N_22576);
nor U28918 (N_28918,N_22339,N_20621);
xnor U28919 (N_28919,N_22229,N_23965);
nor U28920 (N_28920,N_22697,N_20220);
nor U28921 (N_28921,N_20407,N_23385);
xnor U28922 (N_28922,N_22764,N_24641);
and U28923 (N_28923,N_20462,N_24710);
xnor U28924 (N_28924,N_24256,N_24197);
nor U28925 (N_28925,N_23148,N_23996);
nand U28926 (N_28926,N_24952,N_23316);
xnor U28927 (N_28927,N_22317,N_20800);
and U28928 (N_28928,N_21924,N_23683);
nand U28929 (N_28929,N_24700,N_20045);
and U28930 (N_28930,N_20213,N_21971);
nand U28931 (N_28931,N_23618,N_21796);
and U28932 (N_28932,N_23967,N_23602);
nand U28933 (N_28933,N_22318,N_22548);
or U28934 (N_28934,N_20644,N_24193);
xnor U28935 (N_28935,N_23988,N_22927);
xor U28936 (N_28936,N_22651,N_21832);
xnor U28937 (N_28937,N_20168,N_24864);
and U28938 (N_28938,N_21418,N_23480);
xnor U28939 (N_28939,N_20504,N_21931);
and U28940 (N_28940,N_22286,N_20559);
or U28941 (N_28941,N_24937,N_24016);
nand U28942 (N_28942,N_23561,N_23073);
or U28943 (N_28943,N_22427,N_22918);
nand U28944 (N_28944,N_22760,N_24107);
and U28945 (N_28945,N_23139,N_20891);
or U28946 (N_28946,N_21218,N_23473);
and U28947 (N_28947,N_23369,N_21471);
xor U28948 (N_28948,N_21093,N_24801);
nand U28949 (N_28949,N_24983,N_22386);
or U28950 (N_28950,N_23025,N_24771);
and U28951 (N_28951,N_22686,N_22579);
nand U28952 (N_28952,N_23072,N_24673);
xnor U28953 (N_28953,N_22940,N_22345);
xor U28954 (N_28954,N_20789,N_22016);
xnor U28955 (N_28955,N_24156,N_24747);
or U28956 (N_28956,N_23572,N_21346);
and U28957 (N_28957,N_22188,N_20750);
nand U28958 (N_28958,N_21284,N_20578);
or U28959 (N_28959,N_21223,N_23937);
nand U28960 (N_28960,N_20285,N_22440);
nand U28961 (N_28961,N_21710,N_20068);
xnor U28962 (N_28962,N_20183,N_22546);
or U28963 (N_28963,N_24346,N_20167);
nor U28964 (N_28964,N_20872,N_22404);
nand U28965 (N_28965,N_20649,N_23623);
or U28966 (N_28966,N_22637,N_22252);
and U28967 (N_28967,N_24667,N_21225);
xnor U28968 (N_28968,N_24560,N_23108);
nor U28969 (N_28969,N_22911,N_23710);
nand U28970 (N_28970,N_21691,N_21538);
or U28971 (N_28971,N_20015,N_20576);
xnor U28972 (N_28972,N_22469,N_20696);
nand U28973 (N_28973,N_24252,N_24821);
and U28974 (N_28974,N_23254,N_22189);
nand U28975 (N_28975,N_23628,N_20948);
nand U28976 (N_28976,N_24481,N_20163);
and U28977 (N_28977,N_24632,N_23302);
nand U28978 (N_28978,N_22254,N_20285);
nand U28979 (N_28979,N_20076,N_20409);
and U28980 (N_28980,N_24141,N_23552);
xor U28981 (N_28981,N_20433,N_23746);
nor U28982 (N_28982,N_20998,N_20877);
xnor U28983 (N_28983,N_23734,N_22121);
and U28984 (N_28984,N_20681,N_20514);
and U28985 (N_28985,N_21730,N_22153);
nand U28986 (N_28986,N_24503,N_22825);
or U28987 (N_28987,N_21258,N_23629);
nand U28988 (N_28988,N_21290,N_20654);
or U28989 (N_28989,N_24863,N_24628);
and U28990 (N_28990,N_22930,N_23223);
or U28991 (N_28991,N_20038,N_22707);
nor U28992 (N_28992,N_24422,N_23314);
nor U28993 (N_28993,N_22057,N_21288);
or U28994 (N_28994,N_22715,N_23330);
or U28995 (N_28995,N_24989,N_21789);
nand U28996 (N_28996,N_24737,N_22338);
and U28997 (N_28997,N_22278,N_24683);
and U28998 (N_28998,N_20084,N_20687);
or U28999 (N_28999,N_22033,N_24081);
nand U29000 (N_29000,N_24570,N_22037);
nor U29001 (N_29001,N_21324,N_20496);
and U29002 (N_29002,N_23544,N_21078);
nand U29003 (N_29003,N_22637,N_23504);
nor U29004 (N_29004,N_23481,N_21790);
and U29005 (N_29005,N_23800,N_23837);
xnor U29006 (N_29006,N_20148,N_21005);
and U29007 (N_29007,N_21785,N_22154);
and U29008 (N_29008,N_22129,N_21869);
or U29009 (N_29009,N_24417,N_21070);
xnor U29010 (N_29010,N_23326,N_24983);
nand U29011 (N_29011,N_20139,N_22125);
nor U29012 (N_29012,N_20670,N_23756);
nand U29013 (N_29013,N_23421,N_22481);
nor U29014 (N_29014,N_22846,N_20685);
nor U29015 (N_29015,N_21323,N_23144);
xor U29016 (N_29016,N_24961,N_21154);
or U29017 (N_29017,N_23010,N_20604);
and U29018 (N_29018,N_23695,N_24955);
nand U29019 (N_29019,N_21841,N_24353);
or U29020 (N_29020,N_20970,N_21637);
nor U29021 (N_29021,N_24544,N_24680);
or U29022 (N_29022,N_20230,N_21901);
xnor U29023 (N_29023,N_22178,N_24993);
nor U29024 (N_29024,N_21672,N_23531);
nor U29025 (N_29025,N_24931,N_21772);
nand U29026 (N_29026,N_23679,N_23880);
nand U29027 (N_29027,N_24613,N_20927);
and U29028 (N_29028,N_23597,N_20133);
nor U29029 (N_29029,N_21257,N_24594);
and U29030 (N_29030,N_23391,N_21626);
or U29031 (N_29031,N_23660,N_23127);
xor U29032 (N_29032,N_24859,N_22120);
or U29033 (N_29033,N_24969,N_23213);
or U29034 (N_29034,N_23767,N_24358);
or U29035 (N_29035,N_24505,N_24472);
xor U29036 (N_29036,N_23928,N_23689);
xor U29037 (N_29037,N_22164,N_24821);
or U29038 (N_29038,N_22908,N_21404);
xor U29039 (N_29039,N_24251,N_20340);
nand U29040 (N_29040,N_22372,N_23637);
xnor U29041 (N_29041,N_24869,N_24135);
nand U29042 (N_29042,N_20724,N_21687);
and U29043 (N_29043,N_22113,N_22559);
and U29044 (N_29044,N_21228,N_24898);
xor U29045 (N_29045,N_23705,N_24670);
nor U29046 (N_29046,N_23553,N_24641);
nand U29047 (N_29047,N_20100,N_24857);
or U29048 (N_29048,N_24054,N_23148);
and U29049 (N_29049,N_22172,N_20505);
or U29050 (N_29050,N_22371,N_21166);
xor U29051 (N_29051,N_21387,N_23103);
or U29052 (N_29052,N_22093,N_21480);
or U29053 (N_29053,N_20047,N_20594);
nand U29054 (N_29054,N_21997,N_22009);
or U29055 (N_29055,N_20719,N_22486);
xnor U29056 (N_29056,N_24353,N_23627);
nand U29057 (N_29057,N_20075,N_20458);
xnor U29058 (N_29058,N_20655,N_20228);
and U29059 (N_29059,N_23390,N_20201);
xnor U29060 (N_29060,N_22139,N_22165);
xnor U29061 (N_29061,N_22651,N_23710);
nor U29062 (N_29062,N_22990,N_24874);
or U29063 (N_29063,N_24381,N_24316);
and U29064 (N_29064,N_23656,N_20205);
or U29065 (N_29065,N_24212,N_20129);
and U29066 (N_29066,N_22771,N_23687);
nor U29067 (N_29067,N_20539,N_20729);
nand U29068 (N_29068,N_22777,N_24844);
and U29069 (N_29069,N_21327,N_21917);
nand U29070 (N_29070,N_21498,N_21242);
or U29071 (N_29071,N_20394,N_21785);
and U29072 (N_29072,N_20735,N_20581);
nor U29073 (N_29073,N_22748,N_20039);
and U29074 (N_29074,N_23432,N_21999);
nand U29075 (N_29075,N_21429,N_21995);
nand U29076 (N_29076,N_20638,N_22771);
nand U29077 (N_29077,N_21249,N_21032);
xnor U29078 (N_29078,N_21668,N_23037);
or U29079 (N_29079,N_21769,N_23965);
xor U29080 (N_29080,N_21930,N_23101);
xor U29081 (N_29081,N_23321,N_24871);
nand U29082 (N_29082,N_21015,N_21777);
nor U29083 (N_29083,N_21054,N_20674);
xnor U29084 (N_29084,N_21848,N_22011);
nand U29085 (N_29085,N_23545,N_21928);
nand U29086 (N_29086,N_24866,N_20179);
or U29087 (N_29087,N_24411,N_21588);
nand U29088 (N_29088,N_23018,N_22540);
xor U29089 (N_29089,N_20185,N_21142);
nor U29090 (N_29090,N_20111,N_21716);
or U29091 (N_29091,N_20818,N_24103);
nor U29092 (N_29092,N_20854,N_21887);
nor U29093 (N_29093,N_21665,N_24539);
xor U29094 (N_29094,N_24479,N_24550);
or U29095 (N_29095,N_20490,N_23817);
nand U29096 (N_29096,N_22211,N_22702);
and U29097 (N_29097,N_23019,N_23052);
nand U29098 (N_29098,N_21013,N_24509);
nor U29099 (N_29099,N_20337,N_22901);
nor U29100 (N_29100,N_24701,N_20310);
xor U29101 (N_29101,N_23107,N_22860);
xor U29102 (N_29102,N_24911,N_23706);
or U29103 (N_29103,N_20204,N_21898);
nand U29104 (N_29104,N_21007,N_24628);
nand U29105 (N_29105,N_21302,N_20544);
or U29106 (N_29106,N_24662,N_21530);
nor U29107 (N_29107,N_21286,N_20036);
nand U29108 (N_29108,N_24940,N_21220);
and U29109 (N_29109,N_24348,N_21128);
xor U29110 (N_29110,N_23907,N_20944);
nand U29111 (N_29111,N_21978,N_24782);
and U29112 (N_29112,N_21334,N_20073);
and U29113 (N_29113,N_20773,N_22356);
and U29114 (N_29114,N_24426,N_20617);
nor U29115 (N_29115,N_22393,N_24722);
nand U29116 (N_29116,N_24323,N_23724);
and U29117 (N_29117,N_22702,N_23293);
or U29118 (N_29118,N_23509,N_21850);
and U29119 (N_29119,N_23985,N_24787);
nand U29120 (N_29120,N_24462,N_23674);
and U29121 (N_29121,N_20405,N_20187);
and U29122 (N_29122,N_23625,N_21909);
xor U29123 (N_29123,N_23340,N_20177);
xor U29124 (N_29124,N_22554,N_24491);
or U29125 (N_29125,N_23146,N_23047);
nand U29126 (N_29126,N_24827,N_22235);
nor U29127 (N_29127,N_23295,N_20671);
or U29128 (N_29128,N_24300,N_24597);
nor U29129 (N_29129,N_22869,N_22424);
nor U29130 (N_29130,N_24138,N_21233);
nor U29131 (N_29131,N_22408,N_24077);
nand U29132 (N_29132,N_23892,N_20367);
or U29133 (N_29133,N_22529,N_21152);
nor U29134 (N_29134,N_24300,N_24518);
nor U29135 (N_29135,N_20819,N_21018);
nor U29136 (N_29136,N_23859,N_22569);
nor U29137 (N_29137,N_21905,N_23594);
and U29138 (N_29138,N_22170,N_24975);
or U29139 (N_29139,N_22667,N_21555);
xor U29140 (N_29140,N_22079,N_23396);
or U29141 (N_29141,N_20287,N_22578);
xor U29142 (N_29142,N_23788,N_24749);
and U29143 (N_29143,N_20815,N_23907);
and U29144 (N_29144,N_24082,N_22034);
nor U29145 (N_29145,N_21210,N_22458);
xnor U29146 (N_29146,N_20040,N_24503);
xor U29147 (N_29147,N_22463,N_24964);
and U29148 (N_29148,N_22917,N_21728);
xor U29149 (N_29149,N_22356,N_21384);
xor U29150 (N_29150,N_22727,N_24131);
nand U29151 (N_29151,N_20089,N_21639);
or U29152 (N_29152,N_21474,N_23312);
and U29153 (N_29153,N_23916,N_21858);
nand U29154 (N_29154,N_20237,N_24718);
nand U29155 (N_29155,N_20623,N_24251);
nand U29156 (N_29156,N_20889,N_22812);
nand U29157 (N_29157,N_23131,N_23994);
xnor U29158 (N_29158,N_21188,N_21476);
and U29159 (N_29159,N_21303,N_24733);
nor U29160 (N_29160,N_22511,N_23143);
nand U29161 (N_29161,N_22233,N_23585);
nand U29162 (N_29162,N_22314,N_24321);
xor U29163 (N_29163,N_20484,N_24369);
nor U29164 (N_29164,N_24060,N_20608);
and U29165 (N_29165,N_22344,N_23051);
xnor U29166 (N_29166,N_23914,N_20838);
nand U29167 (N_29167,N_24101,N_24390);
nor U29168 (N_29168,N_22877,N_23618);
or U29169 (N_29169,N_20945,N_20418);
and U29170 (N_29170,N_22939,N_20157);
or U29171 (N_29171,N_21129,N_22972);
nand U29172 (N_29172,N_21457,N_24759);
nor U29173 (N_29173,N_23063,N_22134);
xnor U29174 (N_29174,N_20713,N_24366);
nor U29175 (N_29175,N_20348,N_23433);
or U29176 (N_29176,N_23275,N_20515);
or U29177 (N_29177,N_23743,N_21970);
nor U29178 (N_29178,N_24372,N_23581);
nand U29179 (N_29179,N_20578,N_24201);
nor U29180 (N_29180,N_24120,N_23591);
and U29181 (N_29181,N_23341,N_22576);
nor U29182 (N_29182,N_20924,N_22632);
xor U29183 (N_29183,N_20360,N_24188);
nor U29184 (N_29184,N_24511,N_20581);
nor U29185 (N_29185,N_22929,N_23069);
xor U29186 (N_29186,N_24761,N_20930);
nor U29187 (N_29187,N_20556,N_24861);
and U29188 (N_29188,N_21870,N_23138);
nor U29189 (N_29189,N_23338,N_23925);
nand U29190 (N_29190,N_23159,N_24110);
xnor U29191 (N_29191,N_23776,N_22698);
and U29192 (N_29192,N_20922,N_21410);
nand U29193 (N_29193,N_23912,N_20665);
nor U29194 (N_29194,N_22782,N_24859);
xnor U29195 (N_29195,N_23591,N_20622);
nor U29196 (N_29196,N_21584,N_23365);
or U29197 (N_29197,N_20692,N_23005);
xnor U29198 (N_29198,N_24450,N_21644);
xnor U29199 (N_29199,N_24722,N_23577);
and U29200 (N_29200,N_24272,N_24771);
nor U29201 (N_29201,N_23972,N_22670);
nor U29202 (N_29202,N_21905,N_21174);
nand U29203 (N_29203,N_22780,N_22837);
or U29204 (N_29204,N_24290,N_20336);
nand U29205 (N_29205,N_21219,N_21250);
and U29206 (N_29206,N_22605,N_23543);
and U29207 (N_29207,N_22543,N_21583);
or U29208 (N_29208,N_23240,N_21681);
nor U29209 (N_29209,N_23077,N_21697);
or U29210 (N_29210,N_23189,N_21234);
or U29211 (N_29211,N_20335,N_24473);
and U29212 (N_29212,N_21411,N_24270);
nor U29213 (N_29213,N_23930,N_22374);
or U29214 (N_29214,N_20717,N_23033);
xor U29215 (N_29215,N_21920,N_22505);
xnor U29216 (N_29216,N_24609,N_20672);
nand U29217 (N_29217,N_21381,N_21428);
xnor U29218 (N_29218,N_24541,N_22350);
and U29219 (N_29219,N_21454,N_23782);
xor U29220 (N_29220,N_24501,N_23225);
or U29221 (N_29221,N_24191,N_21591);
nor U29222 (N_29222,N_24389,N_20921);
xnor U29223 (N_29223,N_24685,N_22089);
and U29224 (N_29224,N_21807,N_24211);
and U29225 (N_29225,N_23333,N_22958);
or U29226 (N_29226,N_21608,N_20724);
nand U29227 (N_29227,N_22674,N_24402);
and U29228 (N_29228,N_20539,N_22461);
and U29229 (N_29229,N_20284,N_21666);
or U29230 (N_29230,N_23863,N_21102);
or U29231 (N_29231,N_21735,N_21585);
and U29232 (N_29232,N_20706,N_22771);
and U29233 (N_29233,N_23907,N_24971);
nor U29234 (N_29234,N_21997,N_24819);
xor U29235 (N_29235,N_23263,N_22622);
xnor U29236 (N_29236,N_21746,N_20914);
nor U29237 (N_29237,N_20192,N_20150);
nor U29238 (N_29238,N_24516,N_21284);
or U29239 (N_29239,N_23257,N_20096);
or U29240 (N_29240,N_22359,N_23307);
xor U29241 (N_29241,N_23526,N_23593);
and U29242 (N_29242,N_23114,N_21875);
xor U29243 (N_29243,N_21872,N_21585);
and U29244 (N_29244,N_23884,N_23342);
or U29245 (N_29245,N_21081,N_23834);
or U29246 (N_29246,N_23142,N_23813);
nor U29247 (N_29247,N_24384,N_21085);
nor U29248 (N_29248,N_24083,N_23285);
and U29249 (N_29249,N_22604,N_21647);
nand U29250 (N_29250,N_23515,N_23055);
xor U29251 (N_29251,N_21178,N_21203);
xor U29252 (N_29252,N_22445,N_24014);
and U29253 (N_29253,N_20075,N_20023);
nand U29254 (N_29254,N_23478,N_24813);
xnor U29255 (N_29255,N_23320,N_20586);
and U29256 (N_29256,N_22554,N_22854);
or U29257 (N_29257,N_23743,N_24796);
nor U29258 (N_29258,N_21222,N_24246);
and U29259 (N_29259,N_20264,N_20014);
nand U29260 (N_29260,N_24535,N_23845);
xnor U29261 (N_29261,N_24867,N_23853);
nand U29262 (N_29262,N_24194,N_21423);
or U29263 (N_29263,N_23891,N_21017);
nor U29264 (N_29264,N_21012,N_21306);
or U29265 (N_29265,N_21110,N_24122);
nor U29266 (N_29266,N_21064,N_23911);
nor U29267 (N_29267,N_24832,N_22770);
nand U29268 (N_29268,N_21671,N_23653);
nand U29269 (N_29269,N_24251,N_22173);
xor U29270 (N_29270,N_23550,N_22440);
nor U29271 (N_29271,N_24440,N_23456);
nor U29272 (N_29272,N_20218,N_23807);
and U29273 (N_29273,N_20099,N_21721);
or U29274 (N_29274,N_20816,N_21986);
nand U29275 (N_29275,N_22480,N_23692);
nand U29276 (N_29276,N_22881,N_23832);
nand U29277 (N_29277,N_20291,N_22498);
nor U29278 (N_29278,N_22573,N_23110);
nand U29279 (N_29279,N_22102,N_22603);
or U29280 (N_29280,N_24668,N_21237);
or U29281 (N_29281,N_21979,N_21886);
or U29282 (N_29282,N_24372,N_23322);
nand U29283 (N_29283,N_23664,N_24624);
and U29284 (N_29284,N_22960,N_21735);
nor U29285 (N_29285,N_22125,N_22845);
or U29286 (N_29286,N_20854,N_24079);
xnor U29287 (N_29287,N_20659,N_20806);
and U29288 (N_29288,N_23546,N_20487);
nor U29289 (N_29289,N_21557,N_23071);
xor U29290 (N_29290,N_23079,N_21059);
or U29291 (N_29291,N_23635,N_22043);
nand U29292 (N_29292,N_20234,N_24117);
xor U29293 (N_29293,N_20132,N_22169);
nor U29294 (N_29294,N_23652,N_20043);
xnor U29295 (N_29295,N_22558,N_21573);
xor U29296 (N_29296,N_20129,N_24455);
and U29297 (N_29297,N_20588,N_20873);
nand U29298 (N_29298,N_22669,N_22099);
or U29299 (N_29299,N_22792,N_24679);
or U29300 (N_29300,N_23297,N_24985);
nor U29301 (N_29301,N_23569,N_23204);
and U29302 (N_29302,N_22992,N_21268);
or U29303 (N_29303,N_23422,N_24408);
and U29304 (N_29304,N_24626,N_23523);
xnor U29305 (N_29305,N_21721,N_20182);
and U29306 (N_29306,N_22729,N_22255);
nor U29307 (N_29307,N_24368,N_21078);
xor U29308 (N_29308,N_21282,N_22332);
and U29309 (N_29309,N_22725,N_21819);
and U29310 (N_29310,N_23734,N_23252);
and U29311 (N_29311,N_22568,N_24190);
nor U29312 (N_29312,N_24874,N_23791);
and U29313 (N_29313,N_22278,N_22399);
or U29314 (N_29314,N_24319,N_23204);
and U29315 (N_29315,N_21398,N_21620);
nand U29316 (N_29316,N_20721,N_22144);
nor U29317 (N_29317,N_22861,N_23603);
nor U29318 (N_29318,N_20590,N_22410);
nor U29319 (N_29319,N_22929,N_21374);
and U29320 (N_29320,N_22922,N_23579);
nand U29321 (N_29321,N_20071,N_20753);
and U29322 (N_29322,N_24140,N_21589);
or U29323 (N_29323,N_20152,N_23662);
and U29324 (N_29324,N_20101,N_21535);
nand U29325 (N_29325,N_20574,N_21098);
nor U29326 (N_29326,N_24788,N_22977);
and U29327 (N_29327,N_20217,N_21599);
nor U29328 (N_29328,N_24724,N_22840);
or U29329 (N_29329,N_20332,N_24878);
or U29330 (N_29330,N_20972,N_20518);
nand U29331 (N_29331,N_23490,N_23363);
or U29332 (N_29332,N_22276,N_20276);
nor U29333 (N_29333,N_22451,N_20148);
or U29334 (N_29334,N_22108,N_23006);
nand U29335 (N_29335,N_22364,N_24943);
xor U29336 (N_29336,N_22613,N_22423);
and U29337 (N_29337,N_22659,N_22966);
and U29338 (N_29338,N_21347,N_21067);
or U29339 (N_29339,N_24933,N_20698);
xor U29340 (N_29340,N_22921,N_23105);
nor U29341 (N_29341,N_24686,N_24892);
and U29342 (N_29342,N_20409,N_24708);
or U29343 (N_29343,N_21508,N_24713);
xor U29344 (N_29344,N_23951,N_24227);
nor U29345 (N_29345,N_24459,N_21799);
nor U29346 (N_29346,N_21900,N_23816);
nand U29347 (N_29347,N_20895,N_22888);
and U29348 (N_29348,N_24560,N_24608);
and U29349 (N_29349,N_23869,N_20050);
or U29350 (N_29350,N_20495,N_21890);
nor U29351 (N_29351,N_22001,N_21553);
nor U29352 (N_29352,N_24806,N_21049);
or U29353 (N_29353,N_22904,N_24585);
nor U29354 (N_29354,N_24184,N_23022);
xnor U29355 (N_29355,N_24292,N_23476);
and U29356 (N_29356,N_20237,N_21961);
xor U29357 (N_29357,N_24688,N_23618);
and U29358 (N_29358,N_21983,N_24311);
and U29359 (N_29359,N_23686,N_21819);
nand U29360 (N_29360,N_22666,N_21249);
nand U29361 (N_29361,N_21634,N_22076);
and U29362 (N_29362,N_23620,N_21116);
and U29363 (N_29363,N_22070,N_23786);
and U29364 (N_29364,N_21151,N_24315);
nor U29365 (N_29365,N_22091,N_22604);
nor U29366 (N_29366,N_23671,N_24937);
nand U29367 (N_29367,N_22691,N_20291);
xnor U29368 (N_29368,N_22760,N_22195);
or U29369 (N_29369,N_23884,N_23936);
nor U29370 (N_29370,N_22760,N_23442);
nand U29371 (N_29371,N_24541,N_22471);
nor U29372 (N_29372,N_22050,N_22821);
or U29373 (N_29373,N_22222,N_22243);
nand U29374 (N_29374,N_20833,N_22169);
nand U29375 (N_29375,N_21419,N_23844);
nand U29376 (N_29376,N_23539,N_24050);
nand U29377 (N_29377,N_21883,N_22253);
xnor U29378 (N_29378,N_23925,N_24332);
nor U29379 (N_29379,N_23181,N_21838);
xor U29380 (N_29380,N_21232,N_23979);
nand U29381 (N_29381,N_23249,N_24546);
nand U29382 (N_29382,N_21903,N_23149);
or U29383 (N_29383,N_20460,N_21464);
and U29384 (N_29384,N_22452,N_22853);
xnor U29385 (N_29385,N_20697,N_20625);
nand U29386 (N_29386,N_23133,N_21477);
or U29387 (N_29387,N_20555,N_24732);
and U29388 (N_29388,N_24155,N_21893);
and U29389 (N_29389,N_21765,N_24015);
xnor U29390 (N_29390,N_22715,N_24302);
xor U29391 (N_29391,N_24435,N_20520);
xor U29392 (N_29392,N_23067,N_20966);
and U29393 (N_29393,N_20350,N_20696);
or U29394 (N_29394,N_24448,N_21018);
or U29395 (N_29395,N_23649,N_21010);
nor U29396 (N_29396,N_20911,N_21257);
nand U29397 (N_29397,N_23528,N_24943);
and U29398 (N_29398,N_23920,N_21863);
or U29399 (N_29399,N_22388,N_21550);
or U29400 (N_29400,N_23672,N_20070);
nand U29401 (N_29401,N_22495,N_20345);
xor U29402 (N_29402,N_22172,N_24885);
and U29403 (N_29403,N_24869,N_24083);
and U29404 (N_29404,N_24175,N_20139);
nand U29405 (N_29405,N_22403,N_23552);
or U29406 (N_29406,N_22222,N_21212);
nor U29407 (N_29407,N_23292,N_22999);
nor U29408 (N_29408,N_21211,N_24752);
xor U29409 (N_29409,N_24233,N_23928);
xor U29410 (N_29410,N_21798,N_24632);
nor U29411 (N_29411,N_22287,N_21749);
or U29412 (N_29412,N_21032,N_23644);
nor U29413 (N_29413,N_22314,N_21767);
nor U29414 (N_29414,N_22872,N_22994);
xnor U29415 (N_29415,N_22181,N_24184);
nor U29416 (N_29416,N_21343,N_21185);
nand U29417 (N_29417,N_24541,N_20262);
nand U29418 (N_29418,N_24339,N_22862);
and U29419 (N_29419,N_22691,N_23813);
and U29420 (N_29420,N_23259,N_20944);
xnor U29421 (N_29421,N_22159,N_24638);
xnor U29422 (N_29422,N_22117,N_21905);
nand U29423 (N_29423,N_20248,N_24156);
xor U29424 (N_29424,N_21963,N_24863);
nor U29425 (N_29425,N_24316,N_24436);
xor U29426 (N_29426,N_21323,N_22297);
and U29427 (N_29427,N_21962,N_20072);
or U29428 (N_29428,N_22898,N_21647);
nand U29429 (N_29429,N_23414,N_21063);
nor U29430 (N_29430,N_24697,N_24129);
nand U29431 (N_29431,N_20099,N_24696);
or U29432 (N_29432,N_22701,N_22917);
and U29433 (N_29433,N_21916,N_21173);
and U29434 (N_29434,N_23056,N_23136);
or U29435 (N_29435,N_20269,N_22514);
nor U29436 (N_29436,N_23822,N_24342);
and U29437 (N_29437,N_24177,N_20860);
xor U29438 (N_29438,N_21514,N_24406);
nor U29439 (N_29439,N_21599,N_21878);
xnor U29440 (N_29440,N_24691,N_24161);
or U29441 (N_29441,N_24868,N_21213);
and U29442 (N_29442,N_23250,N_24438);
or U29443 (N_29443,N_23089,N_21716);
xnor U29444 (N_29444,N_22817,N_23403);
nor U29445 (N_29445,N_20810,N_23683);
nand U29446 (N_29446,N_24744,N_24310);
xor U29447 (N_29447,N_24377,N_23397);
or U29448 (N_29448,N_22187,N_23950);
nand U29449 (N_29449,N_23732,N_21611);
nor U29450 (N_29450,N_24750,N_20424);
xnor U29451 (N_29451,N_20972,N_24363);
xor U29452 (N_29452,N_24074,N_22305);
nand U29453 (N_29453,N_23472,N_24946);
or U29454 (N_29454,N_20770,N_23954);
nand U29455 (N_29455,N_22522,N_20333);
and U29456 (N_29456,N_23946,N_22533);
and U29457 (N_29457,N_24806,N_24003);
nor U29458 (N_29458,N_24806,N_24752);
nor U29459 (N_29459,N_21950,N_24147);
xor U29460 (N_29460,N_20531,N_21620);
xnor U29461 (N_29461,N_22977,N_24978);
xnor U29462 (N_29462,N_21589,N_24942);
or U29463 (N_29463,N_23202,N_21392);
xnor U29464 (N_29464,N_20544,N_21851);
and U29465 (N_29465,N_22015,N_20500);
xor U29466 (N_29466,N_23737,N_23314);
and U29467 (N_29467,N_20077,N_24234);
nor U29468 (N_29468,N_23556,N_22350);
and U29469 (N_29469,N_22922,N_24579);
xor U29470 (N_29470,N_22675,N_20346);
or U29471 (N_29471,N_24119,N_21240);
xor U29472 (N_29472,N_20319,N_22645);
or U29473 (N_29473,N_21188,N_21326);
and U29474 (N_29474,N_23951,N_21350);
nor U29475 (N_29475,N_21365,N_24178);
nor U29476 (N_29476,N_24848,N_22564);
nor U29477 (N_29477,N_23291,N_23319);
nand U29478 (N_29478,N_21043,N_20501);
nor U29479 (N_29479,N_22932,N_23383);
or U29480 (N_29480,N_22849,N_20092);
nand U29481 (N_29481,N_21276,N_23115);
nand U29482 (N_29482,N_24514,N_21125);
or U29483 (N_29483,N_22318,N_20012);
xnor U29484 (N_29484,N_24627,N_23224);
nand U29485 (N_29485,N_21614,N_23018);
or U29486 (N_29486,N_24767,N_20214);
nand U29487 (N_29487,N_24326,N_20452);
and U29488 (N_29488,N_24791,N_22531);
and U29489 (N_29489,N_24826,N_21197);
nand U29490 (N_29490,N_23584,N_20433);
or U29491 (N_29491,N_21406,N_22460);
and U29492 (N_29492,N_24871,N_24578);
xor U29493 (N_29493,N_22311,N_21706);
or U29494 (N_29494,N_24768,N_24518);
nand U29495 (N_29495,N_24408,N_23760);
and U29496 (N_29496,N_24845,N_22226);
or U29497 (N_29497,N_22968,N_21027);
xnor U29498 (N_29498,N_20514,N_21293);
or U29499 (N_29499,N_22737,N_24320);
xnor U29500 (N_29500,N_24968,N_24615);
xor U29501 (N_29501,N_24472,N_23806);
nor U29502 (N_29502,N_24703,N_22388);
nand U29503 (N_29503,N_23969,N_23032);
and U29504 (N_29504,N_24014,N_24280);
nor U29505 (N_29505,N_24366,N_21200);
and U29506 (N_29506,N_23435,N_23518);
nor U29507 (N_29507,N_20221,N_21365);
or U29508 (N_29508,N_22835,N_23401);
nor U29509 (N_29509,N_21670,N_23550);
or U29510 (N_29510,N_22122,N_23263);
and U29511 (N_29511,N_24835,N_24458);
and U29512 (N_29512,N_22963,N_23338);
xnor U29513 (N_29513,N_22368,N_24475);
or U29514 (N_29514,N_22715,N_24502);
or U29515 (N_29515,N_20545,N_22477);
nor U29516 (N_29516,N_22361,N_21889);
nor U29517 (N_29517,N_24478,N_24630);
xor U29518 (N_29518,N_20434,N_24142);
nor U29519 (N_29519,N_21980,N_23921);
xnor U29520 (N_29520,N_22186,N_22748);
nand U29521 (N_29521,N_22564,N_21860);
or U29522 (N_29522,N_21105,N_21528);
nor U29523 (N_29523,N_20020,N_24148);
nor U29524 (N_29524,N_23560,N_20521);
xnor U29525 (N_29525,N_23251,N_20109);
nand U29526 (N_29526,N_21683,N_21492);
or U29527 (N_29527,N_24389,N_24622);
or U29528 (N_29528,N_23763,N_21095);
or U29529 (N_29529,N_24156,N_22301);
or U29530 (N_29530,N_22816,N_24655);
nor U29531 (N_29531,N_24137,N_23735);
nor U29532 (N_29532,N_22827,N_21075);
and U29533 (N_29533,N_22903,N_23532);
nand U29534 (N_29534,N_21262,N_23573);
nor U29535 (N_29535,N_20557,N_23701);
nand U29536 (N_29536,N_21909,N_24541);
xor U29537 (N_29537,N_21289,N_24281);
nand U29538 (N_29538,N_21395,N_24718);
xnor U29539 (N_29539,N_24508,N_22818);
or U29540 (N_29540,N_20452,N_24292);
nor U29541 (N_29541,N_24398,N_22261);
and U29542 (N_29542,N_23741,N_23222);
nand U29543 (N_29543,N_22289,N_24844);
or U29544 (N_29544,N_22050,N_21721);
and U29545 (N_29545,N_24155,N_23618);
xnor U29546 (N_29546,N_23688,N_23891);
and U29547 (N_29547,N_22970,N_24360);
nand U29548 (N_29548,N_22273,N_22683);
and U29549 (N_29549,N_20826,N_21774);
or U29550 (N_29550,N_24099,N_22251);
nand U29551 (N_29551,N_22300,N_22263);
nand U29552 (N_29552,N_20397,N_20081);
nand U29553 (N_29553,N_23581,N_21630);
or U29554 (N_29554,N_24765,N_21866);
and U29555 (N_29555,N_23685,N_20989);
xnor U29556 (N_29556,N_22537,N_23894);
xor U29557 (N_29557,N_22421,N_24773);
nand U29558 (N_29558,N_24403,N_22436);
xor U29559 (N_29559,N_22919,N_24916);
nor U29560 (N_29560,N_23659,N_22668);
or U29561 (N_29561,N_21324,N_20591);
xnor U29562 (N_29562,N_24462,N_22817);
xnor U29563 (N_29563,N_20784,N_21999);
and U29564 (N_29564,N_20842,N_20885);
nand U29565 (N_29565,N_22027,N_23297);
or U29566 (N_29566,N_24993,N_21414);
nand U29567 (N_29567,N_20806,N_22253);
and U29568 (N_29568,N_20332,N_24603);
nor U29569 (N_29569,N_22019,N_21494);
or U29570 (N_29570,N_23924,N_21672);
nor U29571 (N_29571,N_22627,N_20385);
and U29572 (N_29572,N_20041,N_24492);
nor U29573 (N_29573,N_23086,N_21053);
xor U29574 (N_29574,N_20321,N_23656);
nor U29575 (N_29575,N_23189,N_20168);
or U29576 (N_29576,N_21998,N_24507);
or U29577 (N_29577,N_24347,N_20107);
and U29578 (N_29578,N_24208,N_20347);
and U29579 (N_29579,N_24307,N_20701);
and U29580 (N_29580,N_20295,N_23133);
nand U29581 (N_29581,N_23378,N_21590);
or U29582 (N_29582,N_20048,N_22554);
and U29583 (N_29583,N_23281,N_20015);
xnor U29584 (N_29584,N_24440,N_20267);
nor U29585 (N_29585,N_23586,N_21518);
and U29586 (N_29586,N_23095,N_20697);
and U29587 (N_29587,N_23633,N_24305);
nor U29588 (N_29588,N_23686,N_20797);
nand U29589 (N_29589,N_21122,N_22906);
xor U29590 (N_29590,N_23528,N_21643);
nand U29591 (N_29591,N_20522,N_22579);
or U29592 (N_29592,N_22848,N_23628);
nor U29593 (N_29593,N_22506,N_20778);
xor U29594 (N_29594,N_21771,N_20962);
and U29595 (N_29595,N_21111,N_20790);
nand U29596 (N_29596,N_24821,N_22188);
nand U29597 (N_29597,N_23463,N_20657);
nor U29598 (N_29598,N_23806,N_23997);
xor U29599 (N_29599,N_24383,N_20122);
nand U29600 (N_29600,N_20531,N_22711);
and U29601 (N_29601,N_20568,N_20702);
xor U29602 (N_29602,N_24714,N_20389);
xnor U29603 (N_29603,N_23708,N_24182);
xor U29604 (N_29604,N_22289,N_24548);
nor U29605 (N_29605,N_24963,N_21777);
xor U29606 (N_29606,N_20252,N_22245);
xor U29607 (N_29607,N_22922,N_23801);
and U29608 (N_29608,N_24652,N_24505);
nand U29609 (N_29609,N_23330,N_24178);
xor U29610 (N_29610,N_21747,N_21473);
nand U29611 (N_29611,N_21884,N_24531);
or U29612 (N_29612,N_20480,N_22844);
and U29613 (N_29613,N_21151,N_24199);
or U29614 (N_29614,N_23406,N_22204);
nor U29615 (N_29615,N_20598,N_21013);
or U29616 (N_29616,N_20869,N_20812);
and U29617 (N_29617,N_21313,N_21574);
and U29618 (N_29618,N_21486,N_20429);
nand U29619 (N_29619,N_22526,N_22874);
nand U29620 (N_29620,N_20143,N_22830);
and U29621 (N_29621,N_21597,N_20182);
or U29622 (N_29622,N_23864,N_21648);
or U29623 (N_29623,N_22295,N_20660);
or U29624 (N_29624,N_24445,N_21823);
nor U29625 (N_29625,N_22068,N_21433);
nor U29626 (N_29626,N_22266,N_24149);
or U29627 (N_29627,N_20693,N_22997);
xor U29628 (N_29628,N_22120,N_24360);
nand U29629 (N_29629,N_22127,N_22051);
nand U29630 (N_29630,N_20036,N_24749);
nor U29631 (N_29631,N_23525,N_20293);
or U29632 (N_29632,N_21006,N_20132);
and U29633 (N_29633,N_20812,N_21895);
nor U29634 (N_29634,N_23195,N_24620);
xor U29635 (N_29635,N_24661,N_20666);
xor U29636 (N_29636,N_24428,N_23913);
and U29637 (N_29637,N_23738,N_23679);
or U29638 (N_29638,N_20937,N_20999);
nand U29639 (N_29639,N_24503,N_21372);
nor U29640 (N_29640,N_21231,N_23800);
xor U29641 (N_29641,N_20238,N_20858);
and U29642 (N_29642,N_23991,N_24000);
xor U29643 (N_29643,N_24860,N_23454);
xnor U29644 (N_29644,N_24384,N_23513);
xor U29645 (N_29645,N_20658,N_23228);
nor U29646 (N_29646,N_20495,N_22843);
nor U29647 (N_29647,N_21922,N_24441);
xor U29648 (N_29648,N_21725,N_22808);
and U29649 (N_29649,N_20444,N_23904);
and U29650 (N_29650,N_22130,N_21180);
nand U29651 (N_29651,N_20913,N_22258);
nand U29652 (N_29652,N_20352,N_21045);
nand U29653 (N_29653,N_22821,N_24035);
and U29654 (N_29654,N_22639,N_23911);
and U29655 (N_29655,N_24482,N_22237);
nand U29656 (N_29656,N_22500,N_22702);
nor U29657 (N_29657,N_24373,N_23480);
xor U29658 (N_29658,N_24714,N_23303);
nand U29659 (N_29659,N_20136,N_20513);
nor U29660 (N_29660,N_24159,N_21023);
nand U29661 (N_29661,N_22055,N_23506);
nor U29662 (N_29662,N_22067,N_21409);
nor U29663 (N_29663,N_22131,N_21453);
nand U29664 (N_29664,N_22380,N_21135);
and U29665 (N_29665,N_22314,N_20394);
or U29666 (N_29666,N_22986,N_24806);
and U29667 (N_29667,N_23860,N_20519);
nand U29668 (N_29668,N_22982,N_21593);
xnor U29669 (N_29669,N_21358,N_23013);
nor U29670 (N_29670,N_20287,N_23549);
nor U29671 (N_29671,N_20716,N_23504);
xor U29672 (N_29672,N_20572,N_24544);
nand U29673 (N_29673,N_22005,N_20863);
nand U29674 (N_29674,N_23335,N_23522);
xor U29675 (N_29675,N_23527,N_24305);
xor U29676 (N_29676,N_21966,N_22004);
and U29677 (N_29677,N_24105,N_20379);
and U29678 (N_29678,N_24805,N_20751);
nor U29679 (N_29679,N_21331,N_21734);
xor U29680 (N_29680,N_20246,N_20794);
or U29681 (N_29681,N_24281,N_23127);
or U29682 (N_29682,N_20797,N_22016);
nor U29683 (N_29683,N_23891,N_23274);
nor U29684 (N_29684,N_22683,N_23623);
nand U29685 (N_29685,N_24282,N_21778);
xnor U29686 (N_29686,N_24942,N_23636);
nand U29687 (N_29687,N_22052,N_22790);
nor U29688 (N_29688,N_23346,N_23745);
and U29689 (N_29689,N_20694,N_24986);
nand U29690 (N_29690,N_23244,N_24696);
nor U29691 (N_29691,N_21249,N_24266);
nand U29692 (N_29692,N_24087,N_21715);
nor U29693 (N_29693,N_23863,N_23810);
xnor U29694 (N_29694,N_21572,N_22213);
xor U29695 (N_29695,N_22581,N_20005);
and U29696 (N_29696,N_23523,N_23668);
or U29697 (N_29697,N_22366,N_21318);
nor U29698 (N_29698,N_20982,N_21583);
and U29699 (N_29699,N_22863,N_24908);
or U29700 (N_29700,N_21559,N_20641);
and U29701 (N_29701,N_22817,N_24645);
xor U29702 (N_29702,N_21355,N_22626);
xor U29703 (N_29703,N_24995,N_24970);
xnor U29704 (N_29704,N_23631,N_20451);
nand U29705 (N_29705,N_21177,N_21223);
or U29706 (N_29706,N_22689,N_21796);
nor U29707 (N_29707,N_22295,N_21945);
xnor U29708 (N_29708,N_22980,N_22203);
or U29709 (N_29709,N_23330,N_21464);
or U29710 (N_29710,N_23973,N_20340);
xor U29711 (N_29711,N_21839,N_23651);
nor U29712 (N_29712,N_20884,N_24560);
nor U29713 (N_29713,N_22126,N_22984);
nor U29714 (N_29714,N_20311,N_23554);
nor U29715 (N_29715,N_21261,N_23471);
xor U29716 (N_29716,N_22688,N_22305);
or U29717 (N_29717,N_22196,N_24540);
nor U29718 (N_29718,N_24919,N_21924);
or U29719 (N_29719,N_24298,N_23188);
xor U29720 (N_29720,N_21976,N_23951);
nand U29721 (N_29721,N_20915,N_22593);
xor U29722 (N_29722,N_21714,N_21684);
xnor U29723 (N_29723,N_23533,N_24045);
and U29724 (N_29724,N_22667,N_24346);
nor U29725 (N_29725,N_23662,N_22649);
xnor U29726 (N_29726,N_22305,N_22967);
and U29727 (N_29727,N_20735,N_21775);
and U29728 (N_29728,N_20204,N_24898);
nor U29729 (N_29729,N_20795,N_24560);
nand U29730 (N_29730,N_20785,N_21190);
xor U29731 (N_29731,N_23780,N_24631);
xnor U29732 (N_29732,N_24450,N_20473);
nor U29733 (N_29733,N_21279,N_24039);
or U29734 (N_29734,N_21332,N_23135);
nor U29735 (N_29735,N_23656,N_20166);
and U29736 (N_29736,N_24836,N_24795);
nor U29737 (N_29737,N_23260,N_24651);
nor U29738 (N_29738,N_22657,N_23855);
xor U29739 (N_29739,N_23117,N_21993);
and U29740 (N_29740,N_24776,N_24617);
nor U29741 (N_29741,N_24233,N_20795);
nand U29742 (N_29742,N_23635,N_21550);
xnor U29743 (N_29743,N_22310,N_22455);
or U29744 (N_29744,N_22611,N_22968);
nand U29745 (N_29745,N_22179,N_23535);
nor U29746 (N_29746,N_22346,N_24569);
or U29747 (N_29747,N_22106,N_23597);
or U29748 (N_29748,N_20597,N_22906);
nor U29749 (N_29749,N_24108,N_22717);
nor U29750 (N_29750,N_22413,N_22371);
xnor U29751 (N_29751,N_24136,N_22354);
nand U29752 (N_29752,N_20926,N_22032);
nor U29753 (N_29753,N_21486,N_21609);
xnor U29754 (N_29754,N_23986,N_20882);
or U29755 (N_29755,N_20792,N_24150);
and U29756 (N_29756,N_21194,N_20550);
or U29757 (N_29757,N_24401,N_24625);
nand U29758 (N_29758,N_20693,N_23548);
nand U29759 (N_29759,N_21365,N_21199);
and U29760 (N_29760,N_24491,N_21816);
nor U29761 (N_29761,N_21534,N_23239);
and U29762 (N_29762,N_22230,N_23312);
nand U29763 (N_29763,N_23811,N_24498);
and U29764 (N_29764,N_24161,N_24972);
or U29765 (N_29765,N_22903,N_22420);
xnor U29766 (N_29766,N_21683,N_22495);
nand U29767 (N_29767,N_24177,N_22915);
and U29768 (N_29768,N_22051,N_21246);
and U29769 (N_29769,N_23056,N_20446);
or U29770 (N_29770,N_24499,N_22375);
nand U29771 (N_29771,N_23369,N_24046);
xor U29772 (N_29772,N_21147,N_22346);
nor U29773 (N_29773,N_23750,N_23788);
or U29774 (N_29774,N_20995,N_23665);
and U29775 (N_29775,N_23261,N_23085);
nor U29776 (N_29776,N_23813,N_20520);
nand U29777 (N_29777,N_20898,N_20919);
nand U29778 (N_29778,N_22453,N_24462);
or U29779 (N_29779,N_22518,N_23100);
nand U29780 (N_29780,N_21619,N_21537);
nor U29781 (N_29781,N_20107,N_23834);
nand U29782 (N_29782,N_24481,N_20254);
xnor U29783 (N_29783,N_22687,N_20822);
nand U29784 (N_29784,N_24474,N_23771);
nor U29785 (N_29785,N_20809,N_24289);
xor U29786 (N_29786,N_21749,N_24961);
or U29787 (N_29787,N_24325,N_22564);
nand U29788 (N_29788,N_24522,N_23915);
and U29789 (N_29789,N_24745,N_23430);
nand U29790 (N_29790,N_23016,N_23308);
or U29791 (N_29791,N_20462,N_23018);
nand U29792 (N_29792,N_21925,N_22802);
nor U29793 (N_29793,N_20615,N_21758);
xnor U29794 (N_29794,N_21587,N_24638);
nand U29795 (N_29795,N_20895,N_21860);
nor U29796 (N_29796,N_24662,N_22346);
or U29797 (N_29797,N_22827,N_24361);
and U29798 (N_29798,N_23934,N_23335);
xor U29799 (N_29799,N_23756,N_22197);
nor U29800 (N_29800,N_22845,N_20775);
nand U29801 (N_29801,N_24985,N_23748);
nand U29802 (N_29802,N_20884,N_20999);
nor U29803 (N_29803,N_20396,N_21611);
or U29804 (N_29804,N_21313,N_20023);
nor U29805 (N_29805,N_22704,N_20627);
nand U29806 (N_29806,N_23468,N_22583);
or U29807 (N_29807,N_21182,N_20988);
or U29808 (N_29808,N_23655,N_21832);
xnor U29809 (N_29809,N_21605,N_20412);
xor U29810 (N_29810,N_21009,N_20557);
xor U29811 (N_29811,N_23417,N_20971);
and U29812 (N_29812,N_23783,N_20655);
xnor U29813 (N_29813,N_20762,N_23563);
nand U29814 (N_29814,N_22232,N_21574);
nand U29815 (N_29815,N_21820,N_21016);
and U29816 (N_29816,N_22134,N_22253);
and U29817 (N_29817,N_20813,N_22608);
nand U29818 (N_29818,N_24728,N_24243);
nand U29819 (N_29819,N_21052,N_22119);
nand U29820 (N_29820,N_24522,N_24182);
and U29821 (N_29821,N_20964,N_24422);
or U29822 (N_29822,N_20820,N_24642);
or U29823 (N_29823,N_22019,N_23144);
or U29824 (N_29824,N_23220,N_21203);
nor U29825 (N_29825,N_22504,N_23662);
nand U29826 (N_29826,N_20907,N_23300);
and U29827 (N_29827,N_20288,N_23284);
and U29828 (N_29828,N_20446,N_22358);
nor U29829 (N_29829,N_21647,N_24249);
nand U29830 (N_29830,N_22686,N_21673);
xor U29831 (N_29831,N_23782,N_21865);
xnor U29832 (N_29832,N_20809,N_24382);
xnor U29833 (N_29833,N_20173,N_24406);
or U29834 (N_29834,N_21765,N_24485);
or U29835 (N_29835,N_24225,N_21632);
or U29836 (N_29836,N_20814,N_21630);
and U29837 (N_29837,N_21169,N_20827);
nor U29838 (N_29838,N_21979,N_24872);
and U29839 (N_29839,N_24302,N_23279);
or U29840 (N_29840,N_21911,N_24291);
or U29841 (N_29841,N_21752,N_24288);
and U29842 (N_29842,N_22151,N_22654);
nor U29843 (N_29843,N_22191,N_23540);
and U29844 (N_29844,N_23996,N_23707);
nor U29845 (N_29845,N_22711,N_23825);
xnor U29846 (N_29846,N_20036,N_23990);
nand U29847 (N_29847,N_24883,N_24242);
or U29848 (N_29848,N_24152,N_24271);
or U29849 (N_29849,N_20385,N_23476);
or U29850 (N_29850,N_22823,N_20208);
nand U29851 (N_29851,N_24725,N_23064);
or U29852 (N_29852,N_23065,N_24634);
and U29853 (N_29853,N_20704,N_22527);
nand U29854 (N_29854,N_20822,N_22179);
and U29855 (N_29855,N_24757,N_24609);
and U29856 (N_29856,N_20768,N_24935);
nand U29857 (N_29857,N_21797,N_20510);
nand U29858 (N_29858,N_21093,N_24002);
and U29859 (N_29859,N_21616,N_21195);
or U29860 (N_29860,N_22283,N_21775);
or U29861 (N_29861,N_23320,N_22654);
xor U29862 (N_29862,N_20197,N_22440);
xnor U29863 (N_29863,N_20971,N_20530);
xor U29864 (N_29864,N_21037,N_21254);
and U29865 (N_29865,N_24973,N_23636);
xnor U29866 (N_29866,N_22820,N_23672);
or U29867 (N_29867,N_20343,N_24443);
and U29868 (N_29868,N_23567,N_22361);
nor U29869 (N_29869,N_21511,N_22554);
xor U29870 (N_29870,N_20444,N_21857);
or U29871 (N_29871,N_20203,N_24035);
or U29872 (N_29872,N_23596,N_22402);
and U29873 (N_29873,N_20416,N_23614);
nand U29874 (N_29874,N_21681,N_23331);
nand U29875 (N_29875,N_21082,N_20589);
xnor U29876 (N_29876,N_20508,N_21558);
or U29877 (N_29877,N_22139,N_22390);
or U29878 (N_29878,N_23334,N_23205);
and U29879 (N_29879,N_24368,N_22017);
or U29880 (N_29880,N_23317,N_21771);
and U29881 (N_29881,N_22445,N_21569);
xor U29882 (N_29882,N_20098,N_22972);
or U29883 (N_29883,N_22175,N_24651);
nand U29884 (N_29884,N_24736,N_21691);
or U29885 (N_29885,N_21188,N_22963);
or U29886 (N_29886,N_23295,N_23074);
nand U29887 (N_29887,N_21652,N_21895);
xor U29888 (N_29888,N_24909,N_22581);
nor U29889 (N_29889,N_20819,N_22516);
and U29890 (N_29890,N_23508,N_23881);
or U29891 (N_29891,N_21935,N_22168);
nand U29892 (N_29892,N_24918,N_24742);
or U29893 (N_29893,N_21031,N_22787);
and U29894 (N_29894,N_23189,N_22716);
nand U29895 (N_29895,N_23116,N_23533);
nand U29896 (N_29896,N_21433,N_24174);
or U29897 (N_29897,N_24374,N_20554);
and U29898 (N_29898,N_23317,N_23954);
nand U29899 (N_29899,N_23221,N_22515);
nand U29900 (N_29900,N_22140,N_21129);
nor U29901 (N_29901,N_22559,N_23988);
and U29902 (N_29902,N_23792,N_20082);
and U29903 (N_29903,N_20949,N_24547);
xnor U29904 (N_29904,N_23546,N_20542);
xor U29905 (N_29905,N_21466,N_24282);
nor U29906 (N_29906,N_23967,N_23164);
or U29907 (N_29907,N_23875,N_20397);
nand U29908 (N_29908,N_20158,N_21332);
or U29909 (N_29909,N_24594,N_24010);
nand U29910 (N_29910,N_23708,N_23381);
and U29911 (N_29911,N_21275,N_24432);
nor U29912 (N_29912,N_23711,N_22281);
or U29913 (N_29913,N_22540,N_24577);
nand U29914 (N_29914,N_23568,N_23981);
nand U29915 (N_29915,N_22112,N_21001);
xnor U29916 (N_29916,N_23459,N_20906);
and U29917 (N_29917,N_21627,N_22746);
nand U29918 (N_29918,N_24958,N_22285);
or U29919 (N_29919,N_23379,N_23792);
nand U29920 (N_29920,N_20004,N_23300);
nand U29921 (N_29921,N_24861,N_21906);
nor U29922 (N_29922,N_23901,N_21825);
or U29923 (N_29923,N_24231,N_22411);
and U29924 (N_29924,N_21920,N_24235);
xor U29925 (N_29925,N_20564,N_22341);
nand U29926 (N_29926,N_20509,N_24244);
nor U29927 (N_29927,N_21759,N_23928);
nor U29928 (N_29928,N_23871,N_20627);
xnor U29929 (N_29929,N_20635,N_22722);
xnor U29930 (N_29930,N_20070,N_22910);
and U29931 (N_29931,N_23382,N_23517);
nor U29932 (N_29932,N_20215,N_23018);
nor U29933 (N_29933,N_22465,N_22243);
nor U29934 (N_29934,N_24205,N_21346);
and U29935 (N_29935,N_23570,N_24923);
or U29936 (N_29936,N_20187,N_23080);
or U29937 (N_29937,N_20692,N_21728);
and U29938 (N_29938,N_21334,N_21859);
or U29939 (N_29939,N_20186,N_22774);
nand U29940 (N_29940,N_24933,N_22934);
nor U29941 (N_29941,N_20927,N_21008);
or U29942 (N_29942,N_22114,N_22232);
and U29943 (N_29943,N_22463,N_24644);
and U29944 (N_29944,N_24729,N_22653);
xor U29945 (N_29945,N_23991,N_24710);
or U29946 (N_29946,N_22222,N_21039);
or U29947 (N_29947,N_22644,N_22367);
nor U29948 (N_29948,N_24746,N_20232);
xnor U29949 (N_29949,N_21677,N_23626);
xnor U29950 (N_29950,N_22052,N_22337);
and U29951 (N_29951,N_20228,N_20112);
and U29952 (N_29952,N_21001,N_20626);
and U29953 (N_29953,N_22858,N_21947);
nand U29954 (N_29954,N_22932,N_24577);
nor U29955 (N_29955,N_20806,N_23686);
and U29956 (N_29956,N_22514,N_20005);
xor U29957 (N_29957,N_24005,N_22030);
nor U29958 (N_29958,N_23747,N_24691);
xor U29959 (N_29959,N_20713,N_23519);
or U29960 (N_29960,N_23310,N_20072);
or U29961 (N_29961,N_22910,N_24333);
and U29962 (N_29962,N_21029,N_20137);
and U29963 (N_29963,N_23447,N_22936);
nor U29964 (N_29964,N_24853,N_22653);
or U29965 (N_29965,N_20134,N_23310);
nor U29966 (N_29966,N_20030,N_22955);
nor U29967 (N_29967,N_22823,N_21069);
or U29968 (N_29968,N_24158,N_22778);
and U29969 (N_29969,N_24140,N_20839);
and U29970 (N_29970,N_20643,N_21121);
and U29971 (N_29971,N_21113,N_22412);
and U29972 (N_29972,N_20900,N_23468);
and U29973 (N_29973,N_23994,N_24314);
nand U29974 (N_29974,N_24300,N_22609);
nand U29975 (N_29975,N_24440,N_21114);
nand U29976 (N_29976,N_23716,N_20368);
or U29977 (N_29977,N_20498,N_23858);
or U29978 (N_29978,N_21684,N_22053);
and U29979 (N_29979,N_21413,N_23513);
xnor U29980 (N_29980,N_20208,N_22530);
and U29981 (N_29981,N_24812,N_20127);
nand U29982 (N_29982,N_24271,N_21109);
nand U29983 (N_29983,N_21030,N_24399);
or U29984 (N_29984,N_24065,N_20664);
or U29985 (N_29985,N_21993,N_20881);
nand U29986 (N_29986,N_20554,N_22067);
and U29987 (N_29987,N_21612,N_21324);
nor U29988 (N_29988,N_22947,N_20093);
nand U29989 (N_29989,N_24409,N_20270);
nor U29990 (N_29990,N_20721,N_20491);
nand U29991 (N_29991,N_23319,N_22815);
nand U29992 (N_29992,N_23737,N_21866);
xor U29993 (N_29993,N_20516,N_24241);
nor U29994 (N_29994,N_24157,N_24380);
xnor U29995 (N_29995,N_23877,N_21869);
nor U29996 (N_29996,N_23096,N_23035);
nor U29997 (N_29997,N_20237,N_23228);
xnor U29998 (N_29998,N_20445,N_21686);
or U29999 (N_29999,N_23485,N_22412);
nor U30000 (N_30000,N_27294,N_25836);
nand U30001 (N_30001,N_27101,N_27347);
nor U30002 (N_30002,N_26465,N_29165);
nand U30003 (N_30003,N_27563,N_27244);
nand U30004 (N_30004,N_29097,N_28568);
xor U30005 (N_30005,N_26979,N_27695);
nor U30006 (N_30006,N_25779,N_27595);
nor U30007 (N_30007,N_28999,N_26964);
xnor U30008 (N_30008,N_27431,N_28416);
xor U30009 (N_30009,N_28351,N_27112);
xor U30010 (N_30010,N_29291,N_25337);
and U30011 (N_30011,N_29605,N_27046);
or U30012 (N_30012,N_29975,N_25938);
and U30013 (N_30013,N_29904,N_25731);
and U30014 (N_30014,N_28097,N_26537);
xor U30015 (N_30015,N_26802,N_25065);
nor U30016 (N_30016,N_29689,N_28409);
or U30017 (N_30017,N_28666,N_27470);
nand U30018 (N_30018,N_26395,N_27894);
nor U30019 (N_30019,N_27374,N_28074);
nor U30020 (N_30020,N_28357,N_28191);
or U30021 (N_30021,N_26147,N_25297);
nand U30022 (N_30022,N_25044,N_28225);
and U30023 (N_30023,N_27079,N_27623);
nor U30024 (N_30024,N_28777,N_26246);
and U30025 (N_30025,N_25062,N_26106);
or U30026 (N_30026,N_27909,N_28491);
and U30027 (N_30027,N_29162,N_25041);
xnor U30028 (N_30028,N_27056,N_27759);
or U30029 (N_30029,N_25224,N_28532);
nand U30030 (N_30030,N_25945,N_28885);
or U30031 (N_30031,N_27234,N_26664);
and U30032 (N_30032,N_25621,N_26776);
nand U30033 (N_30033,N_26487,N_28986);
and U30034 (N_30034,N_27031,N_28790);
and U30035 (N_30035,N_29151,N_27673);
nor U30036 (N_30036,N_28541,N_25641);
nand U30037 (N_30037,N_25728,N_25823);
and U30038 (N_30038,N_27153,N_28239);
and U30039 (N_30039,N_26004,N_26604);
nor U30040 (N_30040,N_27076,N_25634);
nor U30041 (N_30041,N_28298,N_26293);
or U30042 (N_30042,N_28236,N_29918);
and U30043 (N_30043,N_25375,N_26583);
and U30044 (N_30044,N_25834,N_29915);
nand U30045 (N_30045,N_26197,N_26286);
nand U30046 (N_30046,N_28242,N_25689);
nand U30047 (N_30047,N_26672,N_28055);
or U30048 (N_30048,N_27457,N_29170);
nor U30049 (N_30049,N_29411,N_28158);
or U30050 (N_30050,N_29383,N_28406);
xor U30051 (N_30051,N_25164,N_28907);
xor U30052 (N_30052,N_29060,N_25220);
nand U30053 (N_30053,N_26712,N_29512);
or U30054 (N_30054,N_27286,N_25829);
or U30055 (N_30055,N_25930,N_28766);
nor U30056 (N_30056,N_27312,N_28270);
nand U30057 (N_30057,N_27151,N_25747);
and U30058 (N_30058,N_29667,N_25825);
xor U30059 (N_30059,N_26685,N_28412);
nor U30060 (N_30060,N_29869,N_28053);
nand U30061 (N_30061,N_26791,N_28827);
nand U30062 (N_30062,N_26140,N_29739);
and U30063 (N_30063,N_27653,N_28060);
nand U30064 (N_30064,N_28340,N_26084);
nor U30065 (N_30065,N_25911,N_25984);
nor U30066 (N_30066,N_27384,N_27096);
and U30067 (N_30067,N_27117,N_27308);
or U30068 (N_30068,N_27259,N_26401);
nor U30069 (N_30069,N_25437,N_28617);
nand U30070 (N_30070,N_28595,N_29310);
nand U30071 (N_30071,N_29846,N_29417);
nand U30072 (N_30072,N_25376,N_28130);
nand U30073 (N_30073,N_28573,N_28194);
and U30074 (N_30074,N_25878,N_28728);
nor U30075 (N_30075,N_28632,N_28170);
xnor U30076 (N_30076,N_27812,N_25471);
nor U30077 (N_30077,N_26539,N_29692);
nor U30078 (N_30078,N_29231,N_25649);
xnor U30079 (N_30079,N_27821,N_29397);
and U30080 (N_30080,N_29150,N_28626);
and U30081 (N_30081,N_25762,N_27020);
xnor U30082 (N_30082,N_27702,N_27647);
nor U30083 (N_30083,N_28774,N_27390);
or U30084 (N_30084,N_25710,N_25599);
nand U30085 (N_30085,N_26740,N_26486);
nor U30086 (N_30086,N_25772,N_26003);
nand U30087 (N_30087,N_28330,N_27837);
or U30088 (N_30088,N_27254,N_27028);
xnor U30089 (N_30089,N_25839,N_25311);
nand U30090 (N_30090,N_28830,N_25391);
or U30091 (N_30091,N_25617,N_29715);
xor U30092 (N_30092,N_26963,N_25629);
nor U30093 (N_30093,N_28017,N_29558);
and U30094 (N_30094,N_28024,N_26173);
nor U30095 (N_30095,N_27646,N_29299);
and U30096 (N_30096,N_26865,N_29652);
and U30097 (N_30097,N_27340,N_27484);
or U30098 (N_30098,N_26602,N_28596);
nor U30099 (N_30099,N_27953,N_25505);
nand U30100 (N_30100,N_27375,N_25462);
and U30101 (N_30101,N_29245,N_26386);
and U30102 (N_30102,N_27570,N_28462);
or U30103 (N_30103,N_25524,N_28968);
or U30104 (N_30104,N_29560,N_29862);
xnor U30105 (N_30105,N_25927,N_25327);
and U30106 (N_30106,N_25926,N_29949);
xor U30107 (N_30107,N_28585,N_29422);
and U30108 (N_30108,N_27852,N_26440);
nor U30109 (N_30109,N_25329,N_26161);
xor U30110 (N_30110,N_27224,N_26909);
and U30111 (N_30111,N_26176,N_26561);
xor U30112 (N_30112,N_28163,N_28865);
nor U30113 (N_30113,N_25607,N_28392);
nand U30114 (N_30114,N_28828,N_25029);
and U30115 (N_30115,N_27229,N_28927);
or U30116 (N_30116,N_27978,N_27104);
and U30117 (N_30117,N_28721,N_28787);
nor U30118 (N_30118,N_29252,N_29164);
xor U30119 (N_30119,N_29214,N_25500);
and U30120 (N_30120,N_27635,N_27630);
xor U30121 (N_30121,N_27580,N_26704);
nor U30122 (N_30122,N_28281,N_25426);
xor U30123 (N_30123,N_25459,N_29349);
and U30124 (N_30124,N_25625,N_25765);
xor U30125 (N_30125,N_28430,N_26476);
xor U30126 (N_30126,N_28183,N_26238);
and U30127 (N_30127,N_28161,N_28711);
or U30128 (N_30128,N_29788,N_26675);
or U30129 (N_30129,N_28495,N_29483);
and U30130 (N_30130,N_26033,N_25814);
or U30131 (N_30131,N_27967,N_26457);
xnor U30132 (N_30132,N_27977,N_25730);
xnor U30133 (N_30133,N_29221,N_27246);
nor U30134 (N_30134,N_28493,N_28373);
nor U30135 (N_30135,N_28886,N_26977);
nor U30136 (N_30136,N_28943,N_28072);
or U30137 (N_30137,N_27189,N_26702);
nand U30138 (N_30138,N_29193,N_29507);
nand U30139 (N_30139,N_26387,N_29554);
or U30140 (N_30140,N_29648,N_29191);
xnor U30141 (N_30141,N_28197,N_25425);
or U30142 (N_30142,N_27777,N_29100);
or U30143 (N_30143,N_27007,N_28915);
nand U30144 (N_30144,N_27337,N_28575);
nand U30145 (N_30145,N_26914,N_27245);
xor U30146 (N_30146,N_29384,N_25248);
or U30147 (N_30147,N_29580,N_25871);
and U30148 (N_30148,N_28807,N_27059);
or U30149 (N_30149,N_25559,N_26768);
nand U30150 (N_30150,N_27736,N_28897);
nor U30151 (N_30151,N_27517,N_26677);
nand U30152 (N_30152,N_27649,N_25897);
and U30153 (N_30153,N_28080,N_28862);
xor U30154 (N_30154,N_29892,N_25113);
and U30155 (N_30155,N_28082,N_27211);
and U30156 (N_30156,N_27146,N_26405);
and U30157 (N_30157,N_25974,N_28376);
xnor U30158 (N_30158,N_25511,N_29099);
or U30159 (N_30159,N_28377,N_27656);
nand U30160 (N_30160,N_29693,N_26576);
nand U30161 (N_30161,N_29913,N_29888);
and U30162 (N_30162,N_25236,N_26563);
nor U30163 (N_30163,N_28372,N_26326);
nand U30164 (N_30164,N_25786,N_26968);
nor U30165 (N_30165,N_29045,N_26463);
xnor U30166 (N_30166,N_28278,N_28136);
xnor U30167 (N_30167,N_29561,N_25484);
and U30168 (N_30168,N_27052,N_26923);
xnor U30169 (N_30169,N_28166,N_25308);
or U30170 (N_30170,N_25388,N_26729);
nor U30171 (N_30171,N_26959,N_27776);
nand U30172 (N_30172,N_29873,N_25396);
nand U30173 (N_30173,N_26365,N_25647);
nand U30174 (N_30174,N_29073,N_26966);
nor U30175 (N_30175,N_28797,N_29457);
xnor U30176 (N_30176,N_25445,N_29189);
and U30177 (N_30177,N_29009,N_29064);
xnor U30178 (N_30178,N_27851,N_27219);
xnor U30179 (N_30179,N_28820,N_26524);
nor U30180 (N_30180,N_27073,N_28224);
nor U30181 (N_30181,N_28567,N_29705);
nand U30182 (N_30182,N_28219,N_25434);
and U30183 (N_30183,N_28508,N_25048);
and U30184 (N_30184,N_29968,N_27983);
nor U30185 (N_30185,N_27678,N_27538);
xor U30186 (N_30186,N_26577,N_26489);
and U30187 (N_30187,N_25700,N_29242);
nor U30188 (N_30188,N_25476,N_28552);
nand U30189 (N_30189,N_29940,N_27813);
or U30190 (N_30190,N_28691,N_28366);
xnor U30191 (N_30191,N_27213,N_26895);
or U30192 (N_30192,N_26887,N_28920);
nor U30193 (N_30193,N_27601,N_29714);
nand U30194 (N_30194,N_25015,N_25146);
xnor U30195 (N_30195,N_28087,N_28824);
nor U30196 (N_30196,N_27618,N_25870);
and U30197 (N_30197,N_28299,N_26253);
nand U30198 (N_30198,N_25133,N_29954);
or U30199 (N_30199,N_29502,N_26133);
and U30200 (N_30200,N_27148,N_25225);
xor U30201 (N_30201,N_25043,N_26634);
xor U30202 (N_30202,N_26321,N_26030);
or U30203 (N_30203,N_26610,N_27632);
and U30204 (N_30204,N_27694,N_28928);
nor U30205 (N_30205,N_27458,N_25850);
and U30206 (N_30206,N_25414,N_27969);
nand U30207 (N_30207,N_29233,N_29264);
nor U30208 (N_30208,N_25746,N_28058);
and U30209 (N_30209,N_26715,N_29763);
xnor U30210 (N_30210,N_27121,N_29497);
xor U30211 (N_30211,N_29066,N_29447);
nor U30212 (N_30212,N_26567,N_28459);
xnor U30213 (N_30213,N_29790,N_26283);
and U30214 (N_30214,N_25017,N_26810);
nand U30215 (N_30215,N_28124,N_25053);
nand U30216 (N_30216,N_25319,N_26936);
and U30217 (N_30217,N_26181,N_27665);
and U30218 (N_30218,N_27469,N_29444);
or U30219 (N_30219,N_29455,N_26965);
xor U30220 (N_30220,N_27515,N_29037);
and U30221 (N_30221,N_26543,N_25679);
xor U30222 (N_30222,N_27970,N_27712);
xor U30223 (N_30223,N_27826,N_29498);
nand U30224 (N_30224,N_25359,N_25651);
or U30225 (N_30225,N_26038,N_27267);
or U30226 (N_30226,N_27130,N_29570);
xnor U30227 (N_30227,N_26245,N_29036);
nand U30228 (N_30228,N_26573,N_28654);
and U30229 (N_30229,N_27296,N_27547);
xnor U30230 (N_30230,N_29459,N_25522);
and U30231 (N_30231,N_27562,N_28308);
or U30232 (N_30232,N_29318,N_29596);
or U30233 (N_30233,N_29813,N_29988);
nand U30234 (N_30234,N_28908,N_28794);
and U30235 (N_30235,N_27086,N_28761);
nor U30236 (N_30236,N_26931,N_29838);
nand U30237 (N_30237,N_28380,N_25761);
nor U30238 (N_30238,N_28816,N_27237);
or U30239 (N_30239,N_25623,N_25760);
nand U30240 (N_30240,N_25783,N_29607);
xor U30241 (N_30241,N_28584,N_26952);
xor U30242 (N_30242,N_28063,N_25211);
or U30243 (N_30243,N_26194,N_27863);
and U30244 (N_30244,N_29978,N_29859);
nor U30245 (N_30245,N_25936,N_26973);
nor U30246 (N_30246,N_29365,N_29129);
nand U30247 (N_30247,N_26836,N_29442);
or U30248 (N_30248,N_29861,N_28850);
nor U30249 (N_30249,N_27015,N_28334);
nand U30250 (N_30250,N_27212,N_27496);
nor U30251 (N_30251,N_26377,N_25399);
nand U30252 (N_30252,N_29981,N_27610);
nor U30253 (N_30253,N_28519,N_28718);
or U30254 (N_30254,N_28640,N_29726);
and U30255 (N_30255,N_25219,N_27316);
nand U30256 (N_30256,N_28333,N_26803);
nor U30257 (N_30257,N_26124,N_25801);
xor U30258 (N_30258,N_28178,N_25238);
and U30259 (N_30259,N_26739,N_25910);
nand U30260 (N_30260,N_27014,N_27218);
and U30261 (N_30261,N_28663,N_25348);
xnor U30262 (N_30262,N_27961,N_25032);
xor U30263 (N_30263,N_25279,N_29974);
and U30264 (N_30264,N_29499,N_26589);
nor U30265 (N_30265,N_27434,N_25357);
or U30266 (N_30266,N_29001,N_27060);
or U30267 (N_30267,N_28440,N_25943);
xnor U30268 (N_30268,N_27985,N_29382);
nor U30269 (N_30269,N_26051,N_26427);
nand U30270 (N_30270,N_28838,N_28045);
and U30271 (N_30271,N_28026,N_27957);
nand U30272 (N_30272,N_27114,N_27235);
xor U30273 (N_30273,N_25004,N_28487);
nand U30274 (N_30274,N_27701,N_26301);
nor U30275 (N_30275,N_27956,N_25237);
xor U30276 (N_30276,N_25270,N_29355);
xnor U30277 (N_30277,N_26688,N_25817);
nand U30278 (N_30278,N_25957,N_28696);
or U30279 (N_30279,N_28076,N_28747);
nand U30280 (N_30280,N_25347,N_29079);
nor U30281 (N_30281,N_27719,N_29420);
nor U30282 (N_30282,N_28798,N_28982);
and U30283 (N_30283,N_27718,N_26266);
nand U30284 (N_30284,N_28506,N_25266);
nor U30285 (N_30285,N_29248,N_29078);
and U30286 (N_30286,N_25545,N_27179);
and U30287 (N_30287,N_28529,N_27169);
xor U30288 (N_30288,N_25941,N_26698);
nor U30289 (N_30289,N_28998,N_25867);
or U30290 (N_30290,N_28699,N_27201);
nor U30291 (N_30291,N_26690,N_28503);
or U30292 (N_30292,N_29311,N_26913);
nor U30293 (N_30293,N_26990,N_26296);
nor U30294 (N_30294,N_28038,N_29931);
xor U30295 (N_30295,N_29908,N_27559);
nand U30296 (N_30296,N_25781,N_28818);
and U30297 (N_30297,N_25780,N_27558);
or U30298 (N_30298,N_28892,N_29977);
xor U30299 (N_30299,N_29807,N_27279);
xor U30300 (N_30300,N_25530,N_26705);
xnor U30301 (N_30301,N_25883,N_26587);
xor U30302 (N_30302,N_26532,N_29932);
or U30303 (N_30303,N_28027,N_25893);
xor U30304 (N_30304,N_29208,N_28420);
xor U30305 (N_30305,N_28645,N_26098);
nor U30306 (N_30306,N_25365,N_26734);
and U30307 (N_30307,N_26426,N_28160);
nor U30308 (N_30308,N_28840,N_25708);
and U30309 (N_30309,N_29563,N_25230);
nor U30310 (N_30310,N_28393,N_26155);
and U30311 (N_30311,N_25451,N_28675);
xor U30312 (N_30312,N_27541,N_27241);
nand U30313 (N_30313,N_27487,N_25727);
xnor U30314 (N_30314,N_26416,N_27998);
nor U30315 (N_30315,N_26789,N_27709);
or U30316 (N_30316,N_26531,N_28132);
xnor U30317 (N_30317,N_29456,N_29251);
nor U30318 (N_30318,N_25600,N_25610);
nand U30319 (N_30319,N_29140,N_29947);
nor U30320 (N_30320,N_27247,N_28108);
or U30321 (N_30321,N_26272,N_27184);
nor U30322 (N_30322,N_26320,N_26498);
and U30323 (N_30323,N_29758,N_27488);
nor U30324 (N_30324,N_25975,N_27236);
xor U30325 (N_30325,N_25296,N_29520);
nor U30326 (N_30326,N_27895,N_27342);
xnor U30327 (N_30327,N_29631,N_27960);
xor U30328 (N_30328,N_29372,N_28591);
xor U30329 (N_30329,N_28492,N_26812);
nand U30330 (N_30330,N_25778,N_25676);
nor U30331 (N_30331,N_29562,N_28930);
nand U30332 (N_30332,N_27089,N_28627);
and U30333 (N_30333,N_25643,N_25566);
or U30334 (N_30334,N_28859,N_26411);
nand U30335 (N_30335,N_26580,N_27951);
or U30336 (N_30336,N_29549,N_28648);
or U30337 (N_30337,N_27942,N_29274);
or U30338 (N_30338,N_27898,N_29709);
nand U30339 (N_30339,N_25812,N_29360);
and U30340 (N_30340,N_26466,N_25831);
nand U30341 (N_30341,N_28203,N_29821);
nor U30342 (N_30342,N_28339,N_25227);
xor U30343 (N_30343,N_27954,N_25134);
or U30344 (N_30344,N_25572,N_28463);
xnor U30345 (N_30345,N_27448,N_29408);
nand U30346 (N_30346,N_28601,N_29332);
nand U30347 (N_30347,N_28951,N_28399);
nand U30348 (N_30348,N_29335,N_25395);
xor U30349 (N_30349,N_26697,N_25038);
or U30350 (N_30350,N_25416,N_25400);
or U30351 (N_30351,N_29398,N_26547);
and U30352 (N_30352,N_28831,N_29088);
nand U30353 (N_30353,N_26854,N_26615);
xnor U30354 (N_30354,N_25925,N_29080);
xnor U30355 (N_30355,N_29999,N_25087);
nand U30356 (N_30356,N_27068,N_25204);
xor U30357 (N_30357,N_29490,N_28477);
xor U30358 (N_30358,N_25869,N_29897);
nand U30359 (N_30359,N_26733,N_25094);
nor U30360 (N_30360,N_29261,N_29096);
and U30361 (N_30361,N_29247,N_25672);
or U30362 (N_30362,N_27664,N_28371);
nor U30363 (N_30363,N_28290,N_29109);
nor U30364 (N_30364,N_25430,N_29229);
and U30365 (N_30365,N_27569,N_29308);
xnor U30366 (N_30366,N_28866,N_27940);
and U30367 (N_30367,N_27808,N_25756);
nand U30368 (N_30368,N_28105,N_28252);
or U30369 (N_30369,N_27395,N_27289);
xor U30370 (N_30370,N_25962,N_28829);
nand U30371 (N_30371,N_27639,N_28029);
xor U30372 (N_30372,N_27544,N_28050);
nand U30373 (N_30373,N_27318,N_26857);
xnor U30374 (N_30374,N_25023,N_26094);
nor U30375 (N_30375,N_27636,N_29865);
nor U30376 (N_30376,N_28015,N_29115);
xor U30377 (N_30377,N_25615,N_29776);
nor U30378 (N_30378,N_28535,N_27276);
nand U30379 (N_30379,N_26350,N_27684);
or U30380 (N_30380,N_27535,N_25758);
or U30381 (N_30381,N_26838,N_26027);
or U30382 (N_30382,N_25235,N_26957);
nand U30383 (N_30383,N_26823,N_29941);
or U30384 (N_30384,N_28559,N_25422);
and U30385 (N_30385,N_29568,N_25276);
and U30386 (N_30386,N_29930,N_29674);
or U30387 (N_30387,N_25320,N_29035);
or U30388 (N_30388,N_25587,N_27402);
nor U30389 (N_30389,N_26681,N_28003);
or U30390 (N_30390,N_26522,N_27346);
and U30391 (N_30391,N_29132,N_29023);
and U30392 (N_30392,N_27176,N_27598);
or U30393 (N_30393,N_25531,N_28327);
nor U30394 (N_30394,N_28799,N_28125);
or U30395 (N_30395,N_27376,N_29260);
xnor U30396 (N_30396,N_28451,N_29149);
nor U30397 (N_30397,N_25152,N_28096);
and U30398 (N_30398,N_27240,N_29683);
xnor U30399 (N_30399,N_28182,N_25967);
nand U30400 (N_30400,N_28300,N_29278);
and U30401 (N_30401,N_27676,N_27857);
or U30402 (N_30402,N_29959,N_27409);
nand U30403 (N_30403,N_27533,N_28836);
nand U30404 (N_30404,N_29569,N_27163);
nor U30405 (N_30405,N_26314,N_26417);
xor U30406 (N_30406,N_25895,N_26288);
and U30407 (N_30407,N_28963,N_29837);
nand U30408 (N_30408,N_26485,N_27847);
and U30409 (N_30409,N_25674,N_29671);
nand U30410 (N_30410,N_28822,N_26654);
nand U30411 (N_30411,N_28417,N_29222);
and U30412 (N_30412,N_28414,N_25837);
nor U30413 (N_30413,N_25265,N_29298);
xor U30414 (N_30414,N_29472,N_26581);
nor U30415 (N_30415,N_28556,N_25554);
xor U30416 (N_30416,N_28620,N_26383);
nand U30417 (N_30417,N_29956,N_27343);
xnor U30418 (N_30418,N_29026,N_27914);
nand U30419 (N_30419,N_25696,N_25924);
xnor U30420 (N_30420,N_27849,N_29878);
nor U30421 (N_30421,N_27751,N_29152);
and U30422 (N_30422,N_29273,N_25285);
and U30423 (N_30423,N_28039,N_25128);
nand U30424 (N_30424,N_27572,N_29526);
xor U30425 (N_30425,N_26040,N_28693);
nor U30426 (N_30426,N_26527,N_25616);
nand U30427 (N_30427,N_25173,N_28682);
xnor U30428 (N_30428,N_28589,N_29505);
nor U30429 (N_30429,N_29346,N_27310);
xor U30430 (N_30430,N_25636,N_26076);
nor U30431 (N_30431,N_25171,N_25860);
or U30432 (N_30432,N_29236,N_27905);
nor U30433 (N_30433,N_26323,N_27309);
or U30434 (N_30434,N_29532,N_29077);
and U30435 (N_30435,N_28092,N_25774);
and U30436 (N_30436,N_25614,N_27422);
xnor U30437 (N_30437,N_27322,N_28335);
nor U30438 (N_30438,N_28378,N_28243);
nor U30439 (N_30439,N_27107,N_26662);
and U30440 (N_30440,N_28176,N_26657);
xor U30441 (N_30441,N_28989,N_28984);
nor U30442 (N_30442,N_29439,N_26452);
nor U30443 (N_30443,N_29018,N_29920);
nor U30444 (N_30444,N_26031,N_28369);
and U30445 (N_30445,N_25503,N_25948);
xor U30446 (N_30446,N_29590,N_29849);
or U30447 (N_30447,N_27220,N_27010);
or U30448 (N_30448,N_29326,N_25859);
nor U30449 (N_30449,N_27711,N_28733);
and U30450 (N_30450,N_29694,N_27165);
nor U30451 (N_30451,N_27738,N_29230);
nand U30452 (N_30452,N_25880,N_27504);
xor U30453 (N_30453,N_26046,N_26745);
and U30454 (N_30454,N_29210,N_26458);
or U30455 (N_30455,N_26209,N_28249);
nand U30456 (N_30456,N_28204,N_27740);
nor U30457 (N_30457,N_25260,N_26833);
and U30458 (N_30458,N_26503,N_25077);
or U30459 (N_30459,N_25026,N_27904);
or U30460 (N_30460,N_29618,N_26398);
or U30461 (N_30461,N_26709,N_25294);
nand U30462 (N_30462,N_25821,N_28312);
or U30463 (N_30463,N_25050,N_29271);
nor U30464 (N_30464,N_29808,N_25682);
and U30465 (N_30465,N_28792,N_27980);
and U30466 (N_30466,N_29463,N_25148);
nor U30467 (N_30467,N_26840,N_28857);
nor U30468 (N_30468,N_28067,N_27824);
or U30469 (N_30469,N_28397,N_29806);
and U30470 (N_30470,N_26382,N_28916);
xnor U30471 (N_30471,N_28360,N_29292);
nand U30472 (N_30472,N_29093,N_28169);
xnor U30473 (N_30473,N_26327,N_27698);
nand U30474 (N_30474,N_29642,N_27924);
nor U30475 (N_30475,N_26175,N_26855);
nand U30476 (N_30476,N_28073,N_29983);
and U30477 (N_30477,N_25848,N_28744);
xor U30478 (N_30478,N_29509,N_28549);
xnor U30479 (N_30479,N_25989,N_25199);
nor U30480 (N_30480,N_26738,N_29262);
and U30481 (N_30481,N_29190,N_29361);
nand U30482 (N_30482,N_28650,N_28844);
xor U30483 (N_30483,N_28713,N_25513);
xor U30484 (N_30484,N_25141,N_28961);
nor U30485 (N_30485,N_26437,N_26508);
and U30486 (N_30486,N_25011,N_25678);
or U30487 (N_30487,N_26831,N_27939);
nor U30488 (N_30488,N_25586,N_25664);
and U30489 (N_30489,N_26351,N_25517);
or U30490 (N_30490,N_25378,N_29348);
nand U30491 (N_30491,N_29468,N_28426);
nor U30492 (N_30492,N_25169,N_27590);
nand U30493 (N_30493,N_25769,N_27773);
nand U30494 (N_30494,N_27135,N_25157);
xor U30495 (N_30495,N_25570,N_27560);
and U30496 (N_30496,N_28572,N_25424);
and U30497 (N_30497,N_27903,N_28520);
xnor U30498 (N_30498,N_26020,N_29102);
nand U30499 (N_30499,N_28561,N_25949);
xnor U30500 (N_30500,N_26079,N_26955);
or U30501 (N_30501,N_26077,N_29712);
or U30502 (N_30502,N_27999,N_26325);
xnor U30503 (N_30503,N_26271,N_29676);
or U30504 (N_30504,N_29433,N_27314);
xnor U30505 (N_30505,N_25256,N_28692);
nor U30506 (N_30506,N_29557,N_26944);
xor U30507 (N_30507,N_29823,N_29945);
xor U30508 (N_30508,N_27654,N_27748);
nor U30509 (N_30509,N_26262,N_28684);
xor U30510 (N_30510,N_26706,N_27779);
or U30511 (N_30511,N_27879,N_26067);
and U30512 (N_30512,N_27147,N_27780);
nor U30513 (N_30513,N_28405,N_29126);
nor U30514 (N_30514,N_27804,N_25218);
nor U30515 (N_30515,N_28867,N_29270);
nor U30516 (N_30516,N_26287,N_26773);
xor U30517 (N_30517,N_26198,N_29901);
nor U30518 (N_30518,N_27173,N_27152);
and U30519 (N_30519,N_28931,N_27627);
xnor U30520 (N_30520,N_29253,N_29434);
nand U30521 (N_30521,N_29522,N_25852);
or U30522 (N_30522,N_27607,N_26462);
or U30523 (N_30523,N_27689,N_26156);
and U30524 (N_30524,N_26771,N_28958);
or U30525 (N_30525,N_27238,N_27265);
or U30526 (N_30526,N_27193,N_28973);
nand U30527 (N_30527,N_27003,N_29535);
nor U30528 (N_30528,N_27379,N_27626);
and U30529 (N_30529,N_29733,N_26608);
or U30530 (N_30530,N_25777,N_28863);
or U30531 (N_30531,N_25030,N_27297);
or U30532 (N_30532,N_28286,N_28064);
nand U30533 (N_30533,N_26607,N_28135);
nor U30534 (N_30534,N_29400,N_28202);
or U30535 (N_30535,N_29283,N_27935);
nor U30536 (N_30536,N_26041,N_28211);
or U30537 (N_30537,N_26391,N_26331);
nand U30538 (N_30538,N_25591,N_27793);
nor U30539 (N_30539,N_25063,N_25797);
xnor U30540 (N_30540,N_26022,N_26333);
nand U30541 (N_30541,N_26817,N_27958);
xor U30542 (N_30542,N_28906,N_25489);
nand U30543 (N_30543,N_29789,N_27026);
nor U30544 (N_30544,N_26985,N_29199);
nor U30545 (N_30545,N_29943,N_29818);
or U30546 (N_30546,N_25160,N_26029);
or U30547 (N_30547,N_26559,N_27393);
or U30548 (N_30548,N_28938,N_28126);
or U30549 (N_30549,N_26920,N_26361);
or U30550 (N_30550,N_25703,N_25232);
nor U30551 (N_30551,N_26804,N_29844);
nand U30552 (N_30552,N_27944,N_29907);
nor U30553 (N_30553,N_26760,N_25452);
xor U30554 (N_30554,N_29760,N_28240);
nor U30555 (N_30555,N_29288,N_28749);
or U30556 (N_30556,N_28670,N_28538);
or U30557 (N_30557,N_27693,N_25239);
nand U30558 (N_30558,N_29551,N_29976);
xor U30559 (N_30559,N_26392,N_29148);
xnor U30560 (N_30560,N_28422,N_25201);
xor U30561 (N_30561,N_27185,N_29857);
xor U30562 (N_30562,N_25138,N_29581);
xnor U30563 (N_30563,N_28113,N_27506);
nor U30564 (N_30564,N_26919,N_28560);
nand U30565 (N_30565,N_26055,N_25012);
xor U30566 (N_30566,N_26343,N_28075);
and U30567 (N_30567,N_25033,N_28768);
nor U30568 (N_30568,N_28647,N_29534);
nand U30569 (N_30569,N_28320,N_27652);
xnor U30570 (N_30570,N_27691,N_25619);
nand U30571 (N_30571,N_26829,N_29385);
nand U30572 (N_30572,N_25415,N_27622);
and U30573 (N_30573,N_28301,N_27327);
or U30574 (N_30574,N_29048,N_26885);
xnor U30575 (N_30575,N_29929,N_29727);
or U30576 (N_30576,N_26663,N_25963);
nor U30577 (N_30577,N_28077,N_27194);
xnor U30578 (N_30578,N_27521,N_25577);
xor U30579 (N_30579,N_25222,N_28390);
or U30580 (N_30580,N_26669,N_29123);
xnor U30581 (N_30581,N_28146,N_27129);
xnor U30582 (N_30582,N_27067,N_27330);
or U30583 (N_30583,N_25208,N_29953);
nor U30584 (N_30584,N_26859,N_25051);
nand U30585 (N_30585,N_28141,N_27729);
xor U30586 (N_30586,N_29307,N_25109);
or U30587 (N_30587,N_28021,N_28494);
or U30588 (N_30588,N_26065,N_27302);
xor U30589 (N_30589,N_26748,N_29816);
xor U30590 (N_30590,N_26216,N_29660);
xor U30591 (N_30591,N_27805,N_28686);
or U30592 (N_30592,N_27583,N_29363);
xnor U30593 (N_30593,N_28386,N_28444);
or U30594 (N_30594,N_26090,N_25548);
xor U30595 (N_30595,N_27100,N_28165);
nand U30596 (N_30596,N_29634,N_27534);
nor U30597 (N_30597,N_27971,N_26670);
or U30598 (N_30598,N_29391,N_28917);
nor U30599 (N_30599,N_28537,N_26951);
xnor U30600 (N_30600,N_27476,N_27889);
or U30601 (N_30601,N_29407,N_27281);
and U30602 (N_30602,N_29996,N_26335);
xor U30603 (N_30603,N_29029,N_28656);
nand U30604 (N_30604,N_25166,N_26666);
or U30605 (N_30605,N_26158,N_25118);
nand U30606 (N_30606,N_29373,N_26092);
nor U30607 (N_30607,N_27768,N_25001);
xor U30608 (N_30608,N_25069,N_26215);
nand U30609 (N_30609,N_28172,N_26316);
or U30610 (N_30610,N_29998,N_27024);
xnor U30611 (N_30611,N_29055,N_28016);
nor U30612 (N_30612,N_25709,N_26661);
nand U30613 (N_30613,N_27091,N_27451);
and U30614 (N_30614,N_29529,N_28813);
nand U30615 (N_30615,N_25333,N_25828);
xnor U30616 (N_30616,N_28815,N_26300);
and U30617 (N_30617,N_28687,N_29312);
nand U30618 (N_30618,N_27001,N_25460);
xnor U30619 (N_30619,N_28133,N_25744);
nor U30620 (N_30620,N_28277,N_28002);
xor U30621 (N_30621,N_26475,N_26884);
xnor U30622 (N_30622,N_29470,N_25690);
xor U30623 (N_30623,N_27036,N_26477);
and U30624 (N_30624,N_27045,N_27388);
nor U30625 (N_30625,N_26512,N_27252);
and U30626 (N_30626,N_28904,N_28037);
or U30627 (N_30627,N_28151,N_26624);
nand U30628 (N_30628,N_25991,N_26641);
xnor U30629 (N_30629,N_29378,N_26588);
or U30630 (N_30630,N_26758,N_26535);
nand U30631 (N_30631,N_28022,N_25132);
or U30632 (N_30632,N_26444,N_25492);
nand U30633 (N_30633,N_27075,N_25955);
nand U30634 (N_30634,N_28442,N_27708);
or U30635 (N_30635,N_27554,N_27690);
nor U30636 (N_30636,N_25805,N_26143);
or U30637 (N_30637,N_28708,N_25808);
xor U30638 (N_30638,N_28590,N_27631);
and U30639 (N_30639,N_27617,N_29666);
and U30640 (N_30640,N_26815,N_29445);
and U30641 (N_30641,N_28257,N_25663);
nor U30642 (N_30642,N_27110,N_28564);
nand U30643 (N_30643,N_28122,N_25475);
nor U30644 (N_30644,N_25246,N_28343);
or U30645 (N_30645,N_25334,N_29624);
and U30646 (N_30646,N_27587,N_25292);
and U30647 (N_30647,N_27878,N_27392);
xnor U30648 (N_30648,N_27144,N_27463);
nand U30649 (N_30649,N_29973,N_29575);
nor U30650 (N_30650,N_26116,N_26490);
nor U30651 (N_30651,N_29112,N_29366);
nor U30652 (N_30652,N_25979,N_25163);
xor U30653 (N_30653,N_28880,N_28266);
nor U30654 (N_30654,N_29178,N_27177);
nor U30655 (N_30655,N_27655,N_28232);
and U30656 (N_30656,N_28152,N_29147);
or U30657 (N_30657,N_28896,N_27526);
nor U30658 (N_30658,N_26894,N_27397);
xor U30659 (N_30659,N_27065,N_27284);
xor U30660 (N_30660,N_26464,N_27982);
nand U30661 (N_30661,N_25719,N_25473);
and U30662 (N_30662,N_29718,N_26843);
nand U30663 (N_30663,N_26342,N_27828);
nor U30664 (N_30664,N_27365,N_25691);
nor U30665 (N_30665,N_26557,N_29637);
xor U30666 (N_30666,N_26584,N_27261);
and U30667 (N_30667,N_27071,N_28638);
xnor U30668 (N_30668,N_29574,N_25449);
nor U30669 (N_30669,N_28116,N_26809);
nand U30670 (N_30670,N_26969,N_29834);
or U30671 (N_30671,N_29380,N_27430);
or U30672 (N_30672,N_29898,N_25342);
nor U30673 (N_30673,N_28909,N_26742);
or U30674 (N_30674,N_28190,N_26127);
nand U30675 (N_30675,N_29516,N_25908);
xor U30676 (N_30676,N_26019,N_28307);
and U30677 (N_30677,N_28571,N_27203);
nor U30678 (N_30678,N_28834,N_29314);
and U30679 (N_30679,N_26769,N_28737);
xnor U30680 (N_30680,N_27609,N_25182);
nor U30681 (N_30681,N_28367,N_29041);
nor U30682 (N_30682,N_28434,N_29935);
or U30683 (N_30683,N_29955,N_25872);
xnor U30684 (N_30684,N_28419,N_25198);
or U30685 (N_30685,N_29244,N_26455);
nand U30686 (N_30686,N_25579,N_26647);
nor U30687 (N_30687,N_27019,N_27818);
nor U30688 (N_30688,N_29668,N_26026);
nand U30689 (N_30689,N_25108,N_27292);
nand U30690 (N_30690,N_27934,N_28275);
xor U30691 (N_30691,N_28706,N_26710);
or U30692 (N_30692,N_29345,N_25481);
or U30693 (N_30693,N_27133,N_26231);
xor U30694 (N_30694,N_28625,N_25662);
nand U30695 (N_30695,N_26991,N_28597);
nand U30696 (N_30696,N_26892,N_28881);
nor U30697 (N_30697,N_29002,N_28009);
nor U30698 (N_30698,N_29950,N_25510);
and U30699 (N_30699,N_28156,N_28913);
and U30700 (N_30700,N_26924,N_25770);
or U30701 (N_30701,N_25862,N_27734);
xor U30702 (N_30702,N_25576,N_25914);
or U30703 (N_30703,N_27323,N_29256);
nand U30704 (N_30704,N_27436,N_27171);
or U30705 (N_30705,N_29141,N_26783);
or U30706 (N_30706,N_25626,N_28662);
xnor U30707 (N_30707,N_29393,N_25303);
xor U30708 (N_30708,N_28731,N_29396);
nand U30709 (N_30709,N_27705,N_27710);
nand U30710 (N_30710,N_29105,N_29095);
nor U30711 (N_30711,N_26713,N_25251);
nand U30712 (N_30712,N_26218,N_28767);
and U30713 (N_30713,N_28510,N_26927);
or U30714 (N_30714,N_29182,N_29128);
and U30715 (N_30715,N_25024,N_28926);
or U30716 (N_30716,N_26877,N_25997);
or U30717 (N_30717,N_28396,N_25317);
and U30718 (N_30718,N_26400,N_27127);
nand U30719 (N_30719,N_29577,N_28615);
or U30720 (N_30720,N_25768,N_29124);
or U30721 (N_30721,N_29698,N_29167);
nor U30722 (N_30722,N_28363,N_27539);
or U30723 (N_30723,N_27513,N_28119);
nand U30724 (N_30724,N_28255,N_26793);
or U30725 (N_30725,N_29188,N_27124);
nand U30726 (N_30726,N_26364,N_25668);
xor U30727 (N_30727,N_26737,N_27105);
and U30728 (N_30728,N_29536,N_26304);
and U30729 (N_30729,N_29194,N_29168);
xor U30730 (N_30730,N_27215,N_28933);
nand U30731 (N_30731,N_27433,N_28715);
or U30732 (N_30732,N_29721,N_25006);
xor U30733 (N_30733,N_29906,N_29275);
nand U30734 (N_30734,N_28606,N_25806);
and U30735 (N_30735,N_28004,N_27025);
or U30736 (N_30736,N_29492,N_25159);
and U30737 (N_30737,N_29062,N_26616);
xnor U30738 (N_30738,N_28311,N_26043);
and U30739 (N_30739,N_26572,N_26898);
or U30740 (N_30740,N_27154,N_26188);
and U30741 (N_30741,N_29226,N_27441);
or U30742 (N_30742,N_29068,N_28317);
nor U30743 (N_30743,N_28899,N_29586);
nor U30744 (N_30744,N_29290,N_29485);
and U30745 (N_30745,N_28523,N_29625);
xor U30746 (N_30746,N_26901,N_26558);
and U30747 (N_30747,N_29430,N_25580);
and U30748 (N_30748,N_27331,N_27263);
or U30749 (N_30749,N_25268,N_25630);
nor U30750 (N_30750,N_28179,N_27902);
nor U30751 (N_30751,N_25267,N_27027);
xor U30752 (N_30752,N_26942,N_25512);
or U30753 (N_30753,N_29795,N_27283);
nand U30754 (N_30754,N_29848,N_29802);
xnor U30755 (N_30755,N_26367,N_27868);
and U30756 (N_30756,N_26759,N_26071);
nor U30757 (N_30757,N_25764,N_28539);
and U30758 (N_30758,N_27317,N_25119);
xor U30759 (N_30759,N_28149,N_29804);
nor U30760 (N_30760,N_26097,N_26394);
xor U30761 (N_30761,N_25624,N_28234);
xnor U30762 (N_30762,N_25882,N_29427);
or U30763 (N_30763,N_28895,N_29473);
or U30764 (N_30764,N_26635,N_26480);
xor U30765 (N_30765,N_27792,N_28145);
nand U30766 (N_30766,N_25968,N_25929);
nand U30767 (N_30767,N_26203,N_26408);
nor U30768 (N_30768,N_26775,N_29057);
xor U30769 (N_30769,N_28258,N_26312);
xnor U30770 (N_30770,N_26640,N_29235);
and U30771 (N_30771,N_28604,N_28769);
xor U30772 (N_30772,N_25330,N_27187);
or U30773 (N_30773,N_25083,N_27134);
nand U30774 (N_30774,N_29539,N_25428);
or U30775 (N_30775,N_27022,N_28732);
nor U30776 (N_30776,N_29757,N_28128);
nor U30777 (N_30777,N_29934,N_28893);
xor U30778 (N_30778,N_29351,N_25519);
or U30779 (N_30779,N_26606,N_29154);
xnor U30780 (N_30780,N_28902,N_26541);
or U30781 (N_30781,N_27989,N_28944);
nand U30782 (N_30782,N_25145,N_29227);
and U30783 (N_30783,N_27275,N_26294);
or U30784 (N_30784,N_26496,N_26206);
or U30785 (N_30785,N_29681,N_28407);
or U30786 (N_30786,N_26310,N_26208);
and U30787 (N_30787,N_26623,N_28826);
nor U30788 (N_30788,N_26566,N_26474);
xnor U30789 (N_30789,N_29313,N_29053);
nor U30790 (N_30790,N_28710,N_29923);
or U30791 (N_30791,N_28355,N_28791);
nor U30792 (N_30792,N_28196,N_27862);
xnor U30793 (N_30793,N_25813,N_28903);
xnor U30794 (N_30794,N_26389,N_28697);
xor U30795 (N_30795,N_26534,N_27795);
nor U30796 (N_30796,N_28621,N_28901);
and U30797 (N_30797,N_29610,N_26191);
and U30798 (N_30798,N_28521,N_26413);
or U30799 (N_30799,N_28782,N_25405);
and U30800 (N_30800,N_29330,N_26945);
and U30801 (N_30801,N_25995,N_26180);
or U30802 (N_30802,N_28384,N_26178);
nor U30803 (N_30803,N_29081,N_27637);
nor U30804 (N_30804,N_28566,N_28667);
nand U30805 (N_30805,N_26751,N_26123);
or U30806 (N_30806,N_25126,N_25757);
or U30807 (N_30807,N_28576,N_25111);
and U30808 (N_30808,N_29749,N_27396);
nor U30809 (N_30809,N_29649,N_29357);
xnor U30810 (N_30810,N_26182,N_28629);
nor U30811 (N_30811,N_27696,N_29883);
xor U30812 (N_30812,N_27928,N_25816);
and U30813 (N_30813,N_25440,N_29309);
nand U30814 (N_30814,N_29719,N_25715);
xor U30815 (N_30815,N_26552,N_26863);
or U30816 (N_30816,N_28162,N_25463);
xor U30817 (N_30817,N_25421,N_28382);
or U30818 (N_30818,N_28383,N_28177);
nand U30819 (N_30819,N_26441,N_27401);
nor U30820 (N_30820,N_29665,N_26190);
nand U30821 (N_30821,N_25288,N_25085);
xnor U30822 (N_30822,N_27157,N_26495);
nor U30823 (N_30823,N_27875,N_25645);
and U30824 (N_30824,N_28425,N_27910);
xnor U30825 (N_30825,N_26109,N_25262);
nor U30826 (N_30826,N_25532,N_27992);
nand U30827 (N_30827,N_25811,N_28514);
nand U30828 (N_30828,N_25382,N_25595);
and U30829 (N_30829,N_29900,N_28467);
nand U30830 (N_30830,N_29225,N_27658);
nand U30831 (N_30831,N_28763,N_26891);
nand U30832 (N_30832,N_25495,N_29803);
and U30833 (N_30833,N_29155,N_25234);
nand U30834 (N_30834,N_27799,N_29003);
nor U30835 (N_30835,N_28762,N_25504);
or U30836 (N_30836,N_26151,N_28527);
or U30837 (N_30837,N_29623,N_29090);
nor U30838 (N_30838,N_25380,N_26826);
nor U30839 (N_30839,N_25341,N_29477);
nor U30840 (N_30840,N_26192,N_27304);
nand U30841 (N_30841,N_25901,N_27606);
nand U30842 (N_30842,N_28910,N_26757);
or U30843 (N_30843,N_29843,N_27564);
or U30844 (N_30844,N_26499,N_29166);
and U30845 (N_30845,N_29729,N_25840);
nor U30846 (N_30846,N_29690,N_27399);
xor U30847 (N_30847,N_26575,N_27338);
or U30848 (N_30848,N_28631,N_27537);
nor U30849 (N_30849,N_26975,N_28465);
xnor U30850 (N_30850,N_25980,N_27510);
and U30851 (N_30851,N_28069,N_27575);
nand U30852 (N_30852,N_25602,N_28634);
nor U30853 (N_30853,N_28233,N_29493);
and U30854 (N_30854,N_26850,N_28241);
nand U30855 (N_30855,N_26523,N_25328);
and U30856 (N_30856,N_25324,N_29216);
xnor U30857 (N_30857,N_28872,N_27881);
and U30858 (N_30858,N_28001,N_28385);
xnor U30859 (N_30859,N_29616,N_26867);
or U30860 (N_30860,N_26388,N_29541);
nand U30861 (N_30861,N_29601,N_25439);
nand U30862 (N_30862,N_29158,N_28683);
and U30863 (N_30863,N_27620,N_28285);
or U30864 (N_30864,N_28869,N_28974);
nor U30865 (N_30865,N_29413,N_26755);
nand U30866 (N_30866,N_26984,N_27499);
and U30867 (N_30867,N_25558,N_29323);
or U30868 (N_30868,N_29890,N_26450);
and U30869 (N_30869,N_25340,N_26852);
nand U30870 (N_30870,N_28328,N_29630);
or U30871 (N_30871,N_29747,N_29567);
nor U30872 (N_30872,N_28238,N_25107);
nand U30873 (N_30873,N_27044,N_26525);
or U30874 (N_30874,N_25371,N_26308);
nand U30875 (N_30875,N_25478,N_27298);
or U30876 (N_30876,N_25002,N_27747);
nand U30877 (N_30877,N_29588,N_26282);
or U30878 (N_30878,N_25861,N_25665);
xnor U30879 (N_30879,N_27249,N_25287);
xor U30880 (N_30880,N_28342,N_25877);
xor U30881 (N_30881,N_25597,N_25453);
and U30882 (N_30882,N_26719,N_25734);
or U30883 (N_30883,N_29171,N_27832);
or U30884 (N_30884,N_29638,N_28470);
nand U30885 (N_30885,N_26570,N_29025);
and U30886 (N_30886,N_26146,N_25596);
nor U30887 (N_30887,N_25282,N_29994);
xor U30888 (N_30888,N_25653,N_29828);
and U30889 (N_30889,N_28181,N_25406);
nand U30890 (N_30890,N_28526,N_29957);
nand U30891 (N_30891,N_26660,N_29316);
or U30892 (N_30892,N_25441,N_25561);
nand U30893 (N_30893,N_27162,N_26774);
nor U30894 (N_30894,N_26380,N_26746);
nor U30895 (N_30895,N_27037,N_25254);
nor U30896 (N_30896,N_25018,N_25656);
and U30897 (N_30897,N_25047,N_27625);
or U30898 (N_30898,N_26375,N_25755);
xor U30899 (N_30899,N_28086,N_28187);
nor U30900 (N_30900,N_28644,N_25309);
nor U30901 (N_30901,N_26258,N_29305);
or U30902 (N_30902,N_27012,N_29604);
and U30903 (N_30903,N_27226,N_27180);
xnor U30904 (N_30904,N_27158,N_26792);
or U30905 (N_30905,N_26318,N_27516);
nand U30906 (N_30906,N_25325,N_28137);
xnor U30907 (N_30907,N_28438,N_29234);
nor U30908 (N_30908,N_29742,N_25670);
nor U30909 (N_30909,N_29737,N_29553);
nor U30910 (N_30910,N_25429,N_27873);
or U30911 (N_30911,N_28264,N_29324);
xor U30912 (N_30912,N_25835,N_25969);
and U30913 (N_30913,N_29571,N_28051);
xor U30914 (N_30914,N_29530,N_27072);
nand U30915 (N_30915,N_26750,N_28099);
nor U30916 (N_30916,N_29617,N_26243);
nand U30917 (N_30917,N_26423,N_26981);
nor U30918 (N_30918,N_27650,N_25907);
or U30919 (N_30919,N_27477,N_28094);
and U30920 (N_30920,N_28505,N_26306);
nor U30921 (N_30921,N_27816,N_27325);
or U30922 (N_30922,N_25020,N_27253);
nor U30923 (N_30923,N_25027,N_27485);
nor U30924 (N_30924,N_26048,N_25386);
or U30925 (N_30925,N_26061,N_26636);
nand U30926 (N_30926,N_28484,N_26032);
xor U30927 (N_30927,N_26585,N_29017);
or U30928 (N_30928,N_29942,N_29893);
or U30929 (N_30929,N_27744,N_27511);
or U30930 (N_30930,N_29927,N_27483);
and U30931 (N_30931,N_25986,N_26073);
xor U30932 (N_30932,N_28402,N_27336);
or U30933 (N_30933,N_26005,N_28779);
nor U30934 (N_30934,N_27937,N_28658);
or U30935 (N_30935,N_25180,N_25402);
and U30936 (N_30936,N_27965,N_26772);
and U30937 (N_30937,N_26467,N_29756);
nor U30938 (N_30938,N_28500,N_29783);
nor U30939 (N_30939,N_28297,N_27945);
nand U30940 (N_30940,N_29964,N_27006);
and U30941 (N_30941,N_27051,N_25802);
nor U30942 (N_30942,N_27077,N_26518);
or U30943 (N_30943,N_25187,N_25858);
nand U30944 (N_30944,N_28665,N_27256);
xor U30945 (N_30945,N_29566,N_27915);
nor U30946 (N_30946,N_28877,N_29673);
nor U30947 (N_30947,N_25789,N_28013);
nand U30948 (N_30948,N_29651,N_25355);
nor U30949 (N_30949,N_25695,N_28025);
and U30950 (N_30950,N_25154,N_28609);
and U30951 (N_30951,N_26153,N_27131);
or U30952 (N_30952,N_25131,N_28011);
or U30953 (N_30953,N_28448,N_29131);
or U30954 (N_30954,N_25436,N_27479);
xnor U30955 (N_30955,N_25660,N_29771);
xor U30956 (N_30956,N_25312,N_25068);
or U30957 (N_30957,N_29595,N_27313);
nor U30958 (N_30958,N_29933,N_29282);
nor U30959 (N_30959,N_28805,N_28900);
nor U30960 (N_30960,N_29089,N_27762);
and U30961 (N_30961,N_29369,N_25921);
or U30962 (N_30962,N_27756,N_26554);
or U30963 (N_30963,N_26784,N_25892);
nor U30964 (N_30964,N_27896,N_28457);
nor U30965 (N_30965,N_26261,N_29451);
nor U30966 (N_30966,N_26352,N_27291);
and U30967 (N_30967,N_28851,N_26360);
nor U30968 (N_30968,N_28408,N_25494);
xnor U30969 (N_30969,N_25638,N_27761);
xor U30970 (N_30970,N_27404,N_28812);
and U30971 (N_30971,N_25724,N_28748);
and U30972 (N_30972,N_25827,N_26949);
nand U30973 (N_30973,N_29829,N_27929);
nand U30974 (N_30974,N_28624,N_25547);
nand U30975 (N_30975,N_29428,N_27827);
or U30976 (N_30976,N_28231,N_26896);
nor U30977 (N_30977,N_27542,N_25074);
nand U30978 (N_30978,N_28410,N_28960);
nand U30979 (N_30979,N_29327,N_25557);
nor U30980 (N_30980,N_28639,N_29854);
nand U30981 (N_30981,N_26471,N_27720);
xor U30982 (N_30982,N_26947,N_29565);
nor U30983 (N_30983,N_26520,N_26269);
xnor U30984 (N_30984,N_28324,N_27000);
nor U30985 (N_30985,N_25589,N_25932);
or U30986 (N_30986,N_27486,N_28649);
or U30987 (N_30987,N_26841,N_29548);
nand U30988 (N_30988,N_26528,N_26727);
nor U30989 (N_30989,N_29005,N_28954);
or U30990 (N_30990,N_28855,N_26667);
xnor U30991 (N_30991,N_28935,N_25274);
and U30992 (N_30992,N_29979,N_25370);
xor U30993 (N_30993,N_27796,N_25259);
xor U30994 (N_30994,N_25091,N_27123);
nand U30995 (N_30995,N_26371,N_28449);
or U30996 (N_30996,N_26908,N_27443);
nand U30997 (N_30997,N_28678,N_25585);
or U30998 (N_30998,N_27920,N_28719);
xor U30999 (N_30999,N_28142,N_27789);
nand U31000 (N_31000,N_26988,N_26149);
or U31001 (N_31001,N_27641,N_28586);
xnor U31002 (N_31002,N_27682,N_29240);
or U31003 (N_31003,N_27207,N_29340);
nand U31004 (N_31004,N_29364,N_28443);
xor U31005 (N_31005,N_28956,N_27557);
xor U31006 (N_31006,N_26433,N_28427);
and U31007 (N_31007,N_26393,N_25306);
nand U31008 (N_31008,N_29180,N_28466);
nor U31009 (N_31009,N_27836,N_26217);
or U31010 (N_31010,N_27228,N_27766);
xor U31011 (N_31011,N_26630,N_27608);
nand U31012 (N_31012,N_29052,N_29917);
nand U31013 (N_31013,N_26196,N_27150);
xor U31014 (N_31014,N_27446,N_25844);
or U31015 (N_31015,N_27271,N_29495);
or U31016 (N_31016,N_25978,N_28753);
and U31017 (N_31017,N_29232,N_26057);
nand U31018 (N_31018,N_26780,N_29421);
and U31019 (N_31019,N_29769,N_27491);
nor U31020 (N_31020,N_28008,N_28995);
or U31021 (N_31021,N_28879,N_29218);
and U31022 (N_31022,N_26911,N_27921);
xnor U31023 (N_31023,N_28100,N_27930);
nand U31024 (N_31024,N_27728,N_26403);
xnor U31025 (N_31025,N_28251,N_27576);
or U31026 (N_31026,N_26502,N_29847);
xnor U31027 (N_31027,N_26967,N_27385);
xnor U31028 (N_31028,N_26211,N_28296);
xor U31029 (N_31029,N_27258,N_25275);
nor U31030 (N_31030,N_29728,N_25736);
or U31031 (N_31031,N_26016,N_28929);
or U31032 (N_31032,N_27175,N_27018);
nor U31033 (N_31033,N_26878,N_29049);
nand U31034 (N_31034,N_29889,N_29710);
xnor U31035 (N_31035,N_25098,N_28534);
xor U31036 (N_31036,N_26551,N_26717);
and U31037 (N_31037,N_29195,N_29860);
nor U31038 (N_31038,N_25706,N_26599);
xnor U31039 (N_31039,N_29338,N_25448);
or U31040 (N_31040,N_28134,N_29640);
or U31041 (N_31041,N_29339,N_29653);
nand U31042 (N_31042,N_28081,N_25271);
nand U31043 (N_31043,N_29402,N_25658);
and U31044 (N_31044,N_28413,N_25322);
and U31045 (N_31045,N_27668,N_27913);
nor U31046 (N_31046,N_27700,N_29951);
xor U31047 (N_31047,N_28788,N_26359);
xor U31048 (N_31048,N_27389,N_26096);
nor U31049 (N_31049,N_25290,N_26671);
or U31050 (N_31050,N_26399,N_26072);
and U31051 (N_31051,N_29467,N_29644);
xnor U31052 (N_31052,N_26972,N_25261);
xnor U31053 (N_31053,N_27842,N_28415);
or U31054 (N_31054,N_28659,N_26553);
nand U31055 (N_31055,N_25244,N_26940);
nand U31056 (N_31056,N_27893,N_26813);
xnor U31057 (N_31057,N_27421,N_28437);
nand U31058 (N_31058,N_25987,N_29238);
and U31059 (N_31059,N_29435,N_25920);
or U31060 (N_31060,N_26997,N_27507);
and U31061 (N_31061,N_28418,N_28603);
or U31062 (N_31062,N_29636,N_28388);
xor U31063 (N_31063,N_28946,N_26226);
or U31064 (N_31064,N_28789,N_26284);
and U31065 (N_31065,N_26171,N_28932);
or U31066 (N_31066,N_25443,N_27613);
xnor U31067 (N_31067,N_27030,N_27428);
xnor U31068 (N_31068,N_26989,N_28282);
and U31069 (N_31069,N_29700,N_27615);
nor U31070 (N_31070,N_28979,N_27119);
or U31071 (N_31071,N_27041,N_28823);
and U31072 (N_31072,N_26732,N_27508);
xnor U31073 (N_31073,N_26313,N_27648);
xor U31074 (N_31074,N_27679,N_26340);
and U31075 (N_31075,N_25064,N_26808);
or U31076 (N_31076,N_27686,N_28483);
or U31077 (N_31077,N_28248,N_25162);
and U31078 (N_31078,N_26207,N_29995);
nand U31079 (N_31079,N_27611,N_28260);
xnor U31080 (N_31080,N_27109,N_29186);
or U31081 (N_31081,N_29061,N_25393);
xnor U31082 (N_31082,N_27355,N_27619);
nor U31083 (N_31083,N_25167,N_29241);
xnor U31084 (N_31084,N_26730,N_28280);
nand U31085 (N_31085,N_29611,N_29916);
or U31086 (N_31086,N_29778,N_27716);
xnor U31087 (N_31087,N_27855,N_27574);
nand U31088 (N_31088,N_25501,N_26939);
xor U31089 (N_31089,N_27326,N_25384);
and U31090 (N_31090,N_25799,N_27372);
or U31091 (N_31091,N_28362,N_28295);
and U31092 (N_31092,N_26276,N_29851);
nand U31093 (N_31093,N_28112,N_28971);
or U31094 (N_31094,N_26074,N_28883);
and U31095 (N_31095,N_27502,N_28924);
nand U31096 (N_31096,N_27867,N_28680);
xnor U31097 (N_31097,N_28587,N_25568);
nand U31098 (N_31098,N_28522,N_28208);
or U31099 (N_31099,N_26298,N_25996);
nand U31100 (N_31100,N_26130,N_26385);
and U31101 (N_31101,N_27183,N_27200);
or U31102 (N_31102,N_25699,N_27791);
and U31103 (N_31103,N_26396,N_25331);
xnor U31104 (N_31104,N_25692,N_26638);
xor U31105 (N_31105,N_25161,N_29775);
nand U31106 (N_31106,N_29518,N_26007);
xnor U31107 (N_31107,N_26257,N_28918);
and U31108 (N_31108,N_26435,N_27783);
and U31109 (N_31109,N_29621,N_26818);
or U31110 (N_31110,N_27724,N_26801);
xor U31111 (N_31111,N_29014,N_26070);
or U31112 (N_31112,N_29297,N_29880);
nor U31113 (N_31113,N_25093,N_29258);
xnor U31114 (N_31114,N_29268,N_26434);
nor U31115 (N_31115,N_26888,N_26432);
xor U31116 (N_31116,N_27860,N_25135);
or U31117 (N_31117,N_26220,N_29863);
or U31118 (N_31118,N_27106,N_28259);
nor U31119 (N_31119,N_28200,N_29895);
nand U31120 (N_31120,N_27268,N_26083);
nor U31121 (N_31121,N_29127,N_27723);
and U31122 (N_31122,N_26141,N_25469);
or U31123 (N_31123,N_29013,N_29320);
nand U31124 (N_31124,N_28101,N_29966);
and U31125 (N_31125,N_27358,N_25884);
and U31126 (N_31126,N_25578,N_26728);
and U31127 (N_31127,N_29752,N_27988);
nor U31128 (N_31128,N_29967,N_29333);
nand U31129 (N_31129,N_25200,N_26782);
nand U31130 (N_31130,N_26493,N_26104);
and U31131 (N_31131,N_25345,N_28188);
nor U31132 (N_31132,N_27936,N_25740);
nor U31133 (N_31133,N_26468,N_27032);
nor U31134 (N_31134,N_25875,N_28599);
or U31135 (N_31135,N_27132,N_26805);
nand U31136 (N_31136,N_28174,N_26542);
or U31137 (N_31137,N_26880,N_25352);
and U31138 (N_31138,N_26039,N_28143);
nand U31139 (N_31139,N_26254,N_27850);
xor U31140 (N_31140,N_26918,N_29894);
xor U31141 (N_31141,N_25657,N_25776);
nand U31142 (N_31142,N_29285,N_26627);
nand U31143 (N_31143,N_29572,N_29970);
nor U31144 (N_31144,N_25563,N_28819);
or U31145 (N_31145,N_26037,N_26056);
or U31146 (N_31146,N_27191,N_29347);
and U31147 (N_31147,N_25104,N_28111);
xnor U31148 (N_31148,N_26451,N_28884);
nor U31149 (N_31149,N_26131,N_28198);
nor U31150 (N_31150,N_28394,N_27332);
nand U31151 (N_31151,N_25851,N_25899);
xor U31152 (N_31152,N_26332,N_26714);
and U31153 (N_31153,N_27408,N_26060);
or U31154 (N_31154,N_26446,N_29058);
xnor U31155 (N_31155,N_27661,N_26105);
or U31156 (N_31156,N_25933,N_27391);
nor U31157 (N_31157,N_29198,N_29555);
nor U31158 (N_31158,N_27964,N_27787);
xnor U31159 (N_31159,N_27122,N_29867);
or U31160 (N_31160,N_29965,N_28952);
or U31161 (N_31161,N_28262,N_29304);
and U31162 (N_31162,N_28433,N_29547);
nand U31163 (N_31163,N_27280,N_29593);
or U31164 (N_31164,N_29460,N_26929);
nor U31165 (N_31165,N_25904,N_28574);
or U31166 (N_31166,N_29629,N_27049);
nand U31167 (N_31167,N_25007,N_29696);
nor U31168 (N_31168,N_25608,N_29243);
or U31169 (N_31169,N_29751,N_26749);
or U31170 (N_31170,N_28690,N_29881);
xor U31171 (N_31171,N_26594,N_26569);
and U31172 (N_31172,N_28289,N_27232);
nand U31173 (N_31173,N_29793,N_25605);
or U31174 (N_31174,N_25881,N_27398);
nand U31175 (N_31175,N_27429,N_26837);
nand U31176 (N_31176,N_26971,N_27675);
nand U31177 (N_31177,N_28752,N_27745);
or U31178 (N_31178,N_27523,N_25465);
nand U31179 (N_31179,N_26650,N_28533);
xnor U31180 (N_31180,N_27349,N_29662);
xnor U31181 (N_31181,N_29885,N_25346);
xor U31182 (N_31182,N_25876,N_27973);
nand U31183 (N_31183,N_28922,N_29585);
xnor U31184 (N_31184,N_28358,N_26665);
nor U31185 (N_31185,N_26036,N_26484);
and U31186 (N_31186,N_29713,N_28619);
xnor U31187 (N_31187,N_28936,N_29223);
nor U31188 (N_31188,N_29489,N_26234);
nor U31189 (N_31189,N_26414,N_25103);
xnor U31190 (N_31190,N_29118,N_25298);
nand U31191 (N_31191,N_25456,N_26506);
nand U31192 (N_31192,N_25507,N_28159);
nor U31193 (N_31193,N_29910,N_26905);
or U31194 (N_31194,N_26483,N_29627);
nand U31195 (N_31195,N_26142,N_25097);
nand U31196 (N_31196,N_25336,N_29504);
and U31197 (N_31197,N_25114,N_26869);
or U31198 (N_31198,N_29280,N_26049);
nand U31199 (N_31199,N_25467,N_27161);
nor U31200 (N_31200,N_27605,N_28184);
xnor U31201 (N_31201,N_26538,N_25934);
xnor U31202 (N_31202,N_28089,N_26926);
and U31203 (N_31203,N_27782,N_28993);
xor U31204 (N_31204,N_28147,N_29767);
nor U31205 (N_31205,N_28273,N_25076);
nand U31206 (N_31206,N_25354,N_29352);
xor U31207 (N_31207,N_27418,N_26747);
or U31208 (N_31208,N_25603,N_29337);
xnor U31209 (N_31209,N_25338,N_25723);
or U31210 (N_31210,N_29087,N_27442);
nand U31211 (N_31211,N_26676,N_28652);
or U31212 (N_31212,N_25286,N_26726);
nand U31213 (N_31213,N_29204,N_27581);
xor U31214 (N_31214,N_26986,N_25039);
xor U31215 (N_31215,N_28353,N_29842);
xor U31216 (N_31216,N_26601,N_26346);
nor U31217 (N_31217,N_26871,N_27290);
and U31218 (N_31218,N_25123,N_29711);
and U31219 (N_31219,N_26941,N_26052);
nand U31220 (N_31220,N_29546,N_25677);
nand U31221 (N_31221,N_26184,N_29759);
and U31222 (N_31222,N_26509,N_25189);
or U31223 (N_31223,N_28040,N_26907);
xnor U31224 (N_31224,N_29990,N_25096);
xor U31225 (N_31225,N_27876,N_29114);
nor U31226 (N_31226,N_25994,N_25854);
and U31227 (N_31227,N_29432,N_29511);
or U31228 (N_31228,N_26126,N_28972);
nand U31229 (N_31229,N_29688,N_26983);
and U31230 (N_31230,N_28379,N_25818);
or U31231 (N_31231,N_28223,N_25206);
and U31232 (N_31232,N_29303,N_25241);
nor U31233 (N_31233,N_29609,N_25061);
or U31234 (N_31234,N_27335,N_29669);
nand U31235 (N_31235,N_29237,N_28776);
and U31236 (N_31236,N_25711,N_26241);
nor U31237 (N_31237,N_25301,N_28227);
xnor U31238 (N_31238,N_29379,N_27489);
nor U31239 (N_31239,N_25803,N_27315);
or U31240 (N_31240,N_27767,N_26917);
and U31241 (N_31241,N_28801,N_25733);
nand U31242 (N_31242,N_25712,N_28007);
nand U31243 (N_31243,N_29284,N_27093);
xnor U31244 (N_31244,N_25184,N_28110);
xnor U31245 (N_31245,N_27529,N_27663);
and U31246 (N_31246,N_26136,N_29301);
nand U31247 (N_31247,N_28635,N_27594);
and U31248 (N_31248,N_28061,N_29358);
nor U31249 (N_31249,N_25909,N_29207);
nand U31250 (N_31250,N_28446,N_25289);
and U31251 (N_31251,N_28657,N_26363);
nand U31252 (N_31252,N_27901,N_26322);
nand U31253 (N_31253,N_29980,N_25196);
or U31254 (N_31254,N_25633,N_29386);
and U31255 (N_31255,N_25903,N_26889);
nor U31256 (N_31256,N_27819,N_27042);
nor U31257 (N_31257,N_29134,N_26612);
xor U31258 (N_31258,N_26613,N_28992);
nor U31259 (N_31259,N_25036,N_28953);
and U31260 (N_31260,N_29635,N_25457);
and U31261 (N_31261,N_27667,N_26054);
nor U31262 (N_31262,N_29810,N_26864);
nand U31263 (N_31263,N_27505,N_29564);
or U31264 (N_31264,N_27987,N_27543);
nand U31265 (N_31265,N_28291,N_26112);
or U31266 (N_31266,N_26592,N_28579);
and U31267 (N_31267,N_25205,N_28889);
nand U31268 (N_31268,N_27083,N_29508);
nor U31269 (N_31269,N_27164,N_29576);
or U31270 (N_31270,N_26795,N_29809);
or U31271 (N_31271,N_25528,N_25800);
or U31272 (N_31272,N_27473,N_29730);
xor U31273 (N_31273,N_26213,N_25446);
or U31274 (N_31274,N_28806,N_26903);
nor U31275 (N_31275,N_26418,N_27230);
and U31276 (N_31276,N_26107,N_26827);
xor U31277 (N_31277,N_27859,N_27588);
and U31278 (N_31278,N_26274,N_28490);
and U31279 (N_31279,N_27403,N_27592);
and U31280 (N_31280,N_27807,N_28945);
or U31281 (N_31281,N_25158,N_27412);
xor U31282 (N_31282,N_28672,N_28403);
nor U31283 (N_31283,N_26358,N_29815);
nand U31284 (N_31284,N_26167,N_27742);
nor U31285 (N_31285,N_29594,N_29819);
nor U31286 (N_31286,N_25525,N_25951);
xor U31287 (N_31287,N_26439,N_25153);
xnor U31288 (N_31288,N_28352,N_29031);
or U31289 (N_31289,N_29069,N_25659);
nand U31290 (N_31290,N_28012,N_27167);
nand U31291 (N_31291,N_25549,N_27257);
or U31292 (N_31292,N_28959,N_25863);
or U31293 (N_31293,N_25953,N_25488);
nor U31294 (N_31294,N_28269,N_29315);
nand U31295 (N_31295,N_27974,N_25533);
nand U31296 (N_31296,N_26279,N_27248);
and U31297 (N_31297,N_27199,N_29924);
xnor U31298 (N_31298,N_28660,N_27344);
xnor U31299 (N_31299,N_26355,N_25520);
xor U31300 (N_31300,N_28852,N_27447);
and U31301 (N_31301,N_29046,N_29921);
and U31302 (N_31302,N_26404,N_26928);
and U31303 (N_31303,N_28365,N_26546);
xor U31304 (N_31304,N_27482,N_25856);
nand U31305 (N_31305,N_28359,N_27897);
and U31306 (N_31306,N_29040,N_29750);
nor U31307 (N_31307,N_29766,N_27550);
and U31308 (N_31308,N_28095,N_29556);
nand U31309 (N_31309,N_29042,N_27730);
or U31310 (N_31310,N_29925,N_25988);
xnor U31311 (N_31311,N_27501,N_29675);
nand U31312 (N_31312,N_25628,N_29962);
nand U31313 (N_31313,N_29106,N_27380);
xnor U31314 (N_31314,N_26716,N_26118);
nand U31315 (N_31315,N_25435,N_27674);
xor U31316 (N_31316,N_26017,N_27949);
nand U31317 (N_31317,N_28809,N_25374);
xnor U31318 (N_31318,N_28602,N_28485);
nor U31319 (N_31319,N_25364,N_26035);
nor U31320 (N_31320,N_29381,N_25976);
or U31321 (N_31321,N_29725,N_26299);
nor U31322 (N_31322,N_28305,N_28569);
xnor U31323 (N_31323,N_29608,N_25193);
and U31324 (N_31324,N_27231,N_26736);
or U31325 (N_31325,N_26814,N_25667);
xor U31326 (N_31326,N_26994,N_25042);
and U31327 (N_31327,N_28876,N_25280);
and U31328 (N_31328,N_25387,N_28966);
nor U31329 (N_31329,N_29050,N_28997);
or U31330 (N_31330,N_27009,N_25705);
nand U31331 (N_31331,N_29117,N_29466);
and U31332 (N_31332,N_28704,N_26309);
nor U31333 (N_31333,N_25420,N_28544);
or U31334 (N_31334,N_28709,N_26469);
nand U31335 (N_31335,N_27087,N_28070);
or U31336 (N_31336,N_26006,N_28157);
nand U31337 (N_31337,N_25010,N_26680);
xor U31338 (N_31338,N_28793,N_28722);
xor U31339 (N_31339,N_27552,N_28391);
nand U31340 (N_31340,N_27753,N_27239);
xnor U31341 (N_31341,N_26796,N_27938);
nor U31342 (N_31342,N_28600,N_29481);
and U31343 (N_31343,N_26128,N_25898);
and U31344 (N_31344,N_28835,N_29989);
or U31345 (N_31345,N_29074,N_28033);
or U31346 (N_31346,N_26515,N_25965);
or U31347 (N_31347,N_27074,N_25916);
nor U31348 (N_31348,N_29736,N_26078);
nor U31349 (N_31349,N_26381,N_26866);
xnor U31350 (N_31350,N_25707,N_27426);
xor U31351 (N_31351,N_26868,N_25919);
and U31352 (N_31352,N_29448,N_26139);
nor U31353 (N_31353,N_28349,N_27764);
nand U31354 (N_31354,N_28139,N_26582);
xor U31355 (N_31355,N_25366,N_27305);
and U31356 (N_31356,N_29032,N_28481);
and U31357 (N_31357,N_25168,N_26295);
and U31358 (N_31358,N_25129,N_27069);
nor U31359 (N_31359,N_25479,N_29476);
xor U31360 (N_31360,N_26622,N_28209);
nor U31361 (N_31361,N_25257,N_26406);
nor U31362 (N_31362,N_29276,N_25737);
xnor U31363 (N_31363,N_29059,N_28471);
or U31364 (N_31364,N_29552,N_26119);
nor U31365 (N_31365,N_28180,N_26409);
or U31366 (N_31366,N_27092,N_26013);
or U31367 (N_31367,N_27371,N_29007);
and U31368 (N_31368,N_27556,N_29130);
nor U31369 (N_31369,N_26014,N_28594);
nor U31370 (N_31370,N_28854,N_26724);
nor U31371 (N_31371,N_27520,N_27677);
xor U31372 (N_31372,N_27721,N_25470);
nor U31373 (N_31373,N_27198,N_26080);
nor U31374 (N_31374,N_28760,N_26148);
nor U31375 (N_31375,N_26397,N_29317);
nor U31376 (N_31376,N_27478,N_25209);
xor U31377 (N_31377,N_25830,N_25973);
nand U31378 (N_31378,N_27604,N_28127);
nand U31379 (N_31379,N_28173,N_28887);
nor U31380 (N_31380,N_29452,N_27085);
and U31381 (N_31381,N_26064,N_25046);
nor U31382 (N_31382,N_28669,N_27681);
or U31383 (N_31383,N_28253,N_29768);
nor U31384 (N_31384,N_27467,N_28705);
nor U31385 (N_31385,N_28745,N_25417);
or U31386 (N_31386,N_25474,N_29197);
or U31387 (N_31387,N_29043,N_26174);
or U31388 (N_31388,N_28607,N_29462);
xnor U31389 (N_31389,N_29879,N_28332);
nor U31390 (N_31390,N_29543,N_26443);
and U31391 (N_31391,N_27416,N_29657);
and U31392 (N_31392,N_27749,N_28725);
or U31393 (N_31393,N_25409,N_27307);
and U31394 (N_31394,N_25174,N_26341);
nor U31395 (N_31395,N_28302,N_26456);
nor U31396 (N_31396,N_26424,N_27035);
xnor U31397 (N_31397,N_25609,N_27645);
nor U31398 (N_31398,N_28811,N_29781);
xor U31399 (N_31399,N_29746,N_25824);
nor U31400 (N_31400,N_27223,N_29614);
nor U31401 (N_31401,N_26845,N_26162);
nor U31402 (N_31402,N_29480,N_29173);
nor U31403 (N_31403,N_26562,N_26233);
and U31404 (N_31404,N_25516,N_28726);
and U31405 (N_31405,N_29334,N_29909);
nand U31406 (N_31406,N_29835,N_28502);
or U31407 (N_31407,N_28582,N_29732);
nor U31408 (N_31408,N_29871,N_29145);
and U31409 (N_31409,N_26160,N_25655);
and U31410 (N_31410,N_29503,N_27364);
nor U31411 (N_31411,N_26872,N_28131);
nand U31412 (N_31412,N_28375,N_28154);
nor U31413 (N_31413,N_28256,N_25833);
nand U31414 (N_31414,N_25798,N_28681);
or U31415 (N_31415,N_29738,N_27023);
nand U31416 (N_31416,N_29792,N_27004);
xor U31417 (N_31417,N_29533,N_27099);
and U31418 (N_31418,N_29525,N_28723);
nand U31419 (N_31419,N_25413,N_26374);
or U31420 (N_31420,N_25842,N_27111);
xnor U31421 (N_31421,N_25807,N_27800);
and U31422 (N_31422,N_29322,N_27334);
nor U31423 (N_31423,N_27293,N_26125);
nand U31424 (N_31424,N_28447,N_27614);
nor U31425 (N_31425,N_29394,N_28937);
nor U31426 (N_31426,N_25982,N_29745);
or U31427 (N_31427,N_25358,N_27120);
nor U31428 (N_31428,N_28565,N_25124);
and U31429 (N_31429,N_25125,N_28192);
and U31430 (N_31430,N_26858,N_27243);
or U31431 (N_31431,N_28750,N_28247);
xor U31432 (N_31432,N_27727,N_28775);
nand U31433 (N_31433,N_28168,N_26472);
nor U31434 (N_31434,N_27208,N_25508);
nor U31435 (N_31435,N_29429,N_27671);
nand U31436 (N_31436,N_25611,N_28345);
xnor U31437 (N_31437,N_27803,N_27891);
xnor U31438 (N_31438,N_29010,N_26229);
nand U31439 (N_31439,N_29984,N_28453);
nor U31440 (N_31440,N_26428,N_29410);
nor U31441 (N_31441,N_29791,N_29325);
nand U31442 (N_31442,N_28983,N_28235);
or U31443 (N_31443,N_28293,N_29886);
and U31444 (N_31444,N_29139,N_29156);
xnor U31445 (N_31445,N_25178,N_26743);
and U31446 (N_31446,N_26744,N_25389);
nand U31447 (N_31447,N_25790,N_25081);
xor U31448 (N_31448,N_28950,N_28215);
xor U31449 (N_31449,N_28237,N_27786);
nor U31450 (N_31450,N_28432,N_29519);
and U31451 (N_31451,N_28861,N_29082);
nor U31452 (N_31452,N_25886,N_28795);
or U31453 (N_31453,N_25845,N_28044);
or U31454 (N_31454,N_25079,N_28536);
xor U31455 (N_31455,N_27790,N_25444);
nand U31456 (N_31456,N_28871,N_27527);
nand U31457 (N_31457,N_27274,N_29302);
nor U31458 (N_31458,N_27061,N_26214);
and U31459 (N_31459,N_29840,N_25546);
or U31460 (N_31460,N_29948,N_25538);
and U31461 (N_31461,N_28263,N_28980);
or U31462 (N_31462,N_28153,N_25931);
xnor U31463 (N_31463,N_28942,N_26479);
or U31464 (N_31464,N_29362,N_25560);
and U31465 (N_31465,N_28474,N_28802);
and U31466 (N_31466,N_25433,N_27359);
and U31467 (N_31467,N_28845,N_27439);
nor U31468 (N_31468,N_26075,N_26478);
or U31469 (N_31469,N_27844,N_28315);
nor U31470 (N_31470,N_26115,N_26344);
or U31471 (N_31471,N_28842,N_29579);
and U31472 (N_31472,N_29388,N_28978);
xnor U31473 (N_31473,N_29328,N_26536);
xor U31474 (N_31474,N_25025,N_26205);
nor U31475 (N_31475,N_25482,N_27743);
nand U31476 (N_31476,N_27285,N_29438);
and U31477 (N_31477,N_28695,N_25540);
xnor U31478 (N_31478,N_27435,N_29153);
and U31479 (N_31479,N_28062,N_27038);
or U31480 (N_31480,N_25021,N_27021);
or U31481 (N_31481,N_29697,N_26777);
or U31482 (N_31482,N_25543,N_26883);
nand U31483 (N_31483,N_29101,N_28511);
xor U31484 (N_31484,N_29033,N_26765);
nor U31485 (N_31485,N_26247,N_26844);
and U31486 (N_31486,N_29319,N_27578);
xnor U31487 (N_31487,N_27603,N_28389);
and U31488 (N_31488,N_25472,N_29723);
or U31489 (N_31489,N_26519,N_29646);
nand U31490 (N_31490,N_29655,N_29764);
nor U31491 (N_31491,N_29874,N_29743);
or U31492 (N_31492,N_28730,N_25120);
or U31493 (N_31493,N_27494,N_27098);
or U31494 (N_31494,N_26862,N_27174);
xnor U31495 (N_31495,N_29488,N_28714);
and U31496 (N_31496,N_29527,N_27034);
nand U31497 (N_31497,N_27480,N_25506);
nor U31498 (N_31498,N_27853,N_29598);
xnor U31499 (N_31499,N_28268,N_26059);
and U31500 (N_31500,N_27490,N_26906);
and U31501 (N_31501,N_29019,N_26545);
nand U31502 (N_31502,N_29296,N_28284);
nand U31503 (N_31503,N_28400,N_29960);
or U31504 (N_31504,N_27492,N_26461);
xnor U31505 (N_31505,N_27845,N_27990);
nor U31506 (N_31506,N_27378,N_27966);
or U31507 (N_31507,N_27159,N_27209);
and U31508 (N_31508,N_28220,N_26251);
nand U31509 (N_31509,N_29628,N_29239);
or U31510 (N_31510,N_26311,N_29306);
nand U31511 (N_31511,N_29219,N_28455);
nor U31512 (N_31512,N_26058,N_27555);
nand U31513 (N_31513,N_26053,N_29703);
or U31514 (N_31514,N_25575,N_28117);
xnor U31515 (N_31515,N_29761,N_25729);
or U31516 (N_31516,N_26447,N_27933);
nor U31517 (N_31517,N_25745,N_25110);
nand U31518 (N_31518,N_28515,N_25000);
nor U31519 (N_31519,N_27357,N_26199);
nand U31520 (N_31520,N_28306,N_26649);
nand U31521 (N_31521,N_28319,N_25701);
nor U31522 (N_31522,N_25650,N_27156);
xnor U31523 (N_31523,N_25142,N_26846);
nor U31524 (N_31524,N_29992,N_29187);
and U31525 (N_31525,N_26766,N_29626);
nor U31526 (N_31526,N_28079,N_29414);
nor U31527 (N_31527,N_29136,N_29331);
nand U31528 (N_31528,N_28368,N_27713);
xor U31529 (N_31529,N_25972,N_27993);
xnor U31530 (N_31530,N_25229,N_25115);
nor U31531 (N_31531,N_26491,N_25939);
nor U31532 (N_31532,N_28592,N_29820);
and U31533 (N_31533,N_29092,N_27524);
nand U31534 (N_31534,N_28054,N_28642);
nor U31535 (N_31535,N_27586,N_25080);
xnor U31536 (N_31536,N_25143,N_29479);
xor U31537 (N_31537,N_28702,N_29478);
xnor U31538 (N_31538,N_26629,N_27368);
xnor U31539 (N_31539,N_28653,N_29664);
nand U31540 (N_31540,N_25360,N_28948);
nand U31541 (N_31541,N_26324,N_29161);
or U31542 (N_31542,N_28608,N_26659);
nand U31543 (N_31543,N_25590,N_29643);
and U31544 (N_31544,N_29392,N_26267);
nor U31545 (N_31545,N_27568,N_25480);
nand U31546 (N_31546,N_25618,N_26275);
or U31547 (N_31547,N_26937,N_26494);
nand U31548 (N_31548,N_27005,N_29006);
xor U31549 (N_31549,N_28949,N_29887);
and U31550 (N_31550,N_28271,N_26305);
xor U31551 (N_31551,N_26121,N_26009);
xnor U31552 (N_31552,N_25486,N_25273);
or U31553 (N_31553,N_27287,N_29876);
or U31554 (N_31554,N_29371,N_29510);
and U31555 (N_31555,N_28784,N_29801);
or U31556 (N_31556,N_28716,N_29469);
nand U31557 (N_31557,N_27994,N_27781);
and U31558 (N_31558,N_29423,N_28267);
and U31559 (N_31559,N_25498,N_27840);
nor U31560 (N_31560,N_26259,N_28783);
or U31561 (N_31561,N_25592,N_26024);
or U31562 (N_31562,N_27108,N_27497);
xor U31563 (N_31563,N_26644,N_29782);
or U31564 (N_31564,N_26658,N_29699);
xnor U31565 (N_31565,N_25685,N_28957);
or U31566 (N_31566,N_25299,N_28965);
nor U31567 (N_31567,N_27996,N_25228);
nor U31568 (N_31568,N_26822,N_26353);
nand U31569 (N_31569,N_27697,N_28098);
xnor U31570 (N_31570,N_28250,N_28083);
nor U31571 (N_31571,N_29985,N_26230);
or U31572 (N_31572,N_28646,N_27809);
nor U31573 (N_31573,N_25407,N_28431);
nand U31574 (N_31574,N_25092,N_27871);
nand U31575 (N_31575,N_27266,N_26510);
nor U31576 (N_31576,N_28630,N_29603);
xnor U31577 (N_31577,N_27125,N_26699);
or U31578 (N_31578,N_29133,N_29903);
or U31579 (N_31579,N_25369,N_25652);
xnor U31580 (N_31580,N_29744,N_26179);
nand U31581 (N_31581,N_28614,N_26093);
and U31582 (N_31582,N_27168,N_27445);
xnor U31583 (N_31583,N_29722,N_28387);
and U31584 (N_31584,N_26835,N_28279);
and U31585 (N_31585,N_25738,N_29403);
xnor U31586 (N_31586,N_27582,N_29735);
nand U31587 (N_31587,N_25016,N_27333);
xor U31588 (N_31588,N_28517,N_29911);
nor U31589 (N_31589,N_26110,N_28764);
nor U31590 (N_31590,N_29376,N_28048);
and U31591 (N_31591,N_28071,N_28216);
nor U31592 (N_31592,N_25477,N_27865);
xor U31593 (N_31593,N_28701,N_25304);
or U31594 (N_31594,N_25088,N_29707);
nand U31595 (N_31595,N_29072,N_29368);
or U31596 (N_31596,N_26099,N_29039);
nand U31597 (N_31597,N_26376,N_28578);
nand U31598 (N_31598,N_27814,N_28611);
nand U31599 (N_31599,N_26421,N_29174);
nor U31600 (N_31600,N_27830,N_25156);
nand U31601 (N_31601,N_28261,N_29926);
and U31602 (N_31602,N_29464,N_29826);
xnor U31603 (N_31603,N_26756,N_27838);
xor U31604 (N_31604,N_25964,N_29436);
xor U31605 (N_31605,N_27916,N_25644);
nand U31606 (N_31606,N_26345,N_27817);
and U31607 (N_31607,N_29678,N_25573);
nand U31608 (N_31608,N_28109,N_26849);
xnor U31609 (N_31609,N_27908,N_26982);
and U31610 (N_31610,N_26779,N_26689);
xnor U31611 (N_31611,N_26786,N_26431);
nor U31612 (N_31612,N_26799,N_26821);
and U31613 (N_31613,N_29599,N_27324);
or U31614 (N_31614,N_25666,N_26289);
nand U31615 (N_31615,N_27975,N_28047);
nand U31616 (N_31616,N_25049,N_29855);
and U31617 (N_31617,N_25240,N_25847);
nor U31618 (N_31618,N_28919,N_27097);
nand U31619 (N_31619,N_28057,N_26100);
and U31620 (N_31620,N_29200,N_28991);
nand U31621 (N_31621,N_27771,N_26221);
xor U31622 (N_31622,N_26904,N_28000);
and U31623 (N_31623,N_26169,N_26185);
nand U31624 (N_31624,N_25742,N_27899);
or U31625 (N_31625,N_25058,N_28395);
xor U31626 (N_31626,N_28498,N_25362);
nand U31627 (N_31627,N_25099,N_25793);
and U31628 (N_31628,N_25302,N_25373);
xnor U31629 (N_31629,N_28028,N_28115);
or U31630 (N_31630,N_25752,N_26001);
nor U31631 (N_31631,N_28066,N_29680);
nor U31632 (N_31632,N_28294,N_25601);
nor U31633 (N_31633,N_25197,N_26992);
or U31634 (N_31634,N_27644,N_27797);
nand U31635 (N_31635,N_26794,N_27394);
and U31636 (N_31636,N_28605,N_27186);
nor U31637 (N_31637,N_29687,N_26086);
nand U31638 (N_31638,N_29780,N_28513);
xor U31639 (N_31639,N_25054,N_26237);
nand U31640 (N_31640,N_26605,N_29656);
and U31641 (N_31641,N_28458,N_28344);
xnor U31642 (N_31642,N_25826,N_29453);
xor U31643 (N_31643,N_27227,N_28428);
and U31644 (N_31644,N_26617,N_25116);
nand U31645 (N_31645,N_25791,N_26614);
nor U31646 (N_31646,N_26529,N_25888);
xor U31647 (N_31647,N_28610,N_28059);
or U31648 (N_31648,N_26621,N_25082);
nor U31649 (N_31649,N_25913,N_28186);
and U31650 (N_31650,N_29067,N_25466);
and U31651 (N_31651,N_25144,N_27103);
nand U31652 (N_31652,N_26626,N_25332);
xnor U31653 (N_31653,N_26548,N_28381);
or U31654 (N_31654,N_29833,N_28019);
and U31655 (N_31655,N_27054,N_27925);
or U31656 (N_31656,N_28773,N_28994);
nand U31657 (N_31657,N_28864,N_25620);
and U31658 (N_31658,N_25086,N_25468);
or U31659 (N_31659,N_25725,N_29159);
nor U31660 (N_31660,N_26195,N_27181);
nand U31661 (N_31661,N_28870,N_25857);
nor U31662 (N_31662,N_26329,N_29641);
and U31663 (N_31663,N_26069,N_27948);
nor U31664 (N_31664,N_29125,N_25221);
nor U31665 (N_31665,N_27856,N_25631);
nand U31666 (N_31666,N_29076,N_27063);
or U31667 (N_31667,N_27532,N_27116);
nor U31668 (N_31668,N_27084,N_27839);
and U31669 (N_31669,N_29135,N_25944);
nor U31670 (N_31670,N_25316,N_26958);
and U31671 (N_31671,N_26264,N_25766);
or U31672 (N_31672,N_26252,N_28868);
xnor U31673 (N_31673,N_28581,N_28171);
nor U31674 (N_31674,N_25450,N_27062);
and U31675 (N_31675,N_28356,N_25139);
or U31676 (N_31676,N_28700,N_26002);
and U31677 (N_31677,N_27772,N_28244);
nor U31678 (N_31678,N_29412,N_27760);
nor U31679 (N_31679,N_29220,N_27573);
xor U31680 (N_31680,N_25217,N_25233);
nand U31681 (N_31681,N_29786,N_25606);
nand U31682 (N_31682,N_28914,N_26370);
xnor U31683 (N_31683,N_29513,N_28756);
nand U31684 (N_31684,N_25175,N_29021);
and U31685 (N_31685,N_27880,N_27320);
nor U31686 (N_31686,N_28010,N_25066);
nand U31687 (N_31687,N_29176,N_26280);
xor U31688 (N_31688,N_27221,N_29494);
xor U31689 (N_31689,N_28551,N_27128);
nor U31690 (N_31690,N_26379,N_27596);
nor U31691 (N_31691,N_28229,N_28468);
and U31692 (N_31692,N_26824,N_29583);
nand U31693 (N_31693,N_29138,N_25242);
or U31694 (N_31694,N_27672,N_26088);
and U31695 (N_31695,N_27968,N_28254);
nor U31696 (N_31696,N_25720,N_28814);
and U31697 (N_31697,N_28411,N_26619);
and U31698 (N_31698,N_27735,N_27741);
nand U31699 (N_31699,N_29343,N_27013);
xnor U31700 (N_31700,N_26696,N_25937);
xor U31701 (N_31701,N_29796,N_28441);
or U31702 (N_31702,N_26102,N_26204);
xnor U31703 (N_31703,N_28843,N_28618);
nand U31704 (N_31704,N_25150,N_28489);
nor U31705 (N_31705,N_29203,N_25693);
nand U31706 (N_31706,N_29587,N_28546);
xor U31707 (N_31707,N_26764,N_26290);
nor U31708 (N_31708,N_28287,N_25037);
nand U31709 (N_31709,N_27785,N_26683);
xnor U31710 (N_31710,N_26025,N_28847);
xnor U31711 (N_31711,N_27946,N_29254);
and U31712 (N_31712,N_29224,N_27685);
and U31713 (N_31713,N_29269,N_28651);
xnor U31714 (N_31714,N_29259,N_29501);
xor U31715 (N_31715,N_29202,N_27612);
nor U31716 (N_31716,N_27754,N_25521);
or U31717 (N_31717,N_29864,N_27118);
and U31718 (N_31718,N_29286,N_28796);
nor U31719 (N_31719,N_26212,N_28736);
nand U31720 (N_31720,N_28480,N_25588);
xnor U31721 (N_31721,N_28304,N_29702);
xnor U31722 (N_31722,N_29389,N_28246);
xnor U31723 (N_31723,N_29279,N_29437);
and U31724 (N_31724,N_26449,N_27113);
nand U31725 (N_31725,N_27688,N_27386);
nand U31726 (N_31726,N_29212,N_25716);
or U31727 (N_31727,N_26113,N_28735);
and U31728 (N_31728,N_25263,N_28207);
or U31729 (N_31729,N_26996,N_26228);
or U31730 (N_31730,N_26651,N_28213);
or U31731 (N_31731,N_28496,N_29589);
or U31732 (N_31732,N_26921,N_26620);
xnor U31733 (N_31733,N_26933,N_25671);
or U31734 (N_31734,N_27986,N_27566);
or U31735 (N_31735,N_25122,N_26082);
or U31736 (N_31736,N_25019,N_28475);
nand U31737 (N_31737,N_27474,N_29993);
nor U31738 (N_31738,N_27050,N_29875);
nor U31739 (N_31739,N_26631,N_27820);
or U31740 (N_31740,N_29578,N_27757);
or U31741 (N_31741,N_27138,N_27381);
xnor U31742 (N_31742,N_27774,N_27115);
or U31743 (N_31743,N_25321,N_27251);
xnor U31744 (N_31744,N_26224,N_26609);
and U31745 (N_31745,N_29405,N_25998);
or U31746 (N_31746,N_29137,N_27890);
and U31747 (N_31747,N_25269,N_25669);
nor U31748 (N_31748,N_27752,N_25754);
and U31749 (N_31749,N_25935,N_29559);
or U31750 (N_31750,N_26673,N_29257);
or U31751 (N_31751,N_26642,N_29777);
and U31752 (N_31752,N_27419,N_27455);
and U31753 (N_31753,N_26962,N_29004);
or U31754 (N_31754,N_26899,N_27633);
nand U31755 (N_31755,N_26095,N_27406);
nand U31756 (N_31756,N_25542,N_25377);
nand U31757 (N_31757,N_28780,N_25313);
nor U31758 (N_31758,N_26454,N_28743);
xor U31759 (N_31759,N_26708,N_29521);
nand U31760 (N_31760,N_29169,N_27088);
or U31761 (N_31761,N_25961,N_28374);
or U31762 (N_31762,N_29211,N_27545);
nand U31763 (N_31763,N_25894,N_26473);
nor U31764 (N_31764,N_28088,N_25952);
and U31765 (N_31765,N_25959,N_26047);
and U31766 (N_31766,N_25732,N_26390);
nand U31767 (N_31767,N_28613,N_28084);
xor U31768 (N_31768,N_28689,N_27600);
or U31769 (N_31769,N_26170,N_25447);
or U31770 (N_31770,N_25009,N_26526);
xor U31771 (N_31771,N_27047,N_27811);
or U31772 (N_31772,N_29531,N_25784);
xor U31773 (N_31773,N_27217,N_26674);
nand U31774 (N_31774,N_27311,N_28542);
xnor U31775 (N_31775,N_25750,N_25410);
nor U31776 (N_31776,N_25106,N_27660);
and U31777 (N_31777,N_25526,N_27549);
or U31778 (N_31778,N_25454,N_29246);
nand U31779 (N_31779,N_25985,N_26807);
nand U31780 (N_31780,N_29986,N_27270);
and U31781 (N_31781,N_27947,N_26193);
or U31782 (N_31782,N_27643,N_27941);
nand U31783 (N_31783,N_25216,N_25956);
and U31784 (N_31784,N_29015,N_26091);
nor U31785 (N_31785,N_26445,N_26735);
nor U31786 (N_31786,N_25529,N_29877);
and U31787 (N_31787,N_25291,N_29661);
and U31788 (N_31788,N_29762,N_27531);
xnor U31789 (N_31789,N_29443,N_27048);
or U31790 (N_31790,N_29573,N_29249);
and U31791 (N_31791,N_26134,N_28123);
and U31792 (N_31792,N_25773,N_25418);
and U31793 (N_31793,N_26042,N_26767);
xor U31794 (N_31794,N_25284,N_26960);
and U31795 (N_31795,N_26618,N_28325);
xor U31796 (N_31796,N_25688,N_26101);
nor U31797 (N_31797,N_27033,N_28206);
nand U31798 (N_31798,N_29831,N_26788);
xnor U31799 (N_31799,N_29856,N_28724);
or U31800 (N_31800,N_28274,N_27449);
and U31801 (N_31801,N_27551,N_29209);
nor U31802 (N_31802,N_25089,N_28189);
xor U31803 (N_31803,N_25571,N_26168);
nor U31804 (N_31804,N_25442,N_28633);
nand U31805 (N_31805,N_29677,N_27707);
xnor U31806 (N_31806,N_27210,N_25635);
nor U31807 (N_31807,N_25014,N_28509);
nor U31808 (N_31808,N_28464,N_25335);
or U31809 (N_31809,N_29839,N_28329);
nand U31810 (N_31810,N_25551,N_29647);
xnor U31811 (N_31811,N_26686,N_25084);
nand U31812 (N_31812,N_25874,N_25458);
nand U31813 (N_31813,N_26278,N_26741);
nand U31814 (N_31814,N_27737,N_25515);
xor U31815 (N_31815,N_27616,N_28150);
nand U31816 (N_31816,N_25686,N_26183);
and U31817 (N_31817,N_27299,N_28734);
or U31818 (N_31818,N_28272,N_29056);
xnor U31819 (N_31819,N_28524,N_25698);
xnor U31820 (N_31820,N_29370,N_25210);
and U31821 (N_31821,N_27778,N_27872);
xnor U31822 (N_31822,N_27155,N_29800);
xnor U31823 (N_31823,N_28326,N_27352);
or U31824 (N_31824,N_25283,N_29841);
and U31825 (N_31825,N_28548,N_26731);
and U31826 (N_31826,N_28898,N_25598);
xnor U31827 (N_31827,N_26481,N_26873);
nand U31828 (N_31828,N_28436,N_26860);
xor U31829 (N_31829,N_26999,N_29597);
nor U31830 (N_31830,N_26268,N_25697);
and U31831 (N_31831,N_28563,N_27269);
nand U31832 (N_31832,N_29659,N_26861);
or U31833 (N_31833,N_26819,N_25536);
or U31834 (N_31834,N_25993,N_29377);
xnor U31835 (N_31835,N_28042,N_25149);
nor U31836 (N_31836,N_29496,N_26085);
nor U31837 (N_31837,N_27160,N_28934);
nand U31838 (N_31838,N_27039,N_25202);
xor U31839 (N_31839,N_25179,N_28641);
nor U31840 (N_31840,N_25868,N_26948);
nor U31841 (N_31841,N_27329,N_26050);
xor U31842 (N_31842,N_28217,N_28185);
xnor U31843 (N_31843,N_27382,N_28107);
and U31844 (N_31844,N_27417,N_25095);
nor U31845 (N_31845,N_29024,N_25264);
xor U31846 (N_31846,N_28364,N_26163);
xor U31847 (N_31847,N_29958,N_26430);
nand U31848 (N_31848,N_29650,N_26132);
nand U31849 (N_31849,N_26263,N_28138);
nand U31850 (N_31850,N_28452,N_25318);
and U31851 (N_31851,N_26643,N_28288);
xnor U31852 (N_31852,N_29110,N_25419);
and U31853 (N_31853,N_29982,N_25075);
xor U31854 (N_31854,N_27861,N_25353);
and U31855 (N_31855,N_29866,N_26560);
xor U31856 (N_31856,N_27536,N_27703);
or U31857 (N_31857,N_29329,N_27823);
or U31858 (N_31858,N_25339,N_29034);
nand U31859 (N_31859,N_26368,N_27997);
xor U31860 (N_31860,N_27810,N_29450);
xnor U31861 (N_31861,N_27078,N_27634);
xor U31862 (N_31862,N_29868,N_26103);
or U31863 (N_31863,N_27670,N_29491);
xor U31864 (N_31864,N_26790,N_28817);
nor U31865 (N_31865,N_27715,N_25277);
nand U31866 (N_31866,N_25535,N_27869);
xor U31867 (N_31867,N_28469,N_26839);
xnor U31868 (N_31868,N_29205,N_29287);
or U31869 (N_31869,N_26114,N_25694);
and U31870 (N_31870,N_27931,N_27341);
and U31871 (N_31871,N_28970,N_26800);
xor U31872 (N_31872,N_29602,N_26900);
nor U31873 (N_31873,N_26603,N_29882);
xor U31874 (N_31874,N_26201,N_27094);
xor U31875 (N_31875,N_26540,N_27264);
or U31876 (N_31876,N_26150,N_29103);
nand U31877 (N_31877,N_27493,N_27991);
nor U31878 (N_31878,N_28486,N_29691);
nor U31879 (N_31879,N_27770,N_27706);
xnor U31880 (N_31880,N_28228,N_29418);
nand U31881 (N_31881,N_25879,N_28129);
or U31882 (N_31882,N_26785,N_25295);
and U31883 (N_31883,N_29000,N_28516);
and U31884 (N_31884,N_27260,N_29544);
nor U31885 (N_31885,N_25379,N_26828);
or U31886 (N_31886,N_27471,N_25815);
xnor U31887 (N_31887,N_25226,N_28577);
and U31888 (N_31888,N_25243,N_25464);
nor U31889 (N_31889,N_26797,N_28314);
xor U31890 (N_31890,N_25681,N_28093);
or U31891 (N_31891,N_29592,N_29591);
xnor U31892 (N_31892,N_28318,N_26339);
and U31893 (N_31893,N_26366,N_27170);
or U31894 (N_31894,N_25127,N_28031);
nor U31895 (N_31895,N_27053,N_25432);
and U31896 (N_31896,N_28102,N_27567);
xor U31897 (N_31897,N_28661,N_29144);
nor U31898 (N_31898,N_26910,N_26922);
nand U31899 (N_31899,N_25981,N_25195);
or U31900 (N_31900,N_29658,N_29196);
nor U31901 (N_31901,N_25245,N_27095);
and U31902 (N_31902,N_28104,N_29670);
or U31903 (N_31903,N_26930,N_25212);
and U31904 (N_31904,N_28195,N_25185);
and U31905 (N_31905,N_28911,N_26565);
and U31906 (N_31906,N_27196,N_25992);
xnor U31907 (N_31907,N_25794,N_25809);
xor U31908 (N_31908,N_26419,N_27815);
or U31909 (N_31909,N_26177,N_25183);
or U31910 (N_31910,N_29359,N_28518);
xnor U31911 (N_31911,N_28020,N_27464);
nand U31912 (N_31912,N_29939,N_27440);
or U31913 (N_31913,N_25583,N_27145);
or U31914 (N_31914,N_28321,N_27205);
and U31915 (N_31915,N_25673,N_28987);
nor U31916 (N_31916,N_26505,N_29827);
xor U31917 (N_31917,N_26628,N_29845);
and U31918 (N_31918,N_26501,N_29770);
xor U31919 (N_31919,N_29120,N_28554);
or U31920 (N_31920,N_29679,N_27906);
or U31921 (N_31921,N_25885,N_28990);
and U31922 (N_31922,N_28846,N_25923);
or U31923 (N_31923,N_27886,N_28758);
nand U31924 (N_31924,N_29160,N_28424);
nor U31925 (N_31925,N_29905,N_27011);
nand U31926 (N_31926,N_29755,N_27651);
or U31927 (N_31927,N_27407,N_26521);
nor U31928 (N_31928,N_28772,N_27415);
xor U31929 (N_31929,N_28482,N_29912);
nor U31930 (N_31930,N_27835,N_28065);
and U31931 (N_31931,N_25155,N_25702);
nor U31932 (N_31932,N_27599,N_26222);
nand U31933 (N_31933,N_27917,N_26916);
nand U31934 (N_31934,N_29419,N_27370);
nor U31935 (N_31935,N_26165,N_27277);
nor U31936 (N_31936,N_27769,N_28276);
xor U31937 (N_31937,N_26886,N_26530);
nor U31938 (N_31938,N_26087,N_27943);
nand U31939 (N_31939,N_25999,N_25073);
nor U31940 (N_31940,N_29022,N_26574);
nor U31941 (N_31941,N_28540,N_29794);
or U31942 (N_31942,N_26062,N_26187);
nand U31943 (N_31943,N_25090,N_27657);
xnor U31944 (N_31944,N_25121,N_27798);
or U31945 (N_31945,N_29772,N_26692);
nor U31946 (N_31946,N_29682,N_25846);
or U31947 (N_31947,N_28106,N_26954);
nor U31948 (N_31948,N_25640,N_26348);
nand U31949 (N_31949,N_28874,N_27242);
xor U31950 (N_31950,N_29870,N_26317);
nand U31951 (N_31951,N_25890,N_27090);
or U31952 (N_31952,N_27353,N_26117);
nor U31953 (N_31953,N_29094,N_25188);
xnor U31954 (N_31954,N_25194,N_25034);
xnor U31955 (N_31955,N_25604,N_29217);
and U31956 (N_31956,N_26723,N_25372);
and U31957 (N_31957,N_26159,N_26045);
nor U31958 (N_31958,N_27669,N_28347);
nand U31959 (N_31959,N_27739,N_26319);
and U31960 (N_31960,N_29179,N_28114);
xor U31961 (N_31961,N_27638,N_26646);
or U31962 (N_31962,N_26235,N_25661);
or U31963 (N_31963,N_25181,N_29404);
nand U31964 (N_31964,N_25553,N_25960);
or U31965 (N_31965,N_27907,N_25562);
or U31966 (N_31966,N_26648,N_25411);
or U31967 (N_31967,N_27043,N_29613);
nand U31968 (N_31968,N_25102,N_29836);
nand U31969 (N_31969,N_25255,N_26902);
or U31970 (N_31970,N_28593,N_27016);
and U31971 (N_31971,N_27366,N_26442);
nand U31972 (N_31972,N_25887,N_27427);
or U31973 (N_31973,N_25743,N_28205);
nand U31974 (N_31974,N_26961,N_25787);
nor U31975 (N_31975,N_25722,N_27456);
nand U31976 (N_31976,N_26292,N_26244);
and U31977 (N_31977,N_28860,N_26533);
and U31978 (N_31978,N_26834,N_25137);
nor U31979 (N_31979,N_26875,N_29774);
or U31980 (N_31980,N_26876,N_27843);
and U31981 (N_31981,N_27475,N_28461);
nor U31982 (N_31982,N_25186,N_27834);
or U31983 (N_31983,N_29293,N_27411);
nand U31984 (N_31984,N_26632,N_25215);
and U31985 (N_31985,N_25954,N_29695);
and U31986 (N_31986,N_28962,N_28310);
xnor U31987 (N_31987,N_27195,N_28803);
nand U31988 (N_31988,N_28439,N_25739);
or U31989 (N_31989,N_27182,N_29946);
xor U31990 (N_31990,N_29012,N_26420);
or U31991 (N_31991,N_28988,N_27178);
xor U31992 (N_31992,N_27680,N_26556);
and U31993 (N_31993,N_26223,N_27058);
xor U31994 (N_31994,N_28875,N_27848);
xnor U31995 (N_31995,N_28923,N_27750);
or U31996 (N_31996,N_27950,N_26172);
nand U31997 (N_31997,N_29734,N_28810);
and U31998 (N_31998,N_26953,N_28841);
nand U31999 (N_31999,N_28175,N_25067);
or U32000 (N_32000,N_28140,N_27444);
and U32001 (N_32001,N_25820,N_28230);
or U32002 (N_32002,N_25147,N_28068);
nand U32003 (N_32003,N_25627,N_26682);
xor U32004 (N_32004,N_26639,N_28562);
or U32005 (N_32005,N_27081,N_27363);
or U32006 (N_32006,N_28858,N_28612);
nor U32007 (N_32007,N_28856,N_27642);
or U32008 (N_32008,N_26595,N_28941);
and U32009 (N_32009,N_29446,N_28046);
or U32010 (N_32010,N_26459,N_29263);
nand U32011 (N_32011,N_28837,N_25363);
nor U32012 (N_32012,N_27593,N_29524);
nand U32013 (N_32013,N_28398,N_26504);
and U32014 (N_32014,N_27801,N_27295);
xnor U32015 (N_32015,N_25541,N_26853);
nor U32016 (N_32016,N_25782,N_28755);
and U32017 (N_32017,N_29474,N_26349);
nand U32018 (N_32018,N_26410,N_28742);
and U32019 (N_32019,N_25632,N_25788);
and U32020 (N_32020,N_27354,N_29425);
nand U32021 (N_32021,N_29295,N_25713);
nor U32022 (N_32022,N_27082,N_26028);
nand U32023 (N_32023,N_29896,N_25639);
xor U32024 (N_32024,N_29122,N_28155);
nor U32025 (N_32025,N_26701,N_27278);
and U32026 (N_32026,N_27413,N_26678);
and U32027 (N_32027,N_28570,N_27142);
nor U32028 (N_32028,N_28685,N_29104);
and U32029 (N_32029,N_29914,N_25900);
nand U32030 (N_32030,N_26781,N_28976);
or U32031 (N_32031,N_25249,N_28370);
or U32032 (N_32032,N_28504,N_26307);
nor U32033 (N_32033,N_27414,N_25368);
nand U32034 (N_32034,N_29294,N_26516);
xor U32035 (N_32035,N_25759,N_26425);
nor U32036 (N_32036,N_29401,N_25749);
or U32037 (N_32037,N_26995,N_29884);
xor U32038 (N_32038,N_29321,N_27188);
nand U32039 (N_32039,N_28322,N_27377);
xor U32040 (N_32040,N_29799,N_25753);
nor U32041 (N_32041,N_25490,N_27854);
nand U32042 (N_32042,N_29814,N_25207);
and U32043 (N_32043,N_25940,N_28530);
or U32044 (N_32044,N_26407,N_25534);
nor U32045 (N_32045,N_26436,N_27995);
nand U32046 (N_32046,N_29811,N_28712);
nand U32047 (N_32047,N_26507,N_26720);
nand U32048 (N_32048,N_27066,N_28967);
and U32049 (N_32049,N_29645,N_27197);
and U32050 (N_32050,N_28759,N_26825);
or U32051 (N_32051,N_29785,N_26240);
nand U32052 (N_32052,N_25487,N_27190);
nor U32053 (N_32053,N_29853,N_25078);
nor U32054 (N_32054,N_27900,N_25683);
xnor U32055 (N_32055,N_29454,N_26250);
or U32056 (N_32056,N_28499,N_28346);
xor U32057 (N_32057,N_28292,N_28636);
nand U32058 (N_32058,N_26338,N_27057);
nor U32059 (N_32059,N_29399,N_28890);
and U32060 (N_32060,N_29944,N_26633);
and U32061 (N_32061,N_29184,N_26372);
and U32062 (N_32062,N_28616,N_26303);
nand U32063 (N_32063,N_29390,N_28771);
nor U32064 (N_32064,N_28821,N_25100);
nor U32065 (N_32065,N_29201,N_27202);
nand U32066 (N_32066,N_27926,N_26544);
or U32067 (N_32067,N_26655,N_27466);
and U32068 (N_32068,N_25544,N_29528);
and U32069 (N_32069,N_28338,N_27345);
nand U32070 (N_32070,N_27319,N_29858);
or U32071 (N_32071,N_26138,N_28035);
xnor U32072 (N_32072,N_26596,N_25431);
xor U32073 (N_32073,N_27571,N_27139);
xor U32074 (N_32074,N_27548,N_25918);
xor U32075 (N_32075,N_27866,N_27731);
nand U32076 (N_32076,N_29487,N_28103);
and U32077 (N_32077,N_29465,N_27102);
nor U32078 (N_32078,N_28043,N_28404);
xor U32079 (N_32079,N_25958,N_29086);
nand U32080 (N_32080,N_29506,N_29584);
xor U32081 (N_32081,N_25804,N_26811);
nor U32082 (N_32082,N_28120,N_28555);
or U32083 (N_32083,N_28558,N_28476);
and U32084 (N_32084,N_26488,N_29441);
xnor U32085 (N_32085,N_28996,N_26402);
or U32086 (N_32086,N_28507,N_26034);
nor U32087 (N_32087,N_25356,N_28676);
nand U32088 (N_32088,N_25305,N_25741);
and U32089 (N_32089,N_25408,N_27514);
xor U32090 (N_32090,N_27522,N_29545);
nor U32091 (N_32091,N_29272,N_27481);
nand U32092 (N_32092,N_26514,N_28036);
or U32093 (N_32093,N_28401,N_29065);
nor U32094 (N_32094,N_25140,N_26881);
nand U32095 (N_32095,N_25567,N_26874);
xor U32096 (N_32096,N_27699,N_29266);
xor U32097 (N_32097,N_28741,N_26330);
nand U32098 (N_32098,N_28655,N_26429);
xnor U32099 (N_32099,N_25556,N_27714);
xnor U32100 (N_32100,N_26347,N_26225);
or U32101 (N_32101,N_25637,N_29773);
nand U32102 (N_32102,N_26008,N_25569);
and U32103 (N_32103,N_27192,N_29716);
or U32104 (N_32104,N_27450,N_29108);
nand U32105 (N_32105,N_29206,N_29724);
and U32106 (N_32106,N_26265,N_27577);
xor U32107 (N_32107,N_29825,N_26718);
and U32108 (N_32108,N_28740,N_25527);
or U32109 (N_32109,N_29027,N_29500);
or U32110 (N_32110,N_28832,N_25101);
and U32111 (N_32111,N_28201,N_25165);
xnor U32112 (N_32112,N_28030,N_28598);
nand U32113 (N_32113,N_27002,N_26357);
and U32114 (N_32114,N_28023,N_26373);
and U32115 (N_32115,N_25170,N_25013);
or U32116 (N_32116,N_27923,N_27565);
and U32117 (N_32117,N_27459,N_26202);
and U32118 (N_32118,N_26227,N_25574);
xor U32119 (N_32119,N_27591,N_28528);
and U32120 (N_32120,N_27452,N_26711);
nor U32121 (N_32121,N_26934,N_27584);
xnor U32122 (N_32122,N_26851,N_29704);
and U32123 (N_32123,N_27659,N_26816);
nor U32124 (N_32124,N_25581,N_27423);
and U32125 (N_32125,N_28144,N_28226);
xor U32126 (N_32126,N_29672,N_29622);
and U32127 (N_32127,N_26021,N_27303);
and U32128 (N_32128,N_27602,N_27784);
nor U32129 (N_32129,N_26693,N_27206);
xnor U32130 (N_32130,N_27687,N_26023);
nor U32131 (N_32131,N_28034,N_25381);
and U32132 (N_32132,N_28283,N_27255);
or U32133 (N_32133,N_26753,N_29424);
xor U32134 (N_32134,N_26315,N_27288);
or U32135 (N_32135,N_27233,N_27858);
or U32136 (N_32136,N_25795,N_28454);
nand U32137 (N_32137,N_25343,N_29899);
and U32138 (N_32138,N_29969,N_27282);
nor U32139 (N_32139,N_25622,N_25300);
and U32140 (N_32140,N_29084,N_28912);
and U32141 (N_32141,N_26337,N_28164);
or U32142 (N_32142,N_29812,N_27763);
nor U32143 (N_32143,N_29020,N_25059);
nand U32144 (N_32144,N_26256,N_26787);
xnor U32145 (N_32145,N_26415,N_26882);
xnor U32146 (N_32146,N_28751,N_26700);
and U32147 (N_32147,N_27339,N_27460);
or U32148 (N_32148,N_28679,N_28090);
or U32149 (N_32149,N_28668,N_27495);
nand U32150 (N_32150,N_26879,N_26668);
or U32151 (N_32151,N_28757,N_28460);
nor U32152 (N_32152,N_27733,N_26761);
nand U32153 (N_32153,N_26511,N_27420);
xnor U32154 (N_32154,N_29971,N_25819);
xor U32155 (N_32155,N_25203,N_29797);
xor U32156 (N_32156,N_28981,N_25057);
or U32157 (N_32157,N_29919,N_28894);
or U32158 (N_32158,N_27927,N_29615);
xnor U32159 (N_32159,N_29030,N_26842);
nor U32160 (N_32160,N_27755,N_25838);
nor U32161 (N_32161,N_26513,N_27666);
nor U32162 (N_32162,N_27405,N_27746);
and U32163 (N_32163,N_27628,N_26645);
nor U32164 (N_32164,N_29720,N_29375);
xnor U32165 (N_32165,N_29997,N_27692);
nor U32166 (N_32166,N_27952,N_28688);
or U32167 (N_32167,N_25775,N_26691);
or U32168 (N_32168,N_28781,N_28348);
nor U32169 (N_32169,N_27704,N_25889);
or U32170 (N_32170,N_29582,N_26166);
nand U32171 (N_32171,N_29471,N_26277);
and U32172 (N_32172,N_25983,N_28720);
xnor U32173 (N_32173,N_25231,N_28435);
or U32174 (N_32174,N_28707,N_25539);
nand U32175 (N_32175,N_29542,N_29832);
nand U32176 (N_32176,N_25537,N_28049);
xnor U32177 (N_32177,N_29779,N_27955);
nor U32178 (N_32178,N_29523,N_29091);
xor U32179 (N_32179,N_29731,N_26297);
nor U32180 (N_32180,N_28664,N_27509);
xnor U32181 (N_32181,N_26591,N_25582);
xnor U32182 (N_32182,N_29517,N_27831);
and U32183 (N_32183,N_27932,N_29537);
or U32184 (N_32184,N_27979,N_26798);
nor U32185 (N_32185,N_26590,N_29054);
or U32186 (N_32186,N_26763,N_28018);
or U32187 (N_32187,N_25947,N_28350);
xor U32188 (N_32188,N_26334,N_29409);
or U32189 (N_32189,N_25060,N_27717);
and U32190 (N_32190,N_28545,N_25849);
and U32191 (N_32191,N_28939,N_26725);
or U32192 (N_32192,N_25721,N_28765);
nand U32193 (N_32193,N_25252,N_25748);
and U32194 (N_32194,N_27725,N_25253);
nand U32195 (N_32195,N_26762,N_25307);
nor U32196 (N_32196,N_25771,N_27528);
nand U32197 (N_32197,N_26232,N_25853);
and U32198 (N_32198,N_25272,N_25151);
and U32199 (N_32199,N_26362,N_28553);
or U32200 (N_32200,N_25687,N_26946);
xor U32201 (N_32201,N_28085,N_28473);
xnor U32202 (N_32202,N_27962,N_27272);
nand U32203 (N_32203,N_28167,N_29119);
nand U32204 (N_32204,N_29461,N_26137);
and U32205 (N_32205,N_29639,N_25350);
nor U32206 (N_32206,N_25552,N_27546);
xor U32207 (N_32207,N_26111,N_28583);
nor U32208 (N_32208,N_28148,N_25905);
nand U32209 (N_32209,N_26336,N_25726);
and U32210 (N_32210,N_29341,N_28091);
nor U32211 (N_32211,N_29753,N_26993);
or U32212 (N_32212,N_26285,N_29620);
or U32213 (N_32213,N_28873,N_25035);
nand U32214 (N_32214,N_28925,N_28221);
and U32215 (N_32215,N_25564,N_25785);
and U32216 (N_32216,N_25314,N_26369);
or U32217 (N_32217,N_28839,N_29902);
and U32218 (N_32218,N_28309,N_27579);
nand U32219 (N_32219,N_27328,N_28738);
nor U32220 (N_32220,N_25864,N_26186);
nand U32221 (N_32221,N_29098,N_29686);
and U32222 (N_32222,N_29484,N_25680);
nor U32223 (N_32223,N_27373,N_26679);
or U32224 (N_32224,N_25942,N_25767);
xnor U32225 (N_32225,N_29426,N_28512);
nor U32226 (N_32226,N_27166,N_27348);
and U32227 (N_32227,N_28331,N_26890);
or U32228 (N_32228,N_27369,N_29344);
nor U32229 (N_32229,N_26925,N_29354);
nor U32230 (N_32230,N_26652,N_28445);
or U32231 (N_32231,N_27624,N_27383);
xnor U32232 (N_32232,N_28488,N_27136);
nand U32233 (N_32233,N_25642,N_29047);
nand U32234 (N_32234,N_26145,N_29215);
or U32235 (N_32235,N_29143,N_28754);
xor U32236 (N_32236,N_27472,N_25404);
or U32237 (N_32237,N_26242,N_26239);
nor U32238 (N_32238,N_25684,N_25483);
nand U32239 (N_32239,N_25176,N_29633);
or U32240 (N_32240,N_27683,N_29663);
xnor U32241 (N_32241,N_27775,N_27976);
xnor U32242 (N_32242,N_28785,N_29928);
xnor U32243 (N_32243,N_25258,N_29415);
nand U32244 (N_32244,N_25214,N_29961);
xor U32245 (N_32245,N_28703,N_26210);
or U32246 (N_32246,N_28323,N_25438);
xnor U32247 (N_32247,N_27468,N_26135);
xor U32248 (N_32248,N_26980,N_29824);
or U32249 (N_32249,N_25971,N_25326);
and U32250 (N_32250,N_29952,N_25654);
nand U32251 (N_32251,N_27585,N_28739);
or U32252 (N_32252,N_29336,N_25990);
or U32253 (N_32253,N_25792,N_29289);
or U32254 (N_32254,N_27640,N_26770);
nor U32255 (N_32255,N_25055,N_28580);
and U32256 (N_32256,N_25003,N_25367);
and U32257 (N_32257,N_26422,N_28199);
and U32258 (N_32258,N_28525,N_25461);
or U32259 (N_32259,N_25315,N_27250);
xnor U32260 (N_32260,N_27806,N_26637);
xor U32261 (N_32261,N_28698,N_28550);
nand U32262 (N_32262,N_25323,N_25928);
xor U32263 (N_32263,N_26108,N_28717);
or U32264 (N_32264,N_27911,N_25247);
nor U32265 (N_32265,N_26273,N_27262);
xnor U32266 (N_32266,N_26010,N_26270);
nor U32267 (N_32267,N_25344,N_27225);
nand U32268 (N_32268,N_29872,N_27214);
or U32269 (N_32269,N_26066,N_26453);
xor U32270 (N_32270,N_25966,N_26611);
nand U32271 (N_32271,N_25646,N_26848);
xor U32272 (N_32272,N_29011,N_28905);
nor U32273 (N_32273,N_26806,N_28673);
nor U32274 (N_32274,N_27589,N_29514);
xnor U32275 (N_32275,N_25584,N_27029);
and U32276 (N_32276,N_26412,N_27438);
nand U32277 (N_32277,N_29701,N_28947);
and U32278 (N_32278,N_29991,N_25523);
and U32279 (N_32279,N_27864,N_29817);
nor U32280 (N_32280,N_29250,N_29612);
and U32281 (N_32281,N_26943,N_27561);
nor U32282 (N_32282,N_29181,N_28969);
xor U32283 (N_32283,N_29085,N_29028);
and U32284 (N_32284,N_26328,N_29177);
and U32285 (N_32285,N_26164,N_28975);
or U32286 (N_32286,N_26856,N_28833);
nor U32287 (N_32287,N_29550,N_29157);
nand U32288 (N_32288,N_27204,N_25310);
and U32289 (N_32289,N_25866,N_25896);
or U32290 (N_32290,N_27972,N_29475);
nor U32291 (N_32291,N_28214,N_27892);
nand U32292 (N_32292,N_26378,N_27884);
or U32293 (N_32293,N_25648,N_26893);
nor U32294 (N_32294,N_27143,N_29822);
xor U32295 (N_32295,N_27360,N_25455);
nor U32296 (N_32296,N_27726,N_28727);
xor U32297 (N_32297,N_25514,N_25398);
xnor U32298 (N_32298,N_29146,N_25040);
xnor U32299 (N_32299,N_27732,N_26687);
nor U32300 (N_32300,N_25351,N_26120);
nand U32301 (N_32301,N_26754,N_25281);
and U32302 (N_32302,N_25502,N_29486);
nand U32303 (N_32303,N_28940,N_29350);
or U32304 (N_32304,N_28193,N_27454);
nand U32305 (N_32305,N_27503,N_26236);
and U32306 (N_32306,N_29850,N_28955);
nand U32307 (N_32307,N_29044,N_25223);
nand U32308 (N_32308,N_26935,N_25891);
nor U32309 (N_32309,N_28472,N_28337);
xnor U32310 (N_32310,N_28623,N_27883);
nor U32311 (N_32311,N_27300,N_27350);
xnor U32312 (N_32312,N_27351,N_27530);
and U32313 (N_32313,N_25070,N_29741);
nand U32314 (N_32314,N_25843,N_26281);
xnor U32315 (N_32315,N_29116,N_27540);
xor U32316 (N_32316,N_26012,N_29267);
nand U32317 (N_32317,N_25970,N_27453);
xnor U32318 (N_32318,N_26157,N_27461);
nand U32319 (N_32319,N_29619,N_27141);
or U32320 (N_32320,N_27888,N_26976);
nor U32321 (N_32321,N_25190,N_27518);
nor U32322 (N_32322,N_29070,N_25250);
nand U32323 (N_32323,N_28501,N_29632);
nand U32324 (N_32324,N_29228,N_25946);
nand U32325 (N_32325,N_28056,N_26778);
nor U32326 (N_32326,N_28336,N_28361);
and U32327 (N_32327,N_29356,N_26707);
xor U32328 (N_32328,N_27919,N_25130);
or U32329 (N_32329,N_27498,N_28746);
nand U32330 (N_32330,N_25841,N_27870);
nand U32331 (N_32331,N_29265,N_29852);
nor U32332 (N_32332,N_26625,N_26550);
nand U32333 (N_32333,N_28786,N_27356);
nor U32334 (N_32334,N_27662,N_26015);
nor U32335 (N_32335,N_27465,N_27846);
xor U32336 (N_32336,N_26129,N_26249);
or U32337 (N_32337,N_29431,N_29787);
and U32338 (N_32338,N_25045,N_29038);
xor U32339 (N_32339,N_26564,N_28643);
xor U32340 (N_32340,N_25390,N_26081);
nand U32341 (N_32341,N_28800,N_28778);
nor U32342 (N_32342,N_29606,N_26579);
xnor U32343 (N_32343,N_25555,N_29922);
nand U32344 (N_32344,N_26830,N_25832);
nand U32345 (N_32345,N_25192,N_27140);
nand U32346 (N_32346,N_25550,N_29798);
or U32347 (N_32347,N_26915,N_28265);
or U32348 (N_32348,N_28891,N_29540);
xor U32349 (N_32349,N_25361,N_26998);
xnor U32350 (N_32350,N_28637,N_26571);
nand U32351 (N_32351,N_27137,N_25950);
and U32352 (N_32352,N_26694,N_25136);
and U32353 (N_32353,N_26448,N_25718);
xnor U32354 (N_32354,N_26089,N_27222);
xor U32355 (N_32355,N_27424,N_27885);
nor U32356 (N_32356,N_29538,N_25499);
nand U32357 (N_32357,N_28479,N_27273);
or U32358 (N_32358,N_27621,N_29051);
nand U32359 (N_32359,N_25349,N_25855);
nand U32360 (N_32360,N_27822,N_26722);
xor U32361 (N_32361,N_27922,N_27008);
xor U32362 (N_32362,N_25385,N_25392);
nand U32363 (N_32363,N_28006,N_26018);
nor U32364 (N_32364,N_26987,N_28450);
nand U32365 (N_32365,N_28313,N_29185);
nand U32366 (N_32366,N_27070,N_25704);
or U32367 (N_32367,N_27984,N_25191);
nand U32368 (N_32368,N_25675,N_26832);
nor U32369 (N_32369,N_26500,N_26820);
xor U32370 (N_32370,N_27829,N_25509);
nand U32371 (N_32371,N_25401,N_26656);
or U32372 (N_32372,N_29353,N_29300);
xnor U32373 (N_32373,N_29685,N_25278);
xnor U32374 (N_32374,N_29183,N_29213);
and U32375 (N_32375,N_29515,N_25613);
and U32376 (N_32376,N_25865,N_27306);
nor U32377 (N_32377,N_26950,N_29111);
nor U32378 (N_32378,N_26438,N_29163);
and U32379 (N_32379,N_28118,N_25031);
and U32380 (N_32380,N_29406,N_29449);
nor U32381 (N_32381,N_27597,N_29936);
nor U32382 (N_32382,N_27301,N_28878);
nand U32383 (N_32383,N_26200,N_28341);
xnor U32384 (N_32384,N_26248,N_25427);
or U32385 (N_32385,N_29708,N_27055);
or U32386 (N_32386,N_29938,N_26978);
xor U32387 (N_32387,N_29717,N_26260);
nor U32388 (N_32388,N_29107,N_27462);
or U32389 (N_32389,N_25172,N_29600);
or U32390 (N_32390,N_27410,N_29440);
and U32391 (N_32391,N_27126,N_28694);
nand U32392 (N_32392,N_29113,N_25397);
or U32393 (N_32393,N_29706,N_29784);
nor U32394 (N_32394,N_29016,N_28888);
xnor U32395 (N_32395,N_28848,N_29395);
nand U32396 (N_32396,N_26870,N_27064);
xnor U32397 (N_32397,N_26122,N_28497);
and U32398 (N_32398,N_26653,N_26000);
nand U32399 (N_32399,N_27758,N_28770);
nand U32400 (N_32400,N_26063,N_25496);
xor U32401 (N_32401,N_26586,N_26154);
nor U32402 (N_32402,N_29754,N_25491);
nand U32403 (N_32403,N_25915,N_28052);
nor U32404 (N_32404,N_27629,N_28078);
nand U32405 (N_32405,N_25412,N_27080);
and U32406 (N_32406,N_26044,N_26497);
and U32407 (N_32407,N_29805,N_26460);
nand U32408 (N_32408,N_28218,N_25493);
xor U32409 (N_32409,N_28543,N_27553);
nor U32410 (N_32410,N_28121,N_26600);
and U32411 (N_32411,N_27981,N_28005);
and U32412 (N_32412,N_25873,N_29008);
nand U32413 (N_32413,N_27765,N_26354);
nor U32414 (N_32414,N_25028,N_27874);
nand U32415 (N_32415,N_28825,N_28212);
nor U32416 (N_32416,N_27437,N_26517);
xor U32417 (N_32417,N_29342,N_26684);
or U32418 (N_32418,N_28964,N_27788);
nor U32419 (N_32419,N_27794,N_25518);
or U32420 (N_32420,N_27833,N_27500);
xnor U32421 (N_32421,N_29277,N_26721);
and U32422 (N_32422,N_27887,N_26482);
or U32423 (N_32423,N_25177,N_26189);
and U32424 (N_32424,N_26695,N_28849);
nor U32425 (N_32425,N_26974,N_25071);
and U32426 (N_32426,N_26752,N_27841);
nor U32427 (N_32427,N_29765,N_25912);
nand U32428 (N_32428,N_27400,N_28853);
xnor U32429 (N_32429,N_25917,N_26384);
nand U32430 (N_32430,N_29654,N_29972);
and U32431 (N_32431,N_29374,N_26302);
and U32432 (N_32432,N_29255,N_26356);
nor U32433 (N_32433,N_29740,N_27040);
nand U32434 (N_32434,N_29684,N_26011);
xnor U32435 (N_32435,N_28671,N_25714);
and U32436 (N_32436,N_27149,N_26470);
nor U32437 (N_32437,N_27918,N_27367);
xnor U32438 (N_32438,N_27519,N_25105);
or U32439 (N_32439,N_28303,N_25394);
or U32440 (N_32440,N_29458,N_26703);
xnor U32441 (N_32441,N_26549,N_26492);
or U32442 (N_32442,N_25022,N_26068);
and U32443 (N_32443,N_25922,N_29175);
or U32444 (N_32444,N_28531,N_25902);
and U32445 (N_32445,N_27825,N_28882);
and U32446 (N_32446,N_25594,N_25485);
and U32447 (N_32447,N_28628,N_29367);
nand U32448 (N_32448,N_25213,N_27525);
nor U32449 (N_32449,N_26938,N_25565);
and U32450 (N_32450,N_29387,N_26144);
xor U32451 (N_32451,N_28985,N_27722);
nor U32452 (N_32452,N_26597,N_27017);
nor U32453 (N_32453,N_29937,N_25008);
nor U32454 (N_32454,N_25751,N_28316);
xnor U32455 (N_32455,N_28222,N_28041);
nor U32456 (N_32456,N_26897,N_29192);
xor U32457 (N_32457,N_25112,N_28423);
nor U32458 (N_32458,N_28421,N_28354);
or U32459 (N_32459,N_28674,N_26593);
or U32460 (N_32460,N_28677,N_25717);
xnor U32461 (N_32461,N_27362,N_25977);
nor U32462 (N_32462,N_27912,N_25052);
nand U32463 (N_32463,N_28729,N_27387);
xor U32464 (N_32464,N_26568,N_27802);
and U32465 (N_32465,N_27512,N_29963);
nor U32466 (N_32466,N_26555,N_28245);
xnor U32467 (N_32467,N_28804,N_27963);
xnor U32468 (N_32468,N_25796,N_29830);
nor U32469 (N_32469,N_29482,N_26152);
nor U32470 (N_32470,N_25056,N_27877);
nand U32471 (N_32471,N_25763,N_29987);
and U32472 (N_32472,N_27882,N_25383);
and U32473 (N_32473,N_28588,N_29142);
nor U32474 (N_32474,N_29281,N_29891);
and U32475 (N_32475,N_28808,N_29416);
nand U32476 (N_32476,N_27216,N_26255);
or U32477 (N_32477,N_28977,N_26291);
and U32478 (N_32478,N_28032,N_28921);
nand U32479 (N_32479,N_29075,N_28456);
nand U32480 (N_32480,N_29071,N_26970);
or U32481 (N_32481,N_25612,N_25810);
or U32482 (N_32482,N_26578,N_29172);
nor U32483 (N_32483,N_29083,N_27361);
xnor U32484 (N_32484,N_28429,N_28557);
and U32485 (N_32485,N_27172,N_25072);
or U32486 (N_32486,N_27425,N_28210);
xor U32487 (N_32487,N_27959,N_26956);
nor U32488 (N_32488,N_25423,N_26847);
nand U32489 (N_32489,N_29121,N_25497);
xor U32490 (N_32490,N_28014,N_25735);
and U32491 (N_32491,N_26912,N_25293);
nor U32492 (N_32492,N_25822,N_25403);
and U32493 (N_32493,N_26598,N_27432);
xor U32494 (N_32494,N_26932,N_29063);
and U32495 (N_32495,N_28622,N_29748);
xnor U32496 (N_32496,N_28547,N_25005);
nor U32497 (N_32497,N_25593,N_28478);
and U32498 (N_32498,N_25117,N_25906);
xnor U32499 (N_32499,N_27321,N_26219);
and U32500 (N_32500,N_28183,N_27126);
nor U32501 (N_32501,N_26636,N_27456);
nand U32502 (N_32502,N_27821,N_29890);
nor U32503 (N_32503,N_28957,N_25047);
nand U32504 (N_32504,N_29644,N_25670);
or U32505 (N_32505,N_25187,N_28348);
nand U32506 (N_32506,N_28388,N_29705);
or U32507 (N_32507,N_26159,N_28147);
xnor U32508 (N_32508,N_29364,N_27001);
or U32509 (N_32509,N_26607,N_25961);
xor U32510 (N_32510,N_26577,N_29845);
or U32511 (N_32511,N_28396,N_29588);
xnor U32512 (N_32512,N_28214,N_26410);
nor U32513 (N_32513,N_25433,N_29677);
nand U32514 (N_32514,N_29802,N_25752);
nand U32515 (N_32515,N_25012,N_26893);
and U32516 (N_32516,N_29500,N_27207);
and U32517 (N_32517,N_29796,N_28541);
nor U32518 (N_32518,N_28592,N_29618);
xnor U32519 (N_32519,N_28132,N_26708);
xor U32520 (N_32520,N_28205,N_27517);
and U32521 (N_32521,N_27984,N_28191);
or U32522 (N_32522,N_28511,N_26388);
xnor U32523 (N_32523,N_29221,N_27393);
or U32524 (N_32524,N_26912,N_27632);
xnor U32525 (N_32525,N_25749,N_28194);
and U32526 (N_32526,N_26269,N_28823);
nand U32527 (N_32527,N_28548,N_27616);
xor U32528 (N_32528,N_26404,N_27311);
or U32529 (N_32529,N_27145,N_27790);
nor U32530 (N_32530,N_28056,N_27629);
and U32531 (N_32531,N_26918,N_27039);
nand U32532 (N_32532,N_25579,N_29719);
or U32533 (N_32533,N_28141,N_25027);
xnor U32534 (N_32534,N_27105,N_27768);
xor U32535 (N_32535,N_29052,N_25160);
nor U32536 (N_32536,N_27632,N_29560);
and U32537 (N_32537,N_28788,N_26390);
xnor U32538 (N_32538,N_27927,N_27722);
nor U32539 (N_32539,N_26525,N_28804);
and U32540 (N_32540,N_28948,N_26689);
or U32541 (N_32541,N_25692,N_25973);
nor U32542 (N_32542,N_27084,N_25646);
nor U32543 (N_32543,N_29338,N_25273);
nor U32544 (N_32544,N_27720,N_28154);
xor U32545 (N_32545,N_27109,N_29725);
nor U32546 (N_32546,N_28917,N_28722);
or U32547 (N_32547,N_29501,N_25395);
nand U32548 (N_32548,N_25112,N_25376);
nand U32549 (N_32549,N_29529,N_27222);
nand U32550 (N_32550,N_25787,N_26738);
or U32551 (N_32551,N_26759,N_25094);
or U32552 (N_32552,N_29322,N_28883);
nor U32553 (N_32553,N_29041,N_26509);
xnor U32554 (N_32554,N_27604,N_28953);
nor U32555 (N_32555,N_27970,N_28536);
nor U32556 (N_32556,N_27659,N_26453);
or U32557 (N_32557,N_28462,N_28956);
and U32558 (N_32558,N_26042,N_25336);
nand U32559 (N_32559,N_29045,N_28095);
and U32560 (N_32560,N_27204,N_25636);
nand U32561 (N_32561,N_25222,N_26761);
nand U32562 (N_32562,N_28467,N_29879);
and U32563 (N_32563,N_29493,N_27898);
or U32564 (N_32564,N_29683,N_29484);
and U32565 (N_32565,N_29129,N_29593);
nor U32566 (N_32566,N_28189,N_25922);
and U32567 (N_32567,N_28457,N_29853);
and U32568 (N_32568,N_26589,N_29351);
and U32569 (N_32569,N_29617,N_25216);
xnor U32570 (N_32570,N_27069,N_25490);
nor U32571 (N_32571,N_27528,N_26535);
and U32572 (N_32572,N_27978,N_29904);
and U32573 (N_32573,N_25147,N_27059);
or U32574 (N_32574,N_26824,N_25843);
nand U32575 (N_32575,N_27356,N_27525);
xnor U32576 (N_32576,N_26557,N_26808);
or U32577 (N_32577,N_27830,N_28578);
nor U32578 (N_32578,N_27845,N_25985);
or U32579 (N_32579,N_29244,N_27793);
nor U32580 (N_32580,N_25930,N_26641);
and U32581 (N_32581,N_28500,N_27439);
nand U32582 (N_32582,N_26975,N_26344);
or U32583 (N_32583,N_25221,N_29594);
and U32584 (N_32584,N_26192,N_29304);
nand U32585 (N_32585,N_25543,N_26448);
or U32586 (N_32586,N_29008,N_29152);
and U32587 (N_32587,N_27610,N_27331);
xnor U32588 (N_32588,N_27356,N_29725);
or U32589 (N_32589,N_28288,N_28124);
and U32590 (N_32590,N_26820,N_25202);
or U32591 (N_32591,N_27173,N_28736);
nand U32592 (N_32592,N_28093,N_28230);
nand U32593 (N_32593,N_27377,N_26121);
and U32594 (N_32594,N_29339,N_29961);
nand U32595 (N_32595,N_28853,N_25691);
xor U32596 (N_32596,N_25803,N_27237);
xnor U32597 (N_32597,N_27901,N_28146);
and U32598 (N_32598,N_27133,N_29681);
nand U32599 (N_32599,N_28210,N_29328);
nor U32600 (N_32600,N_27341,N_27751);
xnor U32601 (N_32601,N_25481,N_26431);
or U32602 (N_32602,N_26639,N_28818);
nor U32603 (N_32603,N_26184,N_26663);
or U32604 (N_32604,N_26197,N_26725);
nor U32605 (N_32605,N_26104,N_26715);
or U32606 (N_32606,N_27537,N_26649);
nor U32607 (N_32607,N_26805,N_27848);
or U32608 (N_32608,N_29565,N_29329);
and U32609 (N_32609,N_26099,N_25643);
nor U32610 (N_32610,N_25088,N_25612);
or U32611 (N_32611,N_26873,N_26077);
and U32612 (N_32612,N_26012,N_25162);
xnor U32613 (N_32613,N_29340,N_27892);
xor U32614 (N_32614,N_28115,N_26734);
nor U32615 (N_32615,N_27694,N_26369);
nand U32616 (N_32616,N_27745,N_26042);
and U32617 (N_32617,N_29775,N_29069);
or U32618 (N_32618,N_28521,N_26407);
nor U32619 (N_32619,N_28579,N_28760);
or U32620 (N_32620,N_29585,N_29611);
and U32621 (N_32621,N_26731,N_29114);
nand U32622 (N_32622,N_29291,N_27140);
nor U32623 (N_32623,N_29478,N_27494);
nor U32624 (N_32624,N_26378,N_25304);
and U32625 (N_32625,N_28142,N_28625);
nor U32626 (N_32626,N_28247,N_28099);
nand U32627 (N_32627,N_26138,N_28987);
and U32628 (N_32628,N_25171,N_26416);
nor U32629 (N_32629,N_25928,N_25878);
xnor U32630 (N_32630,N_29324,N_28408);
or U32631 (N_32631,N_28726,N_29688);
xnor U32632 (N_32632,N_27395,N_27723);
and U32633 (N_32633,N_25852,N_25973);
and U32634 (N_32634,N_26521,N_29398);
nand U32635 (N_32635,N_29514,N_25536);
or U32636 (N_32636,N_25419,N_29142);
nand U32637 (N_32637,N_29948,N_25464);
and U32638 (N_32638,N_25519,N_28738);
nor U32639 (N_32639,N_25999,N_28120);
xor U32640 (N_32640,N_25307,N_26069);
or U32641 (N_32641,N_25799,N_26788);
or U32642 (N_32642,N_28630,N_26700);
nor U32643 (N_32643,N_25503,N_28522);
and U32644 (N_32644,N_26219,N_28888);
xnor U32645 (N_32645,N_28919,N_27358);
xnor U32646 (N_32646,N_26611,N_27416);
nor U32647 (N_32647,N_29266,N_27062);
or U32648 (N_32648,N_25102,N_26119);
or U32649 (N_32649,N_29199,N_27880);
nand U32650 (N_32650,N_29479,N_28255);
nor U32651 (N_32651,N_27512,N_25886);
xor U32652 (N_32652,N_28799,N_26238);
xor U32653 (N_32653,N_26501,N_29362);
nor U32654 (N_32654,N_28812,N_28829);
xnor U32655 (N_32655,N_25837,N_25916);
nand U32656 (N_32656,N_28018,N_27622);
and U32657 (N_32657,N_25933,N_29843);
nor U32658 (N_32658,N_25089,N_26813);
nand U32659 (N_32659,N_25384,N_25884);
nor U32660 (N_32660,N_28624,N_25745);
nor U32661 (N_32661,N_25401,N_27959);
nor U32662 (N_32662,N_28571,N_27979);
or U32663 (N_32663,N_27967,N_29474);
nor U32664 (N_32664,N_28593,N_28183);
and U32665 (N_32665,N_27926,N_28021);
nand U32666 (N_32666,N_27172,N_28136);
and U32667 (N_32667,N_27090,N_25371);
xnor U32668 (N_32668,N_25729,N_28329);
and U32669 (N_32669,N_25138,N_26059);
and U32670 (N_32670,N_27826,N_28878);
or U32671 (N_32671,N_26447,N_25477);
nor U32672 (N_32672,N_25716,N_28285);
and U32673 (N_32673,N_28811,N_28264);
xnor U32674 (N_32674,N_29392,N_28345);
and U32675 (N_32675,N_29157,N_26502);
or U32676 (N_32676,N_26281,N_28011);
nor U32677 (N_32677,N_27517,N_27121);
nand U32678 (N_32678,N_26880,N_26323);
or U32679 (N_32679,N_25282,N_25017);
nand U32680 (N_32680,N_27086,N_27743);
nand U32681 (N_32681,N_27401,N_27781);
and U32682 (N_32682,N_29933,N_25838);
nor U32683 (N_32683,N_29712,N_26681);
or U32684 (N_32684,N_26939,N_28881);
xor U32685 (N_32685,N_29508,N_28714);
xnor U32686 (N_32686,N_28772,N_28248);
nand U32687 (N_32687,N_25287,N_26899);
or U32688 (N_32688,N_25098,N_25712);
or U32689 (N_32689,N_29151,N_26994);
nor U32690 (N_32690,N_26451,N_29884);
xor U32691 (N_32691,N_28831,N_29860);
xnor U32692 (N_32692,N_25992,N_25043);
or U32693 (N_32693,N_26011,N_25729);
or U32694 (N_32694,N_29447,N_26379);
or U32695 (N_32695,N_25835,N_28698);
xnor U32696 (N_32696,N_29460,N_29144);
and U32697 (N_32697,N_28227,N_26322);
or U32698 (N_32698,N_25868,N_26685);
xnor U32699 (N_32699,N_27643,N_29975);
and U32700 (N_32700,N_26786,N_26868);
xor U32701 (N_32701,N_25020,N_26096);
nor U32702 (N_32702,N_28790,N_27789);
xnor U32703 (N_32703,N_29076,N_29348);
xor U32704 (N_32704,N_28141,N_26208);
xor U32705 (N_32705,N_29672,N_25471);
and U32706 (N_32706,N_25320,N_26579);
nand U32707 (N_32707,N_28230,N_25409);
nor U32708 (N_32708,N_26327,N_25542);
nor U32709 (N_32709,N_26429,N_27088);
nand U32710 (N_32710,N_29682,N_26911);
nor U32711 (N_32711,N_25032,N_25300);
and U32712 (N_32712,N_29261,N_27530);
xor U32713 (N_32713,N_28743,N_29259);
xor U32714 (N_32714,N_29926,N_25442);
or U32715 (N_32715,N_27402,N_26691);
nand U32716 (N_32716,N_26657,N_27190);
xnor U32717 (N_32717,N_28374,N_27962);
or U32718 (N_32718,N_28426,N_29693);
nor U32719 (N_32719,N_26788,N_27132);
nor U32720 (N_32720,N_28349,N_26280);
and U32721 (N_32721,N_26447,N_29669);
and U32722 (N_32722,N_29791,N_26650);
xor U32723 (N_32723,N_28407,N_28956);
and U32724 (N_32724,N_28736,N_25367);
nor U32725 (N_32725,N_25850,N_26769);
xnor U32726 (N_32726,N_26194,N_28794);
nand U32727 (N_32727,N_25259,N_29253);
or U32728 (N_32728,N_27076,N_29162);
nand U32729 (N_32729,N_29360,N_25129);
nand U32730 (N_32730,N_27865,N_29434);
and U32731 (N_32731,N_29289,N_25171);
nor U32732 (N_32732,N_25466,N_29877);
or U32733 (N_32733,N_25816,N_25461);
or U32734 (N_32734,N_28914,N_27766);
or U32735 (N_32735,N_29523,N_28630);
xnor U32736 (N_32736,N_26729,N_25941);
or U32737 (N_32737,N_27656,N_25111);
or U32738 (N_32738,N_29830,N_26591);
and U32739 (N_32739,N_28000,N_26591);
and U32740 (N_32740,N_26213,N_29653);
and U32741 (N_32741,N_26289,N_25187);
and U32742 (N_32742,N_26481,N_25184);
xor U32743 (N_32743,N_26952,N_28162);
nand U32744 (N_32744,N_26624,N_25188);
nor U32745 (N_32745,N_28207,N_26051);
nor U32746 (N_32746,N_28861,N_29858);
and U32747 (N_32747,N_26670,N_29528);
nor U32748 (N_32748,N_27920,N_25367);
and U32749 (N_32749,N_29083,N_25008);
or U32750 (N_32750,N_25455,N_27507);
or U32751 (N_32751,N_29185,N_27559);
nand U32752 (N_32752,N_26992,N_27835);
and U32753 (N_32753,N_29496,N_28884);
nor U32754 (N_32754,N_29313,N_27135);
xor U32755 (N_32755,N_28408,N_26250);
nor U32756 (N_32756,N_26895,N_27725);
or U32757 (N_32757,N_25774,N_26400);
xnor U32758 (N_32758,N_29904,N_29641);
nor U32759 (N_32759,N_25903,N_26176);
and U32760 (N_32760,N_26424,N_29000);
nor U32761 (N_32761,N_28466,N_28130);
nor U32762 (N_32762,N_27871,N_26973);
xor U32763 (N_32763,N_29988,N_27164);
xnor U32764 (N_32764,N_27106,N_26220);
and U32765 (N_32765,N_29417,N_28152);
and U32766 (N_32766,N_27641,N_28444);
and U32767 (N_32767,N_28717,N_25982);
nand U32768 (N_32768,N_25332,N_26789);
xor U32769 (N_32769,N_28758,N_25819);
xor U32770 (N_32770,N_26485,N_27791);
nor U32771 (N_32771,N_25816,N_25968);
nor U32772 (N_32772,N_26504,N_25237);
nand U32773 (N_32773,N_28669,N_26640);
nand U32774 (N_32774,N_25578,N_29970);
xor U32775 (N_32775,N_28876,N_26355);
nor U32776 (N_32776,N_27180,N_29119);
nor U32777 (N_32777,N_28315,N_25284);
xnor U32778 (N_32778,N_28241,N_26907);
or U32779 (N_32779,N_29123,N_28838);
xnor U32780 (N_32780,N_25014,N_26062);
xnor U32781 (N_32781,N_25286,N_29426);
or U32782 (N_32782,N_28064,N_25857);
and U32783 (N_32783,N_26271,N_25225);
and U32784 (N_32784,N_25801,N_29457);
or U32785 (N_32785,N_28959,N_27253);
nor U32786 (N_32786,N_28870,N_25218);
nor U32787 (N_32787,N_29874,N_28875);
nand U32788 (N_32788,N_29024,N_28680);
xor U32789 (N_32789,N_29937,N_25509);
or U32790 (N_32790,N_27231,N_26204);
or U32791 (N_32791,N_26598,N_28444);
xnor U32792 (N_32792,N_25243,N_25437);
and U32793 (N_32793,N_25709,N_27467);
xnor U32794 (N_32794,N_28269,N_29401);
nor U32795 (N_32795,N_25821,N_26248);
and U32796 (N_32796,N_29201,N_26160);
or U32797 (N_32797,N_29971,N_26579);
or U32798 (N_32798,N_25683,N_25624);
or U32799 (N_32799,N_28473,N_26066);
xnor U32800 (N_32800,N_28467,N_27384);
nor U32801 (N_32801,N_25711,N_27983);
nand U32802 (N_32802,N_29766,N_26726);
or U32803 (N_32803,N_26928,N_28959);
nor U32804 (N_32804,N_25395,N_25067);
xor U32805 (N_32805,N_27216,N_29717);
nor U32806 (N_32806,N_26290,N_27406);
xnor U32807 (N_32807,N_26439,N_27217);
or U32808 (N_32808,N_29427,N_28050);
and U32809 (N_32809,N_29738,N_27669);
nand U32810 (N_32810,N_25577,N_25414);
nor U32811 (N_32811,N_29177,N_26516);
and U32812 (N_32812,N_26930,N_27104);
nand U32813 (N_32813,N_27700,N_26614);
nand U32814 (N_32814,N_25147,N_27190);
and U32815 (N_32815,N_28756,N_28203);
or U32816 (N_32816,N_26703,N_29898);
nand U32817 (N_32817,N_27944,N_29400);
and U32818 (N_32818,N_28888,N_29444);
or U32819 (N_32819,N_27782,N_25507);
and U32820 (N_32820,N_25628,N_28075);
nand U32821 (N_32821,N_29080,N_27878);
and U32822 (N_32822,N_27507,N_26467);
nor U32823 (N_32823,N_26035,N_27929);
or U32824 (N_32824,N_25183,N_29405);
nor U32825 (N_32825,N_25027,N_29795);
nand U32826 (N_32826,N_25650,N_25658);
xor U32827 (N_32827,N_25348,N_27722);
nand U32828 (N_32828,N_28752,N_27658);
nor U32829 (N_32829,N_25623,N_28629);
nor U32830 (N_32830,N_25655,N_27261);
nand U32831 (N_32831,N_26851,N_26441);
nor U32832 (N_32832,N_27319,N_26242);
and U32833 (N_32833,N_29633,N_25782);
nor U32834 (N_32834,N_25926,N_28274);
nor U32835 (N_32835,N_27535,N_26613);
nand U32836 (N_32836,N_28393,N_29452);
or U32837 (N_32837,N_27110,N_29260);
xnor U32838 (N_32838,N_25943,N_29387);
xor U32839 (N_32839,N_25061,N_29019);
or U32840 (N_32840,N_26501,N_25124);
nor U32841 (N_32841,N_28568,N_29089);
nand U32842 (N_32842,N_25390,N_29216);
or U32843 (N_32843,N_26705,N_25457);
nand U32844 (N_32844,N_27383,N_28631);
or U32845 (N_32845,N_26155,N_28941);
nor U32846 (N_32846,N_29913,N_25244);
nand U32847 (N_32847,N_25221,N_27705);
or U32848 (N_32848,N_27799,N_29701);
nand U32849 (N_32849,N_26662,N_27432);
nand U32850 (N_32850,N_26030,N_26605);
or U32851 (N_32851,N_29366,N_28273);
and U32852 (N_32852,N_27703,N_27331);
xnor U32853 (N_32853,N_27644,N_25862);
or U32854 (N_32854,N_26460,N_26384);
and U32855 (N_32855,N_28537,N_26474);
and U32856 (N_32856,N_29558,N_26363);
or U32857 (N_32857,N_26584,N_29343);
nor U32858 (N_32858,N_29380,N_28048);
and U32859 (N_32859,N_29714,N_27880);
or U32860 (N_32860,N_29840,N_29498);
or U32861 (N_32861,N_25805,N_28926);
and U32862 (N_32862,N_25540,N_29809);
nand U32863 (N_32863,N_29918,N_27573);
nor U32864 (N_32864,N_28852,N_28807);
and U32865 (N_32865,N_29625,N_25022);
and U32866 (N_32866,N_27588,N_28350);
nand U32867 (N_32867,N_29180,N_26921);
and U32868 (N_32868,N_28506,N_25167);
nor U32869 (N_32869,N_28365,N_25229);
xor U32870 (N_32870,N_27015,N_28959);
nor U32871 (N_32871,N_29889,N_27395);
xor U32872 (N_32872,N_29150,N_29720);
nor U32873 (N_32873,N_27896,N_28928);
nor U32874 (N_32874,N_25402,N_25668);
nand U32875 (N_32875,N_26953,N_29384);
nand U32876 (N_32876,N_26245,N_29733);
or U32877 (N_32877,N_25778,N_27651);
xor U32878 (N_32878,N_25707,N_26615);
or U32879 (N_32879,N_25092,N_27410);
nand U32880 (N_32880,N_26673,N_29504);
nand U32881 (N_32881,N_27409,N_27435);
nand U32882 (N_32882,N_28962,N_26201);
xor U32883 (N_32883,N_25184,N_28395);
and U32884 (N_32884,N_29111,N_29198);
nor U32885 (N_32885,N_28469,N_26513);
nand U32886 (N_32886,N_25330,N_29871);
and U32887 (N_32887,N_28377,N_27901);
xor U32888 (N_32888,N_25423,N_29652);
nor U32889 (N_32889,N_27558,N_29702);
nand U32890 (N_32890,N_26753,N_28365);
or U32891 (N_32891,N_26793,N_26362);
or U32892 (N_32892,N_27647,N_28114);
nand U32893 (N_32893,N_28875,N_29642);
or U32894 (N_32894,N_27470,N_29398);
xnor U32895 (N_32895,N_27417,N_28388);
or U32896 (N_32896,N_26297,N_28822);
nand U32897 (N_32897,N_25128,N_26012);
xnor U32898 (N_32898,N_29757,N_28934);
nor U32899 (N_32899,N_28982,N_28126);
and U32900 (N_32900,N_27398,N_29647);
xnor U32901 (N_32901,N_25846,N_25252);
xnor U32902 (N_32902,N_25676,N_29862);
nand U32903 (N_32903,N_26376,N_29411);
or U32904 (N_32904,N_29670,N_29050);
nand U32905 (N_32905,N_26894,N_28152);
xnor U32906 (N_32906,N_26261,N_29363);
xnor U32907 (N_32907,N_27742,N_29828);
or U32908 (N_32908,N_25807,N_28957);
nand U32909 (N_32909,N_26476,N_28057);
nor U32910 (N_32910,N_28863,N_26828);
or U32911 (N_32911,N_28861,N_25420);
nor U32912 (N_32912,N_29437,N_29105);
nand U32913 (N_32913,N_27914,N_28066);
nor U32914 (N_32914,N_28937,N_27327);
nor U32915 (N_32915,N_25648,N_25857);
nand U32916 (N_32916,N_26736,N_27395);
nor U32917 (N_32917,N_27308,N_27475);
nor U32918 (N_32918,N_26071,N_27771);
xnor U32919 (N_32919,N_29650,N_25388);
or U32920 (N_32920,N_28631,N_27299);
nand U32921 (N_32921,N_27688,N_28358);
nand U32922 (N_32922,N_25063,N_27652);
and U32923 (N_32923,N_26025,N_28747);
xnor U32924 (N_32924,N_26296,N_27327);
nor U32925 (N_32925,N_25269,N_25704);
and U32926 (N_32926,N_25884,N_29132);
xor U32927 (N_32927,N_27258,N_26616);
xnor U32928 (N_32928,N_26772,N_26512);
xor U32929 (N_32929,N_25204,N_27003);
or U32930 (N_32930,N_28871,N_26303);
and U32931 (N_32931,N_28343,N_25902);
and U32932 (N_32932,N_26045,N_29420);
or U32933 (N_32933,N_27842,N_28709);
nand U32934 (N_32934,N_28012,N_25666);
nor U32935 (N_32935,N_27619,N_29065);
xnor U32936 (N_32936,N_29711,N_26453);
nand U32937 (N_32937,N_28193,N_28080);
or U32938 (N_32938,N_29303,N_28883);
or U32939 (N_32939,N_25184,N_27871);
or U32940 (N_32940,N_27811,N_26185);
or U32941 (N_32941,N_27605,N_26948);
xor U32942 (N_32942,N_29060,N_28104);
and U32943 (N_32943,N_27909,N_26134);
nor U32944 (N_32944,N_28808,N_26538);
and U32945 (N_32945,N_29839,N_27390);
and U32946 (N_32946,N_26908,N_29236);
nor U32947 (N_32947,N_25900,N_25649);
or U32948 (N_32948,N_26579,N_28220);
and U32949 (N_32949,N_29393,N_25567);
or U32950 (N_32950,N_27101,N_27884);
nand U32951 (N_32951,N_28383,N_28998);
or U32952 (N_32952,N_25472,N_27344);
and U32953 (N_32953,N_28965,N_27605);
xnor U32954 (N_32954,N_26963,N_25658);
nor U32955 (N_32955,N_28563,N_25187);
or U32956 (N_32956,N_25587,N_28820);
and U32957 (N_32957,N_29768,N_28202);
nand U32958 (N_32958,N_29179,N_27112);
or U32959 (N_32959,N_26911,N_27484);
or U32960 (N_32960,N_28041,N_27523);
nand U32961 (N_32961,N_28229,N_29982);
or U32962 (N_32962,N_28622,N_29957);
and U32963 (N_32963,N_27268,N_27296);
nor U32964 (N_32964,N_25751,N_29501);
xor U32965 (N_32965,N_25916,N_27645);
xor U32966 (N_32966,N_28739,N_26326);
xor U32967 (N_32967,N_25265,N_27757);
nand U32968 (N_32968,N_28105,N_28852);
nor U32969 (N_32969,N_28532,N_25048);
nor U32970 (N_32970,N_26200,N_27488);
nor U32971 (N_32971,N_25364,N_25557);
or U32972 (N_32972,N_27185,N_26949);
or U32973 (N_32973,N_28898,N_27573);
or U32974 (N_32974,N_28623,N_25085);
nand U32975 (N_32975,N_25401,N_28506);
nand U32976 (N_32976,N_28336,N_26442);
xor U32977 (N_32977,N_27228,N_28830);
nor U32978 (N_32978,N_29312,N_27143);
xnor U32979 (N_32979,N_26115,N_27422);
nor U32980 (N_32980,N_25767,N_25607);
nand U32981 (N_32981,N_28392,N_26484);
nand U32982 (N_32982,N_26321,N_26575);
and U32983 (N_32983,N_27793,N_27062);
nand U32984 (N_32984,N_27422,N_25287);
and U32985 (N_32985,N_27100,N_27134);
or U32986 (N_32986,N_27362,N_27796);
nor U32987 (N_32987,N_28646,N_29150);
nand U32988 (N_32988,N_28963,N_25480);
or U32989 (N_32989,N_27647,N_25866);
and U32990 (N_32990,N_28088,N_27253);
nand U32991 (N_32991,N_26041,N_29272);
xnor U32992 (N_32992,N_27335,N_28768);
or U32993 (N_32993,N_29248,N_27391);
and U32994 (N_32994,N_29042,N_26174);
xnor U32995 (N_32995,N_29506,N_27830);
xnor U32996 (N_32996,N_28518,N_25717);
nand U32997 (N_32997,N_28992,N_28131);
or U32998 (N_32998,N_29783,N_26850);
xnor U32999 (N_32999,N_29195,N_26684);
nand U33000 (N_33000,N_27905,N_29418);
nand U33001 (N_33001,N_27404,N_26630);
and U33002 (N_33002,N_26491,N_27948);
xor U33003 (N_33003,N_29199,N_25872);
xnor U33004 (N_33004,N_27467,N_27698);
nor U33005 (N_33005,N_28239,N_27204);
xnor U33006 (N_33006,N_28595,N_25822);
nand U33007 (N_33007,N_26396,N_27518);
nand U33008 (N_33008,N_26452,N_27370);
xor U33009 (N_33009,N_28744,N_29002);
or U33010 (N_33010,N_27808,N_28864);
xor U33011 (N_33011,N_25670,N_26118);
xnor U33012 (N_33012,N_26210,N_27756);
or U33013 (N_33013,N_28777,N_28367);
or U33014 (N_33014,N_28218,N_29555);
or U33015 (N_33015,N_26473,N_26474);
nor U33016 (N_33016,N_27451,N_25725);
xnor U33017 (N_33017,N_25150,N_27503);
xor U33018 (N_33018,N_28589,N_27887);
or U33019 (N_33019,N_27973,N_27038);
or U33020 (N_33020,N_29053,N_26948);
nor U33021 (N_33021,N_27317,N_27516);
and U33022 (N_33022,N_29597,N_25299);
xnor U33023 (N_33023,N_29013,N_28434);
xor U33024 (N_33024,N_26097,N_27829);
and U33025 (N_33025,N_27212,N_26566);
and U33026 (N_33026,N_26819,N_28073);
and U33027 (N_33027,N_28693,N_28687);
and U33028 (N_33028,N_27662,N_29495);
xnor U33029 (N_33029,N_25456,N_27719);
or U33030 (N_33030,N_27058,N_29109);
and U33031 (N_33031,N_28500,N_27489);
nor U33032 (N_33032,N_28360,N_26927);
nor U33033 (N_33033,N_27811,N_27594);
or U33034 (N_33034,N_26472,N_25364);
nand U33035 (N_33035,N_26241,N_28757);
and U33036 (N_33036,N_29515,N_27421);
xnor U33037 (N_33037,N_25202,N_28450);
or U33038 (N_33038,N_29931,N_26504);
or U33039 (N_33039,N_28790,N_29354);
or U33040 (N_33040,N_27199,N_29674);
nor U33041 (N_33041,N_26544,N_27356);
nand U33042 (N_33042,N_27594,N_27677);
nand U33043 (N_33043,N_27217,N_27906);
nand U33044 (N_33044,N_25919,N_26760);
nand U33045 (N_33045,N_25127,N_27484);
xnor U33046 (N_33046,N_28598,N_27653);
and U33047 (N_33047,N_29452,N_27149);
or U33048 (N_33048,N_28094,N_29223);
nor U33049 (N_33049,N_27947,N_25912);
xor U33050 (N_33050,N_28471,N_27450);
nand U33051 (N_33051,N_26001,N_29668);
xor U33052 (N_33052,N_27995,N_27731);
nand U33053 (N_33053,N_28213,N_25478);
xnor U33054 (N_33054,N_25765,N_29546);
or U33055 (N_33055,N_29857,N_29783);
nor U33056 (N_33056,N_25525,N_28789);
and U33057 (N_33057,N_28202,N_25369);
nor U33058 (N_33058,N_26940,N_29722);
nand U33059 (N_33059,N_29936,N_28163);
nand U33060 (N_33060,N_26546,N_25144);
and U33061 (N_33061,N_25705,N_26734);
or U33062 (N_33062,N_29676,N_26883);
and U33063 (N_33063,N_29608,N_28168);
and U33064 (N_33064,N_25167,N_29454);
and U33065 (N_33065,N_26439,N_27592);
and U33066 (N_33066,N_27387,N_29746);
xor U33067 (N_33067,N_28321,N_25190);
nor U33068 (N_33068,N_27498,N_25017);
nor U33069 (N_33069,N_29596,N_29926);
nor U33070 (N_33070,N_27261,N_29147);
or U33071 (N_33071,N_26394,N_26295);
xor U33072 (N_33072,N_25232,N_29028);
nor U33073 (N_33073,N_29060,N_27874);
nand U33074 (N_33074,N_28178,N_26316);
and U33075 (N_33075,N_27559,N_28711);
nor U33076 (N_33076,N_25963,N_28752);
and U33077 (N_33077,N_26941,N_29783);
and U33078 (N_33078,N_29865,N_26427);
nor U33079 (N_33079,N_25762,N_28285);
nor U33080 (N_33080,N_26070,N_26084);
xor U33081 (N_33081,N_25948,N_29874);
nand U33082 (N_33082,N_25995,N_29412);
nor U33083 (N_33083,N_25986,N_28368);
and U33084 (N_33084,N_28990,N_27318);
or U33085 (N_33085,N_25598,N_29333);
or U33086 (N_33086,N_25311,N_25613);
or U33087 (N_33087,N_27837,N_25302);
nand U33088 (N_33088,N_27286,N_27650);
xnor U33089 (N_33089,N_28695,N_26802);
nor U33090 (N_33090,N_25075,N_25775);
or U33091 (N_33091,N_27213,N_25822);
nand U33092 (N_33092,N_29385,N_29072);
or U33093 (N_33093,N_27850,N_29705);
xnor U33094 (N_33094,N_26731,N_26657);
and U33095 (N_33095,N_28772,N_27933);
xnor U33096 (N_33096,N_28111,N_27139);
and U33097 (N_33097,N_26334,N_25721);
nand U33098 (N_33098,N_28543,N_28350);
and U33099 (N_33099,N_29990,N_25972);
nor U33100 (N_33100,N_25796,N_26344);
or U33101 (N_33101,N_25195,N_28764);
xor U33102 (N_33102,N_26908,N_25947);
or U33103 (N_33103,N_26411,N_25367);
nand U33104 (N_33104,N_27381,N_28100);
nor U33105 (N_33105,N_25503,N_25074);
nand U33106 (N_33106,N_26756,N_29671);
nor U33107 (N_33107,N_27574,N_28110);
and U33108 (N_33108,N_27561,N_28575);
xor U33109 (N_33109,N_26262,N_25542);
or U33110 (N_33110,N_29814,N_29114);
or U33111 (N_33111,N_27948,N_26167);
and U33112 (N_33112,N_25975,N_28410);
nor U33113 (N_33113,N_28537,N_29079);
nor U33114 (N_33114,N_25215,N_26934);
or U33115 (N_33115,N_26896,N_25265);
and U33116 (N_33116,N_26989,N_29274);
nand U33117 (N_33117,N_28544,N_25785);
nor U33118 (N_33118,N_29562,N_29146);
xnor U33119 (N_33119,N_27372,N_29249);
nand U33120 (N_33120,N_26077,N_26662);
and U33121 (N_33121,N_29096,N_26151);
xnor U33122 (N_33122,N_25860,N_28145);
nand U33123 (N_33123,N_26355,N_28627);
and U33124 (N_33124,N_28244,N_26286);
nand U33125 (N_33125,N_28455,N_28826);
xnor U33126 (N_33126,N_28806,N_26312);
nand U33127 (N_33127,N_27172,N_25270);
and U33128 (N_33128,N_28837,N_25278);
and U33129 (N_33129,N_29225,N_27471);
or U33130 (N_33130,N_28093,N_28852);
and U33131 (N_33131,N_28336,N_29134);
nand U33132 (N_33132,N_27090,N_29059);
xor U33133 (N_33133,N_28510,N_28675);
xor U33134 (N_33134,N_27929,N_29735);
xnor U33135 (N_33135,N_25760,N_27638);
nand U33136 (N_33136,N_29353,N_28685);
nand U33137 (N_33137,N_28021,N_28601);
or U33138 (N_33138,N_27456,N_29240);
or U33139 (N_33139,N_27134,N_26308);
nor U33140 (N_33140,N_29965,N_28024);
nand U33141 (N_33141,N_29737,N_29881);
nand U33142 (N_33142,N_28745,N_26644);
xnor U33143 (N_33143,N_27416,N_28591);
or U33144 (N_33144,N_26543,N_26213);
nand U33145 (N_33145,N_28530,N_29797);
nand U33146 (N_33146,N_25393,N_29619);
nand U33147 (N_33147,N_28783,N_29763);
xor U33148 (N_33148,N_28945,N_26770);
nand U33149 (N_33149,N_26897,N_26951);
nand U33150 (N_33150,N_28593,N_25628);
and U33151 (N_33151,N_25139,N_28283);
or U33152 (N_33152,N_26743,N_27002);
or U33153 (N_33153,N_27499,N_28680);
nor U33154 (N_33154,N_25461,N_27812);
or U33155 (N_33155,N_26620,N_27573);
and U33156 (N_33156,N_28836,N_29159);
and U33157 (N_33157,N_26371,N_29255);
and U33158 (N_33158,N_28890,N_29448);
nor U33159 (N_33159,N_27825,N_28533);
nor U33160 (N_33160,N_28540,N_28699);
nand U33161 (N_33161,N_26006,N_27601);
nor U33162 (N_33162,N_27807,N_25624);
nor U33163 (N_33163,N_26905,N_28585);
or U33164 (N_33164,N_26423,N_26838);
and U33165 (N_33165,N_29056,N_28159);
or U33166 (N_33166,N_26788,N_26920);
xnor U33167 (N_33167,N_29570,N_28650);
nor U33168 (N_33168,N_25067,N_27886);
nor U33169 (N_33169,N_28056,N_25147);
nand U33170 (N_33170,N_25745,N_29754);
xor U33171 (N_33171,N_25207,N_27231);
xor U33172 (N_33172,N_29764,N_25905);
nor U33173 (N_33173,N_29858,N_27800);
xor U33174 (N_33174,N_28714,N_27122);
nand U33175 (N_33175,N_25168,N_27359);
xnor U33176 (N_33176,N_26671,N_25507);
nor U33177 (N_33177,N_27474,N_25289);
nand U33178 (N_33178,N_27094,N_26260);
and U33179 (N_33179,N_25170,N_27941);
nor U33180 (N_33180,N_25630,N_27279);
xnor U33181 (N_33181,N_27181,N_28718);
and U33182 (N_33182,N_27384,N_29454);
nor U33183 (N_33183,N_29305,N_28103);
nand U33184 (N_33184,N_26924,N_28172);
and U33185 (N_33185,N_28621,N_28715);
nand U33186 (N_33186,N_26668,N_26018);
nor U33187 (N_33187,N_25031,N_26707);
and U33188 (N_33188,N_29556,N_26891);
nand U33189 (N_33189,N_29833,N_27183);
xnor U33190 (N_33190,N_27245,N_28183);
nor U33191 (N_33191,N_28061,N_26377);
or U33192 (N_33192,N_28792,N_28069);
nand U33193 (N_33193,N_25930,N_27729);
and U33194 (N_33194,N_25853,N_25696);
nand U33195 (N_33195,N_28536,N_26669);
nand U33196 (N_33196,N_28758,N_25025);
xnor U33197 (N_33197,N_29693,N_25200);
xor U33198 (N_33198,N_29670,N_27287);
or U33199 (N_33199,N_25578,N_26260);
xnor U33200 (N_33200,N_29163,N_27979);
and U33201 (N_33201,N_25157,N_28617);
or U33202 (N_33202,N_26134,N_25694);
nand U33203 (N_33203,N_27320,N_26693);
nand U33204 (N_33204,N_25416,N_25978);
or U33205 (N_33205,N_27553,N_26564);
or U33206 (N_33206,N_28590,N_26076);
nor U33207 (N_33207,N_26455,N_28783);
nand U33208 (N_33208,N_29193,N_27644);
or U33209 (N_33209,N_28796,N_26401);
nand U33210 (N_33210,N_28578,N_28917);
nand U33211 (N_33211,N_27512,N_28648);
or U33212 (N_33212,N_28304,N_28882);
xnor U33213 (N_33213,N_28427,N_26963);
nand U33214 (N_33214,N_26224,N_29940);
and U33215 (N_33215,N_25493,N_27315);
or U33216 (N_33216,N_27770,N_29953);
and U33217 (N_33217,N_26577,N_29409);
xnor U33218 (N_33218,N_28894,N_29040);
nor U33219 (N_33219,N_29597,N_28894);
or U33220 (N_33220,N_26777,N_27621);
nor U33221 (N_33221,N_28976,N_25974);
and U33222 (N_33222,N_26064,N_29096);
xnor U33223 (N_33223,N_27882,N_25233);
nor U33224 (N_33224,N_27784,N_27476);
xor U33225 (N_33225,N_26177,N_27294);
and U33226 (N_33226,N_26456,N_26412);
nor U33227 (N_33227,N_26862,N_25835);
nor U33228 (N_33228,N_25777,N_28545);
nand U33229 (N_33229,N_29157,N_29778);
nor U33230 (N_33230,N_29413,N_29705);
nand U33231 (N_33231,N_28860,N_25661);
or U33232 (N_33232,N_26621,N_28235);
and U33233 (N_33233,N_25674,N_29158);
and U33234 (N_33234,N_25521,N_25637);
and U33235 (N_33235,N_26899,N_26092);
nand U33236 (N_33236,N_25796,N_25078);
nor U33237 (N_33237,N_27601,N_28404);
and U33238 (N_33238,N_26097,N_29480);
and U33239 (N_33239,N_26395,N_27470);
nor U33240 (N_33240,N_25562,N_27207);
and U33241 (N_33241,N_28016,N_27727);
or U33242 (N_33242,N_27227,N_26908);
xnor U33243 (N_33243,N_25858,N_25226);
nor U33244 (N_33244,N_25652,N_25010);
nor U33245 (N_33245,N_28358,N_27574);
xor U33246 (N_33246,N_26775,N_29101);
or U33247 (N_33247,N_25980,N_28204);
or U33248 (N_33248,N_27254,N_25487);
xor U33249 (N_33249,N_29670,N_25011);
and U33250 (N_33250,N_26567,N_27199);
or U33251 (N_33251,N_26014,N_29435);
and U33252 (N_33252,N_29338,N_25930);
or U33253 (N_33253,N_25822,N_28292);
xnor U33254 (N_33254,N_29509,N_27843);
nor U33255 (N_33255,N_29371,N_29009);
and U33256 (N_33256,N_25599,N_27451);
or U33257 (N_33257,N_26303,N_26517);
xor U33258 (N_33258,N_26757,N_26045);
and U33259 (N_33259,N_26063,N_25414);
and U33260 (N_33260,N_28713,N_25672);
nor U33261 (N_33261,N_26958,N_25833);
and U33262 (N_33262,N_25434,N_28488);
and U33263 (N_33263,N_26612,N_27919);
and U33264 (N_33264,N_25809,N_28152);
nand U33265 (N_33265,N_25239,N_25335);
or U33266 (N_33266,N_26633,N_25267);
xor U33267 (N_33267,N_27933,N_27132);
and U33268 (N_33268,N_29480,N_29158);
nand U33269 (N_33269,N_27008,N_29073);
or U33270 (N_33270,N_27600,N_26934);
nor U33271 (N_33271,N_25677,N_29861);
nor U33272 (N_33272,N_25308,N_26173);
xnor U33273 (N_33273,N_25124,N_28350);
or U33274 (N_33274,N_27120,N_28463);
nor U33275 (N_33275,N_26320,N_25670);
or U33276 (N_33276,N_27155,N_28119);
xor U33277 (N_33277,N_25488,N_27934);
and U33278 (N_33278,N_29704,N_26869);
nor U33279 (N_33279,N_28964,N_28460);
xnor U33280 (N_33280,N_26564,N_25716);
xor U33281 (N_33281,N_26334,N_29247);
xor U33282 (N_33282,N_26259,N_25223);
and U33283 (N_33283,N_29204,N_29384);
xnor U33284 (N_33284,N_26669,N_25393);
nor U33285 (N_33285,N_25079,N_28353);
and U33286 (N_33286,N_27115,N_26199);
or U33287 (N_33287,N_28608,N_29786);
and U33288 (N_33288,N_25145,N_29988);
xor U33289 (N_33289,N_27551,N_26461);
nand U33290 (N_33290,N_28112,N_25745);
and U33291 (N_33291,N_26211,N_27333);
nor U33292 (N_33292,N_26225,N_25581);
or U33293 (N_33293,N_29718,N_25449);
nor U33294 (N_33294,N_28118,N_29801);
or U33295 (N_33295,N_27963,N_26431);
or U33296 (N_33296,N_29069,N_25765);
xnor U33297 (N_33297,N_26688,N_29112);
and U33298 (N_33298,N_25310,N_27911);
or U33299 (N_33299,N_27585,N_29923);
xor U33300 (N_33300,N_29112,N_27456);
nand U33301 (N_33301,N_26150,N_26264);
and U33302 (N_33302,N_29732,N_29276);
nand U33303 (N_33303,N_28198,N_28732);
xor U33304 (N_33304,N_26561,N_26543);
and U33305 (N_33305,N_27725,N_25845);
xor U33306 (N_33306,N_29383,N_26634);
or U33307 (N_33307,N_29828,N_28162);
xnor U33308 (N_33308,N_26802,N_25079);
xor U33309 (N_33309,N_28100,N_26007);
nor U33310 (N_33310,N_26477,N_29992);
xnor U33311 (N_33311,N_29521,N_27694);
or U33312 (N_33312,N_26114,N_29456);
and U33313 (N_33313,N_27292,N_25853);
or U33314 (N_33314,N_26556,N_27088);
and U33315 (N_33315,N_29859,N_29098);
nor U33316 (N_33316,N_26878,N_28485);
and U33317 (N_33317,N_29731,N_29397);
nor U33318 (N_33318,N_28329,N_26979);
nand U33319 (N_33319,N_25590,N_29410);
nor U33320 (N_33320,N_26230,N_29715);
nor U33321 (N_33321,N_25520,N_27877);
nor U33322 (N_33322,N_26004,N_26094);
xnor U33323 (N_33323,N_29460,N_25715);
or U33324 (N_33324,N_28950,N_27349);
xor U33325 (N_33325,N_27893,N_28785);
nand U33326 (N_33326,N_26235,N_26973);
nand U33327 (N_33327,N_29547,N_28769);
nor U33328 (N_33328,N_27602,N_27006);
nor U33329 (N_33329,N_28773,N_26396);
and U33330 (N_33330,N_25462,N_27507);
and U33331 (N_33331,N_28717,N_29526);
or U33332 (N_33332,N_28641,N_29428);
nand U33333 (N_33333,N_29972,N_27071);
xnor U33334 (N_33334,N_26555,N_26706);
and U33335 (N_33335,N_28350,N_27823);
nor U33336 (N_33336,N_25657,N_26446);
and U33337 (N_33337,N_29977,N_28942);
nor U33338 (N_33338,N_28255,N_29390);
and U33339 (N_33339,N_25602,N_27699);
or U33340 (N_33340,N_27606,N_25627);
xor U33341 (N_33341,N_28691,N_27544);
nor U33342 (N_33342,N_27520,N_28405);
or U33343 (N_33343,N_28985,N_25088);
nor U33344 (N_33344,N_26069,N_27128);
and U33345 (N_33345,N_28730,N_28417);
and U33346 (N_33346,N_27985,N_28713);
nor U33347 (N_33347,N_25042,N_26777);
or U33348 (N_33348,N_28500,N_25597);
nor U33349 (N_33349,N_29031,N_28007);
nor U33350 (N_33350,N_26084,N_27294);
and U33351 (N_33351,N_29864,N_25788);
nor U33352 (N_33352,N_26491,N_28213);
xnor U33353 (N_33353,N_26349,N_29114);
nand U33354 (N_33354,N_27679,N_29102);
nor U33355 (N_33355,N_28687,N_27957);
nand U33356 (N_33356,N_29142,N_28727);
nor U33357 (N_33357,N_25611,N_25456);
xnor U33358 (N_33358,N_28223,N_25166);
or U33359 (N_33359,N_25024,N_28283);
nor U33360 (N_33360,N_25281,N_28289);
nand U33361 (N_33361,N_27771,N_29982);
or U33362 (N_33362,N_27403,N_25319);
or U33363 (N_33363,N_28084,N_27451);
nand U33364 (N_33364,N_27393,N_28575);
and U33365 (N_33365,N_28365,N_28054);
nor U33366 (N_33366,N_27157,N_27589);
nor U33367 (N_33367,N_25264,N_29771);
nor U33368 (N_33368,N_26645,N_26063);
nor U33369 (N_33369,N_25606,N_29618);
nand U33370 (N_33370,N_28641,N_27255);
nor U33371 (N_33371,N_26075,N_25357);
xor U33372 (N_33372,N_28448,N_25708);
or U33373 (N_33373,N_26726,N_26867);
and U33374 (N_33374,N_28111,N_28048);
or U33375 (N_33375,N_27667,N_28316);
xnor U33376 (N_33376,N_27741,N_26528);
xnor U33377 (N_33377,N_26009,N_28157);
xnor U33378 (N_33378,N_28432,N_27274);
and U33379 (N_33379,N_26747,N_29758);
or U33380 (N_33380,N_29317,N_28688);
xor U33381 (N_33381,N_27468,N_27495);
or U33382 (N_33382,N_25689,N_29750);
nand U33383 (N_33383,N_25208,N_27273);
nor U33384 (N_33384,N_29256,N_26319);
or U33385 (N_33385,N_25726,N_28391);
or U33386 (N_33386,N_29792,N_26558);
xnor U33387 (N_33387,N_27751,N_29043);
or U33388 (N_33388,N_28204,N_29939);
xnor U33389 (N_33389,N_27903,N_29862);
or U33390 (N_33390,N_26420,N_29029);
nor U33391 (N_33391,N_28345,N_27258);
and U33392 (N_33392,N_27432,N_25278);
nand U33393 (N_33393,N_28481,N_27009);
and U33394 (N_33394,N_25503,N_28598);
nor U33395 (N_33395,N_29661,N_27924);
and U33396 (N_33396,N_27755,N_28528);
or U33397 (N_33397,N_29589,N_28893);
or U33398 (N_33398,N_27815,N_26085);
xnor U33399 (N_33399,N_25672,N_25371);
or U33400 (N_33400,N_27912,N_29358);
or U33401 (N_33401,N_27486,N_26722);
nand U33402 (N_33402,N_28932,N_27216);
xnor U33403 (N_33403,N_27304,N_29565);
nand U33404 (N_33404,N_29385,N_29106);
nand U33405 (N_33405,N_28915,N_29953);
or U33406 (N_33406,N_28846,N_27900);
or U33407 (N_33407,N_28656,N_26736);
and U33408 (N_33408,N_26929,N_25392);
and U33409 (N_33409,N_26789,N_29795);
or U33410 (N_33410,N_26618,N_28315);
xnor U33411 (N_33411,N_28504,N_27173);
and U33412 (N_33412,N_29945,N_28322);
nand U33413 (N_33413,N_29327,N_28099);
nor U33414 (N_33414,N_29205,N_27985);
or U33415 (N_33415,N_25370,N_26705);
nand U33416 (N_33416,N_25945,N_27445);
nor U33417 (N_33417,N_28690,N_28411);
xnor U33418 (N_33418,N_28991,N_28874);
xor U33419 (N_33419,N_28156,N_26587);
nand U33420 (N_33420,N_28599,N_27756);
and U33421 (N_33421,N_25480,N_29663);
and U33422 (N_33422,N_26918,N_26225);
nand U33423 (N_33423,N_25910,N_29805);
and U33424 (N_33424,N_29103,N_27618);
xor U33425 (N_33425,N_29642,N_25258);
xnor U33426 (N_33426,N_29592,N_26533);
or U33427 (N_33427,N_28535,N_28735);
and U33428 (N_33428,N_28405,N_29810);
and U33429 (N_33429,N_29627,N_25505);
nand U33430 (N_33430,N_29018,N_27171);
and U33431 (N_33431,N_27539,N_26596);
nand U33432 (N_33432,N_26246,N_29563);
xnor U33433 (N_33433,N_25903,N_27257);
and U33434 (N_33434,N_26923,N_26863);
nor U33435 (N_33435,N_27692,N_28803);
xor U33436 (N_33436,N_25953,N_26594);
nand U33437 (N_33437,N_25442,N_25739);
xnor U33438 (N_33438,N_27534,N_27144);
xnor U33439 (N_33439,N_28219,N_26374);
nand U33440 (N_33440,N_28506,N_29781);
nand U33441 (N_33441,N_28160,N_29429);
xnor U33442 (N_33442,N_28396,N_29338);
and U33443 (N_33443,N_28010,N_29406);
and U33444 (N_33444,N_25940,N_25983);
nand U33445 (N_33445,N_26659,N_29044);
nand U33446 (N_33446,N_25372,N_29998);
nor U33447 (N_33447,N_25458,N_29486);
or U33448 (N_33448,N_29449,N_26612);
nor U33449 (N_33449,N_25253,N_25697);
nor U33450 (N_33450,N_27567,N_29956);
xnor U33451 (N_33451,N_26895,N_28634);
nand U33452 (N_33452,N_27847,N_27624);
nand U33453 (N_33453,N_26617,N_26999);
nand U33454 (N_33454,N_29463,N_29356);
or U33455 (N_33455,N_25734,N_29620);
nand U33456 (N_33456,N_26625,N_25800);
nor U33457 (N_33457,N_26949,N_25663);
nor U33458 (N_33458,N_28229,N_26984);
nor U33459 (N_33459,N_29597,N_28722);
or U33460 (N_33460,N_26853,N_26340);
and U33461 (N_33461,N_25762,N_25587);
nor U33462 (N_33462,N_25217,N_28047);
nor U33463 (N_33463,N_26638,N_29972);
or U33464 (N_33464,N_25698,N_25221);
or U33465 (N_33465,N_28899,N_29098);
nor U33466 (N_33466,N_25580,N_26974);
or U33467 (N_33467,N_28106,N_29557);
xnor U33468 (N_33468,N_28104,N_27614);
nor U33469 (N_33469,N_26299,N_27541);
and U33470 (N_33470,N_27766,N_29146);
or U33471 (N_33471,N_26488,N_26779);
or U33472 (N_33472,N_29010,N_28236);
nand U33473 (N_33473,N_25375,N_25903);
nand U33474 (N_33474,N_29506,N_25352);
xor U33475 (N_33475,N_29251,N_25966);
and U33476 (N_33476,N_29136,N_25381);
nand U33477 (N_33477,N_28681,N_29440);
nor U33478 (N_33478,N_29120,N_25661);
xnor U33479 (N_33479,N_27700,N_25662);
nor U33480 (N_33480,N_27319,N_28650);
nand U33481 (N_33481,N_27192,N_26523);
or U33482 (N_33482,N_26619,N_25417);
or U33483 (N_33483,N_29231,N_28348);
and U33484 (N_33484,N_28075,N_27719);
and U33485 (N_33485,N_26205,N_26891);
and U33486 (N_33486,N_28992,N_26133);
or U33487 (N_33487,N_29477,N_29534);
xnor U33488 (N_33488,N_28979,N_25538);
and U33489 (N_33489,N_25780,N_27661);
nand U33490 (N_33490,N_27768,N_27712);
and U33491 (N_33491,N_26869,N_28475);
nand U33492 (N_33492,N_25787,N_28890);
and U33493 (N_33493,N_28582,N_29565);
xnor U33494 (N_33494,N_27821,N_27127);
or U33495 (N_33495,N_26528,N_27877);
or U33496 (N_33496,N_28150,N_26485);
nand U33497 (N_33497,N_25925,N_28430);
and U33498 (N_33498,N_29757,N_26346);
nor U33499 (N_33499,N_28405,N_25998);
nand U33500 (N_33500,N_25948,N_28512);
or U33501 (N_33501,N_25418,N_29145);
nand U33502 (N_33502,N_28830,N_25241);
and U33503 (N_33503,N_27675,N_29581);
nor U33504 (N_33504,N_27687,N_26960);
and U33505 (N_33505,N_28847,N_25187);
nand U33506 (N_33506,N_29330,N_28666);
nand U33507 (N_33507,N_29555,N_27099);
and U33508 (N_33508,N_28523,N_28018);
or U33509 (N_33509,N_27136,N_28517);
xor U33510 (N_33510,N_29573,N_25581);
or U33511 (N_33511,N_29203,N_27224);
and U33512 (N_33512,N_29101,N_28949);
nand U33513 (N_33513,N_28032,N_26357);
xnor U33514 (N_33514,N_27099,N_29491);
and U33515 (N_33515,N_25041,N_26813);
xor U33516 (N_33516,N_26909,N_27719);
or U33517 (N_33517,N_26449,N_25326);
nor U33518 (N_33518,N_25807,N_28838);
xor U33519 (N_33519,N_26660,N_25780);
nand U33520 (N_33520,N_27240,N_25113);
xnor U33521 (N_33521,N_29757,N_29377);
xor U33522 (N_33522,N_25026,N_26192);
nand U33523 (N_33523,N_26354,N_28192);
nand U33524 (N_33524,N_25076,N_28286);
xnor U33525 (N_33525,N_27864,N_27214);
nand U33526 (N_33526,N_26016,N_25078);
nor U33527 (N_33527,N_27692,N_27202);
xnor U33528 (N_33528,N_28572,N_29218);
and U33529 (N_33529,N_28370,N_25606);
and U33530 (N_33530,N_26788,N_25596);
or U33531 (N_33531,N_26372,N_25914);
nand U33532 (N_33532,N_26029,N_27948);
xor U33533 (N_33533,N_28583,N_28043);
nor U33534 (N_33534,N_26661,N_28722);
or U33535 (N_33535,N_28470,N_25439);
and U33536 (N_33536,N_27991,N_29456);
and U33537 (N_33537,N_26363,N_26896);
xnor U33538 (N_33538,N_27866,N_25754);
nor U33539 (N_33539,N_29244,N_26057);
xor U33540 (N_33540,N_28971,N_26791);
nand U33541 (N_33541,N_25240,N_27974);
nor U33542 (N_33542,N_25223,N_25545);
and U33543 (N_33543,N_27736,N_29763);
xnor U33544 (N_33544,N_27534,N_27860);
nand U33545 (N_33545,N_27304,N_28232);
or U33546 (N_33546,N_28231,N_25507);
nor U33547 (N_33547,N_27176,N_28339);
xnor U33548 (N_33548,N_28861,N_29702);
or U33549 (N_33549,N_27780,N_27969);
nor U33550 (N_33550,N_28689,N_29085);
and U33551 (N_33551,N_26293,N_28681);
or U33552 (N_33552,N_29962,N_27555);
nor U33553 (N_33553,N_25883,N_29962);
xnor U33554 (N_33554,N_26668,N_27816);
xnor U33555 (N_33555,N_29606,N_25604);
nand U33556 (N_33556,N_29045,N_26850);
or U33557 (N_33557,N_27763,N_26899);
nand U33558 (N_33558,N_27483,N_28419);
or U33559 (N_33559,N_28163,N_26183);
nor U33560 (N_33560,N_29806,N_28479);
and U33561 (N_33561,N_26939,N_29457);
or U33562 (N_33562,N_28523,N_29637);
nand U33563 (N_33563,N_28454,N_26507);
nand U33564 (N_33564,N_28737,N_25377);
and U33565 (N_33565,N_27747,N_26819);
nand U33566 (N_33566,N_29922,N_28381);
nand U33567 (N_33567,N_26080,N_27462);
or U33568 (N_33568,N_25409,N_29609);
nand U33569 (N_33569,N_26680,N_29395);
and U33570 (N_33570,N_26364,N_26244);
xnor U33571 (N_33571,N_25237,N_25032);
xor U33572 (N_33572,N_28309,N_26222);
nor U33573 (N_33573,N_28529,N_27580);
xor U33574 (N_33574,N_29260,N_28511);
nand U33575 (N_33575,N_28262,N_27261);
nand U33576 (N_33576,N_26437,N_28107);
xor U33577 (N_33577,N_27830,N_29891);
or U33578 (N_33578,N_25795,N_26442);
nand U33579 (N_33579,N_29019,N_26603);
or U33580 (N_33580,N_28992,N_29619);
and U33581 (N_33581,N_26163,N_25643);
and U33582 (N_33582,N_29998,N_28813);
nand U33583 (N_33583,N_27424,N_26266);
nand U33584 (N_33584,N_29005,N_28799);
nor U33585 (N_33585,N_25312,N_27759);
or U33586 (N_33586,N_26000,N_26145);
nor U33587 (N_33587,N_25129,N_25135);
nor U33588 (N_33588,N_27007,N_26221);
or U33589 (N_33589,N_29350,N_29787);
nand U33590 (N_33590,N_25638,N_27450);
nand U33591 (N_33591,N_27876,N_27030);
xor U33592 (N_33592,N_28554,N_27059);
or U33593 (N_33593,N_26677,N_28403);
xor U33594 (N_33594,N_29738,N_25020);
nand U33595 (N_33595,N_25058,N_26990);
nor U33596 (N_33596,N_28698,N_27221);
and U33597 (N_33597,N_28164,N_29637);
and U33598 (N_33598,N_29226,N_25958);
nand U33599 (N_33599,N_27593,N_26312);
or U33600 (N_33600,N_25240,N_27770);
or U33601 (N_33601,N_29658,N_27766);
xnor U33602 (N_33602,N_27414,N_25091);
and U33603 (N_33603,N_28520,N_29007);
and U33604 (N_33604,N_26403,N_25761);
nor U33605 (N_33605,N_25051,N_29722);
xor U33606 (N_33606,N_26725,N_28723);
nor U33607 (N_33607,N_25059,N_29042);
and U33608 (N_33608,N_28835,N_25283);
and U33609 (N_33609,N_26513,N_26287);
nand U33610 (N_33610,N_29294,N_28451);
or U33611 (N_33611,N_28989,N_27550);
or U33612 (N_33612,N_26338,N_26752);
nand U33613 (N_33613,N_26558,N_25350);
nor U33614 (N_33614,N_26271,N_26331);
and U33615 (N_33615,N_28800,N_28703);
nand U33616 (N_33616,N_27246,N_29500);
or U33617 (N_33617,N_27225,N_28190);
xor U33618 (N_33618,N_26314,N_25504);
or U33619 (N_33619,N_26263,N_26628);
nand U33620 (N_33620,N_28785,N_25302);
xnor U33621 (N_33621,N_29899,N_27667);
nand U33622 (N_33622,N_26002,N_29687);
and U33623 (N_33623,N_26655,N_26423);
xnor U33624 (N_33624,N_26951,N_26345);
xnor U33625 (N_33625,N_26391,N_26141);
and U33626 (N_33626,N_26991,N_27227);
nand U33627 (N_33627,N_29283,N_25205);
and U33628 (N_33628,N_25967,N_28993);
or U33629 (N_33629,N_26310,N_26450);
xor U33630 (N_33630,N_27233,N_28389);
or U33631 (N_33631,N_29188,N_25321);
nand U33632 (N_33632,N_25345,N_26726);
nand U33633 (N_33633,N_25009,N_27200);
and U33634 (N_33634,N_29966,N_25440);
nor U33635 (N_33635,N_26173,N_28037);
xnor U33636 (N_33636,N_25879,N_25831);
nand U33637 (N_33637,N_27814,N_25203);
nand U33638 (N_33638,N_29994,N_25355);
xnor U33639 (N_33639,N_28234,N_28472);
nand U33640 (N_33640,N_27006,N_28509);
and U33641 (N_33641,N_28300,N_25743);
and U33642 (N_33642,N_29090,N_29348);
or U33643 (N_33643,N_25881,N_26546);
xnor U33644 (N_33644,N_27453,N_28965);
nor U33645 (N_33645,N_29804,N_26329);
nor U33646 (N_33646,N_29425,N_26636);
xor U33647 (N_33647,N_25226,N_26871);
and U33648 (N_33648,N_25992,N_29849);
and U33649 (N_33649,N_26944,N_29367);
and U33650 (N_33650,N_25703,N_25370);
xnor U33651 (N_33651,N_28008,N_29320);
and U33652 (N_33652,N_26051,N_25500);
xor U33653 (N_33653,N_28644,N_28789);
nand U33654 (N_33654,N_27081,N_29916);
nand U33655 (N_33655,N_27130,N_29239);
or U33656 (N_33656,N_29073,N_25006);
nor U33657 (N_33657,N_27693,N_26214);
nand U33658 (N_33658,N_26773,N_27178);
and U33659 (N_33659,N_25958,N_28340);
nor U33660 (N_33660,N_27248,N_25612);
xor U33661 (N_33661,N_25435,N_27537);
nand U33662 (N_33662,N_28141,N_28761);
and U33663 (N_33663,N_25837,N_27056);
or U33664 (N_33664,N_27889,N_27964);
nor U33665 (N_33665,N_29918,N_28595);
nand U33666 (N_33666,N_28601,N_27847);
nand U33667 (N_33667,N_29653,N_25271);
and U33668 (N_33668,N_29139,N_28705);
and U33669 (N_33669,N_27477,N_28998);
or U33670 (N_33670,N_29618,N_25550);
or U33671 (N_33671,N_29888,N_27904);
xnor U33672 (N_33672,N_26651,N_28525);
xor U33673 (N_33673,N_26083,N_28410);
nand U33674 (N_33674,N_25139,N_28392);
nand U33675 (N_33675,N_28289,N_26032);
or U33676 (N_33676,N_28627,N_25316);
nand U33677 (N_33677,N_28917,N_25028);
nand U33678 (N_33678,N_26179,N_28161);
or U33679 (N_33679,N_27489,N_27868);
and U33680 (N_33680,N_27692,N_27493);
and U33681 (N_33681,N_28795,N_27842);
and U33682 (N_33682,N_25344,N_28946);
nand U33683 (N_33683,N_25283,N_27987);
nand U33684 (N_33684,N_28047,N_25029);
xnor U33685 (N_33685,N_29577,N_27973);
nor U33686 (N_33686,N_25992,N_25815);
or U33687 (N_33687,N_28371,N_27394);
nor U33688 (N_33688,N_29232,N_26462);
xnor U33689 (N_33689,N_29433,N_27965);
or U33690 (N_33690,N_29847,N_28627);
and U33691 (N_33691,N_27390,N_25427);
or U33692 (N_33692,N_25153,N_27897);
xnor U33693 (N_33693,N_25807,N_28348);
and U33694 (N_33694,N_26634,N_26709);
and U33695 (N_33695,N_25501,N_25317);
and U33696 (N_33696,N_29091,N_25378);
and U33697 (N_33697,N_25064,N_29853);
and U33698 (N_33698,N_27894,N_28501);
or U33699 (N_33699,N_28808,N_28382);
nand U33700 (N_33700,N_25706,N_25790);
and U33701 (N_33701,N_29132,N_27802);
nand U33702 (N_33702,N_29331,N_26028);
or U33703 (N_33703,N_26929,N_29132);
xnor U33704 (N_33704,N_26862,N_27486);
nor U33705 (N_33705,N_26722,N_25119);
nand U33706 (N_33706,N_26326,N_25874);
and U33707 (N_33707,N_27589,N_26733);
nand U33708 (N_33708,N_25712,N_28189);
nand U33709 (N_33709,N_28602,N_27967);
or U33710 (N_33710,N_26643,N_29923);
nor U33711 (N_33711,N_29610,N_26351);
nor U33712 (N_33712,N_26581,N_25794);
nor U33713 (N_33713,N_25341,N_25390);
or U33714 (N_33714,N_25394,N_29063);
and U33715 (N_33715,N_25398,N_28140);
nand U33716 (N_33716,N_27863,N_25243);
xnor U33717 (N_33717,N_28397,N_25276);
and U33718 (N_33718,N_29525,N_27495);
or U33719 (N_33719,N_26862,N_26206);
nor U33720 (N_33720,N_27299,N_29051);
nor U33721 (N_33721,N_25010,N_26429);
xor U33722 (N_33722,N_27374,N_29645);
and U33723 (N_33723,N_27953,N_25200);
nor U33724 (N_33724,N_26929,N_26361);
xnor U33725 (N_33725,N_29162,N_25511);
nand U33726 (N_33726,N_27814,N_29684);
or U33727 (N_33727,N_25485,N_28954);
nor U33728 (N_33728,N_28586,N_28620);
nand U33729 (N_33729,N_26012,N_25769);
xor U33730 (N_33730,N_26578,N_26067);
and U33731 (N_33731,N_29518,N_28355);
nand U33732 (N_33732,N_26019,N_26513);
xnor U33733 (N_33733,N_25271,N_27714);
or U33734 (N_33734,N_25263,N_26755);
or U33735 (N_33735,N_25316,N_26765);
or U33736 (N_33736,N_27485,N_26461);
nor U33737 (N_33737,N_26857,N_28924);
or U33738 (N_33738,N_26670,N_25829);
nor U33739 (N_33739,N_26323,N_29110);
nor U33740 (N_33740,N_27115,N_26241);
or U33741 (N_33741,N_26281,N_25327);
nand U33742 (N_33742,N_26613,N_25156);
xor U33743 (N_33743,N_26482,N_29075);
xnor U33744 (N_33744,N_28551,N_28393);
xor U33745 (N_33745,N_28889,N_29089);
and U33746 (N_33746,N_29583,N_29050);
xor U33747 (N_33747,N_26563,N_28053);
xnor U33748 (N_33748,N_25054,N_28150);
or U33749 (N_33749,N_29747,N_28105);
xnor U33750 (N_33750,N_25588,N_29399);
nand U33751 (N_33751,N_27168,N_25028);
nor U33752 (N_33752,N_28875,N_28540);
xnor U33753 (N_33753,N_25559,N_27701);
and U33754 (N_33754,N_27074,N_27101);
or U33755 (N_33755,N_28754,N_28486);
and U33756 (N_33756,N_27541,N_25783);
nor U33757 (N_33757,N_25343,N_27140);
or U33758 (N_33758,N_26854,N_28652);
nor U33759 (N_33759,N_29943,N_27307);
nor U33760 (N_33760,N_29290,N_26301);
and U33761 (N_33761,N_29354,N_26444);
or U33762 (N_33762,N_25260,N_27234);
xnor U33763 (N_33763,N_29794,N_25470);
nand U33764 (N_33764,N_27248,N_25090);
xnor U33765 (N_33765,N_28195,N_29095);
nand U33766 (N_33766,N_25072,N_28571);
nor U33767 (N_33767,N_27044,N_28296);
or U33768 (N_33768,N_25675,N_25926);
nor U33769 (N_33769,N_29363,N_25231);
xor U33770 (N_33770,N_26084,N_25718);
or U33771 (N_33771,N_28123,N_27102);
or U33772 (N_33772,N_28645,N_25442);
and U33773 (N_33773,N_28779,N_27582);
nor U33774 (N_33774,N_25169,N_27787);
nor U33775 (N_33775,N_29467,N_28051);
nand U33776 (N_33776,N_26278,N_29590);
nand U33777 (N_33777,N_26929,N_29656);
nor U33778 (N_33778,N_28869,N_27202);
xor U33779 (N_33779,N_26884,N_28256);
and U33780 (N_33780,N_25311,N_29691);
and U33781 (N_33781,N_29525,N_26100);
xnor U33782 (N_33782,N_29582,N_26570);
or U33783 (N_33783,N_25999,N_27748);
xnor U33784 (N_33784,N_27654,N_27502);
xnor U33785 (N_33785,N_27086,N_28046);
or U33786 (N_33786,N_27301,N_29363);
or U33787 (N_33787,N_28185,N_28786);
nor U33788 (N_33788,N_28155,N_26388);
and U33789 (N_33789,N_25418,N_28735);
nand U33790 (N_33790,N_27135,N_25657);
or U33791 (N_33791,N_26754,N_29121);
nand U33792 (N_33792,N_28587,N_29594);
and U33793 (N_33793,N_29871,N_25165);
or U33794 (N_33794,N_27591,N_26373);
nor U33795 (N_33795,N_28076,N_27552);
xor U33796 (N_33796,N_29691,N_27452);
nor U33797 (N_33797,N_27601,N_29566);
and U33798 (N_33798,N_28429,N_25215);
nand U33799 (N_33799,N_27950,N_25805);
nand U33800 (N_33800,N_26315,N_29048);
or U33801 (N_33801,N_26777,N_27557);
xor U33802 (N_33802,N_27359,N_28110);
or U33803 (N_33803,N_28088,N_26458);
nand U33804 (N_33804,N_26474,N_25400);
nand U33805 (N_33805,N_25845,N_25611);
nand U33806 (N_33806,N_28715,N_28531);
nor U33807 (N_33807,N_29446,N_28754);
or U33808 (N_33808,N_25184,N_27809);
nor U33809 (N_33809,N_28110,N_29409);
or U33810 (N_33810,N_26526,N_28859);
and U33811 (N_33811,N_29746,N_26916);
and U33812 (N_33812,N_25582,N_26978);
nor U33813 (N_33813,N_28834,N_26496);
nor U33814 (N_33814,N_29018,N_27085);
nand U33815 (N_33815,N_28935,N_26684);
or U33816 (N_33816,N_25552,N_28029);
nor U33817 (N_33817,N_29198,N_25086);
and U33818 (N_33818,N_25900,N_29846);
and U33819 (N_33819,N_28249,N_29491);
nand U33820 (N_33820,N_25210,N_28442);
nand U33821 (N_33821,N_28729,N_27864);
nor U33822 (N_33822,N_25521,N_27254);
and U33823 (N_33823,N_26331,N_25917);
nand U33824 (N_33824,N_27115,N_28929);
or U33825 (N_33825,N_25651,N_28959);
nor U33826 (N_33826,N_28007,N_28459);
nor U33827 (N_33827,N_27062,N_27513);
nor U33828 (N_33828,N_27212,N_27975);
xnor U33829 (N_33829,N_27406,N_27591);
or U33830 (N_33830,N_28851,N_27017);
nand U33831 (N_33831,N_25786,N_26314);
nand U33832 (N_33832,N_27917,N_27981);
and U33833 (N_33833,N_26965,N_29956);
or U33834 (N_33834,N_27734,N_25659);
xnor U33835 (N_33835,N_29749,N_25477);
nand U33836 (N_33836,N_29471,N_27382);
and U33837 (N_33837,N_27556,N_28239);
nor U33838 (N_33838,N_26448,N_27182);
nor U33839 (N_33839,N_26952,N_28151);
nor U33840 (N_33840,N_28302,N_27702);
xnor U33841 (N_33841,N_26246,N_25851);
or U33842 (N_33842,N_25615,N_25296);
and U33843 (N_33843,N_29290,N_25087);
nand U33844 (N_33844,N_25264,N_25899);
and U33845 (N_33845,N_28244,N_26425);
xnor U33846 (N_33846,N_27930,N_29034);
xor U33847 (N_33847,N_28149,N_25247);
xnor U33848 (N_33848,N_26201,N_27468);
xnor U33849 (N_33849,N_25824,N_25859);
nor U33850 (N_33850,N_27693,N_28215);
xnor U33851 (N_33851,N_29913,N_26306);
nand U33852 (N_33852,N_27416,N_25737);
nor U33853 (N_33853,N_25749,N_25266);
nand U33854 (N_33854,N_28859,N_28764);
xor U33855 (N_33855,N_26593,N_26851);
nor U33856 (N_33856,N_29971,N_29825);
xnor U33857 (N_33857,N_29056,N_27477);
nand U33858 (N_33858,N_25253,N_26658);
and U33859 (N_33859,N_27306,N_28093);
nand U33860 (N_33860,N_26471,N_26210);
xor U33861 (N_33861,N_28786,N_29418);
nand U33862 (N_33862,N_27930,N_29063);
nor U33863 (N_33863,N_26489,N_27201);
or U33864 (N_33864,N_25267,N_25447);
nor U33865 (N_33865,N_27096,N_27505);
nor U33866 (N_33866,N_25025,N_25014);
nor U33867 (N_33867,N_27725,N_27879);
or U33868 (N_33868,N_28377,N_28202);
and U33869 (N_33869,N_29314,N_28195);
or U33870 (N_33870,N_27755,N_25937);
nand U33871 (N_33871,N_25901,N_28362);
or U33872 (N_33872,N_25931,N_26801);
nand U33873 (N_33873,N_29503,N_27546);
xnor U33874 (N_33874,N_25904,N_29994);
and U33875 (N_33875,N_28147,N_25198);
or U33876 (N_33876,N_28017,N_25456);
xnor U33877 (N_33877,N_29193,N_28262);
or U33878 (N_33878,N_29650,N_29892);
and U33879 (N_33879,N_26147,N_27497);
or U33880 (N_33880,N_29850,N_27237);
or U33881 (N_33881,N_29875,N_27771);
nor U33882 (N_33882,N_27353,N_27771);
nor U33883 (N_33883,N_26292,N_28015);
xnor U33884 (N_33884,N_29115,N_27684);
nand U33885 (N_33885,N_29659,N_26009);
nor U33886 (N_33886,N_25913,N_28630);
or U33887 (N_33887,N_27074,N_27024);
or U33888 (N_33888,N_25400,N_29718);
nor U33889 (N_33889,N_25451,N_28961);
or U33890 (N_33890,N_28139,N_25823);
nand U33891 (N_33891,N_28660,N_29789);
xnor U33892 (N_33892,N_27498,N_28964);
and U33893 (N_33893,N_26331,N_27582);
and U33894 (N_33894,N_29806,N_29589);
xor U33895 (N_33895,N_25478,N_28143);
nand U33896 (N_33896,N_27790,N_28801);
and U33897 (N_33897,N_28191,N_25130);
xor U33898 (N_33898,N_27658,N_25624);
nor U33899 (N_33899,N_29507,N_27470);
and U33900 (N_33900,N_27105,N_29081);
xnor U33901 (N_33901,N_27780,N_25502);
nand U33902 (N_33902,N_27379,N_26725);
nor U33903 (N_33903,N_29939,N_27918);
and U33904 (N_33904,N_27858,N_29075);
and U33905 (N_33905,N_28335,N_29002);
xor U33906 (N_33906,N_27383,N_28229);
or U33907 (N_33907,N_29253,N_25553);
and U33908 (N_33908,N_25359,N_25863);
and U33909 (N_33909,N_26307,N_28770);
or U33910 (N_33910,N_28323,N_29501);
xnor U33911 (N_33911,N_27541,N_29989);
nand U33912 (N_33912,N_26208,N_28154);
xnor U33913 (N_33913,N_28845,N_29039);
and U33914 (N_33914,N_27872,N_25734);
xor U33915 (N_33915,N_27741,N_29322);
xor U33916 (N_33916,N_26943,N_27472);
xnor U33917 (N_33917,N_26195,N_25151);
or U33918 (N_33918,N_27205,N_25358);
and U33919 (N_33919,N_26719,N_26660);
nor U33920 (N_33920,N_27195,N_25800);
nor U33921 (N_33921,N_27025,N_26461);
and U33922 (N_33922,N_28078,N_25116);
xnor U33923 (N_33923,N_28179,N_27511);
nor U33924 (N_33924,N_28824,N_28298);
xor U33925 (N_33925,N_27819,N_25429);
xor U33926 (N_33926,N_28093,N_27328);
nor U33927 (N_33927,N_25412,N_27631);
nand U33928 (N_33928,N_26949,N_29315);
or U33929 (N_33929,N_29279,N_27053);
xor U33930 (N_33930,N_28444,N_25370);
or U33931 (N_33931,N_25056,N_27150);
and U33932 (N_33932,N_29201,N_29326);
and U33933 (N_33933,N_27826,N_25693);
or U33934 (N_33934,N_25579,N_28770);
nor U33935 (N_33935,N_26277,N_27196);
nand U33936 (N_33936,N_26285,N_28819);
and U33937 (N_33937,N_25280,N_26987);
or U33938 (N_33938,N_25601,N_25392);
xnor U33939 (N_33939,N_29059,N_29968);
nor U33940 (N_33940,N_27996,N_29710);
or U33941 (N_33941,N_29369,N_26960);
nor U33942 (N_33942,N_26119,N_29403);
nand U33943 (N_33943,N_27245,N_25699);
and U33944 (N_33944,N_25255,N_29517);
or U33945 (N_33945,N_25933,N_25282);
nor U33946 (N_33946,N_26209,N_26947);
nor U33947 (N_33947,N_25947,N_25238);
nand U33948 (N_33948,N_29612,N_26369);
nor U33949 (N_33949,N_26604,N_26089);
nand U33950 (N_33950,N_29814,N_29895);
and U33951 (N_33951,N_26119,N_25398);
nor U33952 (N_33952,N_28584,N_29521);
nor U33953 (N_33953,N_28720,N_27300);
and U33954 (N_33954,N_25255,N_26293);
and U33955 (N_33955,N_26156,N_27303);
nand U33956 (N_33956,N_26143,N_29783);
nand U33957 (N_33957,N_28953,N_26524);
and U33958 (N_33958,N_27159,N_28837);
nor U33959 (N_33959,N_29955,N_29720);
nand U33960 (N_33960,N_27169,N_26815);
nand U33961 (N_33961,N_29709,N_25296);
xor U33962 (N_33962,N_28561,N_28528);
xnor U33963 (N_33963,N_26725,N_27485);
or U33964 (N_33964,N_25944,N_28532);
nand U33965 (N_33965,N_28567,N_27766);
nand U33966 (N_33966,N_26543,N_25611);
and U33967 (N_33967,N_29142,N_28721);
nand U33968 (N_33968,N_26066,N_27439);
nand U33969 (N_33969,N_28437,N_25048);
xor U33970 (N_33970,N_26323,N_25174);
nor U33971 (N_33971,N_26654,N_29369);
xor U33972 (N_33972,N_25249,N_25683);
nor U33973 (N_33973,N_25379,N_25394);
nand U33974 (N_33974,N_27915,N_26330);
and U33975 (N_33975,N_28620,N_28274);
and U33976 (N_33976,N_25302,N_26713);
nor U33977 (N_33977,N_27348,N_25072);
and U33978 (N_33978,N_25125,N_27690);
or U33979 (N_33979,N_28152,N_29746);
nand U33980 (N_33980,N_27589,N_28291);
nand U33981 (N_33981,N_25497,N_26789);
or U33982 (N_33982,N_25486,N_27084);
and U33983 (N_33983,N_25503,N_29298);
xor U33984 (N_33984,N_27558,N_26323);
xnor U33985 (N_33985,N_26187,N_27654);
xnor U33986 (N_33986,N_29955,N_26561);
nor U33987 (N_33987,N_26031,N_27040);
nor U33988 (N_33988,N_27975,N_29387);
xnor U33989 (N_33989,N_28141,N_28398);
and U33990 (N_33990,N_29882,N_26970);
nand U33991 (N_33991,N_26728,N_26018);
xor U33992 (N_33992,N_29263,N_26435);
and U33993 (N_33993,N_25445,N_29444);
and U33994 (N_33994,N_25374,N_25187);
nor U33995 (N_33995,N_25816,N_27313);
nor U33996 (N_33996,N_25321,N_26872);
nand U33997 (N_33997,N_27826,N_27187);
xor U33998 (N_33998,N_25333,N_26940);
and U33999 (N_33999,N_25313,N_27417);
nand U34000 (N_34000,N_27355,N_26435);
xor U34001 (N_34001,N_27128,N_27451);
nor U34002 (N_34002,N_28868,N_27620);
xor U34003 (N_34003,N_28295,N_29498);
or U34004 (N_34004,N_25731,N_27622);
nor U34005 (N_34005,N_27809,N_25183);
nor U34006 (N_34006,N_27209,N_28986);
or U34007 (N_34007,N_29229,N_26179);
nor U34008 (N_34008,N_27874,N_26391);
nand U34009 (N_34009,N_28503,N_26585);
xor U34010 (N_34010,N_29110,N_28843);
xor U34011 (N_34011,N_25022,N_27793);
and U34012 (N_34012,N_27555,N_29109);
nor U34013 (N_34013,N_26983,N_27362);
and U34014 (N_34014,N_27945,N_26784);
nand U34015 (N_34015,N_26381,N_27896);
and U34016 (N_34016,N_28658,N_25670);
nor U34017 (N_34017,N_29035,N_25465);
xnor U34018 (N_34018,N_27793,N_27508);
nor U34019 (N_34019,N_25259,N_29337);
or U34020 (N_34020,N_29886,N_25832);
and U34021 (N_34021,N_27091,N_26570);
nor U34022 (N_34022,N_29439,N_26623);
or U34023 (N_34023,N_25501,N_25157);
xnor U34024 (N_34024,N_29924,N_27747);
xor U34025 (N_34025,N_29705,N_29629);
nor U34026 (N_34026,N_25965,N_27088);
nor U34027 (N_34027,N_28163,N_28287);
nand U34028 (N_34028,N_27840,N_26024);
nor U34029 (N_34029,N_27643,N_28091);
xnor U34030 (N_34030,N_29513,N_25485);
nor U34031 (N_34031,N_29090,N_25359);
xnor U34032 (N_34032,N_26760,N_26618);
or U34033 (N_34033,N_29887,N_28519);
and U34034 (N_34034,N_25537,N_26591);
xnor U34035 (N_34035,N_28954,N_25975);
nand U34036 (N_34036,N_28504,N_27044);
or U34037 (N_34037,N_29189,N_27129);
or U34038 (N_34038,N_27983,N_25303);
xor U34039 (N_34039,N_26472,N_28339);
nand U34040 (N_34040,N_26982,N_27564);
and U34041 (N_34041,N_26287,N_28937);
xor U34042 (N_34042,N_27646,N_28704);
or U34043 (N_34043,N_29630,N_25928);
nand U34044 (N_34044,N_25603,N_28240);
nor U34045 (N_34045,N_29815,N_26283);
nand U34046 (N_34046,N_27075,N_26128);
nand U34047 (N_34047,N_25361,N_25878);
or U34048 (N_34048,N_29135,N_29252);
xor U34049 (N_34049,N_27663,N_26456);
and U34050 (N_34050,N_29747,N_26598);
and U34051 (N_34051,N_26483,N_27417);
nand U34052 (N_34052,N_25037,N_28634);
or U34053 (N_34053,N_25870,N_25860);
nor U34054 (N_34054,N_26190,N_29128);
xnor U34055 (N_34055,N_29566,N_26880);
and U34056 (N_34056,N_29501,N_25252);
nand U34057 (N_34057,N_26592,N_29539);
xor U34058 (N_34058,N_28417,N_28370);
nor U34059 (N_34059,N_28752,N_25995);
or U34060 (N_34060,N_29246,N_27925);
or U34061 (N_34061,N_25437,N_26447);
and U34062 (N_34062,N_29565,N_28103);
nand U34063 (N_34063,N_26944,N_28706);
and U34064 (N_34064,N_26108,N_26958);
nand U34065 (N_34065,N_25589,N_27454);
nor U34066 (N_34066,N_29775,N_27665);
xnor U34067 (N_34067,N_29508,N_27239);
xnor U34068 (N_34068,N_26186,N_29620);
and U34069 (N_34069,N_25553,N_25065);
nor U34070 (N_34070,N_26253,N_28172);
and U34071 (N_34071,N_26362,N_29185);
and U34072 (N_34072,N_27582,N_28380);
nor U34073 (N_34073,N_26219,N_29515);
and U34074 (N_34074,N_25947,N_26183);
xnor U34075 (N_34075,N_25225,N_26707);
and U34076 (N_34076,N_28109,N_27194);
nand U34077 (N_34077,N_25927,N_25745);
and U34078 (N_34078,N_28947,N_25520);
xnor U34079 (N_34079,N_28095,N_27612);
nand U34080 (N_34080,N_27440,N_25271);
nor U34081 (N_34081,N_27604,N_26949);
or U34082 (N_34082,N_29475,N_28085);
and U34083 (N_34083,N_25983,N_28040);
nand U34084 (N_34084,N_25388,N_25331);
and U34085 (N_34085,N_29018,N_25016);
nand U34086 (N_34086,N_29292,N_25080);
nand U34087 (N_34087,N_27385,N_28392);
and U34088 (N_34088,N_26018,N_27600);
or U34089 (N_34089,N_26068,N_29648);
nor U34090 (N_34090,N_29547,N_25913);
and U34091 (N_34091,N_27724,N_26336);
nor U34092 (N_34092,N_29001,N_28217);
nand U34093 (N_34093,N_29544,N_28097);
xor U34094 (N_34094,N_25911,N_25584);
nor U34095 (N_34095,N_27543,N_26624);
xnor U34096 (N_34096,N_29422,N_27677);
or U34097 (N_34097,N_28336,N_26052);
nand U34098 (N_34098,N_28328,N_27342);
and U34099 (N_34099,N_28643,N_28426);
or U34100 (N_34100,N_25071,N_26631);
and U34101 (N_34101,N_27991,N_29157);
nor U34102 (N_34102,N_25099,N_25060);
nand U34103 (N_34103,N_27454,N_27657);
or U34104 (N_34104,N_28661,N_27875);
nand U34105 (N_34105,N_25878,N_25116);
nor U34106 (N_34106,N_27550,N_27148);
xor U34107 (N_34107,N_27062,N_25952);
xnor U34108 (N_34108,N_26394,N_27053);
and U34109 (N_34109,N_28096,N_27496);
or U34110 (N_34110,N_29518,N_29469);
or U34111 (N_34111,N_26669,N_29543);
xor U34112 (N_34112,N_29427,N_27118);
xnor U34113 (N_34113,N_27625,N_29527);
xnor U34114 (N_34114,N_27506,N_28887);
nand U34115 (N_34115,N_27516,N_25549);
nor U34116 (N_34116,N_28228,N_27413);
nand U34117 (N_34117,N_28320,N_26907);
nand U34118 (N_34118,N_28037,N_25038);
and U34119 (N_34119,N_28037,N_25369);
nand U34120 (N_34120,N_28784,N_25109);
or U34121 (N_34121,N_25410,N_25914);
and U34122 (N_34122,N_28130,N_27456);
nor U34123 (N_34123,N_27504,N_28060);
nor U34124 (N_34124,N_25227,N_27734);
nor U34125 (N_34125,N_28258,N_29348);
nand U34126 (N_34126,N_29466,N_29305);
nand U34127 (N_34127,N_29667,N_26657);
xor U34128 (N_34128,N_29768,N_29143);
and U34129 (N_34129,N_26130,N_29404);
and U34130 (N_34130,N_25762,N_25081);
nand U34131 (N_34131,N_25470,N_26063);
xor U34132 (N_34132,N_27654,N_29325);
xor U34133 (N_34133,N_29747,N_27096);
nor U34134 (N_34134,N_28275,N_25637);
nor U34135 (N_34135,N_27948,N_29872);
xor U34136 (N_34136,N_27345,N_28221);
nand U34137 (N_34137,N_28353,N_29247);
nor U34138 (N_34138,N_27520,N_25121);
xnor U34139 (N_34139,N_28808,N_25424);
xnor U34140 (N_34140,N_25369,N_25405);
nor U34141 (N_34141,N_27308,N_25648);
nand U34142 (N_34142,N_28412,N_25272);
xor U34143 (N_34143,N_26252,N_25190);
xnor U34144 (N_34144,N_26372,N_29690);
nand U34145 (N_34145,N_27902,N_28565);
or U34146 (N_34146,N_29855,N_25606);
xnor U34147 (N_34147,N_27168,N_29375);
xor U34148 (N_34148,N_29225,N_29136);
xnor U34149 (N_34149,N_26443,N_27344);
nor U34150 (N_34150,N_29710,N_26350);
nand U34151 (N_34151,N_25688,N_25078);
or U34152 (N_34152,N_29904,N_29284);
xnor U34153 (N_34153,N_25598,N_28903);
or U34154 (N_34154,N_26213,N_26274);
nor U34155 (N_34155,N_26316,N_28933);
xor U34156 (N_34156,N_28049,N_28273);
xnor U34157 (N_34157,N_29395,N_27129);
xnor U34158 (N_34158,N_28006,N_29546);
or U34159 (N_34159,N_28835,N_26730);
and U34160 (N_34160,N_25837,N_26785);
xnor U34161 (N_34161,N_25646,N_28252);
nor U34162 (N_34162,N_25511,N_28924);
or U34163 (N_34163,N_26420,N_25497);
xor U34164 (N_34164,N_27794,N_29055);
and U34165 (N_34165,N_27314,N_27266);
or U34166 (N_34166,N_25239,N_25336);
nor U34167 (N_34167,N_26693,N_28069);
or U34168 (N_34168,N_28948,N_25123);
or U34169 (N_34169,N_25079,N_26888);
nor U34170 (N_34170,N_26334,N_28242);
nand U34171 (N_34171,N_25739,N_25135);
and U34172 (N_34172,N_25511,N_29247);
xnor U34173 (N_34173,N_26809,N_27165);
nor U34174 (N_34174,N_25323,N_28071);
and U34175 (N_34175,N_26537,N_29521);
nor U34176 (N_34176,N_25988,N_29546);
or U34177 (N_34177,N_29481,N_27314);
or U34178 (N_34178,N_27054,N_25497);
or U34179 (N_34179,N_25438,N_28282);
or U34180 (N_34180,N_29929,N_28847);
and U34181 (N_34181,N_29326,N_25267);
xor U34182 (N_34182,N_26952,N_26132);
and U34183 (N_34183,N_29440,N_25376);
nand U34184 (N_34184,N_27165,N_25557);
xnor U34185 (N_34185,N_28977,N_27079);
or U34186 (N_34186,N_27032,N_29689);
or U34187 (N_34187,N_26349,N_26792);
and U34188 (N_34188,N_25454,N_27366);
or U34189 (N_34189,N_26661,N_29907);
xor U34190 (N_34190,N_26156,N_27742);
nand U34191 (N_34191,N_26037,N_25852);
xnor U34192 (N_34192,N_28617,N_26307);
xnor U34193 (N_34193,N_26555,N_26320);
nand U34194 (N_34194,N_25130,N_29343);
nand U34195 (N_34195,N_29044,N_27017);
nor U34196 (N_34196,N_29389,N_27946);
nand U34197 (N_34197,N_29901,N_27292);
and U34198 (N_34198,N_28189,N_28642);
xnor U34199 (N_34199,N_28375,N_27965);
nand U34200 (N_34200,N_26725,N_25179);
or U34201 (N_34201,N_29517,N_28040);
and U34202 (N_34202,N_29582,N_25660);
or U34203 (N_34203,N_27719,N_28280);
xnor U34204 (N_34204,N_28571,N_29822);
or U34205 (N_34205,N_25256,N_26088);
and U34206 (N_34206,N_27362,N_27131);
and U34207 (N_34207,N_29178,N_27378);
nand U34208 (N_34208,N_25274,N_29669);
nor U34209 (N_34209,N_26368,N_25575);
xnor U34210 (N_34210,N_26009,N_29501);
or U34211 (N_34211,N_26056,N_26639);
and U34212 (N_34212,N_27540,N_27005);
xnor U34213 (N_34213,N_29384,N_29904);
and U34214 (N_34214,N_26035,N_27658);
nand U34215 (N_34215,N_26395,N_27889);
nand U34216 (N_34216,N_26997,N_27932);
nand U34217 (N_34217,N_25771,N_29814);
nand U34218 (N_34218,N_29271,N_26885);
nor U34219 (N_34219,N_27393,N_26398);
xnor U34220 (N_34220,N_25432,N_26924);
xor U34221 (N_34221,N_29197,N_26146);
xor U34222 (N_34222,N_27835,N_28173);
nand U34223 (N_34223,N_26111,N_28835);
nand U34224 (N_34224,N_25605,N_29789);
and U34225 (N_34225,N_29813,N_27279);
xnor U34226 (N_34226,N_25474,N_27609);
and U34227 (N_34227,N_27478,N_28346);
or U34228 (N_34228,N_25860,N_28471);
nand U34229 (N_34229,N_29990,N_29039);
nand U34230 (N_34230,N_25421,N_26450);
nor U34231 (N_34231,N_25676,N_26241);
or U34232 (N_34232,N_27692,N_29722);
xor U34233 (N_34233,N_25849,N_26834);
or U34234 (N_34234,N_27332,N_27555);
or U34235 (N_34235,N_29855,N_29943);
nand U34236 (N_34236,N_27841,N_29367);
and U34237 (N_34237,N_29467,N_28611);
nor U34238 (N_34238,N_28425,N_28785);
nand U34239 (N_34239,N_26418,N_27544);
nor U34240 (N_34240,N_29672,N_26205);
xnor U34241 (N_34241,N_29550,N_29709);
xnor U34242 (N_34242,N_27627,N_26340);
nor U34243 (N_34243,N_28989,N_26009);
or U34244 (N_34244,N_29992,N_29286);
xnor U34245 (N_34245,N_26572,N_29102);
and U34246 (N_34246,N_26532,N_29897);
or U34247 (N_34247,N_27026,N_28996);
or U34248 (N_34248,N_28153,N_26288);
nor U34249 (N_34249,N_25178,N_27581);
and U34250 (N_34250,N_29657,N_27518);
nand U34251 (N_34251,N_26066,N_26129);
xnor U34252 (N_34252,N_29492,N_26868);
or U34253 (N_34253,N_29199,N_28895);
nor U34254 (N_34254,N_28045,N_26057);
nor U34255 (N_34255,N_29872,N_28215);
nor U34256 (N_34256,N_25806,N_27453);
nor U34257 (N_34257,N_27008,N_28604);
or U34258 (N_34258,N_28367,N_29128);
xor U34259 (N_34259,N_27058,N_29154);
nand U34260 (N_34260,N_25993,N_28832);
and U34261 (N_34261,N_26674,N_26356);
nand U34262 (N_34262,N_29532,N_27275);
and U34263 (N_34263,N_26534,N_27999);
xnor U34264 (N_34264,N_27786,N_28427);
nor U34265 (N_34265,N_27628,N_29467);
and U34266 (N_34266,N_27966,N_28283);
xor U34267 (N_34267,N_28940,N_25275);
nor U34268 (N_34268,N_26158,N_28063);
and U34269 (N_34269,N_27707,N_29024);
or U34270 (N_34270,N_26254,N_25327);
nand U34271 (N_34271,N_27932,N_29758);
or U34272 (N_34272,N_26629,N_29737);
and U34273 (N_34273,N_28009,N_29122);
or U34274 (N_34274,N_25294,N_27838);
nor U34275 (N_34275,N_26987,N_26779);
nor U34276 (N_34276,N_26637,N_26438);
nand U34277 (N_34277,N_26757,N_26297);
and U34278 (N_34278,N_28601,N_29460);
or U34279 (N_34279,N_27402,N_27944);
xor U34280 (N_34280,N_25034,N_29502);
nand U34281 (N_34281,N_27023,N_27795);
and U34282 (N_34282,N_26632,N_25421);
or U34283 (N_34283,N_27240,N_25441);
nand U34284 (N_34284,N_27878,N_26148);
nor U34285 (N_34285,N_29749,N_29869);
nor U34286 (N_34286,N_26183,N_28881);
xor U34287 (N_34287,N_27316,N_27503);
nor U34288 (N_34288,N_29092,N_27495);
xnor U34289 (N_34289,N_29712,N_26468);
and U34290 (N_34290,N_26678,N_25493);
nand U34291 (N_34291,N_28338,N_27761);
nor U34292 (N_34292,N_27006,N_27592);
nor U34293 (N_34293,N_25524,N_25142);
nor U34294 (N_34294,N_29514,N_26362);
and U34295 (N_34295,N_26157,N_25179);
xor U34296 (N_34296,N_27068,N_29653);
nor U34297 (N_34297,N_29805,N_25202);
and U34298 (N_34298,N_29123,N_28574);
nand U34299 (N_34299,N_25166,N_25941);
nor U34300 (N_34300,N_27891,N_28508);
and U34301 (N_34301,N_25732,N_27795);
nor U34302 (N_34302,N_25610,N_28286);
or U34303 (N_34303,N_26139,N_25597);
nand U34304 (N_34304,N_27778,N_29069);
nand U34305 (N_34305,N_29665,N_29884);
nor U34306 (N_34306,N_25109,N_25173);
or U34307 (N_34307,N_25214,N_27524);
nor U34308 (N_34308,N_29572,N_29746);
nor U34309 (N_34309,N_29479,N_27401);
and U34310 (N_34310,N_27130,N_27567);
and U34311 (N_34311,N_27558,N_29278);
nand U34312 (N_34312,N_28719,N_29125);
xnor U34313 (N_34313,N_27952,N_27433);
and U34314 (N_34314,N_29746,N_25990);
nand U34315 (N_34315,N_29584,N_26455);
xnor U34316 (N_34316,N_27975,N_25350);
nor U34317 (N_34317,N_25276,N_29908);
or U34318 (N_34318,N_25983,N_25966);
nor U34319 (N_34319,N_27381,N_27525);
nor U34320 (N_34320,N_29479,N_29957);
and U34321 (N_34321,N_29551,N_26564);
xnor U34322 (N_34322,N_26180,N_29445);
xnor U34323 (N_34323,N_25428,N_28452);
or U34324 (N_34324,N_25980,N_27431);
and U34325 (N_34325,N_27862,N_25693);
xor U34326 (N_34326,N_25419,N_25523);
or U34327 (N_34327,N_26339,N_26564);
xor U34328 (N_34328,N_25343,N_28268);
nand U34329 (N_34329,N_26403,N_29261);
and U34330 (N_34330,N_25957,N_28386);
nand U34331 (N_34331,N_27587,N_25491);
nor U34332 (N_34332,N_25333,N_27942);
nand U34333 (N_34333,N_26630,N_26860);
nor U34334 (N_34334,N_28329,N_27205);
or U34335 (N_34335,N_29920,N_27131);
nor U34336 (N_34336,N_29832,N_27429);
and U34337 (N_34337,N_26700,N_26276);
and U34338 (N_34338,N_29059,N_28614);
nor U34339 (N_34339,N_26098,N_29188);
or U34340 (N_34340,N_26496,N_29995);
or U34341 (N_34341,N_29630,N_27179);
and U34342 (N_34342,N_28161,N_28676);
xor U34343 (N_34343,N_27834,N_26545);
nor U34344 (N_34344,N_26226,N_27926);
or U34345 (N_34345,N_28539,N_28947);
or U34346 (N_34346,N_27331,N_29261);
nor U34347 (N_34347,N_25954,N_27438);
nor U34348 (N_34348,N_28206,N_27760);
and U34349 (N_34349,N_25360,N_26569);
xor U34350 (N_34350,N_25729,N_28645);
or U34351 (N_34351,N_26633,N_28063);
xor U34352 (N_34352,N_26782,N_28620);
nor U34353 (N_34353,N_26650,N_26977);
xor U34354 (N_34354,N_29486,N_28990);
nor U34355 (N_34355,N_28799,N_25802);
nand U34356 (N_34356,N_27330,N_25659);
xor U34357 (N_34357,N_25625,N_27055);
nor U34358 (N_34358,N_29823,N_26062);
nand U34359 (N_34359,N_25439,N_26323);
or U34360 (N_34360,N_28577,N_27671);
nand U34361 (N_34361,N_27516,N_26022);
or U34362 (N_34362,N_26008,N_28965);
xnor U34363 (N_34363,N_28829,N_27559);
xnor U34364 (N_34364,N_27910,N_29001);
nand U34365 (N_34365,N_29680,N_29486);
or U34366 (N_34366,N_27480,N_26223);
and U34367 (N_34367,N_28424,N_28819);
nor U34368 (N_34368,N_26567,N_29475);
nand U34369 (N_34369,N_27133,N_27838);
and U34370 (N_34370,N_28379,N_26932);
and U34371 (N_34371,N_26786,N_28478);
or U34372 (N_34372,N_28757,N_27690);
xor U34373 (N_34373,N_29200,N_26859);
nand U34374 (N_34374,N_27496,N_26159);
or U34375 (N_34375,N_26028,N_27585);
nor U34376 (N_34376,N_26815,N_29100);
nand U34377 (N_34377,N_29420,N_28043);
or U34378 (N_34378,N_28930,N_26091);
xor U34379 (N_34379,N_28112,N_27543);
nor U34380 (N_34380,N_29997,N_27706);
nor U34381 (N_34381,N_28340,N_28305);
xnor U34382 (N_34382,N_27366,N_27728);
or U34383 (N_34383,N_28483,N_26923);
or U34384 (N_34384,N_29898,N_29363);
nor U34385 (N_34385,N_25337,N_26325);
nand U34386 (N_34386,N_25520,N_25080);
xnor U34387 (N_34387,N_29622,N_28452);
nand U34388 (N_34388,N_25551,N_28440);
nor U34389 (N_34389,N_29393,N_29181);
and U34390 (N_34390,N_29462,N_26717);
nand U34391 (N_34391,N_29082,N_26837);
nor U34392 (N_34392,N_29944,N_25310);
nand U34393 (N_34393,N_26523,N_28958);
or U34394 (N_34394,N_25752,N_29023);
or U34395 (N_34395,N_28325,N_27553);
xor U34396 (N_34396,N_28064,N_27739);
nor U34397 (N_34397,N_28158,N_29763);
nor U34398 (N_34398,N_29602,N_28978);
or U34399 (N_34399,N_28590,N_25803);
and U34400 (N_34400,N_28650,N_29965);
xnor U34401 (N_34401,N_27017,N_27493);
nor U34402 (N_34402,N_25993,N_28792);
or U34403 (N_34403,N_25818,N_25921);
xnor U34404 (N_34404,N_27907,N_29864);
or U34405 (N_34405,N_25275,N_25509);
or U34406 (N_34406,N_27550,N_29899);
or U34407 (N_34407,N_27208,N_29553);
nor U34408 (N_34408,N_26848,N_26571);
and U34409 (N_34409,N_28969,N_25105);
or U34410 (N_34410,N_26808,N_28306);
and U34411 (N_34411,N_25083,N_28123);
nor U34412 (N_34412,N_25145,N_29518);
xnor U34413 (N_34413,N_25717,N_27281);
or U34414 (N_34414,N_26052,N_25050);
nand U34415 (N_34415,N_27611,N_25486);
and U34416 (N_34416,N_28893,N_28626);
or U34417 (N_34417,N_28614,N_29526);
xor U34418 (N_34418,N_29743,N_25466);
nor U34419 (N_34419,N_25329,N_27432);
nand U34420 (N_34420,N_27246,N_27504);
xor U34421 (N_34421,N_29529,N_27430);
nand U34422 (N_34422,N_27676,N_28255);
xnor U34423 (N_34423,N_27528,N_28216);
xor U34424 (N_34424,N_26407,N_26823);
xnor U34425 (N_34425,N_26190,N_29178);
nor U34426 (N_34426,N_29703,N_26887);
or U34427 (N_34427,N_29576,N_29057);
nand U34428 (N_34428,N_26275,N_29902);
nand U34429 (N_34429,N_28821,N_26147);
nand U34430 (N_34430,N_25881,N_25089);
or U34431 (N_34431,N_25922,N_28624);
or U34432 (N_34432,N_28491,N_27994);
nand U34433 (N_34433,N_26627,N_28931);
and U34434 (N_34434,N_26811,N_25036);
nor U34435 (N_34435,N_25820,N_29798);
nand U34436 (N_34436,N_25939,N_25188);
or U34437 (N_34437,N_27374,N_28349);
or U34438 (N_34438,N_29881,N_26310);
and U34439 (N_34439,N_25451,N_28269);
xnor U34440 (N_34440,N_25104,N_29783);
and U34441 (N_34441,N_28339,N_25317);
and U34442 (N_34442,N_25931,N_29108);
xor U34443 (N_34443,N_29652,N_25546);
and U34444 (N_34444,N_26640,N_25887);
nor U34445 (N_34445,N_25888,N_26196);
nand U34446 (N_34446,N_28241,N_26838);
xnor U34447 (N_34447,N_29526,N_29120);
nor U34448 (N_34448,N_25560,N_28421);
nand U34449 (N_34449,N_25803,N_26378);
or U34450 (N_34450,N_29584,N_25589);
or U34451 (N_34451,N_28525,N_25137);
xnor U34452 (N_34452,N_29504,N_25951);
or U34453 (N_34453,N_25720,N_27802);
and U34454 (N_34454,N_28783,N_28525);
or U34455 (N_34455,N_28538,N_26854);
xor U34456 (N_34456,N_28379,N_29327);
and U34457 (N_34457,N_25256,N_25745);
and U34458 (N_34458,N_28321,N_27595);
and U34459 (N_34459,N_25448,N_28116);
nor U34460 (N_34460,N_29877,N_25104);
nor U34461 (N_34461,N_28748,N_25326);
or U34462 (N_34462,N_25432,N_29915);
and U34463 (N_34463,N_28418,N_28549);
nand U34464 (N_34464,N_25416,N_27036);
and U34465 (N_34465,N_28925,N_29763);
nand U34466 (N_34466,N_29755,N_27317);
xnor U34467 (N_34467,N_26461,N_28633);
nand U34468 (N_34468,N_25237,N_25828);
and U34469 (N_34469,N_28092,N_26918);
nor U34470 (N_34470,N_27631,N_28077);
nor U34471 (N_34471,N_28674,N_27632);
and U34472 (N_34472,N_26018,N_28967);
nand U34473 (N_34473,N_27252,N_29084);
and U34474 (N_34474,N_29183,N_25840);
xor U34475 (N_34475,N_28220,N_25189);
or U34476 (N_34476,N_28527,N_28339);
and U34477 (N_34477,N_25264,N_27997);
nand U34478 (N_34478,N_27115,N_29263);
nand U34479 (N_34479,N_28559,N_29936);
nor U34480 (N_34480,N_28657,N_26965);
and U34481 (N_34481,N_28909,N_29049);
or U34482 (N_34482,N_26000,N_26127);
nand U34483 (N_34483,N_28631,N_27638);
xor U34484 (N_34484,N_27708,N_29431);
and U34485 (N_34485,N_28235,N_25010);
xnor U34486 (N_34486,N_29083,N_27016);
xnor U34487 (N_34487,N_25599,N_25676);
nand U34488 (N_34488,N_26552,N_29093);
and U34489 (N_34489,N_28423,N_27658);
or U34490 (N_34490,N_29132,N_27877);
and U34491 (N_34491,N_25232,N_28344);
nor U34492 (N_34492,N_29145,N_29294);
and U34493 (N_34493,N_25971,N_26697);
or U34494 (N_34494,N_29022,N_25146);
xor U34495 (N_34495,N_25244,N_27583);
xnor U34496 (N_34496,N_25636,N_28778);
nor U34497 (N_34497,N_25504,N_25034);
and U34498 (N_34498,N_28484,N_28487);
or U34499 (N_34499,N_27524,N_29455);
or U34500 (N_34500,N_27771,N_27616);
nand U34501 (N_34501,N_27616,N_25013);
and U34502 (N_34502,N_29989,N_29623);
nor U34503 (N_34503,N_29429,N_29989);
and U34504 (N_34504,N_25694,N_27305);
xnor U34505 (N_34505,N_25737,N_25256);
xnor U34506 (N_34506,N_29563,N_29545);
nor U34507 (N_34507,N_29399,N_25365);
xor U34508 (N_34508,N_28996,N_26646);
xor U34509 (N_34509,N_25858,N_27830);
nand U34510 (N_34510,N_27043,N_29981);
xnor U34511 (N_34511,N_28521,N_27579);
nor U34512 (N_34512,N_25055,N_29037);
xnor U34513 (N_34513,N_28822,N_25234);
nor U34514 (N_34514,N_25969,N_26688);
or U34515 (N_34515,N_26934,N_27419);
or U34516 (N_34516,N_27141,N_29951);
nand U34517 (N_34517,N_29725,N_27751);
nor U34518 (N_34518,N_29300,N_29371);
xnor U34519 (N_34519,N_25614,N_28681);
nand U34520 (N_34520,N_26330,N_28275);
nor U34521 (N_34521,N_28108,N_25696);
nor U34522 (N_34522,N_25667,N_25443);
nor U34523 (N_34523,N_27040,N_25432);
nand U34524 (N_34524,N_29087,N_28384);
nand U34525 (N_34525,N_25311,N_25899);
or U34526 (N_34526,N_28601,N_28155);
and U34527 (N_34527,N_26291,N_26162);
xnor U34528 (N_34528,N_26940,N_27983);
nor U34529 (N_34529,N_27014,N_28357);
nor U34530 (N_34530,N_27806,N_25791);
xor U34531 (N_34531,N_29585,N_29095);
nor U34532 (N_34532,N_26782,N_29191);
or U34533 (N_34533,N_27140,N_28348);
or U34534 (N_34534,N_28120,N_26927);
and U34535 (N_34535,N_27812,N_27734);
nand U34536 (N_34536,N_28275,N_26124);
and U34537 (N_34537,N_29069,N_27719);
or U34538 (N_34538,N_27038,N_26324);
nor U34539 (N_34539,N_28642,N_26968);
and U34540 (N_34540,N_28281,N_29809);
or U34541 (N_34541,N_28851,N_25030);
xor U34542 (N_34542,N_29183,N_26416);
nor U34543 (N_34543,N_28641,N_26293);
xnor U34544 (N_34544,N_29460,N_27055);
or U34545 (N_34545,N_28474,N_26263);
or U34546 (N_34546,N_25543,N_28676);
xnor U34547 (N_34547,N_27921,N_28185);
nor U34548 (N_34548,N_25426,N_26299);
or U34549 (N_34549,N_27466,N_28678);
nand U34550 (N_34550,N_26435,N_27874);
nor U34551 (N_34551,N_29603,N_28669);
nand U34552 (N_34552,N_29284,N_25472);
xnor U34553 (N_34553,N_26020,N_27015);
xor U34554 (N_34554,N_26055,N_26777);
xor U34555 (N_34555,N_25232,N_28986);
and U34556 (N_34556,N_25944,N_26545);
or U34557 (N_34557,N_25168,N_29348);
xnor U34558 (N_34558,N_29363,N_25428);
nand U34559 (N_34559,N_29488,N_27210);
xor U34560 (N_34560,N_29428,N_28770);
xor U34561 (N_34561,N_26411,N_25371);
xor U34562 (N_34562,N_27080,N_25227);
nor U34563 (N_34563,N_25224,N_29745);
and U34564 (N_34564,N_25443,N_25653);
nor U34565 (N_34565,N_28570,N_26397);
and U34566 (N_34566,N_27150,N_27112);
nand U34567 (N_34567,N_28024,N_27014);
nand U34568 (N_34568,N_26111,N_29902);
nor U34569 (N_34569,N_27180,N_26643);
xnor U34570 (N_34570,N_28972,N_28011);
xnor U34571 (N_34571,N_27829,N_25054);
nand U34572 (N_34572,N_27295,N_25438);
xnor U34573 (N_34573,N_26707,N_28827);
nand U34574 (N_34574,N_26535,N_25535);
and U34575 (N_34575,N_27119,N_28460);
nand U34576 (N_34576,N_27931,N_25655);
or U34577 (N_34577,N_25803,N_28985);
or U34578 (N_34578,N_28629,N_27435);
or U34579 (N_34579,N_27273,N_29470);
and U34580 (N_34580,N_29529,N_25998);
nor U34581 (N_34581,N_26775,N_29041);
xnor U34582 (N_34582,N_25038,N_29430);
or U34583 (N_34583,N_26545,N_27640);
and U34584 (N_34584,N_29733,N_25658);
xnor U34585 (N_34585,N_29244,N_28913);
xnor U34586 (N_34586,N_28816,N_29264);
or U34587 (N_34587,N_27770,N_25036);
or U34588 (N_34588,N_27711,N_25387);
nand U34589 (N_34589,N_28586,N_25579);
or U34590 (N_34590,N_29824,N_29194);
or U34591 (N_34591,N_29436,N_25064);
xnor U34592 (N_34592,N_28528,N_28877);
or U34593 (N_34593,N_25491,N_25862);
nand U34594 (N_34594,N_26273,N_25543);
nand U34595 (N_34595,N_27295,N_28056);
xor U34596 (N_34596,N_28509,N_26460);
and U34597 (N_34597,N_28792,N_25605);
xor U34598 (N_34598,N_25066,N_29944);
nor U34599 (N_34599,N_26924,N_28764);
xor U34600 (N_34600,N_25783,N_27894);
nor U34601 (N_34601,N_29814,N_28962);
or U34602 (N_34602,N_27840,N_28192);
xor U34603 (N_34603,N_26856,N_28660);
xnor U34604 (N_34604,N_25155,N_26181);
or U34605 (N_34605,N_26661,N_25658);
xor U34606 (N_34606,N_28442,N_29367);
xor U34607 (N_34607,N_25737,N_26218);
nor U34608 (N_34608,N_29393,N_25996);
or U34609 (N_34609,N_29080,N_28071);
nor U34610 (N_34610,N_28363,N_25531);
nand U34611 (N_34611,N_26576,N_28058);
and U34612 (N_34612,N_28601,N_28418);
and U34613 (N_34613,N_29026,N_27783);
or U34614 (N_34614,N_26042,N_27819);
nand U34615 (N_34615,N_29880,N_27187);
nor U34616 (N_34616,N_29616,N_25862);
nor U34617 (N_34617,N_28718,N_26324);
nand U34618 (N_34618,N_28626,N_29549);
nand U34619 (N_34619,N_28645,N_25779);
or U34620 (N_34620,N_28129,N_26211);
and U34621 (N_34621,N_29781,N_25711);
and U34622 (N_34622,N_27995,N_29272);
xnor U34623 (N_34623,N_25517,N_25710);
nor U34624 (N_34624,N_28853,N_27607);
and U34625 (N_34625,N_29054,N_25134);
or U34626 (N_34626,N_25683,N_26503);
nand U34627 (N_34627,N_29463,N_29482);
xor U34628 (N_34628,N_26080,N_29485);
nand U34629 (N_34629,N_27775,N_26980);
and U34630 (N_34630,N_25042,N_27454);
nand U34631 (N_34631,N_28857,N_25287);
or U34632 (N_34632,N_25067,N_27155);
xnor U34633 (N_34633,N_29893,N_26525);
and U34634 (N_34634,N_25757,N_25183);
nand U34635 (N_34635,N_28278,N_26354);
xnor U34636 (N_34636,N_29805,N_27811);
xor U34637 (N_34637,N_28500,N_26537);
xor U34638 (N_34638,N_25237,N_25819);
nor U34639 (N_34639,N_27167,N_25736);
nor U34640 (N_34640,N_25334,N_25761);
nand U34641 (N_34641,N_27276,N_25274);
xor U34642 (N_34642,N_25520,N_27155);
nor U34643 (N_34643,N_29668,N_25585);
nand U34644 (N_34644,N_25616,N_29863);
and U34645 (N_34645,N_25728,N_27373);
nand U34646 (N_34646,N_29382,N_26327);
nor U34647 (N_34647,N_26756,N_26587);
and U34648 (N_34648,N_25466,N_25078);
nand U34649 (N_34649,N_28868,N_25349);
nor U34650 (N_34650,N_26994,N_29476);
and U34651 (N_34651,N_29502,N_27399);
nand U34652 (N_34652,N_25405,N_28544);
or U34653 (N_34653,N_28280,N_25433);
nand U34654 (N_34654,N_28937,N_28209);
xor U34655 (N_34655,N_28036,N_26047);
or U34656 (N_34656,N_27695,N_28295);
or U34657 (N_34657,N_25257,N_27166);
or U34658 (N_34658,N_26794,N_28444);
nand U34659 (N_34659,N_26574,N_29413);
nand U34660 (N_34660,N_28349,N_27860);
and U34661 (N_34661,N_26473,N_26820);
and U34662 (N_34662,N_26998,N_29029);
nand U34663 (N_34663,N_28833,N_26688);
nor U34664 (N_34664,N_25471,N_29996);
xnor U34665 (N_34665,N_28967,N_25734);
and U34666 (N_34666,N_28403,N_27585);
and U34667 (N_34667,N_25742,N_25642);
xnor U34668 (N_34668,N_26196,N_28598);
nand U34669 (N_34669,N_28814,N_26847);
nand U34670 (N_34670,N_25271,N_25027);
xor U34671 (N_34671,N_28360,N_29822);
and U34672 (N_34672,N_26380,N_29613);
nand U34673 (N_34673,N_26312,N_28644);
xnor U34674 (N_34674,N_27394,N_27154);
xnor U34675 (N_34675,N_27702,N_28258);
and U34676 (N_34676,N_29442,N_26433);
and U34677 (N_34677,N_27552,N_28130);
and U34678 (N_34678,N_26570,N_26288);
xor U34679 (N_34679,N_25295,N_26379);
xor U34680 (N_34680,N_28925,N_29410);
nor U34681 (N_34681,N_28715,N_27544);
or U34682 (N_34682,N_25807,N_25599);
xor U34683 (N_34683,N_28370,N_28278);
and U34684 (N_34684,N_27744,N_25967);
xnor U34685 (N_34685,N_26333,N_29370);
or U34686 (N_34686,N_25627,N_28435);
and U34687 (N_34687,N_25418,N_25915);
xnor U34688 (N_34688,N_28547,N_26050);
or U34689 (N_34689,N_29480,N_28022);
nor U34690 (N_34690,N_25061,N_29740);
nor U34691 (N_34691,N_27078,N_29168);
or U34692 (N_34692,N_26422,N_29053);
and U34693 (N_34693,N_29074,N_28476);
nor U34694 (N_34694,N_28670,N_25957);
xor U34695 (N_34695,N_26103,N_26454);
or U34696 (N_34696,N_29836,N_27365);
or U34697 (N_34697,N_29098,N_26753);
or U34698 (N_34698,N_29201,N_27383);
or U34699 (N_34699,N_25198,N_26687);
or U34700 (N_34700,N_27125,N_27439);
or U34701 (N_34701,N_26571,N_26961);
nand U34702 (N_34702,N_26390,N_29527);
nand U34703 (N_34703,N_25209,N_27967);
nor U34704 (N_34704,N_29950,N_29611);
nor U34705 (N_34705,N_28375,N_28205);
nand U34706 (N_34706,N_28298,N_28591);
and U34707 (N_34707,N_27417,N_25829);
or U34708 (N_34708,N_27859,N_26691);
xor U34709 (N_34709,N_26849,N_25647);
or U34710 (N_34710,N_28175,N_25338);
nand U34711 (N_34711,N_27536,N_29218);
nor U34712 (N_34712,N_26113,N_28711);
nor U34713 (N_34713,N_29425,N_25781);
and U34714 (N_34714,N_29710,N_26715);
and U34715 (N_34715,N_26604,N_26795);
or U34716 (N_34716,N_27860,N_29242);
and U34717 (N_34717,N_27286,N_25985);
xnor U34718 (N_34718,N_28156,N_27587);
nor U34719 (N_34719,N_29431,N_28024);
or U34720 (N_34720,N_25922,N_28034);
nor U34721 (N_34721,N_26576,N_27328);
nand U34722 (N_34722,N_28172,N_26011);
and U34723 (N_34723,N_27788,N_26269);
nor U34724 (N_34724,N_28374,N_29102);
or U34725 (N_34725,N_28934,N_27037);
xnor U34726 (N_34726,N_26096,N_27021);
and U34727 (N_34727,N_25249,N_28642);
nor U34728 (N_34728,N_27186,N_26129);
xnor U34729 (N_34729,N_28236,N_25744);
xor U34730 (N_34730,N_28754,N_27216);
and U34731 (N_34731,N_28751,N_28966);
nand U34732 (N_34732,N_27142,N_25300);
xor U34733 (N_34733,N_28668,N_29469);
xor U34734 (N_34734,N_25725,N_27866);
xor U34735 (N_34735,N_28947,N_26733);
or U34736 (N_34736,N_29606,N_25441);
xor U34737 (N_34737,N_27912,N_28805);
xor U34738 (N_34738,N_26886,N_29435);
and U34739 (N_34739,N_27389,N_25793);
and U34740 (N_34740,N_29811,N_25895);
nand U34741 (N_34741,N_29008,N_27225);
and U34742 (N_34742,N_27506,N_28512);
and U34743 (N_34743,N_29344,N_25835);
and U34744 (N_34744,N_25879,N_25091);
or U34745 (N_34745,N_29333,N_26615);
nand U34746 (N_34746,N_25236,N_27753);
nor U34747 (N_34747,N_27365,N_25084);
and U34748 (N_34748,N_26899,N_25354);
nor U34749 (N_34749,N_29997,N_26007);
nand U34750 (N_34750,N_27673,N_28190);
nor U34751 (N_34751,N_29560,N_27891);
xor U34752 (N_34752,N_26724,N_27752);
or U34753 (N_34753,N_27361,N_25021);
or U34754 (N_34754,N_29488,N_26932);
xnor U34755 (N_34755,N_29335,N_26379);
or U34756 (N_34756,N_29152,N_29697);
or U34757 (N_34757,N_27085,N_25747);
nor U34758 (N_34758,N_25750,N_25387);
xnor U34759 (N_34759,N_29430,N_29392);
and U34760 (N_34760,N_25278,N_26492);
nor U34761 (N_34761,N_29204,N_27678);
nand U34762 (N_34762,N_27239,N_27394);
or U34763 (N_34763,N_25804,N_25330);
nor U34764 (N_34764,N_27883,N_26259);
or U34765 (N_34765,N_29357,N_29354);
and U34766 (N_34766,N_25880,N_29352);
and U34767 (N_34767,N_29168,N_26603);
and U34768 (N_34768,N_27192,N_29187);
xor U34769 (N_34769,N_26908,N_27285);
nor U34770 (N_34770,N_26869,N_25109);
nor U34771 (N_34771,N_27232,N_26230);
xnor U34772 (N_34772,N_25854,N_26330);
nor U34773 (N_34773,N_27703,N_29761);
xnor U34774 (N_34774,N_29235,N_25914);
or U34775 (N_34775,N_28192,N_27671);
and U34776 (N_34776,N_28254,N_27403);
and U34777 (N_34777,N_27625,N_27797);
nand U34778 (N_34778,N_25212,N_29074);
nor U34779 (N_34779,N_26833,N_25570);
and U34780 (N_34780,N_25788,N_26680);
nand U34781 (N_34781,N_27850,N_27090);
and U34782 (N_34782,N_27121,N_27188);
and U34783 (N_34783,N_27975,N_28652);
nor U34784 (N_34784,N_25766,N_28582);
nand U34785 (N_34785,N_29724,N_26751);
or U34786 (N_34786,N_28689,N_28417);
nor U34787 (N_34787,N_29141,N_29697);
nor U34788 (N_34788,N_25127,N_26331);
xnor U34789 (N_34789,N_29263,N_27601);
or U34790 (N_34790,N_28726,N_28626);
nor U34791 (N_34791,N_29243,N_26226);
xor U34792 (N_34792,N_27692,N_27020);
or U34793 (N_34793,N_27649,N_29299);
and U34794 (N_34794,N_26415,N_27296);
nor U34795 (N_34795,N_25960,N_28565);
and U34796 (N_34796,N_28860,N_28457);
or U34797 (N_34797,N_25121,N_29561);
xor U34798 (N_34798,N_27189,N_28900);
or U34799 (N_34799,N_25301,N_26506);
xor U34800 (N_34800,N_26320,N_27297);
nor U34801 (N_34801,N_25208,N_28463);
or U34802 (N_34802,N_29960,N_29768);
or U34803 (N_34803,N_25295,N_25325);
or U34804 (N_34804,N_29796,N_27271);
xnor U34805 (N_34805,N_27367,N_26160);
or U34806 (N_34806,N_28078,N_29022);
and U34807 (N_34807,N_28281,N_27081);
and U34808 (N_34808,N_25027,N_26580);
and U34809 (N_34809,N_25497,N_26478);
nand U34810 (N_34810,N_28180,N_27614);
and U34811 (N_34811,N_25228,N_26381);
nand U34812 (N_34812,N_26771,N_25981);
or U34813 (N_34813,N_29911,N_25371);
nand U34814 (N_34814,N_28371,N_29262);
nand U34815 (N_34815,N_26750,N_29572);
or U34816 (N_34816,N_28947,N_28497);
nor U34817 (N_34817,N_27765,N_27892);
and U34818 (N_34818,N_26717,N_26777);
xor U34819 (N_34819,N_29161,N_26872);
nand U34820 (N_34820,N_27512,N_28358);
nor U34821 (N_34821,N_27952,N_27877);
nand U34822 (N_34822,N_26320,N_25419);
nand U34823 (N_34823,N_27370,N_27068);
xor U34824 (N_34824,N_26624,N_28446);
and U34825 (N_34825,N_27090,N_29379);
nand U34826 (N_34826,N_26775,N_28066);
or U34827 (N_34827,N_27813,N_27004);
xnor U34828 (N_34828,N_25502,N_29496);
nand U34829 (N_34829,N_28647,N_28989);
xor U34830 (N_34830,N_29982,N_28164);
xnor U34831 (N_34831,N_29062,N_25940);
xor U34832 (N_34832,N_27355,N_26835);
and U34833 (N_34833,N_27739,N_25121);
xor U34834 (N_34834,N_26247,N_27925);
or U34835 (N_34835,N_25896,N_29575);
nor U34836 (N_34836,N_25384,N_28570);
nor U34837 (N_34837,N_28383,N_28695);
xor U34838 (N_34838,N_26073,N_25666);
and U34839 (N_34839,N_25911,N_26578);
nand U34840 (N_34840,N_29566,N_28584);
nand U34841 (N_34841,N_28633,N_29784);
or U34842 (N_34842,N_29513,N_25146);
nand U34843 (N_34843,N_26873,N_29017);
xor U34844 (N_34844,N_28100,N_25725);
nand U34845 (N_34845,N_28245,N_29763);
nand U34846 (N_34846,N_26826,N_28120);
nand U34847 (N_34847,N_26891,N_28263);
xnor U34848 (N_34848,N_26886,N_27657);
nand U34849 (N_34849,N_25328,N_29481);
nand U34850 (N_34850,N_27388,N_27707);
nor U34851 (N_34851,N_29933,N_29094);
nand U34852 (N_34852,N_28370,N_29529);
nand U34853 (N_34853,N_26586,N_28384);
and U34854 (N_34854,N_28274,N_29914);
nand U34855 (N_34855,N_25701,N_26627);
nand U34856 (N_34856,N_26714,N_27029);
or U34857 (N_34857,N_28226,N_28295);
xnor U34858 (N_34858,N_29440,N_29172);
or U34859 (N_34859,N_29239,N_28862);
nand U34860 (N_34860,N_29288,N_27624);
xnor U34861 (N_34861,N_27035,N_25401);
xor U34862 (N_34862,N_27535,N_26489);
nand U34863 (N_34863,N_26201,N_29146);
and U34864 (N_34864,N_25038,N_29932);
nand U34865 (N_34865,N_29403,N_25349);
or U34866 (N_34866,N_27230,N_29929);
and U34867 (N_34867,N_26744,N_26665);
nor U34868 (N_34868,N_28244,N_29564);
xor U34869 (N_34869,N_29391,N_25749);
nor U34870 (N_34870,N_29244,N_25084);
nand U34871 (N_34871,N_27194,N_27029);
and U34872 (N_34872,N_26455,N_26753);
and U34873 (N_34873,N_26203,N_29026);
nor U34874 (N_34874,N_27681,N_28724);
nor U34875 (N_34875,N_27382,N_29497);
nand U34876 (N_34876,N_29442,N_25896);
xor U34877 (N_34877,N_27268,N_25104);
and U34878 (N_34878,N_26825,N_26806);
nor U34879 (N_34879,N_28170,N_26340);
xor U34880 (N_34880,N_27845,N_29200);
nor U34881 (N_34881,N_27858,N_26660);
or U34882 (N_34882,N_28925,N_27479);
or U34883 (N_34883,N_26875,N_27938);
and U34884 (N_34884,N_28355,N_28568);
or U34885 (N_34885,N_25265,N_29317);
and U34886 (N_34886,N_27129,N_28432);
nand U34887 (N_34887,N_29488,N_26573);
xnor U34888 (N_34888,N_27289,N_25819);
nand U34889 (N_34889,N_28812,N_28956);
nor U34890 (N_34890,N_25986,N_26315);
xor U34891 (N_34891,N_25998,N_29770);
xnor U34892 (N_34892,N_27117,N_26195);
or U34893 (N_34893,N_26680,N_28972);
xor U34894 (N_34894,N_27508,N_25937);
nor U34895 (N_34895,N_28735,N_29796);
xnor U34896 (N_34896,N_26463,N_29375);
nor U34897 (N_34897,N_26871,N_27453);
or U34898 (N_34898,N_26119,N_26621);
nand U34899 (N_34899,N_29310,N_29946);
nor U34900 (N_34900,N_25274,N_25397);
and U34901 (N_34901,N_25557,N_27459);
and U34902 (N_34902,N_27406,N_26840);
or U34903 (N_34903,N_28352,N_25418);
and U34904 (N_34904,N_27776,N_29213);
xor U34905 (N_34905,N_26803,N_29576);
xnor U34906 (N_34906,N_28991,N_25286);
or U34907 (N_34907,N_29668,N_26546);
and U34908 (N_34908,N_26039,N_28121);
or U34909 (N_34909,N_26860,N_27353);
xnor U34910 (N_34910,N_29108,N_28560);
or U34911 (N_34911,N_25131,N_27556);
or U34912 (N_34912,N_27563,N_29452);
and U34913 (N_34913,N_28681,N_28609);
nand U34914 (N_34914,N_29688,N_28358);
and U34915 (N_34915,N_26860,N_25222);
nor U34916 (N_34916,N_29585,N_28784);
and U34917 (N_34917,N_29541,N_28425);
nor U34918 (N_34918,N_29107,N_29489);
xor U34919 (N_34919,N_26056,N_28481);
xor U34920 (N_34920,N_27222,N_28574);
nand U34921 (N_34921,N_25763,N_25703);
nor U34922 (N_34922,N_26228,N_28322);
or U34923 (N_34923,N_29964,N_27345);
nand U34924 (N_34924,N_29328,N_25619);
or U34925 (N_34925,N_28583,N_27804);
xor U34926 (N_34926,N_28861,N_29602);
xor U34927 (N_34927,N_28333,N_28861);
and U34928 (N_34928,N_25579,N_28179);
nand U34929 (N_34929,N_25209,N_27940);
nor U34930 (N_34930,N_25836,N_29843);
and U34931 (N_34931,N_26293,N_28740);
and U34932 (N_34932,N_29097,N_28102);
nor U34933 (N_34933,N_28671,N_29359);
nor U34934 (N_34934,N_27837,N_27522);
or U34935 (N_34935,N_28260,N_27920);
nand U34936 (N_34936,N_27628,N_27101);
xnor U34937 (N_34937,N_25522,N_27935);
or U34938 (N_34938,N_29723,N_29933);
nor U34939 (N_34939,N_28486,N_28649);
xor U34940 (N_34940,N_28792,N_28176);
and U34941 (N_34941,N_25809,N_28930);
xor U34942 (N_34942,N_29717,N_26458);
xnor U34943 (N_34943,N_29198,N_28581);
or U34944 (N_34944,N_26986,N_28802);
nor U34945 (N_34945,N_26636,N_28303);
nand U34946 (N_34946,N_29105,N_27176);
and U34947 (N_34947,N_27877,N_27855);
nand U34948 (N_34948,N_29743,N_28187);
and U34949 (N_34949,N_28384,N_25416);
xnor U34950 (N_34950,N_28304,N_25054);
nor U34951 (N_34951,N_26996,N_25440);
nand U34952 (N_34952,N_25674,N_26591);
and U34953 (N_34953,N_25073,N_27788);
and U34954 (N_34954,N_26620,N_26210);
xnor U34955 (N_34955,N_25276,N_27788);
nor U34956 (N_34956,N_27311,N_25850);
and U34957 (N_34957,N_26643,N_29465);
nor U34958 (N_34958,N_25354,N_25364);
nand U34959 (N_34959,N_28159,N_27735);
nor U34960 (N_34960,N_25685,N_27131);
and U34961 (N_34961,N_26814,N_26188);
or U34962 (N_34962,N_27516,N_27824);
or U34963 (N_34963,N_25782,N_26073);
nand U34964 (N_34964,N_27521,N_29337);
or U34965 (N_34965,N_26350,N_27469);
and U34966 (N_34966,N_26535,N_29215);
xor U34967 (N_34967,N_26696,N_27944);
xor U34968 (N_34968,N_27303,N_26987);
and U34969 (N_34969,N_25565,N_29342);
xor U34970 (N_34970,N_27083,N_25898);
nand U34971 (N_34971,N_26195,N_25000);
xor U34972 (N_34972,N_26303,N_26267);
xor U34973 (N_34973,N_25395,N_26812);
nor U34974 (N_34974,N_28361,N_27098);
xor U34975 (N_34975,N_28754,N_29909);
nor U34976 (N_34976,N_26074,N_27075);
xnor U34977 (N_34977,N_29127,N_26579);
nor U34978 (N_34978,N_29928,N_25702);
nand U34979 (N_34979,N_27759,N_27131);
and U34980 (N_34980,N_29196,N_25476);
nor U34981 (N_34981,N_27169,N_28889);
nand U34982 (N_34982,N_28574,N_25213);
and U34983 (N_34983,N_28746,N_28400);
and U34984 (N_34984,N_25392,N_25414);
nand U34985 (N_34985,N_27501,N_27114);
or U34986 (N_34986,N_25022,N_29128);
nor U34987 (N_34987,N_25600,N_27330);
or U34988 (N_34988,N_25644,N_25524);
nor U34989 (N_34989,N_27592,N_28316);
and U34990 (N_34990,N_29022,N_29964);
or U34991 (N_34991,N_25636,N_27019);
nand U34992 (N_34992,N_29663,N_29295);
nand U34993 (N_34993,N_26716,N_27315);
or U34994 (N_34994,N_29479,N_25327);
and U34995 (N_34995,N_28873,N_28422);
xnor U34996 (N_34996,N_28402,N_29290);
nor U34997 (N_34997,N_28337,N_28668);
xor U34998 (N_34998,N_29754,N_28727);
xor U34999 (N_34999,N_27625,N_29819);
and U35000 (N_35000,N_32453,N_30193);
nor U35001 (N_35001,N_34710,N_34999);
nand U35002 (N_35002,N_32837,N_30207);
or U35003 (N_35003,N_31692,N_33993);
or U35004 (N_35004,N_34731,N_30325);
or U35005 (N_35005,N_31982,N_30400);
or U35006 (N_35006,N_33487,N_34524);
xnor U35007 (N_35007,N_34118,N_30503);
nand U35008 (N_35008,N_31937,N_34860);
xnor U35009 (N_35009,N_32415,N_32478);
nor U35010 (N_35010,N_34475,N_31671);
nand U35011 (N_35011,N_32222,N_33722);
nor U35012 (N_35012,N_32368,N_30203);
and U35013 (N_35013,N_31260,N_34983);
xnor U35014 (N_35014,N_34187,N_33201);
xor U35015 (N_35015,N_34142,N_32545);
nor U35016 (N_35016,N_34541,N_30313);
xor U35017 (N_35017,N_32060,N_34743);
xnor U35018 (N_35018,N_32558,N_30577);
nand U35019 (N_35019,N_31546,N_33358);
or U35020 (N_35020,N_33910,N_30861);
nor U35021 (N_35021,N_30172,N_33405);
nor U35022 (N_35022,N_31928,N_34090);
or U35023 (N_35023,N_33447,N_34153);
or U35024 (N_35024,N_31664,N_33871);
or U35025 (N_35025,N_34096,N_30608);
nor U35026 (N_35026,N_30891,N_33788);
nor U35027 (N_35027,N_33591,N_33991);
nand U35028 (N_35028,N_34627,N_32312);
xor U35029 (N_35029,N_30461,N_33978);
or U35030 (N_35030,N_30789,N_34181);
nand U35031 (N_35031,N_31477,N_30285);
or U35032 (N_35032,N_31027,N_33980);
xor U35033 (N_35033,N_34098,N_32143);
nand U35034 (N_35034,N_33678,N_30087);
nand U35035 (N_35035,N_31392,N_34990);
or U35036 (N_35036,N_31321,N_34659);
xor U35037 (N_35037,N_34300,N_31087);
or U35038 (N_35038,N_30790,N_33459);
or U35039 (N_35039,N_34389,N_32433);
nor U35040 (N_35040,N_34135,N_30564);
nand U35041 (N_35041,N_33250,N_30659);
nor U35042 (N_35042,N_33887,N_30668);
nand U35043 (N_35043,N_32903,N_31641);
nand U35044 (N_35044,N_34776,N_31877);
nor U35045 (N_35045,N_31694,N_31874);
nand U35046 (N_35046,N_33835,N_31850);
nand U35047 (N_35047,N_31881,N_33061);
nor U35048 (N_35048,N_31515,N_31174);
or U35049 (N_35049,N_31701,N_31279);
or U35050 (N_35050,N_34255,N_33840);
nand U35051 (N_35051,N_33660,N_33771);
nand U35052 (N_35052,N_34604,N_32546);
nor U35053 (N_35053,N_31512,N_30093);
nor U35054 (N_35054,N_31047,N_31401);
xor U35055 (N_35055,N_32543,N_34958);
nor U35056 (N_35056,N_32844,N_33396);
nor U35057 (N_35057,N_31151,N_34801);
nand U35058 (N_35058,N_30883,N_31436);
nor U35059 (N_35059,N_33412,N_34863);
xor U35060 (N_35060,N_30271,N_32646);
or U35061 (N_35061,N_32010,N_34257);
xnor U35062 (N_35062,N_30769,N_31788);
or U35063 (N_35063,N_32330,N_33424);
and U35064 (N_35064,N_31537,N_32776);
xnor U35065 (N_35065,N_31291,N_32264);
and U35066 (N_35066,N_32030,N_32740);
nand U35067 (N_35067,N_31536,N_34649);
nor U35068 (N_35068,N_30282,N_30167);
and U35069 (N_35069,N_34073,N_34772);
or U35070 (N_35070,N_33570,N_31767);
or U35071 (N_35071,N_31562,N_32825);
nand U35072 (N_35072,N_34719,N_33033);
or U35073 (N_35073,N_32781,N_33812);
nand U35074 (N_35074,N_30099,N_30135);
xnor U35075 (N_35075,N_33902,N_34965);
or U35076 (N_35076,N_32452,N_33572);
and U35077 (N_35077,N_30950,N_33365);
nand U35078 (N_35078,N_34907,N_33782);
nor U35079 (N_35079,N_32022,N_34109);
nor U35080 (N_35080,N_31831,N_30191);
or U35081 (N_35081,N_31393,N_31670);
xor U35082 (N_35082,N_30027,N_32340);
or U35083 (N_35083,N_31544,N_34929);
xnor U35084 (N_35084,N_34394,N_30005);
or U35085 (N_35085,N_31449,N_33411);
or U35086 (N_35086,N_33014,N_30677);
and U35087 (N_35087,N_32018,N_30540);
nor U35088 (N_35088,N_32462,N_30066);
xor U35089 (N_35089,N_30386,N_33325);
nor U35090 (N_35090,N_33148,N_31832);
and U35091 (N_35091,N_34516,N_34511);
and U35092 (N_35092,N_34635,N_34206);
or U35093 (N_35093,N_32738,N_32386);
xor U35094 (N_35094,N_31905,N_31265);
nand U35095 (N_35095,N_31303,N_30121);
xnor U35096 (N_35096,N_33481,N_33512);
xnor U35097 (N_35097,N_34613,N_33057);
nor U35098 (N_35098,N_31068,N_30017);
and U35099 (N_35099,N_30770,N_33287);
and U35100 (N_35100,N_34520,N_34736);
nand U35101 (N_35101,N_31507,N_34882);
nand U35102 (N_35102,N_34575,N_31467);
or U35103 (N_35103,N_31417,N_33097);
or U35104 (N_35104,N_30049,N_32498);
or U35105 (N_35105,N_30717,N_32783);
xor U35106 (N_35106,N_33364,N_34551);
xnor U35107 (N_35107,N_30615,N_31471);
nor U35108 (N_35108,N_30148,N_31454);
nor U35109 (N_35109,N_32073,N_34884);
nor U35110 (N_35110,N_32761,N_31330);
xnor U35111 (N_35111,N_33584,N_30817);
xnor U35112 (N_35112,N_32145,N_32810);
nor U35113 (N_35113,N_32434,N_31722);
and U35114 (N_35114,N_31560,N_32667);
and U35115 (N_35115,N_30595,N_31697);
xnor U35116 (N_35116,N_34016,N_31196);
nor U35117 (N_35117,N_33898,N_31295);
nand U35118 (N_35118,N_31731,N_31166);
or U35119 (N_35119,N_30437,N_30844);
nor U35120 (N_35120,N_31215,N_34108);
and U35121 (N_35121,N_31128,N_33431);
nor U35122 (N_35122,N_30843,N_32489);
xor U35123 (N_35123,N_30574,N_32942);
nor U35124 (N_35124,N_30641,N_31751);
xnor U35125 (N_35125,N_33836,N_34332);
xor U35126 (N_35126,N_31820,N_30962);
nand U35127 (N_35127,N_33905,N_32304);
xnor U35128 (N_35128,N_30990,N_30040);
xor U35129 (N_35129,N_34532,N_30479);
and U35130 (N_35130,N_32081,N_32767);
nor U35131 (N_35131,N_33995,N_30913);
nor U35132 (N_35132,N_31833,N_33720);
nand U35133 (N_35133,N_32564,N_34879);
or U35134 (N_35134,N_33370,N_34764);
nor U35135 (N_35135,N_33864,N_31704);
or U35136 (N_35136,N_33024,N_32590);
nand U35137 (N_35137,N_32834,N_34998);
and U35138 (N_35138,N_30170,N_34028);
xor U35139 (N_35139,N_31341,N_30477);
xnor U35140 (N_35140,N_30162,N_31849);
and U35141 (N_35141,N_32124,N_30886);
xor U35142 (N_35142,N_34839,N_32683);
and U35143 (N_35143,N_34468,N_33952);
or U35144 (N_35144,N_32083,N_31106);
or U35145 (N_35145,N_32284,N_33425);
and U35146 (N_35146,N_34423,N_30853);
or U35147 (N_35147,N_32554,N_30002);
xor U35148 (N_35148,N_30096,N_32913);
xor U35149 (N_35149,N_33826,N_34451);
nand U35150 (N_35150,N_32552,N_32529);
xor U35151 (N_35151,N_30445,N_32713);
xnor U35152 (N_35152,N_30083,N_31712);
xor U35153 (N_35153,N_32128,N_34518);
nand U35154 (N_35154,N_33217,N_30364);
and U35155 (N_35155,N_34288,N_30436);
or U35156 (N_35156,N_34192,N_34357);
or U35157 (N_35157,N_33805,N_34159);
nor U35158 (N_35158,N_34131,N_33649);
nand U35159 (N_35159,N_32146,N_31839);
and U35160 (N_35160,N_33529,N_34132);
nor U35161 (N_35161,N_33658,N_33214);
or U35162 (N_35162,N_31551,N_34012);
xor U35163 (N_35163,N_31953,N_30752);
and U35164 (N_35164,N_32806,N_33762);
nor U35165 (N_35165,N_33443,N_30555);
nor U35166 (N_35166,N_31034,N_34703);
xor U35167 (N_35167,N_34770,N_34121);
or U35168 (N_35168,N_31838,N_30820);
nand U35169 (N_35169,N_31325,N_32162);
and U35170 (N_35170,N_34393,N_30430);
xnor U35171 (N_35171,N_30932,N_30596);
xor U35172 (N_35172,N_32596,N_32390);
nand U35173 (N_35173,N_32011,N_34538);
and U35174 (N_35174,N_32585,N_31131);
nor U35175 (N_35175,N_31711,N_34818);
and U35176 (N_35176,N_32673,N_33379);
nor U35177 (N_35177,N_33809,N_32303);
nor U35178 (N_35178,N_34277,N_34535);
or U35179 (N_35179,N_33693,N_32294);
nand U35180 (N_35180,N_33011,N_30695);
xnor U35181 (N_35181,N_30665,N_31164);
xor U35182 (N_35182,N_34139,N_30388);
nor U35183 (N_35183,N_32720,N_31738);
or U35184 (N_35184,N_30954,N_32947);
or U35185 (N_35185,N_34714,N_32601);
or U35186 (N_35186,N_32748,N_30651);
and U35187 (N_35187,N_30701,N_33622);
xnor U35188 (N_35188,N_31760,N_32698);
or U35189 (N_35189,N_33093,N_32510);
nand U35190 (N_35190,N_33575,N_32805);
nor U35191 (N_35191,N_31787,N_30289);
xnor U35192 (N_35192,N_32047,N_31177);
xor U35193 (N_35193,N_34697,N_32054);
or U35194 (N_35194,N_34085,N_33844);
xor U35195 (N_35195,N_31038,N_34447);
nor U35196 (N_35196,N_31159,N_32762);
or U35197 (N_35197,N_31792,N_34563);
xor U35198 (N_35198,N_34439,N_32912);
nand U35199 (N_35199,N_33091,N_31887);
xnor U35200 (N_35200,N_32615,N_31286);
xor U35201 (N_35201,N_34773,N_33331);
nand U35202 (N_35202,N_33099,N_32387);
and U35203 (N_35203,N_33707,N_31059);
xnor U35204 (N_35204,N_33558,N_31688);
and U35205 (N_35205,N_31564,N_33779);
nand U35206 (N_35206,N_34238,N_33874);
nor U35207 (N_35207,N_30860,N_34996);
xnor U35208 (N_35208,N_31271,N_31799);
nand U35209 (N_35209,N_31500,N_31568);
nand U35210 (N_35210,N_30635,N_34299);
nor U35211 (N_35211,N_31331,N_32192);
or U35212 (N_35212,N_33078,N_30048);
nor U35213 (N_35213,N_34632,N_31635);
and U35214 (N_35214,N_33685,N_30463);
and U35215 (N_35215,N_31980,N_34750);
or U35216 (N_35216,N_33556,N_34642);
xnor U35217 (N_35217,N_31413,N_33476);
nor U35218 (N_35218,N_33967,N_32256);
or U35219 (N_35219,N_31834,N_32205);
nand U35220 (N_35220,N_33113,N_30457);
or U35221 (N_35221,N_32451,N_33798);
nor U35222 (N_35222,N_30404,N_34313);
xnor U35223 (N_35223,N_33907,N_33408);
nor U35224 (N_35224,N_33672,N_34136);
nor U35225 (N_35225,N_30622,N_32741);
and U35226 (N_35226,N_32933,N_33582);
xnor U35227 (N_35227,N_30109,N_31472);
or U35228 (N_35228,N_33847,N_30165);
xor U35229 (N_35229,N_30812,N_30984);
nor U35230 (N_35230,N_32905,N_31315);
nor U35231 (N_35231,N_32332,N_33765);
or U35232 (N_35232,N_31109,N_33116);
nor U35233 (N_35233,N_30697,N_33532);
nor U35234 (N_35234,N_31680,N_33718);
nor U35235 (N_35235,N_32640,N_30290);
nand U35236 (N_35236,N_34284,N_32426);
and U35237 (N_35237,N_33248,N_30973);
or U35238 (N_35238,N_31238,N_33210);
or U35239 (N_35239,N_34278,N_34221);
nand U35240 (N_35240,N_33657,N_31960);
nand U35241 (N_35241,N_33445,N_33708);
nor U35242 (N_35242,N_31050,N_34452);
nand U35243 (N_35243,N_34115,N_30722);
nand U35244 (N_35244,N_34218,N_31894);
nor U35245 (N_35245,N_32027,N_33258);
or U35246 (N_35246,N_34816,N_30827);
xor U35247 (N_35247,N_34976,N_30119);
xor U35248 (N_35248,N_32109,N_33252);
or U35249 (N_35249,N_32780,N_31922);
xnor U35250 (N_35250,N_32105,N_31936);
nor U35251 (N_35251,N_31004,N_31989);
and U35252 (N_35252,N_30971,N_32820);
xnor U35253 (N_35253,N_33682,N_30323);
nor U35254 (N_35254,N_32021,N_34696);
or U35255 (N_35255,N_34807,N_33262);
nand U35256 (N_35256,N_33702,N_31645);
or U35257 (N_35257,N_31088,N_30204);
and U35258 (N_35258,N_31354,N_34345);
nor U35259 (N_35259,N_30340,N_30934);
nor U35260 (N_35260,N_32964,N_34590);
nor U35261 (N_35261,N_33913,N_34715);
and U35262 (N_35262,N_32370,N_32194);
nor U35263 (N_35263,N_32526,N_31236);
nor U35264 (N_35264,N_32463,N_34078);
and U35265 (N_35265,N_33456,N_31157);
nor U35266 (N_35266,N_34975,N_31510);
and U35267 (N_35267,N_33251,N_33772);
nor U35268 (N_35268,N_30928,N_33780);
xor U35269 (N_35269,N_32324,N_31229);
nand U35270 (N_35270,N_33673,N_32659);
and U35271 (N_35271,N_30643,N_34995);
nand U35272 (N_35272,N_34971,N_34403);
xnor U35273 (N_35273,N_31559,N_30345);
nand U35274 (N_35274,N_32454,N_30147);
or U35275 (N_35275,N_33796,N_32005);
xor U35276 (N_35276,N_33477,N_30508);
xnor U35277 (N_35277,N_32042,N_32393);
nand U35278 (N_35278,N_30945,N_33583);
or U35279 (N_35279,N_31235,N_30519);
and U35280 (N_35280,N_30702,N_30684);
and U35281 (N_35281,N_33401,N_30254);
and U35282 (N_35282,N_30588,N_30989);
nor U35283 (N_35283,N_31304,N_30112);
nor U35284 (N_35284,N_30260,N_31520);
nor U35285 (N_35285,N_32189,N_34411);
and U35286 (N_35286,N_30797,N_33155);
or U35287 (N_35287,N_31594,N_30840);
nand U35288 (N_35288,N_31979,N_32736);
and U35289 (N_35289,N_32098,N_33827);
and U35290 (N_35290,N_33923,N_30038);
nor U35291 (N_35291,N_32425,N_30590);
xnor U35292 (N_35292,N_30884,N_33684);
or U35293 (N_35293,N_31789,N_31365);
or U35294 (N_35294,N_33800,N_33164);
nor U35295 (N_35295,N_30486,N_33280);
or U35296 (N_35296,N_31959,N_33467);
nand U35297 (N_35297,N_34500,N_34230);
nor U35298 (N_35298,N_33222,N_34289);
or U35299 (N_35299,N_30452,N_32220);
xnor U35300 (N_35300,N_34112,N_30614);
nor U35301 (N_35301,N_32862,N_30360);
nor U35302 (N_35302,N_32063,N_34396);
nand U35303 (N_35303,N_33752,N_34418);
nor U35304 (N_35304,N_31795,N_32871);
nand U35305 (N_35305,N_33038,N_32519);
nand U35306 (N_35306,N_31517,N_31278);
nor U35307 (N_35307,N_30266,N_31097);
or U35308 (N_35308,N_30763,N_34173);
nor U35309 (N_35309,N_30513,N_32313);
and U35310 (N_35310,N_30502,N_30799);
and U35311 (N_35311,N_31290,N_34082);
and U35312 (N_35312,N_34088,N_30210);
or U35313 (N_35313,N_33122,N_34638);
or U35314 (N_35314,N_31987,N_31913);
xnor U35315 (N_35315,N_34549,N_33434);
nor U35316 (N_35316,N_32556,N_30440);
xor U35317 (N_35317,N_30379,N_34513);
nor U35318 (N_35318,N_34398,N_32274);
xnor U35319 (N_35319,N_30794,N_32833);
nor U35320 (N_35320,N_31843,N_34137);
nor U35321 (N_35321,N_34461,N_33430);
nand U35322 (N_35322,N_34470,N_31175);
and U35323 (N_35323,N_33349,N_30025);
xor U35324 (N_35324,N_34576,N_33621);
and U35325 (N_35325,N_33409,N_31138);
xnor U35326 (N_35326,N_34526,N_34387);
nand U35327 (N_35327,N_32316,N_34509);
and U35328 (N_35328,N_34486,N_30972);
and U35329 (N_35329,N_34992,N_34503);
and U35330 (N_35330,N_34480,N_31276);
or U35331 (N_35331,N_33186,N_32832);
or U35332 (N_35332,N_34189,N_30725);
nor U35333 (N_35333,N_33877,N_31726);
nor U35334 (N_35334,N_33323,N_34856);
xor U35335 (N_35335,N_32375,N_34204);
xnor U35336 (N_35336,N_31983,N_31412);
or U35337 (N_35337,N_33489,N_30350);
or U35338 (N_35338,N_32594,N_32961);
xnor U35339 (N_35339,N_30324,N_30571);
and U35340 (N_35340,N_33573,N_32608);
nor U35341 (N_35341,N_31919,N_31317);
or U35342 (N_35342,N_30784,N_32447);
xor U35343 (N_35343,N_31149,N_32191);
nand U35344 (N_35344,N_32287,N_30868);
or U35345 (N_35345,N_31375,N_33839);
xnor U35346 (N_35346,N_30196,N_33979);
xnor U35347 (N_35347,N_34399,N_32217);
xor U35348 (N_35348,N_33090,N_33492);
nand U35349 (N_35349,N_33883,N_33807);
xnor U35350 (N_35350,N_34831,N_33441);
nand U35351 (N_35351,N_34401,N_34711);
nor U35352 (N_35352,N_31039,N_30804);
and U35353 (N_35353,N_32759,N_34249);
nor U35354 (N_35354,N_33638,N_31285);
nor U35355 (N_35355,N_30339,N_30123);
nor U35356 (N_35356,N_34803,N_30830);
nor U35357 (N_35357,N_31240,N_33664);
xor U35358 (N_35358,N_32889,N_34652);
or U35359 (N_35359,N_34824,N_34309);
and U35360 (N_35360,N_33983,N_34848);
and U35361 (N_35361,N_31347,N_34682);
and U35362 (N_35362,N_34057,N_33015);
xor U35363 (N_35363,N_32900,N_30561);
xor U35364 (N_35364,N_34643,N_34436);
xnor U35365 (N_35365,N_32605,N_33667);
and U35366 (N_35366,N_34471,N_30438);
or U35367 (N_35367,N_32482,N_32369);
and U35368 (N_35368,N_32811,N_30831);
or U35369 (N_35369,N_31732,N_34458);
nor U35370 (N_35370,N_31561,N_30462);
and U35371 (N_35371,N_33951,N_33420);
nand U35372 (N_35372,N_33639,N_31576);
xor U35373 (N_35373,N_34852,N_34004);
nor U35374 (N_35374,N_33209,N_32764);
nor U35375 (N_35375,N_32481,N_32859);
nand U35376 (N_35376,N_33009,N_33310);
xor U35377 (N_35377,N_30174,N_30366);
xnor U35378 (N_35378,N_31659,N_30180);
xor U35379 (N_35379,N_30008,N_30669);
xor U35380 (N_35380,N_34699,N_31848);
or U35381 (N_35381,N_32935,N_33865);
nand U35382 (N_35382,N_31163,N_32861);
and U35383 (N_35383,N_31297,N_30036);
nor U35384 (N_35384,N_31606,N_34322);
and U35385 (N_35385,N_30742,N_34523);
and U35386 (N_35386,N_30481,N_30259);
xnor U35387 (N_35387,N_32789,N_32937);
nand U35388 (N_35388,N_32568,N_31064);
and U35389 (N_35389,N_33036,N_34672);
nor U35390 (N_35390,N_33867,N_30593);
nand U35391 (N_35391,N_33647,N_32491);
and U35392 (N_35392,N_31143,N_33890);
nand U35393 (N_35393,N_33277,N_31464);
and U35394 (N_35394,N_31809,N_33833);
nor U35395 (N_35395,N_32579,N_33471);
or U35396 (N_35396,N_32279,N_32921);
xor U35397 (N_35397,N_31268,N_30068);
nor U35398 (N_35398,N_33650,N_31676);
xor U35399 (N_35399,N_34562,N_30131);
nand U35400 (N_35400,N_34352,N_34290);
xnor U35401 (N_35401,N_33738,N_31085);
nor U35402 (N_35402,N_33893,N_30160);
and U35403 (N_35403,N_34060,N_30060);
or U35404 (N_35404,N_31372,N_31955);
or U35405 (N_35405,N_31535,N_32896);
and U35406 (N_35406,N_34383,N_31150);
and U35407 (N_35407,N_32975,N_34530);
nor U35408 (N_35408,N_34431,N_33936);
nor U35409 (N_35409,N_30585,N_32638);
and U35410 (N_35410,N_32708,N_31119);
nand U35411 (N_35411,N_31626,N_30139);
nand U35412 (N_35412,N_31228,N_32293);
xnor U35413 (N_35413,N_34039,N_34937);
and U35414 (N_35414,N_32229,N_30120);
xnor U35415 (N_35415,N_32051,N_31884);
nor U35416 (N_35416,N_34242,N_31349);
or U35417 (N_35417,N_34633,N_30337);
xnor U35418 (N_35418,N_30300,N_32744);
or U35419 (N_35419,N_34495,N_32301);
xnor U35420 (N_35420,N_33544,N_34164);
nor U35421 (N_35421,N_32350,N_31473);
or U35422 (N_35422,N_32496,N_33949);
and U35423 (N_35423,N_34297,N_33075);
nand U35424 (N_35424,N_34656,N_32050);
nand U35425 (N_35425,N_31161,N_34694);
nand U35426 (N_35426,N_30331,N_30785);
or U35427 (N_35427,N_32650,N_31804);
or U35428 (N_35428,N_33924,N_31643);
nor U35429 (N_35429,N_31010,N_34560);
and U35430 (N_35430,N_33595,N_34813);
xnor U35431 (N_35431,N_32980,N_31842);
or U35432 (N_35432,N_33552,N_34913);
xor U35433 (N_35433,N_32403,N_32441);
xor U35434 (N_35434,N_30236,N_32891);
nor U35435 (N_35435,N_31373,N_31045);
and U35436 (N_35436,N_31390,N_33727);
nor U35437 (N_35437,N_31735,N_33095);
nor U35438 (N_35438,N_34333,N_31357);
nand U35439 (N_35439,N_33754,N_30740);
nor U35440 (N_35440,N_30611,N_31429);
and U35441 (N_35441,N_30741,N_32881);
nor U35442 (N_35442,N_31811,N_33618);
nand U35443 (N_35443,N_34104,N_31169);
and U35444 (N_35444,N_30143,N_30334);
xnor U35445 (N_35445,N_34499,N_32544);
or U35446 (N_35446,N_32012,N_32732);
or U35447 (N_35447,N_34712,N_33596);
nand U35448 (N_35448,N_30177,N_33985);
nand U35449 (N_35449,N_32419,N_33452);
xor U35450 (N_35450,N_32911,N_33410);
nand U35451 (N_35451,N_33926,N_33499);
and U35452 (N_35452,N_30354,N_33637);
and U35453 (N_35453,N_32267,N_33619);
xnor U35454 (N_35454,N_33555,N_30495);
or U35455 (N_35455,N_33783,N_33320);
xor U35456 (N_35456,N_32254,N_31435);
nand U35457 (N_35457,N_33760,N_31513);
or U35458 (N_35458,N_33750,N_33005);
xnor U35459 (N_35459,N_33468,N_33540);
nor U35460 (N_35460,N_30432,N_31430);
and U35461 (N_35461,N_31403,N_30826);
nor U35462 (N_35462,N_32632,N_30140);
nor U35463 (N_35463,N_32039,N_34654);
or U35464 (N_35464,N_32826,N_34919);
nand U35465 (N_35465,N_31459,N_33763);
and U35466 (N_35466,N_32726,N_34832);
nand U35467 (N_35467,N_31094,N_34338);
nor U35468 (N_35468,N_31727,N_34202);
nor U35469 (N_35469,N_34556,N_33538);
nor U35470 (N_35470,N_32629,N_30488);
nand U35471 (N_35471,N_34955,N_32917);
and U35472 (N_35472,N_33549,N_31530);
or U35473 (N_35473,N_34328,N_32406);
nor U35474 (N_35474,N_32772,N_32684);
or U35475 (N_35475,N_34724,N_33382);
nor U35476 (N_35476,N_33136,N_33478);
nor U35477 (N_35477,N_30245,N_34648);
or U35478 (N_35478,N_32927,N_32232);
nand U35479 (N_35479,N_33318,N_31545);
or U35480 (N_35480,N_30936,N_31052);
nor U35481 (N_35481,N_30621,N_32719);
nor U35482 (N_35482,N_33243,N_33086);
nor U35483 (N_35483,N_34928,N_31259);
nor U35484 (N_35484,N_33212,N_32758);
nand U35485 (N_35485,N_33972,N_33021);
and U35486 (N_35486,N_33421,N_30534);
nand U35487 (N_35487,N_32342,N_34018);
or U35488 (N_35488,N_30610,N_32863);
nand U35489 (N_35489,N_34402,N_31216);
nand U35490 (N_35490,N_32384,N_33774);
and U35491 (N_35491,N_33915,N_31076);
xor U35492 (N_35492,N_33679,N_31592);
nor U35493 (N_35493,N_32427,N_30887);
nand U35494 (N_35494,N_32703,N_33119);
nor U35495 (N_35495,N_31493,N_31650);
nand U35496 (N_35496,N_30708,N_30943);
nand U35497 (N_35497,N_33143,N_33987);
nand U35498 (N_35498,N_30650,N_33881);
xnor U35499 (N_35499,N_30253,N_32565);
nand U35500 (N_35500,N_30662,N_31311);
nand U35501 (N_35501,N_31053,N_34540);
and U35502 (N_35502,N_31289,N_34762);
and U35503 (N_35503,N_31210,N_32751);
nand U35504 (N_35504,N_30711,N_30490);
nand U35505 (N_35505,N_30320,N_34002);
xnor U35506 (N_35506,N_31827,N_34533);
nand U35507 (N_35507,N_33715,N_31497);
nand U35508 (N_35508,N_31857,N_33680);
and U35509 (N_35509,N_32094,N_30391);
or U35510 (N_35510,N_30216,N_34370);
nand U35511 (N_35511,N_31091,N_34915);
xor U35512 (N_35512,N_30498,N_30387);
nor U35513 (N_35513,N_32540,N_30398);
xor U35514 (N_35514,N_31845,N_30511);
nor U35515 (N_35515,N_33747,N_34122);
nand U35516 (N_35516,N_32134,N_32381);
nand U35517 (N_35517,N_34572,N_32597);
xor U35518 (N_35518,N_31771,N_33001);
nand U35519 (N_35519,N_33894,N_34072);
nand U35520 (N_35520,N_30649,N_33537);
nand U35521 (N_35521,N_33878,N_33511);
xnor U35522 (N_35522,N_33837,N_32144);
or U35523 (N_35523,N_31486,N_30834);
or U35524 (N_35524,N_34679,N_31651);
or U35525 (N_35525,N_34688,N_33608);
nor U35526 (N_35526,N_34885,N_33686);
nand U35527 (N_35527,N_32551,N_31538);
nand U35528 (N_35528,N_33567,N_34988);
nand U35529 (N_35529,N_33474,N_33539);
nor U35530 (N_35530,N_31057,N_31168);
nand U35531 (N_35531,N_34449,N_30762);
nand U35532 (N_35532,N_32129,N_31005);
and U35533 (N_35533,N_32954,N_33901);
and U35534 (N_35534,N_30756,N_30549);
nand U35535 (N_35535,N_32665,N_30019);
nor U35536 (N_35536,N_30414,N_34916);
and U35537 (N_35537,N_31377,N_32331);
xnor U35538 (N_35538,N_31019,N_32052);
xor U35539 (N_35539,N_32930,N_31223);
xnor U35540 (N_35540,N_32345,N_32204);
or U35541 (N_35541,N_30507,N_32062);
xnor U35542 (N_35542,N_33734,N_32691);
xnor U35543 (N_35543,N_34896,N_34751);
or U35544 (N_35544,N_33981,N_30920);
nand U35545 (N_35545,N_34178,N_33518);
xor U35546 (N_35546,N_33272,N_30125);
xor U35547 (N_35547,N_32309,N_34281);
xnor U35548 (N_35548,N_34140,N_32260);
or U35549 (N_35549,N_34594,N_34769);
xor U35550 (N_35550,N_34849,N_30359);
nand U35551 (N_35551,N_33742,N_32497);
nand U35552 (N_35552,N_32243,N_31523);
and U35553 (N_35553,N_33241,N_32509);
nor U35554 (N_35554,N_32268,N_33292);
xnor U35555 (N_35555,N_33386,N_32113);
xor U35556 (N_35556,N_30773,N_30656);
xor U35557 (N_35557,N_30925,N_31639);
and U35558 (N_35558,N_32186,N_32668);
nor U35559 (N_35559,N_31399,N_32261);
and U35560 (N_35560,N_31628,N_34100);
and U35561 (N_35561,N_31963,N_30178);
nor U35562 (N_35562,N_34817,N_32308);
xor U35563 (N_35563,N_31622,N_31114);
and U35564 (N_35564,N_33034,N_33632);
and U35565 (N_35565,N_34364,N_34827);
xnor U35566 (N_35566,N_30532,N_30541);
and U35567 (N_35567,N_32068,N_31961);
and U35568 (N_35568,N_31720,N_33157);
or U35569 (N_35569,N_33289,N_34144);
nor U35570 (N_35570,N_32500,N_30000);
nor U35571 (N_35571,N_32716,N_34116);
or U35572 (N_35572,N_34303,N_31755);
nand U35573 (N_35573,N_34163,N_30793);
nand U35574 (N_35574,N_31499,N_33694);
or U35575 (N_35575,N_34834,N_32009);
nand U35576 (N_35576,N_33145,N_33601);
xnor U35577 (N_35577,N_30394,N_33308);
and U35578 (N_35578,N_33263,N_34180);
or U35579 (N_35579,N_34527,N_31653);
nand U35580 (N_35580,N_31746,N_33035);
nor U35581 (N_35581,N_34330,N_31288);
nor U35582 (N_35582,N_33088,N_32956);
nand U35583 (N_35583,N_33652,N_32843);
nor U35584 (N_35584,N_30301,N_32743);
xnor U35585 (N_35585,N_31305,N_34268);
xnor U35586 (N_35586,N_34315,N_31404);
or U35587 (N_35587,N_33051,N_31171);
nand U35588 (N_35588,N_33945,N_31888);
nor U35589 (N_35589,N_33990,N_32628);
xnor U35590 (N_35590,N_34780,N_30241);
nand U35591 (N_35591,N_32215,N_34240);
or U35592 (N_35592,N_32966,N_30181);
or U35593 (N_35593,N_33098,N_34061);
nor U35594 (N_35594,N_30559,N_31871);
or U35595 (N_35595,N_30858,N_32779);
and U35596 (N_35596,N_32695,N_31930);
nand U35597 (N_35597,N_30613,N_33794);
nor U35598 (N_35598,N_30351,N_33018);
nand U35599 (N_35599,N_31761,N_34209);
nor U35600 (N_35600,N_33196,N_31753);
xnor U35601 (N_35601,N_30539,N_33640);
and U35602 (N_35602,N_33984,N_34709);
or U35603 (N_35603,N_34946,N_30377);
xor U35604 (N_35604,N_30098,N_32356);
nor U35605 (N_35605,N_32353,N_33395);
or U35606 (N_35606,N_32535,N_30715);
xnor U35607 (N_35607,N_33000,N_33602);
and U35608 (N_35608,N_33104,N_34545);
or U35609 (N_35609,N_33600,N_30892);
xnor U35610 (N_35610,N_32539,N_34037);
and U35611 (N_35611,N_32734,N_31803);
nand U35612 (N_35612,N_31693,N_30531);
xor U35613 (N_35613,N_34918,N_34464);
or U35614 (N_35614,N_34903,N_30022);
nor U35615 (N_35615,N_31371,N_31226);
or U35616 (N_35616,N_31077,N_33111);
and U35617 (N_35617,N_32456,N_32577);
nand U35618 (N_35618,N_33886,N_33536);
and U35619 (N_35619,N_31313,N_34515);
nor U35620 (N_35620,N_32033,N_31909);
and U35621 (N_35621,N_30654,N_30995);
xnor U35622 (N_35622,N_30837,N_33789);
xnor U35623 (N_35623,N_32670,N_33184);
and U35624 (N_35624,N_31394,N_32163);
nor U35625 (N_35625,N_33028,N_34858);
nor U35626 (N_35626,N_30342,N_31379);
and U35627 (N_35627,N_30256,N_32409);
nand U35628 (N_35628,N_32757,N_34508);
xnor U35629 (N_35629,N_31966,N_30453);
or U35630 (N_35630,N_34800,N_31972);
or U35631 (N_35631,N_33108,N_34029);
nor U35632 (N_35632,N_34273,N_31041);
nand U35633 (N_35633,N_30933,N_30333);
nor U35634 (N_35634,N_33698,N_32263);
or U35635 (N_35635,N_34054,N_31968);
nor U35636 (N_35636,N_31179,N_34959);
nor U35637 (N_35637,N_34481,N_34138);
xor U35638 (N_35638,N_33436,N_32960);
nand U35639 (N_35639,N_30619,N_31668);
xor U35640 (N_35640,N_34855,N_30202);
nand U35641 (N_35641,N_33485,N_31496);
xnor U35642 (N_35642,N_33233,N_32355);
nand U35643 (N_35643,N_34747,N_30718);
xor U35644 (N_35644,N_33778,N_30317);
or U35645 (N_35645,N_31176,N_30020);
xor U35646 (N_35646,N_30460,N_32501);
nor U35647 (N_35647,N_33071,N_34256);
nor U35648 (N_35648,N_33317,N_33362);
or U35649 (N_35649,N_33373,N_30921);
nor U35650 (N_35650,N_31648,N_34270);
nand U35651 (N_35651,N_30171,N_34695);
nor U35652 (N_35652,N_30661,N_30319);
nand U35653 (N_35653,N_33414,N_34894);
xor U35654 (N_35654,N_33156,N_32173);
or U35655 (N_35655,N_33857,N_33592);
nand U35656 (N_35656,N_34176,N_34231);
nand U35657 (N_35657,N_30912,N_33958);
nand U35658 (N_35658,N_31024,N_30062);
and U35659 (N_35659,N_32193,N_32445);
and U35660 (N_35660,N_33896,N_31136);
and U35661 (N_35661,N_33187,N_33235);
xor U35662 (N_35662,N_30581,N_33882);
or U35663 (N_35663,N_32346,N_31718);
and U35664 (N_35664,N_31604,N_30105);
nor U35665 (N_35665,N_32344,N_34390);
or U35666 (N_35666,N_30698,N_34733);
nand U35667 (N_35667,N_32547,N_33293);
xor U35668 (N_35668,N_30609,N_32226);
nand U35669 (N_35669,N_32814,N_30451);
nor U35670 (N_35670,N_30117,N_31237);
nand U35671 (N_35671,N_32784,N_32016);
nand U35672 (N_35672,N_32775,N_30122);
or U35673 (N_35673,N_32778,N_31605);
and U35674 (N_35674,N_34141,N_34437);
or U35675 (N_35675,N_30355,N_34748);
nand U35676 (N_35676,N_34577,N_34292);
xnor U35677 (N_35677,N_34317,N_33513);
nand U35678 (N_35678,N_31725,N_31870);
or U35679 (N_35679,N_30908,N_31386);
and U35680 (N_35680,N_30510,N_33975);
and U35681 (N_35681,N_33027,N_31935);
and U35682 (N_35682,N_31976,N_30124);
nor U35683 (N_35683,N_33026,N_33043);
or U35684 (N_35684,N_30263,N_34409);
nand U35685 (N_35685,N_34797,N_34716);
and U35686 (N_35686,N_34271,N_34828);
and U35687 (N_35687,N_32792,N_32430);
xor U35688 (N_35688,N_32460,N_30448);
or U35689 (N_35689,N_30284,N_32643);
and U35690 (N_35690,N_34047,N_32932);
nor U35691 (N_35691,N_34543,N_32208);
xor U35692 (N_35692,N_32252,N_32379);
or U35693 (N_35693,N_30153,N_33307);
or U35694 (N_35694,N_34941,N_31184);
xor U35695 (N_35695,N_33710,N_32449);
xor U35696 (N_35696,N_34227,N_31841);
and U35697 (N_35697,N_31865,N_31340);
or U35698 (N_35698,N_32787,N_31710);
and U35699 (N_35699,N_30110,N_32877);
or U35700 (N_35700,N_33671,N_32587);
nand U35701 (N_35701,N_32442,N_31768);
xor U35702 (N_35702,N_31116,N_33493);
nand U35703 (N_35703,N_30003,N_33246);
and U35704 (N_35704,N_31553,N_31687);
and U35705 (N_35705,N_34195,N_34835);
nand U35706 (N_35706,N_33695,N_34717);
nand U35707 (N_35707,N_31344,N_33301);
xnor U35708 (N_35708,N_34977,N_30968);
xor U35709 (N_35709,N_30631,N_34705);
xnor U35710 (N_35710,N_34637,N_30618);
or U35711 (N_35711,N_33213,N_30280);
nand U35712 (N_35712,N_32253,N_32654);
xor U35713 (N_35713,N_32297,N_33804);
or U35714 (N_35714,N_34220,N_30094);
nand U35715 (N_35715,N_33054,N_30937);
and U35716 (N_35716,N_32221,N_31234);
and U35717 (N_35717,N_31819,N_31446);
or U35718 (N_35718,N_33988,N_33190);
nor U35719 (N_35719,N_32682,N_34435);
and U35720 (N_35720,N_34430,N_30466);
or U35721 (N_35721,N_33643,N_32008);
and U35722 (N_35722,N_31462,N_34089);
and U35723 (N_35723,N_34779,N_30053);
nand U35724 (N_35724,N_32056,N_34062);
nor U35725 (N_35725,N_34578,N_33131);
or U35726 (N_35726,N_30712,N_34969);
and U35727 (N_35727,N_30031,N_30230);
xor U35728 (N_35728,N_31301,N_34492);
and U35729 (N_35729,N_34377,N_31338);
nor U35730 (N_35730,N_34601,N_32195);
xnor U35731 (N_35731,N_32976,N_34968);
xnor U35732 (N_35732,N_32123,N_32328);
nand U35733 (N_35733,N_33058,N_34902);
and U35734 (N_35734,N_33699,N_32371);
xor U35735 (N_35735,N_30288,N_33279);
or U35736 (N_35736,N_30012,N_31992);
nand U35737 (N_35737,N_33971,N_31656);
or U35738 (N_35738,N_31514,N_31418);
nor U35739 (N_35739,N_30808,N_31914);
nand U35740 (N_35740,N_30189,N_31990);
nand U35741 (N_35741,N_31111,N_34252);
and U35742 (N_35742,N_33953,N_30988);
nand U35743 (N_35743,N_30332,N_31941);
or U35744 (N_35744,N_34161,N_33831);
and U35745 (N_35745,N_30034,N_32166);
xor U35746 (N_35746,N_34685,N_30949);
nand U35747 (N_35747,N_32656,N_30580);
nand U35748 (N_35748,N_32766,N_33125);
xor U35749 (N_35749,N_31790,N_31443);
xnor U35750 (N_35750,N_30059,N_31054);
xnor U35751 (N_35751,N_30602,N_34978);
nor U35752 (N_35752,N_34280,N_30184);
or U35753 (N_35753,N_30258,N_30166);
nand U35754 (N_35754,N_32282,N_30419);
or U35755 (N_35755,N_30417,N_30900);
xor U35756 (N_35756,N_32079,N_34706);
nand U35757 (N_35757,N_31448,N_32503);
or U35758 (N_35758,N_31434,N_30727);
nand U35759 (N_35759,N_33462,N_33245);
or U35760 (N_35760,N_34279,N_30413);
nor U35761 (N_35761,N_31230,N_34032);
nand U35762 (N_35762,N_33655,N_33050);
and U35763 (N_35763,N_30576,N_34455);
nand U35764 (N_35764,N_34113,N_33037);
or U35765 (N_35765,N_33264,N_32043);
xor U35766 (N_35766,N_31944,N_31723);
or U35767 (N_35767,N_32617,N_30897);
and U35768 (N_35768,N_34547,N_32159);
xnor U35769 (N_35769,N_32731,N_32972);
nor U35770 (N_35770,N_30876,N_34498);
or U35771 (N_35771,N_32169,N_32785);
or U35772 (N_35772,N_30044,N_33966);
or U35773 (N_35773,N_34561,N_33525);
xor U35774 (N_35774,N_32616,N_30090);
nand U35775 (N_35775,N_32663,N_33957);
nand U35776 (N_35776,N_30169,N_34384);
and U35777 (N_35777,N_32323,N_31655);
xnor U35778 (N_35778,N_30399,N_30294);
xor U35779 (N_35779,N_33588,N_33316);
nor U35780 (N_35780,N_33351,N_31355);
nand U35781 (N_35781,N_31970,N_33249);
or U35782 (N_35782,N_33048,N_33121);
and U35783 (N_35783,N_31170,N_31610);
and U35784 (N_35784,N_31636,N_34241);
nand U35785 (N_35785,N_31996,N_31534);
nand U35786 (N_35786,N_30268,N_33117);
nand U35787 (N_35787,N_31391,N_33466);
or U35788 (N_35788,N_30278,N_34901);
and U35789 (N_35789,N_34584,N_31783);
or U35790 (N_35790,N_31118,N_32566);
nand U35791 (N_35791,N_33404,N_30318);
nand U35792 (N_35792,N_33319,N_34267);
and U35793 (N_35793,N_33268,N_33597);
nor U35794 (N_35794,N_33675,N_31033);
nor U35795 (N_35795,N_30052,N_32652);
nand U35796 (N_35796,N_34448,N_31563);
nor U35797 (N_35797,N_33653,N_30429);
nand U35798 (N_35798,N_33908,N_31046);
nor U35799 (N_35799,N_31547,N_32435);
nand U35800 (N_35800,N_34316,N_32883);
and U35801 (N_35801,N_32710,N_34276);
nor U35802 (N_35802,N_34446,N_32439);
and U35803 (N_35803,N_32755,N_34980);
nand U35804 (N_35804,N_32394,N_33817);
nand U35805 (N_35805,N_30182,N_34045);
xnor U35806 (N_35806,N_34356,N_31717);
xor U35807 (N_35807,N_32518,N_32351);
nor U35808 (N_35808,N_34056,N_31000);
nor U35809 (N_35809,N_31021,N_31048);
xor U35810 (N_35810,N_34111,N_30776);
xnor U35811 (N_35811,N_33851,N_31779);
nor U35812 (N_35812,N_32687,N_33764);
or U35813 (N_35813,N_30009,N_32300);
and U35814 (N_35814,N_33944,N_33146);
or U35815 (N_35815,N_34985,N_31569);
or U35816 (N_35816,N_32291,N_34704);
or U35817 (N_35817,N_30786,N_30601);
and U35818 (N_35818,N_30929,N_33589);
xnor U35819 (N_35819,N_31812,N_33267);
nand U35820 (N_35820,N_34160,N_31907);
and U35821 (N_35821,N_31844,N_31225);
nor U35822 (N_35822,N_31549,N_31642);
xnor U35823 (N_35823,N_34781,N_31825);
nand U35824 (N_35824,N_30365,N_30130);
or U35825 (N_35825,N_32157,N_32470);
and U35826 (N_35826,N_33665,N_34732);
nor U35827 (N_35827,N_30475,N_31784);
nand U35828 (N_35828,N_30520,N_30129);
nand U35829 (N_35829,N_32283,N_34358);
nand U35830 (N_35830,N_34564,N_34759);
or U35831 (N_35831,N_30273,N_34865);
and U35832 (N_35832,N_30723,N_32690);
and U35833 (N_35833,N_33083,N_31369);
xnor U35834 (N_35834,N_30341,N_33868);
and U35835 (N_35835,N_30251,N_30085);
nand U35836 (N_35836,N_34691,N_33194);
nand U35837 (N_35837,N_32846,N_31927);
and U35838 (N_35838,N_34166,N_33457);
nor U35839 (N_35839,N_31599,N_34342);
or U35840 (N_35840,N_31837,N_31543);
xnor U35841 (N_35841,N_33389,N_33355);
nor U35842 (N_35842,N_34191,N_31479);
xnor U35843 (N_35843,N_31020,N_31946);
or U35844 (N_35844,N_32841,N_31095);
or U35845 (N_35845,N_32943,N_33483);
xor U35846 (N_35846,N_34871,N_30223);
or U35847 (N_35847,N_30390,N_31529);
nand U35848 (N_35848,N_33284,N_30078);
and U35849 (N_35849,N_31861,N_34211);
nand U35850 (N_35850,N_32400,N_31765);
nor U35851 (N_35851,N_30045,N_32604);
nand U35852 (N_35852,N_31608,N_32963);
and U35853 (N_35853,N_31902,N_33342);
nor U35854 (N_35854,N_32135,N_33123);
and U35855 (N_35855,N_31703,N_31358);
nor U35856 (N_35856,N_30295,N_32924);
and U35857 (N_35857,N_33746,N_32359);
nor U35858 (N_35858,N_34067,N_31840);
xnor U35859 (N_35859,N_30227,N_30821);
or U35860 (N_35860,N_30942,N_32181);
nor U35861 (N_35861,N_31915,N_30567);
nand U35862 (N_35862,N_33714,N_32512);
nand U35863 (N_35863,N_31879,N_33010);
and U35864 (N_35864,N_33056,N_34375);
and U35865 (N_35865,N_30418,N_32874);
nor U35866 (N_35866,N_34947,N_30097);
xnor U35867 (N_35867,N_34617,N_31912);
xnor U35868 (N_35868,N_31986,N_31425);
nor U35869 (N_35869,N_32101,N_31954);
xnor U35870 (N_35870,N_32630,N_34063);
nor U35871 (N_35871,N_32360,N_34319);
or U35872 (N_35872,N_33161,N_34608);
nor U35873 (N_35873,N_33559,N_32842);
nand U35874 (N_35874,N_30856,N_32315);
and U35875 (N_35875,N_30370,N_30403);
or U35876 (N_35876,N_31058,N_31433);
nor U35877 (N_35877,N_34199,N_32809);
and U35878 (N_35878,N_30724,N_32914);
xor U35879 (N_35879,N_32310,N_31669);
and U35880 (N_35880,N_30582,N_31332);
nand U35881 (N_35881,N_30575,N_32474);
nor U35882 (N_35882,N_33068,N_30546);
or U35883 (N_35883,N_32388,N_31082);
and U35884 (N_35884,N_30924,N_32184);
and U35885 (N_35885,N_31273,N_31588);
nor U35886 (N_35886,N_30881,N_34982);
nor U35887 (N_35887,N_33598,N_33135);
nor U35888 (N_35888,N_34700,N_30563);
or U35889 (N_35889,N_34049,N_34571);
nand U35890 (N_35890,N_33751,N_31485);
nor U35891 (N_35891,N_31885,N_32669);
or U35892 (N_35892,N_31447,N_31333);
and U35893 (N_35893,N_34641,N_30233);
nor U35894 (N_35894,N_30969,N_30806);
nor U35895 (N_35895,N_34809,N_31194);
nand U35896 (N_35896,N_34840,N_30485);
nand U35897 (N_35897,N_33889,N_30693);
and U35898 (N_35898,N_33723,N_34555);
nand U35899 (N_35899,N_33189,N_30822);
xnor U35900 (N_35900,N_32156,N_32377);
and U35901 (N_35901,N_34071,N_32055);
or U35902 (N_35902,N_34592,N_33482);
or U35903 (N_35903,N_32655,N_30849);
nor U35904 (N_35904,N_32017,N_30516);
nand U35905 (N_35905,N_30796,N_30226);
or U35906 (N_35906,N_30091,N_33892);
and U35907 (N_35907,N_34190,N_34812);
nor U35908 (N_35908,N_33480,N_33059);
or U35909 (N_35909,N_32907,N_32203);
nor U35910 (N_35910,N_30905,N_32959);
xnor U35911 (N_35911,N_32599,N_34811);
or U35912 (N_35912,N_33603,N_31908);
or U35913 (N_35913,N_32165,N_33885);
or U35914 (N_35914,N_31453,N_32092);
nor U35915 (N_35915,N_30246,N_31186);
or U35916 (N_35916,N_32213,N_33276);
and U35917 (N_35917,N_32830,N_30205);
xnor U35918 (N_35918,N_33238,N_31619);
xnor U35919 (N_35919,N_34467,N_33053);
and U35920 (N_35920,N_30573,N_33286);
nor U35921 (N_35921,N_32378,N_30745);
or U35922 (N_35922,N_34559,N_33031);
and U35923 (N_35923,N_34320,N_31734);
and U35924 (N_35924,N_30863,N_34354);
and U35925 (N_35925,N_34906,N_30454);
nand U35926 (N_35926,N_33825,N_32086);
nor U35927 (N_35927,N_33174,N_30750);
or U35928 (N_35928,N_31793,N_30314);
nor U35929 (N_35929,N_33508,N_30896);
xnor U35930 (N_35930,N_32170,N_33100);
nor U35931 (N_35931,N_31140,N_34531);
nor U35932 (N_35932,N_30073,N_30710);
nand U35933 (N_35933,N_34395,N_34891);
and U35934 (N_35934,N_31878,N_31707);
or U35935 (N_35935,N_31475,N_30274);
and U35936 (N_35936,N_34441,N_31519);
or U35937 (N_35937,N_34912,N_34251);
xor U35938 (N_35938,N_33960,N_30835);
xnor U35939 (N_35939,N_34616,N_30063);
or U35940 (N_35940,N_32882,N_33534);
nand U35941 (N_35941,N_31892,N_33777);
xor U35942 (N_35942,N_32367,N_31900);
nand U35943 (N_35943,N_33663,N_30474);
and U35944 (N_35944,N_32969,N_32866);
xor U35945 (N_35945,N_34728,N_33884);
and U35946 (N_35946,N_32754,N_30380);
or U35947 (N_35947,N_31994,N_33935);
nand U35948 (N_35948,N_32110,N_34185);
nand U35949 (N_35949,N_32197,N_34629);
nand U35950 (N_35950,N_30688,N_33315);
xor U35951 (N_35951,N_32953,N_30281);
nor U35952 (N_35952,N_34768,N_34542);
xnor U35953 (N_35953,N_30190,N_30759);
and U35954 (N_35954,N_33367,N_31255);
nand U35955 (N_35955,N_33669,N_34940);
and U35956 (N_35956,N_31488,N_30569);
and U35957 (N_35957,N_33625,N_30412);
nor U35958 (N_35958,N_32521,N_30628);
nor U35959 (N_35959,N_30517,N_32750);
and U35960 (N_35960,N_34099,N_31440);
nor U35961 (N_35961,N_34822,N_30766);
xnor U35962 (N_35962,N_31201,N_32515);
xnor U35963 (N_35963,N_34611,N_31595);
or U35964 (N_35964,N_30570,N_34727);
or U35965 (N_35965,N_34948,N_33458);
nand U35966 (N_35966,N_34749,N_34225);
or U35967 (N_35967,N_32918,N_34110);
and U35968 (N_35968,N_30598,N_34146);
and U35969 (N_35969,N_33770,N_33560);
and U35970 (N_35970,N_32443,N_30634);
nand U35971 (N_35971,N_33756,N_30716);
nor U35972 (N_35972,N_32251,N_32609);
nor U35973 (N_35973,N_30551,N_34607);
or U35974 (N_35974,N_31299,N_31056);
and U35975 (N_35975,N_30299,N_32305);
xnor U35976 (N_35976,N_30389,N_31193);
nand U35977 (N_35977,N_30501,N_30603);
nor U35978 (N_35978,N_30705,N_32702);
and U35979 (N_35979,N_30018,N_30838);
xnor U35980 (N_35980,N_34888,N_30816);
nand U35981 (N_35981,N_34790,N_34986);
nor U35982 (N_35982,N_30687,N_30704);
or U35983 (N_35983,N_30671,N_34754);
nor U35984 (N_35984,N_32525,N_32909);
nand U35985 (N_35985,N_31763,N_30158);
xor U35986 (N_35986,N_34307,N_30807);
xor U35987 (N_35987,N_32014,N_32677);
nand U35988 (N_35988,N_31199,N_34598);
nor U35989 (N_35989,N_32973,N_34960);
nand U35990 (N_35990,N_32089,N_32770);
nand U35991 (N_35991,N_31736,N_30304);
and U35992 (N_35992,N_30014,N_30410);
nor U35993 (N_35993,N_33644,N_33469);
nand U35994 (N_35994,N_30478,N_34566);
or U35995 (N_35995,N_30480,N_31880);
nand U35996 (N_35996,N_33919,N_31702);
or U35997 (N_35997,N_31353,N_30686);
and U35998 (N_35998,N_34213,N_32389);
and U35999 (N_35999,N_33787,N_30220);
xnor U36000 (N_36000,N_32520,N_30447);
or U36001 (N_36001,N_33941,N_32723);
nand U36002 (N_36002,N_32459,N_31366);
xnor U36003 (N_36003,N_31901,N_33842);
or U36004 (N_36004,N_34485,N_30967);
or U36005 (N_36005,N_32502,N_33442);
and U36006 (N_36006,N_32292,N_34838);
or U36007 (N_36007,N_32307,N_30335);
or U36008 (N_36008,N_31115,N_32196);
nor U36009 (N_36009,N_32250,N_32828);
or U36010 (N_36010,N_33530,N_30733);
nand U36011 (N_36011,N_30970,N_33464);
or U36012 (N_36012,N_33278,N_34102);
xnor U36013 (N_36013,N_30188,N_34836);
and U36014 (N_36014,N_32555,N_32096);
nor U36015 (N_36015,N_33562,N_32678);
xnor U36016 (N_36016,N_30780,N_30683);
nor U36017 (N_36017,N_31167,N_30142);
nor U36018 (N_36018,N_34782,N_31612);
nor U36019 (N_36019,N_32249,N_34841);
and U36020 (N_36020,N_30867,N_34009);
nor U36021 (N_36021,N_30037,N_31183);
xor U36022 (N_36022,N_33215,N_31999);
xor U36023 (N_36023,N_31350,N_34134);
xnor U36024 (N_36024,N_33939,N_31778);
xor U36025 (N_36025,N_32281,N_33326);
and U36026 (N_36026,N_30811,N_32132);
nand U36027 (N_36027,N_34407,N_32709);
and U36028 (N_36028,N_32745,N_34802);
and U36029 (N_36029,N_34157,N_32090);
and U36030 (N_36030,N_30956,N_31920);
xor U36031 (N_36031,N_33353,N_31466);
nand U36032 (N_36032,N_32962,N_32200);
nor U36033 (N_36033,N_30352,N_30470);
xnor U36034 (N_36034,N_31202,N_33938);
nor U36035 (N_36035,N_32484,N_30302);
nor U36036 (N_36036,N_32153,N_32207);
nor U36037 (N_36037,N_31719,N_32126);
xnor U36038 (N_36038,N_30874,N_31133);
xor U36039 (N_36039,N_34014,N_30810);
and U36040 (N_36040,N_32533,N_30529);
xor U36041 (N_36041,N_30678,N_34169);
and U36042 (N_36042,N_34510,N_33689);
nand U36043 (N_36043,N_30548,N_30664);
xnor U36044 (N_36044,N_33265,N_32432);
xor U36045 (N_36045,N_30675,N_32155);
and U36046 (N_36046,N_33986,N_32799);
xnor U36047 (N_36047,N_33620,N_34019);
or U36048 (N_36048,N_31112,N_32450);
nand U36049 (N_36049,N_32906,N_32644);
and U36050 (N_36050,N_30537,N_32602);
xor U36051 (N_36051,N_34810,N_31739);
and U36052 (N_36052,N_30163,N_30940);
xor U36053 (N_36053,N_32855,N_34143);
nand U36054 (N_36054,N_31756,N_31750);
nor U36055 (N_36055,N_30552,N_34675);
nor U36056 (N_36056,N_31195,N_32240);
and U36057 (N_36057,N_31733,N_33580);
and U36058 (N_36058,N_31188,N_34433);
xnor U36059 (N_36059,N_34587,N_32718);
nor U36060 (N_36060,N_34610,N_33927);
xnor U36061 (N_36061,N_34867,N_33973);
or U36062 (N_36062,N_34820,N_34219);
nand U36063 (N_36063,N_30409,N_33432);
nand U36064 (N_36064,N_30264,N_32685);
and U36065 (N_36065,N_32314,N_32981);
or U36066 (N_36066,N_32864,N_32680);
xnor U36067 (N_36067,N_31638,N_30629);
nand U36068 (N_36068,N_34051,N_33683);
and U36069 (N_36069,N_33294,N_33384);
or U36070 (N_36070,N_32633,N_32624);
nor U36071 (N_36071,N_33740,N_33646);
nor U36072 (N_36072,N_30102,N_32106);
or U36073 (N_36073,N_32357,N_31574);
and U36074 (N_36074,N_33855,N_30033);
nand U36075 (N_36075,N_33321,N_31402);
nor U36076 (N_36076,N_34155,N_31490);
and U36077 (N_36077,N_30591,N_33311);
nor U36078 (N_36078,N_33449,N_34424);
nand U36079 (N_36079,N_31343,N_32383);
nor U36080 (N_36080,N_34568,N_31074);
and U36081 (N_36081,N_34077,N_33744);
or U36082 (N_36082,N_30795,N_32401);
and U36083 (N_36083,N_32506,N_31457);
nor U36084 (N_36084,N_32993,N_30214);
or U36085 (N_36085,N_33312,N_34909);
nand U36086 (N_36086,N_33182,N_31585);
nand U36087 (N_36087,N_32955,N_31093);
nand U36088 (N_36088,N_31629,N_32569);
xnor U36089 (N_36089,N_31924,N_32397);
and U36090 (N_36090,N_33514,N_34482);
nand U36091 (N_36091,N_31644,N_31474);
or U36092 (N_36092,N_34286,N_30218);
or U36093 (N_36093,N_31063,N_30774);
nand U36094 (N_36094,N_34406,N_33240);
nand U36095 (N_36095,N_34171,N_32472);
xor U36096 (N_36096,N_33828,N_32015);
nor U36097 (N_36097,N_31624,N_34020);
and U36098 (N_36098,N_33419,N_33862);
nor U36099 (N_36099,N_30572,N_31762);
and U36100 (N_36100,N_34591,N_33074);
nor U36101 (N_36101,N_33343,N_31652);
nor U36102 (N_36102,N_30694,N_32020);
nor U36103 (N_36103,N_31308,N_30152);
and U36104 (N_36104,N_32464,N_32915);
or U36105 (N_36105,N_34454,N_31104);
xnor U36106 (N_36106,N_31984,N_33269);
or U36107 (N_36107,N_30221,N_33335);
nor U36108 (N_36108,N_32641,N_34504);
nand U36109 (N_36109,N_33191,N_33200);
nand U36110 (N_36110,N_34861,N_34128);
or U36111 (N_36111,N_31573,N_31824);
and U36112 (N_36112,N_30941,N_30828);
and U36113 (N_36113,N_33948,N_34521);
or U36114 (N_36114,N_34934,N_33743);
and U36115 (N_36115,N_31501,N_30058);
nor U36116 (N_36116,N_33261,N_34886);
nor U36117 (N_36117,N_30164,N_34620);
nand U36118 (N_36118,N_34973,N_33577);
nor U36119 (N_36119,N_32247,N_33627);
nand U36120 (N_36120,N_31044,N_33587);
or U36121 (N_36121,N_32696,N_31715);
nor U36122 (N_36122,N_33961,N_32034);
or U36123 (N_36123,N_32839,N_34392);
xor U36124 (N_36124,N_34927,N_34548);
xnor U36125 (N_36125,N_31309,N_33234);
xor U36126 (N_36126,N_34767,N_30035);
nand U36127 (N_36127,N_32413,N_32625);
nand U36128 (N_36128,N_33142,N_30249);
and U36129 (N_36129,N_32373,N_34325);
and U36130 (N_36130,N_34964,N_31411);
or U36131 (N_36131,N_31421,N_34823);
nor U36132 (N_36132,N_34376,N_32049);
xnor U36133 (N_36133,N_32983,N_33888);
xor U36134 (N_36134,N_31567,N_32422);
nand U36135 (N_36135,N_31780,N_34363);
or U36136 (N_36136,N_32890,N_34600);
nor U36137 (N_36137,N_33374,N_31527);
and U36138 (N_36138,N_33604,N_32108);
or U36139 (N_36139,N_32835,N_32306);
or U36140 (N_36140,N_31249,N_31988);
nor U36141 (N_36141,N_32475,N_33931);
nand U36142 (N_36142,N_30728,N_33724);
nor U36143 (N_36143,N_33999,N_33522);
nand U36144 (N_36144,N_32548,N_32595);
or U36145 (N_36145,N_33666,N_32095);
xnor U36146 (N_36146,N_34368,N_33725);
and U36147 (N_36147,N_30594,N_30367);
and U36148 (N_36148,N_31246,N_30882);
nor U36149 (N_36149,N_32908,N_34536);
or U36150 (N_36150,N_33934,N_32122);
nor U36151 (N_36151,N_31741,N_32550);
nor U36152 (N_36152,N_31009,N_32610);
xnor U36153 (N_36153,N_31387,N_33674);
and U36154 (N_36154,N_33516,N_32176);
nand U36155 (N_36155,N_31951,N_30781);
nor U36156 (N_36156,N_33348,N_30222);
and U36157 (N_36157,N_33863,N_31658);
nor U36158 (N_36158,N_33435,N_32329);
nor U36159 (N_36159,N_31681,N_30873);
or U36160 (N_36160,N_30007,N_32729);
nor U36161 (N_36161,N_30904,N_32658);
or U36162 (N_36162,N_31952,N_34582);
and U36163 (N_36163,N_34887,N_33391);
or U36164 (N_36164,N_33609,N_33129);
nand U36165 (N_36165,N_30243,N_30737);
and U36166 (N_36166,N_32420,N_33585);
or U36167 (N_36167,N_31090,N_31406);
nor U36168 (N_36168,N_32137,N_34175);
nand U36169 (N_36169,N_30547,N_31101);
xnor U36170 (N_36170,N_34304,N_30543);
xor U36171 (N_36171,N_30316,N_34318);
and U36172 (N_36172,N_32416,N_32440);
and U36173 (N_36173,N_33109,N_31508);
or U36174 (N_36174,N_30505,N_34825);
or U36175 (N_36175,N_34042,N_34795);
nor U36176 (N_36176,N_31001,N_30648);
or U36177 (N_36177,N_34956,N_33231);
and U36178 (N_36178,N_33630,N_30527);
nor U36179 (N_36179,N_34558,N_32455);
nand U36180 (N_36180,N_32335,N_32150);
nor U36181 (N_36181,N_32850,N_31502);
and U36182 (N_36182,N_34366,N_34625);
and U36183 (N_36183,N_30960,N_34721);
nor U36184 (N_36184,N_33956,N_30327);
nand U36185 (N_36185,N_31690,N_30154);
and U36186 (N_36186,N_31858,N_34235);
nor U36187 (N_36187,N_30071,N_30660);
nor U36188 (N_36188,N_32285,N_31540);
and U36189 (N_36189,N_34645,N_34156);
nand U36190 (N_36190,N_34623,N_33256);
nand U36191 (N_36191,N_34312,N_34258);
nor U36192 (N_36192,N_32857,N_31040);
nor U36193 (N_36193,N_31808,N_30134);
or U36194 (N_36194,N_34247,N_33103);
and U36195 (N_36195,N_33848,N_31525);
xor U36196 (N_36196,N_30151,N_33422);
nor U36197 (N_36197,N_32530,N_34479);
nor U36198 (N_36198,N_34745,N_31121);
and U36199 (N_36199,N_32606,N_33610);
and U36200 (N_36200,N_31943,N_31897);
nand U36201 (N_36201,N_30894,N_30384);
or U36202 (N_36202,N_31821,N_34758);
or U36203 (N_36203,N_32182,N_31185);
and U36204 (N_36204,N_34938,N_33303);
and U36205 (N_36205,N_34784,N_30265);
and U36206 (N_36206,N_33295,N_31035);
nor U36207 (N_36207,N_30425,N_33124);
or U36208 (N_36208,N_32576,N_33218);
nand U36209 (N_36209,N_34729,N_34331);
or U36210 (N_36210,N_33110,N_34391);
nor U36211 (N_36211,N_30493,N_34693);
and U36212 (N_36212,N_30783,N_33922);
and U36213 (N_36213,N_31294,N_33427);
nor U36214 (N_36214,N_32582,N_30754);
nand U36215 (N_36215,N_31740,N_32836);
xor U36216 (N_36216,N_31209,N_33818);
xor U36217 (N_36217,N_30043,N_33557);
and U36218 (N_36218,N_31191,N_31314);
xnor U36219 (N_36219,N_30416,N_31565);
xor U36220 (N_36220,N_30267,N_34869);
nand U36221 (N_36221,N_30681,N_34323);
nor U36222 (N_36222,N_30185,N_32074);
nor U36223 (N_36223,N_33861,N_32705);
and U36224 (N_36224,N_34546,N_33615);
xnor U36225 (N_36225,N_30446,N_33322);
and U36226 (N_36226,N_30015,N_31967);
nand U36227 (N_36227,N_31015,N_31316);
or U36228 (N_36228,N_33563,N_34055);
or U36229 (N_36229,N_33749,N_30981);
xnor U36230 (N_36230,N_30747,N_32798);
xnor U36231 (N_36231,N_33383,N_33345);
nor U36232 (N_36232,N_33645,N_34463);
nand U36233 (N_36233,N_33705,N_32149);
nor U36234 (N_36234,N_33461,N_31198);
and U36235 (N_36235,N_30298,N_30026);
nand U36236 (N_36236,N_34413,N_33834);
nor U36237 (N_36237,N_33823,N_30738);
and U36238 (N_36238,N_31409,N_32302);
nand U36239 (N_36239,N_32724,N_32125);
nor U36240 (N_36240,N_33205,N_33551);
nor U36241 (N_36241,N_32737,N_33072);
xor U36242 (N_36242,N_30865,N_33378);
xor U36243 (N_36243,N_34537,N_31012);
nand U36244 (N_36244,N_30556,N_32504);
nand U36245 (N_36245,N_32031,N_31439);
xnor U36246 (N_36246,N_31851,N_34412);
xnor U36247 (N_36247,N_31007,N_33158);
or U36248 (N_36248,N_32428,N_30343);
and U36249 (N_36249,N_32349,N_31398);
or U36250 (N_36250,N_31632,N_34864);
or U36251 (N_36251,N_34074,N_34740);
nand U36252 (N_36252,N_32486,N_32317);
or U36253 (N_36253,N_31242,N_33429);
nor U36254 (N_36254,N_31591,N_32262);
or U36255 (N_36255,N_34692,N_33025);
or U36256 (N_36256,N_32749,N_30680);
and U36257 (N_36257,N_34796,N_33841);
or U36258 (N_36258,N_34720,N_34404);
nor U36259 (N_36259,N_31218,N_31127);
nor U36260 (N_36260,N_30847,N_32948);
nand U36261 (N_36261,N_30361,N_33729);
xor U36262 (N_36262,N_32214,N_33970);
and U36263 (N_36263,N_32380,N_31873);
xor U36264 (N_36264,N_31389,N_30291);
nor U36265 (N_36265,N_31272,N_33282);
or U36266 (N_36266,N_32326,N_33107);
nand U36267 (N_36267,N_33101,N_34640);
or U36268 (N_36268,N_32614,N_32116);
xnor U36269 (N_36269,N_31197,N_30270);
nor U36270 (N_36270,N_32111,N_33703);
nand U36271 (N_36271,N_33291,N_30919);
xnor U36272 (N_36272,N_31667,N_34013);
and U36273 (N_36273,N_32206,N_33237);
nor U36274 (N_36274,N_34766,N_30427);
or U36275 (N_36275,N_31855,N_33509);
nand U36276 (N_36276,N_31621,N_34586);
and U36277 (N_36277,N_34127,N_31431);
xor U36278 (N_36278,N_31998,N_33060);
nor U36279 (N_36279,N_34669,N_32733);
nor U36280 (N_36280,N_30647,N_31298);
nand U36281 (N_36281,N_30922,N_31997);
and U36282 (N_36282,N_34321,N_33080);
or U36283 (N_36283,N_30262,N_34265);
and U36284 (N_36284,N_33691,N_32651);
and U36285 (N_36285,N_30497,N_30778);
nand U36286 (N_36286,N_33352,N_34579);
and U36287 (N_36287,N_31575,N_31539);
and U36288 (N_36288,N_34793,N_34043);
or U36289 (N_36289,N_30239,N_32103);
nand U36290 (N_36290,N_33506,N_32537);
or U36291 (N_36291,N_34228,N_30473);
xor U36292 (N_36292,N_30732,N_32557);
or U36293 (N_36293,N_32338,N_34657);
nand U36294 (N_36294,N_30088,N_31465);
or U36295 (N_36295,N_31665,N_32408);
xor U36296 (N_36296,N_32788,N_30194);
or U36297 (N_36297,N_30948,N_33962);
and U36298 (N_36298,N_30911,N_32522);
xor U36299 (N_36299,N_30719,N_33290);
xor U36300 (N_36300,N_34259,N_30653);
nand U36301 (N_36301,N_32269,N_31339);
and U36302 (N_36302,N_30168,N_34488);
nor U36303 (N_36303,N_30492,N_30926);
nand U36304 (N_36304,N_33503,N_33989);
xnor U36305 (N_36305,N_33329,N_34914);
or U36306 (N_36306,N_30871,N_30224);
nor U36307 (N_36307,N_32848,N_33846);
xor U36308 (N_36308,N_34168,N_32934);
or U36309 (N_36309,N_34269,N_32711);
and U36310 (N_36310,N_32807,N_34308);
nor U36311 (N_36311,N_33713,N_30211);
nand U36312 (N_36312,N_32583,N_32077);
nand U36313 (N_36313,N_31205,N_34125);
and U36314 (N_36314,N_32875,N_32800);
or U36315 (N_36315,N_32071,N_34792);
or U36316 (N_36316,N_34408,N_31120);
and U36317 (N_36317,N_32974,N_30179);
or U36318 (N_36318,N_31816,N_31146);
or U36319 (N_36319,N_30823,N_30604);
nor U36320 (N_36320,N_31281,N_31081);
xnor U36321 (N_36321,N_30381,N_32880);
nand U36322 (N_36322,N_31442,N_31590);
and U36323 (N_36323,N_30067,N_30791);
nand U36324 (N_36324,N_30714,N_32722);
nand U36325 (N_36325,N_32045,N_33791);
or U36326 (N_36326,N_33565,N_30292);
nand U36327 (N_36327,N_31204,N_31141);
or U36328 (N_36328,N_33140,N_32940);
xnor U36329 (N_36329,N_32468,N_34935);
or U36330 (N_36330,N_30231,N_32593);
or U36331 (N_36331,N_31494,N_34846);
and U36332 (N_36332,N_30930,N_34006);
and U36333 (N_36333,N_30506,N_32563);
xnor U36334 (N_36334,N_34210,N_32573);
nor U36335 (N_36335,N_32541,N_32671);
xnor U36336 (N_36336,N_31657,N_32598);
or U36337 (N_36337,N_32412,N_30599);
nand U36338 (N_36338,N_34899,N_32536);
or U36339 (N_36339,N_30512,N_34388);
nand U36340 (N_36340,N_31775,N_34008);
and U36341 (N_36341,N_34674,N_31689);
xnor U36342 (N_36342,N_31006,N_34124);
xor U36343 (N_36343,N_30893,N_32611);
nor U36344 (N_36344,N_33220,N_32485);
and U36345 (N_36345,N_30805,N_31661);
nand U36346 (N_36346,N_30663,N_33670);
and U36347 (N_36347,N_32492,N_30965);
or U36348 (N_36348,N_33594,N_32717);
nor U36349 (N_36349,N_34890,N_34619);
nand U36350 (N_36350,N_31918,N_31145);
or U36351 (N_36351,N_34478,N_33859);
nor U36352 (N_36352,N_34945,N_34942);
nand U36353 (N_36353,N_33229,N_32951);
and U36354 (N_36354,N_34529,N_31470);
nor U36355 (N_36355,N_31388,N_32391);
and U36356 (N_36356,N_34234,N_33144);
xor U36357 (N_36357,N_34783,N_31326);
and U36358 (N_36358,N_33977,N_33875);
or U36359 (N_36359,N_30499,N_33020);
or U36360 (N_36360,N_34761,N_32892);
and U36361 (N_36361,N_33533,N_32538);
nand U36362 (N_36362,N_30985,N_34474);
xor U36363 (N_36363,N_30999,N_34040);
and U36364 (N_36364,N_34058,N_31152);
or U36365 (N_36365,N_32532,N_31934);
and U36366 (N_36366,N_34603,N_30753);
nand U36367 (N_36367,N_30434,N_30483);
and U36368 (N_36368,N_33965,N_31863);
or U36369 (N_36369,N_33745,N_34117);
xnor U36370 (N_36370,N_34612,N_32158);
and U36371 (N_36371,N_34680,N_33112);
xor U36372 (N_36372,N_30276,N_30392);
xnor U36373 (N_36373,N_31868,N_33413);
xor U36374 (N_36374,N_31721,N_30006);
and U36375 (N_36375,N_34044,N_31969);
nand U36376 (N_36376,N_34615,N_33141);
nand U36377 (N_36377,N_33055,N_30336);
xor U36378 (N_36378,N_30850,N_34229);
xor U36379 (N_36379,N_33568,N_34440);
nor U36380 (N_36380,N_31257,N_32465);
or U36381 (N_36381,N_33531,N_34369);
or U36382 (N_36382,N_30175,N_31423);
nand U36383 (N_36383,N_30888,N_34930);
or U36384 (N_36384,N_32179,N_31801);
and U36385 (N_36385,N_32998,N_34184);
or U36386 (N_36386,N_31142,N_31346);
nand U36387 (N_36387,N_32591,N_33545);
nor U36388 (N_36388,N_33904,N_32884);
nand U36389 (N_36389,N_30219,N_34760);
xnor U36390 (N_36390,N_31947,N_34022);
and U36391 (N_36391,N_33377,N_32476);
and U36392 (N_36392,N_33799,N_31002);
nor U36393 (N_36393,N_31853,N_33741);
nand U36394 (N_36394,N_32808,N_33761);
and U36395 (N_36395,N_34989,N_31950);
and U36396 (N_36396,N_32988,N_30465);
xor U36397 (N_36397,N_31245,N_32141);
nand U36398 (N_36398,N_34459,N_31484);
xor U36399 (N_36399,N_33811,N_34152);
or U36400 (N_36400,N_34327,N_34661);
nand U36401 (N_36401,N_33677,N_32997);
nor U36402 (N_36402,N_31706,N_33415);
or U36403 (N_36403,N_31896,N_33773);
nor U36404 (N_36404,N_33106,N_31293);
and U36405 (N_36405,N_32364,N_30667);
nand U36406 (N_36406,N_33084,N_31649);
xor U36407 (N_36407,N_31818,N_33273);
or U36408 (N_36408,N_30442,N_31451);
xor U36409 (N_36409,N_30315,N_30411);
nand U36410 (N_36410,N_30917,N_33402);
or U36411 (N_36411,N_34372,N_34662);
or U36412 (N_36412,N_31815,N_31617);
nand U36413 (N_36413,N_30699,N_31444);
or U36414 (N_36414,N_31957,N_33937);
nand U36415 (N_36415,N_33153,N_32574);
nor U36416 (N_36416,N_34505,N_30305);
nand U36417 (N_36417,N_34514,N_33940);
xor U36418 (N_36418,N_34302,N_32093);
or U36419 (N_36419,N_34583,N_31310);
nor U36420 (N_36420,N_30638,N_33338);
nor U36421 (N_36421,N_32560,N_34908);
and U36422 (N_36422,N_32634,N_31522);
xor U36423 (N_36423,N_30013,N_30443);
nand U36424 (N_36424,N_30137,N_30378);
or U36425 (N_36425,N_33376,N_30803);
and U36426 (N_36426,N_34670,N_33314);
and U36427 (N_36427,N_32199,N_30010);
nor U36428 (N_36428,N_31327,N_32080);
and U36429 (N_36429,N_32278,N_33795);
and U36430 (N_36430,N_34397,N_30061);
or U36431 (N_36431,N_33755,N_34491);
or U36432 (N_36432,N_31062,N_30187);
or U36433 (N_36433,N_32421,N_30004);
xor U36434 (N_36434,N_32794,N_31807);
and U36435 (N_36435,N_33046,N_33073);
nand U36436 (N_36436,N_34829,N_33717);
nor U36437 (N_36437,N_31254,N_33226);
xnor U36438 (N_36438,N_33824,N_30777);
and U36439 (N_36439,N_32167,N_31830);
or U36440 (N_36440,N_34207,N_30075);
and U36441 (N_36441,N_34671,N_30484);
xor U36442 (N_36442,N_34158,N_32230);
nor U36443 (N_36443,N_32765,N_34494);
nand U36444 (N_36444,N_32626,N_30371);
xnor U36445 (N_36445,N_32856,N_32070);
nand U36446 (N_36446,N_30670,N_32423);
nor U36447 (N_36447,N_30767,N_32007);
nand U36448 (N_36448,N_34845,N_30030);
nand U36449 (N_36449,N_34059,N_30372);
or U36450 (N_36450,N_32697,N_30250);
nor U36451 (N_36451,N_32612,N_34851);
and U36452 (N_36452,N_33876,N_33023);
nor U36453 (N_36453,N_33406,N_33633);
nand U36454 (N_36454,N_30491,N_30974);
and U36455 (N_36455,N_34621,N_31073);
nand U36456 (N_36456,N_34993,N_33381);
nand U36457 (N_36457,N_34644,N_33891);
and U36458 (N_36458,N_31852,N_34429);
xor U36459 (N_36459,N_30356,N_32248);
or U36460 (N_36460,N_31018,N_33496);
nor U36461 (N_36461,N_31495,N_30373);
and U36462 (N_36462,N_34910,N_30617);
xor U36463 (N_36463,N_34484,N_31876);
nor U36464 (N_36464,N_31032,N_31548);
xor U36465 (N_36465,N_32152,N_34742);
xor U36466 (N_36466,N_31233,N_34105);
and U36467 (N_36467,N_31370,N_31263);
or U36468 (N_36468,N_34774,N_33064);
or U36469 (N_36469,N_33852,N_31029);
or U36470 (N_36470,N_34922,N_32929);
or U36471 (N_36471,N_32742,N_32728);
xor U36472 (N_36472,N_30982,N_32853);
xor U36473 (N_36473,N_30813,N_30544);
or U36474 (N_36474,N_32818,N_31300);
nor U36475 (N_36475,N_34664,N_34381);
nand U36476 (N_36476,N_30456,N_33275);
xnor U36477 (N_36477,N_32023,N_34723);
nand U36478 (N_36478,N_30779,N_33605);
nand U36479 (N_36479,N_33895,N_32978);
and U36480 (N_36480,N_32242,N_32160);
nand U36481 (N_36481,N_32414,N_31730);
and U36482 (N_36482,N_30633,N_31031);
nand U36483 (N_36483,N_32363,N_30927);
nand U36484 (N_36484,N_34216,N_31579);
nand U36485 (N_36485,N_33793,N_33454);
and U36486 (N_36486,N_31682,N_34093);
xor U36487 (N_36487,N_32238,N_30297);
xnor U36488 (N_36488,N_34933,N_34961);
nor U36489 (N_36489,N_33309,N_33451);
or U36490 (N_36490,N_30176,N_33688);
and U36491 (N_36491,N_34246,N_33330);
or U36492 (N_36492,N_34310,N_30526);
nand U36493 (N_36493,N_33260,N_32210);
nor U36494 (N_36494,N_34830,N_33757);
nand U36495 (N_36495,N_32188,N_30994);
or U36496 (N_36496,N_31282,N_30542);
and U36497 (N_36497,N_33571,N_34033);
and U36498 (N_36498,N_34194,N_30630);
nand U36499 (N_36499,N_33120,N_33850);
nor U36500 (N_36500,N_33473,N_33013);
nor U36501 (N_36501,N_33994,N_34683);
and U36502 (N_36502,N_33202,N_32968);
or U36503 (N_36503,N_31598,N_32865);
and U36504 (N_36504,N_30269,N_30758);
or U36505 (N_36505,N_30393,N_33974);
and U36506 (N_36506,N_34690,N_34870);
and U36507 (N_36507,N_31904,N_32121);
nor U36508 (N_36508,N_34974,N_34952);
or U36509 (N_36509,N_33527,N_30818);
nand U36510 (N_36510,N_31509,N_30872);
nand U36511 (N_36511,N_34469,N_30279);
and U36512 (N_36512,N_34799,N_30983);
or U36513 (N_36513,N_32944,N_34339);
nor U36514 (N_36514,N_32025,N_30127);
nor U36515 (N_36515,N_33819,N_34777);
and U36516 (N_36516,N_32627,N_32679);
nand U36517 (N_36517,N_33736,N_30107);
or U36518 (N_36518,N_32382,N_30001);
nand U36519 (N_36519,N_34068,N_34875);
xnor U36520 (N_36520,N_32223,N_31724);
nor U36521 (N_36521,N_31835,N_34466);
and U36522 (N_36522,N_32819,N_31817);
nand U36523 (N_36523,N_32407,N_33337);
nand U36524 (N_36524,N_32994,N_30089);
nand U36525 (N_36525,N_32869,N_33726);
xnor U36526 (N_36526,N_30217,N_33221);
and U36527 (N_36527,N_31328,N_33681);
nand U36528 (N_36528,N_34668,N_31971);
and U36529 (N_36529,N_30455,N_31296);
nand U36530 (N_36530,N_33505,N_32241);
nand U36531 (N_36531,N_33266,N_33334);
nand U36532 (N_36532,N_32688,N_30931);
and U36533 (N_36533,N_32822,N_30944);
xor U36534 (N_36534,N_31445,N_33768);
or U36535 (N_36535,N_32763,N_30859);
nand U36536 (N_36536,N_34639,N_31348);
nand U36537 (N_36537,N_34422,N_30666);
and U36538 (N_36538,N_34065,N_32985);
and U36539 (N_36539,N_31672,N_31678);
xor U36540 (N_36540,N_32114,N_31117);
and U36541 (N_36541,N_30407,N_34170);
xnor U36542 (N_36542,N_31587,N_32299);
nand U36543 (N_36543,N_34203,N_32773);
nand U36544 (N_36544,N_34778,N_33706);
nor U36545 (N_36545,N_33354,N_30363);
nand U36546 (N_36546,N_32358,N_31974);
nand U36547 (N_36547,N_34120,N_34380);
xor U36548 (N_36548,N_31714,N_33400);
and U36549 (N_36549,N_30225,N_34924);
nand U36550 (N_36550,N_31028,N_30344);
and U36551 (N_36551,N_32860,N_34296);
nand U36552 (N_36552,N_30557,N_34771);
and U36553 (N_36553,N_33236,N_33283);
nand U36554 (N_36554,N_30065,N_33163);
or U36555 (N_36555,N_32603,N_33810);
nand U36556 (N_36556,N_30423,N_32657);
xnor U36557 (N_36557,N_31616,N_30459);
or U36558 (N_36558,N_33803,N_30528);
or U36559 (N_36559,N_34361,N_33486);
nor U36560 (N_36560,N_31147,N_33344);
nand U36561 (N_36561,N_34589,N_34326);
or U36562 (N_36562,N_32035,N_34805);
and U36563 (N_36563,N_34667,N_34005);
or U36564 (N_36564,N_33285,N_32712);
nand U36565 (N_36565,N_34926,N_32660);
and U36566 (N_36566,N_33169,N_30612);
and U36567 (N_36567,N_30782,N_30197);
nand U36568 (N_36568,N_30032,N_33739);
or U36569 (N_36569,N_32840,N_32234);
nor U36570 (N_36570,N_30842,N_33052);
and U36571 (N_36571,N_32352,N_31011);
nand U36572 (N_36572,N_34472,N_33550);
nor U36573 (N_36573,N_31415,N_32318);
xnor U36574 (N_36574,N_34544,N_33102);
nor U36575 (N_36575,N_33019,N_34944);
or U36576 (N_36576,N_32280,N_33579);
xor U36577 (N_36577,N_33969,N_34442);
nor U36578 (N_36578,N_32674,N_30050);
or U36579 (N_36579,N_33830,N_33346);
nor U36580 (N_36580,N_34434,N_31180);
or U36581 (N_36581,N_34003,N_30729);
and U36582 (N_36582,N_34687,N_31601);
and U36583 (N_36583,N_30764,N_30746);
xor U36584 (N_36584,N_34528,N_33166);
nand U36585 (N_36585,N_32561,N_31580);
nor U36586 (N_36586,N_34814,N_31352);
or U36587 (N_36587,N_32168,N_33067);
nor U36588 (N_36588,N_34416,N_34552);
xnor U36589 (N_36589,N_31975,N_34030);
nor U36590 (N_36590,N_33728,N_34493);
and U36591 (N_36591,N_31777,N_31875);
nor U36592 (N_36592,N_31307,N_33648);
xor U36593 (N_36593,N_31921,N_33821);
xnor U36594 (N_36594,N_31487,N_32607);
and U36595 (N_36595,N_31124,N_33239);
and U36596 (N_36596,N_34673,N_32029);
xnor U36597 (N_36597,N_32072,N_33340);
nand U36598 (N_36598,N_31432,N_30809);
and U36599 (N_36599,N_32567,N_33687);
nand U36600 (N_36600,N_30787,N_32469);
and U36601 (N_36601,N_32038,N_34086);
xnor U36602 (N_36602,N_34808,N_32436);
nand U36603 (N_36603,N_32686,N_34091);
nor U36604 (N_36604,N_34585,N_31898);
nand U36605 (N_36605,N_33032,N_31075);
nand U36606 (N_36606,N_30554,N_33361);
and U36607 (N_36607,N_33082,N_30885);
xnor U36608 (N_36608,N_33925,N_30645);
xor U36609 (N_36609,N_34432,N_32571);
or U36610 (N_36610,N_33081,N_33479);
and U36611 (N_36611,N_32553,N_34651);
and U36612 (N_36612,N_32255,N_33371);
and U36613 (N_36613,N_33298,N_30525);
and U36614 (N_36614,N_32895,N_32140);
nand U36615 (N_36615,N_34686,N_34981);
nand U36616 (N_36616,N_31744,N_32886);
nand U36617 (N_36617,N_30877,N_31363);
nand U36618 (N_36618,N_34525,N_33047);
or U36619 (N_36619,N_34920,N_30607);
or U36620 (N_36620,N_30739,N_31287);
nand U36621 (N_36621,N_34739,N_30848);
nor U36622 (N_36622,N_32600,N_32931);
and U36623 (N_36623,N_31306,N_34465);
xor U36624 (N_36624,N_32581,N_32037);
nand U36625 (N_36625,N_34502,N_30382);
and U36626 (N_36626,N_32621,N_30408);
nand U36627 (N_36627,N_33299,N_34031);
or U36628 (N_36628,N_31557,N_34752);
and U36629 (N_36629,N_34066,N_32562);
nor U36630 (N_36630,N_30039,N_34897);
nand U36631 (N_36631,N_31134,N_31113);
nor U36632 (N_36632,N_34702,N_34385);
nor U36633 (N_36633,N_31620,N_32958);
nand U36634 (N_36634,N_32867,N_33203);
xor U36635 (N_36635,N_30730,N_34614);
and U36636 (N_36636,N_33912,N_34932);
nor U36637 (N_36637,N_33360,N_34034);
nand U36638 (N_36638,N_34631,N_31797);
and U36639 (N_36639,N_34348,N_32019);
nor U36640 (N_36640,N_33748,N_31895);
or U36641 (N_36641,N_32666,N_33599);
nor U36642 (N_36642,N_30329,N_31261);
nor U36643 (N_36643,N_34239,N_32231);
and U36644 (N_36644,N_32524,N_31356);
and U36645 (N_36645,N_32559,N_30159);
nand U36646 (N_36646,N_32648,N_34678);
and U36647 (N_36647,N_31408,N_30422);
nor U36648 (N_36648,N_34755,N_30707);
nor U36649 (N_36649,N_32801,N_31938);
or U36650 (N_36650,N_31222,N_30869);
xor U36651 (N_36651,N_32746,N_31360);
xnor U36652 (N_36652,N_30584,N_34374);
nand U36653 (N_36653,N_30997,N_30735);
nand U36654 (N_36654,N_31794,N_34951);
or U36655 (N_36655,N_34565,N_34263);
and U36656 (N_36656,N_30358,N_30689);
xnor U36657 (N_36657,N_32693,N_33998);
or U36658 (N_36658,N_31345,N_30074);
nor U36659 (N_36659,N_34898,N_32756);
or U36660 (N_36660,N_34226,N_31397);
nand U36661 (N_36661,N_30899,N_33085);
nand U36662 (N_36662,N_33390,N_33460);
xor U36663 (N_36663,N_31367,N_34208);
and U36664 (N_36664,N_34605,N_31933);
or U36665 (N_36665,N_30524,N_33651);
xnor U36666 (N_36666,N_33488,N_34282);
and U36667 (N_36667,N_32804,N_33133);
and U36668 (N_36668,N_30426,N_34367);
and U36669 (N_36669,N_32004,N_30441);
or U36670 (N_36670,N_32580,N_30589);
xor U36671 (N_36671,N_34837,N_34744);
nor U36672 (N_36672,N_34351,N_32699);
nor U36673 (N_36673,N_32858,N_31864);
nand U36674 (N_36674,N_31189,N_32237);
nand U36675 (N_36675,N_32172,N_31258);
nand U36676 (N_36676,N_34097,N_34237);
and U36677 (N_36677,N_31153,N_30144);
xnor U36678 (N_36678,N_30275,N_33063);
and U36679 (N_36679,N_30935,N_33903);
nor U36680 (N_36680,N_32952,N_31770);
nor U36681 (N_36681,N_31008,N_30244);
nand U36682 (N_36682,N_33440,N_31320);
xnor U36683 (N_36683,N_34676,N_32493);
or U36684 (N_36684,N_34123,N_34911);
or U36685 (N_36685,N_32692,N_31096);
or U36686 (N_36686,N_30420,N_30118);
or U36687 (N_36687,N_30898,N_31100);
xor U36688 (N_36688,N_33007,N_33259);
and U36689 (N_36689,N_33553,N_33854);
xnor U36690 (N_36690,N_33712,N_34295);
nand U36691 (N_36691,N_34666,N_33179);
and U36692 (N_36692,N_32174,N_33154);
nand U36693 (N_36693,N_31208,N_32235);
xor U36694 (N_36694,N_33029,N_31985);
nand U36695 (N_36695,N_31182,N_30047);
nor U36696 (N_36696,N_30916,N_34881);
nor U36697 (N_36697,N_32078,N_31489);
nor U36698 (N_36698,N_30975,N_31505);
nand U36699 (N_36699,N_31400,N_33398);
nor U36700 (N_36700,N_31069,N_31103);
nand U36701 (N_36701,N_31125,N_34477);
and U36702 (N_36702,N_34378,N_32466);
or U36703 (N_36703,N_32048,N_34789);
xor U36704 (N_36704,N_30600,N_31917);
xor U36705 (N_36705,N_30114,N_30992);
or U36706 (N_36706,N_32899,N_31107);
nor U36707 (N_36707,N_30951,N_31190);
nor U36708 (N_36708,N_31593,N_32266);
nor U36709 (N_36709,N_32642,N_34001);
nor U36710 (N_36710,N_32494,N_30155);
xor U36711 (N_36711,N_30252,N_31958);
nand U36712 (N_36712,N_32233,N_31491);
xor U36713 (N_36713,N_32938,N_32437);
nor U36714 (N_36714,N_32361,N_33227);
nor U36715 (N_36715,N_34580,N_33134);
and U36716 (N_36716,N_31772,N_32619);
nor U36717 (N_36717,N_33450,N_32258);
or U36718 (N_36718,N_31531,N_31072);
nand U36719 (N_36719,N_32322,N_32321);
nand U36720 (N_36720,N_30632,N_33178);
and U36721 (N_36721,N_30195,N_34350);
nor U36722 (N_36722,N_30106,N_34877);
nor U36723 (N_36723,N_30910,N_34636);
and U36724 (N_36724,N_33128,N_33933);
or U36725 (N_36725,N_30347,N_33149);
xnor U36726 (N_36726,N_32897,N_34298);
nand U36727 (N_36727,N_30691,N_30720);
nand U36728 (N_36728,N_30272,N_32620);
nor U36729 (N_36729,N_32893,N_33470);
xnor U36730 (N_36730,N_34015,N_32715);
or U36731 (N_36731,N_30509,N_33079);
xnor U36732 (N_36732,N_34349,N_31122);
and U36733 (N_36733,N_33500,N_34038);
xor U36734 (N_36734,N_34305,N_30449);
nand U36735 (N_36735,N_30915,N_33207);
and U36736 (N_36736,N_31312,N_34129);
xor U36737 (N_36737,N_30545,N_32374);
nor U36738 (N_36738,N_31890,N_30713);
nand U36739 (N_36739,N_32218,N_30072);
or U36740 (N_36740,N_32584,N_34386);
xnor U36741 (N_36741,N_30642,N_33719);
nand U36742 (N_36742,N_34923,N_33873);
nor U36743 (N_36743,N_30242,N_31437);
nor U36744 (N_36744,N_32334,N_33704);
nor U36745 (N_36745,N_30518,N_31631);
nand U36746 (N_36746,N_34151,N_30108);
nand U36747 (N_36747,N_30082,N_31275);
nor U36748 (N_36748,N_30136,N_33611);
and U36749 (N_36749,N_32528,N_33332);
and U36750 (N_36750,N_34214,N_33407);
nand U36751 (N_36751,N_34876,N_30903);
and U36752 (N_36752,N_32664,N_30353);
nand U36753 (N_36753,N_34630,N_33065);
nand U36754 (N_36754,N_32992,N_34713);
nand U36755 (N_36755,N_33566,N_32514);
nor U36756 (N_36756,N_31663,N_32919);
xnor U36757 (N_36757,N_31498,N_32639);
nand U36758 (N_36758,N_30312,N_30751);
or U36759 (N_36759,N_30104,N_30306);
nand U36760 (N_36760,N_31051,N_34931);
xnor U36761 (N_36761,N_32112,N_34420);
xnor U36762 (N_36762,N_32588,N_30113);
xnor U36763 (N_36763,N_32148,N_30444);
and U36764 (N_36764,N_31283,N_33465);
or U36765 (N_36765,N_33170,N_31483);
nand U36766 (N_36766,N_34197,N_30801);
and U36767 (N_36767,N_30963,N_31187);
xor U36768 (N_36768,N_33701,N_32987);
nand U36769 (N_36769,N_31776,N_34785);
and U36770 (N_36770,N_32508,N_30521);
xor U36771 (N_36771,N_33946,N_31805);
xnor U36772 (N_36772,N_33198,N_31037);
nand U36773 (N_36773,N_31212,N_33423);
or U36774 (N_36774,N_33206,N_30376);
or U36775 (N_36775,N_31049,N_30765);
nand U36776 (N_36776,N_33247,N_32405);
nand U36777 (N_36777,N_34950,N_32675);
xnor U36778 (N_36778,N_30889,N_32097);
xnor U36779 (N_36779,N_30832,N_33045);
or U36780 (N_36780,N_33162,N_34285);
or U36781 (N_36781,N_33448,N_31463);
nor U36782 (N_36782,N_32925,N_34046);
nor U36783 (N_36783,N_31965,N_34593);
nor U36784 (N_36784,N_33444,N_33495);
nor U36785 (N_36785,N_32676,N_34994);
and U36786 (N_36786,N_32185,N_30679);
and U36787 (N_36787,N_33180,N_32171);
and U36788 (N_36788,N_31836,N_34757);
or U36789 (N_36789,N_31698,N_33008);
xor U36790 (N_36790,N_34048,N_30961);
or U36791 (N_36791,N_33668,N_31108);
nor U36792 (N_36792,N_32333,N_34373);
nor U36793 (N_36793,N_30996,N_34275);
or U36794 (N_36794,N_32395,N_30161);
nor U36795 (N_36795,N_32296,N_32142);
nand U36796 (N_36796,N_32661,N_33498);
and U36797 (N_36797,N_32339,N_33433);
or U36798 (N_36798,N_32198,N_32823);
or U36799 (N_36799,N_30116,N_32385);
xnor U36800 (N_36800,N_31516,N_30644);
xor U36801 (N_36801,N_34756,N_31099);
xor U36802 (N_36802,N_32084,N_33302);
nor U36803 (N_36803,N_30307,N_33507);
nand U36804 (N_36804,N_31244,N_34106);
nor U36805 (N_36805,N_31995,N_34821);
nor U36806 (N_36806,N_30792,N_31181);
xnor U36807 (N_36807,N_33964,N_33947);
nor U36808 (N_36808,N_33176,N_32922);
nor U36809 (N_36809,N_30700,N_33044);
or U36810 (N_36810,N_34962,N_33832);
and U36811 (N_36811,N_34550,N_34337);
or U36812 (N_36812,N_31589,N_32187);
or U36813 (N_36813,N_33347,N_33735);
nor U36814 (N_36814,N_32517,N_31679);
or U36815 (N_36815,N_33062,N_32714);
xnor U36816 (N_36816,N_30240,N_34539);
nor U36817 (N_36817,N_31043,N_33968);
nand U36818 (N_36818,N_30775,N_30362);
xor U36819 (N_36819,N_30620,N_30421);
xnor U36820 (N_36820,N_32480,N_34622);
or U36821 (N_36821,N_32786,N_33185);
or U36822 (N_36822,N_30200,N_31292);
or U36823 (N_36823,N_31217,N_32327);
nand U36824 (N_36824,N_30862,N_32028);
or U36825 (N_36825,N_33426,N_33012);
or U36826 (N_36826,N_31550,N_32707);
xor U36827 (N_36827,N_32270,N_34365);
nor U36828 (N_36828,N_31582,N_34957);
and U36829 (N_36829,N_30141,N_34573);
nor U36830 (N_36830,N_32067,N_34336);
nand U36831 (N_36831,N_30566,N_34798);
xnor U36832 (N_36832,N_32161,N_33526);
or U36833 (N_36833,N_32854,N_31826);
xnor U36834 (N_36834,N_30824,N_32216);
nand U36835 (N_36835,N_32774,N_32549);
xor U36836 (N_36836,N_31110,N_31419);
and U36837 (N_36837,N_34301,N_32649);
nor U36838 (N_36838,N_34069,N_34588);
nand U36839 (N_36839,N_30051,N_33463);
and U36840 (N_36840,N_30046,N_32298);
nand U36841 (N_36841,N_30069,N_32989);
nor U36842 (N_36842,N_31675,N_33204);
and U36843 (N_36843,N_34507,N_33328);
nand U36844 (N_36844,N_32024,N_30150);
nand U36845 (N_36845,N_34425,N_33403);
and U36846 (N_36846,N_30133,N_34196);
and U36847 (N_36847,N_31856,N_34972);
nand U36848 (N_36848,N_30640,N_30029);
and U36849 (N_36849,N_30800,N_32265);
and U36850 (N_36850,N_32059,N_30755);
nor U36851 (N_36851,N_34554,N_31973);
xor U36852 (N_36852,N_33659,N_34900);
xor U36853 (N_36853,N_33716,N_33930);
nor U36854 (N_36854,N_33242,N_34147);
nand U36855 (N_36855,N_33942,N_32341);
nor U36856 (N_36856,N_33578,N_31748);
nand U36857 (N_36857,N_31854,N_30772);
nand U36858 (N_36858,N_31407,N_31227);
nor U36859 (N_36859,N_32002,N_32672);
xor U36860 (N_36860,N_32201,N_34949);
nand U36861 (N_36861,N_33297,N_31893);
and U36862 (N_36862,N_31716,N_34150);
xnor U36863 (N_36863,N_33661,N_34293);
xnor U36864 (N_36864,N_34232,N_34400);
nand U36865 (N_36865,N_31503,N_31132);
nor U36866 (N_36866,N_33333,N_32151);
and U36867 (N_36867,N_31823,N_30979);
xnor U36868 (N_36868,N_30958,N_32887);
or U36869 (N_36869,N_31441,N_31428);
nor U36870 (N_36870,N_34883,N_34183);
nor U36871 (N_36871,N_31910,N_34287);
nor U36872 (N_36872,N_30918,N_30703);
or U36873 (N_36873,N_33909,N_31737);
xnor U36874 (N_36874,N_32026,N_32131);
or U36875 (N_36875,N_34880,N_33856);
xnor U36876 (N_36876,N_31336,N_31086);
nand U36877 (N_36877,N_30383,N_34857);
and U36878 (N_36878,N_31860,N_33223);
and U36879 (N_36879,N_33866,N_32821);
or U36880 (N_36880,N_33612,N_33049);
and U36881 (N_36881,N_33388,N_32273);
or U36882 (N_36882,N_33631,N_30991);
or U36883 (N_36883,N_30310,N_30845);
and U36884 (N_36884,N_31981,N_30998);
and U36885 (N_36885,N_30855,N_32102);
and U36886 (N_36886,N_31906,N_31302);
or U36887 (N_36887,N_31929,N_34730);
and U36888 (N_36888,N_31078,N_31155);
xor U36889 (N_36889,N_32410,N_32211);
nor U36890 (N_36890,N_34362,N_32100);
nand U36891 (N_36891,N_30439,N_33077);
nand U36892 (N_36892,N_33094,N_33017);
nand U36893 (N_36893,N_32499,N_30627);
and U36894 (N_36894,N_32289,N_32495);
and U36895 (N_36895,N_31480,N_34487);
or U36896 (N_36896,N_31055,N_33814);
or U36897 (N_36897,N_34462,N_30435);
and U36898 (N_36898,N_30819,N_32689);
nor U36899 (N_36899,N_32531,N_32645);
and U36900 (N_36900,N_34217,N_33357);
nor U36901 (N_36901,N_33253,N_30056);
nand U36902 (N_36902,N_33569,N_33521);
and U36903 (N_36903,N_32311,N_30084);
nor U36904 (N_36904,N_32725,N_33041);
nand U36905 (N_36905,N_30212,N_32228);
nor U36906 (N_36906,N_34359,N_34853);
nor U36907 (N_36907,N_33792,N_32791);
nand U36908 (N_36908,N_32694,N_33801);
nand U36909 (N_36909,N_30938,N_33288);
xor U36910 (N_36910,N_31422,N_34145);
xor U36911 (N_36911,N_30406,N_30215);
or U36912 (N_36912,N_34343,N_31683);
and U36913 (N_36913,N_33629,N_33137);
nand U36914 (N_36914,N_33996,N_34450);
nand U36915 (N_36915,N_31552,N_33193);
and U36916 (N_36916,N_33642,N_30993);
nor U36917 (N_36917,N_33159,N_30606);
nand U36918 (N_36918,N_32700,N_30815);
nand U36919 (N_36919,N_34198,N_30024);
nand U36920 (N_36920,N_31769,N_31342);
and U36921 (N_36921,N_33016,N_30476);
xnor U36922 (N_36922,N_31627,N_32392);
nand U36923 (N_36923,N_34224,N_33167);
or U36924 (N_36924,N_33118,N_31250);
xor U36925 (N_36925,N_33399,N_31329);
nor U36926 (N_36926,N_34553,N_31615);
nand U36927 (N_36927,N_34698,N_33175);
nor U36928 (N_36928,N_30081,N_30213);
or U36929 (N_36929,N_31962,N_31532);
nand U36930 (N_36930,N_31158,N_32239);
xnor U36931 (N_36931,N_30851,N_33271);
nor U36932 (N_36932,N_32398,N_31916);
and U36933 (N_36933,N_31705,N_30248);
nor U36934 (N_36934,N_30947,N_30064);
and U36935 (N_36935,N_33126,N_30757);
nand U36936 (N_36936,N_31978,N_31461);
nor U36937 (N_36937,N_34283,N_33790);
and U36938 (N_36938,N_33324,N_32589);
nor U36939 (N_36939,N_34490,N_32613);
and U36940 (N_36940,N_33590,N_33208);
nand U36941 (N_36941,N_34188,N_30829);
xnor U36942 (N_36942,N_34786,N_32320);
and U36943 (N_36943,N_34741,N_32790);
nand U36944 (N_36944,N_34245,N_34426);
xnor U36945 (N_36945,N_34272,N_31709);
nor U36946 (N_36946,N_32212,N_30076);
and U36947 (N_36947,N_33838,N_31886);
nor U36948 (N_36948,N_30011,N_30706);
nor U36949 (N_36949,N_33879,N_31478);
nand U36950 (N_36950,N_31758,N_33339);
and U36951 (N_36951,N_34460,N_34483);
nor U36952 (N_36952,N_32803,N_30906);
or U36953 (N_36953,N_30057,N_31156);
xor U36954 (N_36954,N_30472,N_30626);
nor U36955 (N_36955,N_31481,N_31686);
nor U36956 (N_36956,N_31337,N_31882);
xnor U36957 (N_36957,N_33501,N_33030);
xnor U36958 (N_36958,N_33350,N_30023);
xnor U36959 (N_36959,N_32984,N_33418);
and U36960 (N_36960,N_31213,N_33943);
nor U36961 (N_36961,N_31533,N_30657);
xnor U36962 (N_36962,N_34567,N_34079);
nand U36963 (N_36963,N_32635,N_30500);
xnor U36964 (N_36964,N_34254,N_32570);
xor U36965 (N_36965,N_30396,N_30428);
nand U36966 (N_36966,N_34445,N_31742);
nor U36967 (N_36967,N_32044,N_32847);
and U36968 (N_36968,N_30255,N_34868);
or U36969 (N_36969,N_31266,N_33528);
xnor U36970 (N_36970,N_31528,N_32971);
nor U36971 (N_36971,N_32319,N_30369);
nor U36972 (N_36972,N_32527,N_31361);
xor U36973 (N_36973,N_32637,N_33040);
xnor U36974 (N_36974,N_33484,N_31695);
nand U36975 (N_36975,N_33543,N_33911);
nor U36976 (N_36976,N_32075,N_31382);
xnor U36977 (N_36977,N_32507,N_34201);
and U36978 (N_36978,N_34842,N_32076);
xnor U36979 (N_36979,N_33296,N_31949);
or U36980 (N_36980,N_31030,N_31224);
nand U36981 (N_36981,N_31458,N_33096);
or U36982 (N_36982,N_32286,N_31786);
and U36983 (N_36983,N_33515,N_34172);
nor U36984 (N_36984,N_33274,N_32796);
xnor U36985 (N_36985,N_31129,N_30639);
and U36986 (N_36986,N_32999,N_34076);
or U36987 (N_36987,N_34624,N_34457);
xor U36988 (N_36988,N_34334,N_30042);
nand U36989 (N_36989,N_31469,N_33359);
xnor U36990 (N_36990,N_30397,N_31685);
and U36991 (N_36991,N_31699,N_33069);
or U36992 (N_36992,N_30283,N_31023);
or U36993 (N_36993,N_33797,N_31752);
and U36994 (N_36994,N_31274,N_33225);
nand U36995 (N_36995,N_31178,N_30939);
nor U36996 (N_36996,N_32473,N_33375);
and U36997 (N_36997,N_33455,N_33733);
or U36998 (N_36998,N_32244,N_33767);
or U36999 (N_36999,N_31754,N_30533);
nor U37000 (N_37000,N_34248,N_31492);
nand U37001 (N_37001,N_32936,N_33954);
or U37002 (N_37002,N_31696,N_30535);
xnor U37003 (N_37003,N_34264,N_31646);
and U37004 (N_37004,N_30748,N_33542);
nand U37005 (N_37005,N_34917,N_30328);
or U37006 (N_37006,N_30768,N_33105);
and U37007 (N_37007,N_33690,N_31555);
nor U37008 (N_37008,N_34094,N_30976);
xor U37009 (N_37009,N_34663,N_33257);
xor U37010 (N_37010,N_32979,N_33950);
nor U37011 (N_37011,N_33439,N_30115);
nor U37012 (N_37012,N_34443,N_30652);
or U37013 (N_37013,N_32488,N_31796);
nand U37014 (N_37014,N_32739,N_30395);
or U37015 (N_37015,N_34083,N_34360);
xnor U37016 (N_37016,N_31232,N_32849);
and U37017 (N_37017,N_30103,N_30690);
and U37018 (N_37018,N_31759,N_30980);
nand U37019 (N_37019,N_32511,N_34193);
nor U37020 (N_37020,N_34177,N_32177);
xnor U37021 (N_37021,N_31673,N_31247);
or U37022 (N_37022,N_30568,N_32701);
nor U37023 (N_37023,N_30309,N_34154);
xnor U37024 (N_37024,N_32295,N_30247);
nor U37025 (N_37025,N_32505,N_31829);
nor U37026 (N_37026,N_32065,N_30237);
and U37027 (N_37027,N_30866,N_33510);
or U37028 (N_37028,N_32926,N_31438);
xor U37029 (N_37029,N_30833,N_30798);
nor U37030 (N_37030,N_34340,N_31728);
or U37031 (N_37031,N_31172,N_32898);
nor U37032 (N_37032,N_33626,N_33636);
nand U37033 (N_37033,N_31633,N_33089);
nor U37034 (N_37034,N_33453,N_34602);
and U37035 (N_37035,N_33921,N_30946);
xnor U37036 (N_37036,N_34765,N_34428);
xor U37037 (N_37037,N_30709,N_31420);
and U37038 (N_37038,N_33785,N_34306);
and U37039 (N_37039,N_32138,N_30579);
or U37040 (N_37040,N_32418,N_31359);
and U37041 (N_37041,N_30966,N_34597);
nand U37042 (N_37042,N_32180,N_30879);
nor U37043 (N_37043,N_33216,N_34341);
or U37044 (N_37044,N_32246,N_31602);
or U37045 (N_37045,N_34052,N_33387);
or U37046 (N_37046,N_32448,N_32399);
and U37047 (N_37047,N_31764,N_34826);
nand U37048 (N_37048,N_33042,N_30734);
nor U37049 (N_37049,N_32219,N_34294);
or U37050 (N_37050,N_34130,N_31623);
nand U37051 (N_37051,N_31810,N_33270);
nor U37052 (N_37052,N_32133,N_30132);
and U37053 (N_37053,N_30028,N_33753);
and U37054 (N_37054,N_32753,N_31221);
xnor U37055 (N_37055,N_31828,N_31380);
xnor U37056 (N_37056,N_34347,N_31662);
nor U37057 (N_37057,N_34379,N_33662);
xnor U37058 (N_37058,N_33392,N_31931);
nand U37059 (N_37059,N_33963,N_31883);
xnor U37060 (N_37060,N_34734,N_32704);
or U37061 (N_37061,N_33813,N_32542);
and U37062 (N_37062,N_34149,N_31578);
nand U37063 (N_37063,N_34970,N_34634);
nor U37064 (N_37064,N_31603,N_32417);
or U37065 (N_37065,N_32040,N_31993);
or U37066 (N_37066,N_33177,N_33696);
or U37067 (N_37067,N_33076,N_30857);
and U37068 (N_37068,N_33758,N_32876);
xor U37069 (N_37069,N_31597,N_32888);
and U37070 (N_37070,N_34410,N_32795);
nand U37071 (N_37071,N_34519,N_31583);
xnor U37072 (N_37072,N_31554,N_34866);
and U37073 (N_37073,N_32592,N_32939);
nand U37074 (N_37074,N_32923,N_34405);
nor U37075 (N_37075,N_31092,N_30515);
nand U37076 (N_37076,N_32402,N_34081);
or U37077 (N_37077,N_30415,N_32950);
and U37078 (N_37078,N_34677,N_34243);
xor U37079 (N_37079,N_32878,N_30100);
and U37080 (N_37080,N_32901,N_34179);
xor U37081 (N_37081,N_30308,N_34753);
nor U37082 (N_37082,N_30560,N_30330);
nand U37083 (N_37083,N_32236,N_32458);
or U37084 (N_37084,N_30229,N_33654);
or U37085 (N_37085,N_32376,N_32245);
nor U37086 (N_37086,N_34506,N_33356);
and U37087 (N_37087,N_34534,N_32816);
xnor U37088 (N_37088,N_33327,N_32272);
nor U37089 (N_37089,N_33581,N_33769);
or U37090 (N_37090,N_30846,N_30550);
xor U37091 (N_37091,N_34921,N_34889);
and U37092 (N_37092,N_30286,N_32438);
nand U37093 (N_37093,N_32107,N_32479);
nand U37094 (N_37094,N_34943,N_31079);
xnor U37095 (N_37095,N_33368,N_30623);
nor U37096 (N_37096,N_33776,N_33916);
nand U37097 (N_37097,N_30199,N_30987);
nand U37098 (N_37098,N_31925,N_34233);
or U37099 (N_37099,N_32064,N_33547);
nand U37100 (N_37100,N_30111,N_34522);
nand U37101 (N_37101,N_31192,N_31745);
nand U37102 (N_37102,N_33244,N_32431);
nor U37103 (N_37103,N_33173,N_32343);
xor U37104 (N_37104,N_34987,N_32424);
xor U37105 (N_37105,N_30685,N_33737);
nor U37106 (N_37106,N_31584,N_30978);
or U37107 (N_37107,N_34476,N_34895);
nand U37108 (N_37108,N_32404,N_32467);
and U37109 (N_37109,N_30637,N_34335);
or U37110 (N_37110,N_31126,N_34114);
and U37111 (N_37111,N_31362,N_34872);
nand U37112 (N_37112,N_30016,N_32957);
nand U37113 (N_37113,N_33880,N_31381);
nor U37114 (N_37114,N_33300,N_31570);
nand U37115 (N_37115,N_33574,N_31504);
nor U37116 (N_37116,N_32061,N_31160);
nand U37117 (N_37117,N_31162,N_33417);
xnor U37118 (N_37118,N_34261,N_34819);
nor U37119 (N_37119,N_32057,N_32904);
nor U37120 (N_37120,N_31640,N_31067);
or U37121 (N_37121,N_33517,N_30238);
nand U37122 (N_37122,N_34427,N_32916);
and U37123 (N_37123,N_32873,N_31596);
and U37124 (N_37124,N_31526,N_31600);
xor U37125 (N_37125,N_33815,N_33497);
or U37126 (N_37126,N_32991,N_33188);
xor U37127 (N_37127,N_34344,N_33211);
nor U37128 (N_37128,N_31252,N_32115);
nand U37129 (N_37129,N_33416,N_34126);
and U37130 (N_37130,N_33168,N_34936);
nand U37131 (N_37131,N_33132,N_31572);
nand U37132 (N_37132,N_33586,N_33336);
xnor U37133 (N_37133,N_32290,N_31749);
and U37134 (N_37134,N_30646,N_32066);
or U37135 (N_37135,N_30077,N_32769);
or U37136 (N_37136,N_30902,N_31577);
and U37137 (N_37137,N_32257,N_31647);
or U37138 (N_37138,N_30235,N_32797);
or U37139 (N_37139,N_34444,N_33152);
and U37140 (N_37140,N_33997,N_32411);
nor U37141 (N_37141,N_30957,N_32490);
and U37142 (N_37142,N_34291,N_31165);
xor U37143 (N_37143,N_32575,N_30696);
xor U37144 (N_37144,N_30208,N_33607);
nand U37145 (N_37145,N_33394,N_32457);
nand U37146 (N_37146,N_34456,N_30578);
nand U37147 (N_37147,N_31956,N_33932);
nor U37148 (N_37148,N_33160,N_34726);
or U37149 (N_37149,N_30401,N_32190);
nor U37150 (N_37150,N_32362,N_33548);
or U37151 (N_37151,N_30055,N_33535);
and U37152 (N_37152,N_31016,N_31521);
nor U37153 (N_37153,N_32396,N_31269);
xor U37154 (N_37154,N_32768,N_31456);
or U37155 (N_37155,N_30870,N_33502);
nor U37156 (N_37156,N_34489,N_34804);
and U37157 (N_37157,N_30424,N_32069);
or U37158 (N_37158,N_30496,N_34833);
xnor U37159 (N_37159,N_33366,N_33635);
nand U37160 (N_37160,N_31932,N_30405);
nand U37161 (N_37161,N_31335,N_32946);
nor U37162 (N_37162,N_31251,N_34653);
xnor U37163 (N_37163,N_31859,N_32802);
nor U37164 (N_37164,N_34103,N_33472);
nor U37165 (N_37165,N_34212,N_32949);
nor U37166 (N_37166,N_33150,N_33593);
xnor U37167 (N_37167,N_30530,N_34419);
or U37168 (N_37168,N_34162,N_30095);
xnor U37169 (N_37169,N_30021,N_31071);
nor U37170 (N_37170,N_34737,N_33576);
nand U37171 (N_37171,N_32970,N_32986);
or U37172 (N_37172,N_30209,N_32471);
nand U37173 (N_37173,N_31911,N_30760);
nand U37174 (N_37174,N_33066,N_33199);
xor U37175 (N_37175,N_31070,N_33171);
or U37176 (N_37176,N_31677,N_31708);
or U37177 (N_37177,N_33692,N_34570);
nand U37178 (N_37178,N_31416,N_31277);
xor U37179 (N_37179,N_30880,N_33541);
nand U37180 (N_37180,N_32271,N_31889);
nand U37181 (N_37181,N_30692,N_30431);
xnor U37182 (N_37182,N_33634,N_34119);
nand U37183 (N_37183,N_30206,N_32087);
or U37184 (N_37184,N_33181,N_32910);
and U37185 (N_37185,N_31374,N_30952);
or U37186 (N_37186,N_31847,N_30450);
or U37187 (N_37187,N_30814,N_30895);
xnor U37188 (N_37188,N_33731,N_31684);
or U37189 (N_37189,N_34473,N_31395);
nor U37190 (N_37190,N_33192,N_32088);
and U37191 (N_37191,N_30676,N_33491);
nor U37192 (N_37192,N_34991,N_33899);
and U37193 (N_37193,N_31558,N_32202);
and U37194 (N_37194,N_33759,N_33822);
nand U37195 (N_37195,N_30736,N_34496);
xor U37196 (N_37196,N_33524,N_31066);
and U37197 (N_37197,N_34847,N_30494);
nand U37198 (N_37198,N_30836,N_30489);
xnor U37199 (N_37199,N_32058,N_34101);
nor U37200 (N_37200,N_31084,N_32120);
nor U37201 (N_37201,N_31206,N_33920);
nor U37202 (N_37202,N_33816,N_32928);
and U37203 (N_37203,N_33554,N_33281);
nor U37204 (N_37204,N_30101,N_33917);
xnor U37205 (N_37205,N_30955,N_33700);
xnor U37206 (N_37206,N_33224,N_31614);
nand U37207 (N_37207,N_31524,N_34371);
nand U37208 (N_37208,N_34414,N_30458);
and U37209 (N_37209,N_30538,N_34963);
nand U37210 (N_37210,N_33955,N_34718);
xor U37211 (N_37211,N_31991,N_30907);
and U37212 (N_37212,N_31609,N_34569);
nand U37213 (N_37213,N_34595,N_34353);
and U37214 (N_37214,N_30368,N_33849);
nor U37215 (N_37215,N_34036,N_32336);
or U37216 (N_37216,N_31243,N_34701);
or U37217 (N_37217,N_31253,N_34650);
or U37218 (N_37218,N_33197,N_34260);
and U37219 (N_37219,N_31130,N_34581);
nor U37220 (N_37220,N_30605,N_30293);
xor U37221 (N_37221,N_34904,N_30864);
nor U37222 (N_37222,N_31036,N_31891);
or U37223 (N_37223,N_32681,N_32747);
nand U37224 (N_37224,N_30232,N_32147);
and U37225 (N_37225,N_34027,N_31396);
or U37226 (N_37226,N_32831,N_31666);
xnor U37227 (N_37227,N_32277,N_34080);
or U37228 (N_37228,N_32578,N_34859);
nand U37229 (N_37229,N_31654,N_34010);
nor U37230 (N_37230,N_30672,N_34274);
and U37231 (N_37231,N_33546,N_31691);
or U37232 (N_37232,N_34557,N_32534);
nor U37233 (N_37233,N_34266,N_32130);
nand U37234 (N_37234,N_32885,N_33992);
and U37235 (N_37235,N_34722,N_34087);
nand U37236 (N_37236,N_34873,N_33845);
xnor U37237 (N_37237,N_33475,N_31607);
nand U37238 (N_37238,N_34628,N_31713);
xor U37239 (N_37239,N_31476,N_30597);
nand U37240 (N_37240,N_34512,N_31256);
nand U37241 (N_37241,N_33976,N_33380);
nand U37242 (N_37242,N_33305,N_32365);
xor U37243 (N_37243,N_32041,N_34165);
nor U37244 (N_37244,N_31867,N_33802);
xor U37245 (N_37245,N_33564,N_32706);
nand U37246 (N_37246,N_34205,N_31383);
and U37247 (N_37247,N_32827,N_30149);
xnor U37248 (N_37248,N_32276,N_34417);
or U37249 (N_37249,N_31262,N_32872);
xnor U37250 (N_37250,N_30374,N_34000);
and U37251 (N_37251,N_33494,N_31280);
xnor U37252 (N_37252,N_34200,N_31241);
nor U37253 (N_37253,N_33959,N_32348);
xnor U37254 (N_37254,N_30854,N_32894);
or U37255 (N_37255,N_31173,N_30080);
nor U37256 (N_37256,N_31866,N_32006);
nand U37257 (N_37257,N_34684,N_34738);
nor U37258 (N_37258,N_33004,N_30349);
and U37259 (N_37259,N_31869,N_33372);
nor U37260 (N_37260,N_30146,N_30192);
xnor U37261 (N_37261,N_30471,N_34501);
or U37262 (N_37262,N_31785,N_31270);
or U37263 (N_37263,N_31351,N_34070);
xor U37264 (N_37264,N_31219,N_31248);
nor U37265 (N_37265,N_33858,N_32444);
or U37266 (N_37266,N_31800,N_33313);
nor U37267 (N_37267,N_30682,N_30092);
or U37268 (N_37268,N_31899,N_31089);
xnor U37269 (N_37269,N_34314,N_33906);
nor U37270 (N_37270,N_31414,N_30553);
and U37271 (N_37271,N_30079,N_30586);
nor U37272 (N_37272,N_32817,N_31743);
nor U37273 (N_37273,N_34415,N_33614);
and U37274 (N_37274,N_34939,N_33914);
nor U37275 (N_37275,N_30953,N_31556);
and U37276 (N_37276,N_30357,N_31518);
nor U37277 (N_37277,N_31846,N_31376);
nor U37278 (N_37278,N_33306,N_32046);
and U37279 (N_37279,N_32636,N_32516);
nand U37280 (N_37280,N_34997,N_33697);
or U37281 (N_37281,N_30788,N_30070);
xor U37282 (N_37282,N_34355,N_34346);
or U37283 (N_37283,N_31806,N_32996);
nand U37284 (N_37284,N_34893,N_33172);
nor U37285 (N_37285,N_30673,N_31700);
nand U37286 (N_37286,N_31017,N_32920);
and U37287 (N_37287,N_30959,N_32870);
and U37288 (N_37288,N_32977,N_32995);
nor U37289 (N_37289,N_32586,N_31506);
xor U37290 (N_37290,N_32325,N_32845);
xnor U37291 (N_37291,N_34787,N_31964);
nand U37292 (N_37292,N_31105,N_31080);
or U37293 (N_37293,N_33006,N_31942);
or U37294 (N_37294,N_31013,N_34791);
nor U37295 (N_37295,N_30802,N_33151);
and U37296 (N_37296,N_32053,N_33709);
and U37297 (N_37297,N_34453,N_32647);
xnor U37298 (N_37298,N_32990,N_31948);
or U37299 (N_37299,N_33872,N_33613);
nand U37300 (N_37300,N_33369,N_33397);
xnor U37301 (N_37301,N_34874,N_32117);
nor U37302 (N_37302,N_34708,N_30201);
nand U37303 (N_37303,N_33623,N_32119);
nand U37304 (N_37304,N_34107,N_33039);
xnor U37305 (N_37305,N_30841,N_33115);
nor U37306 (N_37306,N_34647,N_30338);
nand U37307 (N_37307,N_31613,N_31098);
nand U37308 (N_37308,N_34023,N_33428);
nor U37309 (N_37309,N_34050,N_33929);
nor U37310 (N_37310,N_30583,N_30625);
xnor U37311 (N_37311,N_34746,N_31660);
or U37312 (N_37312,N_31923,N_30326);
nand U37313 (N_37313,N_33523,N_32225);
or U37314 (N_37314,N_33003,N_31822);
xor U37315 (N_37315,N_31813,N_34095);
xnor U37316 (N_37316,N_33130,N_32366);
xnor U37317 (N_37317,N_30852,N_31061);
xnor U37318 (N_37318,N_34892,N_32851);
nand U37319 (N_37319,N_33561,N_31450);
xnor U37320 (N_37320,N_33676,N_34262);
and U37321 (N_37321,N_33087,N_32003);
and U37322 (N_37322,N_32354,N_30156);
nor U37323 (N_37323,N_34626,N_31729);
xnor U37324 (N_37324,N_32000,N_31637);
and U37325 (N_37325,N_32945,N_31634);
nand U37326 (N_37326,N_32838,N_31926);
nand U37327 (N_37327,N_30749,N_34133);
xor U37328 (N_37328,N_34788,N_31323);
and U37329 (N_37329,N_31239,N_34606);
nand U37330 (N_37330,N_30592,N_33254);
nand U37331 (N_37331,N_34186,N_31214);
or U37332 (N_37332,N_34311,N_30562);
and U37333 (N_37333,N_32013,N_31042);
xor U37334 (N_37334,N_30467,N_32793);
nor U37335 (N_37335,N_31334,N_30726);
and U37336 (N_37336,N_34007,N_30731);
nand U37337 (N_37337,N_34725,N_33070);
nand U37338 (N_37338,N_33617,N_32209);
and U37339 (N_37339,N_33711,N_30522);
nand U37340 (N_37340,N_31318,N_31364);
xor U37341 (N_37341,N_31123,N_32288);
nand U37342 (N_37342,N_31026,N_30126);
nand U37343 (N_37343,N_34236,N_34223);
xor U37344 (N_37344,N_32965,N_32735);
nor U37345 (N_37345,N_31378,N_34148);
nand U37346 (N_37346,N_31814,N_34053);
nand U37347 (N_37347,N_34775,N_31802);
nor U37348 (N_37348,N_31872,N_31611);
xnor U37349 (N_37349,N_31674,N_33784);
and U37350 (N_37350,N_33147,N_30616);
nand U37351 (N_37351,N_31319,N_31782);
nand U37352 (N_37352,N_30086,N_33255);
nor U37353 (N_37353,N_34660,N_33853);
nand U37354 (N_37354,N_34084,N_30901);
nand U37355 (N_37355,N_30433,N_34574);
xor U37356 (N_37356,N_33022,N_33341);
xor U37357 (N_37357,N_32771,N_32752);
or U37358 (N_37358,N_34854,N_32813);
nor U37359 (N_37359,N_30514,N_33982);
or U37360 (N_37360,N_33616,N_33820);
xnor U37361 (N_37361,N_34222,N_32164);
or U37362 (N_37362,N_32618,N_33114);
nor U37363 (N_37363,N_30041,N_32523);
or U37364 (N_37364,N_30721,N_33628);
or U37365 (N_37365,N_30228,N_31773);
and U37366 (N_37366,N_31455,N_33490);
nor U37367 (N_37367,N_30482,N_33829);
nor U37368 (N_37368,N_34681,N_33504);
xor U37369 (N_37369,N_34253,N_33363);
or U37370 (N_37370,N_31482,N_30565);
and U37371 (N_37371,N_33002,N_31468);
and U37372 (N_37372,N_33127,N_34167);
and U37373 (N_37373,N_34618,N_34026);
xnor U37374 (N_37374,N_31541,N_33897);
and U37375 (N_37375,N_33606,N_31511);
nor U37376 (N_37376,N_34862,N_32178);
and U37377 (N_37377,N_32347,N_31025);
and U37378 (N_37378,N_30674,N_32941);
nor U37379 (N_37379,N_30878,N_32001);
xor U37380 (N_37380,N_34329,N_34215);
xor U37381 (N_37381,N_32662,N_31144);
nor U37382 (N_37382,N_34596,N_30321);
and U37383 (N_37383,N_34707,N_33775);
and U37384 (N_37384,N_32777,N_34646);
or U37385 (N_37385,N_33228,N_30322);
and U37386 (N_37386,N_33385,N_32902);
nand U37387 (N_37387,N_32085,N_34382);
xnor U37388 (N_37388,N_32372,N_31903);
and U37389 (N_37389,N_30875,N_31137);
or U37390 (N_37390,N_32513,N_30624);
or U37391 (N_37391,N_31083,N_31939);
nor U37392 (N_37392,N_31862,N_30234);
or U37393 (N_37393,N_30977,N_30186);
and U37394 (N_37394,N_33860,N_30173);
or U37395 (N_37395,N_34599,N_32224);
and U37396 (N_37396,N_34665,N_33438);
and U37397 (N_37397,N_30771,N_33732);
and U37398 (N_37398,N_32982,N_31766);
nand U37399 (N_37399,N_34905,N_32824);
nand U37400 (N_37400,N_31385,N_31940);
and U37401 (N_37401,N_31405,N_34021);
nor U37402 (N_37402,N_34815,N_30261);
or U37403 (N_37403,N_32967,N_31211);
nand U37404 (N_37404,N_30348,N_31424);
or U37405 (N_37405,N_33437,N_30145);
nand U37406 (N_37406,N_31284,N_32782);
nand U37407 (N_37407,N_32815,N_32477);
or U37408 (N_37408,N_33870,N_33918);
or U37409 (N_37409,N_32727,N_33786);
nor U37410 (N_37410,N_31586,N_32032);
or U37411 (N_37411,N_30346,N_30287);
and U37412 (N_37412,N_31426,N_30587);
nand U37413 (N_37413,N_34689,N_33928);
or U37414 (N_37414,N_31060,N_31791);
nor U37415 (N_37415,N_31220,N_30636);
nor U37416 (N_37416,N_33656,N_33446);
and U37417 (N_37417,N_32091,N_32082);
or U37418 (N_37418,N_32259,N_31427);
nor U37419 (N_37419,N_32461,N_31630);
nand U37420 (N_37420,N_31139,N_30311);
or U37421 (N_37421,N_30128,N_30487);
and U37422 (N_37422,N_34843,N_31022);
xnor U37423 (N_37423,N_30909,N_30914);
and U37424 (N_37424,N_33195,N_32175);
nor U37425 (N_37425,N_33304,N_34658);
and U37426 (N_37426,N_33138,N_34794);
nand U37427 (N_37427,N_30655,N_30468);
nor U37428 (N_37428,N_33230,N_34984);
xnor U37429 (N_37429,N_33869,N_30385);
or U37430 (N_37430,N_30839,N_30054);
nand U37431 (N_37431,N_34421,N_31566);
nand U37432 (N_37432,N_32730,N_32868);
and U37433 (N_37433,N_31065,N_32760);
nor U37434 (N_37434,N_32721,N_32852);
or U37435 (N_37435,N_30504,N_34011);
xnor U37436 (N_37436,N_31757,N_32118);
and U37437 (N_37437,N_34966,N_31203);
and U37438 (N_37438,N_30257,N_32337);
and U37439 (N_37439,N_34655,N_32036);
and U37440 (N_37440,N_34953,N_32483);
xnor U37441 (N_37441,N_30890,N_33519);
and U37442 (N_37442,N_31774,N_30296);
nor U37443 (N_37443,N_31148,N_30761);
xnor U37444 (N_37444,N_30402,N_32623);
nand U37445 (N_37445,N_32136,N_31384);
or U37446 (N_37446,N_33900,N_33843);
xnor U37447 (N_37447,N_34035,N_34967);
xor U37448 (N_37448,N_33624,N_34844);
nand U37449 (N_37449,N_30964,N_33219);
nor U37450 (N_37450,N_32812,N_31452);
xor U37451 (N_37451,N_32622,N_31135);
xnor U37452 (N_37452,N_34174,N_31200);
nand U37453 (N_37453,N_30375,N_31977);
nor U37454 (N_37454,N_34250,N_30536);
or U37455 (N_37455,N_31571,N_33393);
or U37456 (N_37456,N_34609,N_32631);
xor U37457 (N_37457,N_30138,N_34064);
or U37458 (N_37458,N_34497,N_34438);
and U37459 (N_37459,N_33183,N_31410);
nand U37460 (N_37460,N_31154,N_31542);
or U37461 (N_37461,N_30303,N_31781);
nor U37462 (N_37462,N_34024,N_33806);
or U37463 (N_37463,N_33092,N_34182);
and U37464 (N_37464,N_32487,N_33808);
and U37465 (N_37465,N_30469,N_32879);
or U37466 (N_37466,N_31267,N_34850);
nor U37467 (N_37467,N_30558,N_31747);
nor U37468 (N_37468,N_30923,N_32829);
nand U37469 (N_37469,N_31368,N_30744);
xnor U37470 (N_37470,N_34925,N_32183);
nor U37471 (N_37471,N_30658,N_34954);
nor U37472 (N_37472,N_33520,N_30183);
nand U37473 (N_37473,N_31003,N_31322);
xnor U37474 (N_37474,N_30825,N_34017);
and U37475 (N_37475,N_32227,N_30464);
nand U37476 (N_37476,N_34025,N_32099);
and U37477 (N_37477,N_32429,N_30523);
nor U37478 (N_37478,N_32446,N_31207);
and U37479 (N_37479,N_31264,N_32653);
and U37480 (N_37480,N_32572,N_31581);
nor U37481 (N_37481,N_30198,N_30157);
or U37482 (N_37482,N_34244,N_31798);
nand U37483 (N_37483,N_34806,N_31231);
or U37484 (N_37484,N_31460,N_32127);
nand U37485 (N_37485,N_33232,N_34517);
nor U37486 (N_37486,N_33730,N_32275);
or U37487 (N_37487,N_34878,N_34041);
nor U37488 (N_37488,N_32154,N_34979);
xnor U37489 (N_37489,N_33781,N_32104);
nor U37490 (N_37490,N_30986,N_31324);
nor U37491 (N_37491,N_33766,N_31014);
xor U37492 (N_37492,N_34092,N_31618);
nor U37493 (N_37493,N_34735,N_31625);
xnor U37494 (N_37494,N_33139,N_32139);
nand U37495 (N_37495,N_31102,N_34075);
and U37496 (N_37496,N_30743,N_33641);
or U37497 (N_37497,N_34763,N_30277);
nand U37498 (N_37498,N_33165,N_34324);
xor U37499 (N_37499,N_31945,N_33721);
nand U37500 (N_37500,N_30366,N_31698);
and U37501 (N_37501,N_32238,N_30460);
nand U37502 (N_37502,N_34641,N_31597);
nand U37503 (N_37503,N_30402,N_33498);
or U37504 (N_37504,N_30379,N_31317);
xnor U37505 (N_37505,N_30506,N_31385);
or U37506 (N_37506,N_31433,N_32870);
nand U37507 (N_37507,N_34580,N_30002);
nor U37508 (N_37508,N_30146,N_32750);
and U37509 (N_37509,N_34636,N_33381);
or U37510 (N_37510,N_33767,N_34988);
nor U37511 (N_37511,N_34110,N_31336);
xor U37512 (N_37512,N_31711,N_30307);
xnor U37513 (N_37513,N_32296,N_34337);
xor U37514 (N_37514,N_31346,N_33072);
and U37515 (N_37515,N_31706,N_32943);
nor U37516 (N_37516,N_33951,N_34387);
or U37517 (N_37517,N_34161,N_33411);
xnor U37518 (N_37518,N_31507,N_34407);
nor U37519 (N_37519,N_31690,N_32660);
nor U37520 (N_37520,N_30886,N_30466);
xnor U37521 (N_37521,N_30099,N_30833);
xor U37522 (N_37522,N_32871,N_31480);
nor U37523 (N_37523,N_34700,N_31280);
and U37524 (N_37524,N_30546,N_33548);
xnor U37525 (N_37525,N_31024,N_31992);
xnor U37526 (N_37526,N_31394,N_33391);
or U37527 (N_37527,N_31812,N_30902);
nand U37528 (N_37528,N_33370,N_34656);
and U37529 (N_37529,N_33354,N_31243);
nor U37530 (N_37530,N_33530,N_33088);
nand U37531 (N_37531,N_32744,N_30109);
xnor U37532 (N_37532,N_32340,N_34713);
nor U37533 (N_37533,N_30758,N_34771);
xor U37534 (N_37534,N_31143,N_34969);
nor U37535 (N_37535,N_30942,N_31220);
xnor U37536 (N_37536,N_34461,N_32229);
and U37537 (N_37537,N_33496,N_32620);
nor U37538 (N_37538,N_32657,N_32246);
nand U37539 (N_37539,N_30365,N_34896);
and U37540 (N_37540,N_30098,N_34233);
nor U37541 (N_37541,N_34419,N_33493);
nor U37542 (N_37542,N_33564,N_33623);
nor U37543 (N_37543,N_34139,N_30179);
or U37544 (N_37544,N_32280,N_33828);
and U37545 (N_37545,N_34125,N_33734);
nand U37546 (N_37546,N_33863,N_30357);
xnor U37547 (N_37547,N_32545,N_32685);
nor U37548 (N_37548,N_33609,N_30459);
xor U37549 (N_37549,N_33376,N_31546);
nand U37550 (N_37550,N_30252,N_30264);
nor U37551 (N_37551,N_34851,N_31418);
xor U37552 (N_37552,N_34149,N_33538);
nor U37553 (N_37553,N_34676,N_34904);
and U37554 (N_37554,N_30784,N_32826);
xnor U37555 (N_37555,N_32539,N_32664);
nand U37556 (N_37556,N_32232,N_32723);
xnor U37557 (N_37557,N_33034,N_31980);
or U37558 (N_37558,N_31900,N_32916);
or U37559 (N_37559,N_30605,N_31480);
xor U37560 (N_37560,N_30871,N_31661);
or U37561 (N_37561,N_32133,N_31713);
xor U37562 (N_37562,N_33476,N_31159);
xor U37563 (N_37563,N_34390,N_32680);
nand U37564 (N_37564,N_30392,N_33799);
xor U37565 (N_37565,N_31065,N_32327);
nor U37566 (N_37566,N_31569,N_33842);
nor U37567 (N_37567,N_33524,N_31499);
or U37568 (N_37568,N_30853,N_31035);
nand U37569 (N_37569,N_31073,N_31185);
nand U37570 (N_37570,N_34213,N_34152);
nor U37571 (N_37571,N_33096,N_31298);
xnor U37572 (N_37572,N_33519,N_30855);
nor U37573 (N_37573,N_34150,N_33836);
nand U37574 (N_37574,N_30196,N_30414);
nor U37575 (N_37575,N_30784,N_31098);
or U37576 (N_37576,N_33466,N_30964);
nand U37577 (N_37577,N_33016,N_32951);
and U37578 (N_37578,N_32072,N_33878);
nand U37579 (N_37579,N_34915,N_33307);
nand U37580 (N_37580,N_33567,N_31531);
xor U37581 (N_37581,N_33010,N_33014);
and U37582 (N_37582,N_31942,N_32315);
nor U37583 (N_37583,N_32801,N_34293);
and U37584 (N_37584,N_33589,N_34883);
and U37585 (N_37585,N_32892,N_31775);
nor U37586 (N_37586,N_31768,N_32570);
and U37587 (N_37587,N_30574,N_32909);
or U37588 (N_37588,N_33566,N_30220);
xor U37589 (N_37589,N_30619,N_33736);
nor U37590 (N_37590,N_34348,N_30738);
xor U37591 (N_37591,N_30521,N_31655);
and U37592 (N_37592,N_33570,N_33572);
nand U37593 (N_37593,N_34187,N_33132);
and U37594 (N_37594,N_31121,N_31498);
xor U37595 (N_37595,N_32408,N_33867);
xor U37596 (N_37596,N_34448,N_33065);
xnor U37597 (N_37597,N_30209,N_33270);
xor U37598 (N_37598,N_33654,N_34760);
nor U37599 (N_37599,N_34704,N_30343);
nand U37600 (N_37600,N_34605,N_30504);
and U37601 (N_37601,N_31413,N_32441);
or U37602 (N_37602,N_34364,N_34209);
nand U37603 (N_37603,N_33481,N_30049);
or U37604 (N_37604,N_30503,N_31775);
or U37605 (N_37605,N_31327,N_33247);
nand U37606 (N_37606,N_34942,N_34146);
xnor U37607 (N_37607,N_32017,N_30932);
nand U37608 (N_37608,N_31861,N_31175);
nand U37609 (N_37609,N_33477,N_34798);
and U37610 (N_37610,N_33821,N_33028);
nand U37611 (N_37611,N_34408,N_32738);
or U37612 (N_37612,N_33302,N_30431);
nor U37613 (N_37613,N_34586,N_32504);
xnor U37614 (N_37614,N_30157,N_31385);
and U37615 (N_37615,N_30412,N_33752);
nand U37616 (N_37616,N_30151,N_34743);
nor U37617 (N_37617,N_31494,N_30714);
nor U37618 (N_37618,N_34808,N_30569);
and U37619 (N_37619,N_30741,N_31882);
and U37620 (N_37620,N_32369,N_33917);
or U37621 (N_37621,N_34962,N_31060);
xor U37622 (N_37622,N_33151,N_33939);
xnor U37623 (N_37623,N_31248,N_31824);
xnor U37624 (N_37624,N_32042,N_34161);
nand U37625 (N_37625,N_33278,N_32227);
nand U37626 (N_37626,N_30514,N_33551);
and U37627 (N_37627,N_32826,N_30421);
nor U37628 (N_37628,N_33406,N_30207);
nand U37629 (N_37629,N_30852,N_32076);
or U37630 (N_37630,N_30093,N_33451);
and U37631 (N_37631,N_31542,N_34342);
and U37632 (N_37632,N_34245,N_33868);
nand U37633 (N_37633,N_30250,N_33459);
nor U37634 (N_37634,N_33236,N_34402);
nand U37635 (N_37635,N_31922,N_34061);
nand U37636 (N_37636,N_32745,N_32661);
xnor U37637 (N_37637,N_31583,N_33125);
xnor U37638 (N_37638,N_30350,N_31578);
nand U37639 (N_37639,N_33217,N_30072);
nor U37640 (N_37640,N_34504,N_30631);
and U37641 (N_37641,N_31638,N_34729);
nor U37642 (N_37642,N_31791,N_32064);
xnor U37643 (N_37643,N_34665,N_32112);
nor U37644 (N_37644,N_31712,N_30864);
and U37645 (N_37645,N_30964,N_32397);
xor U37646 (N_37646,N_34699,N_30617);
or U37647 (N_37647,N_34895,N_34181);
and U37648 (N_37648,N_31647,N_32518);
xnor U37649 (N_37649,N_33062,N_34687);
or U37650 (N_37650,N_33587,N_33462);
xnor U37651 (N_37651,N_32108,N_30657);
or U37652 (N_37652,N_34272,N_33081);
and U37653 (N_37653,N_31906,N_34666);
xor U37654 (N_37654,N_34190,N_33474);
nand U37655 (N_37655,N_34107,N_30365);
or U37656 (N_37656,N_30813,N_33647);
nand U37657 (N_37657,N_33074,N_34458);
and U37658 (N_37658,N_32633,N_32488);
or U37659 (N_37659,N_33542,N_31994);
xor U37660 (N_37660,N_30381,N_33804);
nand U37661 (N_37661,N_33996,N_34890);
nor U37662 (N_37662,N_32293,N_34807);
or U37663 (N_37663,N_31324,N_33503);
and U37664 (N_37664,N_33940,N_34538);
or U37665 (N_37665,N_31750,N_34884);
xnor U37666 (N_37666,N_32054,N_33121);
or U37667 (N_37667,N_34996,N_31373);
and U37668 (N_37668,N_32874,N_34075);
or U37669 (N_37669,N_34713,N_32220);
xnor U37670 (N_37670,N_31485,N_34105);
xnor U37671 (N_37671,N_31051,N_31273);
and U37672 (N_37672,N_31514,N_31787);
nor U37673 (N_37673,N_30814,N_32620);
and U37674 (N_37674,N_31758,N_30211);
or U37675 (N_37675,N_30826,N_30430);
or U37676 (N_37676,N_32529,N_30193);
nor U37677 (N_37677,N_34131,N_34553);
or U37678 (N_37678,N_30770,N_30426);
xor U37679 (N_37679,N_30487,N_33127);
and U37680 (N_37680,N_31830,N_33950);
and U37681 (N_37681,N_34879,N_33904);
nor U37682 (N_37682,N_31775,N_31617);
nor U37683 (N_37683,N_32530,N_34869);
and U37684 (N_37684,N_32335,N_30059);
nor U37685 (N_37685,N_31672,N_31130);
or U37686 (N_37686,N_33588,N_32285);
nor U37687 (N_37687,N_32886,N_32650);
or U37688 (N_37688,N_32721,N_30237);
or U37689 (N_37689,N_31242,N_30390);
nor U37690 (N_37690,N_30264,N_34945);
xnor U37691 (N_37691,N_32835,N_30586);
or U37692 (N_37692,N_32517,N_33292);
or U37693 (N_37693,N_31728,N_30372);
xor U37694 (N_37694,N_31560,N_31634);
nand U37695 (N_37695,N_34467,N_33208);
or U37696 (N_37696,N_32849,N_31891);
nor U37697 (N_37697,N_33880,N_31506);
nand U37698 (N_37698,N_31821,N_32656);
or U37699 (N_37699,N_33208,N_34845);
and U37700 (N_37700,N_30179,N_31945);
or U37701 (N_37701,N_30587,N_30207);
or U37702 (N_37702,N_33865,N_30135);
xor U37703 (N_37703,N_34992,N_32636);
xor U37704 (N_37704,N_32220,N_31890);
nand U37705 (N_37705,N_31961,N_31199);
nand U37706 (N_37706,N_31292,N_33244);
xnor U37707 (N_37707,N_33906,N_31239);
and U37708 (N_37708,N_31526,N_30018);
xor U37709 (N_37709,N_31739,N_32800);
and U37710 (N_37710,N_32489,N_31961);
xor U37711 (N_37711,N_31507,N_30156);
nor U37712 (N_37712,N_33089,N_33989);
or U37713 (N_37713,N_32835,N_32505);
nor U37714 (N_37714,N_33759,N_33698);
nand U37715 (N_37715,N_32816,N_30630);
nor U37716 (N_37716,N_34997,N_30548);
or U37717 (N_37717,N_31241,N_30402);
and U37718 (N_37718,N_33647,N_33809);
xor U37719 (N_37719,N_30312,N_32305);
nand U37720 (N_37720,N_34083,N_34782);
and U37721 (N_37721,N_32608,N_31974);
nand U37722 (N_37722,N_30712,N_32277);
or U37723 (N_37723,N_34033,N_30996);
nand U37724 (N_37724,N_34922,N_30946);
or U37725 (N_37725,N_34830,N_32001);
nor U37726 (N_37726,N_31643,N_33903);
nor U37727 (N_37727,N_33317,N_30216);
xor U37728 (N_37728,N_32849,N_33970);
nor U37729 (N_37729,N_32311,N_31140);
and U37730 (N_37730,N_31881,N_34880);
xnor U37731 (N_37731,N_33101,N_32489);
nor U37732 (N_37732,N_30809,N_31821);
or U37733 (N_37733,N_30920,N_31884);
or U37734 (N_37734,N_31851,N_32055);
nand U37735 (N_37735,N_31080,N_31522);
nor U37736 (N_37736,N_32494,N_30178);
nor U37737 (N_37737,N_32087,N_30102);
or U37738 (N_37738,N_33664,N_34514);
or U37739 (N_37739,N_32762,N_32892);
and U37740 (N_37740,N_33399,N_31140);
nor U37741 (N_37741,N_33643,N_32460);
nor U37742 (N_37742,N_33683,N_32827);
or U37743 (N_37743,N_34721,N_32049);
and U37744 (N_37744,N_34858,N_33151);
nor U37745 (N_37745,N_33486,N_33278);
nand U37746 (N_37746,N_30412,N_31958);
xor U37747 (N_37747,N_32016,N_30237);
and U37748 (N_37748,N_31748,N_34881);
or U37749 (N_37749,N_30191,N_33496);
nand U37750 (N_37750,N_34194,N_31306);
nand U37751 (N_37751,N_31285,N_30977);
nor U37752 (N_37752,N_31784,N_31658);
nor U37753 (N_37753,N_32437,N_33496);
nor U37754 (N_37754,N_33825,N_32614);
nor U37755 (N_37755,N_30692,N_33157);
nor U37756 (N_37756,N_30444,N_30869);
and U37757 (N_37757,N_34872,N_32402);
and U37758 (N_37758,N_32020,N_33991);
and U37759 (N_37759,N_32207,N_30619);
xnor U37760 (N_37760,N_31513,N_30143);
nand U37761 (N_37761,N_33467,N_34075);
or U37762 (N_37762,N_30300,N_33612);
or U37763 (N_37763,N_34550,N_33308);
nor U37764 (N_37764,N_33903,N_30439);
nor U37765 (N_37765,N_31166,N_31716);
nor U37766 (N_37766,N_32413,N_32478);
xnor U37767 (N_37767,N_30574,N_34763);
nor U37768 (N_37768,N_30919,N_31734);
xor U37769 (N_37769,N_33685,N_34572);
nor U37770 (N_37770,N_31748,N_34345);
nor U37771 (N_37771,N_32682,N_30097);
nand U37772 (N_37772,N_30098,N_34050);
nor U37773 (N_37773,N_30905,N_33809);
nand U37774 (N_37774,N_31445,N_30694);
nand U37775 (N_37775,N_34953,N_30882);
xor U37776 (N_37776,N_34215,N_34703);
nor U37777 (N_37777,N_30680,N_33979);
nand U37778 (N_37778,N_33914,N_30655);
and U37779 (N_37779,N_31541,N_34812);
nand U37780 (N_37780,N_31783,N_33637);
xor U37781 (N_37781,N_31690,N_31583);
and U37782 (N_37782,N_33543,N_34770);
xnor U37783 (N_37783,N_30595,N_33413);
nor U37784 (N_37784,N_33388,N_33576);
nor U37785 (N_37785,N_34477,N_32901);
xor U37786 (N_37786,N_34262,N_33896);
nand U37787 (N_37787,N_30272,N_34231);
nor U37788 (N_37788,N_32401,N_30912);
nand U37789 (N_37789,N_32452,N_32838);
and U37790 (N_37790,N_31513,N_33610);
nor U37791 (N_37791,N_30697,N_33339);
xor U37792 (N_37792,N_30150,N_33738);
or U37793 (N_37793,N_33882,N_33269);
nand U37794 (N_37794,N_33439,N_32554);
xnor U37795 (N_37795,N_32640,N_33746);
and U37796 (N_37796,N_32177,N_32026);
nor U37797 (N_37797,N_31678,N_32511);
xnor U37798 (N_37798,N_33644,N_34044);
xnor U37799 (N_37799,N_34373,N_33130);
and U37800 (N_37800,N_31542,N_31069);
nor U37801 (N_37801,N_33745,N_30757);
and U37802 (N_37802,N_31786,N_33796);
or U37803 (N_37803,N_31176,N_33693);
or U37804 (N_37804,N_32659,N_30303);
nor U37805 (N_37805,N_32488,N_32123);
or U37806 (N_37806,N_31991,N_34795);
xnor U37807 (N_37807,N_31490,N_33729);
nand U37808 (N_37808,N_30021,N_32212);
and U37809 (N_37809,N_31956,N_31715);
nor U37810 (N_37810,N_34390,N_32075);
nor U37811 (N_37811,N_34974,N_32938);
and U37812 (N_37812,N_34455,N_32633);
or U37813 (N_37813,N_31441,N_34266);
or U37814 (N_37814,N_32467,N_31312);
nand U37815 (N_37815,N_34816,N_34612);
nand U37816 (N_37816,N_34130,N_34103);
nand U37817 (N_37817,N_34894,N_31488);
or U37818 (N_37818,N_30202,N_31920);
or U37819 (N_37819,N_30582,N_31100);
nor U37820 (N_37820,N_33556,N_32778);
and U37821 (N_37821,N_32066,N_31797);
xor U37822 (N_37822,N_34683,N_30228);
and U37823 (N_37823,N_32529,N_33883);
xnor U37824 (N_37824,N_30556,N_34186);
and U37825 (N_37825,N_31278,N_30787);
xor U37826 (N_37826,N_34749,N_31841);
and U37827 (N_37827,N_32179,N_34600);
nor U37828 (N_37828,N_32650,N_33485);
and U37829 (N_37829,N_31594,N_32499);
or U37830 (N_37830,N_34455,N_31545);
xor U37831 (N_37831,N_32033,N_34686);
and U37832 (N_37832,N_30443,N_30290);
xor U37833 (N_37833,N_32818,N_31800);
nand U37834 (N_37834,N_30244,N_31221);
nor U37835 (N_37835,N_32305,N_30912);
and U37836 (N_37836,N_30034,N_31556);
or U37837 (N_37837,N_30882,N_32698);
and U37838 (N_37838,N_30251,N_32422);
xor U37839 (N_37839,N_30537,N_30055);
nand U37840 (N_37840,N_33962,N_34234);
and U37841 (N_37841,N_30030,N_30180);
and U37842 (N_37842,N_32823,N_32985);
and U37843 (N_37843,N_32214,N_33126);
nor U37844 (N_37844,N_31804,N_33719);
nor U37845 (N_37845,N_30105,N_31859);
nor U37846 (N_37846,N_34028,N_33550);
and U37847 (N_37847,N_34818,N_30672);
nor U37848 (N_37848,N_33090,N_30246);
xor U37849 (N_37849,N_31115,N_32254);
and U37850 (N_37850,N_33860,N_32736);
and U37851 (N_37851,N_34916,N_33750);
nand U37852 (N_37852,N_33252,N_33642);
nor U37853 (N_37853,N_30052,N_30702);
and U37854 (N_37854,N_32544,N_31421);
nor U37855 (N_37855,N_34429,N_33808);
nor U37856 (N_37856,N_33711,N_31848);
xor U37857 (N_37857,N_34384,N_31018);
or U37858 (N_37858,N_33689,N_31142);
nand U37859 (N_37859,N_31692,N_33574);
or U37860 (N_37860,N_33766,N_34324);
or U37861 (N_37861,N_33797,N_33169);
and U37862 (N_37862,N_34378,N_34611);
and U37863 (N_37863,N_33061,N_33984);
nand U37864 (N_37864,N_33256,N_32305);
and U37865 (N_37865,N_34619,N_32477);
or U37866 (N_37866,N_33186,N_32526);
nand U37867 (N_37867,N_33636,N_30658);
and U37868 (N_37868,N_33047,N_32281);
xor U37869 (N_37869,N_34389,N_30661);
or U37870 (N_37870,N_30217,N_30463);
and U37871 (N_37871,N_33532,N_32000);
xnor U37872 (N_37872,N_30817,N_30598);
nand U37873 (N_37873,N_34040,N_30415);
or U37874 (N_37874,N_30768,N_31855);
or U37875 (N_37875,N_33075,N_30485);
and U37876 (N_37876,N_33197,N_30233);
or U37877 (N_37877,N_31787,N_30890);
nor U37878 (N_37878,N_32171,N_31548);
and U37879 (N_37879,N_33317,N_33538);
nand U37880 (N_37880,N_33226,N_34262);
and U37881 (N_37881,N_33007,N_32195);
xnor U37882 (N_37882,N_31516,N_31401);
nand U37883 (N_37883,N_33180,N_30992);
and U37884 (N_37884,N_33105,N_30454);
nand U37885 (N_37885,N_33665,N_34863);
or U37886 (N_37886,N_34970,N_32523);
xnor U37887 (N_37887,N_33158,N_32555);
or U37888 (N_37888,N_34638,N_34318);
nor U37889 (N_37889,N_32924,N_33669);
and U37890 (N_37890,N_30564,N_31326);
and U37891 (N_37891,N_34175,N_32320);
nor U37892 (N_37892,N_33697,N_33543);
and U37893 (N_37893,N_31426,N_30521);
and U37894 (N_37894,N_33293,N_32718);
and U37895 (N_37895,N_33850,N_31958);
and U37896 (N_37896,N_31841,N_33253);
nand U37897 (N_37897,N_33502,N_33964);
nor U37898 (N_37898,N_30622,N_31369);
xnor U37899 (N_37899,N_34986,N_31720);
nor U37900 (N_37900,N_30721,N_31948);
nor U37901 (N_37901,N_34929,N_30640);
xnor U37902 (N_37902,N_33927,N_33971);
and U37903 (N_37903,N_34625,N_33249);
nand U37904 (N_37904,N_30373,N_34049);
and U37905 (N_37905,N_32878,N_32375);
xor U37906 (N_37906,N_34472,N_33165);
or U37907 (N_37907,N_33452,N_30271);
nand U37908 (N_37908,N_32754,N_34288);
nor U37909 (N_37909,N_32483,N_33098);
and U37910 (N_37910,N_33393,N_33941);
nand U37911 (N_37911,N_30196,N_34281);
nand U37912 (N_37912,N_34154,N_33810);
or U37913 (N_37913,N_31379,N_31543);
or U37914 (N_37914,N_34396,N_33752);
nor U37915 (N_37915,N_33910,N_31188);
or U37916 (N_37916,N_31694,N_34114);
or U37917 (N_37917,N_30017,N_31859);
nor U37918 (N_37918,N_34372,N_30855);
xor U37919 (N_37919,N_31061,N_32701);
or U37920 (N_37920,N_30958,N_34627);
or U37921 (N_37921,N_30071,N_31717);
nand U37922 (N_37922,N_33940,N_34895);
nor U37923 (N_37923,N_31386,N_31266);
xnor U37924 (N_37924,N_33008,N_30393);
xor U37925 (N_37925,N_34083,N_30282);
xor U37926 (N_37926,N_32623,N_32282);
and U37927 (N_37927,N_32284,N_33905);
xor U37928 (N_37928,N_30818,N_31282);
and U37929 (N_37929,N_30008,N_33530);
nor U37930 (N_37930,N_33353,N_31541);
and U37931 (N_37931,N_34434,N_32382);
xor U37932 (N_37932,N_31777,N_30759);
and U37933 (N_37933,N_31432,N_33356);
or U37934 (N_37934,N_33500,N_30119);
nor U37935 (N_37935,N_33662,N_31992);
or U37936 (N_37936,N_30768,N_32874);
or U37937 (N_37937,N_34932,N_33852);
nor U37938 (N_37938,N_34776,N_33169);
xor U37939 (N_37939,N_30585,N_34305);
or U37940 (N_37940,N_34734,N_31144);
or U37941 (N_37941,N_34594,N_30629);
or U37942 (N_37942,N_30641,N_32615);
xor U37943 (N_37943,N_34859,N_32983);
and U37944 (N_37944,N_30705,N_31583);
nand U37945 (N_37945,N_32572,N_32026);
nand U37946 (N_37946,N_34077,N_31021);
or U37947 (N_37947,N_31116,N_34258);
nor U37948 (N_37948,N_34734,N_32649);
and U37949 (N_37949,N_34781,N_30417);
or U37950 (N_37950,N_30653,N_30392);
and U37951 (N_37951,N_31324,N_34563);
and U37952 (N_37952,N_34682,N_33031);
and U37953 (N_37953,N_32106,N_33494);
nor U37954 (N_37954,N_33674,N_32759);
or U37955 (N_37955,N_34025,N_33054);
xor U37956 (N_37956,N_31533,N_31040);
and U37957 (N_37957,N_34055,N_32472);
xor U37958 (N_37958,N_30515,N_31727);
xnor U37959 (N_37959,N_34977,N_33467);
and U37960 (N_37960,N_34937,N_34400);
xnor U37961 (N_37961,N_31605,N_30222);
xor U37962 (N_37962,N_31479,N_31776);
or U37963 (N_37963,N_33125,N_30603);
nor U37964 (N_37964,N_32681,N_30664);
nor U37965 (N_37965,N_31802,N_33929);
or U37966 (N_37966,N_31922,N_34896);
and U37967 (N_37967,N_31188,N_30091);
nand U37968 (N_37968,N_31306,N_31131);
xnor U37969 (N_37969,N_34768,N_33799);
or U37970 (N_37970,N_34468,N_32965);
nor U37971 (N_37971,N_33789,N_33261);
nand U37972 (N_37972,N_34473,N_30215);
and U37973 (N_37973,N_31165,N_30249);
and U37974 (N_37974,N_34237,N_34265);
nand U37975 (N_37975,N_30478,N_30079);
nand U37976 (N_37976,N_31467,N_33056);
and U37977 (N_37977,N_33352,N_34261);
nor U37978 (N_37978,N_31943,N_33380);
nand U37979 (N_37979,N_30553,N_30321);
or U37980 (N_37980,N_33270,N_32960);
or U37981 (N_37981,N_30365,N_31748);
or U37982 (N_37982,N_32852,N_33171);
and U37983 (N_37983,N_34421,N_32404);
nand U37984 (N_37984,N_30017,N_33401);
nor U37985 (N_37985,N_32918,N_31550);
or U37986 (N_37986,N_30771,N_32631);
nand U37987 (N_37987,N_34862,N_32718);
or U37988 (N_37988,N_34510,N_31491);
nand U37989 (N_37989,N_32131,N_34886);
and U37990 (N_37990,N_34075,N_34353);
nand U37991 (N_37991,N_30117,N_33413);
xor U37992 (N_37992,N_33495,N_31535);
and U37993 (N_37993,N_32322,N_31369);
and U37994 (N_37994,N_34502,N_32563);
xnor U37995 (N_37995,N_31102,N_34776);
and U37996 (N_37996,N_32322,N_32290);
or U37997 (N_37997,N_30931,N_32014);
nor U37998 (N_37998,N_32799,N_33116);
nand U37999 (N_37999,N_30035,N_33370);
or U38000 (N_38000,N_33067,N_30693);
nand U38001 (N_38001,N_34547,N_33468);
or U38002 (N_38002,N_33284,N_33193);
nor U38003 (N_38003,N_30065,N_34481);
nor U38004 (N_38004,N_31771,N_32947);
nand U38005 (N_38005,N_33261,N_31772);
nor U38006 (N_38006,N_30920,N_32425);
xor U38007 (N_38007,N_30038,N_30640);
and U38008 (N_38008,N_34678,N_31212);
xnor U38009 (N_38009,N_32155,N_33024);
xor U38010 (N_38010,N_30060,N_31211);
or U38011 (N_38011,N_31143,N_31262);
and U38012 (N_38012,N_33335,N_33574);
or U38013 (N_38013,N_34509,N_31967);
or U38014 (N_38014,N_30162,N_31056);
nor U38015 (N_38015,N_34263,N_34758);
nand U38016 (N_38016,N_33256,N_30432);
nand U38017 (N_38017,N_31236,N_30338);
and U38018 (N_38018,N_33330,N_34281);
and U38019 (N_38019,N_32244,N_30426);
or U38020 (N_38020,N_32836,N_33043);
nand U38021 (N_38021,N_31008,N_30840);
nand U38022 (N_38022,N_33421,N_33650);
and U38023 (N_38023,N_33012,N_31803);
and U38024 (N_38024,N_31113,N_32700);
nor U38025 (N_38025,N_30237,N_32435);
xnor U38026 (N_38026,N_32079,N_30111);
and U38027 (N_38027,N_33563,N_33359);
xor U38028 (N_38028,N_31398,N_31952);
nor U38029 (N_38029,N_34116,N_31424);
or U38030 (N_38030,N_30808,N_30332);
or U38031 (N_38031,N_33529,N_32677);
nor U38032 (N_38032,N_31800,N_31655);
nor U38033 (N_38033,N_30842,N_32590);
nor U38034 (N_38034,N_33562,N_31639);
or U38035 (N_38035,N_33015,N_34094);
nor U38036 (N_38036,N_30007,N_30205);
xnor U38037 (N_38037,N_34343,N_33166);
nor U38038 (N_38038,N_30234,N_32230);
or U38039 (N_38039,N_33390,N_33019);
nand U38040 (N_38040,N_31808,N_33536);
nand U38041 (N_38041,N_30609,N_33022);
nor U38042 (N_38042,N_34754,N_30369);
and U38043 (N_38043,N_32568,N_33232);
or U38044 (N_38044,N_30066,N_31003);
and U38045 (N_38045,N_32829,N_32126);
nand U38046 (N_38046,N_30238,N_31170);
nor U38047 (N_38047,N_33279,N_31975);
nand U38048 (N_38048,N_30114,N_30504);
or U38049 (N_38049,N_31189,N_32456);
xor U38050 (N_38050,N_30041,N_30836);
nor U38051 (N_38051,N_31253,N_33265);
nand U38052 (N_38052,N_31708,N_33383);
or U38053 (N_38053,N_34436,N_30116);
nand U38054 (N_38054,N_33236,N_31652);
and U38055 (N_38055,N_34247,N_32701);
nand U38056 (N_38056,N_32279,N_31382);
and U38057 (N_38057,N_33262,N_33445);
and U38058 (N_38058,N_31441,N_34420);
and U38059 (N_38059,N_34146,N_32746);
nand U38060 (N_38060,N_31007,N_30058);
nor U38061 (N_38061,N_31523,N_30449);
xor U38062 (N_38062,N_32805,N_34739);
or U38063 (N_38063,N_32898,N_30848);
xor U38064 (N_38064,N_31124,N_34324);
and U38065 (N_38065,N_31043,N_31169);
nor U38066 (N_38066,N_30475,N_33900);
nand U38067 (N_38067,N_30936,N_30385);
nor U38068 (N_38068,N_33508,N_30606);
and U38069 (N_38069,N_32335,N_30112);
xnor U38070 (N_38070,N_31301,N_30010);
or U38071 (N_38071,N_31003,N_33172);
xnor U38072 (N_38072,N_32918,N_30060);
or U38073 (N_38073,N_33063,N_30654);
xor U38074 (N_38074,N_30249,N_32570);
nor U38075 (N_38075,N_32721,N_33626);
nand U38076 (N_38076,N_33092,N_33008);
nor U38077 (N_38077,N_33859,N_30103);
nand U38078 (N_38078,N_31504,N_30466);
nand U38079 (N_38079,N_30862,N_30369);
nor U38080 (N_38080,N_34018,N_34637);
xnor U38081 (N_38081,N_30920,N_33082);
nor U38082 (N_38082,N_30251,N_32404);
xnor U38083 (N_38083,N_32724,N_30025);
xor U38084 (N_38084,N_30051,N_33286);
and U38085 (N_38085,N_31763,N_31621);
nand U38086 (N_38086,N_31934,N_32524);
and U38087 (N_38087,N_31629,N_31569);
nand U38088 (N_38088,N_30262,N_32935);
xnor U38089 (N_38089,N_34003,N_33563);
xor U38090 (N_38090,N_34636,N_30397);
nand U38091 (N_38091,N_30285,N_32174);
nand U38092 (N_38092,N_32006,N_31537);
or U38093 (N_38093,N_32800,N_33383);
xor U38094 (N_38094,N_34925,N_32798);
or U38095 (N_38095,N_33172,N_34610);
or U38096 (N_38096,N_32648,N_31235);
and U38097 (N_38097,N_34512,N_34910);
or U38098 (N_38098,N_32967,N_32485);
nand U38099 (N_38099,N_34223,N_30757);
nand U38100 (N_38100,N_31250,N_33248);
xnor U38101 (N_38101,N_30474,N_34215);
nor U38102 (N_38102,N_30765,N_30382);
xnor U38103 (N_38103,N_30910,N_30816);
nand U38104 (N_38104,N_31539,N_32418);
or U38105 (N_38105,N_33242,N_33526);
nand U38106 (N_38106,N_34562,N_34189);
nor U38107 (N_38107,N_33420,N_31470);
nand U38108 (N_38108,N_31476,N_32660);
xor U38109 (N_38109,N_32519,N_31059);
xnor U38110 (N_38110,N_32881,N_33373);
or U38111 (N_38111,N_34215,N_32231);
or U38112 (N_38112,N_34252,N_32839);
nor U38113 (N_38113,N_32273,N_32906);
and U38114 (N_38114,N_34299,N_31468);
or U38115 (N_38115,N_32036,N_31655);
or U38116 (N_38116,N_34106,N_32258);
nor U38117 (N_38117,N_34352,N_34777);
or U38118 (N_38118,N_30892,N_33793);
nor U38119 (N_38119,N_32187,N_33770);
and U38120 (N_38120,N_34364,N_32568);
nand U38121 (N_38121,N_34671,N_32763);
nand U38122 (N_38122,N_34435,N_31002);
nor U38123 (N_38123,N_32735,N_33435);
and U38124 (N_38124,N_33692,N_33703);
or U38125 (N_38125,N_34432,N_30352);
or U38126 (N_38126,N_31833,N_30663);
or U38127 (N_38127,N_34168,N_30548);
nor U38128 (N_38128,N_34701,N_31869);
xor U38129 (N_38129,N_34379,N_32492);
nand U38130 (N_38130,N_31896,N_32996);
and U38131 (N_38131,N_30197,N_30243);
and U38132 (N_38132,N_31525,N_34360);
and U38133 (N_38133,N_32969,N_34042);
or U38134 (N_38134,N_30128,N_32147);
nor U38135 (N_38135,N_32272,N_31522);
or U38136 (N_38136,N_32883,N_30510);
xnor U38137 (N_38137,N_34457,N_31445);
and U38138 (N_38138,N_31696,N_33981);
xnor U38139 (N_38139,N_33736,N_30400);
xnor U38140 (N_38140,N_33494,N_30460);
or U38141 (N_38141,N_31196,N_34126);
and U38142 (N_38142,N_33498,N_32388);
xor U38143 (N_38143,N_30471,N_30608);
or U38144 (N_38144,N_32329,N_33277);
nor U38145 (N_38145,N_34635,N_32406);
xnor U38146 (N_38146,N_33059,N_30931);
or U38147 (N_38147,N_34433,N_30622);
nand U38148 (N_38148,N_32728,N_32753);
nor U38149 (N_38149,N_30716,N_31379);
and U38150 (N_38150,N_31478,N_30436);
nor U38151 (N_38151,N_34562,N_30799);
and U38152 (N_38152,N_34784,N_30704);
nor U38153 (N_38153,N_31656,N_32647);
and U38154 (N_38154,N_33910,N_32203);
nand U38155 (N_38155,N_34572,N_32774);
or U38156 (N_38156,N_30346,N_32854);
or U38157 (N_38157,N_31433,N_30614);
nand U38158 (N_38158,N_33396,N_34655);
xnor U38159 (N_38159,N_33776,N_31174);
or U38160 (N_38160,N_30765,N_34118);
or U38161 (N_38161,N_31546,N_31729);
nor U38162 (N_38162,N_33317,N_32959);
nand U38163 (N_38163,N_30734,N_31288);
xor U38164 (N_38164,N_33805,N_34338);
and U38165 (N_38165,N_33621,N_33498);
xnor U38166 (N_38166,N_34759,N_31485);
nand U38167 (N_38167,N_34561,N_33527);
nand U38168 (N_38168,N_31712,N_32097);
or U38169 (N_38169,N_30617,N_34964);
nor U38170 (N_38170,N_32185,N_34166);
and U38171 (N_38171,N_33601,N_32331);
and U38172 (N_38172,N_32347,N_31632);
nor U38173 (N_38173,N_34836,N_32792);
nor U38174 (N_38174,N_31800,N_31280);
or U38175 (N_38175,N_30688,N_34548);
xnor U38176 (N_38176,N_31967,N_31456);
or U38177 (N_38177,N_34856,N_34612);
nand U38178 (N_38178,N_33898,N_32001);
or U38179 (N_38179,N_33454,N_32856);
xnor U38180 (N_38180,N_34084,N_34538);
or U38181 (N_38181,N_31828,N_32607);
and U38182 (N_38182,N_34373,N_34245);
or U38183 (N_38183,N_31819,N_32077);
nand U38184 (N_38184,N_32734,N_34399);
nand U38185 (N_38185,N_32238,N_30496);
nand U38186 (N_38186,N_33948,N_31314);
or U38187 (N_38187,N_34134,N_30117);
and U38188 (N_38188,N_34509,N_31833);
xnor U38189 (N_38189,N_33600,N_33697);
nor U38190 (N_38190,N_31615,N_32384);
nand U38191 (N_38191,N_31431,N_31565);
nor U38192 (N_38192,N_33900,N_32676);
nor U38193 (N_38193,N_30690,N_30811);
and U38194 (N_38194,N_32122,N_32615);
nor U38195 (N_38195,N_30401,N_33474);
xnor U38196 (N_38196,N_32871,N_33069);
or U38197 (N_38197,N_31586,N_30363);
nand U38198 (N_38198,N_30918,N_32564);
nor U38199 (N_38199,N_32623,N_30822);
nor U38200 (N_38200,N_31372,N_32602);
or U38201 (N_38201,N_31667,N_31650);
and U38202 (N_38202,N_31995,N_34250);
and U38203 (N_38203,N_34172,N_31788);
nand U38204 (N_38204,N_34826,N_31052);
xnor U38205 (N_38205,N_31089,N_30279);
or U38206 (N_38206,N_31100,N_33180);
and U38207 (N_38207,N_33432,N_34712);
or U38208 (N_38208,N_31380,N_30922);
or U38209 (N_38209,N_30378,N_33781);
nor U38210 (N_38210,N_34322,N_32703);
or U38211 (N_38211,N_32041,N_30093);
nor U38212 (N_38212,N_30709,N_31430);
and U38213 (N_38213,N_31793,N_32307);
nand U38214 (N_38214,N_34818,N_31973);
nand U38215 (N_38215,N_33482,N_33637);
nand U38216 (N_38216,N_34777,N_34796);
nor U38217 (N_38217,N_34162,N_33658);
xor U38218 (N_38218,N_32990,N_33955);
nand U38219 (N_38219,N_33144,N_32507);
nor U38220 (N_38220,N_30541,N_31267);
nor U38221 (N_38221,N_34014,N_32260);
nor U38222 (N_38222,N_32623,N_31516);
nor U38223 (N_38223,N_33573,N_30553);
nand U38224 (N_38224,N_33540,N_30203);
nor U38225 (N_38225,N_31616,N_33093);
and U38226 (N_38226,N_32171,N_33455);
xnor U38227 (N_38227,N_34725,N_32909);
and U38228 (N_38228,N_31719,N_30511);
or U38229 (N_38229,N_30478,N_33919);
or U38230 (N_38230,N_32616,N_34671);
xnor U38231 (N_38231,N_34260,N_31712);
nor U38232 (N_38232,N_31110,N_34655);
nand U38233 (N_38233,N_30507,N_32571);
nand U38234 (N_38234,N_32446,N_33579);
or U38235 (N_38235,N_33060,N_34878);
nor U38236 (N_38236,N_30808,N_31585);
nor U38237 (N_38237,N_32453,N_30576);
or U38238 (N_38238,N_31874,N_34087);
or U38239 (N_38239,N_34989,N_34588);
nor U38240 (N_38240,N_32407,N_34864);
nor U38241 (N_38241,N_31196,N_30194);
nand U38242 (N_38242,N_31874,N_31915);
or U38243 (N_38243,N_30674,N_33282);
nor U38244 (N_38244,N_30288,N_31260);
xnor U38245 (N_38245,N_32151,N_32028);
and U38246 (N_38246,N_31256,N_30800);
or U38247 (N_38247,N_30520,N_30413);
nand U38248 (N_38248,N_33424,N_34390);
nor U38249 (N_38249,N_30333,N_30304);
and U38250 (N_38250,N_30218,N_32304);
nand U38251 (N_38251,N_31116,N_32675);
nor U38252 (N_38252,N_33586,N_32951);
nand U38253 (N_38253,N_31625,N_31800);
nor U38254 (N_38254,N_34350,N_32256);
and U38255 (N_38255,N_31410,N_31495);
and U38256 (N_38256,N_32083,N_33054);
or U38257 (N_38257,N_34303,N_32734);
nor U38258 (N_38258,N_32818,N_32348);
or U38259 (N_38259,N_33239,N_34817);
xnor U38260 (N_38260,N_31517,N_31123);
and U38261 (N_38261,N_32148,N_30883);
and U38262 (N_38262,N_30294,N_33642);
nor U38263 (N_38263,N_34617,N_32990);
and U38264 (N_38264,N_33709,N_32107);
nand U38265 (N_38265,N_31209,N_34468);
or U38266 (N_38266,N_32271,N_33061);
xor U38267 (N_38267,N_32985,N_33894);
and U38268 (N_38268,N_33368,N_30916);
nand U38269 (N_38269,N_31660,N_32244);
or U38270 (N_38270,N_32569,N_33307);
or U38271 (N_38271,N_31987,N_34613);
and U38272 (N_38272,N_32865,N_32732);
or U38273 (N_38273,N_32717,N_32171);
xor U38274 (N_38274,N_31381,N_34747);
xor U38275 (N_38275,N_31441,N_30573);
nor U38276 (N_38276,N_33628,N_32318);
xor U38277 (N_38277,N_30933,N_32016);
xor U38278 (N_38278,N_32206,N_33181);
or U38279 (N_38279,N_33253,N_32333);
xor U38280 (N_38280,N_34767,N_31321);
nor U38281 (N_38281,N_34517,N_33290);
nand U38282 (N_38282,N_34449,N_33916);
nor U38283 (N_38283,N_32048,N_32226);
xnor U38284 (N_38284,N_31804,N_33887);
and U38285 (N_38285,N_32836,N_33544);
nand U38286 (N_38286,N_31179,N_31340);
nand U38287 (N_38287,N_33479,N_33729);
or U38288 (N_38288,N_34910,N_30052);
xor U38289 (N_38289,N_31634,N_33779);
and U38290 (N_38290,N_31301,N_34993);
nor U38291 (N_38291,N_34105,N_31115);
xor U38292 (N_38292,N_33578,N_33699);
nand U38293 (N_38293,N_34476,N_32694);
xor U38294 (N_38294,N_32907,N_34663);
xnor U38295 (N_38295,N_32138,N_31723);
or U38296 (N_38296,N_30060,N_31264);
or U38297 (N_38297,N_33985,N_30958);
and U38298 (N_38298,N_31291,N_30315);
and U38299 (N_38299,N_33706,N_30255);
nor U38300 (N_38300,N_31544,N_33511);
or U38301 (N_38301,N_31601,N_31298);
or U38302 (N_38302,N_32138,N_32123);
and U38303 (N_38303,N_34291,N_33558);
and U38304 (N_38304,N_31514,N_30821);
or U38305 (N_38305,N_32413,N_32824);
nand U38306 (N_38306,N_31086,N_32510);
nor U38307 (N_38307,N_33363,N_31417);
or U38308 (N_38308,N_34294,N_33276);
xnor U38309 (N_38309,N_33217,N_33304);
xnor U38310 (N_38310,N_32203,N_33281);
nand U38311 (N_38311,N_31070,N_31126);
xor U38312 (N_38312,N_33640,N_33013);
nand U38313 (N_38313,N_34812,N_31434);
and U38314 (N_38314,N_32201,N_32301);
xnor U38315 (N_38315,N_32303,N_31559);
xor U38316 (N_38316,N_33508,N_30099);
and U38317 (N_38317,N_32603,N_30018);
or U38318 (N_38318,N_32107,N_32696);
nand U38319 (N_38319,N_30961,N_30159);
nor U38320 (N_38320,N_33127,N_30949);
nand U38321 (N_38321,N_34177,N_31193);
xor U38322 (N_38322,N_33773,N_34913);
nor U38323 (N_38323,N_33766,N_33603);
or U38324 (N_38324,N_30071,N_32896);
nand U38325 (N_38325,N_34890,N_30603);
nand U38326 (N_38326,N_33281,N_33443);
and U38327 (N_38327,N_31318,N_34693);
nor U38328 (N_38328,N_30105,N_31420);
nor U38329 (N_38329,N_30005,N_31885);
and U38330 (N_38330,N_30681,N_33276);
or U38331 (N_38331,N_34920,N_33996);
xnor U38332 (N_38332,N_31891,N_33421);
or U38333 (N_38333,N_34508,N_32606);
nor U38334 (N_38334,N_30970,N_34089);
nor U38335 (N_38335,N_34865,N_34154);
xnor U38336 (N_38336,N_32346,N_32511);
or U38337 (N_38337,N_31280,N_34560);
nor U38338 (N_38338,N_30747,N_31220);
xor U38339 (N_38339,N_32221,N_34167);
nor U38340 (N_38340,N_30828,N_31070);
nor U38341 (N_38341,N_34666,N_33538);
or U38342 (N_38342,N_34694,N_30345);
xor U38343 (N_38343,N_32609,N_31905);
nor U38344 (N_38344,N_32892,N_31973);
nand U38345 (N_38345,N_31262,N_31957);
nand U38346 (N_38346,N_31682,N_33194);
xnor U38347 (N_38347,N_32881,N_31576);
xor U38348 (N_38348,N_30377,N_30126);
nor U38349 (N_38349,N_32724,N_30930);
xnor U38350 (N_38350,N_34976,N_33007);
nand U38351 (N_38351,N_30322,N_34756);
and U38352 (N_38352,N_33303,N_31793);
or U38353 (N_38353,N_34637,N_32886);
nand U38354 (N_38354,N_30355,N_31009);
xor U38355 (N_38355,N_32048,N_32992);
and U38356 (N_38356,N_34437,N_32345);
nand U38357 (N_38357,N_31038,N_33567);
and U38358 (N_38358,N_30734,N_32474);
nor U38359 (N_38359,N_30241,N_32889);
and U38360 (N_38360,N_34876,N_34436);
xor U38361 (N_38361,N_32344,N_30582);
or U38362 (N_38362,N_30324,N_32669);
nand U38363 (N_38363,N_30864,N_32675);
nor U38364 (N_38364,N_30779,N_30185);
or U38365 (N_38365,N_32116,N_33438);
and U38366 (N_38366,N_31097,N_32553);
and U38367 (N_38367,N_32025,N_34996);
or U38368 (N_38368,N_32009,N_34520);
nor U38369 (N_38369,N_31819,N_31320);
nor U38370 (N_38370,N_31322,N_34240);
nor U38371 (N_38371,N_30068,N_31393);
xnor U38372 (N_38372,N_30809,N_30802);
nand U38373 (N_38373,N_32702,N_34034);
or U38374 (N_38374,N_33063,N_33417);
and U38375 (N_38375,N_32538,N_33430);
nand U38376 (N_38376,N_33199,N_31788);
nor U38377 (N_38377,N_34260,N_31705);
nor U38378 (N_38378,N_31300,N_34973);
and U38379 (N_38379,N_33437,N_30889);
or U38380 (N_38380,N_33787,N_33318);
or U38381 (N_38381,N_31180,N_32818);
or U38382 (N_38382,N_30233,N_33217);
or U38383 (N_38383,N_32110,N_30175);
nand U38384 (N_38384,N_31161,N_34610);
and U38385 (N_38385,N_30048,N_34648);
nor U38386 (N_38386,N_32631,N_34657);
nand U38387 (N_38387,N_30202,N_34929);
xor U38388 (N_38388,N_31341,N_33723);
xor U38389 (N_38389,N_30982,N_30631);
xor U38390 (N_38390,N_32834,N_32337);
and U38391 (N_38391,N_33801,N_33748);
or U38392 (N_38392,N_33172,N_30122);
xor U38393 (N_38393,N_31056,N_34927);
xor U38394 (N_38394,N_32223,N_32465);
xor U38395 (N_38395,N_33429,N_31921);
xor U38396 (N_38396,N_30106,N_32097);
nand U38397 (N_38397,N_31096,N_31594);
xnor U38398 (N_38398,N_33363,N_30595);
nand U38399 (N_38399,N_34249,N_31588);
nor U38400 (N_38400,N_31212,N_33752);
nor U38401 (N_38401,N_34759,N_33343);
and U38402 (N_38402,N_31243,N_30992);
nor U38403 (N_38403,N_32243,N_34917);
nor U38404 (N_38404,N_32001,N_34066);
nand U38405 (N_38405,N_31558,N_33228);
or U38406 (N_38406,N_31241,N_33529);
xnor U38407 (N_38407,N_32907,N_33997);
or U38408 (N_38408,N_34010,N_32302);
nand U38409 (N_38409,N_31467,N_33386);
nor U38410 (N_38410,N_32832,N_33934);
nor U38411 (N_38411,N_32733,N_31007);
nor U38412 (N_38412,N_33487,N_34755);
xnor U38413 (N_38413,N_34918,N_31366);
nor U38414 (N_38414,N_31129,N_34383);
nand U38415 (N_38415,N_34810,N_32883);
or U38416 (N_38416,N_32788,N_31005);
nand U38417 (N_38417,N_31733,N_34696);
xor U38418 (N_38418,N_30248,N_33640);
xor U38419 (N_38419,N_32067,N_33832);
nand U38420 (N_38420,N_30571,N_32011);
and U38421 (N_38421,N_34663,N_33066);
and U38422 (N_38422,N_32031,N_30314);
or U38423 (N_38423,N_33842,N_34614);
or U38424 (N_38424,N_32648,N_31340);
nand U38425 (N_38425,N_33586,N_33611);
xor U38426 (N_38426,N_32003,N_32316);
nand U38427 (N_38427,N_33970,N_31046);
xor U38428 (N_38428,N_33995,N_32051);
or U38429 (N_38429,N_32328,N_34648);
nand U38430 (N_38430,N_33490,N_34900);
nor U38431 (N_38431,N_34551,N_32729);
and U38432 (N_38432,N_31989,N_30776);
or U38433 (N_38433,N_31544,N_31039);
nor U38434 (N_38434,N_32939,N_34655);
or U38435 (N_38435,N_30254,N_31971);
xor U38436 (N_38436,N_34531,N_34456);
nor U38437 (N_38437,N_34858,N_32864);
and U38438 (N_38438,N_34849,N_34629);
and U38439 (N_38439,N_31054,N_34837);
and U38440 (N_38440,N_32956,N_30477);
xnor U38441 (N_38441,N_30431,N_31465);
and U38442 (N_38442,N_31591,N_30669);
or U38443 (N_38443,N_32406,N_31476);
and U38444 (N_38444,N_31642,N_32143);
nand U38445 (N_38445,N_32872,N_30366);
or U38446 (N_38446,N_34109,N_30798);
or U38447 (N_38447,N_34718,N_31664);
xnor U38448 (N_38448,N_30561,N_34730);
and U38449 (N_38449,N_33831,N_31719);
and U38450 (N_38450,N_34442,N_30674);
nand U38451 (N_38451,N_32405,N_30405);
nand U38452 (N_38452,N_31576,N_34260);
xnor U38453 (N_38453,N_32420,N_30057);
nor U38454 (N_38454,N_32948,N_33578);
and U38455 (N_38455,N_33152,N_31071);
xnor U38456 (N_38456,N_31687,N_33698);
or U38457 (N_38457,N_31751,N_32010);
xnor U38458 (N_38458,N_33244,N_33436);
nand U38459 (N_38459,N_32082,N_30674);
or U38460 (N_38460,N_34043,N_30956);
or U38461 (N_38461,N_34813,N_31162);
nand U38462 (N_38462,N_32550,N_34723);
and U38463 (N_38463,N_30762,N_33410);
or U38464 (N_38464,N_34180,N_34345);
or U38465 (N_38465,N_34822,N_31727);
xor U38466 (N_38466,N_31659,N_31712);
nand U38467 (N_38467,N_30130,N_34620);
and U38468 (N_38468,N_30322,N_33541);
xor U38469 (N_38469,N_34332,N_31639);
nor U38470 (N_38470,N_31849,N_31367);
nand U38471 (N_38471,N_33788,N_34101);
nor U38472 (N_38472,N_30304,N_34969);
xor U38473 (N_38473,N_31357,N_33800);
nand U38474 (N_38474,N_31742,N_32433);
nand U38475 (N_38475,N_32024,N_33667);
nor U38476 (N_38476,N_30656,N_34875);
or U38477 (N_38477,N_34715,N_32461);
xnor U38478 (N_38478,N_34254,N_32437);
xor U38479 (N_38479,N_34563,N_34595);
nand U38480 (N_38480,N_34914,N_30402);
xnor U38481 (N_38481,N_34105,N_30581);
xnor U38482 (N_38482,N_31412,N_32512);
nand U38483 (N_38483,N_32295,N_34072);
or U38484 (N_38484,N_30172,N_33360);
nor U38485 (N_38485,N_34607,N_32686);
xor U38486 (N_38486,N_31721,N_30875);
nor U38487 (N_38487,N_31342,N_31314);
or U38488 (N_38488,N_31616,N_31252);
or U38489 (N_38489,N_34802,N_32960);
and U38490 (N_38490,N_31856,N_33044);
xnor U38491 (N_38491,N_34897,N_33214);
or U38492 (N_38492,N_32394,N_34411);
nand U38493 (N_38493,N_31564,N_32527);
or U38494 (N_38494,N_31911,N_34261);
or U38495 (N_38495,N_30658,N_31168);
or U38496 (N_38496,N_31079,N_34459);
xnor U38497 (N_38497,N_32225,N_30834);
and U38498 (N_38498,N_30751,N_31171);
and U38499 (N_38499,N_32702,N_34245);
or U38500 (N_38500,N_30318,N_32064);
xor U38501 (N_38501,N_34051,N_32359);
or U38502 (N_38502,N_30785,N_31020);
nor U38503 (N_38503,N_32671,N_34642);
xnor U38504 (N_38504,N_31365,N_33126);
or U38505 (N_38505,N_30619,N_33875);
nor U38506 (N_38506,N_32723,N_31839);
and U38507 (N_38507,N_34406,N_32010);
and U38508 (N_38508,N_31838,N_34436);
xor U38509 (N_38509,N_31104,N_30756);
xnor U38510 (N_38510,N_32237,N_34429);
and U38511 (N_38511,N_30670,N_30693);
nand U38512 (N_38512,N_31288,N_34969);
and U38513 (N_38513,N_34433,N_30528);
nor U38514 (N_38514,N_31651,N_33353);
and U38515 (N_38515,N_32497,N_31441);
and U38516 (N_38516,N_31219,N_33615);
nand U38517 (N_38517,N_34986,N_33206);
or U38518 (N_38518,N_34237,N_33730);
and U38519 (N_38519,N_30348,N_30035);
or U38520 (N_38520,N_34315,N_33701);
and U38521 (N_38521,N_33182,N_32564);
xor U38522 (N_38522,N_30766,N_34118);
nand U38523 (N_38523,N_33163,N_33098);
nand U38524 (N_38524,N_31757,N_34672);
nor U38525 (N_38525,N_33059,N_31626);
xor U38526 (N_38526,N_34342,N_34716);
nand U38527 (N_38527,N_31597,N_30401);
and U38528 (N_38528,N_31514,N_30076);
and U38529 (N_38529,N_34639,N_32901);
xor U38530 (N_38530,N_33116,N_30861);
nand U38531 (N_38531,N_33401,N_31528);
xor U38532 (N_38532,N_34932,N_32588);
xor U38533 (N_38533,N_32079,N_30497);
or U38534 (N_38534,N_33250,N_33208);
xnor U38535 (N_38535,N_34948,N_32118);
and U38536 (N_38536,N_34336,N_32082);
nor U38537 (N_38537,N_32597,N_32172);
nand U38538 (N_38538,N_31044,N_33162);
xnor U38539 (N_38539,N_34200,N_32860);
nand U38540 (N_38540,N_32488,N_31298);
nand U38541 (N_38541,N_31848,N_33123);
xor U38542 (N_38542,N_32632,N_33740);
and U38543 (N_38543,N_32436,N_33602);
nand U38544 (N_38544,N_31769,N_30850);
and U38545 (N_38545,N_34400,N_30011);
nand U38546 (N_38546,N_33918,N_31595);
xnor U38547 (N_38547,N_30903,N_34651);
nand U38548 (N_38548,N_32266,N_34090);
nor U38549 (N_38549,N_31840,N_30737);
nor U38550 (N_38550,N_30394,N_34033);
or U38551 (N_38551,N_30958,N_30797);
and U38552 (N_38552,N_32167,N_31595);
xor U38553 (N_38553,N_32817,N_34888);
and U38554 (N_38554,N_30262,N_34173);
xnor U38555 (N_38555,N_30577,N_31165);
and U38556 (N_38556,N_31508,N_32706);
nor U38557 (N_38557,N_30417,N_33393);
and U38558 (N_38558,N_34829,N_32452);
nor U38559 (N_38559,N_31952,N_34957);
or U38560 (N_38560,N_30133,N_31605);
nor U38561 (N_38561,N_34769,N_32542);
nor U38562 (N_38562,N_31334,N_33432);
xnor U38563 (N_38563,N_31981,N_33460);
xnor U38564 (N_38564,N_32952,N_34654);
nor U38565 (N_38565,N_30651,N_31632);
and U38566 (N_38566,N_34100,N_31973);
and U38567 (N_38567,N_33913,N_33363);
nand U38568 (N_38568,N_33276,N_33358);
nand U38569 (N_38569,N_30179,N_33848);
nor U38570 (N_38570,N_30493,N_31681);
xor U38571 (N_38571,N_33821,N_32483);
xnor U38572 (N_38572,N_30369,N_31951);
and U38573 (N_38573,N_30133,N_34319);
or U38574 (N_38574,N_31909,N_31289);
or U38575 (N_38575,N_33117,N_34400);
and U38576 (N_38576,N_33365,N_31649);
nand U38577 (N_38577,N_33397,N_33614);
or U38578 (N_38578,N_32266,N_34466);
or U38579 (N_38579,N_31007,N_32070);
nand U38580 (N_38580,N_32589,N_31803);
nor U38581 (N_38581,N_34789,N_34549);
xnor U38582 (N_38582,N_32866,N_30150);
xnor U38583 (N_38583,N_31848,N_33561);
nand U38584 (N_38584,N_33269,N_33428);
xnor U38585 (N_38585,N_31928,N_33233);
nand U38586 (N_38586,N_33741,N_32504);
and U38587 (N_38587,N_34265,N_32993);
nand U38588 (N_38588,N_33305,N_30803);
nor U38589 (N_38589,N_32669,N_32869);
nand U38590 (N_38590,N_34919,N_32028);
and U38591 (N_38591,N_32145,N_33382);
xnor U38592 (N_38592,N_32628,N_30070);
or U38593 (N_38593,N_31558,N_31938);
and U38594 (N_38594,N_32129,N_30124);
or U38595 (N_38595,N_32675,N_34539);
xor U38596 (N_38596,N_34359,N_34345);
nand U38597 (N_38597,N_31536,N_30528);
or U38598 (N_38598,N_30552,N_33725);
xnor U38599 (N_38599,N_32319,N_32427);
nor U38600 (N_38600,N_30596,N_32020);
xor U38601 (N_38601,N_31467,N_33311);
or U38602 (N_38602,N_33568,N_32350);
xnor U38603 (N_38603,N_33264,N_34896);
nor U38604 (N_38604,N_34041,N_33985);
nand U38605 (N_38605,N_33766,N_31869);
xnor U38606 (N_38606,N_30811,N_33147);
nor U38607 (N_38607,N_33499,N_34244);
or U38608 (N_38608,N_34536,N_34799);
and U38609 (N_38609,N_32986,N_34124);
nor U38610 (N_38610,N_32318,N_32090);
nor U38611 (N_38611,N_32852,N_30638);
nor U38612 (N_38612,N_33727,N_33946);
nor U38613 (N_38613,N_30403,N_30363);
or U38614 (N_38614,N_33520,N_31704);
and U38615 (N_38615,N_30310,N_33351);
and U38616 (N_38616,N_31660,N_34318);
and U38617 (N_38617,N_32580,N_33392);
or U38618 (N_38618,N_34365,N_34747);
nand U38619 (N_38619,N_31655,N_32024);
and U38620 (N_38620,N_30631,N_33471);
nor U38621 (N_38621,N_31874,N_34464);
nand U38622 (N_38622,N_32380,N_32651);
xor U38623 (N_38623,N_30812,N_30610);
nor U38624 (N_38624,N_30219,N_30575);
and U38625 (N_38625,N_34962,N_33739);
xnor U38626 (N_38626,N_34252,N_33782);
nand U38627 (N_38627,N_30002,N_34023);
xor U38628 (N_38628,N_30085,N_34431);
nor U38629 (N_38629,N_33414,N_30405);
xnor U38630 (N_38630,N_31122,N_30861);
xnor U38631 (N_38631,N_34172,N_31588);
or U38632 (N_38632,N_33985,N_31499);
and U38633 (N_38633,N_31855,N_34184);
nand U38634 (N_38634,N_33762,N_32514);
xor U38635 (N_38635,N_31221,N_33205);
nand U38636 (N_38636,N_30532,N_32731);
nand U38637 (N_38637,N_32545,N_31506);
nor U38638 (N_38638,N_30808,N_33118);
or U38639 (N_38639,N_34668,N_32556);
nand U38640 (N_38640,N_33665,N_30607);
or U38641 (N_38641,N_34092,N_34670);
nor U38642 (N_38642,N_32413,N_34101);
xnor U38643 (N_38643,N_31865,N_31450);
nand U38644 (N_38644,N_32177,N_31437);
or U38645 (N_38645,N_30583,N_32469);
or U38646 (N_38646,N_33860,N_31858);
or U38647 (N_38647,N_33661,N_34694);
xor U38648 (N_38648,N_33981,N_30923);
nand U38649 (N_38649,N_31359,N_30427);
xor U38650 (N_38650,N_32756,N_34834);
nor U38651 (N_38651,N_34589,N_31830);
nor U38652 (N_38652,N_34767,N_34681);
xnor U38653 (N_38653,N_34039,N_32502);
or U38654 (N_38654,N_33795,N_30776);
nor U38655 (N_38655,N_34367,N_30686);
nand U38656 (N_38656,N_32844,N_30870);
nand U38657 (N_38657,N_34024,N_34000);
xnor U38658 (N_38658,N_33262,N_31719);
nand U38659 (N_38659,N_33266,N_31140);
nor U38660 (N_38660,N_30048,N_30800);
nor U38661 (N_38661,N_33772,N_34796);
and U38662 (N_38662,N_34611,N_32407);
nand U38663 (N_38663,N_33518,N_32122);
nand U38664 (N_38664,N_32262,N_33128);
nor U38665 (N_38665,N_34627,N_30051);
and U38666 (N_38666,N_31904,N_31398);
nand U38667 (N_38667,N_31913,N_33540);
or U38668 (N_38668,N_32784,N_31710);
and U38669 (N_38669,N_32277,N_33388);
xor U38670 (N_38670,N_33119,N_32710);
xnor U38671 (N_38671,N_32648,N_34384);
nor U38672 (N_38672,N_30824,N_32835);
or U38673 (N_38673,N_33197,N_31642);
xnor U38674 (N_38674,N_34226,N_30612);
or U38675 (N_38675,N_34777,N_30344);
and U38676 (N_38676,N_30499,N_34378);
or U38677 (N_38677,N_34698,N_33309);
and U38678 (N_38678,N_32545,N_30512);
nand U38679 (N_38679,N_31505,N_34939);
and U38680 (N_38680,N_30358,N_33242);
xnor U38681 (N_38681,N_33937,N_33094);
nor U38682 (N_38682,N_32170,N_31457);
xnor U38683 (N_38683,N_30556,N_33533);
xor U38684 (N_38684,N_32467,N_32512);
and U38685 (N_38685,N_34721,N_30405);
xor U38686 (N_38686,N_31121,N_31160);
nand U38687 (N_38687,N_33964,N_33635);
nor U38688 (N_38688,N_30782,N_34918);
nor U38689 (N_38689,N_34630,N_30560);
or U38690 (N_38690,N_31854,N_32912);
or U38691 (N_38691,N_31505,N_32397);
or U38692 (N_38692,N_31391,N_32556);
or U38693 (N_38693,N_31294,N_30535);
nand U38694 (N_38694,N_30257,N_34192);
and U38695 (N_38695,N_30448,N_31618);
and U38696 (N_38696,N_34388,N_30469);
xor U38697 (N_38697,N_33535,N_32037);
and U38698 (N_38698,N_34664,N_33037);
xnor U38699 (N_38699,N_31671,N_31015);
or U38700 (N_38700,N_34431,N_31368);
or U38701 (N_38701,N_31333,N_32058);
nor U38702 (N_38702,N_31274,N_31306);
xor U38703 (N_38703,N_33866,N_31852);
xor U38704 (N_38704,N_32662,N_31789);
xor U38705 (N_38705,N_32920,N_30563);
nor U38706 (N_38706,N_33485,N_30569);
xor U38707 (N_38707,N_33914,N_31146);
xnor U38708 (N_38708,N_31160,N_30770);
nand U38709 (N_38709,N_33638,N_32860);
nand U38710 (N_38710,N_31217,N_31019);
xor U38711 (N_38711,N_32427,N_33119);
xor U38712 (N_38712,N_34632,N_32090);
xor U38713 (N_38713,N_31907,N_34238);
or U38714 (N_38714,N_30936,N_30051);
and U38715 (N_38715,N_30494,N_30053);
xnor U38716 (N_38716,N_34523,N_33538);
or U38717 (N_38717,N_32618,N_34215);
and U38718 (N_38718,N_32198,N_31293);
xor U38719 (N_38719,N_34390,N_32626);
and U38720 (N_38720,N_32622,N_31898);
and U38721 (N_38721,N_30912,N_34967);
nor U38722 (N_38722,N_32205,N_31374);
xor U38723 (N_38723,N_33008,N_33523);
and U38724 (N_38724,N_34070,N_33808);
xor U38725 (N_38725,N_32454,N_31908);
and U38726 (N_38726,N_30785,N_30629);
or U38727 (N_38727,N_32193,N_30470);
nand U38728 (N_38728,N_33919,N_31917);
or U38729 (N_38729,N_31010,N_33701);
and U38730 (N_38730,N_33675,N_31244);
and U38731 (N_38731,N_34285,N_30067);
and U38732 (N_38732,N_33489,N_34604);
or U38733 (N_38733,N_30952,N_33521);
nand U38734 (N_38734,N_30252,N_32193);
and U38735 (N_38735,N_32863,N_32548);
and U38736 (N_38736,N_30908,N_30197);
nor U38737 (N_38737,N_31608,N_32301);
nor U38738 (N_38738,N_34272,N_34069);
and U38739 (N_38739,N_31160,N_33369);
and U38740 (N_38740,N_34336,N_32269);
or U38741 (N_38741,N_33636,N_31544);
xnor U38742 (N_38742,N_30639,N_32189);
xor U38743 (N_38743,N_34414,N_32946);
and U38744 (N_38744,N_33939,N_31026);
and U38745 (N_38745,N_33459,N_30800);
and U38746 (N_38746,N_31645,N_33361);
xor U38747 (N_38747,N_31628,N_33473);
or U38748 (N_38748,N_31442,N_34622);
or U38749 (N_38749,N_32325,N_33216);
nand U38750 (N_38750,N_34333,N_33013);
nand U38751 (N_38751,N_34887,N_33990);
and U38752 (N_38752,N_32960,N_33669);
or U38753 (N_38753,N_30238,N_31324);
nand U38754 (N_38754,N_32960,N_32681);
and U38755 (N_38755,N_32254,N_30414);
or U38756 (N_38756,N_34944,N_31128);
nor U38757 (N_38757,N_33267,N_30314);
xnor U38758 (N_38758,N_31783,N_33413);
or U38759 (N_38759,N_32389,N_33582);
or U38760 (N_38760,N_31050,N_34264);
xor U38761 (N_38761,N_33631,N_33451);
xor U38762 (N_38762,N_33585,N_31568);
nand U38763 (N_38763,N_32285,N_30887);
nand U38764 (N_38764,N_33548,N_31622);
and U38765 (N_38765,N_34134,N_33790);
or U38766 (N_38766,N_32223,N_32733);
and U38767 (N_38767,N_32471,N_33735);
xor U38768 (N_38768,N_33122,N_30202);
nand U38769 (N_38769,N_31736,N_34456);
nand U38770 (N_38770,N_32603,N_31237);
nand U38771 (N_38771,N_32259,N_30396);
nand U38772 (N_38772,N_34739,N_32641);
and U38773 (N_38773,N_30054,N_33438);
nor U38774 (N_38774,N_30286,N_31783);
nand U38775 (N_38775,N_32977,N_34192);
nand U38776 (N_38776,N_31980,N_30188);
nand U38777 (N_38777,N_30591,N_34343);
xnor U38778 (N_38778,N_30924,N_30490);
nand U38779 (N_38779,N_31581,N_30993);
and U38780 (N_38780,N_31772,N_32616);
xor U38781 (N_38781,N_33722,N_31877);
or U38782 (N_38782,N_33599,N_30413);
or U38783 (N_38783,N_32315,N_33972);
nand U38784 (N_38784,N_34400,N_33510);
xnor U38785 (N_38785,N_33880,N_32689);
and U38786 (N_38786,N_34142,N_31855);
xnor U38787 (N_38787,N_34741,N_33112);
and U38788 (N_38788,N_32010,N_30592);
or U38789 (N_38789,N_31940,N_31702);
nor U38790 (N_38790,N_32789,N_33892);
and U38791 (N_38791,N_32118,N_34375);
and U38792 (N_38792,N_34157,N_34199);
and U38793 (N_38793,N_30566,N_31005);
or U38794 (N_38794,N_34783,N_32965);
and U38795 (N_38795,N_34319,N_31683);
and U38796 (N_38796,N_31269,N_31569);
nand U38797 (N_38797,N_31815,N_32012);
nand U38798 (N_38798,N_30608,N_32887);
nand U38799 (N_38799,N_33853,N_34213);
nand U38800 (N_38800,N_32422,N_30280);
and U38801 (N_38801,N_34743,N_30437);
or U38802 (N_38802,N_34404,N_30689);
xnor U38803 (N_38803,N_33730,N_30074);
nor U38804 (N_38804,N_33731,N_34773);
nor U38805 (N_38805,N_34675,N_31127);
or U38806 (N_38806,N_34860,N_33961);
xor U38807 (N_38807,N_33356,N_32430);
nand U38808 (N_38808,N_32090,N_31432);
nand U38809 (N_38809,N_32699,N_31451);
or U38810 (N_38810,N_32339,N_33637);
and U38811 (N_38811,N_32775,N_31704);
nand U38812 (N_38812,N_31396,N_30707);
and U38813 (N_38813,N_32612,N_33798);
and U38814 (N_38814,N_32838,N_32864);
nor U38815 (N_38815,N_30478,N_34230);
nor U38816 (N_38816,N_32490,N_33911);
nand U38817 (N_38817,N_30725,N_32851);
or U38818 (N_38818,N_33619,N_34722);
or U38819 (N_38819,N_31031,N_32938);
and U38820 (N_38820,N_32707,N_31762);
or U38821 (N_38821,N_30223,N_31771);
or U38822 (N_38822,N_31006,N_32822);
nand U38823 (N_38823,N_34461,N_31449);
nand U38824 (N_38824,N_32615,N_34214);
or U38825 (N_38825,N_34836,N_33179);
nor U38826 (N_38826,N_34667,N_31497);
or U38827 (N_38827,N_33087,N_33973);
xor U38828 (N_38828,N_33055,N_34862);
nor U38829 (N_38829,N_34056,N_32263);
nor U38830 (N_38830,N_32816,N_32810);
nor U38831 (N_38831,N_30946,N_30590);
or U38832 (N_38832,N_30497,N_32475);
nor U38833 (N_38833,N_30257,N_34898);
and U38834 (N_38834,N_31747,N_30840);
and U38835 (N_38835,N_33307,N_31548);
nand U38836 (N_38836,N_30812,N_32473);
nor U38837 (N_38837,N_34298,N_32416);
and U38838 (N_38838,N_33833,N_31499);
or U38839 (N_38839,N_34823,N_31510);
nor U38840 (N_38840,N_32657,N_32421);
nand U38841 (N_38841,N_31139,N_32672);
nor U38842 (N_38842,N_30936,N_33755);
nor U38843 (N_38843,N_31371,N_33036);
xnor U38844 (N_38844,N_30934,N_32544);
nor U38845 (N_38845,N_30552,N_31858);
xnor U38846 (N_38846,N_34367,N_31137);
and U38847 (N_38847,N_30902,N_30768);
xnor U38848 (N_38848,N_34520,N_33874);
or U38849 (N_38849,N_32287,N_33526);
xnor U38850 (N_38850,N_34235,N_33536);
and U38851 (N_38851,N_33020,N_34865);
nand U38852 (N_38852,N_32944,N_30380);
nand U38853 (N_38853,N_32202,N_33025);
and U38854 (N_38854,N_30419,N_30603);
and U38855 (N_38855,N_34856,N_34026);
nand U38856 (N_38856,N_30967,N_30736);
nand U38857 (N_38857,N_31054,N_30121);
nor U38858 (N_38858,N_34603,N_32258);
nand U38859 (N_38859,N_30681,N_33350);
xnor U38860 (N_38860,N_34003,N_31841);
nand U38861 (N_38861,N_34481,N_32022);
nand U38862 (N_38862,N_31801,N_32466);
or U38863 (N_38863,N_34060,N_32852);
xor U38864 (N_38864,N_33179,N_30829);
and U38865 (N_38865,N_32424,N_30568);
or U38866 (N_38866,N_31322,N_33276);
and U38867 (N_38867,N_33221,N_30140);
nor U38868 (N_38868,N_34194,N_33735);
xor U38869 (N_38869,N_33937,N_33321);
and U38870 (N_38870,N_30981,N_32604);
nor U38871 (N_38871,N_34116,N_33003);
nor U38872 (N_38872,N_30773,N_31538);
nor U38873 (N_38873,N_32649,N_31357);
nand U38874 (N_38874,N_31954,N_33627);
and U38875 (N_38875,N_33107,N_32093);
nand U38876 (N_38876,N_30208,N_31976);
nor U38877 (N_38877,N_34916,N_33264);
and U38878 (N_38878,N_30573,N_33271);
or U38879 (N_38879,N_34317,N_34936);
xor U38880 (N_38880,N_33639,N_33432);
or U38881 (N_38881,N_32874,N_32924);
xor U38882 (N_38882,N_31041,N_32700);
or U38883 (N_38883,N_32453,N_32182);
nor U38884 (N_38884,N_31152,N_30775);
or U38885 (N_38885,N_30921,N_31066);
or U38886 (N_38886,N_31963,N_30081);
nor U38887 (N_38887,N_31658,N_32534);
nor U38888 (N_38888,N_33628,N_34525);
nand U38889 (N_38889,N_30498,N_30082);
nand U38890 (N_38890,N_34330,N_32757);
and U38891 (N_38891,N_31287,N_34633);
or U38892 (N_38892,N_30170,N_31449);
nand U38893 (N_38893,N_33981,N_34166);
nand U38894 (N_38894,N_32801,N_32438);
or U38895 (N_38895,N_31498,N_33177);
nor U38896 (N_38896,N_34329,N_33375);
or U38897 (N_38897,N_34016,N_32485);
nand U38898 (N_38898,N_31659,N_34355);
and U38899 (N_38899,N_34271,N_31616);
xnor U38900 (N_38900,N_32330,N_34796);
nand U38901 (N_38901,N_32959,N_30898);
nand U38902 (N_38902,N_33539,N_32999);
and U38903 (N_38903,N_33128,N_33846);
nand U38904 (N_38904,N_30904,N_32239);
xnor U38905 (N_38905,N_32572,N_34751);
xnor U38906 (N_38906,N_34294,N_31443);
or U38907 (N_38907,N_31750,N_31303);
and U38908 (N_38908,N_32082,N_30318);
or U38909 (N_38909,N_31442,N_34935);
and U38910 (N_38910,N_31263,N_31179);
nor U38911 (N_38911,N_33515,N_32769);
or U38912 (N_38912,N_34410,N_31874);
or U38913 (N_38913,N_30570,N_34962);
and U38914 (N_38914,N_34411,N_32809);
nand U38915 (N_38915,N_32890,N_32234);
nor U38916 (N_38916,N_33728,N_34841);
nand U38917 (N_38917,N_31123,N_33039);
or U38918 (N_38918,N_32675,N_34731);
nand U38919 (N_38919,N_30250,N_32392);
xor U38920 (N_38920,N_30079,N_34377);
nor U38921 (N_38921,N_31060,N_30130);
xor U38922 (N_38922,N_30131,N_31108);
xor U38923 (N_38923,N_31811,N_33100);
xor U38924 (N_38924,N_31030,N_31805);
nor U38925 (N_38925,N_33203,N_31760);
and U38926 (N_38926,N_30033,N_34704);
or U38927 (N_38927,N_33235,N_32663);
nand U38928 (N_38928,N_30882,N_33242);
and U38929 (N_38929,N_32902,N_33403);
and U38930 (N_38930,N_32345,N_32544);
nor U38931 (N_38931,N_34913,N_31895);
or U38932 (N_38932,N_32913,N_33033);
nor U38933 (N_38933,N_33139,N_31992);
xor U38934 (N_38934,N_31829,N_30343);
xor U38935 (N_38935,N_31068,N_32125);
nand U38936 (N_38936,N_34046,N_31497);
xnor U38937 (N_38937,N_33313,N_30590);
nand U38938 (N_38938,N_30289,N_34554);
nand U38939 (N_38939,N_30307,N_33230);
and U38940 (N_38940,N_31921,N_31054);
xor U38941 (N_38941,N_33421,N_33613);
nand U38942 (N_38942,N_30244,N_30971);
or U38943 (N_38943,N_32429,N_33187);
xor U38944 (N_38944,N_31767,N_34198);
or U38945 (N_38945,N_30899,N_30892);
or U38946 (N_38946,N_31790,N_31059);
and U38947 (N_38947,N_34673,N_32157);
xor U38948 (N_38948,N_34656,N_32140);
and U38949 (N_38949,N_30721,N_31051);
xnor U38950 (N_38950,N_33901,N_34930);
or U38951 (N_38951,N_33779,N_33817);
nand U38952 (N_38952,N_30291,N_32156);
or U38953 (N_38953,N_33623,N_30420);
or U38954 (N_38954,N_31385,N_31806);
and U38955 (N_38955,N_34445,N_33059);
and U38956 (N_38956,N_30204,N_32971);
nor U38957 (N_38957,N_34336,N_33376);
nor U38958 (N_38958,N_33244,N_30450);
xor U38959 (N_38959,N_34070,N_33338);
and U38960 (N_38960,N_34628,N_30802);
xor U38961 (N_38961,N_32432,N_34843);
xnor U38962 (N_38962,N_34978,N_34226);
and U38963 (N_38963,N_30521,N_32541);
nand U38964 (N_38964,N_34744,N_31676);
xor U38965 (N_38965,N_31401,N_33586);
or U38966 (N_38966,N_33397,N_34245);
nor U38967 (N_38967,N_33412,N_30881);
nand U38968 (N_38968,N_32915,N_30303);
xor U38969 (N_38969,N_34081,N_34210);
xnor U38970 (N_38970,N_30758,N_34660);
and U38971 (N_38971,N_30917,N_31534);
and U38972 (N_38972,N_33654,N_33247);
or U38973 (N_38973,N_34062,N_30152);
nand U38974 (N_38974,N_30726,N_31344);
or U38975 (N_38975,N_34556,N_31344);
xor U38976 (N_38976,N_30358,N_32050);
xnor U38977 (N_38977,N_30418,N_34930);
nor U38978 (N_38978,N_33058,N_32659);
and U38979 (N_38979,N_31917,N_30889);
nand U38980 (N_38980,N_34477,N_31012);
nor U38981 (N_38981,N_31108,N_32848);
and U38982 (N_38982,N_31483,N_34537);
xor U38983 (N_38983,N_31691,N_34218);
xnor U38984 (N_38984,N_34162,N_30193);
nor U38985 (N_38985,N_30208,N_30528);
xnor U38986 (N_38986,N_32786,N_32693);
nor U38987 (N_38987,N_31890,N_33507);
or U38988 (N_38988,N_32885,N_34190);
and U38989 (N_38989,N_33893,N_31888);
and U38990 (N_38990,N_34021,N_34315);
nor U38991 (N_38991,N_31435,N_33056);
and U38992 (N_38992,N_33241,N_34957);
nand U38993 (N_38993,N_30250,N_32943);
or U38994 (N_38994,N_30131,N_33919);
or U38995 (N_38995,N_34893,N_32275);
nor U38996 (N_38996,N_33588,N_34863);
and U38997 (N_38997,N_33961,N_34104);
or U38998 (N_38998,N_34628,N_32944);
and U38999 (N_38999,N_34943,N_33601);
nand U39000 (N_39000,N_30525,N_32718);
and U39001 (N_39001,N_31493,N_31443);
nor U39002 (N_39002,N_30298,N_31348);
nor U39003 (N_39003,N_30711,N_33661);
nor U39004 (N_39004,N_32603,N_33519);
or U39005 (N_39005,N_32122,N_30660);
nor U39006 (N_39006,N_31203,N_34087);
xor U39007 (N_39007,N_33194,N_31277);
or U39008 (N_39008,N_31025,N_31845);
or U39009 (N_39009,N_31080,N_30950);
nor U39010 (N_39010,N_32695,N_31124);
or U39011 (N_39011,N_34065,N_30633);
nor U39012 (N_39012,N_31368,N_33370);
or U39013 (N_39013,N_31254,N_30053);
and U39014 (N_39014,N_32157,N_30250);
nand U39015 (N_39015,N_32304,N_33333);
nand U39016 (N_39016,N_34061,N_34258);
nor U39017 (N_39017,N_31561,N_30780);
or U39018 (N_39018,N_32460,N_30092);
nor U39019 (N_39019,N_34796,N_33928);
nor U39020 (N_39020,N_30903,N_34275);
nor U39021 (N_39021,N_32891,N_34489);
xor U39022 (N_39022,N_30976,N_31414);
and U39023 (N_39023,N_34123,N_32025);
or U39024 (N_39024,N_31067,N_33564);
or U39025 (N_39025,N_33948,N_34974);
nand U39026 (N_39026,N_32896,N_30715);
nand U39027 (N_39027,N_34850,N_32038);
nor U39028 (N_39028,N_30143,N_32591);
nand U39029 (N_39029,N_30403,N_32079);
and U39030 (N_39030,N_30407,N_30273);
nor U39031 (N_39031,N_32772,N_31555);
xor U39032 (N_39032,N_31428,N_34115);
and U39033 (N_39033,N_30443,N_30911);
nand U39034 (N_39034,N_32322,N_33037);
or U39035 (N_39035,N_34602,N_30014);
and U39036 (N_39036,N_30708,N_31154);
xor U39037 (N_39037,N_30937,N_32323);
or U39038 (N_39038,N_32326,N_32456);
and U39039 (N_39039,N_34088,N_30348);
xnor U39040 (N_39040,N_34477,N_31489);
nand U39041 (N_39041,N_33105,N_33745);
and U39042 (N_39042,N_33136,N_31002);
nand U39043 (N_39043,N_34583,N_33958);
and U39044 (N_39044,N_32303,N_32665);
and U39045 (N_39045,N_33918,N_30277);
nand U39046 (N_39046,N_31643,N_30725);
or U39047 (N_39047,N_33347,N_33639);
or U39048 (N_39048,N_33381,N_34876);
xnor U39049 (N_39049,N_33830,N_33119);
and U39050 (N_39050,N_34471,N_33619);
xor U39051 (N_39051,N_34873,N_33739);
nand U39052 (N_39052,N_32154,N_33817);
or U39053 (N_39053,N_30447,N_30150);
xor U39054 (N_39054,N_31423,N_32340);
or U39055 (N_39055,N_33078,N_30639);
nor U39056 (N_39056,N_31716,N_34127);
and U39057 (N_39057,N_31650,N_31974);
or U39058 (N_39058,N_34288,N_32935);
xnor U39059 (N_39059,N_33425,N_31605);
nand U39060 (N_39060,N_30559,N_33038);
nor U39061 (N_39061,N_30319,N_31339);
and U39062 (N_39062,N_34644,N_34173);
nand U39063 (N_39063,N_32338,N_30857);
and U39064 (N_39064,N_34240,N_31440);
nand U39065 (N_39065,N_31497,N_30832);
and U39066 (N_39066,N_30867,N_30609);
nor U39067 (N_39067,N_32609,N_33395);
xnor U39068 (N_39068,N_33268,N_33930);
xnor U39069 (N_39069,N_32703,N_32527);
nor U39070 (N_39070,N_34070,N_30030);
xnor U39071 (N_39071,N_34326,N_32380);
nor U39072 (N_39072,N_32822,N_33236);
nor U39073 (N_39073,N_32364,N_30099);
nor U39074 (N_39074,N_32355,N_31001);
nor U39075 (N_39075,N_31579,N_31091);
nor U39076 (N_39076,N_31845,N_32344);
and U39077 (N_39077,N_30169,N_32203);
nor U39078 (N_39078,N_32486,N_30796);
or U39079 (N_39079,N_33928,N_34407);
nand U39080 (N_39080,N_32556,N_30309);
nor U39081 (N_39081,N_34032,N_31542);
nor U39082 (N_39082,N_34001,N_34315);
or U39083 (N_39083,N_34785,N_32229);
xnor U39084 (N_39084,N_32597,N_30691);
nand U39085 (N_39085,N_30891,N_30900);
or U39086 (N_39086,N_33376,N_31328);
xnor U39087 (N_39087,N_32933,N_31093);
nor U39088 (N_39088,N_31715,N_32281);
or U39089 (N_39089,N_34745,N_31418);
nand U39090 (N_39090,N_33831,N_33584);
and U39091 (N_39091,N_33767,N_34601);
or U39092 (N_39092,N_33884,N_31681);
nor U39093 (N_39093,N_33749,N_30564);
and U39094 (N_39094,N_30927,N_34373);
nor U39095 (N_39095,N_33229,N_30806);
and U39096 (N_39096,N_33883,N_30116);
xnor U39097 (N_39097,N_31381,N_32276);
or U39098 (N_39098,N_34309,N_31112);
xnor U39099 (N_39099,N_30840,N_33397);
or U39100 (N_39100,N_33977,N_31913);
xor U39101 (N_39101,N_30296,N_34234);
nor U39102 (N_39102,N_34127,N_33744);
xnor U39103 (N_39103,N_32303,N_33982);
and U39104 (N_39104,N_31403,N_32616);
xnor U39105 (N_39105,N_30247,N_31422);
nor U39106 (N_39106,N_34374,N_34344);
xor U39107 (N_39107,N_30195,N_30433);
or U39108 (N_39108,N_34324,N_32478);
and U39109 (N_39109,N_30589,N_32114);
nand U39110 (N_39110,N_31957,N_30999);
nor U39111 (N_39111,N_32684,N_30832);
xor U39112 (N_39112,N_31326,N_32640);
nor U39113 (N_39113,N_32456,N_34751);
and U39114 (N_39114,N_33159,N_32516);
or U39115 (N_39115,N_34106,N_32761);
and U39116 (N_39116,N_33302,N_31726);
nand U39117 (N_39117,N_30317,N_34384);
nand U39118 (N_39118,N_34984,N_32119);
nor U39119 (N_39119,N_30126,N_32386);
nor U39120 (N_39120,N_33209,N_32341);
and U39121 (N_39121,N_34982,N_32288);
and U39122 (N_39122,N_31757,N_32166);
nor U39123 (N_39123,N_32113,N_33102);
and U39124 (N_39124,N_34576,N_31851);
nand U39125 (N_39125,N_31299,N_31285);
nor U39126 (N_39126,N_33744,N_33067);
nand U39127 (N_39127,N_34210,N_30094);
nand U39128 (N_39128,N_30277,N_32557);
xor U39129 (N_39129,N_33786,N_31375);
and U39130 (N_39130,N_34255,N_30992);
or U39131 (N_39131,N_32343,N_32251);
and U39132 (N_39132,N_33756,N_32601);
xor U39133 (N_39133,N_31228,N_32909);
nand U39134 (N_39134,N_30784,N_33752);
or U39135 (N_39135,N_34672,N_31092);
xor U39136 (N_39136,N_32793,N_33723);
nand U39137 (N_39137,N_31752,N_34558);
or U39138 (N_39138,N_32627,N_34937);
nand U39139 (N_39139,N_33973,N_30689);
and U39140 (N_39140,N_30507,N_30427);
or U39141 (N_39141,N_33725,N_33514);
and U39142 (N_39142,N_34312,N_30704);
nand U39143 (N_39143,N_33952,N_33752);
and U39144 (N_39144,N_33185,N_34662);
or U39145 (N_39145,N_33491,N_34346);
xor U39146 (N_39146,N_32561,N_32711);
nand U39147 (N_39147,N_30778,N_30675);
and U39148 (N_39148,N_30143,N_32650);
nand U39149 (N_39149,N_32692,N_34505);
nor U39150 (N_39150,N_34383,N_32437);
and U39151 (N_39151,N_33824,N_32584);
or U39152 (N_39152,N_34528,N_32416);
and U39153 (N_39153,N_32761,N_30002);
nor U39154 (N_39154,N_34353,N_34783);
xor U39155 (N_39155,N_33224,N_31679);
and U39156 (N_39156,N_30314,N_30319);
xnor U39157 (N_39157,N_30992,N_30069);
nand U39158 (N_39158,N_34958,N_31011);
and U39159 (N_39159,N_34280,N_31666);
or U39160 (N_39160,N_34092,N_31539);
or U39161 (N_39161,N_33333,N_32880);
or U39162 (N_39162,N_34595,N_30891);
or U39163 (N_39163,N_33158,N_34253);
nor U39164 (N_39164,N_32874,N_34446);
nand U39165 (N_39165,N_31419,N_32134);
and U39166 (N_39166,N_32359,N_32168);
and U39167 (N_39167,N_30298,N_33170);
xnor U39168 (N_39168,N_30249,N_34843);
and U39169 (N_39169,N_33268,N_32968);
and U39170 (N_39170,N_33973,N_31588);
nand U39171 (N_39171,N_30440,N_32350);
and U39172 (N_39172,N_34363,N_33942);
nand U39173 (N_39173,N_30404,N_30610);
and U39174 (N_39174,N_34925,N_33608);
xnor U39175 (N_39175,N_34055,N_34823);
or U39176 (N_39176,N_32330,N_31573);
xor U39177 (N_39177,N_34721,N_33274);
and U39178 (N_39178,N_32004,N_34648);
nand U39179 (N_39179,N_33953,N_31505);
and U39180 (N_39180,N_31521,N_33474);
and U39181 (N_39181,N_31193,N_30015);
nand U39182 (N_39182,N_32799,N_34786);
xnor U39183 (N_39183,N_32709,N_31142);
or U39184 (N_39184,N_33845,N_34314);
and U39185 (N_39185,N_34624,N_30249);
nor U39186 (N_39186,N_30577,N_32921);
nor U39187 (N_39187,N_32300,N_33426);
and U39188 (N_39188,N_31029,N_33810);
nand U39189 (N_39189,N_31133,N_33436);
or U39190 (N_39190,N_31515,N_34706);
or U39191 (N_39191,N_31355,N_31680);
or U39192 (N_39192,N_30981,N_33260);
and U39193 (N_39193,N_34662,N_30901);
or U39194 (N_39194,N_30229,N_32330);
nor U39195 (N_39195,N_34806,N_32211);
or U39196 (N_39196,N_34457,N_32384);
xnor U39197 (N_39197,N_33016,N_32813);
xor U39198 (N_39198,N_30750,N_30220);
nor U39199 (N_39199,N_33189,N_34561);
or U39200 (N_39200,N_34440,N_33866);
and U39201 (N_39201,N_33088,N_31617);
nand U39202 (N_39202,N_33846,N_34871);
xor U39203 (N_39203,N_31479,N_31348);
and U39204 (N_39204,N_34620,N_34897);
and U39205 (N_39205,N_32285,N_30388);
xnor U39206 (N_39206,N_30757,N_34276);
xor U39207 (N_39207,N_30292,N_30676);
xnor U39208 (N_39208,N_32738,N_31711);
and U39209 (N_39209,N_33912,N_32548);
and U39210 (N_39210,N_33303,N_32938);
nand U39211 (N_39211,N_33245,N_32534);
xnor U39212 (N_39212,N_30179,N_30377);
and U39213 (N_39213,N_31130,N_33530);
nand U39214 (N_39214,N_30004,N_33215);
nand U39215 (N_39215,N_32723,N_33009);
nand U39216 (N_39216,N_31805,N_33272);
nand U39217 (N_39217,N_32544,N_34514);
or U39218 (N_39218,N_32243,N_31376);
nor U39219 (N_39219,N_34688,N_34532);
nor U39220 (N_39220,N_30113,N_30670);
or U39221 (N_39221,N_33344,N_34696);
nor U39222 (N_39222,N_34017,N_30027);
nor U39223 (N_39223,N_32819,N_34884);
or U39224 (N_39224,N_34416,N_30158);
xnor U39225 (N_39225,N_32391,N_33640);
nor U39226 (N_39226,N_32498,N_33166);
and U39227 (N_39227,N_32028,N_32608);
nor U39228 (N_39228,N_31303,N_34327);
nand U39229 (N_39229,N_31776,N_33569);
nor U39230 (N_39230,N_30125,N_30731);
or U39231 (N_39231,N_32980,N_31565);
and U39232 (N_39232,N_34509,N_30750);
and U39233 (N_39233,N_32616,N_31195);
or U39234 (N_39234,N_32914,N_30637);
and U39235 (N_39235,N_30506,N_33396);
and U39236 (N_39236,N_33745,N_33246);
xnor U39237 (N_39237,N_31917,N_33664);
xor U39238 (N_39238,N_33566,N_34265);
and U39239 (N_39239,N_30455,N_32584);
and U39240 (N_39240,N_30982,N_33728);
nor U39241 (N_39241,N_30730,N_33278);
nand U39242 (N_39242,N_30266,N_33785);
or U39243 (N_39243,N_31434,N_33887);
nand U39244 (N_39244,N_31944,N_32434);
nor U39245 (N_39245,N_32863,N_30958);
xor U39246 (N_39246,N_34376,N_32959);
and U39247 (N_39247,N_30051,N_33477);
nor U39248 (N_39248,N_34481,N_31096);
and U39249 (N_39249,N_31704,N_31034);
nor U39250 (N_39250,N_30410,N_33164);
or U39251 (N_39251,N_31048,N_34241);
or U39252 (N_39252,N_32499,N_32054);
or U39253 (N_39253,N_30712,N_31514);
and U39254 (N_39254,N_31383,N_34541);
or U39255 (N_39255,N_31915,N_30673);
xnor U39256 (N_39256,N_30569,N_34732);
nand U39257 (N_39257,N_34826,N_31787);
xor U39258 (N_39258,N_31514,N_32395);
nand U39259 (N_39259,N_32512,N_34096);
nor U39260 (N_39260,N_33298,N_31774);
nand U39261 (N_39261,N_30514,N_32958);
and U39262 (N_39262,N_30575,N_31299);
nand U39263 (N_39263,N_31636,N_31362);
xor U39264 (N_39264,N_32992,N_34882);
nand U39265 (N_39265,N_33542,N_32673);
and U39266 (N_39266,N_33572,N_31319);
and U39267 (N_39267,N_34466,N_32713);
nor U39268 (N_39268,N_33245,N_32338);
or U39269 (N_39269,N_30596,N_31762);
nand U39270 (N_39270,N_32931,N_32231);
and U39271 (N_39271,N_31365,N_32682);
and U39272 (N_39272,N_32862,N_34667);
nand U39273 (N_39273,N_33061,N_34852);
and U39274 (N_39274,N_32549,N_34827);
nor U39275 (N_39275,N_34966,N_31987);
and U39276 (N_39276,N_30293,N_30361);
nand U39277 (N_39277,N_32474,N_30278);
and U39278 (N_39278,N_31481,N_30345);
and U39279 (N_39279,N_31027,N_34094);
xor U39280 (N_39280,N_30387,N_31097);
xnor U39281 (N_39281,N_31063,N_34308);
nor U39282 (N_39282,N_31941,N_34500);
nor U39283 (N_39283,N_33224,N_34457);
nand U39284 (N_39284,N_31304,N_34717);
nand U39285 (N_39285,N_33769,N_34653);
or U39286 (N_39286,N_34310,N_30130);
xnor U39287 (N_39287,N_31364,N_33461);
nand U39288 (N_39288,N_31452,N_30179);
or U39289 (N_39289,N_33939,N_32226);
and U39290 (N_39290,N_33048,N_34235);
and U39291 (N_39291,N_33043,N_33422);
and U39292 (N_39292,N_34469,N_30596);
nor U39293 (N_39293,N_31235,N_33490);
or U39294 (N_39294,N_31293,N_34374);
or U39295 (N_39295,N_34675,N_30592);
or U39296 (N_39296,N_31068,N_33244);
or U39297 (N_39297,N_32931,N_33443);
nand U39298 (N_39298,N_30493,N_31818);
xnor U39299 (N_39299,N_33868,N_34175);
or U39300 (N_39300,N_32951,N_30246);
or U39301 (N_39301,N_30274,N_32604);
or U39302 (N_39302,N_31083,N_34275);
nor U39303 (N_39303,N_31264,N_33375);
or U39304 (N_39304,N_34882,N_31040);
and U39305 (N_39305,N_30779,N_33964);
or U39306 (N_39306,N_31787,N_31035);
or U39307 (N_39307,N_30578,N_34646);
nor U39308 (N_39308,N_30187,N_33299);
and U39309 (N_39309,N_32923,N_34755);
nor U39310 (N_39310,N_34235,N_32072);
nand U39311 (N_39311,N_30505,N_33705);
or U39312 (N_39312,N_31945,N_31609);
nor U39313 (N_39313,N_32269,N_34377);
nand U39314 (N_39314,N_32874,N_30531);
xor U39315 (N_39315,N_30595,N_33503);
xor U39316 (N_39316,N_33038,N_30379);
xor U39317 (N_39317,N_32933,N_33233);
or U39318 (N_39318,N_30730,N_31999);
xor U39319 (N_39319,N_31276,N_30028);
or U39320 (N_39320,N_32868,N_34770);
and U39321 (N_39321,N_34797,N_30000);
nor U39322 (N_39322,N_33836,N_34630);
nand U39323 (N_39323,N_31602,N_30506);
and U39324 (N_39324,N_34726,N_34568);
or U39325 (N_39325,N_31381,N_34692);
nand U39326 (N_39326,N_34780,N_31827);
and U39327 (N_39327,N_31746,N_33874);
nor U39328 (N_39328,N_32372,N_32616);
nor U39329 (N_39329,N_30837,N_31070);
and U39330 (N_39330,N_32169,N_30888);
xnor U39331 (N_39331,N_33132,N_34340);
or U39332 (N_39332,N_34199,N_31932);
nor U39333 (N_39333,N_31010,N_31172);
and U39334 (N_39334,N_31029,N_32055);
nand U39335 (N_39335,N_33319,N_34969);
and U39336 (N_39336,N_32097,N_33495);
and U39337 (N_39337,N_30549,N_31210);
nand U39338 (N_39338,N_34039,N_31853);
and U39339 (N_39339,N_34227,N_33456);
or U39340 (N_39340,N_33277,N_31470);
and U39341 (N_39341,N_33038,N_33324);
or U39342 (N_39342,N_32132,N_33269);
and U39343 (N_39343,N_32895,N_33457);
nand U39344 (N_39344,N_33716,N_31656);
xnor U39345 (N_39345,N_33028,N_34041);
nand U39346 (N_39346,N_30349,N_34414);
and U39347 (N_39347,N_32770,N_32040);
or U39348 (N_39348,N_32316,N_32114);
and U39349 (N_39349,N_32524,N_32827);
nor U39350 (N_39350,N_34743,N_31353);
nor U39351 (N_39351,N_32491,N_33519);
nor U39352 (N_39352,N_30276,N_31942);
nor U39353 (N_39353,N_30408,N_33396);
or U39354 (N_39354,N_30866,N_31870);
and U39355 (N_39355,N_33729,N_31466);
nor U39356 (N_39356,N_30800,N_34281);
xnor U39357 (N_39357,N_33791,N_32313);
or U39358 (N_39358,N_33640,N_30245);
or U39359 (N_39359,N_31401,N_32489);
nand U39360 (N_39360,N_33549,N_33249);
nor U39361 (N_39361,N_33585,N_30550);
or U39362 (N_39362,N_30754,N_31026);
xnor U39363 (N_39363,N_30767,N_31832);
or U39364 (N_39364,N_32128,N_34566);
nand U39365 (N_39365,N_30918,N_33124);
xor U39366 (N_39366,N_34338,N_30291);
and U39367 (N_39367,N_31503,N_34578);
and U39368 (N_39368,N_31666,N_31258);
and U39369 (N_39369,N_31533,N_33861);
nand U39370 (N_39370,N_32378,N_30876);
nor U39371 (N_39371,N_30958,N_30485);
or U39372 (N_39372,N_31339,N_33339);
nand U39373 (N_39373,N_34836,N_33503);
xor U39374 (N_39374,N_31198,N_31140);
nor U39375 (N_39375,N_31171,N_34063);
nor U39376 (N_39376,N_30607,N_31003);
xnor U39377 (N_39377,N_31956,N_33507);
nand U39378 (N_39378,N_32583,N_34905);
nor U39379 (N_39379,N_34376,N_34741);
xor U39380 (N_39380,N_30772,N_33523);
nand U39381 (N_39381,N_30581,N_33424);
and U39382 (N_39382,N_33718,N_34105);
and U39383 (N_39383,N_33580,N_33073);
or U39384 (N_39384,N_32527,N_32401);
xnor U39385 (N_39385,N_32677,N_32315);
nor U39386 (N_39386,N_34208,N_30834);
nand U39387 (N_39387,N_30152,N_33024);
xor U39388 (N_39388,N_31577,N_31691);
and U39389 (N_39389,N_34997,N_31725);
and U39390 (N_39390,N_32651,N_31447);
xnor U39391 (N_39391,N_34936,N_31936);
xnor U39392 (N_39392,N_32264,N_31296);
nand U39393 (N_39393,N_32877,N_33343);
nand U39394 (N_39394,N_33478,N_31486);
and U39395 (N_39395,N_34856,N_31241);
nor U39396 (N_39396,N_31841,N_34092);
and U39397 (N_39397,N_30071,N_34863);
nor U39398 (N_39398,N_34504,N_33104);
nor U39399 (N_39399,N_30277,N_30146);
and U39400 (N_39400,N_32709,N_33445);
or U39401 (N_39401,N_33406,N_31867);
nor U39402 (N_39402,N_33079,N_33528);
or U39403 (N_39403,N_30170,N_34163);
or U39404 (N_39404,N_32834,N_34440);
and U39405 (N_39405,N_32152,N_31732);
and U39406 (N_39406,N_33223,N_30989);
nor U39407 (N_39407,N_30655,N_34696);
nand U39408 (N_39408,N_34475,N_30175);
nand U39409 (N_39409,N_31300,N_34243);
or U39410 (N_39410,N_31346,N_31650);
and U39411 (N_39411,N_34100,N_31724);
and U39412 (N_39412,N_32626,N_32273);
or U39413 (N_39413,N_33882,N_34644);
or U39414 (N_39414,N_32107,N_31392);
nand U39415 (N_39415,N_32969,N_31424);
xor U39416 (N_39416,N_33730,N_30152);
xor U39417 (N_39417,N_31952,N_34516);
nand U39418 (N_39418,N_33845,N_33279);
nor U39419 (N_39419,N_32670,N_32104);
nand U39420 (N_39420,N_33925,N_31915);
nor U39421 (N_39421,N_30848,N_32291);
or U39422 (N_39422,N_31129,N_32225);
xor U39423 (N_39423,N_30736,N_34948);
nor U39424 (N_39424,N_34825,N_32255);
and U39425 (N_39425,N_32193,N_33627);
nor U39426 (N_39426,N_33732,N_32989);
nor U39427 (N_39427,N_30503,N_34688);
xor U39428 (N_39428,N_31835,N_30149);
xnor U39429 (N_39429,N_34232,N_32754);
or U39430 (N_39430,N_30689,N_32693);
or U39431 (N_39431,N_32179,N_31514);
nor U39432 (N_39432,N_31533,N_31455);
nor U39433 (N_39433,N_30557,N_32546);
nor U39434 (N_39434,N_32850,N_31005);
xor U39435 (N_39435,N_30495,N_31718);
nand U39436 (N_39436,N_32639,N_31284);
xor U39437 (N_39437,N_32845,N_31099);
and U39438 (N_39438,N_31154,N_34493);
xnor U39439 (N_39439,N_31781,N_32159);
and U39440 (N_39440,N_32905,N_33163);
and U39441 (N_39441,N_34632,N_31328);
nand U39442 (N_39442,N_34397,N_33584);
xnor U39443 (N_39443,N_30370,N_30827);
or U39444 (N_39444,N_34066,N_32922);
or U39445 (N_39445,N_30238,N_30664);
and U39446 (N_39446,N_32416,N_32803);
nor U39447 (N_39447,N_34822,N_33000);
or U39448 (N_39448,N_32873,N_31020);
xnor U39449 (N_39449,N_33421,N_33958);
nand U39450 (N_39450,N_31098,N_31635);
nor U39451 (N_39451,N_32010,N_31436);
xnor U39452 (N_39452,N_33493,N_32946);
or U39453 (N_39453,N_31275,N_34073);
nand U39454 (N_39454,N_34583,N_33252);
nand U39455 (N_39455,N_34013,N_33478);
or U39456 (N_39456,N_32567,N_33543);
nand U39457 (N_39457,N_30664,N_33215);
nor U39458 (N_39458,N_30408,N_33710);
or U39459 (N_39459,N_34003,N_30989);
xor U39460 (N_39460,N_30175,N_33279);
nand U39461 (N_39461,N_33414,N_31685);
and U39462 (N_39462,N_31443,N_34882);
nor U39463 (N_39463,N_30940,N_31790);
nand U39464 (N_39464,N_32657,N_33464);
and U39465 (N_39465,N_33744,N_32311);
nor U39466 (N_39466,N_32285,N_31452);
nor U39467 (N_39467,N_31977,N_32500);
nand U39468 (N_39468,N_30205,N_33744);
xor U39469 (N_39469,N_32148,N_34091);
nor U39470 (N_39470,N_32165,N_30367);
or U39471 (N_39471,N_32507,N_33869);
and U39472 (N_39472,N_31355,N_33682);
or U39473 (N_39473,N_32399,N_32012);
xnor U39474 (N_39474,N_33593,N_33862);
xnor U39475 (N_39475,N_30550,N_31936);
xnor U39476 (N_39476,N_30772,N_31757);
xor U39477 (N_39477,N_32337,N_32006);
nor U39478 (N_39478,N_32337,N_34998);
and U39479 (N_39479,N_30224,N_33866);
or U39480 (N_39480,N_30676,N_30820);
nand U39481 (N_39481,N_32242,N_34825);
or U39482 (N_39482,N_32583,N_31875);
nand U39483 (N_39483,N_31840,N_30169);
and U39484 (N_39484,N_30036,N_33689);
nand U39485 (N_39485,N_32137,N_33014);
and U39486 (N_39486,N_34932,N_31090);
and U39487 (N_39487,N_34982,N_32630);
or U39488 (N_39488,N_32354,N_31004);
xor U39489 (N_39489,N_33808,N_30318);
nand U39490 (N_39490,N_31826,N_33494);
and U39491 (N_39491,N_33286,N_31902);
nor U39492 (N_39492,N_32348,N_31087);
xor U39493 (N_39493,N_33952,N_31456);
nand U39494 (N_39494,N_32124,N_32652);
or U39495 (N_39495,N_32254,N_30305);
nand U39496 (N_39496,N_32611,N_33557);
nand U39497 (N_39497,N_34663,N_32867);
and U39498 (N_39498,N_31131,N_33099);
xnor U39499 (N_39499,N_32946,N_31982);
nor U39500 (N_39500,N_34987,N_30423);
and U39501 (N_39501,N_30121,N_34679);
xnor U39502 (N_39502,N_32632,N_31686);
nand U39503 (N_39503,N_31737,N_31710);
nand U39504 (N_39504,N_32092,N_34631);
xnor U39505 (N_39505,N_32069,N_33677);
nor U39506 (N_39506,N_31802,N_33232);
and U39507 (N_39507,N_30206,N_30924);
nand U39508 (N_39508,N_30648,N_32692);
nor U39509 (N_39509,N_33465,N_34677);
nand U39510 (N_39510,N_32467,N_30736);
nand U39511 (N_39511,N_32542,N_32971);
xor U39512 (N_39512,N_33134,N_34661);
nand U39513 (N_39513,N_30273,N_33288);
or U39514 (N_39514,N_32348,N_33885);
or U39515 (N_39515,N_30989,N_31140);
nor U39516 (N_39516,N_33697,N_30446);
and U39517 (N_39517,N_30287,N_34210);
xnor U39518 (N_39518,N_34930,N_33993);
and U39519 (N_39519,N_32536,N_32799);
and U39520 (N_39520,N_30233,N_30239);
xor U39521 (N_39521,N_32476,N_30835);
nand U39522 (N_39522,N_33395,N_34434);
and U39523 (N_39523,N_30082,N_30463);
nand U39524 (N_39524,N_30769,N_33149);
nand U39525 (N_39525,N_30590,N_30021);
nor U39526 (N_39526,N_30126,N_32635);
nor U39527 (N_39527,N_31318,N_34802);
nor U39528 (N_39528,N_30205,N_34530);
xnor U39529 (N_39529,N_33971,N_31919);
nor U39530 (N_39530,N_31751,N_33257);
xor U39531 (N_39531,N_31662,N_30184);
nand U39532 (N_39532,N_31719,N_34406);
nor U39533 (N_39533,N_32072,N_33614);
or U39534 (N_39534,N_31749,N_31982);
nand U39535 (N_39535,N_34524,N_33428);
nand U39536 (N_39536,N_33151,N_30954);
nand U39537 (N_39537,N_31017,N_30559);
and U39538 (N_39538,N_34611,N_31110);
nor U39539 (N_39539,N_31089,N_33933);
xnor U39540 (N_39540,N_34371,N_32563);
or U39541 (N_39541,N_31060,N_34352);
and U39542 (N_39542,N_32831,N_32496);
nand U39543 (N_39543,N_30394,N_34467);
or U39544 (N_39544,N_34601,N_33564);
or U39545 (N_39545,N_33513,N_30290);
nand U39546 (N_39546,N_34076,N_33892);
nor U39547 (N_39547,N_31708,N_33568);
nor U39548 (N_39548,N_32310,N_34875);
and U39549 (N_39549,N_34999,N_33359);
or U39550 (N_39550,N_31474,N_33643);
or U39551 (N_39551,N_31051,N_31437);
or U39552 (N_39552,N_32310,N_34675);
and U39553 (N_39553,N_34313,N_30008);
or U39554 (N_39554,N_32114,N_33603);
nor U39555 (N_39555,N_31597,N_34430);
xnor U39556 (N_39556,N_33168,N_31322);
and U39557 (N_39557,N_30350,N_31008);
nand U39558 (N_39558,N_34053,N_33459);
nor U39559 (N_39559,N_30334,N_32555);
nor U39560 (N_39560,N_31001,N_31783);
nand U39561 (N_39561,N_30532,N_33585);
nor U39562 (N_39562,N_31546,N_33585);
nand U39563 (N_39563,N_33884,N_30961);
or U39564 (N_39564,N_31528,N_30937);
nor U39565 (N_39565,N_32338,N_33504);
or U39566 (N_39566,N_31629,N_34238);
nor U39567 (N_39567,N_33790,N_32205);
or U39568 (N_39568,N_31480,N_30046);
or U39569 (N_39569,N_34048,N_34680);
and U39570 (N_39570,N_33737,N_31828);
xor U39571 (N_39571,N_30356,N_30803);
and U39572 (N_39572,N_32888,N_33112);
or U39573 (N_39573,N_33130,N_31517);
nor U39574 (N_39574,N_30206,N_34713);
nand U39575 (N_39575,N_33164,N_30796);
nand U39576 (N_39576,N_33101,N_33502);
nor U39577 (N_39577,N_34450,N_32512);
and U39578 (N_39578,N_33749,N_32171);
or U39579 (N_39579,N_30884,N_30150);
xor U39580 (N_39580,N_34188,N_31469);
or U39581 (N_39581,N_31798,N_30837);
xor U39582 (N_39582,N_34691,N_32668);
nand U39583 (N_39583,N_34115,N_32655);
and U39584 (N_39584,N_31191,N_34778);
nor U39585 (N_39585,N_33427,N_31537);
and U39586 (N_39586,N_30285,N_33771);
or U39587 (N_39587,N_33413,N_30983);
xor U39588 (N_39588,N_34407,N_33039);
or U39589 (N_39589,N_33917,N_31210);
and U39590 (N_39590,N_31136,N_31445);
and U39591 (N_39591,N_30629,N_32335);
or U39592 (N_39592,N_30982,N_32038);
xor U39593 (N_39593,N_32026,N_31439);
nand U39594 (N_39594,N_34168,N_34114);
nand U39595 (N_39595,N_32935,N_33683);
xnor U39596 (N_39596,N_33720,N_30054);
xor U39597 (N_39597,N_30029,N_34205);
or U39598 (N_39598,N_33790,N_34573);
nor U39599 (N_39599,N_34837,N_30222);
nand U39600 (N_39600,N_31713,N_32527);
or U39601 (N_39601,N_31004,N_33592);
xnor U39602 (N_39602,N_34816,N_33893);
xnor U39603 (N_39603,N_32762,N_33961);
xor U39604 (N_39604,N_30588,N_33913);
or U39605 (N_39605,N_33812,N_34521);
and U39606 (N_39606,N_30320,N_30090);
and U39607 (N_39607,N_30393,N_31750);
nand U39608 (N_39608,N_34185,N_34513);
or U39609 (N_39609,N_30912,N_30600);
and U39610 (N_39610,N_32286,N_34425);
nand U39611 (N_39611,N_33547,N_33099);
nand U39612 (N_39612,N_30938,N_30247);
or U39613 (N_39613,N_32009,N_33795);
or U39614 (N_39614,N_33113,N_31839);
or U39615 (N_39615,N_31962,N_32901);
nor U39616 (N_39616,N_34257,N_34588);
xnor U39617 (N_39617,N_30193,N_30852);
or U39618 (N_39618,N_32142,N_32132);
xor U39619 (N_39619,N_30211,N_32018);
or U39620 (N_39620,N_30998,N_33317);
nor U39621 (N_39621,N_34149,N_33977);
nor U39622 (N_39622,N_30287,N_30408);
nand U39623 (N_39623,N_32153,N_33081);
xnor U39624 (N_39624,N_30085,N_34043);
xnor U39625 (N_39625,N_34335,N_30642);
or U39626 (N_39626,N_33761,N_34923);
xnor U39627 (N_39627,N_34453,N_34141);
nor U39628 (N_39628,N_30274,N_32699);
nand U39629 (N_39629,N_30069,N_31084);
xnor U39630 (N_39630,N_34742,N_30885);
nor U39631 (N_39631,N_32606,N_33845);
xor U39632 (N_39632,N_34741,N_34136);
or U39633 (N_39633,N_31326,N_34765);
nor U39634 (N_39634,N_34946,N_30825);
nor U39635 (N_39635,N_31204,N_32909);
xor U39636 (N_39636,N_30562,N_32690);
xor U39637 (N_39637,N_34841,N_31364);
or U39638 (N_39638,N_30245,N_31985);
nand U39639 (N_39639,N_34083,N_33000);
and U39640 (N_39640,N_33107,N_30945);
or U39641 (N_39641,N_31215,N_33624);
or U39642 (N_39642,N_32668,N_33306);
or U39643 (N_39643,N_31914,N_34612);
nor U39644 (N_39644,N_34603,N_34082);
and U39645 (N_39645,N_33619,N_34217);
nand U39646 (N_39646,N_32900,N_31049);
and U39647 (N_39647,N_30240,N_30549);
nor U39648 (N_39648,N_32841,N_32091);
xnor U39649 (N_39649,N_34807,N_33315);
or U39650 (N_39650,N_32854,N_33399);
or U39651 (N_39651,N_32590,N_31788);
xor U39652 (N_39652,N_34928,N_33142);
or U39653 (N_39653,N_33485,N_31053);
nor U39654 (N_39654,N_31815,N_31261);
and U39655 (N_39655,N_33303,N_33785);
nand U39656 (N_39656,N_31517,N_31773);
or U39657 (N_39657,N_32294,N_30332);
nand U39658 (N_39658,N_34221,N_33959);
nand U39659 (N_39659,N_33128,N_31250);
or U39660 (N_39660,N_31283,N_30360);
nand U39661 (N_39661,N_33438,N_32183);
xor U39662 (N_39662,N_30397,N_34290);
xor U39663 (N_39663,N_31827,N_31786);
or U39664 (N_39664,N_32057,N_32471);
xor U39665 (N_39665,N_32645,N_31050);
nor U39666 (N_39666,N_34160,N_33115);
and U39667 (N_39667,N_34344,N_31100);
nand U39668 (N_39668,N_34632,N_33424);
xor U39669 (N_39669,N_30955,N_30083);
nor U39670 (N_39670,N_32523,N_30881);
xnor U39671 (N_39671,N_31032,N_30703);
nor U39672 (N_39672,N_31853,N_33784);
nand U39673 (N_39673,N_32161,N_32683);
nor U39674 (N_39674,N_33267,N_33571);
or U39675 (N_39675,N_30753,N_33499);
and U39676 (N_39676,N_31705,N_33300);
nor U39677 (N_39677,N_33060,N_30829);
or U39678 (N_39678,N_34724,N_31445);
nor U39679 (N_39679,N_34388,N_33298);
and U39680 (N_39680,N_32526,N_34955);
xor U39681 (N_39681,N_33513,N_33073);
and U39682 (N_39682,N_32047,N_30716);
nand U39683 (N_39683,N_30540,N_32886);
xnor U39684 (N_39684,N_31022,N_30405);
and U39685 (N_39685,N_31992,N_31647);
or U39686 (N_39686,N_30012,N_33973);
nand U39687 (N_39687,N_34185,N_30922);
nand U39688 (N_39688,N_30418,N_31434);
and U39689 (N_39689,N_33051,N_30551);
or U39690 (N_39690,N_34068,N_34687);
or U39691 (N_39691,N_31373,N_32693);
or U39692 (N_39692,N_34411,N_34762);
or U39693 (N_39693,N_32499,N_31610);
or U39694 (N_39694,N_34236,N_31297);
xor U39695 (N_39695,N_33406,N_33214);
xor U39696 (N_39696,N_31120,N_31863);
xnor U39697 (N_39697,N_34865,N_33769);
xnor U39698 (N_39698,N_34348,N_32902);
or U39699 (N_39699,N_31677,N_34276);
and U39700 (N_39700,N_32538,N_33977);
xnor U39701 (N_39701,N_30416,N_34819);
nor U39702 (N_39702,N_31768,N_31412);
xor U39703 (N_39703,N_32695,N_33606);
xnor U39704 (N_39704,N_30784,N_34945);
nand U39705 (N_39705,N_31159,N_31576);
and U39706 (N_39706,N_31277,N_30733);
nor U39707 (N_39707,N_30274,N_34936);
or U39708 (N_39708,N_33181,N_31135);
nor U39709 (N_39709,N_33349,N_34946);
and U39710 (N_39710,N_30948,N_33956);
xnor U39711 (N_39711,N_30525,N_30423);
nor U39712 (N_39712,N_33710,N_31855);
xor U39713 (N_39713,N_31065,N_30157);
or U39714 (N_39714,N_33006,N_32377);
xnor U39715 (N_39715,N_30411,N_32587);
and U39716 (N_39716,N_31559,N_32174);
xor U39717 (N_39717,N_30478,N_32725);
nand U39718 (N_39718,N_32727,N_33014);
xnor U39719 (N_39719,N_30741,N_32301);
nor U39720 (N_39720,N_31890,N_31789);
nand U39721 (N_39721,N_32682,N_34375);
nor U39722 (N_39722,N_31811,N_31677);
or U39723 (N_39723,N_33911,N_30860);
and U39724 (N_39724,N_31578,N_34485);
nor U39725 (N_39725,N_33744,N_32357);
nand U39726 (N_39726,N_30136,N_32336);
nand U39727 (N_39727,N_33268,N_32590);
nor U39728 (N_39728,N_34040,N_30810);
nor U39729 (N_39729,N_31993,N_31597);
nor U39730 (N_39730,N_33083,N_34885);
nand U39731 (N_39731,N_31815,N_34364);
nor U39732 (N_39732,N_34938,N_30055);
xor U39733 (N_39733,N_31379,N_31897);
or U39734 (N_39734,N_30755,N_31888);
and U39735 (N_39735,N_31282,N_34515);
or U39736 (N_39736,N_33684,N_34999);
xnor U39737 (N_39737,N_31478,N_30541);
nor U39738 (N_39738,N_34474,N_32176);
or U39739 (N_39739,N_32690,N_30276);
nor U39740 (N_39740,N_33737,N_30087);
nor U39741 (N_39741,N_30136,N_32784);
xor U39742 (N_39742,N_33567,N_32569);
xor U39743 (N_39743,N_33734,N_31937);
and U39744 (N_39744,N_30759,N_31061);
xnor U39745 (N_39745,N_30462,N_33842);
nor U39746 (N_39746,N_33042,N_31065);
and U39747 (N_39747,N_32899,N_33815);
or U39748 (N_39748,N_32778,N_32466);
xnor U39749 (N_39749,N_31547,N_34851);
or U39750 (N_39750,N_33833,N_34928);
nor U39751 (N_39751,N_34921,N_33545);
xnor U39752 (N_39752,N_30956,N_34337);
and U39753 (N_39753,N_30670,N_31915);
nor U39754 (N_39754,N_31756,N_32830);
nor U39755 (N_39755,N_33232,N_33927);
and U39756 (N_39756,N_32306,N_33194);
xnor U39757 (N_39757,N_30691,N_34128);
nor U39758 (N_39758,N_30599,N_30954);
or U39759 (N_39759,N_31861,N_30585);
nand U39760 (N_39760,N_33142,N_33617);
or U39761 (N_39761,N_34691,N_33932);
xnor U39762 (N_39762,N_30454,N_34597);
or U39763 (N_39763,N_32521,N_32604);
and U39764 (N_39764,N_30334,N_33137);
xnor U39765 (N_39765,N_33876,N_31964);
xnor U39766 (N_39766,N_34076,N_32259);
nor U39767 (N_39767,N_34304,N_30853);
and U39768 (N_39768,N_34109,N_30189);
nand U39769 (N_39769,N_34757,N_34284);
and U39770 (N_39770,N_33523,N_31644);
nand U39771 (N_39771,N_33736,N_32684);
or U39772 (N_39772,N_33813,N_31205);
xor U39773 (N_39773,N_33388,N_30126);
or U39774 (N_39774,N_31234,N_32495);
and U39775 (N_39775,N_30724,N_34496);
nor U39776 (N_39776,N_34015,N_31358);
nand U39777 (N_39777,N_30879,N_33573);
nor U39778 (N_39778,N_32335,N_31749);
xnor U39779 (N_39779,N_33589,N_32601);
and U39780 (N_39780,N_33002,N_31885);
nand U39781 (N_39781,N_31522,N_32342);
nand U39782 (N_39782,N_32669,N_33688);
or U39783 (N_39783,N_31607,N_31831);
and U39784 (N_39784,N_31040,N_32121);
xor U39785 (N_39785,N_33325,N_33503);
xor U39786 (N_39786,N_34284,N_30593);
nor U39787 (N_39787,N_33169,N_31592);
or U39788 (N_39788,N_33487,N_33969);
and U39789 (N_39789,N_33353,N_31550);
nor U39790 (N_39790,N_34498,N_33120);
or U39791 (N_39791,N_32479,N_31531);
xnor U39792 (N_39792,N_30538,N_34856);
and U39793 (N_39793,N_33236,N_32831);
nand U39794 (N_39794,N_33647,N_30073);
nand U39795 (N_39795,N_34012,N_34072);
nor U39796 (N_39796,N_33446,N_34196);
or U39797 (N_39797,N_30516,N_34376);
nor U39798 (N_39798,N_34420,N_32599);
xor U39799 (N_39799,N_31138,N_31267);
nor U39800 (N_39800,N_30224,N_34690);
and U39801 (N_39801,N_32815,N_33036);
nand U39802 (N_39802,N_30851,N_30784);
nor U39803 (N_39803,N_33758,N_34983);
and U39804 (N_39804,N_30487,N_30109);
nand U39805 (N_39805,N_30496,N_33357);
nor U39806 (N_39806,N_30574,N_30876);
and U39807 (N_39807,N_30852,N_31745);
and U39808 (N_39808,N_34259,N_33341);
nor U39809 (N_39809,N_30939,N_31892);
nor U39810 (N_39810,N_30749,N_34542);
xnor U39811 (N_39811,N_31160,N_33262);
nor U39812 (N_39812,N_34472,N_30083);
nand U39813 (N_39813,N_31381,N_33069);
or U39814 (N_39814,N_31885,N_32772);
xnor U39815 (N_39815,N_31894,N_31498);
and U39816 (N_39816,N_30679,N_32906);
nand U39817 (N_39817,N_31002,N_34806);
nand U39818 (N_39818,N_31355,N_32990);
and U39819 (N_39819,N_32762,N_34199);
nand U39820 (N_39820,N_30374,N_31066);
nor U39821 (N_39821,N_33422,N_30600);
xor U39822 (N_39822,N_32628,N_34317);
xor U39823 (N_39823,N_31130,N_30842);
nor U39824 (N_39824,N_32272,N_33911);
nor U39825 (N_39825,N_31522,N_33708);
nand U39826 (N_39826,N_31892,N_30255);
nor U39827 (N_39827,N_30606,N_32379);
and U39828 (N_39828,N_31682,N_33369);
xor U39829 (N_39829,N_34084,N_33430);
xor U39830 (N_39830,N_34034,N_32632);
or U39831 (N_39831,N_33524,N_33923);
nor U39832 (N_39832,N_34121,N_32072);
or U39833 (N_39833,N_32792,N_31640);
nand U39834 (N_39834,N_33616,N_34010);
or U39835 (N_39835,N_31849,N_31365);
xor U39836 (N_39836,N_30062,N_32587);
nor U39837 (N_39837,N_31904,N_31798);
and U39838 (N_39838,N_32203,N_34969);
and U39839 (N_39839,N_30133,N_32538);
xnor U39840 (N_39840,N_30198,N_31923);
and U39841 (N_39841,N_30793,N_31666);
nand U39842 (N_39842,N_34582,N_34429);
xnor U39843 (N_39843,N_32202,N_34860);
nand U39844 (N_39844,N_31958,N_34476);
xor U39845 (N_39845,N_31375,N_34564);
nor U39846 (N_39846,N_30216,N_30314);
or U39847 (N_39847,N_32252,N_32128);
or U39848 (N_39848,N_32512,N_31843);
xnor U39849 (N_39849,N_32977,N_32254);
nor U39850 (N_39850,N_31106,N_30547);
nand U39851 (N_39851,N_34311,N_32968);
or U39852 (N_39852,N_33152,N_34167);
nand U39853 (N_39853,N_31795,N_34375);
nand U39854 (N_39854,N_30863,N_30239);
or U39855 (N_39855,N_34012,N_31029);
or U39856 (N_39856,N_32174,N_32516);
or U39857 (N_39857,N_34564,N_32946);
or U39858 (N_39858,N_34243,N_31867);
nand U39859 (N_39859,N_32658,N_34383);
nor U39860 (N_39860,N_31586,N_32715);
nand U39861 (N_39861,N_30068,N_32277);
nand U39862 (N_39862,N_33397,N_34265);
or U39863 (N_39863,N_32415,N_30590);
nand U39864 (N_39864,N_32095,N_33259);
and U39865 (N_39865,N_33445,N_30696);
and U39866 (N_39866,N_31942,N_32791);
or U39867 (N_39867,N_30938,N_31430);
nor U39868 (N_39868,N_32726,N_32751);
and U39869 (N_39869,N_33420,N_33703);
and U39870 (N_39870,N_32856,N_34894);
and U39871 (N_39871,N_34059,N_34060);
nand U39872 (N_39872,N_31609,N_34015);
and U39873 (N_39873,N_34927,N_33920);
xor U39874 (N_39874,N_32951,N_34205);
nor U39875 (N_39875,N_33025,N_30770);
nor U39876 (N_39876,N_33169,N_34824);
xor U39877 (N_39877,N_34062,N_33851);
and U39878 (N_39878,N_34505,N_30644);
nor U39879 (N_39879,N_30981,N_32771);
nor U39880 (N_39880,N_34348,N_31460);
xor U39881 (N_39881,N_33808,N_32284);
or U39882 (N_39882,N_31190,N_34622);
nand U39883 (N_39883,N_32983,N_32214);
or U39884 (N_39884,N_33606,N_32498);
and U39885 (N_39885,N_32631,N_32412);
nand U39886 (N_39886,N_30060,N_30862);
nor U39887 (N_39887,N_33962,N_30562);
nor U39888 (N_39888,N_30788,N_34054);
nor U39889 (N_39889,N_32395,N_32882);
nand U39890 (N_39890,N_30270,N_32668);
nand U39891 (N_39891,N_30273,N_31248);
or U39892 (N_39892,N_30908,N_34124);
xnor U39893 (N_39893,N_30466,N_34866);
and U39894 (N_39894,N_32801,N_32992);
and U39895 (N_39895,N_31495,N_30186);
or U39896 (N_39896,N_33768,N_32501);
xor U39897 (N_39897,N_32705,N_32212);
and U39898 (N_39898,N_33019,N_33349);
nand U39899 (N_39899,N_30153,N_34565);
nand U39900 (N_39900,N_31908,N_33649);
and U39901 (N_39901,N_33007,N_34852);
xor U39902 (N_39902,N_32481,N_30529);
and U39903 (N_39903,N_34509,N_31389);
nand U39904 (N_39904,N_34184,N_34036);
or U39905 (N_39905,N_32371,N_33779);
nand U39906 (N_39906,N_33220,N_31598);
nor U39907 (N_39907,N_33198,N_34509);
nor U39908 (N_39908,N_30915,N_34088);
or U39909 (N_39909,N_30777,N_30307);
nor U39910 (N_39910,N_33175,N_30527);
or U39911 (N_39911,N_34604,N_31481);
nand U39912 (N_39912,N_33224,N_33765);
nor U39913 (N_39913,N_30157,N_34558);
nor U39914 (N_39914,N_32505,N_34977);
or U39915 (N_39915,N_30442,N_32445);
xor U39916 (N_39916,N_31165,N_33765);
or U39917 (N_39917,N_30638,N_32121);
xor U39918 (N_39918,N_30101,N_30104);
nor U39919 (N_39919,N_30726,N_34706);
nand U39920 (N_39920,N_32014,N_33360);
or U39921 (N_39921,N_32814,N_33898);
nand U39922 (N_39922,N_31419,N_34659);
and U39923 (N_39923,N_32118,N_32942);
or U39924 (N_39924,N_31129,N_32208);
and U39925 (N_39925,N_34476,N_31733);
nor U39926 (N_39926,N_31825,N_33307);
nor U39927 (N_39927,N_33250,N_31932);
nand U39928 (N_39928,N_31849,N_34702);
xor U39929 (N_39929,N_31994,N_33586);
or U39930 (N_39930,N_32962,N_30578);
and U39931 (N_39931,N_33407,N_33742);
nor U39932 (N_39932,N_31915,N_32271);
and U39933 (N_39933,N_31881,N_32076);
nand U39934 (N_39934,N_32853,N_32517);
xnor U39935 (N_39935,N_34673,N_32740);
nor U39936 (N_39936,N_34273,N_31644);
xnor U39937 (N_39937,N_30667,N_31091);
and U39938 (N_39938,N_34062,N_33416);
or U39939 (N_39939,N_34132,N_32971);
nand U39940 (N_39940,N_32893,N_34635);
and U39941 (N_39941,N_31278,N_30011);
nand U39942 (N_39942,N_30755,N_32284);
xnor U39943 (N_39943,N_33505,N_34862);
nor U39944 (N_39944,N_33399,N_30508);
nor U39945 (N_39945,N_33104,N_30047);
and U39946 (N_39946,N_34926,N_30787);
xnor U39947 (N_39947,N_30254,N_31093);
nor U39948 (N_39948,N_33656,N_32495);
nand U39949 (N_39949,N_32569,N_30643);
xor U39950 (N_39950,N_34727,N_30890);
or U39951 (N_39951,N_33794,N_33562);
nor U39952 (N_39952,N_31535,N_30046);
and U39953 (N_39953,N_30115,N_31187);
xnor U39954 (N_39954,N_32878,N_32864);
or U39955 (N_39955,N_32844,N_32016);
nor U39956 (N_39956,N_31907,N_33308);
and U39957 (N_39957,N_34109,N_32686);
xnor U39958 (N_39958,N_33332,N_33778);
nor U39959 (N_39959,N_34225,N_34487);
or U39960 (N_39960,N_34005,N_34921);
xnor U39961 (N_39961,N_30040,N_30698);
or U39962 (N_39962,N_33695,N_34231);
nand U39963 (N_39963,N_34062,N_30241);
nor U39964 (N_39964,N_34520,N_33774);
or U39965 (N_39965,N_31375,N_33359);
or U39966 (N_39966,N_30659,N_30088);
or U39967 (N_39967,N_33181,N_34964);
nor U39968 (N_39968,N_33931,N_30940);
or U39969 (N_39969,N_30882,N_34594);
xnor U39970 (N_39970,N_34069,N_31550);
or U39971 (N_39971,N_33432,N_30353);
nor U39972 (N_39972,N_33405,N_32796);
or U39973 (N_39973,N_32914,N_32601);
xnor U39974 (N_39974,N_33136,N_33862);
or U39975 (N_39975,N_31617,N_31729);
nor U39976 (N_39976,N_32657,N_33964);
nor U39977 (N_39977,N_33203,N_34626);
or U39978 (N_39978,N_31639,N_32389);
nand U39979 (N_39979,N_31918,N_32169);
nand U39980 (N_39980,N_30561,N_32250);
nand U39981 (N_39981,N_30057,N_32777);
or U39982 (N_39982,N_30018,N_30647);
nand U39983 (N_39983,N_31124,N_30426);
nor U39984 (N_39984,N_31726,N_34007);
or U39985 (N_39985,N_33042,N_34255);
and U39986 (N_39986,N_30247,N_33964);
xor U39987 (N_39987,N_33232,N_32892);
and U39988 (N_39988,N_33797,N_33451);
or U39989 (N_39989,N_32684,N_32683);
nor U39990 (N_39990,N_33678,N_31211);
and U39991 (N_39991,N_33576,N_30839);
nand U39992 (N_39992,N_34633,N_30026);
nor U39993 (N_39993,N_30886,N_31281);
nand U39994 (N_39994,N_34769,N_30813);
nand U39995 (N_39995,N_33139,N_31380);
nand U39996 (N_39996,N_34236,N_30132);
or U39997 (N_39997,N_33014,N_30943);
or U39998 (N_39998,N_31924,N_34680);
nor U39999 (N_39999,N_34808,N_34941);
nand U40000 (N_40000,N_36398,N_38839);
nand U40001 (N_40001,N_37539,N_36290);
nor U40002 (N_40002,N_35669,N_37383);
and U40003 (N_40003,N_37562,N_35073);
or U40004 (N_40004,N_35635,N_38636);
nand U40005 (N_40005,N_39809,N_36320);
xor U40006 (N_40006,N_36709,N_38934);
and U40007 (N_40007,N_35907,N_38215);
or U40008 (N_40008,N_39736,N_36673);
nor U40009 (N_40009,N_35279,N_37196);
nor U40010 (N_40010,N_35020,N_39616);
nor U40011 (N_40011,N_38876,N_39070);
and U40012 (N_40012,N_38416,N_36161);
nand U40013 (N_40013,N_36499,N_36694);
or U40014 (N_40014,N_37857,N_35555);
xor U40015 (N_40015,N_37997,N_37463);
or U40016 (N_40016,N_35963,N_37325);
nand U40017 (N_40017,N_39225,N_37838);
and U40018 (N_40018,N_36753,N_36442);
and U40019 (N_40019,N_35303,N_35546);
nor U40020 (N_40020,N_39502,N_37610);
nor U40021 (N_40021,N_39247,N_37555);
or U40022 (N_40022,N_36867,N_39347);
nand U40023 (N_40023,N_36010,N_35231);
xor U40024 (N_40024,N_36011,N_35184);
nor U40025 (N_40025,N_38570,N_37906);
xor U40026 (N_40026,N_38527,N_35914);
nand U40027 (N_40027,N_37047,N_37337);
nand U40028 (N_40028,N_37314,N_37986);
nand U40029 (N_40029,N_39937,N_37531);
xnor U40030 (N_40030,N_37330,N_35026);
and U40031 (N_40031,N_35648,N_36949);
xor U40032 (N_40032,N_35282,N_37661);
or U40033 (N_40033,N_39729,N_37220);
or U40034 (N_40034,N_39186,N_38703);
nor U40035 (N_40035,N_36569,N_36587);
and U40036 (N_40036,N_36094,N_37454);
and U40037 (N_40037,N_35786,N_35789);
nand U40038 (N_40038,N_36080,N_35512);
xor U40039 (N_40039,N_36558,N_37421);
or U40040 (N_40040,N_37859,N_38093);
or U40041 (N_40041,N_39984,N_38517);
nor U40042 (N_40042,N_36821,N_38159);
and U40043 (N_40043,N_37420,N_39345);
xor U40044 (N_40044,N_36904,N_37429);
and U40045 (N_40045,N_38658,N_39413);
xor U40046 (N_40046,N_39739,N_37790);
nor U40047 (N_40047,N_39865,N_36229);
and U40048 (N_40048,N_35116,N_37427);
or U40049 (N_40049,N_38118,N_38834);
nand U40050 (N_40050,N_35199,N_37450);
nand U40051 (N_40051,N_37213,N_38523);
xnor U40052 (N_40052,N_35081,N_35652);
nor U40053 (N_40053,N_39294,N_38098);
or U40054 (N_40054,N_35079,N_37035);
or U40055 (N_40055,N_37726,N_36150);
xnor U40056 (N_40056,N_37161,N_36259);
nor U40057 (N_40057,N_35050,N_36335);
or U40058 (N_40058,N_36984,N_39105);
and U40059 (N_40059,N_35502,N_35008);
nor U40060 (N_40060,N_37260,N_39101);
and U40061 (N_40061,N_38469,N_38131);
and U40062 (N_40062,N_35978,N_36318);
xnor U40063 (N_40063,N_36960,N_35385);
xor U40064 (N_40064,N_35695,N_37993);
and U40065 (N_40065,N_35513,N_36073);
or U40066 (N_40066,N_35554,N_39781);
xnor U40067 (N_40067,N_37936,N_38544);
nand U40068 (N_40068,N_39769,N_36533);
and U40069 (N_40069,N_39807,N_36248);
and U40070 (N_40070,N_38984,N_37579);
nand U40071 (N_40071,N_38260,N_35010);
nand U40072 (N_40072,N_38513,N_39673);
xor U40073 (N_40073,N_38334,N_36524);
and U40074 (N_40074,N_35196,N_36899);
and U40075 (N_40075,N_35895,N_38535);
and U40076 (N_40076,N_35204,N_37843);
xor U40077 (N_40077,N_39743,N_39987);
xnor U40078 (N_40078,N_36830,N_35739);
xnor U40079 (N_40079,N_36112,N_37322);
or U40080 (N_40080,N_37292,N_35981);
nor U40081 (N_40081,N_36119,N_38370);
nand U40082 (N_40082,N_35037,N_36403);
xor U40083 (N_40083,N_36205,N_35329);
nand U40084 (N_40084,N_39595,N_39112);
nand U40085 (N_40085,N_39530,N_35190);
nand U40086 (N_40086,N_35832,N_38423);
nand U40087 (N_40087,N_35780,N_39857);
nor U40088 (N_40088,N_35818,N_38904);
xor U40089 (N_40089,N_35115,N_35839);
and U40090 (N_40090,N_37987,N_38475);
xor U40091 (N_40091,N_36246,N_39031);
nor U40092 (N_40092,N_36693,N_39237);
nand U40093 (N_40093,N_38805,N_36251);
xnor U40094 (N_40094,N_36141,N_39951);
and U40095 (N_40095,N_38052,N_38936);
nand U40096 (N_40096,N_38433,N_38239);
and U40097 (N_40097,N_38263,N_37373);
and U40098 (N_40098,N_36514,N_35210);
or U40099 (N_40099,N_36828,N_35176);
xnor U40100 (N_40100,N_37946,N_38482);
or U40101 (N_40101,N_35468,N_39024);
xor U40102 (N_40102,N_39864,N_37611);
nor U40103 (N_40103,N_35574,N_36303);
nand U40104 (N_40104,N_36299,N_38476);
and U40105 (N_40105,N_38883,N_36085);
and U40106 (N_40106,N_38025,N_38778);
nand U40107 (N_40107,N_36404,N_38486);
and U40108 (N_40108,N_38672,N_38086);
or U40109 (N_40109,N_35684,N_36545);
nand U40110 (N_40110,N_36738,N_36761);
xnor U40111 (N_40111,N_39917,N_37558);
or U40112 (N_40112,N_38851,N_37564);
nor U40113 (N_40113,N_37310,N_37316);
or U40114 (N_40114,N_38646,N_39722);
nor U40115 (N_40115,N_35972,N_38424);
xnor U40116 (N_40116,N_37074,N_35371);
nor U40117 (N_40117,N_39157,N_36659);
xor U40118 (N_40118,N_35606,N_36104);
and U40119 (N_40119,N_39128,N_37528);
nand U40120 (N_40120,N_37862,N_35382);
xnor U40121 (N_40121,N_36863,N_39171);
nand U40122 (N_40122,N_38706,N_35137);
nand U40123 (N_40123,N_39591,N_38584);
nor U40124 (N_40124,N_37468,N_38384);
nor U40125 (N_40125,N_39188,N_37389);
or U40126 (N_40126,N_35364,N_39215);
nand U40127 (N_40127,N_37797,N_36167);
nor U40128 (N_40128,N_35362,N_37103);
and U40129 (N_40129,N_36736,N_38701);
nor U40130 (N_40130,N_37169,N_36183);
xor U40131 (N_40131,N_36009,N_39652);
or U40132 (N_40132,N_36622,N_37460);
nand U40133 (N_40133,N_39371,N_37118);
and U40134 (N_40134,N_38142,N_35423);
and U40135 (N_40135,N_39922,N_38329);
or U40136 (N_40136,N_36768,N_39478);
nor U40137 (N_40137,N_39427,N_37633);
or U40138 (N_40138,N_38575,N_37930);
and U40139 (N_40139,N_37979,N_38790);
or U40140 (N_40140,N_39683,N_36342);
xnor U40141 (N_40141,N_37445,N_38090);
xnor U40142 (N_40142,N_37925,N_36084);
and U40143 (N_40143,N_35992,N_37822);
nand U40144 (N_40144,N_39764,N_37876);
nor U40145 (N_40145,N_35219,N_39709);
and U40146 (N_40146,N_39222,N_36950);
or U40147 (N_40147,N_36123,N_35367);
xnor U40148 (N_40148,N_38945,N_39156);
nor U40149 (N_40149,N_37263,N_37407);
and U40150 (N_40150,N_38205,N_35339);
and U40151 (N_40151,N_36317,N_39023);
nand U40152 (N_40152,N_36149,N_35658);
nor U40153 (N_40153,N_38234,N_38900);
nor U40154 (N_40154,N_37985,N_37826);
and U40155 (N_40155,N_35634,N_36557);
or U40156 (N_40156,N_39617,N_36102);
or U40157 (N_40157,N_37134,N_35244);
and U40158 (N_40158,N_36628,N_36629);
nand U40159 (N_40159,N_38355,N_38655);
xnor U40160 (N_40160,N_36647,N_38328);
nor U40161 (N_40161,N_38966,N_38866);
and U40162 (N_40162,N_36354,N_36776);
nor U40163 (N_40163,N_35054,N_35350);
xnor U40164 (N_40164,N_38766,N_36348);
and U40165 (N_40165,N_36630,N_35736);
or U40166 (N_40166,N_39445,N_37761);
nand U40167 (N_40167,N_37347,N_39520);
or U40168 (N_40168,N_38878,N_39688);
xor U40169 (N_40169,N_39968,N_35337);
nand U40170 (N_40170,N_36735,N_36646);
nand U40171 (N_40171,N_35173,N_35194);
nor U40172 (N_40172,N_38971,N_39964);
or U40173 (N_40173,N_36593,N_37198);
nor U40174 (N_40174,N_38693,N_35524);
and U40175 (N_40175,N_35482,N_37242);
xnor U40176 (N_40176,N_37493,N_37848);
nand U40177 (N_40177,N_36853,N_38682);
and U40178 (N_40178,N_39077,N_36577);
nand U40179 (N_40179,N_36063,N_36210);
nor U40180 (N_40180,N_38689,N_37350);
or U40181 (N_40181,N_37135,N_38375);
nand U40182 (N_40182,N_38303,N_38942);
nor U40183 (N_40183,N_36395,N_39376);
and U40184 (N_40184,N_36555,N_36717);
or U40185 (N_40185,N_37776,N_36969);
nor U40186 (N_40186,N_36741,N_35436);
or U40187 (N_40187,N_38014,N_39974);
and U40188 (N_40188,N_39515,N_38799);
and U40189 (N_40189,N_36169,N_35563);
and U40190 (N_40190,N_37805,N_35175);
xnor U40191 (N_40191,N_35192,N_36013);
nor U40192 (N_40192,N_35751,N_39369);
or U40193 (N_40193,N_38181,N_37698);
nand U40194 (N_40194,N_36507,N_39009);
or U40195 (N_40195,N_38882,N_37551);
nor U40196 (N_40196,N_39934,N_38922);
xnor U40197 (N_40197,N_35307,N_38187);
and U40198 (N_40198,N_36531,N_39249);
xnor U40199 (N_40199,N_38796,N_37354);
or U40200 (N_40200,N_36605,N_36544);
xor U40201 (N_40201,N_35582,N_35944);
or U40202 (N_40202,N_35363,N_39501);
nor U40203 (N_40203,N_38522,N_39557);
nand U40204 (N_40204,N_38121,N_39287);
nor U40205 (N_40205,N_36083,N_35139);
or U40206 (N_40206,N_37044,N_38925);
nand U40207 (N_40207,N_35141,N_39223);
xor U40208 (N_40208,N_35626,N_37307);
or U40209 (N_40209,N_35263,N_38064);
nand U40210 (N_40210,N_35660,N_37148);
nor U40211 (N_40211,N_39885,N_36105);
or U40212 (N_40212,N_38598,N_36614);
and U40213 (N_40213,N_37875,N_37889);
and U40214 (N_40214,N_37609,N_36196);
nor U40215 (N_40215,N_38609,N_35384);
xor U40216 (N_40216,N_37130,N_35179);
xor U40217 (N_40217,N_38097,N_39882);
and U40218 (N_40218,N_39162,N_36526);
nor U40219 (N_40219,N_37916,N_36539);
nand U40220 (N_40220,N_37825,N_37368);
nand U40221 (N_40221,N_39025,N_36812);
xnor U40222 (N_40222,N_37115,N_39317);
nand U40223 (N_40223,N_37385,N_38286);
or U40224 (N_40224,N_35955,N_39653);
or U40225 (N_40225,N_37750,N_35603);
nor U40226 (N_40226,N_35323,N_39060);
nor U40227 (N_40227,N_35619,N_37442);
nor U40228 (N_40228,N_38002,N_38128);
nand U40229 (N_40229,N_39626,N_36338);
and U40230 (N_40230,N_37593,N_36370);
nand U40231 (N_40231,N_36356,N_39503);
and U40232 (N_40232,N_38694,N_39375);
and U40233 (N_40233,N_37613,N_35998);
nand U40234 (N_40234,N_39842,N_37447);
nor U40235 (N_40235,N_36291,N_35781);
nand U40236 (N_40236,N_39644,N_39126);
xor U40237 (N_40237,N_39867,N_36896);
or U40238 (N_40238,N_36885,N_37273);
or U40239 (N_40239,N_35707,N_36719);
xor U40240 (N_40240,N_35971,N_35728);
xor U40241 (N_40241,N_39786,N_36732);
nor U40242 (N_40242,N_37342,N_37175);
xor U40243 (N_40243,N_38588,N_38039);
or U40244 (N_40244,N_39839,N_35357);
nand U40245 (N_40245,N_36799,N_36315);
nand U40246 (N_40246,N_36176,N_37366);
nor U40247 (N_40247,N_35248,N_36093);
xor U40248 (N_40248,N_35505,N_37785);
nor U40249 (N_40249,N_35968,N_38510);
nor U40250 (N_40250,N_38754,N_36602);
nor U40251 (N_40251,N_39082,N_39311);
nor U40252 (N_40252,N_38688,N_38429);
and U40253 (N_40253,N_38770,N_37305);
nand U40254 (N_40254,N_37861,N_39339);
xor U40255 (N_40255,N_35481,N_39602);
xnor U40256 (N_40256,N_36855,N_39055);
or U40257 (N_40257,N_36683,N_38727);
nor U40258 (N_40258,N_36304,N_37852);
and U40259 (N_40259,N_39872,N_35366);
nor U40260 (N_40260,N_39266,N_35095);
xnor U40261 (N_40261,N_39458,N_38854);
nand U40262 (N_40262,N_38105,N_39122);
and U40263 (N_40263,N_37370,N_36752);
nand U40264 (N_40264,N_38845,N_37332);
xnor U40265 (N_40265,N_36771,N_39746);
or U40266 (N_40266,N_39142,N_38896);
xnor U40267 (N_40267,N_36434,N_35327);
xor U40268 (N_40268,N_39620,N_35819);
xor U40269 (N_40269,N_39147,N_35397);
nor U40270 (N_40270,N_35762,N_36754);
nor U40271 (N_40271,N_38902,N_35683);
or U40272 (N_40272,N_35138,N_36898);
and U40273 (N_40273,N_36826,N_35414);
or U40274 (N_40274,N_37717,N_36405);
and U40275 (N_40275,N_39267,N_36012);
xnor U40276 (N_40276,N_38855,N_37003);
nor U40277 (N_40277,N_37699,N_38255);
and U40278 (N_40278,N_37098,N_39555);
nand U40279 (N_40279,N_35039,N_39404);
nand U40280 (N_40280,N_37070,N_39331);
nand U40281 (N_40281,N_35516,N_37749);
nand U40282 (N_40282,N_35325,N_37662);
xor U40283 (N_40283,N_38911,N_35458);
or U40284 (N_40284,N_38524,N_38521);
or U40285 (N_40285,N_39394,N_39381);
and U40286 (N_40286,N_38982,N_37833);
xor U40287 (N_40287,N_37006,N_37657);
or U40288 (N_40288,N_36854,N_39999);
nand U40289 (N_40289,N_37435,N_39944);
nand U40290 (N_40290,N_37246,N_39732);
and U40291 (N_40291,N_39001,N_36897);
nor U40292 (N_40292,N_39412,N_38626);
xnor U40293 (N_40293,N_38279,N_39076);
nor U40294 (N_40294,N_37894,N_36294);
nand U40295 (N_40295,N_35016,N_38258);
nor U40296 (N_40296,N_39610,N_38846);
and U40297 (N_40297,N_38109,N_38048);
and U40298 (N_40298,N_35617,N_39314);
nand U40299 (N_40299,N_35831,N_37064);
nor U40300 (N_40300,N_39430,N_37667);
xnor U40301 (N_40301,N_36822,N_37267);
nor U40302 (N_40302,N_38226,N_38251);
nand U40303 (N_40303,N_37126,N_39890);
and U40304 (N_40304,N_36877,N_38055);
nor U40305 (N_40305,N_37204,N_36494);
and U40306 (N_40306,N_35668,N_36783);
nand U40307 (N_40307,N_36226,N_38257);
or U40308 (N_40308,N_35561,N_37642);
and U40309 (N_40309,N_35101,N_38027);
xnor U40310 (N_40310,N_37959,N_38530);
or U40311 (N_40311,N_37693,N_37587);
or U40312 (N_40312,N_39093,N_36277);
nand U40313 (N_40313,N_37666,N_39131);
nor U40314 (N_40314,N_38997,N_35270);
nor U40315 (N_40315,N_38087,N_37492);
and U40316 (N_40316,N_36801,N_38946);
xor U40317 (N_40317,N_37380,N_36059);
nand U40318 (N_40318,N_37612,N_38947);
or U40319 (N_40319,N_37628,N_36661);
nor U40320 (N_40320,N_38204,N_38618);
nand U40321 (N_40321,N_38833,N_36037);
xnor U40322 (N_40322,N_39810,N_38478);
xor U40323 (N_40323,N_37835,N_39702);
nor U40324 (N_40324,N_37107,N_36146);
or U40325 (N_40325,N_35065,N_37723);
nand U40326 (N_40326,N_37414,N_38341);
and U40327 (N_40327,N_36839,N_35457);
nor U40328 (N_40328,N_36087,N_37804);
nand U40329 (N_40329,N_37422,N_38276);
and U40330 (N_40330,N_37309,N_36803);
xor U40331 (N_40331,N_35857,N_38421);
nand U40332 (N_40332,N_35551,N_36720);
nand U40333 (N_40333,N_39187,N_39067);
nand U40334 (N_40334,N_38172,N_38309);
xnor U40335 (N_40335,N_38988,N_38981);
nand U40336 (N_40336,N_35718,N_36328);
or U40337 (N_40337,N_39808,N_37919);
and U40338 (N_40338,N_38932,N_35259);
xnor U40339 (N_40339,N_38256,N_37469);
or U40340 (N_40340,N_35509,N_36939);
nand U40341 (N_40341,N_39103,N_39465);
xnor U40342 (N_40342,N_39210,N_38442);
nor U40343 (N_40343,N_39948,N_38508);
nand U40344 (N_40344,N_38100,N_35402);
nand U40345 (N_40345,N_37046,N_36228);
nand U40346 (N_40346,N_36734,N_39166);
xnor U40347 (N_40347,N_37855,N_35461);
xor U40348 (N_40348,N_36814,N_39700);
nand U40349 (N_40349,N_35153,N_39387);
nand U40350 (N_40350,N_38554,N_35009);
nand U40351 (N_40351,N_39561,N_38166);
or U40352 (N_40352,N_36671,N_36561);
and U40353 (N_40353,N_37284,N_38975);
nand U40354 (N_40354,N_37762,N_35926);
nand U40355 (N_40355,N_39179,N_38067);
nor U40356 (N_40356,N_35433,N_35272);
nor U40357 (N_40357,N_38374,N_36053);
nor U40358 (N_40358,N_39470,N_38707);
nand U40359 (N_40359,N_39705,N_35804);
and U40360 (N_40360,N_36536,N_38242);
xor U40361 (N_40361,N_35042,N_35912);
xnor U40362 (N_40362,N_37999,N_37482);
xnor U40363 (N_40363,N_37923,N_39628);
nand U40364 (N_40364,N_38669,N_38488);
nor U40365 (N_40365,N_35790,N_38886);
nand U40366 (N_40366,N_35427,N_39125);
or U40367 (N_40367,N_37224,N_39850);
or U40368 (N_40368,N_39170,N_39203);
or U40369 (N_40369,N_39957,N_36952);
xnor U40370 (N_40370,N_37849,N_39395);
or U40371 (N_40371,N_35390,N_39416);
and U40372 (N_40372,N_36723,N_38280);
xor U40373 (N_40373,N_35149,N_39648);
nor U40374 (N_40374,N_35867,N_39611);
nand U40375 (N_40375,N_36447,N_36810);
nand U40376 (N_40376,N_39059,N_39144);
and U40377 (N_40377,N_35759,N_38663);
nand U40378 (N_40378,N_37245,N_38603);
xor U40379 (N_40379,N_37943,N_39449);
or U40380 (N_40380,N_36745,N_36222);
xnor U40381 (N_40381,N_35150,N_36583);
or U40382 (N_40382,N_35351,N_37568);
and U40383 (N_40383,N_39820,N_37358);
nand U40384 (N_40384,N_39932,N_36065);
xnor U40385 (N_40385,N_39986,N_38901);
nand U40386 (N_40386,N_38681,N_38697);
or U40387 (N_40387,N_38661,N_36714);
xnor U40388 (N_40388,N_38801,N_39967);
xnor U40389 (N_40389,N_36833,N_35993);
nor U40390 (N_40390,N_38017,N_38895);
and U40391 (N_40391,N_39289,N_39747);
and U40392 (N_40392,N_35227,N_39522);
and U40393 (N_40393,N_36932,N_36326);
or U40394 (N_40394,N_35701,N_35534);
nand U40395 (N_40395,N_36766,N_36684);
nand U40396 (N_40396,N_36069,N_37913);
or U40397 (N_40397,N_37372,N_38292);
or U40398 (N_40398,N_35662,N_35594);
nand U40399 (N_40399,N_37105,N_39913);
xnor U40400 (N_40400,N_35726,N_38129);
nand U40401 (N_40401,N_35164,N_38208);
nand U40402 (N_40402,N_35913,N_37183);
xor U40403 (N_40403,N_36159,N_39823);
and U40404 (N_40404,N_36199,N_38459);
and U40405 (N_40405,N_39040,N_37159);
nor U40406 (N_40406,N_38371,N_38505);
nand U40407 (N_40407,N_38147,N_35161);
nand U40408 (N_40408,N_36608,N_37547);
or U40409 (N_40409,N_37145,N_36708);
xnor U40410 (N_40410,N_35833,N_39930);
or U40411 (N_40411,N_39889,N_37343);
and U40412 (N_40412,N_38792,N_38720);
nor U40413 (N_40413,N_36690,N_35166);
xnor U40414 (N_40414,N_39533,N_38216);
and U40415 (N_40415,N_37257,N_37068);
nand U40416 (N_40416,N_36422,N_37841);
or U40417 (N_40417,N_37742,N_35374);
nand U40418 (N_40418,N_39834,N_38124);
nor U40419 (N_40419,N_37449,N_39432);
and U40420 (N_40420,N_39956,N_35247);
nor U40421 (N_40421,N_38311,N_39181);
nand U40422 (N_40422,N_37125,N_35504);
or U40423 (N_40423,N_36120,N_36400);
nand U40424 (N_40424,N_37668,N_38822);
xnor U40425 (N_40425,N_39123,N_39022);
and U40426 (N_40426,N_35454,N_38835);
or U40427 (N_40427,N_36945,N_38927);
nand U40428 (N_40428,N_36194,N_37234);
or U40429 (N_40429,N_36528,N_38293);
and U40430 (N_40430,N_35269,N_38567);
and U40431 (N_40431,N_39288,N_39164);
nor U40432 (N_40432,N_37880,N_39488);
nand U40433 (N_40433,N_36962,N_38321);
nand U40434 (N_40434,N_39783,N_35851);
xnor U40435 (N_40435,N_35290,N_37928);
or U40436 (N_40436,N_36800,N_39468);
xnor U40437 (N_40437,N_39218,N_39609);
xnor U40438 (N_40438,N_37743,N_35964);
nand U40439 (N_40439,N_37099,N_35157);
xnor U40440 (N_40440,N_36364,N_35345);
xnor U40441 (N_40441,N_39075,N_36232);
xnor U40442 (N_40442,N_36110,N_39525);
nand U40443 (N_40443,N_36594,N_38220);
xor U40444 (N_40444,N_38777,N_38036);
nand U40445 (N_40445,N_39970,N_39771);
or U40446 (N_40446,N_37541,N_36079);
nand U40447 (N_40447,N_36679,N_38150);
nand U40448 (N_40448,N_35887,N_35674);
nand U40449 (N_40449,N_35782,N_35407);
xnor U40450 (N_40450,N_38031,N_37081);
or U40451 (N_40451,N_38526,N_37972);
nand U40452 (N_40452,N_35796,N_35375);
nand U40453 (N_40453,N_38477,N_35649);
xor U40454 (N_40454,N_37738,N_37225);
nand U40455 (N_40455,N_38955,N_35168);
xor U40456 (N_40456,N_39719,N_35775);
nand U40457 (N_40457,N_35543,N_35680);
xor U40458 (N_40458,N_38748,N_39466);
nor U40459 (N_40459,N_35040,N_39402);
or U40460 (N_40460,N_35464,N_37878);
xnor U40461 (N_40461,N_38495,N_36115);
or U40462 (N_40462,N_35395,N_37388);
nand U40463 (N_40463,N_37967,N_35178);
and U40464 (N_40464,N_37152,N_38736);
nor U40465 (N_40465,N_39351,N_39028);
and U40466 (N_40466,N_35836,N_38007);
nand U40467 (N_40467,N_38361,N_36100);
and U40468 (N_40468,N_39320,N_35297);
and U40469 (N_40469,N_38959,N_38812);
xnor U40470 (N_40470,N_38960,N_39835);
and U40471 (N_40471,N_38667,N_35428);
xor U40472 (N_40472,N_35693,N_38358);
or U40473 (N_40473,N_36168,N_38921);
nor U40474 (N_40474,N_35240,N_38116);
or U40475 (N_40475,N_36249,N_36691);
nand U40476 (N_40476,N_39753,N_35613);
nand U40477 (N_40477,N_35142,N_39548);
or U40478 (N_40478,N_35156,N_37237);
or U40479 (N_40479,N_38454,N_37032);
and U40480 (N_40480,N_39480,N_37236);
and U40481 (N_40481,N_39265,N_38949);
nor U40482 (N_40482,N_37629,N_39551);
and U40483 (N_40483,N_39507,N_35273);
or U40484 (N_40484,N_37489,N_38101);
xor U40485 (N_40485,N_36770,N_37641);
xor U40486 (N_40486,N_35379,N_38843);
nand U40487 (N_40487,N_37965,N_37259);
or U40488 (N_40488,N_39035,N_39392);
nor U40489 (N_40489,N_39639,N_35041);
nand U40490 (N_40490,N_35003,N_37637);
nor U40491 (N_40491,N_39097,N_39645);
nand U40492 (N_40492,N_38114,N_37129);
and U40493 (N_40493,N_35591,N_36439);
nand U40494 (N_40494,N_39056,N_35144);
nor U40495 (N_40495,N_35152,N_39681);
nor U40496 (N_40496,N_38506,N_38308);
nand U40497 (N_40497,N_38970,N_35201);
or U40498 (N_40498,N_36596,N_38958);
xnor U40499 (N_40499,N_39262,N_38253);
or U40500 (N_40500,N_36490,N_36349);
and U40501 (N_40501,N_39497,N_39316);
or U40502 (N_40502,N_37019,N_36913);
xor U40503 (N_40503,N_38364,N_36293);
nand U40504 (N_40504,N_38288,N_37166);
nor U40505 (N_40505,N_36756,N_37703);
nor U40506 (N_40506,N_38545,N_35999);
nand U40507 (N_40507,N_36762,N_37094);
xnor U40508 (N_40508,N_38553,N_35532);
or U40509 (N_40509,N_37005,N_38687);
xor U40510 (N_40510,N_35062,N_38277);
nor U40511 (N_40511,N_39299,N_38725);
or U40512 (N_40512,N_38231,N_36675);
and U40513 (N_40513,N_36454,N_38373);
xnor U40514 (N_40514,N_35860,N_36262);
nand U40515 (N_40515,N_37526,N_39789);
and U40516 (N_40516,N_35378,N_39763);
and U40517 (N_40517,N_36721,N_39544);
and U40518 (N_40518,N_37926,N_37167);
and U40519 (N_40519,N_35862,N_38704);
xnor U40520 (N_40520,N_36077,N_38192);
nor U40521 (N_40521,N_39061,N_37519);
xnor U40522 (N_40522,N_39421,N_38444);
and U40523 (N_40523,N_39980,N_37440);
nand U40524 (N_40524,N_35341,N_38152);
nand U40525 (N_40525,N_37050,N_37455);
nand U40526 (N_40526,N_37756,N_38432);
xor U40527 (N_40527,N_39037,N_35437);
or U40528 (N_40528,N_35979,N_37556);
or U40529 (N_40529,N_36862,N_39744);
or U40530 (N_40530,N_37004,N_38115);
nor U40531 (N_40531,N_38624,N_38290);
and U40532 (N_40532,N_39148,N_38148);
and U40533 (N_40533,N_35047,N_35729);
nor U40534 (N_40534,N_35438,N_39996);
or U40535 (N_40535,N_35167,N_36298);
and U40536 (N_40536,N_39301,N_35890);
xnor U40537 (N_40537,N_37741,N_35170);
xnor U40538 (N_40538,N_36642,N_39163);
or U40539 (N_40539,N_39879,N_37590);
and U40540 (N_40540,N_36384,N_35291);
nor U40541 (N_40541,N_35479,N_39441);
xor U40542 (N_40542,N_38189,N_35057);
nand U40543 (N_40543,N_35510,N_36886);
and U40544 (N_40544,N_38411,N_38157);
xnor U40545 (N_40545,N_38924,N_37184);
nand U40546 (N_40546,N_37080,N_36296);
xor U40547 (N_40547,N_36153,N_37989);
xnor U40548 (N_40548,N_37932,N_39699);
or U40549 (N_40549,N_39356,N_37977);
nor U40550 (N_40550,N_37614,N_36278);
and U40551 (N_40551,N_38077,N_39933);
and U40552 (N_40552,N_39500,N_36172);
nor U40553 (N_40553,N_39847,N_35946);
nor U40554 (N_40554,N_37287,N_39659);
or U40555 (N_40555,N_36739,N_37786);
xor U40556 (N_40556,N_37747,N_37057);
nand U40557 (N_40557,N_36934,N_39696);
nor U40558 (N_40558,N_39925,N_37122);
nor U40559 (N_40559,N_35490,N_35493);
nor U40560 (N_40560,N_38396,N_36824);
nand U40561 (N_40561,N_38783,N_35788);
and U40562 (N_40562,N_38765,N_38326);
xor U40563 (N_40563,N_37964,N_35130);
or U40564 (N_40564,N_36931,N_37509);
nand U40565 (N_40565,N_35456,N_36385);
nand U40566 (N_40566,N_37278,N_35431);
xnor U40567 (N_40567,N_37009,N_39400);
nand U40568 (N_40568,N_38793,N_38581);
or U40569 (N_40569,N_36912,N_39836);
and U40570 (N_40570,N_38542,N_38434);
or U40571 (N_40571,N_36758,N_38012);
and U40572 (N_40572,N_36529,N_37029);
nand U40573 (N_40573,N_39667,N_39273);
nor U40574 (N_40574,N_36664,N_38096);
or U40575 (N_40575,N_35349,N_37591);
xnor U40576 (N_40576,N_35217,N_38190);
and U40577 (N_40577,N_37045,N_38363);
nand U40578 (N_40578,N_38972,N_39992);
nor U40579 (N_40579,N_37559,N_37694);
xor U40580 (N_40580,N_39141,N_37239);
nand U40581 (N_40581,N_35522,N_36036);
xor U40582 (N_40582,N_37680,N_37501);
or U40583 (N_40583,N_39483,N_35947);
and U40584 (N_40584,N_35443,N_38635);
nand U40585 (N_40585,N_35148,N_36777);
nand U40586 (N_40586,N_36137,N_35255);
and U40587 (N_40587,N_39439,N_38319);
or U40588 (N_40588,N_38177,N_37708);
xnor U40589 (N_40589,N_36302,N_37486);
xor U40590 (N_40590,N_36117,N_37334);
xnor U40591 (N_40591,N_37364,N_35226);
nand U40592 (N_40592,N_39027,N_38015);
nor U40593 (N_40593,N_37384,N_36920);
nor U40594 (N_40594,N_37321,N_37415);
xnor U40595 (N_40595,N_37574,N_38119);
or U40596 (N_40596,N_39923,N_37842);
and U40597 (N_40597,N_38032,N_36961);
and U40598 (N_40598,N_35442,N_36911);
or U40599 (N_40599,N_37798,N_35756);
nand U40600 (N_40600,N_38764,N_36927);
and U40601 (N_40601,N_37031,N_36990);
and U40602 (N_40602,N_36645,N_39274);
and U40603 (N_40603,N_38024,N_38004);
nor U40604 (N_40604,N_35779,N_38059);
nand U40605 (N_40605,N_39876,N_35903);
nor U40606 (N_40606,N_37018,N_38763);
nor U40607 (N_40607,N_39151,N_38587);
or U40608 (N_40608,N_37768,N_37961);
or U40609 (N_40609,N_35055,N_35904);
and U40610 (N_40610,N_35715,N_37137);
nor U40611 (N_40611,N_36916,N_37378);
xnor U40612 (N_40612,N_37048,N_38425);
or U40613 (N_40613,N_39373,N_38752);
nor U40614 (N_40614,N_36511,N_39359);
and U40615 (N_40615,N_38735,N_38897);
and U40616 (N_40616,N_39924,N_36742);
nand U40617 (N_40617,N_35228,N_37565);
and U40618 (N_40618,N_36215,N_36607);
nor U40619 (N_40619,N_39242,N_36523);
nor U40620 (N_40620,N_37203,N_36211);
nor U40621 (N_40621,N_35957,N_37425);
nand U40622 (N_40622,N_39451,N_39536);
and U40623 (N_40623,N_35763,N_35388);
and U40624 (N_40624,N_37024,N_39297);
and U40625 (N_40625,N_36072,N_36773);
or U40626 (N_40626,N_37827,N_39472);
nor U40627 (N_40627,N_38595,N_37810);
nor U40628 (N_40628,N_38200,N_39905);
nor U40629 (N_40629,N_36846,N_35973);
xnor U40630 (N_40630,N_35394,N_39424);
nor U40631 (N_40631,N_36750,N_37712);
and U40632 (N_40632,N_38091,N_37856);
nor U40633 (N_40633,N_35419,N_37866);
or U40634 (N_40634,N_39408,N_38236);
xnor U40635 (N_40635,N_39100,N_36164);
and U40636 (N_40636,N_36937,N_38448);
and U40637 (N_40637,N_38106,N_39637);
or U40638 (N_40638,N_35891,N_38232);
xor U40639 (N_40639,N_36267,N_36957);
xnor U40640 (N_40640,N_35185,N_35793);
nand U40641 (N_40641,N_35538,N_39590);
nand U40642 (N_40642,N_35823,N_37598);
nand U40643 (N_40643,N_38539,N_36667);
xnor U40644 (N_40644,N_38607,N_38228);
nor U40645 (N_40645,N_38823,N_38739);
or U40646 (N_40646,N_38346,N_37724);
and U40647 (N_40647,N_39647,N_39587);
and U40648 (N_40648,N_37689,N_35991);
xor U40649 (N_40649,N_39594,N_36807);
nand U40650 (N_40650,N_37411,N_37147);
xnor U40651 (N_40651,N_36552,N_39665);
nor U40652 (N_40652,N_38178,N_39793);
nand U40653 (N_40653,N_39825,N_38441);
nor U40654 (N_40654,N_36460,N_39000);
or U40655 (N_40655,N_38928,N_37793);
or U40656 (N_40656,N_38998,N_37918);
xor U40657 (N_40657,N_39496,N_35800);
or U40658 (N_40658,N_37144,N_35246);
xnor U40659 (N_40659,N_36250,N_38880);
nor U40660 (N_40660,N_38775,N_35386);
nand U40661 (N_40661,N_35114,N_38435);
xnor U40662 (N_40662,N_38073,N_38296);
nand U40663 (N_40663,N_38497,N_35415);
nand U40664 (N_40664,N_37860,N_35719);
nand U40665 (N_40665,N_36542,N_37060);
nor U40666 (N_40666,N_38391,N_36551);
nand U40667 (N_40667,N_39152,N_39778);
nor U40668 (N_40668,N_36285,N_36574);
or U40669 (N_40669,N_39605,N_39615);
and U40670 (N_40670,N_36208,N_36831);
nor U40671 (N_40671,N_36440,N_39278);
or U40672 (N_40672,N_39815,N_37851);
nor U40673 (N_40673,N_39484,N_36025);
nand U40674 (N_40674,N_35704,N_37266);
xor U40675 (N_40675,N_35723,N_39420);
nand U40676 (N_40676,N_39597,N_35925);
nor U40677 (N_40677,N_35358,N_37706);
nor U40678 (N_40678,N_38571,N_38734);
nand U40679 (N_40679,N_39527,N_35859);
or U40680 (N_40680,N_38362,N_35162);
and U40681 (N_40681,N_37025,N_35506);
xor U40682 (N_40682,N_39229,N_37673);
nand U40683 (N_40683,N_35411,N_35124);
or U40684 (N_40684,N_35100,N_37011);
nor U40685 (N_40685,N_35216,N_36540);
and U40686 (N_40686,N_37417,N_36880);
nand U40687 (N_40687,N_36495,N_37062);
nand U40688 (N_40688,N_35601,N_35314);
and U40689 (N_40689,N_36570,N_39085);
and U40690 (N_40690,N_38999,N_36712);
and U40691 (N_40691,N_38304,N_36725);
xor U40692 (N_40692,N_35870,N_39606);
nor U40693 (N_40693,N_35399,N_39694);
xor U40694 (N_40694,N_39324,N_36955);
nand U40695 (N_40695,N_38630,N_36509);
xor U40696 (N_40696,N_36122,N_36099);
xnor U40697 (N_40697,N_39309,N_38219);
xor U40698 (N_40698,N_36427,N_39053);
or U40699 (N_40699,N_39030,N_39821);
nor U40700 (N_40700,N_37433,N_35893);
nor U40701 (N_40701,N_38393,N_35412);
xor U40702 (N_40702,N_35549,N_38968);
nand U40703 (N_40703,N_35901,N_37684);
or U40704 (N_40704,N_36944,N_37451);
nor U40705 (N_40705,N_37401,N_35583);
nand U40706 (N_40706,N_38183,N_38515);
and U40707 (N_40707,N_36365,N_38871);
xnor U40708 (N_40708,N_35570,N_38606);
nand U40709 (N_40709,N_38577,N_35632);
and U40710 (N_40710,N_37336,N_38246);
xor U40711 (N_40711,N_36744,N_36778);
or U40712 (N_40712,N_39892,N_36409);
nor U40713 (N_40713,N_38699,N_36965);
nand U40714 (N_40714,N_35596,N_39945);
nor U40715 (N_40715,N_38034,N_37594);
nor U40716 (N_40716,N_35084,N_36438);
or U40717 (N_40717,N_37781,N_36582);
nand U40718 (N_40718,N_36935,N_35657);
and U40719 (N_40719,N_35370,N_35806);
and U40720 (N_40720,N_38158,N_35625);
nor U40721 (N_40721,N_38484,N_39552);
or U40722 (N_40722,N_37902,N_35005);
nand U40723 (N_40723,N_35503,N_35752);
xor U40724 (N_40724,N_35581,N_35962);
xor U40725 (N_40725,N_39190,N_38961);
xnor U40726 (N_40726,N_37293,N_37341);
xnor U40727 (N_40727,N_35983,N_35099);
xnor U40728 (N_40728,N_37807,N_38525);
or U40729 (N_40729,N_36914,N_35929);
or U40730 (N_40730,N_37162,N_35917);
nand U40731 (N_40731,N_36682,N_37131);
nor U40732 (N_40732,N_36256,N_36030);
and U40733 (N_40733,N_38768,N_36535);
or U40734 (N_40734,N_35681,N_39078);
xnor U40735 (N_40735,N_36657,N_36258);
or U40736 (N_40736,N_36412,N_35369);
nor U40737 (N_40737,N_35017,N_36128);
nor U40738 (N_40738,N_35197,N_35019);
xnor U40739 (N_40739,N_39177,N_35742);
or U40740 (N_40740,N_36901,N_37991);
nand U40741 (N_40741,N_37431,N_37922);
nand U40742 (N_40742,N_35665,N_35134);
xnor U40743 (N_40743,N_39244,N_36022);
and U40744 (N_40744,N_38746,N_39725);
nor U40745 (N_40745,N_36765,N_38503);
nor U40746 (N_40746,N_35910,N_37867);
or U40747 (N_40747,N_37907,N_35309);
and U40748 (N_40748,N_39569,N_35048);
xor U40749 (N_40749,N_36988,N_35118);
nand U40750 (N_40750,N_36751,N_37811);
nor U40751 (N_40751,N_37095,N_35007);
or U40752 (N_40752,N_36793,N_39086);
and U40753 (N_40753,N_38511,N_36554);
or U40754 (N_40754,N_35425,N_36598);
or U40755 (N_40755,N_35448,N_38909);
and U40756 (N_40756,N_37795,N_39990);
and U40757 (N_40757,N_35842,N_37605);
or U40758 (N_40758,N_36410,N_39907);
and U40759 (N_40759,N_36655,N_37496);
and U40760 (N_40760,N_36113,N_38816);
and U40761 (N_40761,N_36678,N_36368);
nand U40762 (N_40762,N_39270,N_37413);
xnor U40763 (N_40763,N_39321,N_39697);
xnor U40764 (N_40764,N_39799,N_37834);
xnor U40765 (N_40765,N_37498,N_37394);
and U40766 (N_40766,N_38075,N_35441);
or U40767 (N_40767,N_35722,N_35846);
nor U40768 (N_40768,N_36155,N_39726);
or U40769 (N_40769,N_38387,N_39893);
nor U40770 (N_40770,N_38066,N_35974);
nand U40771 (N_40771,N_37671,N_38892);
or U40772 (N_40772,N_36006,N_35696);
and U40773 (N_40773,N_39363,N_37643);
nor U40774 (N_40774,N_36895,N_38638);
nand U40775 (N_40775,N_37620,N_37845);
or U40776 (N_40776,N_35556,N_36534);
or U40777 (N_40777,N_35063,N_36633);
nand U40778 (N_40778,N_38480,N_38837);
nand U40779 (N_40779,N_39545,N_38976);
and U40780 (N_40780,N_36848,N_35706);
nand U40781 (N_40781,N_35492,N_39698);
and U40782 (N_40782,N_37954,N_39760);
or U40783 (N_40783,N_36426,N_36362);
nor U40784 (N_40784,N_35189,N_36595);
nand U40785 (N_40785,N_39189,N_38146);
nand U40786 (N_40786,N_39720,N_36882);
xnor U40787 (N_40787,N_39305,N_37931);
nand U40788 (N_40788,N_36857,N_37211);
nand U40789 (N_40789,N_35877,N_37911);
nand U40790 (N_40790,N_38628,N_35559);
xor U40791 (N_40791,N_39213,N_39981);
or U40792 (N_40792,N_39398,N_35898);
xor U40793 (N_40793,N_35691,N_36715);
or U40794 (N_40794,N_39775,N_36054);
nand U40795 (N_40795,N_35714,N_39539);
xnor U40796 (N_40796,N_36254,N_38543);
xnor U40797 (N_40797,N_36230,N_36860);
nor U40798 (N_40798,N_38332,N_37418);
or U40799 (N_40799,N_37622,N_38041);
or U40800 (N_40800,N_37490,N_38449);
and U40801 (N_40801,N_35485,N_37264);
nor U40802 (N_40802,N_37709,N_38301);
nand U40803 (N_40803,N_37548,N_38094);
nand U40804 (N_40804,N_37772,N_36187);
xnor U40805 (N_40805,N_36567,N_35209);
nor U40806 (N_40806,N_39014,N_35829);
nor U40807 (N_40807,N_37535,N_38548);
xor U40808 (N_40808,N_39209,N_37051);
and U40809 (N_40809,N_37520,N_35765);
xnor U40810 (N_40810,N_35813,N_36553);
or U40811 (N_40811,N_38715,N_38285);
or U40812 (N_40812,N_38283,N_35160);
and U40813 (N_40813,N_37114,N_35778);
or U40814 (N_40814,N_36470,N_36288);
xor U40815 (N_40815,N_36292,N_36129);
xnor U40816 (N_40816,N_36733,N_35755);
and U40817 (N_40817,N_36261,N_39173);
or U40818 (N_40818,N_38498,N_35032);
nand U40819 (N_40819,N_38069,N_39881);
or U40820 (N_40820,N_38652,N_38802);
or U40821 (N_40821,N_39429,N_37595);
nor U40822 (N_40822,N_39549,N_38755);
or U40823 (N_40823,N_39130,N_39588);
nand U40824 (N_40824,N_36780,N_37397);
nor U40825 (N_40825,N_38729,N_39574);
nand U40826 (N_40826,N_35655,N_38576);
and U40827 (N_40827,N_37983,N_38244);
xor U40828 (N_40828,N_38675,N_36189);
and U40829 (N_40829,N_35036,N_35834);
nand U40830 (N_40830,N_35835,N_37697);
and U40831 (N_40831,N_37540,N_36947);
nand U40832 (N_40832,N_36383,N_38040);
nor U40833 (N_40833,N_35949,N_38954);
and U40834 (N_40834,N_36270,N_36203);
or U40835 (N_40835,N_38350,N_36843);
or U40836 (N_40836,N_38436,N_39211);
nor U40837 (N_40837,N_38723,N_36956);
xor U40838 (N_40838,N_39202,N_37096);
or U40839 (N_40839,N_38490,N_38908);
and U40840 (N_40840,N_37419,N_37416);
and U40841 (N_40841,N_36861,N_35171);
nand U40842 (N_40842,N_39295,N_36478);
and U40843 (N_40843,N_36401,N_37430);
nand U40844 (N_40844,N_35439,N_37491);
or U40845 (N_40845,N_39715,N_39455);
xnor U40846 (N_40846,N_39568,N_37194);
nand U40847 (N_40847,N_38103,N_36157);
xor U40848 (N_40848,N_35931,N_37534);
and U40849 (N_40849,N_36959,N_37578);
nand U40850 (N_40850,N_36658,N_36611);
nor U40851 (N_40851,N_35518,N_39660);
xnor U40852 (N_40852,N_36279,N_39064);
nor U40853 (N_40853,N_39537,N_39137);
xnor U40854 (N_40854,N_35106,N_35744);
and U40855 (N_40855,N_39306,N_37374);
xor U40856 (N_40856,N_37942,N_35338);
or U40857 (N_40857,N_36522,N_38776);
nand U40858 (N_40858,N_38985,N_37512);
and U40859 (N_40859,N_38713,N_39851);
or U40860 (N_40860,N_37677,N_37339);
xor U40861 (N_40861,N_38383,N_36784);
xor U40862 (N_40862,N_35140,N_36983);
nand U40863 (N_40863,N_39989,N_37969);
or U40864 (N_40864,N_35151,N_38366);
nor U40865 (N_40865,N_39390,N_36805);
or U40866 (N_40866,N_38071,N_37665);
or U40867 (N_40867,N_36345,N_37543);
nand U40868 (N_40868,N_38144,N_35572);
nor U40869 (N_40869,N_36740,N_38844);
nor U40870 (N_40870,N_38753,N_38193);
nor U40871 (N_40871,N_38003,N_39334);
xor U40872 (N_40872,N_36894,N_39325);
xor U40873 (N_40873,N_35046,N_39406);
or U40874 (N_40874,N_37763,N_38352);
or U40875 (N_40875,N_36713,N_35764);
xnor U40876 (N_40876,N_39367,N_39940);
or U40877 (N_40877,N_36234,N_37319);
nor U40878 (N_40878,N_38771,N_38881);
or U40879 (N_40879,N_39742,N_35785);
nor U40880 (N_40880,N_38291,N_38512);
nand U40881 (N_40881,N_35070,N_39263);
and U40882 (N_40882,N_37079,N_38133);
and U40883 (N_40883,N_37053,N_38759);
xnor U40884 (N_40884,N_38376,N_36143);
xor U40885 (N_40885,N_35035,N_36041);
nor U40886 (N_40886,N_36154,N_35187);
and U40887 (N_40887,N_36889,N_38582);
nor U40888 (N_40888,N_37434,N_38760);
xor U40889 (N_40889,N_38458,N_36493);
nand U40890 (N_40890,N_35571,N_38825);
xnor U40891 (N_40891,N_35432,N_38785);
nand U40892 (N_40892,N_35682,N_37059);
or U40893 (N_40893,N_36480,N_35022);
xnor U40894 (N_40894,N_39794,N_35905);
nor U40895 (N_40895,N_35450,N_38247);
xor U40896 (N_40896,N_35409,N_36387);
nand U40897 (N_40897,N_38038,N_38092);
and U40898 (N_40898,N_38107,N_35772);
or U40899 (N_40899,N_36703,N_35876);
or U40900 (N_40900,N_36455,N_37796);
xor U40901 (N_40901,N_38674,N_38963);
nand U40902 (N_40902,N_39853,N_37037);
nor U40903 (N_40903,N_35875,N_39477);
nor U40904 (N_40904,N_36585,N_35607);
xor U40905 (N_40905,N_38419,N_39344);
and U40906 (N_40906,N_38062,N_38413);
nor U40907 (N_40907,N_39139,N_36566);
nand U40908 (N_40908,N_38632,N_36443);
and U40909 (N_40909,N_38502,N_36506);
or U40910 (N_40910,N_35334,N_35061);
and U40911 (N_40911,N_38861,N_36847);
and U40912 (N_40912,N_36273,N_36575);
nand U40913 (N_40913,N_39414,N_37812);
nor U40914 (N_40914,N_39916,N_37895);
and U40915 (N_40915,N_35348,N_36339);
and U40916 (N_40916,N_36666,N_39863);
and U40917 (N_40917,N_36244,N_37362);
nand U40918 (N_40918,N_38534,N_35553);
xnor U40919 (N_40919,N_35475,N_36995);
nor U40920 (N_40920,N_37748,N_39379);
nand U40921 (N_40921,N_38610,N_39841);
nand U40922 (N_40922,N_36808,N_37659);
nor U40923 (N_40923,N_39463,N_35590);
nor U40924 (N_40924,N_35034,N_38899);
xnor U40925 (N_40925,N_38645,N_38018);
xnor U40926 (N_40926,N_36823,N_36255);
nor U40927 (N_40927,N_37396,N_39510);
nand U40928 (N_40928,N_38992,N_35202);
xnor U40929 (N_40929,N_35749,N_36674);
or U40930 (N_40930,N_39939,N_38519);
nor U40931 (N_40931,N_38648,N_36417);
nor U40932 (N_40932,N_38993,N_35915);
and U40933 (N_40933,N_35471,N_37751);
and U40934 (N_40934,N_39543,N_38060);
and U40935 (N_40935,N_37163,N_36497);
nor U40936 (N_40936,N_35730,N_39630);
nand U40937 (N_40937,N_39550,N_37466);
or U40938 (N_40938,N_35452,N_39904);
and U40939 (N_40939,N_37026,N_37471);
xor U40940 (N_40940,N_36184,N_37573);
nand U40941 (N_40941,N_38379,N_39567);
xnor U40942 (N_40942,N_39909,N_39654);
nor U40943 (N_40943,N_39107,N_35953);
and U40944 (N_40944,N_39366,N_39300);
xnor U40945 (N_40945,N_38451,N_36527);
xnor U40946 (N_40946,N_35302,N_35938);
nor U40947 (N_40947,N_36476,N_38330);
or U40948 (N_40948,N_39418,N_38265);
nor U40949 (N_40949,N_38664,N_38156);
or U40950 (N_40950,N_38078,N_36779);
and U40951 (N_40951,N_36669,N_38827);
nor U40952 (N_40952,N_36411,N_36002);
or U40953 (N_40953,N_35278,N_39282);
nor U40954 (N_40954,N_37714,N_37141);
xnor U40955 (N_40955,N_39517,N_36352);
and U40956 (N_40956,N_38151,N_36516);
or U40957 (N_40957,N_35072,N_39051);
nand U40958 (N_40958,N_37265,N_37317);
nand U40959 (N_40959,N_38962,N_36042);
xor U40960 (N_40960,N_38198,N_36466);
and U40961 (N_40961,N_37515,N_35515);
and U40962 (N_40962,N_37432,N_37286);
nor U40963 (N_40963,N_39514,N_39526);
nor U40964 (N_40964,N_39182,N_36700);
xnor U40965 (N_40965,N_35770,N_37604);
or U40966 (N_40966,N_36560,N_35091);
and U40967 (N_40967,N_39385,N_35214);
and U40968 (N_40968,N_37791,N_37504);
or U40969 (N_40969,N_39735,N_38680);
nor U40970 (N_40970,N_36584,N_38841);
or U40971 (N_40971,N_37608,N_39685);
or U40972 (N_40972,N_39221,N_37563);
nor U40973 (N_40973,N_38828,N_39943);
nand U40974 (N_40974,N_37108,N_35888);
xnor U40975 (N_40975,N_39669,N_36786);
nor U40976 (N_40976,N_38377,N_35679);
nor U40977 (N_40977,N_39224,N_38820);
nand U40978 (N_40978,N_37255,N_36797);
nor U40979 (N_40979,N_39464,N_37582);
nand U40980 (N_40980,N_39434,N_38378);
nor U40981 (N_40981,N_37078,N_36654);
nor U40982 (N_40982,N_36082,N_35486);
nand U40983 (N_40983,N_37853,N_37174);
nand U40984 (N_40984,N_36624,N_36472);
and U40985 (N_40985,N_39498,N_39811);
and U40986 (N_40986,N_35271,N_36309);
nor U40987 (N_40987,N_39576,N_39983);
and U40988 (N_40988,N_35600,N_37970);
xor U40989 (N_40989,N_38614,N_37527);
nand U40990 (N_40990,N_35470,N_39074);
xor U40991 (N_40991,N_36227,N_36265);
xor U40992 (N_40992,N_39585,N_39978);
nor U40993 (N_40993,N_38572,N_38336);
and U40994 (N_40994,N_39340,N_39453);
and U40995 (N_40995,N_37360,N_37745);
or U40996 (N_40996,N_38862,N_36875);
nand U40997 (N_40997,N_35577,N_39354);
nand U40998 (N_40998,N_38249,N_39927);
xnor U40999 (N_40999,N_39423,N_35109);
xor U41000 (N_41000,N_37296,N_39069);
nor U41001 (N_41001,N_36662,N_39754);
nand U41002 (N_41002,N_39607,N_36626);
xor U41003 (N_41003,N_35533,N_37367);
nand U41004 (N_41004,N_39776,N_39136);
and U41005 (N_41005,N_39880,N_36617);
or U41006 (N_41006,N_36482,N_37721);
nor U41007 (N_41007,N_38916,N_38644);
nor U41008 (N_41008,N_38556,N_36716);
and U41009 (N_41009,N_39832,N_36878);
and U41010 (N_41010,N_35198,N_35143);
and U41011 (N_41011,N_37164,N_39264);
and U41012 (N_41012,N_39280,N_39485);
or U41013 (N_41013,N_35713,N_39952);
xor U41014 (N_41014,N_37818,N_37219);
or U41015 (N_41015,N_36488,N_35720);
xor U41016 (N_41016,N_39806,N_38950);
xor U41017 (N_41017,N_36692,N_38991);
or U41018 (N_41018,N_35808,N_36774);
nand U41019 (N_41019,N_38314,N_36864);
nand U41020 (N_41020,N_36537,N_37663);
xnor U41021 (N_41021,N_37681,N_39766);
nand U41022 (N_41022,N_37288,N_39146);
or U41023 (N_41023,N_36500,N_39253);
and U41024 (N_41024,N_35111,N_35566);
nor U41025 (N_41025,N_36212,N_35361);
or U41026 (N_41026,N_36048,N_38026);
or U41027 (N_41027,N_37157,N_38786);
nand U41028 (N_41028,N_35545,N_37576);
nor U41029 (N_41029,N_38817,N_39217);
or U41030 (N_41030,N_39134,N_39902);
xnor U41031 (N_41031,N_39495,N_35646);
and U41032 (N_41032,N_35422,N_38604);
xnor U41033 (N_41033,N_38194,N_36925);
or U41034 (N_41034,N_38915,N_35120);
and U41035 (N_41035,N_35521,N_39969);
nor U41036 (N_41036,N_39357,N_39446);
nor U41037 (N_41037,N_39577,N_37597);
or U41038 (N_41038,N_37649,N_37423);
and U41039 (N_41039,N_39386,N_37253);
and U41040 (N_41040,N_36473,N_36165);
or U41041 (N_41041,N_35805,N_37929);
and U41042 (N_41042,N_38175,N_37361);
xor U41043 (N_41043,N_36588,N_37815);
xnor U41044 (N_41044,N_38331,N_38721);
nor U41045 (N_41045,N_39586,N_38472);
nand U41046 (N_41046,N_39795,N_38163);
or U41047 (N_41047,N_38568,N_35088);
and U41048 (N_41048,N_37160,N_35299);
nor U41049 (N_41049,N_36660,N_37476);
nor U41050 (N_41050,N_36651,N_38428);
nand U41051 (N_41051,N_38798,N_35238);
nor U41052 (N_41052,N_35943,N_39640);
xor U41053 (N_41053,N_39664,N_36057);
nand U41054 (N_41054,N_35579,N_35393);
and U41055 (N_41055,N_36188,N_37550);
nor U41056 (N_41056,N_38028,N_37470);
and U41057 (N_41057,N_39554,N_35988);
xnor U41058 (N_41058,N_37289,N_36519);
nand U41059 (N_41059,N_39573,N_37111);
or U41060 (N_41060,N_38714,N_37924);
nand U41061 (N_41061,N_39358,N_36224);
xnor U41062 (N_41062,N_37988,N_39251);
nor U41063 (N_41063,N_39490,N_39791);
and U41064 (N_41064,N_39604,N_38381);
and U41065 (N_41065,N_38233,N_39624);
or U41066 (N_41066,N_35748,N_37392);
nor U41067 (N_41067,N_36649,N_39582);
or U41068 (N_41068,N_37753,N_39961);
nand U41069 (N_41069,N_38551,N_36837);
xnor U41070 (N_41070,N_35319,N_38110);
and U41071 (N_41071,N_35675,N_35761);
nor U41072 (N_41072,N_38874,N_35803);
and U41073 (N_41073,N_36218,N_39767);
nand U41074 (N_41074,N_37444,N_35235);
nand U41075 (N_41075,N_35221,N_39088);
or U41076 (N_41076,N_36314,N_39950);
and U41077 (N_41077,N_36781,N_36340);
xor U41078 (N_41078,N_37187,N_38013);
nor U41079 (N_41079,N_35256,N_38494);
or U41080 (N_41080,N_38762,N_36140);
nor U41081 (N_41081,N_35853,N_37656);
nor U41082 (N_41082,N_38136,N_36201);
nor U41083 (N_41083,N_35602,N_39079);
nor U41084 (N_41084,N_38456,N_36970);
and U41085 (N_41085,N_37180,N_37240);
xor U41086 (N_41086,N_38196,N_37139);
xnor U41087 (N_41087,N_39580,N_39518);
nor U41088 (N_41088,N_37247,N_39046);
nand U41089 (N_41089,N_38875,N_36852);
or U41090 (N_41090,N_37315,N_39007);
or U41091 (N_41091,N_36782,N_37905);
nand U41092 (N_41092,N_38944,N_35799);
nand U41093 (N_41093,N_38832,N_36609);
nor U41094 (N_41094,N_38879,N_36978);
nand U41095 (N_41095,N_38493,N_38213);
nor U41096 (N_41096,N_39201,N_38111);
xor U41097 (N_41097,N_36998,N_38487);
or U41098 (N_41098,N_35621,N_36127);
and U41099 (N_41099,N_38784,N_35158);
and U41100 (N_41100,N_37705,N_35597);
and U41101 (N_41101,N_39635,N_39682);
and U41102 (N_41102,N_37651,N_35365);
nand U41103 (N_41103,N_37456,N_36174);
nand U41104 (N_41104,N_35593,N_36601);
and U41105 (N_41105,N_38952,N_39875);
and U41106 (N_41106,N_38089,N_38201);
nand U41107 (N_41107,N_36891,N_36926);
or U41108 (N_41108,N_35286,N_37624);
nor U41109 (N_41109,N_35641,N_39856);
nand U41110 (N_41110,N_37909,N_35587);
nor U41111 (N_41111,N_39283,N_35312);
or U41112 (N_41112,N_39433,N_35639);
and U41113 (N_41113,N_35847,N_37438);
nor U41114 (N_41114,N_36386,N_38724);
or U41115 (N_41115,N_35703,N_39703);
and U41116 (N_41116,N_38948,N_38979);
and U41117 (N_41117,N_36727,N_37769);
nand U41118 (N_41118,N_35268,N_38709);
nor U41119 (N_41119,N_35697,N_37484);
or U41120 (N_41120,N_36007,N_39377);
and U41121 (N_41121,N_37975,N_37995);
and U41122 (N_41122,N_38814,N_39336);
and U41123 (N_41123,N_35737,N_39584);
and U41124 (N_41124,N_36220,N_36870);
nand U41125 (N_41125,N_38054,N_37941);
nor U41126 (N_41126,N_39979,N_36656);
and U41127 (N_41127,N_39538,N_39233);
xnor U41128 (N_41128,N_35274,N_35816);
nand U41129 (N_41129,N_36289,N_38241);
and U41130 (N_41130,N_35630,N_35261);
xnor U41131 (N_41131,N_36971,N_38235);
and U41132 (N_41132,N_36639,N_36979);
or U41133 (N_41133,N_35328,N_39745);
nor U41134 (N_41134,N_35177,N_37178);
nor U41135 (N_41135,N_39638,N_38473);
nand U41136 (N_41136,N_36017,N_35410);
xor U41137 (N_41137,N_39994,N_37136);
nor U41138 (N_41138,N_37517,N_39338);
and U41139 (N_41139,N_38640,N_39272);
nand U41140 (N_41140,N_37837,N_38230);
nand U41141 (N_41141,N_37522,N_35304);
nand U41142 (N_41142,N_38917,N_38139);
or U41143 (N_41143,N_37290,N_35301);
or U41144 (N_41144,N_36459,N_36481);
and U41145 (N_41145,N_39337,N_38889);
nor U41146 (N_41146,N_37783,N_35520);
nor U41147 (N_41147,N_38348,N_38218);
nand U41148 (N_41148,N_37968,N_37061);
xnor U41149 (N_41149,N_35133,N_37767);
nor U41150 (N_41150,N_38643,N_35712);
nand U41151 (N_41151,N_37410,N_38898);
and U41152 (N_41152,N_35965,N_39110);
nand U41153 (N_41153,N_39896,N_38914);
or U41154 (N_41154,N_35959,N_39878);
nand U41155 (N_41155,N_36994,N_35791);
nor U41156 (N_41156,N_39570,N_38380);
nor U41157 (N_41157,N_35743,N_38155);
and U41158 (N_41158,N_37625,N_35336);
and U41159 (N_41159,N_37545,N_37701);
or U41160 (N_41160,N_37116,N_35686);
nor U41161 (N_41161,N_39409,N_38051);
nand U41162 (N_41162,N_37917,N_35264);
nand U41163 (N_41163,N_35424,N_38161);
or U41164 (N_41164,N_36501,N_36471);
or U41165 (N_41165,N_39869,N_39460);
and U41166 (N_41166,N_38360,N_39174);
xnor U41167 (N_41167,N_39541,N_36371);
nor U41168 (N_41168,N_37700,N_37800);
xnor U41169 (N_41169,N_35107,N_36031);
nor U41170 (N_41170,N_35218,N_37645);
or U41171 (N_41171,N_37327,N_38123);
xor U41172 (N_41172,N_37974,N_39304);
xor U41173 (N_41173,N_35627,N_38894);
nor U41174 (N_41174,N_39873,N_39284);
nor U41175 (N_41175,N_36028,N_38274);
and U41176 (N_41176,N_38426,N_38673);
xor U41177 (N_41177,N_37675,N_36225);
nand U41178 (N_41178,N_36530,N_35223);
xnor U41179 (N_41179,N_36491,N_39092);
nand U41180 (N_41180,N_37829,N_35030);
xnor U41181 (N_41181,N_38021,N_39450);
and U41182 (N_41182,N_37650,N_37457);
xnor U41183 (N_41183,N_36297,N_35308);
and U41184 (N_41184,N_35817,N_37206);
xor U41185 (N_41185,N_37885,N_36586);
and U41186 (N_41186,N_35225,N_36525);
xor U41187 (N_41187,N_38154,N_38397);
nand U41188 (N_41188,N_38184,N_37424);
or U41189 (N_41189,N_35129,N_35865);
xnor U41190 (N_41190,N_37884,N_36635);
nor U41191 (N_41191,N_35612,N_38072);
nor U41192 (N_41192,N_39243,N_37282);
nor U41193 (N_41193,N_37731,N_37782);
and U41194 (N_41194,N_39874,N_35346);
nor U41195 (N_41195,N_35539,N_36748);
nor U41196 (N_41196,N_38642,N_36458);
xor U41197 (N_41197,N_36953,N_35821);
nor U41198 (N_41198,N_37324,N_35773);
xnor U41199 (N_41199,N_38660,N_38906);
and U41200 (N_41200,N_37536,N_37479);
xnor U41201 (N_41201,N_38500,N_35444);
nand U41202 (N_41202,N_36974,N_39285);
nor U41203 (N_41203,N_35568,N_37391);
xnor U41204 (N_41204,N_36332,N_39852);
xor U41205 (N_41205,N_36361,N_35927);
nand U41206 (N_41206,N_37124,N_39303);
or U41207 (N_41207,N_35750,N_35465);
xnor U41208 (N_41208,N_35711,N_35104);
nor U41209 (N_41209,N_38858,N_39636);
nand U41210 (N_41210,N_35827,N_37233);
nand U41211 (N_41211,N_39391,N_36023);
and U41212 (N_41212,N_36052,N_39094);
or U41213 (N_41213,N_39792,N_36865);
and U41214 (N_41214,N_38831,N_39246);
and U41215 (N_41215,N_39822,N_35689);
xor U41216 (N_41216,N_38108,N_38164);
nand U41217 (N_41217,N_37295,N_35086);
or U41218 (N_41218,N_38112,N_37355);
xor U41219 (N_41219,N_35224,N_37702);
and U41220 (N_41220,N_38063,N_35896);
or U41221 (N_41221,N_37865,N_37027);
or U41222 (N_41222,N_39556,N_38547);
and U41223 (N_41223,N_37179,N_39613);
and U41224 (N_41224,N_36419,N_37892);
nand U41225 (N_41225,N_38939,N_38058);
nor U41226 (N_41226,N_39955,N_37363);
xnor U41227 (N_41227,N_35792,N_35708);
or U41228 (N_41228,N_37500,N_35103);
or U41229 (N_41229,N_37117,N_36576);
nand U41230 (N_41230,N_35609,N_36316);
and U41231 (N_41231,N_35200,N_38633);
nor U41232 (N_41232,N_37802,N_35473);
nand U41233 (N_41233,N_38395,N_39328);
nand U41234 (N_41234,N_35102,N_39124);
nor U41235 (N_41235,N_38639,N_35013);
nor U41236 (N_41236,N_36286,N_38708);
nor U41237 (N_41237,N_38867,N_37274);
nor U41238 (N_41238,N_36615,N_36242);
or U41239 (N_41239,N_39844,N_35517);
or U41240 (N_41240,N_35347,N_36260);
xor U41241 (N_41241,N_37495,N_36005);
nor U41242 (N_41242,N_37789,N_39860);
and U41243 (N_41243,N_35899,N_39019);
nor U41244 (N_41244,N_39005,N_39138);
nor U41245 (N_41245,N_37069,N_39050);
and U41246 (N_41246,N_37228,N_36856);
nor U41247 (N_41247,N_35952,N_35507);
nor U41248 (N_41248,N_37241,N_35321);
and U41249 (N_41249,N_39919,N_36367);
nor U41250 (N_41250,N_35824,N_39765);
nor U41251 (N_41251,N_35254,N_38940);
nand U41252 (N_41252,N_38957,N_37209);
xnor U41253 (N_41253,N_38005,N_36919);
or U41254 (N_41254,N_36940,N_36623);
nand U41255 (N_41255,N_37013,N_37660);
nand U41256 (N_41256,N_36213,N_35976);
xor U41257 (N_41257,N_39461,N_38850);
xnor U41258 (N_41258,N_39846,N_35871);
nor U41259 (N_41259,N_37695,N_36710);
or U41260 (N_41260,N_36257,N_35638);
or U41261 (N_41261,N_35287,N_35077);
and U41262 (N_41262,N_39117,N_35094);
nand U41263 (N_41263,N_38586,N_39928);
nor U41264 (N_41264,N_36590,N_37038);
nand U41265 (N_41265,N_38935,N_39672);
and U41266 (N_41266,N_38143,N_36816);
xnor U41267 (N_41267,N_38068,N_39871);
nor U41268 (N_41268,N_37329,N_37940);
and U41269 (N_41269,N_36905,N_39601);
or U41270 (N_41270,N_35087,N_39650);
nor U41271 (N_41271,N_39603,N_36382);
nand U41272 (N_41272,N_38297,N_38803);
nor U41273 (N_41273,N_36872,N_39689);
and U41274 (N_41274,N_35083,N_37870);
or U41275 (N_41275,N_38081,N_35377);
xnor U41276 (N_41276,N_37566,N_37071);
xnor U41277 (N_41277,N_35501,N_35994);
nand U41278 (N_41278,N_38188,N_38313);
nor U41279 (N_41279,N_39592,N_36849);
or U41280 (N_41280,N_35186,N_36107);
or U41281 (N_41281,N_36216,N_38953);
and U41282 (N_41282,N_35353,N_35794);
xor U41283 (N_41283,N_37215,N_38686);
nand U41284 (N_41284,N_36697,N_38446);
nand U41285 (N_41285,N_39208,N_38813);
and U41286 (N_41286,N_35233,N_38767);
nor U41287 (N_41287,N_39716,N_38907);
xnor U41288 (N_41288,N_38462,N_35942);
xnor U41289 (N_41289,N_36029,N_35417);
or U41290 (N_41290,N_36513,N_37021);
and U41291 (N_41291,N_35043,N_38468);
or U41292 (N_41292,N_39819,N_35121);
and U41293 (N_41293,N_37323,N_37844);
nor U41294 (N_41294,N_38541,N_39578);
or U41295 (N_41295,N_39403,N_35207);
nor U41296 (N_41296,N_35886,N_35687);
nand U41297 (N_41297,N_39768,N_38637);
or U41298 (N_41298,N_37216,N_39816);
nand U41299 (N_41299,N_38728,N_36883);
nand U41300 (N_41300,N_39011,N_35664);
and U41301 (N_41301,N_37250,N_36873);
or U41302 (N_41302,N_39572,N_36869);
xor U41303 (N_41303,N_37621,N_38033);
or U41304 (N_41304,N_35082,N_37487);
and U41305 (N_41305,N_39038,N_37229);
nand U41306 (N_41306,N_35289,N_37012);
nor U41307 (N_41307,N_35645,N_39643);
nand U41308 (N_41308,N_38483,N_36928);
or U41309 (N_41309,N_37497,N_38186);
or U41310 (N_41310,N_37232,N_37639);
and U41311 (N_41311,N_36198,N_38995);
nand U41312 (N_41312,N_37001,N_39252);
xor U41313 (N_41313,N_37311,N_37377);
xnor U41314 (N_41314,N_38008,N_35089);
nor U41315 (N_41315,N_39185,N_35136);
nand U41316 (N_41316,N_35498,N_39350);
nand U41317 (N_41317,N_36000,N_38167);
nand U41318 (N_41318,N_37506,N_37814);
and U41319 (N_41319,N_35310,N_36308);
xor U41320 (N_41320,N_35650,N_39662);
or U41321 (N_41321,N_36414,N_37112);
xnor U41322 (N_41322,N_37518,N_37730);
or U41323 (N_41323,N_39153,N_39954);
nand U41324 (N_41324,N_36967,N_38466);
nor U41325 (N_41325,N_39511,N_39800);
nor U41326 (N_41326,N_39269,N_36027);
or U41327 (N_41327,N_37601,N_36591);
or U41328 (N_41328,N_39532,N_36951);
nand U41329 (N_41329,N_37049,N_36271);
nand U41330 (N_41330,N_38750,N_36858);
nor U41331 (N_41331,N_36064,N_39802);
xor U41332 (N_41332,N_38905,N_39220);
nor U41333 (N_41333,N_38137,N_36677);
xnor U41334 (N_41334,N_37819,N_36284);
nand U41335 (N_41335,N_39491,N_39353);
and U41336 (N_41336,N_38608,N_37872);
or U41337 (N_41337,N_35241,N_38237);
and U41338 (N_41338,N_37008,N_37984);
and U41339 (N_41339,N_39929,N_37406);
xnor U41340 (N_41340,N_38372,N_39583);
nand U41341 (N_41341,N_35984,N_37104);
nor U41342 (N_41342,N_36942,N_37275);
nor U41343 (N_41343,N_38611,N_37110);
or U41344 (N_41344,N_37138,N_35825);
nand U41345 (N_41345,N_35317,N_36578);
nand U41346 (N_41346,N_39279,N_37269);
nand U41347 (N_41347,N_39717,N_37244);
nand U41348 (N_41348,N_36032,N_37054);
and U41349 (N_41349,N_37586,N_39899);
xnor U41350 (N_41350,N_37208,N_39172);
and U41351 (N_41351,N_38211,N_35709);
or U41352 (N_41352,N_35908,N_38599);
xnor U41353 (N_41353,N_37085,N_39438);
or U41354 (N_41354,N_39833,N_35578);
and U41355 (N_41355,N_38826,N_37441);
xor U41356 (N_41356,N_36243,N_35128);
or U41357 (N_41357,N_35733,N_38020);
or U41358 (N_41358,N_37935,N_39302);
nor U41359 (N_41359,N_39938,N_36711);
xor U41360 (N_41360,N_39169,N_36055);
and U41361 (N_41361,N_38001,N_38978);
xnor U41362 (N_41362,N_36281,N_37172);
nor U41363 (N_41363,N_37338,N_37272);
and U41364 (N_41364,N_37927,N_35058);
or U41365 (N_41365,N_35837,N_39184);
or U41366 (N_41366,N_39787,N_39062);
or U41367 (N_41367,N_38179,N_37127);
nor U41368 (N_41368,N_37644,N_38884);
nor U41369 (N_41369,N_37221,N_37636);
or U41370 (N_41370,N_35666,N_38847);
nand U41371 (N_41371,N_37494,N_38176);
nand U41372 (N_41372,N_38849,N_35598);
nor U41373 (N_41373,N_36429,N_38394);
nand U41374 (N_41374,N_35883,N_39231);
and U41375 (N_41375,N_39440,N_38670);
or U41376 (N_41376,N_39782,N_39276);
nand U41377 (N_41377,N_35633,N_37944);
nand U41378 (N_41378,N_35766,N_38354);
and U41379 (N_41379,N_36373,N_39361);
nand U41380 (N_41380,N_38489,N_37546);
nor U41381 (N_41381,N_36026,N_35391);
xnor U41382 (N_41382,N_37335,N_39663);
nand U41383 (N_41383,N_39718,N_35840);
or U41384 (N_41384,N_38270,N_36178);
nand U41385 (N_41385,N_35776,N_38830);
and U41386 (N_41386,N_35828,N_39192);
xor U41387 (N_41387,N_36044,N_38273);
nor U41388 (N_41388,N_38410,N_37400);
nand U41389 (N_41389,N_36091,N_38056);
and U41390 (N_41390,N_37823,N_39310);
or U41391 (N_41391,N_35535,N_39333);
and U41392 (N_41392,N_39711,N_39910);
nand U41393 (N_41393,N_36280,N_38082);
xnor U41394 (N_41394,N_37002,N_38990);
or U41395 (N_41395,N_38272,N_39897);
nand U41396 (N_41396,N_35930,N_35672);
nand U41397 (N_41397,N_39474,N_39486);
nor U41398 (N_41398,N_35928,N_38617);
and U41399 (N_41399,N_36915,N_38243);
nand U41400 (N_41400,N_35462,N_39487);
and U41401 (N_41401,N_36103,N_35097);
or U41402 (N_41402,N_37507,N_38730);
nor U41403 (N_41403,N_35344,N_37488);
nor U41404 (N_41404,N_35434,N_37277);
nand U41405 (N_41405,N_35801,N_36268);
nand U41406 (N_41406,N_39193,N_35941);
or U41407 (N_41407,N_38307,N_38824);
xnor U41408 (N_41408,N_37920,N_35526);
nand U41409 (N_41409,N_37066,N_37132);
or U41410 (N_41410,N_39158,N_37318);
or U41411 (N_41411,N_36247,N_38938);
nand U41412 (N_41412,N_39378,N_37722);
nor U41413 (N_41413,N_35320,N_37382);
xnor U41414 (N_41414,N_37775,N_35987);
and U41415 (N_41415,N_39895,N_37473);
or U41416 (N_41416,N_39045,N_35855);
and U41417 (N_41417,N_38284,N_39661);
and U41418 (N_41418,N_36918,N_37015);
xor U41419 (N_41419,N_35489,N_35966);
xnor U41420 (N_41420,N_39676,N_36109);
and U41421 (N_41421,N_35637,N_38295);
nor U41422 (N_41422,N_39115,N_37168);
nor U41423 (N_41423,N_37231,N_35067);
and U41424 (N_41424,N_38965,N_37412);
nor U41425 (N_41425,N_38926,N_38891);
or U41426 (N_41426,N_36372,N_38757);
nor U41427 (N_41427,N_37508,N_36376);
nand U41428 (N_41428,N_39068,N_35540);
nand U41429 (N_41429,N_35460,N_36610);
and U41430 (N_41430,N_36704,N_39963);
nor U41431 (N_41431,N_35924,N_37197);
nor U41432 (N_41432,N_36921,N_37863);
or U41433 (N_41433,N_39752,N_37755);
nor U41434 (N_41434,N_38781,N_38738);
or U41435 (N_41435,N_37186,N_37285);
or U41436 (N_41436,N_37669,N_38023);
nand U41437 (N_41437,N_36015,N_36749);
xor U41438 (N_41438,N_39563,N_37632);
and U41439 (N_41439,N_38811,N_35195);
nand U41440 (N_41440,N_38559,N_37951);
nor U41441 (N_41441,N_37478,N_35710);
nand U41442 (N_41442,N_35537,N_38135);
nand U41443 (N_41443,N_38684,N_37549);
nand U41444 (N_41444,N_38453,N_35085);
nand U41445 (N_41445,N_36903,N_38696);
and U41446 (N_41446,N_38438,N_38780);
nor U41447 (N_41447,N_35112,N_39524);
xnor U41448 (N_41448,N_38987,N_35982);
nand U41449 (N_41449,N_39261,N_36343);
or U41450 (N_41450,N_38070,N_37910);
xor U41451 (N_41451,N_37542,N_36759);
xor U41452 (N_41452,N_36325,N_39504);
or U41453 (N_41453,N_35011,N_39291);
nand U41454 (N_41454,N_36452,N_35531);
xor U41455 (N_41455,N_36033,N_36879);
or U41456 (N_41456,N_35977,N_36505);
and U41457 (N_41457,N_39724,N_36487);
and U41458 (N_41458,N_39021,N_35809);
nand U41459 (N_41459,N_39106,N_35389);
and U41460 (N_41460,N_36240,N_36804);
xnor U41461 (N_41461,N_37261,N_39167);
nor U41462 (N_41462,N_38666,N_39327);
nand U41463 (N_41463,N_36347,N_37640);
nor U41464 (N_41464,N_36699,N_38566);
nand U41465 (N_41465,N_35629,N_35933);
or U41466 (N_41466,N_38722,N_39388);
nor U41467 (N_41467,N_38840,N_35155);
and U41468 (N_41468,N_38537,N_35033);
and U41469 (N_41469,N_36806,N_37569);
and U41470 (N_41470,N_35738,N_38569);
nor U41471 (N_41471,N_39596,N_39706);
or U41472 (N_41472,N_36016,N_36034);
or U41473 (N_41473,N_35656,N_35787);
nand U41474 (N_41474,N_38460,N_35078);
or U41475 (N_41475,N_37452,N_37063);
nand U41476 (N_41476,N_38011,N_38463);
xor U41477 (N_41477,N_39175,N_35882);
nor U41478 (N_41478,N_35038,N_38171);
or U41479 (N_41479,N_39228,N_37897);
xnor U41480 (N_41480,N_39383,N_36375);
nand U41481 (N_41481,N_38138,N_39962);
and U41482 (N_41482,N_38538,N_38342);
and U41483 (N_41483,N_36071,N_39292);
or U41484 (N_41484,N_39542,N_39008);
or U41485 (N_41485,N_37626,N_39168);
and U41486 (N_41486,N_35420,N_38929);
and U41487 (N_41487,N_35562,N_37784);
nor U41488 (N_41488,N_35740,N_35892);
nand U41489 (N_41489,N_39622,N_39442);
nand U41490 (N_41490,N_38717,N_36841);
nor U41491 (N_41491,N_36938,N_38074);
xnor U41492 (N_41492,N_35295,N_35127);
nor U41493 (N_41493,N_35700,N_39080);
nor U41494 (N_41494,N_38705,N_38185);
nor U41495 (N_41495,N_37912,N_38712);
or U41496 (N_41496,N_38996,N_38620);
nand U41497 (N_41497,N_35868,N_39250);
or U41498 (N_41498,N_36275,N_36827);
nand U41499 (N_41499,N_38061,N_36763);
and U41500 (N_41500,N_36301,N_38113);
xor U41501 (N_41501,N_37746,N_37093);
and U41502 (N_41502,N_39855,N_38791);
nor U41503 (N_41503,N_36479,N_35523);
and U41504 (N_41504,N_38322,N_35586);
xnor U41505 (N_41505,N_38973,N_36997);
nor U41506 (N_41506,N_38619,N_37777);
nor U41507 (N_41507,N_39362,N_39161);
and U41508 (N_41508,N_37439,N_38099);
and U41509 (N_41509,N_35281,N_39089);
and U41510 (N_41510,N_37235,N_38102);
or U41511 (N_41511,N_39528,N_37537);
or U41512 (N_41512,N_39547,N_38758);
or U41513 (N_41513,N_35021,N_36089);
and U41514 (N_41514,N_39479,N_37328);
nor U41515 (N_41515,N_36451,N_36966);
nor U41516 (N_41516,N_38918,N_39684);
or U41517 (N_41517,N_39761,N_36133);
xnor U41518 (N_41518,N_39214,N_36788);
or U41519 (N_41519,N_39393,N_39553);
nand U41520 (N_41520,N_39198,N_38365);
or U41521 (N_41521,N_37976,N_35529);
nand U41522 (N_41522,N_38145,N_38217);
xor U41523 (N_41523,N_35025,N_38049);
or U41524 (N_41524,N_39318,N_36868);
nand U41525 (N_41525,N_36333,N_36223);
or U41526 (N_41526,N_35404,N_35315);
nor U41527 (N_41527,N_36020,N_38289);
or U41528 (N_41528,N_35811,N_38671);
nor U41529 (N_41529,N_35798,N_35006);
nand U41530 (N_41530,N_37592,N_36802);
or U41531 (N_41531,N_38305,N_36850);
and U41532 (N_41532,N_39646,N_35760);
xor U41533 (N_41533,N_36840,N_39670);
and U41534 (N_41534,N_36418,N_35105);
nand U41535 (N_41535,N_35018,N_36547);
and U41536 (N_41536,N_35980,N_36767);
or U41537 (N_41537,N_37736,N_36130);
nor U41538 (N_41538,N_38407,N_36310);
or U41539 (N_41539,N_35753,N_35872);
xnor U41540 (N_41540,N_39671,N_36415);
and U41541 (N_41541,N_38821,N_35918);
nor U41542 (N_41542,N_38597,N_35354);
or U41543 (N_41543,N_38868,N_39238);
xnor U41544 (N_41544,N_35921,N_38594);
nand U41545 (N_41545,N_35826,N_37133);
or U41546 (N_41546,N_39710,N_39489);
and U41547 (N_41547,N_36829,N_36266);
nor U41548 (N_41548,N_36330,N_39425);
nand U41549 (N_41549,N_36707,N_36688);
xor U41550 (N_41550,N_37190,N_35576);
xnor U41551 (N_41551,N_35045,N_35631);
and U41552 (N_41552,N_39205,N_36798);
nor U41553 (N_41553,N_37567,N_35051);
or U41554 (N_41554,N_36388,N_35108);
xor U41555 (N_41555,N_37839,N_35298);
and U41556 (N_41556,N_39401,N_37692);
nand U41557 (N_41557,N_37617,N_39149);
and U41558 (N_41558,N_39788,N_36160);
nor U41559 (N_41559,N_39830,N_37436);
nor U41560 (N_41560,N_35205,N_36772);
nor U41561 (N_41561,N_39212,N_37200);
nor U41562 (N_41562,N_39723,N_37688);
nand U41563 (N_41563,N_37754,N_35416);
nand U41564 (N_41564,N_39618,N_36076);
nor U41565 (N_41565,N_38732,N_37864);
nand U41566 (N_41566,N_38690,N_35864);
and U41567 (N_41567,N_36670,N_36474);
xnor U41568 (N_41568,N_36461,N_37042);
or U41569 (N_41569,N_37149,N_37803);
xnor U41570 (N_41570,N_37718,N_39002);
nor U41571 (N_41571,N_35784,N_39476);
nand U41572 (N_41572,N_37887,N_39868);
nand U41573 (N_41573,N_36836,N_39623);
and U41574 (N_41574,N_36981,N_37571);
or U41575 (N_41575,N_35690,N_35881);
xnor U41576 (N_41576,N_35969,N_39817);
nor U41577 (N_41577,N_37020,N_38347);
xnor U41578 (N_41578,N_39750,N_39625);
xor U41579 (N_41579,N_37303,N_39268);
or U41580 (N_41580,N_39102,N_37113);
nand U41581 (N_41581,N_37634,N_37158);
or U41582 (N_41582,N_37306,N_36597);
and U41583 (N_41583,N_37128,N_36389);
or U41584 (N_41584,N_37557,N_37934);
xnor U41585 (N_41585,N_39858,N_39308);
nor U41586 (N_41586,N_35330,N_36887);
xor U41587 (N_41587,N_39701,N_35401);
or U41588 (N_41588,N_36151,N_38245);
xnor U41589 (N_41589,N_39234,N_38126);
nand U41590 (N_41590,N_36045,N_35313);
nor U41591 (N_41591,N_35754,N_37302);
or U41592 (N_41592,N_39275,N_39405);
nor U41593 (N_41593,N_35182,N_36668);
nand U41594 (N_41594,N_36842,N_35373);
and U41595 (N_41595,N_35769,N_35560);
or U41596 (N_41596,N_36731,N_38344);
xor U41597 (N_41597,N_38859,N_39456);
nor U41598 (N_41598,N_38937,N_39829);
or U41599 (N_41599,N_39926,N_37376);
nand U41600 (N_41600,N_38562,N_35777);
nor U41601 (N_41601,N_35275,N_39772);
or U41602 (N_41602,N_37616,N_37757);
xor U41603 (N_41603,N_36906,N_35698);
or U41604 (N_41604,N_36287,N_35239);
nor U41605 (N_41605,N_39707,N_38887);
xnor U41606 (N_41606,N_38930,N_38737);
nor U41607 (N_41607,N_35478,N_37313);
nand U41608 (N_41608,N_35440,N_39632);
or U41609 (N_41609,N_39513,N_38302);
nor U41610 (N_41610,N_37379,N_38229);
or U41611 (N_41611,N_38259,N_36571);
nand U41612 (N_41612,N_37227,N_37072);
nand U41613 (N_41613,N_38585,N_38264);
xnor U41614 (N_41614,N_35474,N_38340);
xor U41615 (N_41615,N_39374,N_35031);
or U41616 (N_41616,N_39521,N_38612);
or U41617 (N_41617,N_35487,N_39677);
and U41618 (N_41618,N_35266,N_36730);
xnor U41619 (N_41619,N_37387,N_39176);
nor U41620 (N_41620,N_38491,N_36604);
or U41621 (N_41621,N_39758,N_35500);
nand U41622 (N_41622,N_39431,N_39277);
nand U41623 (N_41623,N_37732,N_37381);
nor U41624 (N_41624,N_36976,N_37816);
or U41625 (N_41625,N_37679,N_36702);
nand U41626 (N_41626,N_39629,N_35508);
nor U41627 (N_41627,N_37652,N_39756);
nand U41628 (N_41628,N_39341,N_38540);
xnor U41629 (N_41629,N_35838,N_37214);
and U41630 (N_41630,N_39227,N_39382);
and U41631 (N_41631,N_35243,N_36217);
or U41632 (N_41632,N_38404,N_36982);
and U41633 (N_41633,N_37171,N_39627);
or U41634 (N_41634,N_36933,N_39032);
or U41635 (N_41635,N_38117,N_37945);
nand U41636 (N_41636,N_36757,N_39114);
and U41637 (N_41637,N_39020,N_37584);
nor U41638 (N_41638,N_39034,N_37890);
xnor U41639 (N_41639,N_37530,N_39090);
nand U41640 (N_41640,N_36747,N_36175);
xor U41641 (N_41641,N_35096,N_35623);
or U41642 (N_41642,N_35735,N_38677);
nor U41643 (N_41643,N_39352,N_35575);
nor U41644 (N_41644,N_39831,N_37028);
xor U41645 (N_41645,N_37185,N_35483);
or U41646 (N_41646,N_36075,N_38406);
nor U41647 (N_41647,N_39728,N_38865);
and U41648 (N_41648,N_36353,N_35774);
nand U41649 (N_41649,N_36391,N_38676);
or U41650 (N_41650,N_36652,N_37357);
xor U41651 (N_41651,N_36061,N_37056);
or U41652 (N_41652,N_38349,N_36706);
nor U41653 (N_41653,N_37402,N_35734);
nor U41654 (N_41654,N_37393,N_38923);
and U41655 (N_41655,N_36051,N_36900);
and U41656 (N_41656,N_36423,N_36344);
and U41657 (N_41657,N_36049,N_39993);
nor U41658 (N_41658,N_36341,N_38641);
nor U41659 (N_41659,N_39256,N_36214);
xnor U41660 (N_41660,N_39096,N_35874);
or U41661 (N_41661,N_39010,N_35880);
or U41662 (N_41662,N_38339,N_36322);
xor U41663 (N_41663,N_37153,N_38745);
or U41664 (N_41664,N_37481,N_38656);
or U41665 (N_41665,N_36687,N_37345);
nor U41666 (N_41666,N_36236,N_35343);
nand U41667 (N_41667,N_38810,N_39360);
nand U41668 (N_41668,N_35557,N_36138);
nor U41669 (N_41669,N_36408,N_35429);
and U41670 (N_41670,N_35986,N_35426);
or U41671 (N_41671,N_36021,N_39837);
nand U41672 (N_41672,N_37222,N_37686);
nand U41673 (N_41673,N_36621,N_39649);
nand U41674 (N_41674,N_38531,N_36235);
and U41675 (N_41675,N_37249,N_38437);
xnor U41676 (N_41676,N_37039,N_36685);
nand U41677 (N_41677,N_39194,N_38565);
nand U41678 (N_41678,N_38651,N_36038);
xnor U41679 (N_41679,N_35383,N_37404);
and U41680 (N_41680,N_36306,N_39315);
nand U41681 (N_41681,N_36787,N_38782);
xor U41682 (N_41682,N_39797,N_36179);
xor U41683 (N_41683,N_35208,N_36701);
nand U41684 (N_41684,N_38479,N_35131);
xor U41685 (N_41685,N_37958,N_39232);
nor U41686 (N_41686,N_39988,N_38593);
or U41687 (N_41687,N_37553,N_37348);
nor U41688 (N_41688,N_39047,N_38357);
nand U41689 (N_41689,N_35340,N_38415);
and U41690 (N_41690,N_37635,N_36964);
and U41691 (N_41691,N_37787,N_37603);
nor U41692 (N_41692,N_36559,N_36358);
or U41693 (N_41693,N_35220,N_37408);
nand U41694 (N_41694,N_38870,N_39631);
nor U41695 (N_41695,N_36785,N_35169);
and U41696 (N_41696,N_39459,N_36640);
and U41697 (N_41697,N_35628,N_39827);
and U41698 (N_41698,N_37173,N_35463);
nor U41699 (N_41699,N_36876,N_36627);
nand U41700 (N_41700,N_39959,N_39779);
xor U41701 (N_41701,N_35296,N_39777);
xnor U41702 (N_41702,N_38860,N_39015);
nand U41703 (N_41703,N_35858,N_35950);
and U41704 (N_41704,N_35614,N_37472);
or U41705 (N_41705,N_39727,N_38382);
and U41706 (N_41706,N_38044,N_36366);
and U41707 (N_41707,N_38267,N_35702);
nor U41708 (N_41708,N_37682,N_38240);
xor U41709 (N_41709,N_36512,N_36498);
xnor U41710 (N_41710,N_39448,N_38046);
or U41711 (N_41711,N_39428,N_38740);
or U41712 (N_41712,N_38662,N_36142);
nand U41713 (N_41713,N_37696,N_39036);
nor U41714 (N_41714,N_35381,N_36489);
nor U41715 (N_41715,N_37252,N_38471);
xnor U41716 (N_41716,N_37395,N_39444);
nor U41717 (N_41717,N_38726,N_37356);
nor U41718 (N_41718,N_36468,N_35453);
or U41719 (N_41719,N_35937,N_39734);
and U41720 (N_41720,N_37847,N_38422);
nor U41721 (N_41721,N_36795,N_38282);
xnor U41722 (N_41722,N_35861,N_35573);
nand U41723 (N_41723,N_37886,N_35616);
nand U41724 (N_41724,N_38650,N_38250);
nor U41725 (N_41725,N_38409,N_38398);
nor U41726 (N_41726,N_37403,N_37994);
or U41727 (N_41727,N_38731,N_37100);
nor U41728 (N_41728,N_38122,N_38324);
xor U41729 (N_41729,N_37607,N_38010);
nand U41730 (N_41730,N_38455,N_37683);
or U41731 (N_41731,N_35757,N_35405);
xor U41732 (N_41732,N_37058,N_38047);
nor U41733 (N_41733,N_35863,N_35716);
and U41734 (N_41734,N_36483,N_38716);
nor U41735 (N_41735,N_38431,N_38345);
nand U41736 (N_41736,N_39505,N_39854);
xnor U41737 (N_41737,N_36008,N_38809);
or U41738 (N_41738,N_38977,N_37017);
xor U41739 (N_41739,N_35653,N_39713);
and U41740 (N_41740,N_37102,N_38550);
or U41741 (N_41741,N_36171,N_35954);
and U41742 (N_41742,N_37477,N_37658);
nand U41743 (N_41743,N_36467,N_35661);
nor U41744 (N_41744,N_38080,N_38994);
or U41745 (N_41745,N_35400,N_36943);
nor U41746 (N_41746,N_36040,N_36817);
nand U41747 (N_41747,N_39840,N_38016);
xor U41748 (N_41748,N_37869,N_38367);
xnor U41749 (N_41749,N_36653,N_36634);
nor U41750 (N_41750,N_39958,N_37615);
nor U41751 (N_41751,N_36238,N_39824);
nor U41752 (N_41752,N_39426,N_36755);
nor U41753 (N_41753,N_38931,N_36147);
nand U41754 (N_41754,N_36397,N_36813);
nand U41755 (N_41755,N_37300,N_35237);
and U41756 (N_41756,N_35530,N_36818);
nand U41757 (N_41757,N_38333,N_39135);
and U41758 (N_41758,N_39976,N_38751);
or U41759 (N_41759,N_39346,N_38327);
and U41760 (N_41760,N_37268,N_37735);
or U41761 (N_41761,N_37513,N_36207);
xnor U41762 (N_41762,N_35849,N_35845);
xor U41763 (N_41763,N_38252,N_36648);
nand U41764 (N_41764,N_37973,N_38492);
and U41765 (N_41765,N_37840,N_35180);
xnor U41766 (N_41766,N_37760,N_36269);
and U41767 (N_41767,N_35258,N_37251);
xnor U41768 (N_41768,N_38869,N_37903);
nand U41769 (N_41769,N_36425,N_39049);
and U41770 (N_41770,N_36705,N_36696);
xnor U41771 (N_41771,N_35265,N_37771);
xnor U41772 (N_41772,N_38654,N_38053);
xnor U41773 (N_41773,N_38989,N_35333);
nand U41774 (N_41774,N_39731,N_39219);
nor U41775 (N_41775,N_35074,N_35459);
or U41776 (N_41776,N_39679,N_38261);
or U41777 (N_41777,N_38162,N_35059);
xnor U41778 (N_41778,N_36019,N_38408);
and U41779 (N_41779,N_38564,N_36508);
and U41780 (N_41780,N_35484,N_37142);
nor U41781 (N_41781,N_38789,N_39492);
xnor U41782 (N_41782,N_38130,N_35234);
nor U41783 (N_41783,N_38893,N_36116);
and U41784 (N_41784,N_37618,N_39121);
nand U41785 (N_41785,N_35359,N_37947);
nand U41786 (N_41786,N_36620,N_37369);
xor U41787 (N_41787,N_37453,N_37283);
xor U41788 (N_41788,N_38035,N_39914);
nor U41789 (N_41789,N_35447,N_36549);
nand U41790 (N_41790,N_36760,N_36413);
nand U41791 (N_41791,N_38306,N_39417);
nor U41792 (N_41792,N_39608,N_38806);
xor U41793 (N_41793,N_36726,N_38920);
nand U41794 (N_41794,N_39447,N_35066);
and U41795 (N_41795,N_39564,N_37101);
or U41796 (N_41796,N_39633,N_38315);
and U41797 (N_41797,N_38695,N_36851);
xor U41798 (N_41798,N_35636,N_35455);
and U41799 (N_41799,N_38403,N_35146);
and U41800 (N_41800,N_37933,N_38700);
and U41801 (N_41801,N_36252,N_39329);
and U41802 (N_41802,N_35550,N_37898);
and U41803 (N_41803,N_37146,N_38605);
nand U41804 (N_41804,N_35076,N_38076);
or U41805 (N_41805,N_37067,N_38741);
xor U41806 (N_41806,N_37981,N_36039);
and U41807 (N_41807,N_36058,N_39104);
and U41808 (N_41808,N_36428,N_36074);
nand U41809 (N_41809,N_39748,N_38852);
and U41810 (N_41810,N_36641,N_36181);
nor U41811 (N_41811,N_37950,N_37109);
nand U41812 (N_41812,N_37900,N_38913);
nor U41813 (N_41813,N_36665,N_35316);
nand U41814 (N_41814,N_39226,N_37443);
or U41815 (N_41815,N_36393,N_36448);
nor U41816 (N_41816,N_35469,N_36152);
nor U41817 (N_41817,N_39084,N_39559);
or U41818 (N_41818,N_35123,N_37262);
and U41819 (N_41819,N_38804,N_38877);
nand U41820 (N_41820,N_38779,N_39462);
or U41821 (N_41821,N_37446,N_36135);
xnor U41822 (N_41822,N_37858,N_37301);
or U41823 (N_41823,N_37525,N_36737);
nor U41824 (N_41824,N_37346,N_38298);
nor U41825 (N_41825,N_36070,N_38848);
or U41826 (N_41826,N_36589,N_37788);
or U41827 (N_41827,N_38227,N_39762);
nand U41828 (N_41828,N_39862,N_36550);
and U41829 (N_41829,N_38678,N_38749);
nor U41830 (N_41830,N_38602,N_36910);
nand U41831 (N_41831,N_38050,N_37879);
xor U41832 (N_41832,N_39614,N_39508);
nor U41833 (N_41833,N_35647,N_38206);
nor U41834 (N_41834,N_36565,N_36486);
and U41835 (N_41835,N_39749,N_37371);
or U41836 (N_41836,N_37672,N_38464);
and U41837 (N_41837,N_35213,N_36233);
xor U41838 (N_41838,N_38337,N_39941);
nor U41839 (N_41839,N_36564,N_38769);
or U41840 (N_41840,N_36485,N_37280);
nand U41841 (N_41841,N_38583,N_35527);
nor U41842 (N_41842,N_37033,N_35245);
nor U41843 (N_41843,N_39686,N_35093);
or U41844 (N_41844,N_36616,N_35080);
nor U41845 (N_41845,N_39349,N_37538);
xnor U41846 (N_41846,N_35936,N_37464);
or U41847 (N_41847,N_36180,N_35215);
or U41848 (N_41848,N_39499,N_38325);
nor U41849 (N_41849,N_35873,N_38956);
and U41850 (N_41850,N_37744,N_35768);
nor U41851 (N_41851,N_35589,N_35288);
nor U41852 (N_41852,N_37083,N_37998);
and U41853 (N_41853,N_35671,N_35408);
or U41854 (N_41854,N_39200,N_35528);
or U41855 (N_41855,N_39095,N_39343);
nor U41856 (N_41856,N_37467,N_38499);
and U41857 (N_41857,N_37729,N_36477);
and U41858 (N_41858,N_37523,N_36078);
or U41859 (N_41859,N_35884,N_35932);
and U41860 (N_41860,N_35869,N_35956);
nand U41861 (N_41861,N_37739,N_39183);
and U41862 (N_41862,N_36924,N_35119);
nand U41863 (N_41863,N_35293,N_35995);
nor U41864 (N_41864,N_38174,N_36724);
nand U41865 (N_41865,N_36518,N_36206);
nand U41866 (N_41866,N_39048,N_38903);
xnor U41867 (N_41867,N_35236,N_35193);
nor U41868 (N_41868,N_38853,N_36437);
or U41869 (N_41869,N_36980,N_36185);
nor U41870 (N_41870,N_39997,N_37084);
xnor U41871 (N_41871,N_39770,N_35211);
xor U41872 (N_41872,N_36276,N_38271);
nand U41873 (N_41873,N_39307,N_36874);
xnor U41874 (N_41874,N_36832,N_38000);
nor U41875 (N_41875,N_37461,N_37150);
nand U41876 (N_41876,N_35967,N_36532);
xor U41877 (N_41877,N_37041,N_38665);
or U41878 (N_41878,N_36789,N_38509);
nor U41879 (N_41879,N_36815,N_38359);
and U41880 (N_41880,N_38857,N_37978);
or U41881 (N_41881,N_36619,N_37685);
or U41882 (N_41882,N_39298,N_36686);
or U41883 (N_41883,N_37939,N_36835);
or U41884 (N_41884,N_36435,N_38873);
xor U41885 (N_41885,N_39012,N_38470);
xnor U41886 (N_41886,N_38933,N_38452);
nand U41887 (N_41887,N_36954,N_39113);
and U41888 (N_41888,N_35844,N_38440);
nand U41889 (N_41889,N_39160,N_39780);
nand U41890 (N_41890,N_39348,N_35654);
nand U41891 (N_41891,N_37690,N_38647);
nand U41892 (N_41892,N_36190,N_39946);
nand U41893 (N_41893,N_36272,N_36568);
xnor U41894 (N_41894,N_35909,N_38743);
nor U41895 (N_41895,N_38580,N_38863);
xor U41896 (N_41896,N_35260,N_39072);
xnor U41897 (N_41897,N_36722,N_35396);
nor U41898 (N_41898,N_37765,N_39519);
or U41899 (N_41899,N_39674,N_35705);
xor U41900 (N_41900,N_39296,N_36327);
nand U41901 (N_41901,N_39240,N_36728);
and U41902 (N_41902,N_35519,N_36139);
nor U41903 (N_41903,N_39562,N_35841);
and U41904 (N_41904,N_37780,N_38549);
and U41905 (N_41905,N_36420,N_36282);
or U41906 (N_41906,N_35595,N_38623);
nand U41907 (N_41907,N_37646,N_36820);
nand U41908 (N_41908,N_36088,N_39733);
or U41909 (N_41909,N_35727,N_37606);
nor U41910 (N_41910,N_38269,N_39805);
nand U41911 (N_41911,N_36695,N_37952);
nor U41912 (N_41912,N_39116,N_39668);
or U41913 (N_41913,N_39235,N_36446);
nor U41914 (N_41914,N_39512,N_35355);
nand U41915 (N_41915,N_36193,N_37960);
and U41916 (N_41916,N_39506,N_39342);
nand U41917 (N_41917,N_37140,N_38800);
or U41918 (N_41918,N_38127,N_37304);
nor U41919 (N_41919,N_35807,N_38388);
and U41920 (N_41920,N_39828,N_36202);
and U41921 (N_41921,N_36563,N_39687);
and U41922 (N_41922,N_35203,N_35398);
nand U41923 (N_41923,N_37713,N_39655);
or U41924 (N_41924,N_37899,N_36521);
xnor U41925 (N_41925,N_38625,N_35159);
nand U41926 (N_41926,N_39396,N_36046);
or U41927 (N_41927,N_38389,N_39773);
xnor U41928 (N_41928,N_35961,N_35165);
and U41929 (N_41929,N_39651,N_39365);
nand U41930 (N_41930,N_39712,N_38120);
nand U41931 (N_41931,N_37230,N_35024);
nand U41932 (N_41932,N_39920,N_35856);
nand U41933 (N_41933,N_36433,N_35497);
and U41934 (N_41934,N_39191,N_37297);
or U41935 (N_41935,N_37821,N_35172);
or U41936 (N_41936,N_38872,N_36136);
nor U41937 (N_41937,N_39991,N_38037);
and U41938 (N_41938,N_39751,N_36047);
or U41939 (N_41939,N_38083,N_36637);
and U41940 (N_41940,N_38009,N_39693);
xor U41941 (N_41941,N_36148,N_36987);
nor U41942 (N_41942,N_38774,N_38590);
and U41943 (N_41943,N_38504,N_35332);
and U41944 (N_41944,N_36992,N_37572);
nand U41945 (N_41945,N_39033,N_36124);
nand U41946 (N_41946,N_38248,N_37648);
and U41947 (N_41947,N_36484,N_38275);
nor U41948 (N_41948,N_38912,N_37499);
xnor U41949 (N_41949,N_37022,N_35604);
nand U41950 (N_41950,N_39293,N_39065);
nor U41951 (N_41951,N_37664,N_37817);
nor U41952 (N_41952,N_35467,N_37065);
or U41953 (N_41953,N_36444,N_39814);
nor U41954 (N_41954,N_36092,N_36902);
nand U41955 (N_41955,N_36631,N_39003);
xor U41956 (N_41956,N_37836,N_38659);
and U41957 (N_41957,N_35413,N_37631);
and U41958 (N_41958,N_39271,N_35477);
nor U41959 (N_41959,N_38668,N_35229);
xnor U41960 (N_41960,N_35113,N_36182);
xnor U41961 (N_41961,N_38417,N_37458);
nor U41962 (N_41962,N_35536,N_37176);
nand U41963 (N_41963,N_37524,N_38815);
nor U41964 (N_41964,N_36746,N_35878);
nand U41965 (N_41965,N_35732,N_38202);
nor U41966 (N_41966,N_39207,N_38254);
xor U41967 (N_41967,N_39785,N_39845);
nand U41968 (N_41968,N_36650,N_35565);
nor U41969 (N_41969,N_37181,N_37915);
or U41970 (N_41970,N_38756,N_35191);
nor U41971 (N_41971,N_39389,N_37896);
nand U41972 (N_41972,N_35741,N_39565);
and U41973 (N_41973,N_36283,N_35135);
and U41974 (N_41974,N_36946,N_39818);
and U41975 (N_41975,N_36402,N_39087);
or U41976 (N_41976,N_39804,N_37830);
xnor U41977 (N_41977,N_36004,N_37405);
and U41978 (N_41978,N_35071,N_37308);
nand U41979 (N_41979,N_36324,N_36090);
and U41980 (N_41980,N_39598,N_38141);
xor U41981 (N_41981,N_38299,N_37589);
and U41982 (N_41982,N_35885,N_35585);
and U41983 (N_41983,N_39666,N_38807);
nand U41984 (N_41984,N_39965,N_38132);
xnor U41985 (N_41985,N_35747,N_35640);
nor U41986 (N_41986,N_39132,N_36177);
and U41987 (N_41987,N_38447,N_38134);
and U41988 (N_41988,N_36680,N_35802);
or U41989 (N_41989,N_37485,N_35352);
xnor U41990 (N_41990,N_38318,N_36173);
xnor U41991 (N_41991,N_35280,N_39714);
xor U41992 (N_41992,N_35588,N_36463);
xnor U41993 (N_41993,N_37828,N_38043);
nor U41994 (N_41994,N_39966,N_38450);
nand U41995 (N_41995,N_35028,N_36081);
nor U41996 (N_41996,N_39204,N_39859);
or U41997 (N_41997,N_36541,N_37428);
nand U41998 (N_41998,N_36056,N_37728);
nor U41999 (N_41999,N_36888,N_37092);
xor U42000 (N_42000,N_38225,N_38579);
nand U42001 (N_42001,N_35919,N_36663);
nand U42002 (N_42002,N_38711,N_36329);
nand U42003 (N_42003,N_36359,N_35678);
or U42004 (N_42004,N_39571,N_37480);
or U42005 (N_42005,N_39326,N_37036);
xnor U42006 (N_42006,N_39159,N_37585);
nor U42007 (N_42007,N_39540,N_39678);
nand U42008 (N_42008,N_38222,N_38589);
or U42009 (N_42009,N_37281,N_38557);
xnor U42010 (N_42010,N_37733,N_37691);
nor U42011 (N_42011,N_37217,N_38268);
xnor U42012 (N_42012,N_37710,N_35446);
xor U42013 (N_42013,N_36884,N_39290);
or U42014 (N_42014,N_38443,N_37554);
and U42015 (N_42015,N_35324,N_39245);
and U42016 (N_42016,N_35064,N_35584);
nor U42017 (N_42017,N_36794,N_37577);
nor U42018 (N_42018,N_35848,N_35996);
nand U42019 (N_42019,N_35948,N_36844);
or U42020 (N_42020,N_39482,N_39066);
and U42021 (N_42021,N_36538,N_35250);
xnor U42022 (N_42022,N_39523,N_36197);
xnor U42023 (N_42023,N_37326,N_38195);
or U42024 (N_42024,N_36963,N_36305);
nand U42025 (N_42025,N_38649,N_38197);
xor U42026 (N_42026,N_37199,N_36975);
nand U42027 (N_42027,N_39812,N_37704);
and U42028 (N_42028,N_36162,N_38467);
or U42029 (N_42029,N_36096,N_39949);
nor U42030 (N_42030,N_39411,N_39982);
or U42031 (N_42031,N_37914,N_36264);
and U42032 (N_42032,N_35252,N_37893);
nand U42033 (N_42033,N_35810,N_39108);
xor U42034 (N_42034,N_39407,N_39658);
nor U42035 (N_42035,N_37218,N_35717);
xnor U42036 (N_42036,N_37483,N_36958);
or U42037 (N_42037,N_37375,N_39467);
and U42038 (N_42038,N_37809,N_35331);
or U42039 (N_42039,N_39018,N_37871);
nor U42040 (N_42040,N_35126,N_37734);
and U42041 (N_42041,N_39026,N_35342);
and U42042 (N_42042,N_35663,N_39043);
and U42043 (N_42043,N_36996,N_35676);
xnor U42044 (N_42044,N_37552,N_35387);
and U42045 (N_42045,N_36060,N_39906);
and U42046 (N_42046,N_35012,N_35694);
xor U42047 (N_42047,N_38199,N_35592);
nand U42048 (N_42048,N_37716,N_39589);
nor U42049 (N_42049,N_35724,N_37832);
nand U42050 (N_42050,N_36086,N_37331);
xnor U42051 (N_42051,N_35797,N_38836);
xor U42052 (N_42052,N_39843,N_35822);
and U42053 (N_42053,N_36993,N_35406);
nand U42054 (N_42054,N_37205,N_35356);
nor U42055 (N_42055,N_39675,N_39399);
nand U42056 (N_42056,N_35916,N_38561);
and U42057 (N_42057,N_37359,N_37956);
and U42058 (N_42058,N_39098,N_39041);
xnor U42059 (N_42059,N_38943,N_37073);
xnor U42060 (N_42060,N_38744,N_39801);
nand U42061 (N_42061,N_39165,N_39887);
xnor U42062 (N_42062,N_38182,N_36543);
nand U42063 (N_42063,N_39516,N_38634);
nand U42064 (N_42064,N_39599,N_35558);
and U42065 (N_42065,N_39531,N_37544);
or U42066 (N_42066,N_36067,N_38742);
nand U42067 (N_42067,N_38596,N_39230);
or U42068 (N_42068,N_38592,N_36001);
xnor U42069 (N_42069,N_35911,N_35542);
nand U42070 (N_42070,N_36929,N_35098);
and U42071 (N_42071,N_35495,N_35491);
and U42072 (N_42072,N_36191,N_38427);
or U42073 (N_42073,N_35624,N_39757);
nor U42074 (N_42074,N_39254,N_35644);
and U42075 (N_42075,N_37996,N_38773);
nand U42076 (N_42076,N_36972,N_39755);
xor U42077 (N_42077,N_37014,N_37276);
nor U42078 (N_42078,N_38057,N_39838);
nor U42079 (N_42079,N_37602,N_38165);
nand U42080 (N_42080,N_36764,N_35820);
nor U42081 (N_42081,N_38941,N_39774);
xnor U42082 (N_42082,N_39029,N_35421);
and U42083 (N_42083,N_38710,N_35445);
nor U42084 (N_42084,N_35285,N_39475);
nor U42085 (N_42085,N_37971,N_35814);
or U42086 (N_42086,N_38691,N_35023);
nor U42087 (N_42087,N_39372,N_38601);
or U42088 (N_42088,N_35322,N_39708);
nand U42089 (N_42089,N_36351,N_36441);
or U42090 (N_42090,N_39258,N_39695);
and U42091 (N_42091,N_35318,N_38560);
or U42092 (N_42092,N_37982,N_36504);
and U42093 (N_42093,N_35725,N_35335);
and U42094 (N_42094,N_38474,N_38065);
xor U42095 (N_42095,N_37521,N_36469);
and U42096 (N_42096,N_39443,N_36948);
and U42097 (N_42097,N_39109,N_38351);
nor U42098 (N_42098,N_35670,N_35685);
nor U42099 (N_42099,N_39581,N_36922);
and U42100 (N_42100,N_38169,N_35843);
xnor U42101 (N_42101,N_38679,N_39942);
nor U42102 (N_42102,N_39044,N_38890);
nand U42103 (N_42103,N_36907,N_36592);
and U42104 (N_42104,N_37353,N_39452);
nor U42105 (N_42105,N_36859,N_38518);
or U42106 (N_42106,N_35232,N_39322);
or U42107 (N_42107,N_37238,N_37596);
xor U42108 (N_42108,N_37291,N_38520);
nor U42109 (N_42109,N_37990,N_35230);
xor U42110 (N_42110,N_36465,N_35222);
nor U42111 (N_42111,N_38029,N_35069);
and U42112 (N_42112,N_36156,N_35552);
xor U42113 (N_42113,N_36219,N_36999);
xnor U42114 (N_42114,N_37638,N_39058);
or U42115 (N_42115,N_36114,N_36357);
nor U42116 (N_42116,N_36510,N_35610);
nor U42117 (N_42117,N_36457,N_38203);
and U42118 (N_42118,N_39054,N_39422);
nand U42119 (N_42119,N_38536,N_38390);
nor U42120 (N_42120,N_37846,N_35494);
xnor U42121 (N_42121,N_35283,N_36825);
or U42122 (N_42122,N_38528,N_38485);
nor U42123 (N_42123,N_36346,N_37076);
nand U42124 (N_42124,N_38563,N_36977);
nor U42125 (N_42125,N_36580,N_38546);
nor U42126 (N_42126,N_37561,N_35771);
and U42127 (N_42127,N_36131,N_38439);
xor U42128 (N_42128,N_38529,N_36456);
nand U42129 (N_42129,N_37143,N_39081);
or U42130 (N_42130,N_38533,N_35618);
nor U42131 (N_42131,N_39368,N_38019);
xnor U42132 (N_42132,N_38385,N_36392);
nand U42133 (N_42133,N_36144,N_38591);
nand U42134 (N_42134,N_35181,N_37980);
nand U42135 (N_42135,N_36186,N_36231);
nand U42136 (N_42136,N_37195,N_37474);
or U42137 (N_42137,N_37874,N_36985);
nand U42138 (N_42138,N_37156,N_37599);
nand U42139 (N_42139,N_39740,N_38964);
or U42140 (N_42140,N_36613,N_35075);
nor U42141 (N_42141,N_35430,N_36379);
or U42142 (N_42142,N_36374,N_38095);
and U42143 (N_42143,N_38262,N_38402);
nor U42144 (N_42144,N_39579,N_39977);
xor U42145 (N_42145,N_36377,N_38405);
nor U42146 (N_42146,N_35292,N_35090);
nand U42147 (N_42147,N_36436,N_37192);
or U42148 (N_42148,N_38210,N_39415);
xnor U42149 (N_42149,N_37949,N_39145);
nand U42150 (N_42150,N_38808,N_39216);
or U42151 (N_42151,N_38719,N_37475);
or U42152 (N_42152,N_37707,N_39111);
or U42153 (N_42153,N_37627,N_37007);
or U42154 (N_42154,N_36062,N_36431);
xnor U42155 (N_42155,N_39154,N_38209);
nor U42156 (N_42156,N_37154,N_36769);
xnor U42157 (N_42157,N_36681,N_37090);
nand U42158 (N_42158,N_36399,N_35608);
and U42159 (N_42159,N_38316,N_35257);
nor U42160 (N_42160,N_35548,N_35052);
nor U42161 (N_42161,N_36406,N_37052);
nor U42162 (N_42162,N_37120,N_39236);
nand U42163 (N_42163,N_39013,N_37294);
nor U42164 (N_42164,N_37966,N_39877);
and U42165 (N_42165,N_36743,N_39239);
xnor U42166 (N_42166,N_37948,N_39593);
nand U42167 (N_42167,N_38160,N_38555);
and U42168 (N_42168,N_39612,N_36132);
nand U42169 (N_42169,N_36396,N_38573);
or U42170 (N_42170,N_38317,N_37016);
nor U42171 (N_42171,N_35514,N_35206);
and U42172 (N_42172,N_38392,N_35049);
and U42173 (N_42173,N_35306,N_36014);
nand U42174 (N_42174,N_38191,N_35001);
and U42175 (N_42175,N_35117,N_37963);
nor U42176 (N_42176,N_35906,N_37737);
or U42177 (N_42177,N_37740,N_36125);
nand U42178 (N_42178,N_36908,N_39471);
and U42179 (N_42179,N_36562,N_39935);
or U42180 (N_42180,N_35125,N_37207);
and U42181 (N_42181,N_38281,N_37877);
xor U42182 (N_42182,N_39931,N_37888);
nor U42183 (N_42183,N_39281,N_35951);
nand U42184 (N_42184,N_36546,N_35923);
and U42185 (N_42185,N_39248,N_35499);
nor U42186 (N_42186,N_35815,N_35894);
and U42187 (N_42187,N_36930,N_37575);
nand U42188 (N_42188,N_35000,N_37121);
and U42189 (N_42189,N_39936,N_39575);
or U42190 (N_42190,N_37647,N_36274);
and U42191 (N_42191,N_37448,N_36209);
and U42192 (N_42192,N_37298,N_36515);
xnor U42193 (N_42193,N_39960,N_36917);
and U42194 (N_42194,N_39312,N_36050);
or U42195 (N_42195,N_35451,N_38838);
and U42196 (N_42196,N_39397,N_39355);
xor U42197 (N_42197,N_38338,N_37271);
nor U42198 (N_42198,N_39257,N_37774);
nand U42199 (N_42199,N_38294,N_36424);
xor U42200 (N_42200,N_39975,N_35990);
xor U42201 (N_42201,N_36311,N_39129);
nor U42202 (N_42202,N_36430,N_35300);
or U42203 (N_42203,N_37505,N_37299);
nor U42204 (N_42204,N_37799,N_38006);
nand U42205 (N_42205,N_38238,N_35511);
nand U42206 (N_42206,N_39127,N_37089);
nor U42207 (N_42207,N_37908,N_36579);
and U42208 (N_42208,N_39419,N_36416);
xnor U42209 (N_42209,N_37881,N_37904);
or U42210 (N_42210,N_39370,N_39255);
and U42211 (N_42211,N_37655,N_36600);
nand U42212 (N_42212,N_35277,N_35611);
or U42213 (N_42213,N_36581,N_39436);
nand U42214 (N_42214,N_39558,N_36603);
xnor U42215 (N_42215,N_39319,N_36313);
nor U42216 (N_42216,N_38787,N_36791);
xor U42217 (N_42217,N_37077,N_39657);
xnor U42218 (N_42218,N_37097,N_35745);
and U42219 (N_42219,N_37226,N_37201);
and U42220 (N_42220,N_36612,N_36638);
nor U42221 (N_42221,N_36556,N_35850);
nor U42222 (N_42222,N_35569,N_35060);
and U42223 (N_42223,N_39759,N_38794);
and U42224 (N_42224,N_38856,N_37082);
and U42225 (N_42225,N_36464,N_36936);
or U42226 (N_42226,N_36790,N_38223);
nand U42227 (N_42227,N_38088,N_37465);
nor U42228 (N_42228,N_36369,N_39886);
xnor U42229 (N_42229,N_37778,N_39091);
nand U42230 (N_42230,N_38104,N_37653);
xor U42231 (N_42231,N_37580,N_39870);
and U42232 (N_42232,N_36973,N_38888);
or U42233 (N_42233,N_38369,N_36572);
nor U42234 (N_42234,N_37256,N_35889);
nor U42235 (N_42235,N_35958,N_38983);
xnor U42236 (N_42236,N_38558,N_36245);
or U42237 (N_42237,N_35935,N_38353);
nand U42238 (N_42238,N_35940,N_38967);
or U42239 (N_42239,N_37938,N_37503);
xor U42240 (N_42240,N_39073,N_38910);
and U42241 (N_42241,N_35418,N_36360);
or U42242 (N_42242,N_38343,N_38552);
xnor U42243 (N_42243,N_36221,N_38287);
and U42244 (N_42244,N_39738,N_35326);
nand U42245 (N_42245,N_38919,N_39057);
xnor U42246 (N_42246,N_36625,N_39680);
nand U42247 (N_42247,N_35044,N_37151);
nand U42248 (N_42248,N_36407,N_39704);
nor U42249 (N_42249,N_39260,N_36066);
and U42250 (N_42250,N_37010,N_37801);
and U42251 (N_42251,N_38733,N_39004);
nand U42252 (N_42252,N_39883,N_35154);
nand U42253 (N_42253,N_38214,N_35997);
nand U42254 (N_42254,N_35902,N_36866);
xor U42255 (N_42255,N_39457,N_35934);
nor U42256 (N_42256,N_39898,N_37808);
nor U42257 (N_42257,N_37962,N_39335);
or U42258 (N_42258,N_38335,N_37773);
or U42259 (N_42259,N_39888,N_35580);
nor U42260 (N_42260,N_39560,N_36363);
nand U42261 (N_42261,N_36991,N_36881);
xor U42262 (N_42262,N_38631,N_37630);
xnor U42263 (N_42263,N_39119,N_36126);
nand U42264 (N_42264,N_36095,N_38692);
nand U42265 (N_42265,N_36636,N_35163);
nand U42266 (N_42266,N_35866,N_39849);
or U42267 (N_42267,N_37619,N_38356);
or U42268 (N_42268,N_37766,N_38702);
nor U42269 (N_42269,N_38368,N_35147);
nor U42270 (N_42270,N_35599,N_39323);
and U42271 (N_42271,N_36307,N_37462);
nand U42272 (N_42272,N_37086,N_39120);
nand U42273 (N_42273,N_35002,N_36845);
nand U42274 (N_42274,N_36166,N_38532);
or U42275 (N_42275,N_38030,N_38207);
nor U42276 (N_42276,N_36334,N_37123);
and U42277 (N_42277,N_35449,N_39642);
xor U42278 (N_42278,N_39534,N_37514);
nor U42279 (N_42279,N_35372,N_38153);
nand U42280 (N_42280,N_37752,N_35651);
xor U42281 (N_42281,N_38829,N_39973);
and U42282 (N_42282,N_36170,N_37023);
nor U42283 (N_42283,N_38683,N_37711);
or U42284 (N_42284,N_35212,N_37758);
nand U42285 (N_42285,N_38022,N_39998);
nand U42286 (N_42286,N_39884,N_38085);
nor U42287 (N_42287,N_35183,N_36432);
xnor U42288 (N_42288,N_35699,N_39901);
nor U42289 (N_42289,N_37155,N_36819);
nand U42290 (N_42290,N_38278,N_38516);
nor U42291 (N_42291,N_37674,N_39915);
xor U42292 (N_42292,N_39178,N_35879);
xor U42293 (N_42293,N_35852,N_35525);
or U42294 (N_42294,N_38980,N_39206);
or U42295 (N_42295,N_39195,N_38747);
nor U42296 (N_42296,N_37437,N_36158);
and U42297 (N_42297,N_35472,N_35267);
nor U42298 (N_42298,N_37333,N_39813);
and U42299 (N_42299,N_38418,N_36378);
nand U42300 (N_42300,N_37351,N_37570);
nand U42301 (N_42301,N_39619,N_35970);
xnor U42302 (N_42302,N_35376,N_35132);
xnor U42303 (N_42303,N_36321,N_39866);
or U42304 (N_42304,N_37398,N_39071);
xor U42305 (N_42305,N_37344,N_39972);
or U42306 (N_42306,N_39796,N_38125);
and U42307 (N_42307,N_37725,N_35110);
nand U42308 (N_42308,N_35480,N_35945);
nand U42309 (N_42309,N_38481,N_38797);
or U42310 (N_42310,N_36643,N_36390);
and U42311 (N_42311,N_35767,N_36445);
nand U42312 (N_42312,N_38501,N_37715);
and U42313 (N_42313,N_35251,N_39634);
or U42314 (N_42314,N_37390,N_38842);
nand U42315 (N_42315,N_37854,N_39921);
nand U42316 (N_42316,N_35746,N_39435);
xnor U42317 (N_42317,N_38718,N_38149);
xnor U42318 (N_42318,N_39641,N_39364);
xor U42319 (N_42319,N_38457,N_39803);
xnor U42320 (N_42320,N_36462,N_36118);
and U42321 (N_42321,N_36134,N_35496);
nand U42322 (N_42322,N_39259,N_36003);
xor U42323 (N_42323,N_35360,N_35053);
xnor U42324 (N_42324,N_36237,N_37770);
or U42325 (N_42325,N_38974,N_37727);
nand U42326 (N_42326,N_38622,N_37719);
nand U42327 (N_42327,N_36043,N_37779);
xnor U42328 (N_42328,N_39286,N_36108);
or U42329 (N_42329,N_35488,N_36496);
nand U42330 (N_42330,N_38627,N_37087);
and U42331 (N_42331,N_39535,N_39903);
nor U42332 (N_42332,N_39971,N_39656);
nand U42333 (N_42333,N_37034,N_35758);
or U42334 (N_42334,N_35547,N_35305);
nand U42335 (N_42335,N_39784,N_37243);
and U42336 (N_42336,N_39790,N_36204);
xnor U42337 (N_42337,N_39083,N_37000);
xnor U42338 (N_42338,N_38414,N_35659);
xor U42339 (N_42339,N_39384,N_37623);
nand U42340 (N_42340,N_37075,N_37600);
nor U42341 (N_42341,N_39546,N_37882);
xor U42342 (N_42342,N_38615,N_36548);
nand U42343 (N_42343,N_36300,N_37030);
nor U42344 (N_42344,N_35403,N_35249);
or U42345 (N_42345,N_37399,N_35242);
xnor U42346 (N_42346,N_36644,N_36718);
xor U42347 (N_42347,N_36698,N_37055);
and U42348 (N_42348,N_39140,N_38445);
nor U42349 (N_42349,N_35029,N_38613);
or U42350 (N_42350,N_38600,N_38266);
xor U42351 (N_42351,N_37202,N_39063);
xnor U42352 (N_42352,N_37992,N_38653);
or U42353 (N_42353,N_39410,N_39995);
nor U42354 (N_42354,N_38323,N_39737);
xnor U42355 (N_42355,N_36098,N_37511);
xnor U42356 (N_42356,N_35920,N_37106);
or U42357 (N_42357,N_35004,N_39017);
nor U42358 (N_42358,N_35311,N_38578);
nor U42359 (N_42359,N_37868,N_35544);
or U42360 (N_42360,N_37588,N_38140);
or U42361 (N_42361,N_39918,N_37560);
xor U42362 (N_42362,N_37670,N_36838);
nor U42363 (N_42363,N_35643,N_38795);
xor U42364 (N_42364,N_36097,N_35541);
and U42365 (N_42365,N_36336,N_35466);
or U42366 (N_42366,N_37831,N_39042);
or U42367 (N_42367,N_38788,N_39566);
xor U42368 (N_42368,N_36503,N_36986);
and U42369 (N_42369,N_36893,N_35476);
xor U42370 (N_42370,N_35564,N_35830);
nor U42371 (N_42371,N_36599,N_37529);
or U42372 (N_42372,N_36923,N_36618);
or U42373 (N_42373,N_39721,N_37043);
and U42374 (N_42374,N_39118,N_36068);
or U42375 (N_42375,N_37813,N_37223);
xor U42376 (N_42376,N_36449,N_37248);
nand U42377 (N_42377,N_36195,N_35253);
or U42378 (N_42378,N_38212,N_35567);
and U42379 (N_42379,N_36163,N_39894);
nor U42380 (N_42380,N_35922,N_35015);
or U42381 (N_42381,N_38420,N_39006);
nand U42382 (N_42382,N_38864,N_39052);
nor U42383 (N_42383,N_37676,N_35939);
xor U42384 (N_42384,N_39143,N_35688);
xnor U42385 (N_42385,N_39155,N_39150);
or U42386 (N_42386,N_39730,N_35783);
xnor U42387 (N_42387,N_39690,N_37533);
nor U42388 (N_42388,N_35027,N_35989);
nand U42389 (N_42389,N_36319,N_36792);
and U42390 (N_42390,N_37957,N_36239);
nand U42391 (N_42391,N_38507,N_39313);
xor U42392 (N_42392,N_35014,N_37720);
or U42393 (N_42393,N_39912,N_36573);
nand U42394 (N_42394,N_39197,N_35721);
xor U42395 (N_42395,N_37792,N_36871);
and U42396 (N_42396,N_39241,N_37170);
nor U42397 (N_42397,N_35174,N_38170);
xnor U42398 (N_42398,N_35692,N_38168);
or U42399 (N_42399,N_36502,N_37891);
nor U42400 (N_42400,N_37687,N_35068);
nor U42401 (N_42401,N_37921,N_39493);
nor U42402 (N_42402,N_36312,N_35284);
or U42403 (N_42403,N_37850,N_36811);
nor U42404 (N_42404,N_38042,N_37210);
nand U42405 (N_42405,N_36121,N_39947);
or U42406 (N_42406,N_37212,N_35294);
nand U42407 (N_42407,N_38465,N_39891);
nand U42408 (N_42408,N_39330,N_37312);
nand U42409 (N_42409,N_38772,N_39180);
nand U42410 (N_42410,N_37365,N_36672);
nand U42411 (N_42411,N_36350,N_36380);
or U42412 (N_42412,N_37352,N_38084);
xnor U42413 (N_42413,N_36989,N_38224);
nand U42414 (N_42414,N_36941,N_37502);
nor U42415 (N_42415,N_36192,N_37189);
nor U42416 (N_42416,N_38401,N_38310);
nor U42417 (N_42417,N_38430,N_35960);
xor U42418 (N_42418,N_39199,N_37177);
nor U42419 (N_42419,N_37191,N_39908);
nor U42420 (N_42420,N_38386,N_35854);
xor U42421 (N_42421,N_39039,N_37320);
xor U42422 (N_42422,N_36421,N_39099);
nand U42423 (N_42423,N_36968,N_35122);
xnor U42424 (N_42424,N_38312,N_37678);
nand U42425 (N_42425,N_36676,N_39469);
nand U42426 (N_42426,N_35435,N_39621);
and U42427 (N_42427,N_35615,N_36775);
xnor U42428 (N_42428,N_35667,N_36337);
nand U42429 (N_42429,N_37794,N_39437);
nor U42430 (N_42430,N_35897,N_37340);
and U42431 (N_42431,N_39861,N_38574);
xor U42432 (N_42432,N_36018,N_37165);
nor U42433 (N_42433,N_36632,N_36809);
nor U42434 (N_42434,N_35673,N_35605);
or U42435 (N_42435,N_39600,N_37258);
or U42436 (N_42436,N_38180,N_36520);
nor U42437 (N_42437,N_38818,N_39953);
or U42438 (N_42438,N_39380,N_39911);
or U42439 (N_42439,N_37510,N_37349);
and U42440 (N_42440,N_36796,N_35622);
or U42441 (N_42441,N_38969,N_39481);
or U42442 (N_42442,N_35145,N_39529);
xnor U42443 (N_42443,N_38496,N_37409);
xnor U42444 (N_42444,N_39741,N_36729);
nor U42445 (N_42445,N_37883,N_39509);
xor U42446 (N_42446,N_37937,N_37953);
xor U42447 (N_42447,N_38761,N_38079);
nor U42448 (N_42448,N_36295,N_36035);
or U42449 (N_42449,N_36475,N_38173);
xnor U42450 (N_42450,N_39494,N_36101);
or U42451 (N_42451,N_38986,N_38514);
xor U42452 (N_42452,N_39985,N_37088);
or U42453 (N_42453,N_35188,N_36606);
nand U42454 (N_42454,N_39454,N_38621);
xor U42455 (N_42455,N_37386,N_37581);
nor U42456 (N_42456,N_35677,N_39900);
nor U42457 (N_42457,N_36106,N_36453);
nor U42458 (N_42458,N_35380,N_36834);
xnor U42459 (N_42459,N_36689,N_37759);
and U42460 (N_42460,N_38461,N_38221);
nand U42461 (N_42461,N_39826,N_37188);
nand U42462 (N_42462,N_38400,N_39692);
or U42463 (N_42463,N_37193,N_36111);
nor U42464 (N_42464,N_37426,N_36200);
xnor U42465 (N_42465,N_38616,N_37516);
and U42466 (N_42466,N_38698,N_38951);
or U42467 (N_42467,N_35642,N_36890);
and U42468 (N_42468,N_37459,N_35092);
or U42469 (N_42469,N_37270,N_35731);
nor U42470 (N_42470,N_36394,N_37764);
nand U42471 (N_42471,N_37873,N_38300);
nand U42472 (N_42472,N_39133,N_36331);
nand U42473 (N_42473,N_39196,N_39016);
or U42474 (N_42474,N_38399,N_39798);
xnor U42475 (N_42475,N_37654,N_38885);
and U42476 (N_42476,N_37254,N_35276);
nand U42477 (N_42477,N_37901,N_37955);
nor U42478 (N_42478,N_37824,N_36253);
or U42479 (N_42479,N_39332,N_37532);
and U42480 (N_42480,N_37806,N_39848);
and U42481 (N_42481,N_35985,N_36909);
or U42482 (N_42482,N_36263,N_35392);
nor U42483 (N_42483,N_35812,N_36492);
and U42484 (N_42484,N_38657,N_36892);
nand U42485 (N_42485,N_36381,N_38320);
or U42486 (N_42486,N_37583,N_39473);
nand U42487 (N_42487,N_35900,N_38685);
nand U42488 (N_42488,N_39691,N_35262);
nor U42489 (N_42489,N_36145,N_35620);
or U42490 (N_42490,N_36517,N_38412);
nor U42491 (N_42491,N_35975,N_38629);
and U42492 (N_42492,N_37119,N_37091);
xor U42493 (N_42493,N_37040,N_36355);
or U42494 (N_42494,N_37182,N_35795);
xor U42495 (N_42495,N_37820,N_36241);
xnor U42496 (N_42496,N_38819,N_36323);
and U42497 (N_42497,N_36450,N_37279);
and U42498 (N_42498,N_35056,N_36024);
nor U42499 (N_42499,N_35368,N_38045);
nor U42500 (N_42500,N_38915,N_38427);
nor U42501 (N_42501,N_35450,N_39784);
nor U42502 (N_42502,N_35941,N_37088);
nor U42503 (N_42503,N_39087,N_36416);
or U42504 (N_42504,N_37581,N_39728);
nor U42505 (N_42505,N_38282,N_39951);
nor U42506 (N_42506,N_39531,N_35347);
xor U42507 (N_42507,N_39944,N_35424);
xor U42508 (N_42508,N_38254,N_37520);
nor U42509 (N_42509,N_37630,N_36528);
xor U42510 (N_42510,N_38797,N_38830);
nor U42511 (N_42511,N_38207,N_38980);
nor U42512 (N_42512,N_36008,N_35550);
or U42513 (N_42513,N_36093,N_39746);
and U42514 (N_42514,N_35436,N_39581);
xor U42515 (N_42515,N_36252,N_38762);
nand U42516 (N_42516,N_38824,N_36934);
and U42517 (N_42517,N_37639,N_39419);
nor U42518 (N_42518,N_39669,N_35686);
nor U42519 (N_42519,N_39929,N_35311);
or U42520 (N_42520,N_36065,N_35749);
nand U42521 (N_42521,N_37785,N_35966);
xor U42522 (N_42522,N_37046,N_36190);
nand U42523 (N_42523,N_38845,N_36123);
nand U42524 (N_42524,N_35397,N_39689);
nor U42525 (N_42525,N_36553,N_37727);
nand U42526 (N_42526,N_38796,N_35331);
nand U42527 (N_42527,N_37076,N_36067);
xnor U42528 (N_42528,N_36608,N_35449);
nor U42529 (N_42529,N_36278,N_36819);
nand U42530 (N_42530,N_38549,N_37362);
nor U42531 (N_42531,N_38540,N_35032);
or U42532 (N_42532,N_39187,N_39411);
xor U42533 (N_42533,N_35588,N_37037);
and U42534 (N_42534,N_36592,N_36344);
nand U42535 (N_42535,N_35898,N_39279);
nor U42536 (N_42536,N_39865,N_38460);
nor U42537 (N_42537,N_37096,N_35088);
nor U42538 (N_42538,N_38489,N_38727);
and U42539 (N_42539,N_36976,N_35294);
nand U42540 (N_42540,N_35362,N_35413);
nor U42541 (N_42541,N_37503,N_35046);
xnor U42542 (N_42542,N_35854,N_36008);
nor U42543 (N_42543,N_37905,N_37835);
and U42544 (N_42544,N_38520,N_39917);
xnor U42545 (N_42545,N_35803,N_39297);
or U42546 (N_42546,N_39566,N_37882);
or U42547 (N_42547,N_37787,N_36623);
nand U42548 (N_42548,N_35802,N_35292);
nand U42549 (N_42549,N_37402,N_39841);
and U42550 (N_42550,N_36761,N_37028);
nand U42551 (N_42551,N_36095,N_37686);
nor U42552 (N_42552,N_36197,N_35564);
nor U42553 (N_42553,N_39312,N_38479);
xnor U42554 (N_42554,N_36429,N_37667);
and U42555 (N_42555,N_36067,N_37392);
xor U42556 (N_42556,N_38702,N_35615);
or U42557 (N_42557,N_35029,N_38522);
nor U42558 (N_42558,N_35287,N_39174);
or U42559 (N_42559,N_39325,N_37691);
xor U42560 (N_42560,N_38423,N_36999);
nand U42561 (N_42561,N_39179,N_39028);
xnor U42562 (N_42562,N_35927,N_39482);
or U42563 (N_42563,N_39054,N_38754);
and U42564 (N_42564,N_37267,N_37699);
and U42565 (N_42565,N_37821,N_38494);
nor U42566 (N_42566,N_38779,N_36111);
and U42567 (N_42567,N_37138,N_37276);
xnor U42568 (N_42568,N_36206,N_39873);
xor U42569 (N_42569,N_37499,N_39752);
or U42570 (N_42570,N_38235,N_37123);
or U42571 (N_42571,N_38160,N_35015);
xor U42572 (N_42572,N_38622,N_37632);
xor U42573 (N_42573,N_35174,N_35959);
and U42574 (N_42574,N_39993,N_38702);
or U42575 (N_42575,N_38821,N_39528);
nand U42576 (N_42576,N_39947,N_35851);
nand U42577 (N_42577,N_35887,N_35397);
or U42578 (N_42578,N_38051,N_35693);
nor U42579 (N_42579,N_37702,N_38567);
and U42580 (N_42580,N_37166,N_36751);
or U42581 (N_42581,N_38078,N_37521);
and U42582 (N_42582,N_35570,N_37194);
nand U42583 (N_42583,N_35464,N_37618);
or U42584 (N_42584,N_36638,N_38103);
and U42585 (N_42585,N_39015,N_38737);
xor U42586 (N_42586,N_35212,N_35774);
and U42587 (N_42587,N_36264,N_37379);
and U42588 (N_42588,N_39520,N_37787);
and U42589 (N_42589,N_35749,N_35328);
nand U42590 (N_42590,N_39421,N_39795);
nor U42591 (N_42591,N_35369,N_39933);
nor U42592 (N_42592,N_39982,N_38129);
nand U42593 (N_42593,N_37087,N_36389);
xnor U42594 (N_42594,N_39389,N_38744);
and U42595 (N_42595,N_35096,N_35286);
or U42596 (N_42596,N_35897,N_38553);
and U42597 (N_42597,N_35625,N_35416);
and U42598 (N_42598,N_38587,N_37869);
nor U42599 (N_42599,N_38344,N_38529);
and U42600 (N_42600,N_39584,N_36236);
nor U42601 (N_42601,N_36205,N_35087);
and U42602 (N_42602,N_36359,N_37194);
or U42603 (N_42603,N_35939,N_37592);
xor U42604 (N_42604,N_35974,N_39817);
and U42605 (N_42605,N_36454,N_37917);
or U42606 (N_42606,N_36834,N_35839);
xor U42607 (N_42607,N_38257,N_38352);
xnor U42608 (N_42608,N_37459,N_39464);
xor U42609 (N_42609,N_38929,N_36370);
xor U42610 (N_42610,N_37267,N_35952);
or U42611 (N_42611,N_36581,N_36746);
nand U42612 (N_42612,N_36256,N_37178);
and U42613 (N_42613,N_39757,N_39681);
or U42614 (N_42614,N_36861,N_35642);
or U42615 (N_42615,N_39439,N_39321);
or U42616 (N_42616,N_35277,N_38325);
nand U42617 (N_42617,N_38253,N_36905);
and U42618 (N_42618,N_39408,N_35173);
and U42619 (N_42619,N_35460,N_35044);
or U42620 (N_42620,N_37279,N_35667);
and U42621 (N_42621,N_36745,N_36062);
or U42622 (N_42622,N_35160,N_38163);
xor U42623 (N_42623,N_38251,N_36611);
or U42624 (N_42624,N_37372,N_37032);
nand U42625 (N_42625,N_38015,N_39640);
nand U42626 (N_42626,N_35168,N_37672);
and U42627 (N_42627,N_37514,N_38674);
xnor U42628 (N_42628,N_36940,N_38910);
or U42629 (N_42629,N_37810,N_35136);
nor U42630 (N_42630,N_39959,N_38766);
nand U42631 (N_42631,N_39334,N_37721);
nor U42632 (N_42632,N_36416,N_37285);
nand U42633 (N_42633,N_35217,N_39206);
or U42634 (N_42634,N_37027,N_38432);
nand U42635 (N_42635,N_38043,N_37935);
nor U42636 (N_42636,N_35141,N_36560);
nor U42637 (N_42637,N_38614,N_35103);
or U42638 (N_42638,N_37636,N_35030);
nand U42639 (N_42639,N_38429,N_38399);
nand U42640 (N_42640,N_37712,N_36775);
xor U42641 (N_42641,N_39556,N_38278);
nor U42642 (N_42642,N_39278,N_36103);
or U42643 (N_42643,N_38176,N_35645);
or U42644 (N_42644,N_38139,N_35266);
nand U42645 (N_42645,N_36092,N_38861);
and U42646 (N_42646,N_37177,N_36093);
xnor U42647 (N_42647,N_39634,N_37255);
and U42648 (N_42648,N_37227,N_37368);
or U42649 (N_42649,N_39478,N_38060);
nand U42650 (N_42650,N_39901,N_35581);
nand U42651 (N_42651,N_35190,N_36050);
and U42652 (N_42652,N_39104,N_36095);
xnor U42653 (N_42653,N_38349,N_38029);
nor U42654 (N_42654,N_37864,N_36991);
nor U42655 (N_42655,N_38153,N_39854);
or U42656 (N_42656,N_37296,N_39509);
or U42657 (N_42657,N_36147,N_39506);
xor U42658 (N_42658,N_36575,N_38163);
and U42659 (N_42659,N_35732,N_39789);
xnor U42660 (N_42660,N_38575,N_37387);
or U42661 (N_42661,N_35490,N_37210);
xnor U42662 (N_42662,N_36971,N_35867);
nor U42663 (N_42663,N_37976,N_36482);
xor U42664 (N_42664,N_39343,N_35710);
nand U42665 (N_42665,N_36473,N_35730);
nor U42666 (N_42666,N_38854,N_37286);
xnor U42667 (N_42667,N_35451,N_39253);
nand U42668 (N_42668,N_39295,N_38637);
or U42669 (N_42669,N_36554,N_35634);
nor U42670 (N_42670,N_38970,N_36231);
nor U42671 (N_42671,N_36403,N_36295);
xor U42672 (N_42672,N_37600,N_39958);
xnor U42673 (N_42673,N_39862,N_37041);
and U42674 (N_42674,N_36520,N_36454);
nand U42675 (N_42675,N_36789,N_36980);
nand U42676 (N_42676,N_38829,N_35121);
xor U42677 (N_42677,N_38823,N_39520);
nor U42678 (N_42678,N_35069,N_36189);
nand U42679 (N_42679,N_37439,N_36128);
nand U42680 (N_42680,N_38683,N_37274);
xor U42681 (N_42681,N_37239,N_36587);
or U42682 (N_42682,N_39310,N_39451);
or U42683 (N_42683,N_38895,N_35275);
and U42684 (N_42684,N_37285,N_36764);
nand U42685 (N_42685,N_38737,N_39677);
nand U42686 (N_42686,N_37608,N_35818);
or U42687 (N_42687,N_36352,N_35530);
or U42688 (N_42688,N_37128,N_38738);
nand U42689 (N_42689,N_35191,N_36649);
or U42690 (N_42690,N_36794,N_35780);
xor U42691 (N_42691,N_39000,N_36738);
and U42692 (N_42692,N_38908,N_37741);
xnor U42693 (N_42693,N_38030,N_39048);
nand U42694 (N_42694,N_35125,N_37552);
or U42695 (N_42695,N_39188,N_35562);
nand U42696 (N_42696,N_39390,N_38451);
nand U42697 (N_42697,N_36502,N_37248);
or U42698 (N_42698,N_37500,N_36534);
nor U42699 (N_42699,N_36300,N_35340);
nand U42700 (N_42700,N_37976,N_39636);
or U42701 (N_42701,N_38688,N_36240);
and U42702 (N_42702,N_38859,N_35389);
and U42703 (N_42703,N_35703,N_39866);
nor U42704 (N_42704,N_37786,N_39769);
and U42705 (N_42705,N_36376,N_35188);
xor U42706 (N_42706,N_39360,N_37947);
or U42707 (N_42707,N_36606,N_36907);
nand U42708 (N_42708,N_36026,N_38023);
or U42709 (N_42709,N_38973,N_39794);
nor U42710 (N_42710,N_35597,N_39180);
xnor U42711 (N_42711,N_35622,N_39410);
xnor U42712 (N_42712,N_39112,N_36925);
or U42713 (N_42713,N_35871,N_39964);
xnor U42714 (N_42714,N_36690,N_36898);
nor U42715 (N_42715,N_35443,N_38396);
nand U42716 (N_42716,N_39364,N_39980);
nand U42717 (N_42717,N_39903,N_37257);
nor U42718 (N_42718,N_36763,N_37548);
xnor U42719 (N_42719,N_36366,N_36064);
nand U42720 (N_42720,N_38461,N_35504);
or U42721 (N_42721,N_38883,N_38141);
and U42722 (N_42722,N_37579,N_39328);
xnor U42723 (N_42723,N_39251,N_38439);
and U42724 (N_42724,N_36381,N_37439);
and U42725 (N_42725,N_36490,N_36043);
or U42726 (N_42726,N_37017,N_37225);
xnor U42727 (N_42727,N_35587,N_35307);
nor U42728 (N_42728,N_36457,N_38379);
or U42729 (N_42729,N_39972,N_37995);
xor U42730 (N_42730,N_35474,N_38219);
xor U42731 (N_42731,N_36418,N_38957);
nand U42732 (N_42732,N_39318,N_37023);
nor U42733 (N_42733,N_39297,N_39661);
nand U42734 (N_42734,N_37872,N_38963);
or U42735 (N_42735,N_37990,N_37557);
nor U42736 (N_42736,N_38118,N_39022);
nor U42737 (N_42737,N_35417,N_38756);
nor U42738 (N_42738,N_35521,N_35583);
nand U42739 (N_42739,N_39075,N_37190);
nor U42740 (N_42740,N_37909,N_35984);
or U42741 (N_42741,N_38457,N_36416);
nand U42742 (N_42742,N_38967,N_35128);
xnor U42743 (N_42743,N_37953,N_38507);
nor U42744 (N_42744,N_38474,N_37492);
and U42745 (N_42745,N_37571,N_38177);
and U42746 (N_42746,N_39035,N_39391);
nand U42747 (N_42747,N_36338,N_35928);
or U42748 (N_42748,N_35951,N_38857);
and U42749 (N_42749,N_36010,N_39938);
or U42750 (N_42750,N_38084,N_38338);
or U42751 (N_42751,N_37292,N_39138);
and U42752 (N_42752,N_37828,N_35602);
nand U42753 (N_42753,N_38860,N_37475);
and U42754 (N_42754,N_39608,N_36284);
xor U42755 (N_42755,N_39986,N_35219);
xnor U42756 (N_42756,N_37947,N_35460);
or U42757 (N_42757,N_39576,N_35552);
or U42758 (N_42758,N_35612,N_36927);
nand U42759 (N_42759,N_36871,N_36846);
xnor U42760 (N_42760,N_38135,N_39851);
xnor U42761 (N_42761,N_36573,N_39950);
and U42762 (N_42762,N_37285,N_39967);
xor U42763 (N_42763,N_37456,N_35560);
nor U42764 (N_42764,N_36166,N_38522);
or U42765 (N_42765,N_36458,N_36501);
xnor U42766 (N_42766,N_35915,N_35404);
nor U42767 (N_42767,N_37336,N_35186);
nor U42768 (N_42768,N_39883,N_35227);
nor U42769 (N_42769,N_37217,N_38397);
nor U42770 (N_42770,N_36584,N_36853);
nand U42771 (N_42771,N_37122,N_39449);
nand U42772 (N_42772,N_36391,N_37342);
nor U42773 (N_42773,N_39052,N_39807);
and U42774 (N_42774,N_39128,N_38316);
nand U42775 (N_42775,N_39254,N_36502);
or U42776 (N_42776,N_38714,N_36662);
nor U42777 (N_42777,N_37925,N_38061);
xor U42778 (N_42778,N_36613,N_35291);
or U42779 (N_42779,N_36888,N_38033);
nand U42780 (N_42780,N_38277,N_37474);
nor U42781 (N_42781,N_35407,N_35659);
or U42782 (N_42782,N_37592,N_37297);
nand U42783 (N_42783,N_37756,N_36783);
or U42784 (N_42784,N_36963,N_38439);
nand U42785 (N_42785,N_38066,N_36070);
nor U42786 (N_42786,N_35022,N_38452);
xor U42787 (N_42787,N_37991,N_37368);
nand U42788 (N_42788,N_35707,N_37220);
or U42789 (N_42789,N_36135,N_37669);
xor U42790 (N_42790,N_35621,N_36447);
nand U42791 (N_42791,N_38051,N_36896);
nor U42792 (N_42792,N_37444,N_39287);
or U42793 (N_42793,N_37722,N_38432);
nor U42794 (N_42794,N_35701,N_37438);
xnor U42795 (N_42795,N_39845,N_37556);
xnor U42796 (N_42796,N_37376,N_36883);
or U42797 (N_42797,N_38448,N_36128);
nand U42798 (N_42798,N_39586,N_39434);
xor U42799 (N_42799,N_39652,N_38027);
nor U42800 (N_42800,N_39049,N_35377);
nand U42801 (N_42801,N_35326,N_37047);
and U42802 (N_42802,N_38765,N_36229);
xnor U42803 (N_42803,N_37627,N_35297);
or U42804 (N_42804,N_37396,N_37435);
and U42805 (N_42805,N_39142,N_35945);
xor U42806 (N_42806,N_39575,N_37767);
and U42807 (N_42807,N_36301,N_38102);
xnor U42808 (N_42808,N_36837,N_39103);
nor U42809 (N_42809,N_35429,N_37070);
nor U42810 (N_42810,N_37643,N_39668);
nand U42811 (N_42811,N_35321,N_36931);
nor U42812 (N_42812,N_36394,N_39346);
nand U42813 (N_42813,N_37347,N_38078);
or U42814 (N_42814,N_35439,N_35207);
and U42815 (N_42815,N_37281,N_37528);
xnor U42816 (N_42816,N_36819,N_39374);
and U42817 (N_42817,N_39277,N_39154);
nor U42818 (N_42818,N_36454,N_37200);
and U42819 (N_42819,N_37122,N_35315);
nor U42820 (N_42820,N_37342,N_37466);
and U42821 (N_42821,N_35846,N_36518);
or U42822 (N_42822,N_35985,N_37692);
nand U42823 (N_42823,N_37730,N_38352);
and U42824 (N_42824,N_36556,N_39370);
and U42825 (N_42825,N_35494,N_38682);
and U42826 (N_42826,N_39202,N_36491);
xor U42827 (N_42827,N_35861,N_38833);
nand U42828 (N_42828,N_36994,N_39213);
and U42829 (N_42829,N_39609,N_37744);
or U42830 (N_42830,N_36157,N_39049);
nor U42831 (N_42831,N_38561,N_37010);
nand U42832 (N_42832,N_38383,N_35013);
and U42833 (N_42833,N_36578,N_38111);
or U42834 (N_42834,N_35742,N_36887);
nor U42835 (N_42835,N_35541,N_38943);
and U42836 (N_42836,N_35094,N_39428);
or U42837 (N_42837,N_35191,N_39315);
nand U42838 (N_42838,N_36426,N_36184);
xnor U42839 (N_42839,N_35949,N_35454);
nand U42840 (N_42840,N_38963,N_36104);
xnor U42841 (N_42841,N_38763,N_39658);
xor U42842 (N_42842,N_38697,N_38156);
nor U42843 (N_42843,N_36915,N_36339);
or U42844 (N_42844,N_36024,N_35895);
and U42845 (N_42845,N_38817,N_35568);
or U42846 (N_42846,N_39912,N_39325);
and U42847 (N_42847,N_35409,N_35907);
or U42848 (N_42848,N_38257,N_38412);
nand U42849 (N_42849,N_38953,N_38870);
nor U42850 (N_42850,N_38634,N_37155);
or U42851 (N_42851,N_39152,N_36817);
xor U42852 (N_42852,N_38796,N_37003);
xnor U42853 (N_42853,N_39138,N_36212);
nand U42854 (N_42854,N_39550,N_36053);
and U42855 (N_42855,N_36051,N_35416);
nand U42856 (N_42856,N_39429,N_36156);
nand U42857 (N_42857,N_35085,N_38438);
xor U42858 (N_42858,N_36244,N_38641);
or U42859 (N_42859,N_39955,N_39427);
or U42860 (N_42860,N_39125,N_36351);
nor U42861 (N_42861,N_36435,N_38120);
xnor U42862 (N_42862,N_39360,N_36314);
or U42863 (N_42863,N_36469,N_36836);
xnor U42864 (N_42864,N_35548,N_35879);
and U42865 (N_42865,N_39528,N_36710);
and U42866 (N_42866,N_39320,N_38335);
nor U42867 (N_42867,N_36862,N_39658);
and U42868 (N_42868,N_35900,N_38853);
nor U42869 (N_42869,N_38879,N_36132);
and U42870 (N_42870,N_38116,N_38750);
or U42871 (N_42871,N_39030,N_38754);
xor U42872 (N_42872,N_39233,N_38810);
nand U42873 (N_42873,N_35685,N_37856);
or U42874 (N_42874,N_37873,N_37804);
or U42875 (N_42875,N_37682,N_39368);
nand U42876 (N_42876,N_37406,N_37182);
and U42877 (N_42877,N_39157,N_38969);
or U42878 (N_42878,N_39139,N_36488);
and U42879 (N_42879,N_38665,N_36385);
and U42880 (N_42880,N_35964,N_36079);
xnor U42881 (N_42881,N_36258,N_39400);
xor U42882 (N_42882,N_37170,N_36482);
nand U42883 (N_42883,N_38147,N_36259);
and U42884 (N_42884,N_35666,N_39335);
nor U42885 (N_42885,N_36914,N_39085);
xnor U42886 (N_42886,N_36164,N_38886);
or U42887 (N_42887,N_37126,N_39425);
nand U42888 (N_42888,N_35764,N_36206);
nand U42889 (N_42889,N_38483,N_38848);
and U42890 (N_42890,N_38530,N_37457);
nor U42891 (N_42891,N_35901,N_38086);
nand U42892 (N_42892,N_39137,N_38787);
or U42893 (N_42893,N_36489,N_38989);
nand U42894 (N_42894,N_35157,N_39971);
or U42895 (N_42895,N_35882,N_39476);
nor U42896 (N_42896,N_36040,N_37583);
nor U42897 (N_42897,N_38046,N_39421);
xor U42898 (N_42898,N_35356,N_39063);
xnor U42899 (N_42899,N_38787,N_35542);
nor U42900 (N_42900,N_36711,N_36348);
or U42901 (N_42901,N_35754,N_38496);
or U42902 (N_42902,N_39832,N_38099);
xnor U42903 (N_42903,N_35814,N_39177);
or U42904 (N_42904,N_36046,N_37558);
and U42905 (N_42905,N_37870,N_36859);
and U42906 (N_42906,N_37522,N_35227);
or U42907 (N_42907,N_37837,N_36703);
or U42908 (N_42908,N_38391,N_37824);
nor U42909 (N_42909,N_36869,N_37174);
and U42910 (N_42910,N_36320,N_39780);
or U42911 (N_42911,N_35947,N_37682);
and U42912 (N_42912,N_37592,N_37009);
or U42913 (N_42913,N_38295,N_38476);
or U42914 (N_42914,N_37253,N_38649);
nor U42915 (N_42915,N_38857,N_38632);
xor U42916 (N_42916,N_35949,N_37796);
nor U42917 (N_42917,N_37347,N_38777);
or U42918 (N_42918,N_35946,N_39073);
xnor U42919 (N_42919,N_37650,N_38626);
nand U42920 (N_42920,N_39248,N_38744);
and U42921 (N_42921,N_37319,N_38675);
nor U42922 (N_42922,N_37988,N_37495);
nand U42923 (N_42923,N_35321,N_37648);
and U42924 (N_42924,N_38361,N_37470);
xnor U42925 (N_42925,N_35855,N_39027);
nand U42926 (N_42926,N_37962,N_36348);
or U42927 (N_42927,N_37617,N_39303);
or U42928 (N_42928,N_39612,N_36495);
or U42929 (N_42929,N_37949,N_38264);
nand U42930 (N_42930,N_35137,N_39100);
xnor U42931 (N_42931,N_37308,N_37916);
nand U42932 (N_42932,N_36622,N_35268);
or U42933 (N_42933,N_37717,N_39082);
and U42934 (N_42934,N_36786,N_39905);
nand U42935 (N_42935,N_38240,N_38402);
nor U42936 (N_42936,N_36327,N_39753);
nand U42937 (N_42937,N_36404,N_38245);
xnor U42938 (N_42938,N_36310,N_37406);
nor U42939 (N_42939,N_39628,N_38103);
nor U42940 (N_42940,N_37566,N_35516);
nor U42941 (N_42941,N_36052,N_35051);
nand U42942 (N_42942,N_36526,N_39062);
and U42943 (N_42943,N_39411,N_35886);
nand U42944 (N_42944,N_36302,N_35883);
xnor U42945 (N_42945,N_36522,N_37824);
and U42946 (N_42946,N_38026,N_36543);
xnor U42947 (N_42947,N_37663,N_39680);
nand U42948 (N_42948,N_39829,N_37712);
and U42949 (N_42949,N_35593,N_36308);
nor U42950 (N_42950,N_36903,N_38777);
xor U42951 (N_42951,N_39502,N_38219);
xnor U42952 (N_42952,N_36950,N_39245);
xor U42953 (N_42953,N_37011,N_36783);
nor U42954 (N_42954,N_36964,N_35798);
and U42955 (N_42955,N_36764,N_38800);
nand U42956 (N_42956,N_36376,N_35299);
or U42957 (N_42957,N_37359,N_35584);
or U42958 (N_42958,N_35273,N_39982);
nand U42959 (N_42959,N_36965,N_39005);
nor U42960 (N_42960,N_38216,N_37268);
and U42961 (N_42961,N_38811,N_37884);
nor U42962 (N_42962,N_36584,N_38637);
nor U42963 (N_42963,N_36799,N_39207);
xor U42964 (N_42964,N_38709,N_36135);
and U42965 (N_42965,N_35623,N_35291);
nor U42966 (N_42966,N_37826,N_35423);
or U42967 (N_42967,N_38180,N_39022);
xnor U42968 (N_42968,N_38475,N_37367);
nor U42969 (N_42969,N_37061,N_37450);
or U42970 (N_42970,N_37097,N_37544);
nor U42971 (N_42971,N_35003,N_35261);
nand U42972 (N_42972,N_36734,N_38377);
nor U42973 (N_42973,N_35071,N_37116);
or U42974 (N_42974,N_37288,N_35706);
nand U42975 (N_42975,N_36726,N_35554);
nor U42976 (N_42976,N_35571,N_39693);
nor U42977 (N_42977,N_37726,N_36220);
nand U42978 (N_42978,N_37007,N_38496);
nor U42979 (N_42979,N_38852,N_35565);
xnor U42980 (N_42980,N_37207,N_36296);
xor U42981 (N_42981,N_36573,N_35063);
or U42982 (N_42982,N_36169,N_35866);
or U42983 (N_42983,N_37154,N_37893);
xnor U42984 (N_42984,N_36877,N_35167);
nand U42985 (N_42985,N_36797,N_37134);
nor U42986 (N_42986,N_36543,N_36463);
or U42987 (N_42987,N_35260,N_36956);
nor U42988 (N_42988,N_39819,N_35703);
nor U42989 (N_42989,N_38779,N_38843);
nor U42990 (N_42990,N_35638,N_37911);
nor U42991 (N_42991,N_37565,N_36925);
nor U42992 (N_42992,N_36727,N_38498);
xor U42993 (N_42993,N_36346,N_36845);
nor U42994 (N_42994,N_36746,N_36535);
nand U42995 (N_42995,N_37714,N_37156);
and U42996 (N_42996,N_38823,N_35586);
nand U42997 (N_42997,N_39857,N_35178);
nor U42998 (N_42998,N_37231,N_35204);
nand U42999 (N_42999,N_36348,N_38537);
and U43000 (N_43000,N_38663,N_39954);
or U43001 (N_43001,N_35317,N_36866);
and U43002 (N_43002,N_37081,N_36448);
nand U43003 (N_43003,N_38501,N_39744);
or U43004 (N_43004,N_35312,N_38184);
and U43005 (N_43005,N_35770,N_35593);
nand U43006 (N_43006,N_37530,N_38491);
or U43007 (N_43007,N_36320,N_37823);
nor U43008 (N_43008,N_36725,N_35836);
nand U43009 (N_43009,N_38279,N_37617);
nor U43010 (N_43010,N_37987,N_38334);
or U43011 (N_43011,N_35669,N_37113);
and U43012 (N_43012,N_36444,N_38704);
nor U43013 (N_43013,N_38410,N_36239);
xnor U43014 (N_43014,N_35597,N_38928);
nor U43015 (N_43015,N_35663,N_37216);
and U43016 (N_43016,N_36817,N_37588);
nor U43017 (N_43017,N_36381,N_38450);
and U43018 (N_43018,N_37055,N_39363);
or U43019 (N_43019,N_39851,N_35525);
xnor U43020 (N_43020,N_35360,N_37022);
or U43021 (N_43021,N_39197,N_37338);
and U43022 (N_43022,N_35138,N_38759);
and U43023 (N_43023,N_35914,N_37908);
and U43024 (N_43024,N_38854,N_35661);
xor U43025 (N_43025,N_39713,N_39349);
and U43026 (N_43026,N_38203,N_39557);
nor U43027 (N_43027,N_37213,N_38803);
nor U43028 (N_43028,N_36502,N_35251);
and U43029 (N_43029,N_36302,N_37873);
nor U43030 (N_43030,N_36117,N_39478);
xor U43031 (N_43031,N_39689,N_36402);
xnor U43032 (N_43032,N_37187,N_36664);
or U43033 (N_43033,N_36089,N_35225);
nand U43034 (N_43034,N_37303,N_38958);
and U43035 (N_43035,N_38605,N_37515);
or U43036 (N_43036,N_36148,N_36691);
and U43037 (N_43037,N_38639,N_38394);
nor U43038 (N_43038,N_35815,N_36853);
xor U43039 (N_43039,N_39749,N_35957);
nand U43040 (N_43040,N_37764,N_36701);
nand U43041 (N_43041,N_39229,N_38764);
nand U43042 (N_43042,N_35572,N_36781);
and U43043 (N_43043,N_36142,N_39894);
and U43044 (N_43044,N_37033,N_36276);
xnor U43045 (N_43045,N_39623,N_39983);
nand U43046 (N_43046,N_38190,N_36896);
nor U43047 (N_43047,N_35573,N_35018);
and U43048 (N_43048,N_37851,N_35775);
nor U43049 (N_43049,N_35373,N_36047);
or U43050 (N_43050,N_35446,N_38124);
and U43051 (N_43051,N_37504,N_35778);
and U43052 (N_43052,N_37402,N_36433);
nand U43053 (N_43053,N_37183,N_39092);
nand U43054 (N_43054,N_35388,N_35163);
xor U43055 (N_43055,N_38309,N_39874);
nand U43056 (N_43056,N_37144,N_35460);
xnor U43057 (N_43057,N_37869,N_38403);
nor U43058 (N_43058,N_39121,N_36842);
nand U43059 (N_43059,N_35960,N_39806);
xnor U43060 (N_43060,N_38718,N_39953);
or U43061 (N_43061,N_35170,N_35680);
nor U43062 (N_43062,N_36769,N_36192);
nor U43063 (N_43063,N_37335,N_35479);
nand U43064 (N_43064,N_39616,N_36788);
nand U43065 (N_43065,N_35243,N_35410);
nand U43066 (N_43066,N_35656,N_37047);
xnor U43067 (N_43067,N_37132,N_37788);
nor U43068 (N_43068,N_36522,N_36482);
xnor U43069 (N_43069,N_38335,N_39561);
and U43070 (N_43070,N_35867,N_39297);
xor U43071 (N_43071,N_37582,N_38242);
and U43072 (N_43072,N_39154,N_36807);
nand U43073 (N_43073,N_38209,N_39223);
or U43074 (N_43074,N_38783,N_39462);
nand U43075 (N_43075,N_36019,N_36383);
and U43076 (N_43076,N_38248,N_38667);
xor U43077 (N_43077,N_37546,N_37830);
nand U43078 (N_43078,N_39085,N_36235);
nand U43079 (N_43079,N_35067,N_37404);
nor U43080 (N_43080,N_36281,N_38368);
or U43081 (N_43081,N_36441,N_39631);
nor U43082 (N_43082,N_37266,N_37697);
nand U43083 (N_43083,N_37929,N_38859);
xnor U43084 (N_43084,N_38446,N_38639);
nand U43085 (N_43085,N_38264,N_35993);
xnor U43086 (N_43086,N_37802,N_35952);
and U43087 (N_43087,N_36924,N_37634);
and U43088 (N_43088,N_36023,N_39363);
nor U43089 (N_43089,N_38021,N_38911);
nand U43090 (N_43090,N_38492,N_35167);
nor U43091 (N_43091,N_37241,N_36603);
nand U43092 (N_43092,N_35421,N_35734);
nor U43093 (N_43093,N_38561,N_39200);
xor U43094 (N_43094,N_38430,N_39403);
or U43095 (N_43095,N_37872,N_36408);
and U43096 (N_43096,N_39559,N_35790);
xor U43097 (N_43097,N_39200,N_37107);
or U43098 (N_43098,N_36268,N_39835);
or U43099 (N_43099,N_37532,N_35735);
nor U43100 (N_43100,N_36246,N_39576);
and U43101 (N_43101,N_36020,N_39782);
or U43102 (N_43102,N_37734,N_36578);
and U43103 (N_43103,N_38793,N_38478);
or U43104 (N_43104,N_35652,N_36611);
xnor U43105 (N_43105,N_35125,N_37492);
nand U43106 (N_43106,N_36051,N_39500);
nor U43107 (N_43107,N_37249,N_39388);
nand U43108 (N_43108,N_37086,N_39942);
xnor U43109 (N_43109,N_39399,N_38339);
xor U43110 (N_43110,N_39999,N_35097);
or U43111 (N_43111,N_35293,N_37716);
or U43112 (N_43112,N_39030,N_37281);
or U43113 (N_43113,N_38516,N_37319);
nor U43114 (N_43114,N_35652,N_37525);
nand U43115 (N_43115,N_37282,N_36671);
or U43116 (N_43116,N_35590,N_36730);
and U43117 (N_43117,N_38517,N_37266);
nand U43118 (N_43118,N_38231,N_35949);
nor U43119 (N_43119,N_39654,N_39402);
nand U43120 (N_43120,N_35386,N_35003);
or U43121 (N_43121,N_39594,N_39293);
and U43122 (N_43122,N_36482,N_36572);
nand U43123 (N_43123,N_38926,N_38373);
nor U43124 (N_43124,N_37709,N_38104);
xnor U43125 (N_43125,N_37239,N_37946);
and U43126 (N_43126,N_36175,N_35727);
or U43127 (N_43127,N_39686,N_36214);
or U43128 (N_43128,N_36482,N_35074);
and U43129 (N_43129,N_35098,N_39829);
and U43130 (N_43130,N_39816,N_39480);
nand U43131 (N_43131,N_36298,N_35158);
and U43132 (N_43132,N_39775,N_38271);
nand U43133 (N_43133,N_37831,N_36062);
or U43134 (N_43134,N_37004,N_35776);
or U43135 (N_43135,N_38082,N_38094);
or U43136 (N_43136,N_39739,N_38185);
nand U43137 (N_43137,N_36529,N_35370);
xor U43138 (N_43138,N_35978,N_35713);
and U43139 (N_43139,N_39683,N_37242);
nor U43140 (N_43140,N_38358,N_35160);
or U43141 (N_43141,N_35788,N_39987);
nor U43142 (N_43142,N_38735,N_39626);
xnor U43143 (N_43143,N_39827,N_39959);
xnor U43144 (N_43144,N_35122,N_36841);
nand U43145 (N_43145,N_39771,N_39219);
and U43146 (N_43146,N_37780,N_37367);
nor U43147 (N_43147,N_39927,N_37947);
and U43148 (N_43148,N_38180,N_36095);
or U43149 (N_43149,N_36025,N_36324);
and U43150 (N_43150,N_39626,N_37048);
nand U43151 (N_43151,N_36381,N_38016);
nand U43152 (N_43152,N_38157,N_38760);
nand U43153 (N_43153,N_38456,N_38243);
nor U43154 (N_43154,N_35287,N_36710);
or U43155 (N_43155,N_38414,N_36311);
xnor U43156 (N_43156,N_36495,N_39487);
xor U43157 (N_43157,N_36808,N_39465);
nand U43158 (N_43158,N_39041,N_39165);
nand U43159 (N_43159,N_37157,N_38799);
nand U43160 (N_43160,N_35170,N_39550);
and U43161 (N_43161,N_37164,N_38698);
nand U43162 (N_43162,N_37041,N_38266);
or U43163 (N_43163,N_37028,N_37533);
xnor U43164 (N_43164,N_38115,N_37618);
or U43165 (N_43165,N_37154,N_38503);
nor U43166 (N_43166,N_38600,N_35934);
or U43167 (N_43167,N_36196,N_35012);
or U43168 (N_43168,N_35867,N_35235);
and U43169 (N_43169,N_36281,N_37440);
nor U43170 (N_43170,N_38043,N_35478);
nor U43171 (N_43171,N_38612,N_35017);
nand U43172 (N_43172,N_39272,N_38521);
or U43173 (N_43173,N_36252,N_36574);
and U43174 (N_43174,N_37205,N_36055);
nand U43175 (N_43175,N_35369,N_35086);
xor U43176 (N_43176,N_35053,N_37205);
nand U43177 (N_43177,N_36905,N_35010);
nor U43178 (N_43178,N_35961,N_38283);
nand U43179 (N_43179,N_39191,N_39650);
nand U43180 (N_43180,N_39712,N_37757);
nand U43181 (N_43181,N_36788,N_35501);
nor U43182 (N_43182,N_39356,N_35559);
xnor U43183 (N_43183,N_39583,N_36551);
xor U43184 (N_43184,N_39050,N_38043);
nor U43185 (N_43185,N_38857,N_37943);
or U43186 (N_43186,N_37468,N_38714);
or U43187 (N_43187,N_39798,N_37138);
nand U43188 (N_43188,N_37105,N_35227);
and U43189 (N_43189,N_38280,N_37792);
and U43190 (N_43190,N_38131,N_38982);
nand U43191 (N_43191,N_35400,N_38643);
or U43192 (N_43192,N_37920,N_35210);
nand U43193 (N_43193,N_36566,N_35327);
xnor U43194 (N_43194,N_35868,N_38900);
and U43195 (N_43195,N_39853,N_38485);
nand U43196 (N_43196,N_39387,N_37600);
nand U43197 (N_43197,N_35331,N_36837);
and U43198 (N_43198,N_36921,N_37316);
nor U43199 (N_43199,N_37864,N_36963);
nand U43200 (N_43200,N_37918,N_39348);
or U43201 (N_43201,N_37025,N_35412);
nand U43202 (N_43202,N_37012,N_36386);
xor U43203 (N_43203,N_37936,N_38833);
and U43204 (N_43204,N_39706,N_39742);
or U43205 (N_43205,N_39602,N_35765);
nand U43206 (N_43206,N_39175,N_38164);
nand U43207 (N_43207,N_37729,N_38899);
nand U43208 (N_43208,N_39904,N_37365);
and U43209 (N_43209,N_37981,N_36595);
xnor U43210 (N_43210,N_38751,N_39067);
or U43211 (N_43211,N_37573,N_39978);
nand U43212 (N_43212,N_36276,N_37931);
nand U43213 (N_43213,N_39678,N_37882);
nand U43214 (N_43214,N_39120,N_36130);
or U43215 (N_43215,N_37374,N_35409);
and U43216 (N_43216,N_36509,N_38707);
and U43217 (N_43217,N_35515,N_36594);
or U43218 (N_43218,N_37735,N_37203);
xor U43219 (N_43219,N_39148,N_35822);
nor U43220 (N_43220,N_37492,N_35088);
nand U43221 (N_43221,N_36849,N_38662);
xor U43222 (N_43222,N_36973,N_39849);
xor U43223 (N_43223,N_36390,N_38942);
nand U43224 (N_43224,N_36323,N_37268);
nor U43225 (N_43225,N_35019,N_37776);
and U43226 (N_43226,N_39826,N_35204);
and U43227 (N_43227,N_38514,N_37471);
nor U43228 (N_43228,N_36063,N_39764);
or U43229 (N_43229,N_36398,N_37901);
or U43230 (N_43230,N_37565,N_35479);
nand U43231 (N_43231,N_38927,N_35397);
nand U43232 (N_43232,N_36033,N_35644);
xor U43233 (N_43233,N_38648,N_35824);
nand U43234 (N_43234,N_37436,N_35546);
nand U43235 (N_43235,N_39838,N_39092);
or U43236 (N_43236,N_36861,N_38426);
or U43237 (N_43237,N_38383,N_38223);
and U43238 (N_43238,N_36411,N_35054);
xor U43239 (N_43239,N_35268,N_38747);
xor U43240 (N_43240,N_37336,N_36607);
nor U43241 (N_43241,N_35060,N_37093);
or U43242 (N_43242,N_36204,N_36193);
nand U43243 (N_43243,N_37314,N_38003);
or U43244 (N_43244,N_36053,N_37223);
or U43245 (N_43245,N_35263,N_37203);
nand U43246 (N_43246,N_37112,N_39157);
nand U43247 (N_43247,N_39748,N_39202);
nor U43248 (N_43248,N_39904,N_37062);
xor U43249 (N_43249,N_39167,N_35317);
and U43250 (N_43250,N_37505,N_38464);
nand U43251 (N_43251,N_35870,N_35215);
nand U43252 (N_43252,N_39904,N_36990);
nor U43253 (N_43253,N_39029,N_37450);
xor U43254 (N_43254,N_35408,N_38074);
or U43255 (N_43255,N_39122,N_37671);
nor U43256 (N_43256,N_39419,N_36838);
or U43257 (N_43257,N_35642,N_39507);
and U43258 (N_43258,N_36288,N_36871);
or U43259 (N_43259,N_39626,N_37008);
nand U43260 (N_43260,N_37988,N_35621);
or U43261 (N_43261,N_39697,N_38629);
or U43262 (N_43262,N_35972,N_36755);
or U43263 (N_43263,N_35515,N_39210);
nor U43264 (N_43264,N_35815,N_35769);
and U43265 (N_43265,N_35604,N_39479);
and U43266 (N_43266,N_38788,N_38982);
or U43267 (N_43267,N_37918,N_36013);
nor U43268 (N_43268,N_39624,N_38742);
nand U43269 (N_43269,N_38291,N_36771);
or U43270 (N_43270,N_38471,N_36981);
xor U43271 (N_43271,N_38603,N_38881);
xor U43272 (N_43272,N_35813,N_36232);
nand U43273 (N_43273,N_36185,N_38225);
xnor U43274 (N_43274,N_35618,N_39431);
nor U43275 (N_43275,N_37672,N_39682);
nand U43276 (N_43276,N_35540,N_38602);
and U43277 (N_43277,N_35638,N_39875);
xnor U43278 (N_43278,N_35089,N_35461);
xnor U43279 (N_43279,N_37348,N_35441);
nor U43280 (N_43280,N_35126,N_37878);
nor U43281 (N_43281,N_35354,N_35500);
and U43282 (N_43282,N_36492,N_37328);
xor U43283 (N_43283,N_37105,N_39122);
or U43284 (N_43284,N_38309,N_39913);
nand U43285 (N_43285,N_35159,N_38965);
or U43286 (N_43286,N_39355,N_37941);
nand U43287 (N_43287,N_36792,N_35373);
xor U43288 (N_43288,N_39024,N_39365);
nor U43289 (N_43289,N_39096,N_36314);
nand U43290 (N_43290,N_37233,N_36103);
xnor U43291 (N_43291,N_36742,N_37367);
nand U43292 (N_43292,N_37571,N_35302);
and U43293 (N_43293,N_39385,N_35072);
nor U43294 (N_43294,N_35662,N_36165);
xor U43295 (N_43295,N_38567,N_35115);
and U43296 (N_43296,N_39171,N_37236);
xnor U43297 (N_43297,N_38370,N_38871);
xor U43298 (N_43298,N_35823,N_37970);
or U43299 (N_43299,N_35456,N_39751);
nor U43300 (N_43300,N_37172,N_38482);
or U43301 (N_43301,N_39787,N_35117);
or U43302 (N_43302,N_38180,N_36536);
xor U43303 (N_43303,N_38590,N_35456);
nor U43304 (N_43304,N_39572,N_38755);
nand U43305 (N_43305,N_37323,N_37123);
xnor U43306 (N_43306,N_38677,N_35021);
and U43307 (N_43307,N_38165,N_35287);
and U43308 (N_43308,N_35233,N_36399);
and U43309 (N_43309,N_37001,N_39159);
xnor U43310 (N_43310,N_38004,N_38689);
nor U43311 (N_43311,N_39750,N_37333);
nand U43312 (N_43312,N_37515,N_37934);
xor U43313 (N_43313,N_39445,N_38615);
nor U43314 (N_43314,N_35323,N_37668);
nand U43315 (N_43315,N_38080,N_37780);
or U43316 (N_43316,N_35033,N_35762);
xor U43317 (N_43317,N_39340,N_35655);
xor U43318 (N_43318,N_37703,N_39469);
nor U43319 (N_43319,N_35760,N_38892);
nor U43320 (N_43320,N_36194,N_36643);
or U43321 (N_43321,N_39800,N_37392);
or U43322 (N_43322,N_35180,N_38329);
or U43323 (N_43323,N_37282,N_37907);
nand U43324 (N_43324,N_39394,N_36488);
and U43325 (N_43325,N_35480,N_36186);
or U43326 (N_43326,N_35736,N_37484);
or U43327 (N_43327,N_39667,N_36037);
nor U43328 (N_43328,N_36138,N_38553);
nand U43329 (N_43329,N_36246,N_39677);
xnor U43330 (N_43330,N_36351,N_39387);
and U43331 (N_43331,N_38044,N_39137);
nand U43332 (N_43332,N_35631,N_35234);
or U43333 (N_43333,N_38271,N_35499);
nor U43334 (N_43334,N_38949,N_35410);
xor U43335 (N_43335,N_38010,N_38940);
nand U43336 (N_43336,N_38097,N_36637);
nand U43337 (N_43337,N_39029,N_39531);
nor U43338 (N_43338,N_35047,N_37809);
and U43339 (N_43339,N_36473,N_37185);
nor U43340 (N_43340,N_37099,N_38010);
nor U43341 (N_43341,N_35274,N_39775);
or U43342 (N_43342,N_39936,N_39879);
nor U43343 (N_43343,N_36085,N_38561);
xor U43344 (N_43344,N_35467,N_38807);
xnor U43345 (N_43345,N_36583,N_38655);
and U43346 (N_43346,N_39834,N_36287);
xor U43347 (N_43347,N_36575,N_39548);
and U43348 (N_43348,N_39284,N_37059);
nor U43349 (N_43349,N_38260,N_37937);
nand U43350 (N_43350,N_37450,N_36996);
or U43351 (N_43351,N_36745,N_36686);
and U43352 (N_43352,N_36801,N_39581);
and U43353 (N_43353,N_39693,N_38776);
or U43354 (N_43354,N_39621,N_38050);
or U43355 (N_43355,N_38148,N_37433);
or U43356 (N_43356,N_39223,N_39893);
and U43357 (N_43357,N_36439,N_35966);
xnor U43358 (N_43358,N_35678,N_35545);
or U43359 (N_43359,N_36358,N_37872);
nor U43360 (N_43360,N_37778,N_37708);
and U43361 (N_43361,N_39492,N_37508);
nand U43362 (N_43362,N_37750,N_38358);
or U43363 (N_43363,N_37328,N_35073);
and U43364 (N_43364,N_37401,N_37467);
nand U43365 (N_43365,N_38841,N_38850);
xnor U43366 (N_43366,N_39987,N_36146);
or U43367 (N_43367,N_35476,N_36523);
nand U43368 (N_43368,N_36700,N_37594);
nand U43369 (N_43369,N_38417,N_35172);
xor U43370 (N_43370,N_39642,N_37580);
nand U43371 (N_43371,N_37034,N_37792);
or U43372 (N_43372,N_35426,N_35671);
xor U43373 (N_43373,N_35787,N_37782);
or U43374 (N_43374,N_38513,N_37988);
and U43375 (N_43375,N_36452,N_37691);
and U43376 (N_43376,N_39813,N_37814);
and U43377 (N_43377,N_37343,N_38421);
xor U43378 (N_43378,N_37501,N_39611);
and U43379 (N_43379,N_38301,N_39125);
xor U43380 (N_43380,N_36937,N_39183);
nand U43381 (N_43381,N_39641,N_39509);
nand U43382 (N_43382,N_39965,N_39773);
nor U43383 (N_43383,N_37790,N_37208);
xnor U43384 (N_43384,N_38667,N_35620);
nor U43385 (N_43385,N_39256,N_39860);
nand U43386 (N_43386,N_36945,N_38738);
or U43387 (N_43387,N_38457,N_38641);
nor U43388 (N_43388,N_39376,N_38237);
or U43389 (N_43389,N_37777,N_36086);
nor U43390 (N_43390,N_39903,N_36948);
nor U43391 (N_43391,N_38664,N_39080);
nor U43392 (N_43392,N_35714,N_38050);
and U43393 (N_43393,N_36402,N_39989);
or U43394 (N_43394,N_37912,N_38412);
and U43395 (N_43395,N_39342,N_39300);
xor U43396 (N_43396,N_36374,N_39909);
or U43397 (N_43397,N_38399,N_36760);
or U43398 (N_43398,N_36426,N_35616);
or U43399 (N_43399,N_36443,N_38840);
nand U43400 (N_43400,N_39844,N_37466);
or U43401 (N_43401,N_39147,N_38498);
and U43402 (N_43402,N_39086,N_35997);
or U43403 (N_43403,N_39664,N_36888);
or U43404 (N_43404,N_36192,N_35567);
xor U43405 (N_43405,N_36967,N_39696);
xnor U43406 (N_43406,N_39657,N_38157);
xor U43407 (N_43407,N_37555,N_38770);
and U43408 (N_43408,N_37195,N_38028);
and U43409 (N_43409,N_37267,N_39693);
nor U43410 (N_43410,N_37741,N_37101);
xor U43411 (N_43411,N_36011,N_39162);
nor U43412 (N_43412,N_38807,N_38020);
or U43413 (N_43413,N_37301,N_37149);
xor U43414 (N_43414,N_39987,N_39751);
nand U43415 (N_43415,N_37244,N_38656);
xnor U43416 (N_43416,N_39056,N_36029);
nand U43417 (N_43417,N_36821,N_35103);
or U43418 (N_43418,N_37204,N_35559);
or U43419 (N_43419,N_35317,N_35161);
nor U43420 (N_43420,N_37992,N_39882);
nand U43421 (N_43421,N_36194,N_36044);
xnor U43422 (N_43422,N_38208,N_37511);
nand U43423 (N_43423,N_36268,N_35649);
nor U43424 (N_43424,N_37994,N_38419);
nor U43425 (N_43425,N_35647,N_38667);
or U43426 (N_43426,N_36331,N_36211);
xnor U43427 (N_43427,N_36292,N_38756);
nand U43428 (N_43428,N_37977,N_38520);
or U43429 (N_43429,N_39045,N_37687);
and U43430 (N_43430,N_39287,N_35053);
nand U43431 (N_43431,N_38152,N_35629);
nor U43432 (N_43432,N_37420,N_36037);
or U43433 (N_43433,N_35710,N_35506);
or U43434 (N_43434,N_39221,N_39315);
xor U43435 (N_43435,N_36408,N_37974);
nor U43436 (N_43436,N_38233,N_38194);
and U43437 (N_43437,N_36796,N_37943);
nand U43438 (N_43438,N_39619,N_37946);
nor U43439 (N_43439,N_37158,N_37378);
xnor U43440 (N_43440,N_37811,N_39981);
nand U43441 (N_43441,N_39955,N_35437);
nor U43442 (N_43442,N_39624,N_36624);
nand U43443 (N_43443,N_36232,N_38257);
nor U43444 (N_43444,N_35501,N_38555);
and U43445 (N_43445,N_38925,N_38712);
nor U43446 (N_43446,N_38752,N_35634);
nor U43447 (N_43447,N_38116,N_36497);
nor U43448 (N_43448,N_35171,N_38275);
nor U43449 (N_43449,N_39027,N_38614);
nand U43450 (N_43450,N_38317,N_37197);
xor U43451 (N_43451,N_37360,N_37089);
xor U43452 (N_43452,N_36558,N_35671);
nand U43453 (N_43453,N_39650,N_38940);
or U43454 (N_43454,N_35239,N_38307);
xnor U43455 (N_43455,N_37611,N_35150);
or U43456 (N_43456,N_37372,N_37132);
xnor U43457 (N_43457,N_37180,N_35741);
nor U43458 (N_43458,N_35701,N_35738);
and U43459 (N_43459,N_38418,N_36172);
and U43460 (N_43460,N_39026,N_39910);
or U43461 (N_43461,N_36345,N_36517);
nand U43462 (N_43462,N_37804,N_37493);
or U43463 (N_43463,N_39712,N_37894);
xor U43464 (N_43464,N_36736,N_35344);
and U43465 (N_43465,N_38215,N_37251);
or U43466 (N_43466,N_38345,N_39140);
or U43467 (N_43467,N_36012,N_38853);
nor U43468 (N_43468,N_39447,N_39077);
nor U43469 (N_43469,N_38793,N_36486);
nand U43470 (N_43470,N_37911,N_39929);
nor U43471 (N_43471,N_38709,N_36239);
and U43472 (N_43472,N_35525,N_38825);
nor U43473 (N_43473,N_36878,N_37524);
or U43474 (N_43474,N_35042,N_35602);
nand U43475 (N_43475,N_36683,N_36197);
or U43476 (N_43476,N_36038,N_36921);
nor U43477 (N_43477,N_35337,N_36901);
and U43478 (N_43478,N_35375,N_37547);
nand U43479 (N_43479,N_36264,N_35453);
xor U43480 (N_43480,N_37918,N_37870);
xnor U43481 (N_43481,N_35323,N_35705);
xor U43482 (N_43482,N_36767,N_37547);
or U43483 (N_43483,N_35620,N_38332);
nand U43484 (N_43484,N_39152,N_38950);
nor U43485 (N_43485,N_35632,N_38896);
xnor U43486 (N_43486,N_35496,N_35197);
xor U43487 (N_43487,N_38058,N_36657);
nor U43488 (N_43488,N_39712,N_36763);
and U43489 (N_43489,N_39041,N_36181);
xor U43490 (N_43490,N_37468,N_38798);
and U43491 (N_43491,N_39336,N_35722);
xnor U43492 (N_43492,N_35723,N_37511);
xor U43493 (N_43493,N_36388,N_37434);
xor U43494 (N_43494,N_36155,N_35846);
xnor U43495 (N_43495,N_39936,N_36358);
xnor U43496 (N_43496,N_39880,N_37242);
nand U43497 (N_43497,N_38323,N_36011);
nand U43498 (N_43498,N_39307,N_37943);
and U43499 (N_43499,N_38341,N_36225);
or U43500 (N_43500,N_38891,N_35075);
and U43501 (N_43501,N_35703,N_37761);
nor U43502 (N_43502,N_35366,N_36512);
nand U43503 (N_43503,N_36127,N_36759);
nand U43504 (N_43504,N_37614,N_36122);
nand U43505 (N_43505,N_38246,N_39932);
xnor U43506 (N_43506,N_36939,N_36956);
xnor U43507 (N_43507,N_38558,N_36459);
and U43508 (N_43508,N_37812,N_38887);
nand U43509 (N_43509,N_38203,N_37523);
xnor U43510 (N_43510,N_37992,N_39947);
or U43511 (N_43511,N_37485,N_37461);
and U43512 (N_43512,N_37072,N_38877);
nor U43513 (N_43513,N_39037,N_35054);
or U43514 (N_43514,N_38069,N_38335);
nand U43515 (N_43515,N_39847,N_37896);
and U43516 (N_43516,N_36962,N_39503);
nor U43517 (N_43517,N_38972,N_38678);
nand U43518 (N_43518,N_37157,N_35866);
and U43519 (N_43519,N_35723,N_38609);
and U43520 (N_43520,N_35615,N_35916);
xor U43521 (N_43521,N_35886,N_37319);
nor U43522 (N_43522,N_37341,N_38566);
and U43523 (N_43523,N_38624,N_39836);
xnor U43524 (N_43524,N_38402,N_38556);
xor U43525 (N_43525,N_39210,N_37368);
or U43526 (N_43526,N_36212,N_36026);
nor U43527 (N_43527,N_36432,N_39792);
xor U43528 (N_43528,N_35771,N_35624);
nor U43529 (N_43529,N_35617,N_36993);
or U43530 (N_43530,N_37035,N_35246);
and U43531 (N_43531,N_39916,N_38363);
or U43532 (N_43532,N_36505,N_35124);
or U43533 (N_43533,N_37609,N_35968);
nand U43534 (N_43534,N_35087,N_35378);
nor U43535 (N_43535,N_38039,N_38179);
or U43536 (N_43536,N_39269,N_37833);
xnor U43537 (N_43537,N_39503,N_37039);
and U43538 (N_43538,N_36222,N_36064);
and U43539 (N_43539,N_37084,N_37614);
nor U43540 (N_43540,N_36033,N_35003);
xnor U43541 (N_43541,N_37530,N_39119);
or U43542 (N_43542,N_38069,N_37559);
and U43543 (N_43543,N_37665,N_35386);
nand U43544 (N_43544,N_35988,N_35724);
and U43545 (N_43545,N_39087,N_38002);
nand U43546 (N_43546,N_37386,N_36989);
nand U43547 (N_43547,N_39883,N_35519);
nand U43548 (N_43548,N_36368,N_35870);
nor U43549 (N_43549,N_36325,N_35359);
nor U43550 (N_43550,N_36385,N_39940);
nor U43551 (N_43551,N_36045,N_39190);
or U43552 (N_43552,N_39218,N_36992);
xor U43553 (N_43553,N_37864,N_39360);
and U43554 (N_43554,N_35436,N_35288);
or U43555 (N_43555,N_39611,N_37989);
or U43556 (N_43556,N_37732,N_37795);
xor U43557 (N_43557,N_37447,N_36457);
nor U43558 (N_43558,N_35826,N_39920);
nor U43559 (N_43559,N_37947,N_39373);
nor U43560 (N_43560,N_35740,N_35430);
nand U43561 (N_43561,N_39759,N_39221);
xnor U43562 (N_43562,N_39441,N_35190);
or U43563 (N_43563,N_35554,N_37099);
or U43564 (N_43564,N_39057,N_35919);
nand U43565 (N_43565,N_37638,N_37828);
xnor U43566 (N_43566,N_39307,N_39032);
and U43567 (N_43567,N_36972,N_38323);
or U43568 (N_43568,N_35313,N_38084);
nand U43569 (N_43569,N_35899,N_36037);
nor U43570 (N_43570,N_36801,N_38292);
or U43571 (N_43571,N_36875,N_37396);
or U43572 (N_43572,N_36219,N_36932);
nand U43573 (N_43573,N_39152,N_35385);
nor U43574 (N_43574,N_38740,N_36116);
and U43575 (N_43575,N_39624,N_37137);
xnor U43576 (N_43576,N_37035,N_39896);
and U43577 (N_43577,N_36274,N_35257);
and U43578 (N_43578,N_36237,N_39182);
xor U43579 (N_43579,N_35191,N_39402);
nand U43580 (N_43580,N_37404,N_38808);
and U43581 (N_43581,N_38377,N_36609);
and U43582 (N_43582,N_37211,N_35289);
and U43583 (N_43583,N_36973,N_38152);
or U43584 (N_43584,N_38785,N_37182);
nand U43585 (N_43585,N_39384,N_39696);
nor U43586 (N_43586,N_38145,N_35740);
and U43587 (N_43587,N_38485,N_37802);
or U43588 (N_43588,N_35577,N_36875);
nor U43589 (N_43589,N_35958,N_38770);
xnor U43590 (N_43590,N_35277,N_39631);
and U43591 (N_43591,N_36320,N_36758);
or U43592 (N_43592,N_39001,N_38070);
nand U43593 (N_43593,N_37408,N_37409);
and U43594 (N_43594,N_36872,N_37041);
or U43595 (N_43595,N_38643,N_35904);
nand U43596 (N_43596,N_38801,N_38019);
nand U43597 (N_43597,N_39402,N_36400);
nand U43598 (N_43598,N_39946,N_35847);
or U43599 (N_43599,N_35934,N_35197);
nand U43600 (N_43600,N_36771,N_35788);
and U43601 (N_43601,N_35614,N_36886);
xnor U43602 (N_43602,N_37253,N_38709);
or U43603 (N_43603,N_38353,N_38104);
xnor U43604 (N_43604,N_35634,N_36893);
or U43605 (N_43605,N_37042,N_35283);
xor U43606 (N_43606,N_35329,N_37447);
xnor U43607 (N_43607,N_35296,N_36645);
xor U43608 (N_43608,N_39764,N_36981);
nor U43609 (N_43609,N_37898,N_38840);
and U43610 (N_43610,N_35735,N_35516);
xor U43611 (N_43611,N_37075,N_35734);
xnor U43612 (N_43612,N_39955,N_35720);
or U43613 (N_43613,N_37682,N_38998);
nor U43614 (N_43614,N_38660,N_39430);
nor U43615 (N_43615,N_39746,N_35166);
nand U43616 (N_43616,N_38503,N_38105);
nor U43617 (N_43617,N_39600,N_39965);
nand U43618 (N_43618,N_35199,N_39220);
nor U43619 (N_43619,N_36334,N_37531);
or U43620 (N_43620,N_36446,N_35366);
nand U43621 (N_43621,N_35703,N_37254);
and U43622 (N_43622,N_38141,N_35063);
nor U43623 (N_43623,N_38383,N_36954);
or U43624 (N_43624,N_36949,N_37670);
or U43625 (N_43625,N_36977,N_37212);
xor U43626 (N_43626,N_38504,N_35647);
and U43627 (N_43627,N_37334,N_36190);
nand U43628 (N_43628,N_39035,N_37342);
or U43629 (N_43629,N_36096,N_38074);
nor U43630 (N_43630,N_38087,N_37867);
nand U43631 (N_43631,N_39453,N_36489);
or U43632 (N_43632,N_35754,N_38838);
xor U43633 (N_43633,N_38644,N_38599);
nor U43634 (N_43634,N_38342,N_36752);
nand U43635 (N_43635,N_39288,N_37633);
nand U43636 (N_43636,N_39482,N_38076);
and U43637 (N_43637,N_37710,N_37706);
or U43638 (N_43638,N_39074,N_36789);
or U43639 (N_43639,N_37431,N_37463);
nand U43640 (N_43640,N_36959,N_39573);
nor U43641 (N_43641,N_36514,N_36755);
and U43642 (N_43642,N_37388,N_39897);
nand U43643 (N_43643,N_37869,N_35335);
or U43644 (N_43644,N_37646,N_38859);
nand U43645 (N_43645,N_37815,N_37402);
or U43646 (N_43646,N_37335,N_39113);
and U43647 (N_43647,N_36153,N_37547);
or U43648 (N_43648,N_39482,N_35344);
nand U43649 (N_43649,N_39164,N_35212);
and U43650 (N_43650,N_37931,N_39836);
xnor U43651 (N_43651,N_38477,N_35363);
nor U43652 (N_43652,N_35412,N_39380);
nand U43653 (N_43653,N_39643,N_39073);
xor U43654 (N_43654,N_39545,N_37392);
nand U43655 (N_43655,N_36743,N_39605);
nand U43656 (N_43656,N_37502,N_39881);
nor U43657 (N_43657,N_36300,N_36499);
nand U43658 (N_43658,N_38558,N_36742);
nand U43659 (N_43659,N_37998,N_35439);
nor U43660 (N_43660,N_38394,N_38365);
nor U43661 (N_43661,N_39610,N_37778);
xnor U43662 (N_43662,N_35864,N_39388);
or U43663 (N_43663,N_38769,N_36702);
or U43664 (N_43664,N_39028,N_37068);
nor U43665 (N_43665,N_37966,N_38459);
or U43666 (N_43666,N_37583,N_39046);
and U43667 (N_43667,N_38755,N_37955);
nor U43668 (N_43668,N_36390,N_37775);
and U43669 (N_43669,N_39227,N_37901);
nand U43670 (N_43670,N_35487,N_37110);
or U43671 (N_43671,N_37608,N_36188);
nand U43672 (N_43672,N_38747,N_35256);
nor U43673 (N_43673,N_38324,N_36678);
nand U43674 (N_43674,N_38286,N_38545);
xnor U43675 (N_43675,N_36566,N_37313);
or U43676 (N_43676,N_38976,N_38981);
xor U43677 (N_43677,N_39465,N_37213);
nand U43678 (N_43678,N_35040,N_39496);
nor U43679 (N_43679,N_35998,N_38055);
nand U43680 (N_43680,N_36214,N_39662);
nor U43681 (N_43681,N_36189,N_35176);
nor U43682 (N_43682,N_36563,N_39766);
or U43683 (N_43683,N_37170,N_39687);
xor U43684 (N_43684,N_39706,N_39195);
nand U43685 (N_43685,N_38843,N_36507);
nor U43686 (N_43686,N_39426,N_36804);
or U43687 (N_43687,N_38613,N_39592);
nand U43688 (N_43688,N_37652,N_38065);
or U43689 (N_43689,N_35147,N_36196);
and U43690 (N_43690,N_37784,N_37501);
nor U43691 (N_43691,N_39880,N_37434);
nor U43692 (N_43692,N_38725,N_39965);
or U43693 (N_43693,N_35606,N_39708);
and U43694 (N_43694,N_35249,N_38872);
nor U43695 (N_43695,N_37469,N_36117);
xnor U43696 (N_43696,N_36842,N_39804);
or U43697 (N_43697,N_35198,N_38444);
xor U43698 (N_43698,N_38377,N_38974);
or U43699 (N_43699,N_36955,N_36157);
and U43700 (N_43700,N_37328,N_35938);
nand U43701 (N_43701,N_38520,N_36823);
xnor U43702 (N_43702,N_35781,N_37915);
and U43703 (N_43703,N_37898,N_35431);
and U43704 (N_43704,N_39782,N_36871);
xnor U43705 (N_43705,N_37089,N_38247);
xor U43706 (N_43706,N_38057,N_35131);
or U43707 (N_43707,N_38239,N_37915);
nand U43708 (N_43708,N_36554,N_39686);
xor U43709 (N_43709,N_39938,N_37082);
and U43710 (N_43710,N_37035,N_38582);
nand U43711 (N_43711,N_39388,N_38244);
or U43712 (N_43712,N_37698,N_38961);
nor U43713 (N_43713,N_38724,N_39054);
xor U43714 (N_43714,N_38866,N_39718);
or U43715 (N_43715,N_38569,N_36600);
nand U43716 (N_43716,N_38625,N_35008);
xnor U43717 (N_43717,N_38590,N_39217);
xnor U43718 (N_43718,N_39395,N_37549);
or U43719 (N_43719,N_35765,N_39146);
or U43720 (N_43720,N_36134,N_38377);
nand U43721 (N_43721,N_35816,N_35169);
nor U43722 (N_43722,N_36050,N_35815);
nand U43723 (N_43723,N_39477,N_38531);
nor U43724 (N_43724,N_36379,N_38399);
and U43725 (N_43725,N_35511,N_37383);
xnor U43726 (N_43726,N_35742,N_37696);
and U43727 (N_43727,N_36342,N_35326);
nand U43728 (N_43728,N_36234,N_36476);
xnor U43729 (N_43729,N_35009,N_35564);
and U43730 (N_43730,N_37000,N_39551);
nand U43731 (N_43731,N_35010,N_38484);
nor U43732 (N_43732,N_37432,N_35563);
nand U43733 (N_43733,N_39137,N_39327);
nor U43734 (N_43734,N_35790,N_39012);
and U43735 (N_43735,N_39541,N_38569);
xnor U43736 (N_43736,N_35306,N_37926);
or U43737 (N_43737,N_39641,N_36726);
xor U43738 (N_43738,N_39932,N_38262);
nand U43739 (N_43739,N_36510,N_39734);
and U43740 (N_43740,N_38224,N_35737);
nand U43741 (N_43741,N_38793,N_35942);
nand U43742 (N_43742,N_38552,N_36089);
nand U43743 (N_43743,N_38632,N_35356);
xnor U43744 (N_43744,N_35681,N_36216);
xor U43745 (N_43745,N_35596,N_37042);
xor U43746 (N_43746,N_36774,N_35309);
and U43747 (N_43747,N_39393,N_35883);
nand U43748 (N_43748,N_39086,N_36595);
nand U43749 (N_43749,N_35661,N_39989);
and U43750 (N_43750,N_37895,N_37928);
nor U43751 (N_43751,N_38841,N_38186);
xnor U43752 (N_43752,N_35806,N_38037);
and U43753 (N_43753,N_39820,N_36673);
or U43754 (N_43754,N_36206,N_36436);
xnor U43755 (N_43755,N_36110,N_35372);
nand U43756 (N_43756,N_39132,N_39044);
xnor U43757 (N_43757,N_38024,N_37685);
or U43758 (N_43758,N_37064,N_36318);
xor U43759 (N_43759,N_39621,N_35232);
or U43760 (N_43760,N_36308,N_39883);
and U43761 (N_43761,N_37242,N_36537);
nor U43762 (N_43762,N_35827,N_35418);
or U43763 (N_43763,N_36940,N_36755);
nand U43764 (N_43764,N_36099,N_38715);
and U43765 (N_43765,N_39031,N_37668);
nor U43766 (N_43766,N_37361,N_39982);
or U43767 (N_43767,N_35986,N_35098);
nor U43768 (N_43768,N_35508,N_35164);
nand U43769 (N_43769,N_39261,N_37598);
or U43770 (N_43770,N_39846,N_37209);
and U43771 (N_43771,N_39470,N_38177);
xor U43772 (N_43772,N_37729,N_35244);
and U43773 (N_43773,N_37450,N_35005);
or U43774 (N_43774,N_36706,N_39215);
and U43775 (N_43775,N_39171,N_39213);
nand U43776 (N_43776,N_37403,N_39232);
nand U43777 (N_43777,N_39221,N_38450);
nand U43778 (N_43778,N_37284,N_37781);
or U43779 (N_43779,N_35224,N_37504);
or U43780 (N_43780,N_38521,N_38336);
nand U43781 (N_43781,N_35554,N_36243);
and U43782 (N_43782,N_35089,N_37493);
xor U43783 (N_43783,N_38505,N_35512);
or U43784 (N_43784,N_35313,N_37501);
xor U43785 (N_43785,N_37386,N_35804);
nand U43786 (N_43786,N_39808,N_37854);
nand U43787 (N_43787,N_35259,N_35517);
nor U43788 (N_43788,N_36233,N_36600);
nor U43789 (N_43789,N_39640,N_38867);
and U43790 (N_43790,N_36332,N_38987);
nor U43791 (N_43791,N_37714,N_35994);
and U43792 (N_43792,N_35578,N_35761);
nand U43793 (N_43793,N_35770,N_37667);
nor U43794 (N_43794,N_39865,N_35808);
or U43795 (N_43795,N_35460,N_38676);
and U43796 (N_43796,N_37589,N_37919);
xnor U43797 (N_43797,N_39005,N_37037);
or U43798 (N_43798,N_36056,N_38759);
xnor U43799 (N_43799,N_35636,N_36836);
xnor U43800 (N_43800,N_39269,N_39067);
or U43801 (N_43801,N_35028,N_36594);
nand U43802 (N_43802,N_38264,N_35071);
and U43803 (N_43803,N_36475,N_36407);
nand U43804 (N_43804,N_38861,N_39074);
xor U43805 (N_43805,N_36149,N_38549);
xnor U43806 (N_43806,N_37248,N_39567);
nand U43807 (N_43807,N_39137,N_38531);
or U43808 (N_43808,N_39416,N_35462);
nand U43809 (N_43809,N_37350,N_37615);
nor U43810 (N_43810,N_39330,N_38261);
nand U43811 (N_43811,N_39792,N_35126);
nand U43812 (N_43812,N_39947,N_37633);
or U43813 (N_43813,N_36265,N_39354);
nor U43814 (N_43814,N_36970,N_36041);
xnor U43815 (N_43815,N_37521,N_39620);
xor U43816 (N_43816,N_36299,N_35076);
xor U43817 (N_43817,N_36239,N_37821);
xor U43818 (N_43818,N_39441,N_38431);
nor U43819 (N_43819,N_37468,N_39550);
and U43820 (N_43820,N_36156,N_35797);
and U43821 (N_43821,N_35268,N_39333);
xnor U43822 (N_43822,N_35770,N_37284);
nand U43823 (N_43823,N_36300,N_38136);
xnor U43824 (N_43824,N_35146,N_35424);
xnor U43825 (N_43825,N_37280,N_37105);
xor U43826 (N_43826,N_36953,N_36729);
nor U43827 (N_43827,N_38848,N_37123);
and U43828 (N_43828,N_37657,N_37724);
nand U43829 (N_43829,N_38343,N_35740);
and U43830 (N_43830,N_37855,N_36705);
or U43831 (N_43831,N_37294,N_38135);
nor U43832 (N_43832,N_39892,N_38841);
nor U43833 (N_43833,N_36645,N_38286);
nor U43834 (N_43834,N_37827,N_36388);
xor U43835 (N_43835,N_35664,N_38884);
or U43836 (N_43836,N_36998,N_38014);
and U43837 (N_43837,N_39639,N_37593);
and U43838 (N_43838,N_36275,N_38015);
nand U43839 (N_43839,N_39572,N_39941);
xnor U43840 (N_43840,N_39235,N_36611);
xnor U43841 (N_43841,N_37970,N_36786);
and U43842 (N_43842,N_38438,N_36266);
nor U43843 (N_43843,N_39116,N_39599);
nor U43844 (N_43844,N_35862,N_39403);
xnor U43845 (N_43845,N_36016,N_35859);
xor U43846 (N_43846,N_35416,N_36677);
xor U43847 (N_43847,N_35406,N_39616);
nand U43848 (N_43848,N_38671,N_36359);
nor U43849 (N_43849,N_39072,N_37145);
nor U43850 (N_43850,N_36101,N_35323);
and U43851 (N_43851,N_36326,N_38145);
nand U43852 (N_43852,N_35363,N_37247);
and U43853 (N_43853,N_37482,N_36366);
nor U43854 (N_43854,N_39957,N_35741);
nand U43855 (N_43855,N_37981,N_38760);
nand U43856 (N_43856,N_35019,N_36586);
nor U43857 (N_43857,N_35093,N_39485);
or U43858 (N_43858,N_35674,N_39533);
xor U43859 (N_43859,N_39735,N_37326);
nor U43860 (N_43860,N_37867,N_37570);
nor U43861 (N_43861,N_38635,N_35417);
nor U43862 (N_43862,N_39032,N_38637);
nand U43863 (N_43863,N_37869,N_38894);
and U43864 (N_43864,N_38833,N_37149);
nor U43865 (N_43865,N_35843,N_35327);
xor U43866 (N_43866,N_36545,N_36981);
or U43867 (N_43867,N_36181,N_36745);
nor U43868 (N_43868,N_36715,N_37644);
nand U43869 (N_43869,N_36527,N_37736);
and U43870 (N_43870,N_37878,N_38040);
nor U43871 (N_43871,N_36994,N_35695);
nand U43872 (N_43872,N_39655,N_38921);
xor U43873 (N_43873,N_36826,N_37571);
xnor U43874 (N_43874,N_38303,N_36357);
nand U43875 (N_43875,N_39306,N_36594);
or U43876 (N_43876,N_37065,N_35633);
and U43877 (N_43877,N_36866,N_39868);
and U43878 (N_43878,N_38422,N_39580);
nor U43879 (N_43879,N_38145,N_39362);
or U43880 (N_43880,N_36763,N_36884);
and U43881 (N_43881,N_39396,N_38923);
nand U43882 (N_43882,N_38725,N_36025);
and U43883 (N_43883,N_39983,N_39692);
and U43884 (N_43884,N_36292,N_38869);
xor U43885 (N_43885,N_37379,N_39782);
xnor U43886 (N_43886,N_35738,N_37003);
or U43887 (N_43887,N_38966,N_37740);
or U43888 (N_43888,N_39018,N_36778);
nor U43889 (N_43889,N_37614,N_36923);
and U43890 (N_43890,N_39816,N_39500);
and U43891 (N_43891,N_39202,N_39014);
nand U43892 (N_43892,N_37069,N_36055);
xnor U43893 (N_43893,N_39272,N_37879);
nand U43894 (N_43894,N_36106,N_37269);
and U43895 (N_43895,N_37327,N_37038);
xnor U43896 (N_43896,N_37685,N_35135);
nor U43897 (N_43897,N_37644,N_37570);
nand U43898 (N_43898,N_38858,N_38448);
xor U43899 (N_43899,N_36930,N_39305);
and U43900 (N_43900,N_37964,N_38016);
xor U43901 (N_43901,N_35774,N_39809);
nor U43902 (N_43902,N_36292,N_37225);
nor U43903 (N_43903,N_37158,N_35214);
and U43904 (N_43904,N_35152,N_38123);
nand U43905 (N_43905,N_37889,N_37094);
xor U43906 (N_43906,N_36739,N_38600);
nand U43907 (N_43907,N_36717,N_37233);
nand U43908 (N_43908,N_36439,N_37688);
nand U43909 (N_43909,N_35909,N_37606);
nand U43910 (N_43910,N_35562,N_39004);
xor U43911 (N_43911,N_37872,N_35690);
xor U43912 (N_43912,N_35340,N_36765);
nand U43913 (N_43913,N_37744,N_38312);
and U43914 (N_43914,N_35332,N_39924);
nor U43915 (N_43915,N_38694,N_36720);
xor U43916 (N_43916,N_36120,N_36766);
and U43917 (N_43917,N_35630,N_39180);
nor U43918 (N_43918,N_39539,N_35494);
or U43919 (N_43919,N_36738,N_37981);
xor U43920 (N_43920,N_39911,N_35007);
nor U43921 (N_43921,N_37738,N_35154);
xor U43922 (N_43922,N_35806,N_39993);
nand U43923 (N_43923,N_38067,N_35967);
or U43924 (N_43924,N_36423,N_37981);
or U43925 (N_43925,N_35270,N_39974);
and U43926 (N_43926,N_37061,N_39500);
nand U43927 (N_43927,N_37009,N_36618);
or U43928 (N_43928,N_36579,N_35739);
nand U43929 (N_43929,N_39973,N_38132);
nor U43930 (N_43930,N_35383,N_38656);
or U43931 (N_43931,N_36511,N_37193);
nor U43932 (N_43932,N_37295,N_38541);
xor U43933 (N_43933,N_37221,N_36780);
and U43934 (N_43934,N_37371,N_37825);
or U43935 (N_43935,N_39637,N_36394);
or U43936 (N_43936,N_39116,N_36256);
and U43937 (N_43937,N_38952,N_37951);
nor U43938 (N_43938,N_36917,N_35800);
nand U43939 (N_43939,N_37782,N_36923);
nand U43940 (N_43940,N_36279,N_35151);
or U43941 (N_43941,N_38922,N_35329);
xor U43942 (N_43942,N_37381,N_36796);
or U43943 (N_43943,N_38565,N_36985);
nor U43944 (N_43944,N_36740,N_39377);
xnor U43945 (N_43945,N_38334,N_38951);
nand U43946 (N_43946,N_35007,N_36265);
nor U43947 (N_43947,N_35655,N_39655);
xnor U43948 (N_43948,N_39373,N_35757);
xnor U43949 (N_43949,N_37906,N_35737);
or U43950 (N_43950,N_39656,N_36449);
or U43951 (N_43951,N_35006,N_37072);
or U43952 (N_43952,N_38060,N_38421);
or U43953 (N_43953,N_39366,N_35986);
and U43954 (N_43954,N_38305,N_37658);
nand U43955 (N_43955,N_39274,N_36255);
nand U43956 (N_43956,N_38464,N_38467);
or U43957 (N_43957,N_35630,N_38867);
nand U43958 (N_43958,N_36843,N_39088);
xnor U43959 (N_43959,N_36159,N_39857);
nor U43960 (N_43960,N_36810,N_36098);
or U43961 (N_43961,N_38560,N_39745);
and U43962 (N_43962,N_36275,N_36962);
xor U43963 (N_43963,N_39978,N_35231);
and U43964 (N_43964,N_35130,N_37294);
xnor U43965 (N_43965,N_38830,N_36928);
nor U43966 (N_43966,N_37298,N_35029);
nor U43967 (N_43967,N_38922,N_38474);
nor U43968 (N_43968,N_36245,N_39603);
or U43969 (N_43969,N_38150,N_37488);
xor U43970 (N_43970,N_36972,N_35001);
xor U43971 (N_43971,N_38120,N_38754);
and U43972 (N_43972,N_35253,N_36043);
xnor U43973 (N_43973,N_35876,N_37634);
nor U43974 (N_43974,N_36804,N_37454);
or U43975 (N_43975,N_37674,N_36129);
xnor U43976 (N_43976,N_39310,N_35944);
nand U43977 (N_43977,N_35391,N_35777);
nor U43978 (N_43978,N_38551,N_39898);
nor U43979 (N_43979,N_38154,N_38755);
nand U43980 (N_43980,N_39723,N_37401);
or U43981 (N_43981,N_37658,N_38812);
xor U43982 (N_43982,N_39356,N_37899);
nand U43983 (N_43983,N_38765,N_38480);
and U43984 (N_43984,N_37545,N_37063);
nor U43985 (N_43985,N_38094,N_38558);
nand U43986 (N_43986,N_37566,N_39346);
or U43987 (N_43987,N_36820,N_37593);
nand U43988 (N_43988,N_38713,N_35574);
nor U43989 (N_43989,N_39250,N_36454);
or U43990 (N_43990,N_36254,N_35838);
nand U43991 (N_43991,N_38702,N_37405);
or U43992 (N_43992,N_38311,N_35480);
nand U43993 (N_43993,N_36495,N_35260);
and U43994 (N_43994,N_36574,N_37837);
nand U43995 (N_43995,N_36310,N_39912);
nand U43996 (N_43996,N_39325,N_38106);
xor U43997 (N_43997,N_35226,N_35837);
nand U43998 (N_43998,N_39750,N_38828);
or U43999 (N_43999,N_38945,N_39914);
and U44000 (N_44000,N_36322,N_37494);
nor U44001 (N_44001,N_37522,N_38706);
nor U44002 (N_44002,N_39417,N_36444);
nor U44003 (N_44003,N_38440,N_36743);
nand U44004 (N_44004,N_37437,N_37703);
xor U44005 (N_44005,N_39267,N_36149);
nor U44006 (N_44006,N_35471,N_35461);
nor U44007 (N_44007,N_36708,N_36228);
nand U44008 (N_44008,N_36333,N_39770);
nand U44009 (N_44009,N_39162,N_37610);
xor U44010 (N_44010,N_35460,N_39956);
or U44011 (N_44011,N_38017,N_35626);
and U44012 (N_44012,N_36929,N_39483);
xor U44013 (N_44013,N_36315,N_39318);
nand U44014 (N_44014,N_37567,N_37547);
xor U44015 (N_44015,N_35686,N_36007);
nand U44016 (N_44016,N_36464,N_38670);
nand U44017 (N_44017,N_36151,N_36544);
or U44018 (N_44018,N_38906,N_36168);
or U44019 (N_44019,N_39688,N_36673);
xnor U44020 (N_44020,N_35006,N_35526);
nor U44021 (N_44021,N_37934,N_38421);
nand U44022 (N_44022,N_38877,N_37040);
xnor U44023 (N_44023,N_38967,N_39325);
xnor U44024 (N_44024,N_35118,N_35756);
and U44025 (N_44025,N_38034,N_37284);
or U44026 (N_44026,N_39002,N_36897);
nand U44027 (N_44027,N_37313,N_39285);
or U44028 (N_44028,N_38651,N_39874);
nand U44029 (N_44029,N_36446,N_39205);
nor U44030 (N_44030,N_39376,N_39941);
or U44031 (N_44031,N_39811,N_38007);
nor U44032 (N_44032,N_38183,N_35209);
xnor U44033 (N_44033,N_37232,N_38743);
xnor U44034 (N_44034,N_39195,N_37839);
nor U44035 (N_44035,N_38500,N_38664);
and U44036 (N_44036,N_35221,N_36779);
nor U44037 (N_44037,N_37744,N_39685);
nor U44038 (N_44038,N_36189,N_39130);
xnor U44039 (N_44039,N_38411,N_36482);
and U44040 (N_44040,N_39603,N_39003);
or U44041 (N_44041,N_38332,N_38732);
nand U44042 (N_44042,N_36447,N_39475);
or U44043 (N_44043,N_36692,N_36122);
or U44044 (N_44044,N_36239,N_39417);
nand U44045 (N_44045,N_36987,N_37366);
and U44046 (N_44046,N_36893,N_37034);
nor U44047 (N_44047,N_38136,N_36679);
nor U44048 (N_44048,N_36527,N_35604);
or U44049 (N_44049,N_35702,N_39586);
and U44050 (N_44050,N_37900,N_38234);
nor U44051 (N_44051,N_35252,N_36700);
xnor U44052 (N_44052,N_35289,N_37070);
nand U44053 (N_44053,N_37923,N_39443);
or U44054 (N_44054,N_37307,N_38165);
xor U44055 (N_44055,N_36826,N_39894);
xor U44056 (N_44056,N_36128,N_37997);
nand U44057 (N_44057,N_39687,N_38955);
nand U44058 (N_44058,N_35581,N_39228);
nand U44059 (N_44059,N_35000,N_38543);
nor U44060 (N_44060,N_36928,N_35262);
nand U44061 (N_44061,N_35929,N_37604);
or U44062 (N_44062,N_38757,N_37866);
or U44063 (N_44063,N_38124,N_35856);
xnor U44064 (N_44064,N_38942,N_38509);
or U44065 (N_44065,N_39225,N_39562);
nand U44066 (N_44066,N_35349,N_36882);
nor U44067 (N_44067,N_37069,N_37468);
xor U44068 (N_44068,N_38107,N_35781);
xnor U44069 (N_44069,N_39490,N_35866);
xnor U44070 (N_44070,N_38896,N_38247);
nand U44071 (N_44071,N_38801,N_35657);
nand U44072 (N_44072,N_37432,N_35393);
and U44073 (N_44073,N_36334,N_37347);
xnor U44074 (N_44074,N_39708,N_38693);
or U44075 (N_44075,N_38264,N_38337);
nor U44076 (N_44076,N_36296,N_39911);
and U44077 (N_44077,N_38566,N_39457);
or U44078 (N_44078,N_37750,N_38221);
or U44079 (N_44079,N_35192,N_35048);
nand U44080 (N_44080,N_39904,N_39814);
and U44081 (N_44081,N_36647,N_36575);
or U44082 (N_44082,N_37676,N_36255);
and U44083 (N_44083,N_39241,N_39725);
nand U44084 (N_44084,N_35468,N_38210);
xor U44085 (N_44085,N_36872,N_37820);
and U44086 (N_44086,N_36187,N_38723);
nand U44087 (N_44087,N_38519,N_38741);
xor U44088 (N_44088,N_35068,N_36270);
or U44089 (N_44089,N_38196,N_39058);
and U44090 (N_44090,N_37807,N_39957);
nand U44091 (N_44091,N_35820,N_39016);
and U44092 (N_44092,N_38437,N_37440);
nand U44093 (N_44093,N_38534,N_39768);
and U44094 (N_44094,N_35238,N_39211);
or U44095 (N_44095,N_37739,N_39225);
nor U44096 (N_44096,N_36922,N_38357);
nor U44097 (N_44097,N_35453,N_37299);
and U44098 (N_44098,N_35131,N_36603);
and U44099 (N_44099,N_37366,N_37841);
xor U44100 (N_44100,N_39223,N_39734);
xnor U44101 (N_44101,N_35682,N_35508);
xnor U44102 (N_44102,N_38355,N_39431);
nand U44103 (N_44103,N_37671,N_35839);
nand U44104 (N_44104,N_36786,N_36215);
nand U44105 (N_44105,N_39072,N_36447);
xor U44106 (N_44106,N_38042,N_36109);
nor U44107 (N_44107,N_39374,N_38988);
xor U44108 (N_44108,N_37422,N_36006);
nor U44109 (N_44109,N_39231,N_39265);
nand U44110 (N_44110,N_38063,N_38410);
nand U44111 (N_44111,N_39693,N_38367);
or U44112 (N_44112,N_35807,N_37767);
xnor U44113 (N_44113,N_37938,N_37359);
nand U44114 (N_44114,N_39414,N_37888);
nor U44115 (N_44115,N_38035,N_37163);
nand U44116 (N_44116,N_35533,N_39078);
nand U44117 (N_44117,N_36109,N_39129);
xor U44118 (N_44118,N_38755,N_35036);
xnor U44119 (N_44119,N_38202,N_37612);
nor U44120 (N_44120,N_37098,N_37052);
or U44121 (N_44121,N_38623,N_38657);
or U44122 (N_44122,N_35183,N_36468);
or U44123 (N_44123,N_39068,N_36267);
nor U44124 (N_44124,N_38328,N_38036);
nor U44125 (N_44125,N_35676,N_39645);
xor U44126 (N_44126,N_36961,N_37438);
or U44127 (N_44127,N_39154,N_36212);
or U44128 (N_44128,N_37731,N_39675);
or U44129 (N_44129,N_37914,N_38064);
nand U44130 (N_44130,N_39483,N_36376);
xnor U44131 (N_44131,N_35049,N_36496);
nor U44132 (N_44132,N_38157,N_39006);
and U44133 (N_44133,N_38758,N_38133);
xor U44134 (N_44134,N_38232,N_35415);
xnor U44135 (N_44135,N_39345,N_39601);
or U44136 (N_44136,N_38515,N_38255);
xor U44137 (N_44137,N_38723,N_37629);
and U44138 (N_44138,N_35726,N_38156);
and U44139 (N_44139,N_35325,N_35382);
nand U44140 (N_44140,N_37394,N_39285);
or U44141 (N_44141,N_38327,N_36213);
nand U44142 (N_44142,N_36785,N_37409);
xor U44143 (N_44143,N_38383,N_36744);
nand U44144 (N_44144,N_37969,N_38362);
xnor U44145 (N_44145,N_36717,N_36171);
or U44146 (N_44146,N_38780,N_38199);
nor U44147 (N_44147,N_39704,N_39867);
and U44148 (N_44148,N_37455,N_36837);
nand U44149 (N_44149,N_36297,N_38213);
nand U44150 (N_44150,N_35162,N_36838);
nand U44151 (N_44151,N_39921,N_39196);
and U44152 (N_44152,N_35899,N_39156);
nor U44153 (N_44153,N_38967,N_39599);
or U44154 (N_44154,N_37936,N_35914);
xor U44155 (N_44155,N_38134,N_37206);
nand U44156 (N_44156,N_39471,N_37371);
or U44157 (N_44157,N_35166,N_35924);
nor U44158 (N_44158,N_38169,N_36059);
nand U44159 (N_44159,N_37209,N_38692);
and U44160 (N_44160,N_36346,N_38721);
or U44161 (N_44161,N_36116,N_38010);
nand U44162 (N_44162,N_37027,N_35284);
or U44163 (N_44163,N_39423,N_38027);
nand U44164 (N_44164,N_35347,N_37030);
and U44165 (N_44165,N_37834,N_35692);
and U44166 (N_44166,N_35599,N_35110);
and U44167 (N_44167,N_35161,N_36010);
and U44168 (N_44168,N_37519,N_35127);
nand U44169 (N_44169,N_38824,N_36972);
or U44170 (N_44170,N_37498,N_38126);
and U44171 (N_44171,N_38749,N_39501);
or U44172 (N_44172,N_37285,N_37899);
or U44173 (N_44173,N_37546,N_38134);
xnor U44174 (N_44174,N_36210,N_37007);
nor U44175 (N_44175,N_39622,N_37723);
nor U44176 (N_44176,N_36976,N_39447);
and U44177 (N_44177,N_39269,N_36793);
or U44178 (N_44178,N_35717,N_39496);
nor U44179 (N_44179,N_38521,N_39300);
nor U44180 (N_44180,N_35725,N_38085);
nor U44181 (N_44181,N_36556,N_36070);
or U44182 (N_44182,N_38291,N_35808);
xnor U44183 (N_44183,N_35986,N_38478);
nor U44184 (N_44184,N_38486,N_35608);
or U44185 (N_44185,N_37448,N_38250);
nand U44186 (N_44186,N_37374,N_37443);
xor U44187 (N_44187,N_38449,N_35356);
and U44188 (N_44188,N_37276,N_37660);
nand U44189 (N_44189,N_36542,N_37031);
nor U44190 (N_44190,N_38256,N_36695);
and U44191 (N_44191,N_36094,N_36230);
and U44192 (N_44192,N_38333,N_36678);
xor U44193 (N_44193,N_38166,N_37183);
nand U44194 (N_44194,N_35604,N_38509);
or U44195 (N_44195,N_38684,N_37833);
nand U44196 (N_44196,N_38043,N_36260);
and U44197 (N_44197,N_39478,N_36370);
xnor U44198 (N_44198,N_39211,N_37370);
and U44199 (N_44199,N_37044,N_39347);
xor U44200 (N_44200,N_37090,N_35822);
nor U44201 (N_44201,N_37811,N_36137);
nand U44202 (N_44202,N_35838,N_36193);
xnor U44203 (N_44203,N_39841,N_37222);
and U44204 (N_44204,N_35263,N_38006);
xor U44205 (N_44205,N_39282,N_39353);
nand U44206 (N_44206,N_35070,N_37900);
nand U44207 (N_44207,N_36107,N_36627);
xnor U44208 (N_44208,N_37193,N_36981);
and U44209 (N_44209,N_39079,N_39254);
or U44210 (N_44210,N_37784,N_39005);
and U44211 (N_44211,N_36721,N_39462);
or U44212 (N_44212,N_36184,N_39359);
nand U44213 (N_44213,N_39333,N_35167);
nand U44214 (N_44214,N_37718,N_35935);
or U44215 (N_44215,N_38099,N_36435);
and U44216 (N_44216,N_36464,N_37988);
xnor U44217 (N_44217,N_37757,N_37324);
xnor U44218 (N_44218,N_37752,N_35723);
and U44219 (N_44219,N_35408,N_38995);
nor U44220 (N_44220,N_37759,N_38977);
nor U44221 (N_44221,N_37492,N_38650);
xnor U44222 (N_44222,N_39773,N_35947);
nand U44223 (N_44223,N_39044,N_39145);
and U44224 (N_44224,N_35914,N_36418);
nand U44225 (N_44225,N_39228,N_37818);
or U44226 (N_44226,N_37926,N_39017);
or U44227 (N_44227,N_35601,N_35658);
or U44228 (N_44228,N_39316,N_38819);
and U44229 (N_44229,N_39022,N_36927);
or U44230 (N_44230,N_35355,N_35134);
nand U44231 (N_44231,N_35056,N_39900);
and U44232 (N_44232,N_38551,N_37395);
nor U44233 (N_44233,N_35669,N_36843);
nor U44234 (N_44234,N_37044,N_37488);
or U44235 (N_44235,N_39964,N_36390);
xnor U44236 (N_44236,N_36940,N_37159);
nand U44237 (N_44237,N_39317,N_37959);
nor U44238 (N_44238,N_36694,N_35605);
nand U44239 (N_44239,N_39579,N_38978);
nand U44240 (N_44240,N_38763,N_36441);
xnor U44241 (N_44241,N_39124,N_37028);
or U44242 (N_44242,N_38173,N_39435);
and U44243 (N_44243,N_37125,N_38086);
nor U44244 (N_44244,N_38344,N_35196);
nand U44245 (N_44245,N_36243,N_36026);
xnor U44246 (N_44246,N_37211,N_35106);
or U44247 (N_44247,N_38162,N_37798);
nor U44248 (N_44248,N_36561,N_38819);
or U44249 (N_44249,N_35565,N_36531);
xor U44250 (N_44250,N_39978,N_39665);
nor U44251 (N_44251,N_38924,N_38537);
or U44252 (N_44252,N_35979,N_38128);
xor U44253 (N_44253,N_39484,N_39181);
nor U44254 (N_44254,N_37921,N_38704);
and U44255 (N_44255,N_37145,N_35376);
nor U44256 (N_44256,N_38882,N_37460);
nand U44257 (N_44257,N_37647,N_35995);
nor U44258 (N_44258,N_35073,N_36542);
xor U44259 (N_44259,N_37896,N_37160);
and U44260 (N_44260,N_39359,N_37664);
xnor U44261 (N_44261,N_37618,N_39147);
nor U44262 (N_44262,N_38572,N_36214);
xnor U44263 (N_44263,N_36005,N_39913);
nand U44264 (N_44264,N_39720,N_39578);
nand U44265 (N_44265,N_35292,N_39436);
xor U44266 (N_44266,N_37777,N_37308);
nor U44267 (N_44267,N_35746,N_37639);
or U44268 (N_44268,N_39794,N_38101);
nor U44269 (N_44269,N_39173,N_37058);
nand U44270 (N_44270,N_38660,N_39266);
xnor U44271 (N_44271,N_35636,N_35959);
or U44272 (N_44272,N_37187,N_38939);
xnor U44273 (N_44273,N_39031,N_36440);
nor U44274 (N_44274,N_38763,N_38149);
xnor U44275 (N_44275,N_35474,N_36670);
nor U44276 (N_44276,N_38653,N_36564);
xor U44277 (N_44277,N_38684,N_37070);
nor U44278 (N_44278,N_38320,N_38675);
nor U44279 (N_44279,N_37746,N_39875);
nor U44280 (N_44280,N_36168,N_39768);
nor U44281 (N_44281,N_38025,N_39298);
or U44282 (N_44282,N_37372,N_37795);
nor U44283 (N_44283,N_35085,N_39012);
nand U44284 (N_44284,N_38986,N_37482);
and U44285 (N_44285,N_39137,N_38923);
xor U44286 (N_44286,N_38543,N_39805);
xor U44287 (N_44287,N_39214,N_36662);
nor U44288 (N_44288,N_39704,N_37051);
or U44289 (N_44289,N_36350,N_39911);
or U44290 (N_44290,N_35373,N_38016);
xor U44291 (N_44291,N_37150,N_35335);
nand U44292 (N_44292,N_35866,N_36122);
xnor U44293 (N_44293,N_35776,N_35953);
and U44294 (N_44294,N_36195,N_39995);
and U44295 (N_44295,N_39373,N_35634);
xor U44296 (N_44296,N_38348,N_37184);
nor U44297 (N_44297,N_37957,N_36394);
and U44298 (N_44298,N_35176,N_38853);
nor U44299 (N_44299,N_39598,N_39238);
or U44300 (N_44300,N_35271,N_37031);
and U44301 (N_44301,N_36024,N_39228);
nor U44302 (N_44302,N_36051,N_35968);
nor U44303 (N_44303,N_38565,N_39738);
nor U44304 (N_44304,N_39894,N_37604);
xnor U44305 (N_44305,N_37030,N_37152);
xnor U44306 (N_44306,N_39149,N_39015);
xnor U44307 (N_44307,N_36633,N_38845);
nor U44308 (N_44308,N_35964,N_38280);
and U44309 (N_44309,N_35454,N_37643);
or U44310 (N_44310,N_38269,N_35043);
nand U44311 (N_44311,N_35631,N_38925);
nor U44312 (N_44312,N_36091,N_39863);
nor U44313 (N_44313,N_35714,N_36992);
xnor U44314 (N_44314,N_39069,N_39366);
or U44315 (N_44315,N_38283,N_38922);
xnor U44316 (N_44316,N_35960,N_38958);
and U44317 (N_44317,N_39732,N_38796);
and U44318 (N_44318,N_38863,N_36716);
nand U44319 (N_44319,N_37017,N_36088);
nand U44320 (N_44320,N_37998,N_38839);
nand U44321 (N_44321,N_37999,N_38787);
xor U44322 (N_44322,N_39252,N_37750);
and U44323 (N_44323,N_35484,N_38909);
nor U44324 (N_44324,N_37376,N_37707);
xnor U44325 (N_44325,N_38580,N_39673);
and U44326 (N_44326,N_38152,N_35690);
nor U44327 (N_44327,N_39475,N_37764);
nor U44328 (N_44328,N_36374,N_38027);
xnor U44329 (N_44329,N_38267,N_37837);
nor U44330 (N_44330,N_38068,N_36675);
or U44331 (N_44331,N_36472,N_38716);
xnor U44332 (N_44332,N_38349,N_37636);
nor U44333 (N_44333,N_37690,N_36484);
nor U44334 (N_44334,N_36783,N_35151);
nand U44335 (N_44335,N_35331,N_36311);
or U44336 (N_44336,N_38208,N_38629);
xnor U44337 (N_44337,N_39740,N_36518);
nor U44338 (N_44338,N_38764,N_39231);
xnor U44339 (N_44339,N_36981,N_37807);
nand U44340 (N_44340,N_36766,N_36942);
nand U44341 (N_44341,N_36303,N_36811);
nand U44342 (N_44342,N_39305,N_37881);
nor U44343 (N_44343,N_39390,N_35502);
or U44344 (N_44344,N_36796,N_39629);
nor U44345 (N_44345,N_35730,N_36896);
and U44346 (N_44346,N_35935,N_39558);
nor U44347 (N_44347,N_38383,N_36945);
nand U44348 (N_44348,N_37729,N_35716);
nor U44349 (N_44349,N_39837,N_36207);
xnor U44350 (N_44350,N_38161,N_38293);
and U44351 (N_44351,N_36531,N_37891);
nor U44352 (N_44352,N_38604,N_37565);
xnor U44353 (N_44353,N_35570,N_38702);
or U44354 (N_44354,N_35520,N_35769);
nor U44355 (N_44355,N_35000,N_35458);
and U44356 (N_44356,N_35690,N_36780);
nor U44357 (N_44357,N_39836,N_36569);
or U44358 (N_44358,N_36636,N_37471);
and U44359 (N_44359,N_37458,N_37906);
and U44360 (N_44360,N_36785,N_37599);
and U44361 (N_44361,N_38902,N_36070);
or U44362 (N_44362,N_37673,N_36267);
xor U44363 (N_44363,N_37793,N_38552);
and U44364 (N_44364,N_37789,N_39563);
nor U44365 (N_44365,N_37658,N_39885);
nand U44366 (N_44366,N_35843,N_35680);
nand U44367 (N_44367,N_36869,N_36481);
or U44368 (N_44368,N_37783,N_39343);
xnor U44369 (N_44369,N_36978,N_39049);
xnor U44370 (N_44370,N_37328,N_36688);
nand U44371 (N_44371,N_35745,N_35459);
nand U44372 (N_44372,N_39756,N_38285);
or U44373 (N_44373,N_38457,N_37959);
nor U44374 (N_44374,N_36681,N_37811);
and U44375 (N_44375,N_37184,N_38814);
xnor U44376 (N_44376,N_39473,N_38798);
xnor U44377 (N_44377,N_36356,N_35541);
nand U44378 (N_44378,N_37136,N_37178);
nand U44379 (N_44379,N_38498,N_36822);
xor U44380 (N_44380,N_36880,N_38191);
and U44381 (N_44381,N_37798,N_37293);
nand U44382 (N_44382,N_39573,N_38108);
nor U44383 (N_44383,N_37885,N_38767);
xnor U44384 (N_44384,N_37033,N_35192);
xnor U44385 (N_44385,N_36896,N_37351);
nand U44386 (N_44386,N_38927,N_39599);
and U44387 (N_44387,N_36515,N_38760);
or U44388 (N_44388,N_37043,N_37142);
nand U44389 (N_44389,N_39508,N_35590);
xnor U44390 (N_44390,N_38065,N_35921);
nor U44391 (N_44391,N_37215,N_37801);
nor U44392 (N_44392,N_39321,N_39015);
nand U44393 (N_44393,N_35840,N_36994);
nand U44394 (N_44394,N_38526,N_36344);
xor U44395 (N_44395,N_36221,N_36028);
nor U44396 (N_44396,N_38708,N_36892);
nor U44397 (N_44397,N_38798,N_37328);
xor U44398 (N_44398,N_37789,N_39354);
nor U44399 (N_44399,N_39195,N_38971);
or U44400 (N_44400,N_35531,N_39887);
nor U44401 (N_44401,N_37431,N_38537);
or U44402 (N_44402,N_39834,N_38003);
nand U44403 (N_44403,N_39488,N_35836);
xnor U44404 (N_44404,N_36222,N_35813);
or U44405 (N_44405,N_36950,N_35802);
xor U44406 (N_44406,N_38053,N_35394);
nor U44407 (N_44407,N_38455,N_38205);
nand U44408 (N_44408,N_39671,N_35099);
and U44409 (N_44409,N_37568,N_37535);
and U44410 (N_44410,N_38775,N_39034);
and U44411 (N_44411,N_37238,N_38345);
and U44412 (N_44412,N_36258,N_35210);
or U44413 (N_44413,N_37034,N_39407);
nand U44414 (N_44414,N_39537,N_35481);
xor U44415 (N_44415,N_37603,N_39654);
xnor U44416 (N_44416,N_39158,N_36382);
xnor U44417 (N_44417,N_35882,N_37027);
or U44418 (N_44418,N_35624,N_38275);
and U44419 (N_44419,N_37598,N_36813);
and U44420 (N_44420,N_39781,N_37002);
nand U44421 (N_44421,N_37192,N_38082);
and U44422 (N_44422,N_36948,N_36773);
nor U44423 (N_44423,N_36054,N_37904);
nand U44424 (N_44424,N_38817,N_37004);
or U44425 (N_44425,N_37516,N_35600);
nor U44426 (N_44426,N_35609,N_37703);
nor U44427 (N_44427,N_39258,N_35303);
nor U44428 (N_44428,N_35131,N_35611);
xor U44429 (N_44429,N_35647,N_37770);
and U44430 (N_44430,N_39875,N_36274);
and U44431 (N_44431,N_35545,N_36195);
xor U44432 (N_44432,N_37397,N_37655);
nand U44433 (N_44433,N_38438,N_36099);
nor U44434 (N_44434,N_36800,N_39322);
nor U44435 (N_44435,N_39015,N_39144);
xor U44436 (N_44436,N_38216,N_38006);
nand U44437 (N_44437,N_38891,N_35797);
and U44438 (N_44438,N_39657,N_35357);
or U44439 (N_44439,N_39410,N_35262);
and U44440 (N_44440,N_38737,N_37884);
xnor U44441 (N_44441,N_39292,N_35427);
nand U44442 (N_44442,N_36218,N_37477);
nand U44443 (N_44443,N_37672,N_36881);
and U44444 (N_44444,N_39879,N_36020);
and U44445 (N_44445,N_37651,N_38629);
nand U44446 (N_44446,N_39566,N_35369);
nor U44447 (N_44447,N_39739,N_36536);
and U44448 (N_44448,N_37087,N_37556);
or U44449 (N_44449,N_38962,N_37680);
or U44450 (N_44450,N_37969,N_38477);
nor U44451 (N_44451,N_37000,N_38432);
nand U44452 (N_44452,N_35620,N_38759);
nor U44453 (N_44453,N_39455,N_35316);
and U44454 (N_44454,N_38814,N_39652);
xnor U44455 (N_44455,N_39673,N_39715);
or U44456 (N_44456,N_36290,N_37701);
or U44457 (N_44457,N_38090,N_36982);
nor U44458 (N_44458,N_38604,N_35348);
nor U44459 (N_44459,N_35797,N_37685);
xnor U44460 (N_44460,N_35382,N_37004);
xnor U44461 (N_44461,N_35717,N_39912);
and U44462 (N_44462,N_39222,N_35687);
nand U44463 (N_44463,N_35965,N_36801);
and U44464 (N_44464,N_36234,N_35037);
xnor U44465 (N_44465,N_35167,N_37112);
xnor U44466 (N_44466,N_35120,N_36838);
or U44467 (N_44467,N_38535,N_39375);
xor U44468 (N_44468,N_37208,N_39870);
nor U44469 (N_44469,N_36559,N_38415);
and U44470 (N_44470,N_39296,N_35033);
and U44471 (N_44471,N_38271,N_36852);
nor U44472 (N_44472,N_39465,N_35147);
or U44473 (N_44473,N_35412,N_35229);
nor U44474 (N_44474,N_35266,N_36167);
nand U44475 (N_44475,N_39710,N_36268);
nor U44476 (N_44476,N_37181,N_38909);
nand U44477 (N_44477,N_37601,N_38779);
or U44478 (N_44478,N_39698,N_37197);
nand U44479 (N_44479,N_38920,N_36792);
or U44480 (N_44480,N_36406,N_35825);
nor U44481 (N_44481,N_36768,N_37470);
nor U44482 (N_44482,N_35539,N_35495);
xor U44483 (N_44483,N_38042,N_35563);
or U44484 (N_44484,N_37822,N_36510);
nand U44485 (N_44485,N_36485,N_37435);
or U44486 (N_44486,N_35923,N_39177);
xnor U44487 (N_44487,N_37849,N_39044);
and U44488 (N_44488,N_38077,N_36577);
and U44489 (N_44489,N_36357,N_38556);
nor U44490 (N_44490,N_39267,N_37158);
and U44491 (N_44491,N_38072,N_39543);
nor U44492 (N_44492,N_37214,N_39523);
or U44493 (N_44493,N_36931,N_38953);
xnor U44494 (N_44494,N_37390,N_35248);
or U44495 (N_44495,N_37095,N_37443);
xnor U44496 (N_44496,N_37697,N_37912);
nor U44497 (N_44497,N_36543,N_37761);
or U44498 (N_44498,N_36208,N_36470);
or U44499 (N_44499,N_37927,N_36174);
xor U44500 (N_44500,N_38467,N_36887);
xnor U44501 (N_44501,N_36831,N_35669);
nand U44502 (N_44502,N_36401,N_36515);
or U44503 (N_44503,N_35992,N_35017);
nor U44504 (N_44504,N_35104,N_36955);
or U44505 (N_44505,N_36240,N_35650);
xnor U44506 (N_44506,N_38371,N_39059);
nor U44507 (N_44507,N_38435,N_35031);
xor U44508 (N_44508,N_38808,N_37874);
nor U44509 (N_44509,N_39889,N_39227);
nor U44510 (N_44510,N_38694,N_36725);
or U44511 (N_44511,N_36787,N_35867);
or U44512 (N_44512,N_36850,N_37895);
nand U44513 (N_44513,N_38938,N_39418);
or U44514 (N_44514,N_35866,N_35343);
nor U44515 (N_44515,N_36156,N_38016);
and U44516 (N_44516,N_37668,N_37322);
or U44517 (N_44517,N_38962,N_36607);
nor U44518 (N_44518,N_37417,N_38581);
nand U44519 (N_44519,N_38307,N_37889);
nor U44520 (N_44520,N_38775,N_36252);
and U44521 (N_44521,N_35407,N_37336);
nor U44522 (N_44522,N_37828,N_37559);
xnor U44523 (N_44523,N_35151,N_38393);
or U44524 (N_44524,N_37282,N_35568);
xor U44525 (N_44525,N_35821,N_36441);
xnor U44526 (N_44526,N_37743,N_38425);
or U44527 (N_44527,N_35477,N_37251);
nand U44528 (N_44528,N_38330,N_39007);
nand U44529 (N_44529,N_37467,N_37200);
xor U44530 (N_44530,N_38391,N_35459);
or U44531 (N_44531,N_35280,N_39674);
nand U44532 (N_44532,N_35539,N_35958);
and U44533 (N_44533,N_38266,N_38848);
nand U44534 (N_44534,N_38030,N_39242);
nand U44535 (N_44535,N_35497,N_39808);
nand U44536 (N_44536,N_38967,N_38304);
and U44537 (N_44537,N_39482,N_38883);
and U44538 (N_44538,N_36478,N_37269);
nand U44539 (N_44539,N_35839,N_37334);
xor U44540 (N_44540,N_36409,N_36819);
or U44541 (N_44541,N_37133,N_35463);
nand U44542 (N_44542,N_36816,N_38949);
and U44543 (N_44543,N_36083,N_35573);
xnor U44544 (N_44544,N_38384,N_36368);
xnor U44545 (N_44545,N_38157,N_39663);
nor U44546 (N_44546,N_39354,N_37796);
nor U44547 (N_44547,N_38514,N_38240);
nand U44548 (N_44548,N_36773,N_37701);
nand U44549 (N_44549,N_37230,N_35136);
or U44550 (N_44550,N_39889,N_38241);
nor U44551 (N_44551,N_35152,N_35814);
or U44552 (N_44552,N_38459,N_39693);
xor U44553 (N_44553,N_36711,N_36777);
or U44554 (N_44554,N_38163,N_35492);
or U44555 (N_44555,N_37533,N_37928);
or U44556 (N_44556,N_36379,N_38010);
or U44557 (N_44557,N_35538,N_36753);
xor U44558 (N_44558,N_38966,N_38488);
nor U44559 (N_44559,N_36344,N_39705);
nor U44560 (N_44560,N_36545,N_38659);
and U44561 (N_44561,N_37950,N_37465);
xor U44562 (N_44562,N_35059,N_38904);
nand U44563 (N_44563,N_37182,N_39069);
xnor U44564 (N_44564,N_38918,N_37567);
xor U44565 (N_44565,N_36309,N_35358);
xnor U44566 (N_44566,N_38717,N_37362);
nand U44567 (N_44567,N_36002,N_36105);
and U44568 (N_44568,N_37678,N_38667);
nor U44569 (N_44569,N_35303,N_37475);
nor U44570 (N_44570,N_37642,N_38829);
xor U44571 (N_44571,N_36642,N_39374);
nand U44572 (N_44572,N_38519,N_36580);
nand U44573 (N_44573,N_37915,N_35061);
and U44574 (N_44574,N_36798,N_37894);
nand U44575 (N_44575,N_38356,N_35681);
nor U44576 (N_44576,N_35418,N_37126);
nor U44577 (N_44577,N_36899,N_37512);
nand U44578 (N_44578,N_37211,N_39204);
or U44579 (N_44579,N_39511,N_39683);
nor U44580 (N_44580,N_36947,N_38249);
or U44581 (N_44581,N_36271,N_38083);
and U44582 (N_44582,N_36350,N_37432);
nor U44583 (N_44583,N_38098,N_35629);
nand U44584 (N_44584,N_38156,N_39375);
or U44585 (N_44585,N_35766,N_37962);
or U44586 (N_44586,N_38596,N_37857);
nand U44587 (N_44587,N_36924,N_37668);
nand U44588 (N_44588,N_38246,N_39021);
or U44589 (N_44589,N_36144,N_36711);
or U44590 (N_44590,N_36152,N_35459);
or U44591 (N_44591,N_38212,N_36249);
nand U44592 (N_44592,N_38136,N_36924);
nor U44593 (N_44593,N_38768,N_35842);
nor U44594 (N_44594,N_39598,N_37375);
nor U44595 (N_44595,N_38917,N_35485);
nor U44596 (N_44596,N_38225,N_38655);
or U44597 (N_44597,N_36264,N_35813);
nand U44598 (N_44598,N_35178,N_38630);
and U44599 (N_44599,N_35766,N_39526);
or U44600 (N_44600,N_38703,N_37195);
nor U44601 (N_44601,N_35961,N_37667);
and U44602 (N_44602,N_37396,N_39658);
nor U44603 (N_44603,N_35104,N_36612);
xnor U44604 (N_44604,N_38985,N_35933);
or U44605 (N_44605,N_39515,N_35945);
xnor U44606 (N_44606,N_36493,N_39425);
and U44607 (N_44607,N_38887,N_35727);
or U44608 (N_44608,N_38565,N_38703);
xnor U44609 (N_44609,N_36951,N_39558);
nor U44610 (N_44610,N_38202,N_37072);
and U44611 (N_44611,N_35605,N_37753);
xnor U44612 (N_44612,N_36078,N_35844);
and U44613 (N_44613,N_35796,N_37548);
nand U44614 (N_44614,N_39135,N_35797);
nand U44615 (N_44615,N_39501,N_35574);
or U44616 (N_44616,N_35509,N_38744);
nand U44617 (N_44617,N_37380,N_38425);
or U44618 (N_44618,N_35005,N_36400);
nand U44619 (N_44619,N_38733,N_39305);
or U44620 (N_44620,N_37768,N_36029);
and U44621 (N_44621,N_35369,N_37571);
nor U44622 (N_44622,N_39458,N_35426);
nor U44623 (N_44623,N_38755,N_37212);
nor U44624 (N_44624,N_39260,N_37347);
xor U44625 (N_44625,N_39390,N_38020);
nand U44626 (N_44626,N_37296,N_36236);
xor U44627 (N_44627,N_35724,N_35655);
and U44628 (N_44628,N_39331,N_37041);
or U44629 (N_44629,N_37350,N_36298);
or U44630 (N_44630,N_39810,N_39006);
xnor U44631 (N_44631,N_35016,N_35043);
or U44632 (N_44632,N_38058,N_35248);
and U44633 (N_44633,N_35198,N_37132);
or U44634 (N_44634,N_38038,N_38271);
or U44635 (N_44635,N_37704,N_39754);
xnor U44636 (N_44636,N_39122,N_37745);
nor U44637 (N_44637,N_38489,N_38368);
or U44638 (N_44638,N_38315,N_37850);
or U44639 (N_44639,N_35084,N_38140);
or U44640 (N_44640,N_38873,N_37420);
nor U44641 (N_44641,N_36653,N_39177);
and U44642 (N_44642,N_37017,N_35393);
and U44643 (N_44643,N_35345,N_35597);
nor U44644 (N_44644,N_39930,N_37091);
and U44645 (N_44645,N_36321,N_39051);
nand U44646 (N_44646,N_36591,N_35661);
xor U44647 (N_44647,N_35960,N_36892);
nand U44648 (N_44648,N_35089,N_39201);
xor U44649 (N_44649,N_37668,N_37196);
nand U44650 (N_44650,N_35299,N_38710);
nor U44651 (N_44651,N_37006,N_39272);
xor U44652 (N_44652,N_38053,N_39180);
xnor U44653 (N_44653,N_39931,N_35692);
and U44654 (N_44654,N_36434,N_35336);
xnor U44655 (N_44655,N_36858,N_38945);
nand U44656 (N_44656,N_36637,N_36146);
or U44657 (N_44657,N_36408,N_37660);
or U44658 (N_44658,N_37193,N_37262);
xor U44659 (N_44659,N_37486,N_38591);
or U44660 (N_44660,N_35645,N_36103);
or U44661 (N_44661,N_39600,N_37406);
nand U44662 (N_44662,N_37095,N_35567);
and U44663 (N_44663,N_36658,N_37533);
xnor U44664 (N_44664,N_37402,N_36370);
xnor U44665 (N_44665,N_38779,N_37609);
nand U44666 (N_44666,N_37043,N_39129);
and U44667 (N_44667,N_37415,N_38285);
nor U44668 (N_44668,N_39441,N_36429);
nand U44669 (N_44669,N_36511,N_36640);
and U44670 (N_44670,N_37409,N_36797);
xor U44671 (N_44671,N_35181,N_36694);
nor U44672 (N_44672,N_37998,N_37023);
nand U44673 (N_44673,N_37631,N_38137);
and U44674 (N_44674,N_38165,N_37919);
nor U44675 (N_44675,N_36470,N_35727);
or U44676 (N_44676,N_35677,N_39385);
or U44677 (N_44677,N_37211,N_35217);
xnor U44678 (N_44678,N_35376,N_37274);
nor U44679 (N_44679,N_35970,N_35799);
nand U44680 (N_44680,N_36338,N_39025);
nand U44681 (N_44681,N_36090,N_36857);
xor U44682 (N_44682,N_37870,N_39114);
xor U44683 (N_44683,N_37961,N_39297);
or U44684 (N_44684,N_38710,N_38717);
nor U44685 (N_44685,N_36995,N_35493);
or U44686 (N_44686,N_36062,N_37405);
nand U44687 (N_44687,N_38704,N_35779);
xor U44688 (N_44688,N_38273,N_35802);
or U44689 (N_44689,N_38954,N_39663);
xor U44690 (N_44690,N_36794,N_38056);
xor U44691 (N_44691,N_36554,N_38702);
and U44692 (N_44692,N_39856,N_35954);
nand U44693 (N_44693,N_35795,N_37772);
nand U44694 (N_44694,N_39257,N_38623);
nor U44695 (N_44695,N_38899,N_38592);
xor U44696 (N_44696,N_39873,N_39021);
and U44697 (N_44697,N_36402,N_36903);
nor U44698 (N_44698,N_37117,N_37106);
or U44699 (N_44699,N_38845,N_35772);
nand U44700 (N_44700,N_37269,N_37253);
and U44701 (N_44701,N_36939,N_38313);
or U44702 (N_44702,N_37987,N_38522);
nor U44703 (N_44703,N_38617,N_36437);
and U44704 (N_44704,N_36013,N_36364);
nor U44705 (N_44705,N_35172,N_36567);
nor U44706 (N_44706,N_39191,N_37455);
or U44707 (N_44707,N_38527,N_37981);
nor U44708 (N_44708,N_37043,N_36378);
or U44709 (N_44709,N_38524,N_37980);
xor U44710 (N_44710,N_36145,N_39918);
nand U44711 (N_44711,N_36482,N_37781);
nor U44712 (N_44712,N_37150,N_37060);
and U44713 (N_44713,N_37868,N_38018);
or U44714 (N_44714,N_35776,N_35199);
xor U44715 (N_44715,N_39590,N_36753);
and U44716 (N_44716,N_39537,N_38567);
or U44717 (N_44717,N_38739,N_35123);
and U44718 (N_44718,N_36099,N_37241);
nand U44719 (N_44719,N_39868,N_38015);
xor U44720 (N_44720,N_36610,N_37016);
nand U44721 (N_44721,N_39284,N_39841);
xnor U44722 (N_44722,N_38414,N_39903);
nor U44723 (N_44723,N_35927,N_36921);
xnor U44724 (N_44724,N_35175,N_38646);
nor U44725 (N_44725,N_38008,N_35929);
nor U44726 (N_44726,N_35457,N_39511);
nand U44727 (N_44727,N_36503,N_35339);
or U44728 (N_44728,N_35885,N_35674);
xnor U44729 (N_44729,N_35497,N_35056);
or U44730 (N_44730,N_36915,N_35075);
or U44731 (N_44731,N_36053,N_37156);
and U44732 (N_44732,N_37987,N_35248);
nand U44733 (N_44733,N_35954,N_36375);
and U44734 (N_44734,N_36148,N_38134);
and U44735 (N_44735,N_38249,N_38125);
xnor U44736 (N_44736,N_35275,N_39357);
and U44737 (N_44737,N_35263,N_38536);
or U44738 (N_44738,N_35940,N_38538);
and U44739 (N_44739,N_35939,N_35338);
nor U44740 (N_44740,N_35352,N_39412);
or U44741 (N_44741,N_35745,N_35878);
and U44742 (N_44742,N_39231,N_39109);
or U44743 (N_44743,N_38410,N_37410);
nand U44744 (N_44744,N_38220,N_39737);
nand U44745 (N_44745,N_37470,N_36382);
xnor U44746 (N_44746,N_38879,N_37518);
and U44747 (N_44747,N_36111,N_38293);
or U44748 (N_44748,N_36901,N_35689);
nand U44749 (N_44749,N_36352,N_39389);
nand U44750 (N_44750,N_37942,N_38309);
nand U44751 (N_44751,N_39232,N_35391);
and U44752 (N_44752,N_36820,N_36066);
or U44753 (N_44753,N_36077,N_35558);
and U44754 (N_44754,N_35802,N_35713);
or U44755 (N_44755,N_37155,N_38111);
or U44756 (N_44756,N_37589,N_37754);
or U44757 (N_44757,N_39319,N_37798);
and U44758 (N_44758,N_36803,N_36099);
nor U44759 (N_44759,N_37958,N_35142);
xor U44760 (N_44760,N_36041,N_38248);
or U44761 (N_44761,N_38632,N_35615);
and U44762 (N_44762,N_36464,N_38321);
and U44763 (N_44763,N_38479,N_39494);
or U44764 (N_44764,N_36108,N_36459);
xor U44765 (N_44765,N_39167,N_39911);
nor U44766 (N_44766,N_39033,N_39398);
nand U44767 (N_44767,N_37282,N_37892);
or U44768 (N_44768,N_35394,N_36945);
and U44769 (N_44769,N_39998,N_38803);
nor U44770 (N_44770,N_39741,N_38554);
nand U44771 (N_44771,N_39165,N_38546);
and U44772 (N_44772,N_35506,N_36114);
nand U44773 (N_44773,N_37158,N_38727);
nand U44774 (N_44774,N_35660,N_37310);
nand U44775 (N_44775,N_35909,N_37588);
nand U44776 (N_44776,N_37838,N_35083);
or U44777 (N_44777,N_39211,N_38251);
nand U44778 (N_44778,N_36144,N_35332);
xor U44779 (N_44779,N_36619,N_39907);
and U44780 (N_44780,N_39536,N_39929);
or U44781 (N_44781,N_39365,N_35182);
xnor U44782 (N_44782,N_35267,N_37787);
xor U44783 (N_44783,N_35827,N_36637);
xor U44784 (N_44784,N_37991,N_38544);
nor U44785 (N_44785,N_36693,N_36469);
nand U44786 (N_44786,N_38605,N_38807);
nor U44787 (N_44787,N_39092,N_37371);
xor U44788 (N_44788,N_39584,N_38546);
or U44789 (N_44789,N_35391,N_36989);
xnor U44790 (N_44790,N_39046,N_36041);
xnor U44791 (N_44791,N_35394,N_37464);
nand U44792 (N_44792,N_39455,N_39135);
and U44793 (N_44793,N_37621,N_37232);
nand U44794 (N_44794,N_36413,N_37706);
or U44795 (N_44795,N_37894,N_39866);
nand U44796 (N_44796,N_37668,N_38861);
or U44797 (N_44797,N_36764,N_39496);
or U44798 (N_44798,N_39744,N_35115);
or U44799 (N_44799,N_36284,N_36975);
xnor U44800 (N_44800,N_36101,N_39887);
and U44801 (N_44801,N_39331,N_38578);
and U44802 (N_44802,N_39169,N_37536);
and U44803 (N_44803,N_37911,N_35000);
xor U44804 (N_44804,N_36750,N_36991);
or U44805 (N_44805,N_37934,N_36523);
nor U44806 (N_44806,N_39002,N_36952);
xor U44807 (N_44807,N_38982,N_35401);
xnor U44808 (N_44808,N_36770,N_36178);
nor U44809 (N_44809,N_37485,N_36951);
nor U44810 (N_44810,N_37356,N_37312);
or U44811 (N_44811,N_37348,N_37307);
and U44812 (N_44812,N_39239,N_38855);
nand U44813 (N_44813,N_35141,N_35187);
nor U44814 (N_44814,N_36679,N_36392);
or U44815 (N_44815,N_35449,N_35670);
and U44816 (N_44816,N_35277,N_36967);
xor U44817 (N_44817,N_39571,N_39685);
and U44818 (N_44818,N_37939,N_35989);
xor U44819 (N_44819,N_37109,N_38838);
and U44820 (N_44820,N_35058,N_37549);
or U44821 (N_44821,N_35594,N_35663);
xnor U44822 (N_44822,N_37364,N_36213);
or U44823 (N_44823,N_38689,N_36174);
or U44824 (N_44824,N_37387,N_36659);
nand U44825 (N_44825,N_39237,N_35166);
nand U44826 (N_44826,N_39707,N_38331);
and U44827 (N_44827,N_38121,N_38644);
nor U44828 (N_44828,N_35658,N_35815);
nor U44829 (N_44829,N_37471,N_35663);
and U44830 (N_44830,N_37470,N_36133);
and U44831 (N_44831,N_37053,N_39316);
nand U44832 (N_44832,N_36340,N_37282);
nor U44833 (N_44833,N_36517,N_35262);
nor U44834 (N_44834,N_36941,N_39564);
nor U44835 (N_44835,N_37694,N_35324);
or U44836 (N_44836,N_39505,N_38570);
nand U44837 (N_44837,N_37806,N_36105);
nor U44838 (N_44838,N_37482,N_36723);
xor U44839 (N_44839,N_39024,N_38123);
nor U44840 (N_44840,N_38278,N_37270);
and U44841 (N_44841,N_35115,N_39566);
nor U44842 (N_44842,N_38334,N_35866);
or U44843 (N_44843,N_36992,N_35683);
xor U44844 (N_44844,N_35402,N_39543);
nand U44845 (N_44845,N_37056,N_35984);
nand U44846 (N_44846,N_36326,N_36220);
nand U44847 (N_44847,N_38300,N_36550);
nand U44848 (N_44848,N_35560,N_39215);
nand U44849 (N_44849,N_36087,N_35683);
xor U44850 (N_44850,N_38623,N_37304);
or U44851 (N_44851,N_38545,N_39374);
nand U44852 (N_44852,N_36661,N_36055);
nor U44853 (N_44853,N_37567,N_37695);
and U44854 (N_44854,N_37406,N_38300);
and U44855 (N_44855,N_35514,N_36563);
xor U44856 (N_44856,N_37187,N_39843);
or U44857 (N_44857,N_36471,N_35435);
and U44858 (N_44858,N_36627,N_36506);
or U44859 (N_44859,N_36667,N_35986);
and U44860 (N_44860,N_39816,N_37072);
and U44861 (N_44861,N_38856,N_37971);
or U44862 (N_44862,N_36959,N_37606);
or U44863 (N_44863,N_39151,N_38503);
or U44864 (N_44864,N_36270,N_38589);
and U44865 (N_44865,N_35456,N_36754);
and U44866 (N_44866,N_36519,N_36353);
nor U44867 (N_44867,N_39510,N_37719);
nor U44868 (N_44868,N_39343,N_39935);
nor U44869 (N_44869,N_35424,N_37100);
nand U44870 (N_44870,N_39627,N_36977);
or U44871 (N_44871,N_36117,N_37576);
or U44872 (N_44872,N_36842,N_35964);
xnor U44873 (N_44873,N_38106,N_39590);
xor U44874 (N_44874,N_35713,N_37034);
nand U44875 (N_44875,N_37873,N_38479);
nor U44876 (N_44876,N_35253,N_39121);
nand U44877 (N_44877,N_39344,N_36273);
nor U44878 (N_44878,N_35046,N_39882);
xnor U44879 (N_44879,N_39523,N_39728);
and U44880 (N_44880,N_35558,N_39901);
and U44881 (N_44881,N_37302,N_36339);
or U44882 (N_44882,N_39038,N_37454);
and U44883 (N_44883,N_35357,N_36492);
or U44884 (N_44884,N_37381,N_38698);
xor U44885 (N_44885,N_37625,N_37685);
nand U44886 (N_44886,N_35072,N_39126);
or U44887 (N_44887,N_38160,N_38633);
xor U44888 (N_44888,N_39559,N_38488);
xnor U44889 (N_44889,N_39992,N_36077);
xor U44890 (N_44890,N_38602,N_39915);
xor U44891 (N_44891,N_36501,N_38394);
nor U44892 (N_44892,N_37498,N_35371);
and U44893 (N_44893,N_37763,N_36134);
and U44894 (N_44894,N_36269,N_35861);
or U44895 (N_44895,N_37045,N_36411);
and U44896 (N_44896,N_37846,N_35116);
or U44897 (N_44897,N_39779,N_39894);
or U44898 (N_44898,N_37501,N_36339);
or U44899 (N_44899,N_37986,N_35872);
or U44900 (N_44900,N_39628,N_38730);
and U44901 (N_44901,N_37456,N_36530);
or U44902 (N_44902,N_36063,N_35347);
or U44903 (N_44903,N_38333,N_36437);
nor U44904 (N_44904,N_37297,N_36926);
nor U44905 (N_44905,N_38696,N_36963);
xnor U44906 (N_44906,N_36289,N_37021);
or U44907 (N_44907,N_39756,N_36257);
and U44908 (N_44908,N_36189,N_38245);
or U44909 (N_44909,N_36232,N_38565);
and U44910 (N_44910,N_38974,N_35557);
nand U44911 (N_44911,N_38501,N_36295);
and U44912 (N_44912,N_36147,N_36537);
or U44913 (N_44913,N_36547,N_36200);
nor U44914 (N_44914,N_36903,N_37163);
and U44915 (N_44915,N_38830,N_38141);
and U44916 (N_44916,N_36101,N_36989);
and U44917 (N_44917,N_37963,N_36648);
xor U44918 (N_44918,N_38589,N_39158);
nand U44919 (N_44919,N_39706,N_35282);
or U44920 (N_44920,N_38116,N_35325);
nor U44921 (N_44921,N_38583,N_38427);
nand U44922 (N_44922,N_35399,N_37378);
or U44923 (N_44923,N_35393,N_38382);
nand U44924 (N_44924,N_35252,N_38243);
nor U44925 (N_44925,N_38569,N_35933);
xnor U44926 (N_44926,N_37715,N_36483);
xor U44927 (N_44927,N_38902,N_37383);
and U44928 (N_44928,N_39393,N_35263);
nand U44929 (N_44929,N_39017,N_38572);
xnor U44930 (N_44930,N_36538,N_38565);
xnor U44931 (N_44931,N_38807,N_35485);
nor U44932 (N_44932,N_37441,N_38570);
xnor U44933 (N_44933,N_38019,N_39110);
nor U44934 (N_44934,N_39955,N_37626);
nor U44935 (N_44935,N_39855,N_35839);
nand U44936 (N_44936,N_39426,N_37755);
xnor U44937 (N_44937,N_39474,N_36172);
and U44938 (N_44938,N_38697,N_37661);
nand U44939 (N_44939,N_36115,N_39197);
and U44940 (N_44940,N_39774,N_38193);
and U44941 (N_44941,N_39388,N_36146);
nand U44942 (N_44942,N_35400,N_35261);
nor U44943 (N_44943,N_36247,N_35041);
nand U44944 (N_44944,N_35048,N_37003);
xnor U44945 (N_44945,N_37651,N_36844);
nand U44946 (N_44946,N_35609,N_35588);
and U44947 (N_44947,N_39583,N_37658);
nand U44948 (N_44948,N_35528,N_36088);
or U44949 (N_44949,N_37326,N_35953);
nand U44950 (N_44950,N_35651,N_37117);
nor U44951 (N_44951,N_37715,N_36317);
nand U44952 (N_44952,N_38488,N_35290);
or U44953 (N_44953,N_36888,N_35960);
or U44954 (N_44954,N_38854,N_35945);
nand U44955 (N_44955,N_36332,N_39260);
nor U44956 (N_44956,N_38975,N_39575);
xor U44957 (N_44957,N_36007,N_36094);
nor U44958 (N_44958,N_37199,N_36711);
or U44959 (N_44959,N_38421,N_37644);
xnor U44960 (N_44960,N_36356,N_35424);
and U44961 (N_44961,N_39935,N_37442);
xnor U44962 (N_44962,N_37389,N_36826);
or U44963 (N_44963,N_37320,N_38586);
nor U44964 (N_44964,N_35217,N_39528);
nand U44965 (N_44965,N_36085,N_36005);
xnor U44966 (N_44966,N_37734,N_39275);
and U44967 (N_44967,N_38282,N_36907);
xnor U44968 (N_44968,N_38711,N_37614);
nor U44969 (N_44969,N_39557,N_38723);
nand U44970 (N_44970,N_37295,N_35467);
nor U44971 (N_44971,N_38758,N_38338);
and U44972 (N_44972,N_37775,N_39364);
xnor U44973 (N_44973,N_36373,N_39105);
nand U44974 (N_44974,N_39453,N_36044);
or U44975 (N_44975,N_35354,N_36137);
and U44976 (N_44976,N_35114,N_38225);
or U44977 (N_44977,N_37739,N_38982);
nand U44978 (N_44978,N_38191,N_38177);
nor U44979 (N_44979,N_35042,N_38904);
xnor U44980 (N_44980,N_36587,N_35160);
nor U44981 (N_44981,N_39400,N_38928);
or U44982 (N_44982,N_35480,N_37727);
nor U44983 (N_44983,N_35116,N_36506);
nor U44984 (N_44984,N_35311,N_37641);
nor U44985 (N_44985,N_37978,N_35833);
or U44986 (N_44986,N_35040,N_39995);
nor U44987 (N_44987,N_39879,N_35956);
and U44988 (N_44988,N_35765,N_37675);
and U44989 (N_44989,N_39327,N_38421);
or U44990 (N_44990,N_37356,N_35985);
nor U44991 (N_44991,N_39877,N_38251);
nand U44992 (N_44992,N_39992,N_36234);
nor U44993 (N_44993,N_39551,N_38470);
nor U44994 (N_44994,N_36885,N_35164);
nor U44995 (N_44995,N_39270,N_37084);
or U44996 (N_44996,N_38954,N_35641);
and U44997 (N_44997,N_39268,N_37805);
nand U44998 (N_44998,N_38662,N_35914);
nor U44999 (N_44999,N_37192,N_37863);
nor U45000 (N_45000,N_41803,N_44324);
nor U45001 (N_45001,N_40449,N_43142);
nand U45002 (N_45002,N_40156,N_43727);
nor U45003 (N_45003,N_43716,N_42738);
nor U45004 (N_45004,N_42898,N_40792);
xor U45005 (N_45005,N_44614,N_42355);
nor U45006 (N_45006,N_42585,N_42861);
xnor U45007 (N_45007,N_44077,N_43427);
nor U45008 (N_45008,N_43907,N_42977);
xnor U45009 (N_45009,N_41106,N_43406);
nor U45010 (N_45010,N_41277,N_42157);
nor U45011 (N_45011,N_41767,N_40136);
and U45012 (N_45012,N_44251,N_44790);
or U45013 (N_45013,N_41785,N_41701);
nand U45014 (N_45014,N_42628,N_43107);
nor U45015 (N_45015,N_43238,N_40656);
or U45016 (N_45016,N_44144,N_41759);
and U45017 (N_45017,N_41680,N_40640);
nor U45018 (N_45018,N_41020,N_40161);
and U45019 (N_45019,N_40668,N_42587);
and U45020 (N_45020,N_40070,N_43363);
nor U45021 (N_45021,N_43531,N_43969);
nand U45022 (N_45022,N_40850,N_44892);
nand U45023 (N_45023,N_42349,N_43000);
or U45024 (N_45024,N_43008,N_43063);
nand U45025 (N_45025,N_41225,N_43634);
and U45026 (N_45026,N_40326,N_41597);
nor U45027 (N_45027,N_42932,N_40886);
or U45028 (N_45028,N_41594,N_42900);
nand U45029 (N_45029,N_43143,N_40721);
nand U45030 (N_45030,N_43391,N_40968);
nand U45031 (N_45031,N_44985,N_44793);
and U45032 (N_45032,N_43691,N_43661);
nand U45033 (N_45033,N_42896,N_42950);
xnor U45034 (N_45034,N_40686,N_43185);
nor U45035 (N_45035,N_41426,N_44581);
nor U45036 (N_45036,N_44554,N_43575);
nand U45037 (N_45037,N_44270,N_42528);
and U45038 (N_45038,N_44908,N_42229);
or U45039 (N_45039,N_44692,N_42087);
nor U45040 (N_45040,N_42792,N_42142);
xnor U45041 (N_45041,N_40999,N_44607);
nand U45042 (N_45042,N_42639,N_40025);
nand U45043 (N_45043,N_41578,N_40048);
and U45044 (N_45044,N_43930,N_40678);
nor U45045 (N_45045,N_42652,N_42375);
nor U45046 (N_45046,N_40798,N_42991);
and U45047 (N_45047,N_41044,N_44474);
nor U45048 (N_45048,N_43748,N_44584);
or U45049 (N_45049,N_43120,N_44434);
and U45050 (N_45050,N_40364,N_43830);
nor U45051 (N_45051,N_43042,N_40173);
xor U45052 (N_45052,N_43561,N_40116);
nor U45053 (N_45053,N_42957,N_43591);
nor U45054 (N_45054,N_43933,N_42687);
or U45055 (N_45055,N_40357,N_43659);
or U45056 (N_45056,N_40179,N_42338);
xor U45057 (N_45057,N_42227,N_40024);
nor U45058 (N_45058,N_43781,N_44522);
nand U45059 (N_45059,N_40914,N_40500);
nand U45060 (N_45060,N_43594,N_40995);
and U45061 (N_45061,N_40741,N_41097);
xnor U45062 (N_45062,N_40994,N_40008);
or U45063 (N_45063,N_41949,N_44178);
and U45064 (N_45064,N_43465,N_44127);
and U45065 (N_45065,N_44103,N_43168);
nand U45066 (N_45066,N_40910,N_41994);
xor U45067 (N_45067,N_40300,N_43192);
or U45068 (N_45068,N_44083,N_41929);
nand U45069 (N_45069,N_42303,N_42299);
xor U45070 (N_45070,N_40313,N_44316);
and U45071 (N_45071,N_43570,N_42640);
nand U45072 (N_45072,N_41220,N_43341);
nand U45073 (N_45073,N_41304,N_42678);
nor U45074 (N_45074,N_41454,N_44646);
xor U45075 (N_45075,N_40318,N_42698);
nand U45076 (N_45076,N_42093,N_41029);
nand U45077 (N_45077,N_43383,N_41408);
nand U45078 (N_45078,N_43095,N_41493);
and U45079 (N_45079,N_40354,N_43509);
nor U45080 (N_45080,N_43750,N_44188);
nand U45081 (N_45081,N_44478,N_40906);
xor U45082 (N_45082,N_43652,N_43048);
and U45083 (N_45083,N_40895,N_44571);
nand U45084 (N_45084,N_42966,N_41703);
or U45085 (N_45085,N_43843,N_44219);
nor U45086 (N_45086,N_40029,N_41471);
nor U45087 (N_45087,N_41821,N_41887);
nand U45088 (N_45088,N_43084,N_41572);
and U45089 (N_45089,N_42124,N_40918);
nand U45090 (N_45090,N_40031,N_40998);
xnor U45091 (N_45091,N_40432,N_43963);
and U45092 (N_45092,N_43765,N_44413);
or U45093 (N_45093,N_44123,N_42472);
or U45094 (N_45094,N_43223,N_43773);
xor U45095 (N_45095,N_42336,N_41792);
nor U45096 (N_45096,N_41971,N_41831);
or U45097 (N_45097,N_42503,N_41663);
nand U45098 (N_45098,N_44895,N_40295);
or U45099 (N_45099,N_44021,N_43728);
or U45100 (N_45100,N_43221,N_42507);
nor U45101 (N_45101,N_42421,N_41352);
nor U45102 (N_45102,N_40377,N_41836);
nand U45103 (N_45103,N_40426,N_44559);
xnor U45104 (N_45104,N_44394,N_40080);
nor U45105 (N_45105,N_41183,N_44027);
nor U45106 (N_45106,N_44719,N_41439);
and U45107 (N_45107,N_44408,N_42513);
nor U45108 (N_45108,N_44982,N_44670);
nand U45109 (N_45109,N_43167,N_43187);
nor U45110 (N_45110,N_41835,N_40203);
and U45111 (N_45111,N_42886,N_41468);
or U45112 (N_45112,N_43301,N_40127);
or U45113 (N_45113,N_42965,N_42176);
nor U45114 (N_45114,N_41688,N_41743);
nand U45115 (N_45115,N_41945,N_43605);
nand U45116 (N_45116,N_43190,N_44940);
nor U45117 (N_45117,N_41430,N_41462);
xor U45118 (N_45118,N_43157,N_42582);
nand U45119 (N_45119,N_42137,N_42048);
nand U45120 (N_45120,N_40244,N_41769);
and U45121 (N_45121,N_41478,N_42213);
nand U45122 (N_45122,N_40246,N_41437);
or U45123 (N_45123,N_44582,N_43809);
nand U45124 (N_45124,N_42813,N_43711);
xnor U45125 (N_45125,N_41187,N_42818);
or U45126 (N_45126,N_44966,N_44978);
nand U45127 (N_45127,N_42757,N_42829);
and U45128 (N_45128,N_43239,N_42367);
or U45129 (N_45129,N_41169,N_42429);
nor U45130 (N_45130,N_43184,N_42262);
and U45131 (N_45131,N_40984,N_43318);
nand U45132 (N_45132,N_41240,N_41820);
and U45133 (N_45133,N_42415,N_40261);
nor U45134 (N_45134,N_44296,N_41391);
xor U45135 (N_45135,N_40967,N_41230);
nor U45136 (N_45136,N_44638,N_43483);
nand U45137 (N_45137,N_41376,N_41285);
nor U45138 (N_45138,N_40360,N_42990);
nor U45139 (N_45139,N_44820,N_40302);
nand U45140 (N_45140,N_41823,N_40996);
and U45141 (N_45141,N_41103,N_44004);
nor U45142 (N_45142,N_41637,N_44082);
nor U45143 (N_45143,N_42378,N_43276);
and U45144 (N_45144,N_40617,N_41214);
and U45145 (N_45145,N_41699,N_44336);
nand U45146 (N_45146,N_41907,N_41709);
nor U45147 (N_45147,N_40130,N_41908);
and U45148 (N_45148,N_43090,N_43672);
or U45149 (N_45149,N_42455,N_41655);
nand U45150 (N_45150,N_44859,N_43795);
or U45151 (N_45151,N_43714,N_42023);
or U45152 (N_45152,N_42890,N_40780);
nand U45153 (N_45153,N_43996,N_40233);
xor U45154 (N_45154,N_44403,N_43958);
xor U45155 (N_45155,N_42835,N_43360);
nor U45156 (N_45156,N_44730,N_44871);
and U45157 (N_45157,N_41257,N_42434);
and U45158 (N_45158,N_42233,N_41399);
xnor U45159 (N_45159,N_42959,N_40495);
xor U45160 (N_45160,N_42939,N_42269);
xor U45161 (N_45161,N_41174,N_40832);
nand U45162 (N_45162,N_40503,N_41777);
nand U45163 (N_45163,N_44222,N_41719);
or U45164 (N_45164,N_41824,N_42834);
xnor U45165 (N_45165,N_41969,N_42770);
nor U45166 (N_45166,N_44665,N_44393);
nor U45167 (N_45167,N_41425,N_44079);
nor U45168 (N_45168,N_40180,N_43987);
or U45169 (N_45169,N_40768,N_41898);
and U45170 (N_45170,N_43226,N_40211);
nand U45171 (N_45171,N_43548,N_43989);
and U45172 (N_45172,N_42833,N_43611);
nand U45173 (N_45173,N_41390,N_42481);
or U45174 (N_45174,N_43068,N_44031);
nand U45175 (N_45175,N_41062,N_44532);
and U45176 (N_45176,N_44736,N_42758);
or U45177 (N_45177,N_41291,N_40079);
xor U45178 (N_45178,N_44242,N_40873);
and U45179 (N_45179,N_43701,N_42292);
or U45180 (N_45180,N_43032,N_43447);
and U45181 (N_45181,N_42926,N_42712);
xnor U45182 (N_45182,N_40598,N_42619);
nand U45183 (N_45183,N_40271,N_42419);
and U45184 (N_45184,N_42425,N_41166);
nor U45185 (N_45185,N_40767,N_42032);
or U45186 (N_45186,N_42901,N_42734);
or U45187 (N_45187,N_42380,N_41005);
xor U45188 (N_45188,N_42623,N_40400);
xnor U45189 (N_45189,N_41032,N_44808);
nor U45190 (N_45190,N_43816,N_41923);
nor U45191 (N_45191,N_44570,N_44436);
nand U45192 (N_45192,N_44273,N_43999);
or U45193 (N_45193,N_42632,N_44204);
nand U45194 (N_45194,N_41822,N_42099);
nand U45195 (N_45195,N_43027,N_43094);
or U45196 (N_45196,N_41300,N_44964);
nand U45197 (N_45197,N_41992,N_41617);
or U45198 (N_45198,N_40328,N_43164);
xnor U45199 (N_45199,N_42307,N_43857);
and U45200 (N_45200,N_41316,N_42591);
nand U45201 (N_45201,N_43343,N_42874);
or U45202 (N_45202,N_40698,N_42431);
nand U45203 (N_45203,N_42557,N_40557);
or U45204 (N_45204,N_44851,N_43233);
nand U45205 (N_45205,N_41827,N_43369);
nor U45206 (N_45206,N_42502,N_41515);
and U45207 (N_45207,N_40213,N_43799);
or U45208 (N_45208,N_42613,N_40085);
xor U45209 (N_45209,N_44277,N_42988);
nand U45210 (N_45210,N_44025,N_43662);
nor U45211 (N_45211,N_41560,N_41223);
nand U45212 (N_45212,N_43950,N_41746);
nand U45213 (N_45213,N_41529,N_44564);
nor U45214 (N_45214,N_43904,N_40695);
nand U45215 (N_45215,N_44893,N_41484);
or U45216 (N_45216,N_43956,N_40111);
nand U45217 (N_45217,N_42516,N_42040);
nand U45218 (N_45218,N_40389,N_42746);
nand U45219 (N_45219,N_40565,N_42645);
and U45220 (N_45220,N_41059,N_41903);
or U45221 (N_45221,N_42987,N_42948);
or U45222 (N_45222,N_44843,N_41664);
and U45223 (N_45223,N_42270,N_44090);
nor U45224 (N_45224,N_41446,N_40572);
nand U45225 (N_45225,N_40710,N_43231);
xnor U45226 (N_45226,N_41937,N_40359);
xor U45227 (N_45227,N_40883,N_40724);
xor U45228 (N_45228,N_43050,N_43814);
and U45229 (N_45229,N_44742,N_41299);
and U45230 (N_45230,N_42290,N_40128);
xnor U45231 (N_45231,N_42050,N_44891);
nand U45232 (N_45232,N_43484,N_42410);
nor U45233 (N_45233,N_41555,N_40846);
nand U45234 (N_45234,N_42065,N_40081);
nand U45235 (N_45235,N_42963,N_44124);
nor U45236 (N_45236,N_44604,N_43450);
xor U45237 (N_45237,N_43299,N_44725);
xnor U45238 (N_45238,N_42786,N_42817);
nor U45239 (N_45239,N_40073,N_41619);
or U45240 (N_45240,N_43928,N_44148);
xor U45241 (N_45241,N_42542,N_44252);
or U45242 (N_45242,N_40087,N_41041);
nand U45243 (N_45243,N_44932,N_40441);
or U45244 (N_45244,N_43518,N_43873);
and U45245 (N_45245,N_43466,N_43539);
nor U45246 (N_45246,N_44310,N_43758);
xor U45247 (N_45247,N_42360,N_41412);
nand U45248 (N_45248,N_44331,N_40657);
xor U45249 (N_45249,N_44605,N_44929);
xor U45250 (N_45250,N_41339,N_43644);
nor U45251 (N_45251,N_40607,N_44190);
nand U45252 (N_45252,N_42740,N_41119);
nand U45253 (N_45253,N_42268,N_40763);
and U45254 (N_45254,N_44923,N_43086);
nor U45255 (N_45255,N_44107,N_40017);
nand U45256 (N_45256,N_44187,N_40206);
nor U45257 (N_45257,N_43395,N_42521);
or U45258 (N_45258,N_41802,N_42705);
xor U45259 (N_45259,N_43024,N_43170);
and U45260 (N_45260,N_42531,N_40049);
and U45261 (N_45261,N_42924,N_41142);
or U45262 (N_45262,N_44257,N_44800);
xor U45263 (N_45263,N_42940,N_40866);
xnor U45264 (N_45264,N_41361,N_44563);
or U45265 (N_45265,N_44971,N_42112);
nor U45266 (N_45266,N_41817,N_43625);
and U45267 (N_45267,N_43074,N_44778);
xor U45268 (N_45268,N_43235,N_44879);
nor U45269 (N_45269,N_42524,N_41852);
nand U45270 (N_45270,N_44922,N_43984);
nor U45271 (N_45271,N_40347,N_44530);
xnor U45272 (N_45272,N_42034,N_43284);
nor U45273 (N_45273,N_41837,N_41863);
nor U45274 (N_45274,N_44452,N_44467);
xnor U45275 (N_45275,N_41222,N_43797);
nand U45276 (N_45276,N_40473,N_43475);
and U45277 (N_45277,N_41781,N_40667);
or U45278 (N_45278,N_43257,N_40493);
xor U45279 (N_45279,N_40286,N_41203);
and U45280 (N_45280,N_40920,N_43893);
nor U45281 (N_45281,N_41348,N_40939);
nor U45282 (N_45282,N_42993,N_42201);
nand U45283 (N_45283,N_43455,N_44876);
xor U45284 (N_45284,N_41283,N_40590);
nand U45285 (N_45285,N_43126,N_44295);
nand U45286 (N_45286,N_41089,N_44326);
nor U45287 (N_45287,N_42897,N_41087);
nand U45288 (N_45288,N_41509,N_41268);
nor U45289 (N_45289,N_44873,N_41482);
and U45290 (N_45290,N_41789,N_40799);
xor U45291 (N_45291,N_41301,N_44802);
nand U45292 (N_45292,N_43290,N_43827);
nor U45293 (N_45293,N_44321,N_43583);
or U45294 (N_45294,N_41900,N_42567);
xor U45295 (N_45295,N_44823,N_42188);
nor U45296 (N_45296,N_43708,N_43016);
xnor U45297 (N_45297,N_40163,N_41736);
nor U45298 (N_45298,N_41094,N_40708);
nor U45299 (N_45299,N_41448,N_40988);
xnor U45300 (N_45300,N_43679,N_43053);
and U45301 (N_45301,N_40675,N_40339);
or U45302 (N_45302,N_40228,N_43218);
nor U45303 (N_45303,N_40982,N_41807);
nor U45304 (N_45304,N_40570,N_42830);
nor U45305 (N_45305,N_42782,N_44312);
and U45306 (N_45306,N_44469,N_44958);
and U45307 (N_45307,N_43131,N_44414);
xnor U45308 (N_45308,N_43717,N_43906);
nand U45309 (N_45309,N_42005,N_43327);
nand U45310 (N_45310,N_44780,N_42529);
or U45311 (N_45311,N_41595,N_40153);
nand U45312 (N_45312,N_40577,N_43515);
and U45313 (N_45313,N_42826,N_40759);
xor U45314 (N_45314,N_40146,N_40843);
xor U45315 (N_45315,N_42994,N_43640);
nor U45316 (N_45316,N_42356,N_40809);
nand U45317 (N_45317,N_40453,N_40977);
nand U45318 (N_45318,N_44387,N_42892);
or U45319 (N_45319,N_42092,N_41327);
or U45320 (N_45320,N_40663,N_42559);
and U45321 (N_45321,N_41760,N_44032);
and U45322 (N_45322,N_43490,N_41710);
nor U45323 (N_45323,N_41685,N_42469);
or U45324 (N_45324,N_44239,N_40069);
or U45325 (N_45325,N_42575,N_44629);
or U45326 (N_45326,N_43722,N_42851);
nor U45327 (N_45327,N_40502,N_43771);
nor U45328 (N_45328,N_40641,N_40397);
nor U45329 (N_45329,N_41978,N_43558);
and U45330 (N_45330,N_44630,N_44133);
and U45331 (N_45331,N_43966,N_41137);
nand U45332 (N_45332,N_44608,N_44221);
or U45333 (N_45333,N_42009,N_44975);
or U45334 (N_45334,N_43034,N_40310);
and U45335 (N_45335,N_42372,N_40393);
and U45336 (N_45336,N_43333,N_42018);
nor U45337 (N_45337,N_44134,N_44718);
xnor U45338 (N_45338,N_43638,N_44381);
nand U45339 (N_45339,N_44696,N_40789);
nor U45340 (N_45340,N_44244,N_43039);
nand U45341 (N_45341,N_44363,N_44451);
or U45342 (N_45342,N_43564,N_42797);
xor U45343 (N_45343,N_42553,N_42510);
nand U45344 (N_45344,N_41157,N_42533);
xnor U45345 (N_45345,N_44415,N_41386);
xor U45346 (N_45346,N_41265,N_43791);
xnor U45347 (N_45347,N_44535,N_44442);
and U45348 (N_45348,N_43394,N_42416);
nor U45349 (N_45349,N_43473,N_43277);
nor U45350 (N_45350,N_42703,N_40257);
nand U45351 (N_45351,N_41933,N_44553);
or U45352 (N_45352,N_43497,N_41856);
and U45353 (N_45353,N_44741,N_41093);
nor U45354 (N_45354,N_41770,N_43952);
and U45355 (N_45355,N_42337,N_42848);
nor U45356 (N_45356,N_40838,N_41197);
and U45357 (N_45357,N_43865,N_43668);
nor U45358 (N_45358,N_40512,N_42461);
nor U45359 (N_45359,N_44249,N_44155);
nor U45360 (N_45360,N_42985,N_44946);
nand U45361 (N_45361,N_40330,N_42354);
or U45362 (N_45362,N_44151,N_44831);
nor U45363 (N_45363,N_44645,N_43020);
or U45364 (N_45364,N_42244,N_44115);
or U45365 (N_45365,N_41522,N_41344);
and U45366 (N_45366,N_41828,N_44575);
xnor U45367 (N_45367,N_41422,N_41015);
or U45368 (N_45368,N_42265,N_40777);
xor U45369 (N_45369,N_41131,N_41158);
or U45370 (N_45370,N_40517,N_43424);
xnor U45371 (N_45371,N_41264,N_42891);
and U45372 (N_45372,N_40676,N_40221);
or U45373 (N_45373,N_41645,N_42550);
nor U45374 (N_45374,N_40787,N_41403);
nand U45375 (N_45375,N_41483,N_41566);
or U45376 (N_45376,N_41259,N_43241);
nand U45377 (N_45377,N_40576,N_43596);
and U45378 (N_45378,N_40791,N_40120);
xor U45379 (N_45379,N_42719,N_41204);
xnor U45380 (N_45380,N_42535,N_44139);
nor U45381 (N_45381,N_41512,N_44091);
or U45382 (N_45382,N_40195,N_40134);
nand U45383 (N_45383,N_43295,N_42821);
or U45384 (N_45384,N_41149,N_42970);
xor U45385 (N_45385,N_42181,N_44954);
and U45386 (N_45386,N_40804,N_43098);
nand U45387 (N_45387,N_44158,N_43657);
and U45388 (N_45388,N_41700,N_42011);
nor U45389 (N_45389,N_43001,N_42089);
xnor U45390 (N_45390,N_43478,N_40814);
nand U45391 (N_45391,N_44087,N_40445);
nor U45392 (N_45392,N_40215,N_41748);
and U45393 (N_45393,N_43097,N_44416);
xnor U45394 (N_45394,N_44334,N_43542);
xnor U45395 (N_45395,N_41440,N_40618);
or U45396 (N_45396,N_42444,N_43026);
xnor U45397 (N_45397,N_41254,N_40979);
xnor U45398 (N_45398,N_44437,N_41724);
nand U45399 (N_45399,N_44636,N_44482);
nand U45400 (N_45400,N_43643,N_40496);
nand U45401 (N_45401,N_41884,N_41882);
xor U45402 (N_45402,N_43477,N_44346);
and U45403 (N_45403,N_42175,N_42808);
xnor U45404 (N_45404,N_44086,N_44853);
or U45405 (N_45405,N_43543,N_43352);
or U45406 (N_45406,N_44597,N_40929);
nand U45407 (N_45407,N_41191,N_44981);
xor U45408 (N_45408,N_42390,N_40702);
nor U45409 (N_45409,N_44701,N_43201);
nor U45410 (N_45410,N_42986,N_43410);
and U45411 (N_45411,N_44603,N_41847);
or U45412 (N_45412,N_40363,N_43182);
nand U45413 (N_45413,N_40857,N_41541);
or U45414 (N_45414,N_43140,N_43871);
or U45415 (N_45415,N_44201,N_43313);
xor U45416 (N_45416,N_44766,N_42788);
nor U45417 (N_45417,N_40416,N_40961);
xor U45418 (N_45418,N_40027,N_43066);
xnor U45419 (N_45419,N_41885,N_41378);
and U45420 (N_45420,N_42031,N_44905);
or U45421 (N_45421,N_40946,N_42779);
and U45422 (N_45422,N_44835,N_44506);
and U45423 (N_45423,N_40434,N_42766);
or U45424 (N_45424,N_41894,N_44913);
nand U45425 (N_45425,N_43077,N_43516);
nand U45426 (N_45426,N_41590,N_40872);
nor U45427 (N_45427,N_44776,N_43637);
nor U45428 (N_45428,N_44883,N_42304);
nand U45429 (N_45429,N_44501,N_41346);
nor U45430 (N_45430,N_40683,N_44162);
xor U45431 (N_45431,N_40482,N_42974);
nor U45432 (N_45432,N_42569,N_41369);
nand U45433 (N_45433,N_42106,N_44003);
and U45434 (N_45434,N_40338,N_42715);
and U45435 (N_45435,N_43929,N_41586);
xor U45436 (N_45436,N_44832,N_44305);
nand U45437 (N_45437,N_40608,N_41549);
or U45438 (N_45438,N_40202,N_44611);
or U45439 (N_45439,N_42667,N_43537);
nor U45440 (N_45440,N_44392,N_40964);
nor U45441 (N_45441,N_44283,N_40862);
or U45442 (N_45442,N_44746,N_40187);
xor U45443 (N_45443,N_41311,N_41199);
nor U45444 (N_45444,N_44948,N_42206);
xor U45445 (N_45445,N_40865,N_42036);
and U45446 (N_45446,N_40349,N_40431);
and U45447 (N_45447,N_40372,N_44837);
nor U45448 (N_45448,N_43677,N_43686);
and U45449 (N_45449,N_40537,N_42230);
nor U45450 (N_45450,N_41620,N_44238);
nand U45451 (N_45451,N_42847,N_40278);
and U45452 (N_45452,N_44870,N_42895);
and U45453 (N_45453,N_41442,N_42660);
and U45454 (N_45454,N_42656,N_44752);
nand U45455 (N_45455,N_40481,N_44212);
nand U45456 (N_45456,N_42505,N_40197);
and U45457 (N_45457,N_43739,N_41782);
xor U45458 (N_45458,N_41936,N_43832);
or U45459 (N_45459,N_44796,N_42311);
and U45460 (N_45460,N_42456,N_43111);
nor U45461 (N_45461,N_42998,N_43368);
nand U45462 (N_45462,N_43236,N_44762);
or U45463 (N_45463,N_40299,N_42228);
nor U45464 (N_45464,N_43022,N_40256);
or U45465 (N_45465,N_43180,N_44685);
nor U45466 (N_45466,N_40986,N_41658);
xnor U45467 (N_45467,N_41098,N_44720);
or U45468 (N_45468,N_40797,N_43009);
nor U45469 (N_45469,N_40561,N_42055);
nor U45470 (N_45470,N_44269,N_41647);
and U45471 (N_45471,N_41979,N_44666);
or U45472 (N_45472,N_40619,N_40279);
nand U45473 (N_45473,N_44227,N_41355);
xor U45474 (N_45474,N_40638,N_41527);
nor U45475 (N_45475,N_41622,N_44217);
nand U45476 (N_45476,N_40821,N_42135);
nand U45477 (N_45477,N_40362,N_40424);
or U45478 (N_45478,N_43782,N_43839);
xor U45479 (N_45479,N_44261,N_40855);
nand U45480 (N_45480,N_42702,N_43138);
xor U45481 (N_45481,N_43908,N_41922);
xor U45482 (N_45482,N_44754,N_41871);
nor U45483 (N_45483,N_44423,N_40358);
nor U45484 (N_45484,N_41548,N_42508);
xor U45485 (N_45485,N_40365,N_40823);
or U45486 (N_45486,N_44682,N_42573);
and U45487 (N_45487,N_43064,N_40186);
and U45488 (N_45488,N_44957,N_40788);
and U45489 (N_45489,N_42867,N_40192);
or U45490 (N_45490,N_44229,N_43106);
nand U45491 (N_45491,N_40267,N_43569);
nand U45492 (N_45492,N_40375,N_43715);
nand U45493 (N_45493,N_42643,N_43801);
and U45494 (N_45494,N_42625,N_42723);
or U45495 (N_45495,N_43413,N_44081);
or U45496 (N_45496,N_41668,N_44468);
nor U45497 (N_45497,N_40019,N_40520);
xor U45498 (N_45498,N_43085,N_40505);
or U45499 (N_45499,N_40296,N_41393);
nor U45500 (N_45500,N_42713,N_43041);
xor U45501 (N_45501,N_40485,N_44440);
nand U45502 (N_45502,N_44255,N_42881);
xor U45503 (N_45503,N_44345,N_40930);
nand U45504 (N_45504,N_44919,N_41128);
nor U45505 (N_45505,N_42246,N_40926);
nand U45506 (N_45506,N_42312,N_42611);
nor U45507 (N_45507,N_43471,N_44502);
nor U45508 (N_45508,N_42308,N_40881);
xnor U45509 (N_45509,N_40987,N_42448);
or U45510 (N_45510,N_40867,N_44073);
or U45511 (N_45511,N_43927,N_44174);
nor U45512 (N_45512,N_40610,N_41262);
and U45513 (N_45513,N_42838,N_40553);
and U45514 (N_45514,N_44126,N_41841);
or U45515 (N_45515,N_41049,N_43980);
xnor U45516 (N_45516,N_44199,N_41463);
nand U45517 (N_45517,N_40115,N_42411);
or U45518 (N_45518,N_41771,N_43292);
nand U45519 (N_45519,N_43937,N_44700);
xnor U45520 (N_45520,N_43453,N_42844);
xor U45521 (N_45521,N_44119,N_44196);
and U45522 (N_45522,N_44355,N_43227);
and U45523 (N_45523,N_40046,N_44066);
or U45524 (N_45524,N_40117,N_43486);
or U45525 (N_45525,N_43469,N_42389);
nor U45526 (N_45526,N_41568,N_44484);
and U45527 (N_45527,N_43964,N_44848);
or U45528 (N_45528,N_40697,N_41004);
and U45529 (N_45529,N_40784,N_42856);
and U45530 (N_45530,N_41891,N_44896);
nand U45531 (N_45531,N_42497,N_44030);
or U45532 (N_45532,N_43361,N_41576);
nand U45533 (N_45533,N_42294,N_41684);
and U45534 (N_45534,N_43109,N_44218);
nor U45535 (N_45535,N_44904,N_44325);
and U45536 (N_45536,N_42935,N_41155);
xor U45537 (N_45537,N_43960,N_40971);
or U45538 (N_45538,N_40185,N_43713);
nand U45539 (N_45539,N_41865,N_44005);
nor U45540 (N_45540,N_42382,N_43353);
nand U45541 (N_45541,N_41633,N_44294);
xnor U45542 (N_45542,N_42618,N_44189);
nor U45543 (N_45543,N_44993,N_42215);
nor U45544 (N_45544,N_43630,N_41953);
xnor U45545 (N_45545,N_44552,N_43399);
xnor U45546 (N_45546,N_42754,N_40421);
xor U45547 (N_45547,N_42804,N_43806);
xor U45548 (N_45548,N_41205,N_43513);
or U45549 (N_45549,N_44001,N_41053);
nor U45550 (N_45550,N_42218,N_40074);
nand U45551 (N_45551,N_44263,N_40344);
nand U45552 (N_45552,N_40727,N_41470);
xnor U45553 (N_45553,N_41652,N_42657);
and U45554 (N_45554,N_42622,N_42658);
xnor U45555 (N_45555,N_44592,N_41851);
nor U45556 (N_45556,N_40371,N_44444);
or U45557 (N_45557,N_44536,N_41774);
nand U45558 (N_45558,N_44952,N_43262);
xnor U45559 (N_45559,N_42665,N_41670);
and U45560 (N_45560,N_42605,N_43563);
or U45561 (N_45561,N_44500,N_41513);
xor U45562 (N_45562,N_40616,N_40324);
nor U45563 (N_45563,N_40191,N_44292);
nor U45564 (N_45564,N_40103,N_44276);
nor U45565 (N_45565,N_41031,N_42037);
and U45566 (N_45566,N_40658,N_42743);
and U45567 (N_45567,N_43909,N_41310);
nor U45568 (N_45568,N_43642,N_43196);
nand U45569 (N_45569,N_43636,N_43462);
and U45570 (N_45570,N_42334,N_44191);
and U45571 (N_45571,N_42096,N_40222);
nand U45572 (N_45572,N_43697,N_41564);
or U45573 (N_45573,N_41876,N_40793);
nand U45574 (N_45574,N_43670,N_41069);
nor U45575 (N_45575,N_44590,N_43334);
nor U45576 (N_45576,N_44529,N_44909);
nand U45577 (N_45577,N_44770,N_42841);
or U45578 (N_45578,N_42972,N_42223);
and U45579 (N_45579,N_40735,N_44301);
or U45580 (N_45580,N_40662,N_41245);
nand U45581 (N_45581,N_42546,N_40370);
xnor U45582 (N_45582,N_44105,N_41932);
and U45583 (N_45583,N_41628,N_43061);
nor U45584 (N_45584,N_42954,N_40475);
nor U45585 (N_45585,N_44344,N_43267);
and U45586 (N_45586,N_42919,N_40586);
nor U45587 (N_45587,N_40142,N_43524);
nor U45588 (N_45588,N_44280,N_44361);
xnor U45589 (N_45589,N_42289,N_42365);
nand U45590 (N_45590,N_43379,N_44298);
nand U45591 (N_45591,N_44460,N_42133);
or U45592 (N_45592,N_41196,N_41551);
nor U45593 (N_45593,N_42594,N_44058);
nor U45594 (N_45594,N_41397,N_40852);
xor U45595 (N_45595,N_40086,N_40263);
xor U45596 (N_45596,N_40585,N_41261);
nor U45597 (N_45597,N_44816,N_40593);
nor U45598 (N_45598,N_44372,N_43559);
nor U45599 (N_45599,N_43618,N_42610);
nor U45600 (N_45600,N_41946,N_43199);
xnor U45601 (N_45601,N_42342,N_40670);
and U45602 (N_45602,N_42589,N_41721);
nand U45603 (N_45603,N_43225,N_40054);
nand U45604 (N_45604,N_40224,N_41466);
nand U45605 (N_45605,N_43680,N_40223);
and U45606 (N_45606,N_44250,N_43556);
nand U45607 (N_45607,N_42199,N_41375);
xnor U45608 (N_45608,N_40584,N_42849);
or U45609 (N_45609,N_44568,N_44878);
nor U45610 (N_45610,N_43818,N_42775);
xnor U45611 (N_45611,N_44704,N_41100);
nand U45612 (N_45612,N_40107,N_43141);
and U45613 (N_45613,N_43617,N_40887);
and U45614 (N_45614,N_43738,N_40468);
nand U45615 (N_45615,N_43674,N_42739);
nand U45616 (N_45616,N_42316,N_40808);
and U45617 (N_45617,N_40776,N_44579);
and U45618 (N_45618,N_44495,N_43057);
and U45619 (N_45619,N_43891,N_42864);
xnor U45620 (N_45620,N_40489,N_41113);
and U45621 (N_45621,N_43358,N_41786);
xnor U45622 (N_45622,N_44359,N_40205);
nand U45623 (N_45623,N_40401,N_42080);
or U45624 (N_45624,N_41571,N_42664);
and U45625 (N_45625,N_42068,N_40891);
and U45626 (N_45626,N_44961,N_42061);
or U45627 (N_45627,N_42615,N_43510);
nand U45628 (N_45628,N_40923,N_43994);
and U45629 (N_45629,N_41780,N_43317);
nand U45630 (N_45630,N_40108,N_44547);
or U45631 (N_45631,N_44152,N_41910);
xnor U45632 (N_45632,N_43892,N_43608);
xnor U45633 (N_45633,N_44633,N_41502);
nor U45634 (N_45634,N_43349,N_44877);
or U45635 (N_45635,N_44095,N_42807);
xor U45636 (N_45636,N_44748,N_40309);
and U45637 (N_45637,N_41826,N_43408);
xnor U45638 (N_45638,N_43298,N_42785);
and U45639 (N_45639,N_40497,N_42043);
or U45640 (N_45640,N_41368,N_41606);
xor U45641 (N_45641,N_42899,N_43260);
or U45642 (N_45642,N_42637,N_42200);
nor U45643 (N_45643,N_42725,N_43757);
or U45644 (N_45644,N_43002,N_42801);
and U45645 (N_45645,N_42933,N_41656);
xnor U45646 (N_45646,N_40602,N_41926);
and U45647 (N_45647,N_41123,N_42260);
nor U45648 (N_45648,N_44192,N_44839);
nor U45649 (N_45649,N_44268,N_40249);
xnor U45650 (N_45650,N_44100,N_40169);
xor U45651 (N_45651,N_43663,N_44672);
xor U45652 (N_45652,N_41133,N_43222);
xor U45653 (N_45653,N_40225,N_41194);
nor U45654 (N_45654,N_44690,N_41866);
or U45655 (N_45655,N_40643,N_43500);
xor U45656 (N_45656,N_44247,N_41998);
nor U45657 (N_45657,N_41707,N_44236);
and U45658 (N_45658,N_44002,N_41795);
nand U45659 (N_45659,N_43529,N_42127);
or U45660 (N_45660,N_42267,N_41381);
xnor U45661 (N_45661,N_43894,N_41485);
nand U45662 (N_45662,N_41705,N_40239);
and U45663 (N_45663,N_43848,N_44120);
xor U45664 (N_45664,N_40293,N_42647);
nor U45665 (N_45665,N_42682,N_42937);
nor U45666 (N_45666,N_44914,N_44714);
nor U45667 (N_45667,N_43280,N_40088);
xor U45668 (N_45668,N_40583,N_41218);
xor U45669 (N_45669,N_40292,N_43229);
and U45670 (N_45670,N_44309,N_44850);
or U45671 (N_45671,N_40262,N_40337);
xor U45672 (N_45672,N_41122,N_43501);
and U45673 (N_45673,N_42491,N_40280);
nand U45674 (N_45674,N_43153,N_41279);
xnor U45675 (N_45675,N_44223,N_43756);
nand U45676 (N_45676,N_41959,N_41068);
or U45677 (N_45677,N_43420,N_40738);
nor U45678 (N_45678,N_44572,N_44821);
or U45679 (N_45679,N_44694,N_40283);
and U45680 (N_45680,N_41373,N_43442);
xor U45681 (N_45681,N_40830,N_41110);
or U45682 (N_45682,N_43841,N_42208);
xor U45683 (N_45683,N_44065,N_41109);
and U45684 (N_45684,N_42275,N_43978);
and U45685 (N_45685,N_44388,N_41829);
xor U45686 (N_45686,N_42257,N_44531);
nand U45687 (N_45687,N_40226,N_44404);
xnor U45688 (N_45688,N_41499,N_43942);
or U45689 (N_45689,N_42568,N_40329);
nor U45690 (N_45690,N_41435,N_40290);
or U45691 (N_45691,N_44454,N_42914);
or U45692 (N_45692,N_43967,N_44049);
or U45693 (N_45693,N_44485,N_42744);
xnor U45694 (N_45694,N_40450,N_40022);
nand U45695 (N_45695,N_43945,N_40540);
or U45696 (N_45696,N_41609,N_41858);
and U45697 (N_45697,N_44660,N_40055);
nor U45698 (N_45698,N_41146,N_43823);
nor U45699 (N_45699,N_40509,N_44260);
or U45700 (N_45700,N_41039,N_42747);
xor U45701 (N_45701,N_44654,N_42057);
nand U45702 (N_45702,N_40563,N_41143);
and U45703 (N_45703,N_44279,N_43734);
nor U45704 (N_45704,N_43687,N_44246);
or U45705 (N_45705,N_44234,N_41288);
xor U45706 (N_45706,N_43899,N_40366);
nor U45707 (N_45707,N_42636,N_43308);
and U45708 (N_45708,N_43915,N_41518);
nor U45709 (N_45709,N_41150,N_44953);
nor U45710 (N_45710,N_42493,N_41938);
nor U45711 (N_45711,N_43589,N_43926);
and U45712 (N_45712,N_41981,N_42460);
nand U45713 (N_45713,N_43794,N_41414);
or U45714 (N_45714,N_42820,N_42630);
xor U45715 (N_45715,N_41111,N_44446);
nor U45716 (N_45716,N_41941,N_44979);
and U45717 (N_45717,N_40904,N_42543);
xnor U45718 (N_45718,N_44856,N_41800);
and U45719 (N_45719,N_41216,N_43312);
and U45720 (N_45720,N_44342,N_43777);
or U45721 (N_45721,N_43586,N_44560);
nor U45722 (N_45722,N_44689,N_42520);
and U45723 (N_45723,N_43302,N_40479);
and U45724 (N_45724,N_40148,N_41407);
nand U45725 (N_45725,N_44693,N_42027);
xnor U45726 (N_45726,N_44383,N_43293);
and U45727 (N_45727,N_42250,N_42165);
and U45728 (N_45728,N_40795,N_41694);
nand U45729 (N_45729,N_43335,N_43502);
xnor U45730 (N_45730,N_41968,N_44826);
or U45731 (N_45731,N_44785,N_40527);
nor U45732 (N_45732,N_44874,N_43105);
nand U45733 (N_45733,N_44472,N_42422);
or U45734 (N_45734,N_40320,N_41124);
xnor U45735 (N_45735,N_40885,N_41269);
and U45736 (N_45736,N_44287,N_44070);
nor U45737 (N_45737,N_44898,N_44486);
nor U45738 (N_45738,N_42203,N_44395);
xor U45739 (N_45739,N_43228,N_44959);
nor U45740 (N_45740,N_43046,N_43102);
and U45741 (N_45741,N_42685,N_40611);
or U45742 (N_45742,N_41662,N_41925);
and U45743 (N_45743,N_41392,N_42006);
xor U45744 (N_45744,N_42403,N_41735);
nand U45745 (N_45745,N_43281,N_42710);
xor U45746 (N_45746,N_44172,N_41431);
nand U45747 (N_45747,N_41202,N_41626);
nand U45748 (N_45748,N_42122,N_44622);
xor U45749 (N_45749,N_43761,N_41761);
xor U45750 (N_45750,N_43829,N_43808);
nand U45751 (N_45751,N_41363,N_42400);
nand U45752 (N_45752,N_44202,N_41676);
nor U45753 (N_45753,N_43540,N_42385);
or U45754 (N_45754,N_44206,N_42219);
nor U45755 (N_45755,N_42373,N_42177);
xor U45756 (N_45756,N_40755,N_44180);
nor U45757 (N_45757,N_42247,N_40065);
xnor U45758 (N_45758,N_44947,N_40922);
nor U45759 (N_45759,N_43838,N_42642);
xnor U45760 (N_45760,N_42069,N_44884);
or U45761 (N_45761,N_43807,N_44424);
or U45762 (N_45762,N_42081,N_42449);
xnor U45763 (N_45763,N_40810,N_41754);
or U45764 (N_45764,N_40902,N_41520);
or U45765 (N_45765,N_44051,N_40693);
or U45766 (N_45766,N_42168,N_40773);
nand U45767 (N_45767,N_43404,N_44686);
xor U45768 (N_45768,N_40805,N_43139);
and U45769 (N_45769,N_41830,N_41607);
and U45770 (N_45770,N_44007,N_43940);
nand U45771 (N_45771,N_44200,N_44237);
and U45772 (N_45772,N_40124,N_40308);
nand U45773 (N_45773,N_44606,N_43923);
and U45774 (N_45774,N_44102,N_41862);
or U45775 (N_45775,N_42750,N_44176);
or U45776 (N_45776,N_44396,N_40682);
or U45777 (N_45777,N_43866,N_40899);
and U45778 (N_45778,N_44537,N_40457);
or U45779 (N_45779,N_41542,N_41338);
and U45780 (N_45780,N_42893,N_44181);
or U45781 (N_45781,N_41559,N_43159);
xnor U45782 (N_45782,N_40090,N_43279);
xor U45783 (N_45783,N_42532,N_43660);
xor U45784 (N_45784,N_43072,N_40782);
or U45785 (N_45785,N_40076,N_44936);
and U45786 (N_45786,N_42309,N_44880);
or U45787 (N_45787,N_43519,N_41583);
nand U45788 (N_45788,N_41864,N_41915);
nor U45789 (N_45789,N_43158,N_42466);
nand U45790 (N_45790,N_43590,N_41173);
and U45791 (N_45791,N_43913,N_43031);
or U45792 (N_45792,N_43270,N_43421);
nand U45793 (N_45793,N_40060,N_44000);
xor U45794 (N_45794,N_40905,N_43725);
and U45795 (N_45795,N_40633,N_42210);
xor U45796 (N_45796,N_42799,N_41723);
xnor U45797 (N_45797,N_42151,N_41521);
and U45798 (N_45798,N_44907,N_43300);
nand U45799 (N_45799,N_41043,N_42721);
nor U45800 (N_45800,N_44799,N_44129);
nand U45801 (N_45801,N_43393,N_43081);
xor U45802 (N_45802,N_40251,N_43114);
and U45803 (N_45803,N_42123,N_40002);
xnor U45804 (N_45804,N_42162,N_44576);
or U45805 (N_45805,N_43439,N_41909);
and U45806 (N_45806,N_44935,N_43330);
and U45807 (N_45807,N_40542,N_42166);
or U45808 (N_45808,N_43454,N_41833);
xor U45809 (N_45809,N_42626,N_41930);
nand U45810 (N_45810,N_44639,N_42202);
and U45811 (N_45811,N_40214,N_44110);
and U45812 (N_45812,N_42700,N_43476);
and U45813 (N_45813,N_44632,N_44335);
nor U45814 (N_45814,N_44039,N_41753);
or U45815 (N_45815,N_43155,N_41751);
xnor U45816 (N_45816,N_44577,N_44824);
xnor U45817 (N_45817,N_41233,N_43896);
or U45818 (N_45818,N_44587,N_44315);
or U45819 (N_45819,N_41028,N_43112);
nand U45820 (N_45820,N_44368,N_42912);
nand U45821 (N_45821,N_43177,N_42288);
nor U45822 (N_45822,N_42689,N_43375);
or U45823 (N_45823,N_44328,N_41942);
or U45824 (N_45824,N_44220,N_41367);
xor U45825 (N_45825,N_43073,N_41231);
or U45826 (N_45826,N_44917,N_41244);
and U45827 (N_45827,N_42755,N_41720);
or U45828 (N_45828,N_44950,N_44872);
or U45829 (N_45829,N_40932,N_42178);
xnor U45830 (N_45830,N_42115,N_43036);
and U45831 (N_45831,N_41474,N_41334);
nor U45832 (N_45832,N_43078,N_43283);
or U45833 (N_45833,N_43890,N_42305);
or U45834 (N_45834,N_43331,N_43600);
xor U45835 (N_45835,N_41624,N_40177);
nor U45836 (N_45836,N_41536,N_40621);
and U45837 (N_45837,N_41160,N_40447);
nand U45838 (N_45838,N_42812,N_42116);
and U45839 (N_45839,N_44010,N_40015);
nor U45840 (N_45840,N_40647,N_44565);
nor U45841 (N_45841,N_40764,N_40588);
nand U45842 (N_45842,N_41012,N_42536);
xnor U45843 (N_45843,N_40612,N_40410);
nor U45844 (N_45844,N_40217,N_40137);
nand U45845 (N_45845,N_40614,N_43897);
or U45846 (N_45846,N_42090,N_41794);
and U45847 (N_45847,N_40661,N_44794);
or U45848 (N_45848,N_41729,N_40084);
nand U45849 (N_45849,N_41593,N_40917);
or U45850 (N_45850,N_40168,N_43101);
nor U45851 (N_45851,N_42916,N_42440);
and U45852 (N_45852,N_41883,N_43949);
and U45853 (N_45853,N_42473,N_40413);
xnor U45854 (N_45854,N_42054,N_43536);
nor U45855 (N_45855,N_42371,N_40796);
nand U45856 (N_45856,N_41473,N_43763);
nand U45857 (N_45857,N_40467,N_42126);
xor U45858 (N_45858,N_43265,N_44483);
and U45859 (N_45859,N_44006,N_43146);
nand U45860 (N_45860,N_42364,N_42341);
nor U45861 (N_45861,N_41047,N_42348);
nand U45862 (N_45862,N_40949,N_40403);
nor U45863 (N_45863,N_40164,N_41413);
xor U45864 (N_45864,N_42149,N_40471);
xor U45865 (N_45865,N_44897,N_41940);
or U45866 (N_45866,N_41993,N_44698);
and U45867 (N_45867,N_44758,N_41248);
or U45868 (N_45868,N_41501,N_44744);
nand U45869 (N_45869,N_42405,N_41418);
nand U45870 (N_45870,N_43854,N_43023);
nand U45871 (N_45871,N_40268,N_43415);
and U45872 (N_45872,N_44471,N_44089);
and U45873 (N_45873,N_42692,N_42150);
nor U45874 (N_45874,N_43194,N_43541);
nand U45875 (N_45875,N_44669,N_43766);
and U45876 (N_45876,N_40314,N_43261);
or U45877 (N_45877,N_40427,N_44906);
xnor U45878 (N_45878,N_44792,N_44076);
nor U45879 (N_45879,N_41643,N_41065);
xnor U45880 (N_45880,N_44650,N_44464);
nand U45881 (N_45881,N_40913,N_40849);
or U45882 (N_45882,N_42297,N_43696);
nand U45883 (N_45883,N_43760,N_44818);
xor U45884 (N_45884,N_44509,N_40474);
xnor U45885 (N_45885,N_42109,N_40507);
and U45886 (N_45886,N_43982,N_44781);
xor U45887 (N_45887,N_40150,N_42408);
or U45888 (N_45888,N_44267,N_44097);
nand U45889 (N_45889,N_40840,N_44986);
xor U45890 (N_45890,N_44194,N_43925);
nor U45891 (N_45891,N_44407,N_40630);
or U45892 (N_45892,N_42272,N_44018);
nand U45893 (N_45893,N_44825,N_41345);
nand U45894 (N_45894,N_43702,N_42967);
or U45895 (N_45895,N_44942,N_40119);
xor U45896 (N_45896,N_44293,N_42376);
xnor U45897 (N_45897,N_42949,N_42254);
nor U45898 (N_45898,N_44096,N_44111);
and U45899 (N_45899,N_40709,N_43884);
or U45900 (N_45900,N_41347,N_41860);
or U45901 (N_45901,N_40159,N_44022);
nor U45902 (N_45902,N_43647,N_40216);
or U45903 (N_45903,N_43288,N_41717);
nor U45904 (N_45904,N_44901,N_41477);
or U45905 (N_45905,N_44525,N_43804);
xnor U45906 (N_45906,N_41565,N_42417);
nor U45907 (N_45907,N_41374,N_41024);
xor U45908 (N_45908,N_41073,N_44356);
and U45909 (N_45909,N_43332,N_41995);
and U45910 (N_45910,N_41050,N_44098);
or U45911 (N_45911,N_41846,N_43719);
xnor U45912 (N_45912,N_43247,N_40975);
and U45913 (N_45913,N_44779,N_42999);
and U45914 (N_45914,N_43860,N_42197);
nand U45915 (N_45915,N_43151,N_42066);
or U45916 (N_45916,N_41690,N_40254);
xnor U45917 (N_45917,N_42565,N_43175);
nand U45918 (N_45918,N_43357,N_43723);
and U45919 (N_45919,N_40105,N_41052);
nand U45920 (N_45920,N_43127,N_40719);
nand U45921 (N_45921,N_40543,N_41384);
nand U45922 (N_45922,N_43178,N_41692);
xor U45923 (N_45923,N_41126,N_43428);
xor U45924 (N_45924,N_42079,N_41410);
nor U45925 (N_45925,N_42852,N_43560);
or U45926 (N_45926,N_40976,N_44398);
and U45927 (N_45927,N_41749,N_44732);
and U45928 (N_45928,N_42030,N_43545);
nor U45929 (N_45929,N_44751,N_42730);
and U45930 (N_45930,N_44062,N_42159);
and U45931 (N_45931,N_40859,N_43417);
nand U45932 (N_45932,N_43961,N_42485);
nor U45933 (N_45933,N_41263,N_42982);
nor U45934 (N_45934,N_44771,N_41546);
or U45935 (N_45935,N_44617,N_43612);
or U45936 (N_45936,N_42547,N_44738);
nor U45937 (N_45937,N_42420,N_42953);
and U45938 (N_45938,N_40525,N_40518);
xnor U45939 (N_45939,N_40327,N_40935);
nand U45940 (N_45940,N_40409,N_42638);
or U45941 (N_45941,N_40951,N_41886);
xnor U45942 (N_45942,N_42842,N_42706);
and U45943 (N_45943,N_43321,N_42492);
and U45944 (N_45944,N_42695,N_42022);
and U45945 (N_45945,N_42794,N_40650);
or U45946 (N_45946,N_41983,N_44226);
nand U45947 (N_45947,N_43388,N_42261);
nor U45948 (N_45948,N_41035,N_41008);
nand U45949 (N_45949,N_40515,N_43965);
xnor U45950 (N_45950,N_41017,N_44918);
xor U45951 (N_45951,N_42049,N_40945);
nor U45952 (N_45952,N_43614,N_42154);
or U45953 (N_45953,N_43730,N_40699);
nand U45954 (N_45954,N_43028,N_43834);
nand U45955 (N_45955,N_40958,N_40652);
and U45956 (N_45956,N_41396,N_40336);
and U45957 (N_45957,N_40252,N_41806);
nor U45958 (N_45958,N_42634,N_43336);
xor U45959 (N_45959,N_43093,N_43398);
or U45960 (N_45960,N_41400,N_43264);
nor U45961 (N_45961,N_43867,N_43412);
or U45962 (N_45962,N_42781,N_43709);
nand U45963 (N_45963,N_40096,N_40071);
nor U45964 (N_45964,N_41325,N_40868);
nand U45965 (N_45965,N_42904,N_42504);
nor U45966 (N_45966,N_44951,N_42243);
and U45967 (N_45967,N_44311,N_44011);
nand U45968 (N_45968,N_43113,N_43737);
or U45969 (N_45969,N_44094,N_40816);
nand U45970 (N_45970,N_43895,N_44164);
or U45971 (N_45971,N_43359,N_41669);
and U45972 (N_45972,N_43134,N_43198);
or U45973 (N_45973,N_41693,N_40644);
nor U45974 (N_45974,N_42328,N_44149);
nor U45975 (N_45975,N_43488,N_41321);
nor U45976 (N_45976,N_40691,N_40451);
nor U45977 (N_45977,N_41046,N_41281);
or U45978 (N_45978,N_43234,N_42800);
and U45979 (N_45979,N_43986,N_40713);
nand U45980 (N_45980,N_41129,N_41708);
xor U45981 (N_45981,N_42362,N_42293);
nand U45982 (N_45982,N_41924,N_40839);
xnor U45983 (N_45983,N_43272,N_42614);
nor U45984 (N_45984,N_42160,N_42581);
nand U45985 (N_45985,N_42075,N_42767);
nand U45986 (N_45986,N_42236,N_43514);
nor U45987 (N_45987,N_43431,N_42078);
nand U45988 (N_45988,N_41161,N_40936);
nand U45989 (N_45989,N_40443,N_42596);
nor U45990 (N_45990,N_41164,N_44080);
xor U45991 (N_45991,N_40531,N_40436);
nand U45992 (N_45992,N_44834,N_43315);
nor U45993 (N_45993,N_42612,N_42759);
xnor U45994 (N_45994,N_40654,N_41071);
and U45995 (N_45995,N_44759,N_43525);
and U45996 (N_45996,N_43985,N_42321);
and U45997 (N_45997,N_44716,N_40790);
and U45998 (N_45998,N_41030,N_40231);
nor U45999 (N_45999,N_41297,N_42445);
and U46000 (N_46000,N_42837,N_44858);
or U46001 (N_46001,N_40632,N_42277);
xor U46002 (N_46002,N_40581,N_40528);
nor U46003 (N_46003,N_40944,N_41272);
and U46004 (N_46004,N_43130,N_42968);
and U46005 (N_46005,N_42787,N_43232);
and U46006 (N_46006,N_42980,N_43191);
xnor U46007 (N_46007,N_44245,N_40550);
or U46008 (N_46008,N_43770,N_44447);
nand U46009 (N_46009,N_41677,N_43195);
xnor U46010 (N_46010,N_41511,N_42251);
and U46011 (N_46011,N_41963,N_41427);
or U46012 (N_46012,N_42173,N_42193);
nor U46013 (N_46013,N_40028,N_40005);
xnor U46014 (N_46014,N_43849,N_40289);
nor U46015 (N_46015,N_41854,N_42882);
xor U46016 (N_46016,N_42045,N_42860);
nand U46017 (N_46017,N_42936,N_43817);
xor U46018 (N_46018,N_44262,N_43311);
and U46019 (N_46019,N_43792,N_40193);
nand U46020 (N_46020,N_41090,N_40877);
xor U46021 (N_46021,N_44014,N_40723);
or U46022 (N_46022,N_40412,N_40875);
and U46023 (N_46023,N_42629,N_44112);
xor U46024 (N_46024,N_42071,N_41532);
xnor U46025 (N_46025,N_44806,N_44782);
and U46026 (N_46026,N_40890,N_44697);
or U46027 (N_46027,N_41424,N_40083);
or U46028 (N_46028,N_40938,N_44179);
or U46029 (N_46029,N_40730,N_44811);
or U46030 (N_46030,N_41320,N_44480);
xnor U46031 (N_46031,N_44302,N_42917);
or U46032 (N_46032,N_44847,N_41725);
nor U46033 (N_46033,N_43997,N_40385);
nor U46034 (N_46034,N_41026,N_40733);
and U46035 (N_46035,N_43991,N_42474);
nand U46036 (N_46036,N_44810,N_42583);
xnor U46037 (N_46037,N_41534,N_41314);
and U46038 (N_46038,N_41243,N_42148);
nor U46039 (N_46039,N_44866,N_40321);
nor U46040 (N_46040,N_40687,N_42515);
and U46041 (N_46041,N_40827,N_41526);
or U46042 (N_46042,N_40275,N_41545);
nand U46043 (N_46043,N_44713,N_43627);
and U46044 (N_46044,N_44455,N_42136);
xnor U46045 (N_46045,N_40848,N_43962);
nor U46046 (N_46046,N_44463,N_43874);
nand U46047 (N_46047,N_44036,N_40101);
nand U46048 (N_46048,N_40399,N_43092);
and U46049 (N_46049,N_44117,N_43681);
or U46050 (N_46050,N_42060,N_41326);
or U46051 (N_46051,N_42780,N_41950);
and U46052 (N_46052,N_43571,N_41516);
nand U46053 (N_46053,N_41037,N_41416);
nand U46054 (N_46054,N_44640,N_40807);
nor U46055 (N_46055,N_42017,N_42414);
xor U46056 (N_46056,N_44662,N_43554);
nand U46057 (N_46057,N_41519,N_40847);
xnor U46058 (N_46058,N_42839,N_42042);
and U46059 (N_46059,N_40903,N_43214);
xor U46060 (N_46060,N_42676,N_40234);
and U46061 (N_46061,N_44338,N_41273);
xnor U46062 (N_46062,N_44538,N_44990);
or U46063 (N_46063,N_42194,N_42696);
and U46064 (N_46064,N_44470,N_43859);
or U46065 (N_46065,N_41108,N_42889);
or U46066 (N_46066,N_40626,N_41853);
or U46067 (N_46067,N_42869,N_43811);
xnor U46068 (N_46068,N_43204,N_42944);
xor U46069 (N_46069,N_40240,N_41799);
and U46070 (N_46070,N_42255,N_40317);
nor U46071 (N_46071,N_41388,N_44740);
nand U46072 (N_46072,N_40615,N_42495);
or U46073 (N_46073,N_44926,N_42691);
nand U46074 (N_46074,N_40548,N_44496);
nand U46075 (N_46075,N_42646,N_43129);
nor U46076 (N_46076,N_41712,N_42670);
nor U46077 (N_46077,N_43212,N_42222);
xor U46078 (N_46078,N_43953,N_43268);
nor U46079 (N_46079,N_41165,N_43585);
xor U46080 (N_46080,N_42666,N_42742);
or U46081 (N_46081,N_43504,N_44903);
and U46082 (N_46082,N_42398,N_42487);
nand U46083 (N_46083,N_40568,N_41294);
and U46084 (N_46084,N_44291,N_41117);
nand U46085 (N_46085,N_42709,N_42574);
nor U46086 (N_46086,N_44864,N_42163);
and U46087 (N_46087,N_44631,N_44459);
xor U46088 (N_46088,N_44008,N_42082);
xor U46089 (N_46089,N_44533,N_42720);
nor U46090 (N_46090,N_44655,N_41476);
xnor U46091 (N_46091,N_41934,N_44801);
or U46092 (N_46092,N_44113,N_40573);
or U46093 (N_46093,N_44977,N_40491);
nand U46094 (N_46094,N_42404,N_44135);
xnor U46095 (N_46095,N_40956,N_43056);
xor U46096 (N_46096,N_40369,N_40933);
nand U46097 (N_46097,N_41417,N_42412);
or U46098 (N_46098,N_42942,N_43658);
nand U46099 (N_46099,N_40014,N_40508);
nand U46100 (N_46100,N_42934,N_43154);
nor U46101 (N_46101,N_43220,N_40973);
nor U46102 (N_46102,N_43285,N_42278);
and U46103 (N_46103,N_44722,N_41890);
nor U46104 (N_46104,N_44619,N_41732);
xnor U46105 (N_46105,N_41960,N_44763);
and U46106 (N_46106,N_41897,N_41036);
xnor U46107 (N_46107,N_43435,N_40243);
nor U46108 (N_46108,N_44067,N_41812);
nand U46109 (N_46109,N_40734,N_42534);
nor U46110 (N_46110,N_40605,N_42198);
or U46111 (N_46111,N_43457,N_42015);
xnor U46112 (N_46112,N_42793,N_40504);
and U46113 (N_46113,N_44561,N_40659);
nand U46114 (N_46114,N_44391,N_40704);
nand U46115 (N_46115,N_40030,N_41673);
nand U46116 (N_46116,N_41739,N_42152);
nand U46117 (N_46117,N_40480,N_44527);
nand U46118 (N_46118,N_43215,N_43461);
nand U46119 (N_46119,N_43784,N_44386);
nand U46120 (N_46120,N_42301,N_44093);
xor U46121 (N_46121,N_42377,N_43099);
xnor U46122 (N_46122,N_43729,N_40301);
xnor U46123 (N_46123,N_41745,N_40259);
nor U46124 (N_46124,N_43576,N_44104);
nor U46125 (N_46125,N_44589,N_40672);
nand U46126 (N_46126,N_43122,N_44657);
xnor U46127 (N_46127,N_41246,N_42631);
nand U46128 (N_46128,N_44341,N_40815);
or U46129 (N_46129,N_40623,N_44121);
or U46130 (N_46130,N_44518,N_40781);
and U46131 (N_46131,N_44709,N_40955);
nor U46132 (N_46132,N_42282,N_42164);
or U46133 (N_46133,N_41234,N_44546);
xor U46134 (N_46134,N_43912,N_41975);
nand U46135 (N_46135,N_42083,N_42560);
xnor U46136 (N_46136,N_41523,N_40948);
nand U46137 (N_46137,N_41022,N_42789);
and U46138 (N_46138,N_41716,N_44999);
xor U46139 (N_46139,N_43065,N_44612);
or U46140 (N_46140,N_43675,N_41667);
nand U46141 (N_46141,N_42383,N_40732);
nor U46142 (N_46142,N_40817,N_40407);
nor U46143 (N_46143,N_43382,N_41913);
nor U46144 (N_46144,N_41018,N_43176);
and U46145 (N_46145,N_43698,N_40004);
nor U46146 (N_46146,N_43160,N_42733);
nand U46147 (N_46147,N_42189,N_41130);
or U46148 (N_46148,N_43076,N_41341);
nor U46149 (N_46149,N_42540,N_41340);
nor U46150 (N_46150,N_43619,N_40140);
xnor U46151 (N_46151,N_42130,N_44235);
nand U46152 (N_46152,N_44854,N_40227);
nand U46153 (N_46153,N_42253,N_40405);
nand U46154 (N_46154,N_43875,N_40901);
nor U46155 (N_46155,N_44072,N_43850);
or U46156 (N_46156,N_44272,N_42518);
nor U46157 (N_46157,N_40912,N_41242);
or U46158 (N_46158,N_44846,N_40075);
xnor U46159 (N_46159,N_44938,N_41343);
xnor U46160 (N_46160,N_42186,N_43193);
nor U46161 (N_46161,N_43970,N_44511);
nor U46162 (N_46162,N_43805,N_41464);
xnor U46163 (N_46163,N_43047,N_40603);
xor U46164 (N_46164,N_40072,N_40510);
xnor U46165 (N_46165,N_42204,N_43245);
nand U46166 (N_46166,N_43905,N_44231);
nand U46167 (N_46167,N_44944,N_44987);
xor U46168 (N_46168,N_40052,N_43788);
nand U46169 (N_46169,N_40303,N_41965);
or U46170 (N_46170,N_42675,N_44747);
nor U46171 (N_46171,N_42129,N_41315);
and U46172 (N_46172,N_44330,N_41625);
and U46173 (N_46173,N_41813,N_43744);
or U46174 (N_46174,N_40779,N_40097);
nor U46175 (N_46175,N_43506,N_43511);
and U46176 (N_46176,N_44505,N_40634);
or U46177 (N_46177,N_41672,N_42084);
xor U46178 (N_46178,N_41584,N_40423);
or U46179 (N_46179,N_41184,N_41525);
xor U46180 (N_46180,N_44186,N_43445);
and U46181 (N_46181,N_41599,N_41335);
or U46182 (N_46182,N_40122,N_42727);
nor U46183 (N_46183,N_42761,N_40521);
nor U46184 (N_46184,N_43682,N_42370);
xor U46185 (N_46185,N_41977,N_40044);
or U46186 (N_46186,N_40770,N_41758);
xor U46187 (N_46187,N_44677,N_42214);
or U46188 (N_46188,N_41980,N_41317);
nand U46189 (N_46189,N_43356,N_41554);
xnor U46190 (N_46190,N_42883,N_42028);
and U46191 (N_46191,N_41765,N_41258);
and U46192 (N_46192,N_43503,N_40042);
or U46193 (N_46193,N_41105,N_43163);
or U46194 (N_46194,N_44616,N_40717);
xor U46195 (N_46195,N_40343,N_40541);
or U46196 (N_46196,N_44029,N_40714);
and U46197 (N_46197,N_43344,N_42960);
nand U46198 (N_46198,N_43599,N_42981);
nor U46199 (N_46199,N_42806,N_40151);
nor U46200 (N_46200,N_42478,N_41947);
or U46201 (N_46201,N_42007,N_43448);
xor U46202 (N_46202,N_44343,N_41740);
and U46203 (N_46203,N_44122,N_41256);
xnor U46204 (N_46204,N_43367,N_41175);
nand U46205 (N_46205,N_41811,N_41480);
nand U46206 (N_46206,N_40376,N_40681);
and U46207 (N_46207,N_40677,N_40942);
nor U46208 (N_46208,N_40408,N_42035);
and U46209 (N_46209,N_43508,N_42996);
or U46210 (N_46210,N_42209,N_43732);
or U46211 (N_46211,N_43438,N_42765);
nand U46212 (N_46212,N_41861,N_42798);
or U46213 (N_46213,N_41660,N_43741);
nor U46214 (N_46214,N_43706,N_42418);
or U46215 (N_46215,N_42144,N_42663);
and U46216 (N_46216,N_42484,N_40066);
xor U46217 (N_46217,N_44610,N_41213);
nand U46218 (N_46218,N_40154,N_44441);
and U46219 (N_46219,N_43992,N_41689);
or U46220 (N_46220,N_41377,N_42862);
nor U46221 (N_46221,N_43746,N_43796);
and U46222 (N_46222,N_41472,N_41603);
nor U46223 (N_46223,N_44912,N_44773);
or U46224 (N_46224,N_40559,N_41895);
xor U46225 (N_46225,N_43294,N_42052);
nor U46226 (N_46226,N_40571,N_41547);
xor U46227 (N_46227,N_44479,N_42326);
nor U46228 (N_46228,N_41467,N_41951);
nand U46229 (N_46229,N_42273,N_44333);
nor U46230 (N_46230,N_43303,N_43011);
xnor U46231 (N_46231,N_41491,N_40783);
or U46232 (N_46232,N_43186,N_40034);
xor U46233 (N_46233,N_43411,N_42928);
nor U46234 (N_46234,N_40063,N_40236);
xnor U46235 (N_46235,N_44466,N_43690);
or U46236 (N_46236,N_40141,N_44933);
nor U46237 (N_46237,N_43881,N_40258);
or U46238 (N_46238,N_40786,N_44106);
nor U46239 (N_46239,N_40058,N_44304);
and U46240 (N_46240,N_42119,N_43587);
or U46241 (N_46241,N_41651,N_43845);
nor U46242 (N_46242,N_44651,N_41120);
nand U46243 (N_46243,N_40665,N_41838);
and U46244 (N_46244,N_44075,N_42291);
xnor U46245 (N_46245,N_43495,N_42239);
xor U46246 (N_46246,N_43626,N_42828);
nor U46247 (N_46247,N_43549,N_41078);
xor U46248 (N_46248,N_42649,N_42053);
xor U46249 (N_46249,N_43824,N_42004);
xor U46250 (N_46250,N_41421,N_42956);
or U46251 (N_46251,N_40020,N_42187);
nand U46252 (N_46252,N_41650,N_44737);
or U46253 (N_46253,N_42319,N_41600);
nand U46254 (N_46254,N_41957,N_42590);
nor U46255 (N_46255,N_44707,N_41319);
nand U46256 (N_46256,N_44809,N_44930);
nand U46257 (N_46257,N_43947,N_43671);
and U46258 (N_46258,N_44931,N_42717);
nand U46259 (N_46259,N_41596,N_40558);
nor U46260 (N_46260,N_40888,N_43783);
or U46261 (N_46261,N_40094,N_42266);
xor U46262 (N_46262,N_40538,N_44491);
nor U46263 (N_46263,N_40059,N_40342);
or U46264 (N_46264,N_44435,N_43628);
or U46265 (N_46265,N_41612,N_43855);
nand U46266 (N_46266,N_40785,N_40551);
and U46267 (N_46267,N_43037,N_41101);
nand U46268 (N_46268,N_42141,N_43443);
nor U46269 (N_46269,N_40943,N_41610);
nor U46270 (N_46270,N_40701,N_44899);
nor U46271 (N_46271,N_40291,N_43474);
nand U46272 (N_46272,N_40036,N_43579);
nor U46273 (N_46273,N_40960,N_42238);
and U46274 (N_46274,N_43444,N_40803);
nor U46275 (N_46275,N_40269,N_44400);
nor U46276 (N_46276,N_40165,N_42598);
xnor U46277 (N_46277,N_40757,N_44743);
or U46278 (N_46278,N_42704,N_42033);
nor U46279 (N_46279,N_41804,N_41469);
xnor U46280 (N_46280,N_44402,N_40331);
or U46281 (N_46281,N_43254,N_40718);
nor U46282 (N_46282,N_44875,N_42662);
nand U46283 (N_46283,N_42556,N_40013);
nor U46284 (N_46284,N_43957,N_44925);
xnor U46285 (N_46285,N_41896,N_44955);
and U46286 (N_46286,N_44886,N_40635);
or U46287 (N_46287,N_43623,N_42771);
nand U46288 (N_46288,N_43624,N_44320);
xor U46289 (N_46289,N_44493,N_42973);
xor U46290 (N_46290,N_44703,N_41962);
nor U46291 (N_46291,N_43990,N_44860);
nor U46292 (N_46292,N_43971,N_42396);
or U46293 (N_46293,N_41357,N_44457);
nor U46294 (N_46294,N_41081,N_41303);
and U46295 (N_46295,N_40934,N_44556);
and U46296 (N_46296,N_42245,N_40351);
nand U46297 (N_46297,N_44602,N_44881);
nand U46298 (N_46298,N_40175,N_43263);
nand U46299 (N_46299,N_40744,N_44659);
or U46300 (N_46300,N_42114,N_41902);
and U46301 (N_46301,N_43886,N_44983);
nand U46302 (N_46302,N_43407,N_40740);
xnor U46303 (N_46303,N_42003,N_44015);
nand U46304 (N_46304,N_44210,N_41475);
and U46305 (N_46305,N_40198,N_44609);
nor U46306 (N_46306,N_42686,N_44406);
xor U46307 (N_46307,N_43144,N_43460);
nor U46308 (N_46308,N_42248,N_43593);
and U46309 (N_46309,N_41613,N_44060);
nand U46310 (N_46310,N_43683,N_40692);
and U46311 (N_46311,N_40394,N_41561);
nor U46312 (N_46312,N_43693,N_43710);
nor U46313 (N_46313,N_42441,N_43432);
nor U46314 (N_46314,N_40620,N_42046);
xnor U46315 (N_46315,N_44453,N_40794);
or U46316 (N_46316,N_44350,N_44798);
nor U46317 (N_46317,N_41460,N_40207);
nand U46318 (N_46318,N_42701,N_40965);
or U46319 (N_46319,N_43646,N_43753);
xor U46320 (N_46320,N_41779,N_43631);
xnor U46321 (N_46321,N_43322,N_42384);
nor U46322 (N_46322,N_42633,N_44618);
and U46323 (N_46323,N_41040,N_43253);
nor U46324 (N_46324,N_44037,N_44421);
xnor U46325 (N_46325,N_40919,N_41989);
nand U46326 (N_46326,N_42548,N_40311);
xor U46327 (N_46327,N_44193,N_42586);
and U46328 (N_46328,N_41270,N_41855);
nand U46329 (N_46329,N_40766,N_44271);
nand U46330 (N_46330,N_41021,N_41025);
xor U46331 (N_46331,N_44791,N_41255);
nand U46332 (N_46332,N_44888,N_40834);
or U46333 (N_46333,N_40379,N_40597);
nand U46334 (N_46334,N_44585,N_44492);
nor U46335 (N_46335,N_40492,N_42479);
nand U46336 (N_46336,N_43800,N_44601);
nand U46337 (N_46337,N_40386,N_40690);
or U46338 (N_46338,N_42322,N_41984);
xnor U46339 (N_46339,N_43070,N_43117);
or U46340 (N_46340,N_40438,N_41873);
nand U46341 (N_46341,N_40696,N_44830);
or U46342 (N_46342,N_40769,N_44167);
and U46343 (N_46343,N_42741,N_41567);
or U46344 (N_46344,N_41172,N_43179);
nor U46345 (N_46345,N_44661,N_42310);
or U46346 (N_46346,N_44307,N_42578);
and U46347 (N_46347,N_41495,N_42343);
nand U46348 (N_46348,N_41948,N_41488);
xnor U46349 (N_46349,N_44710,N_43645);
nand U46350 (N_46350,N_42226,N_42564);
nand U46351 (N_46351,N_40962,N_43467);
or U46352 (N_46352,N_40765,N_43622);
xnor U46353 (N_46353,N_41000,N_40276);
nor U46354 (N_46354,N_43128,N_41148);
and U46355 (N_46355,N_43089,N_41481);
xnor U46356 (N_46356,N_41114,N_42094);
nand U46357 (N_46357,N_42514,N_40601);
or U46358 (N_46358,N_41621,N_41045);
nor U46359 (N_46359,N_42323,N_43555);
and U46360 (N_46360,N_41738,N_44541);
xnor U46361 (N_46361,N_41429,N_44627);
xor U46362 (N_46362,N_40762,N_42563);
and U46363 (N_46363,N_43752,N_42462);
or U46364 (N_46364,N_42845,N_43451);
nand U46365 (N_46365,N_40167,N_43440);
or U46366 (N_46366,N_40487,N_44591);
or U46367 (N_46367,N_41251,N_43499);
nor U46368 (N_46368,N_44508,N_43565);
nand U46369 (N_46369,N_42014,N_41444);
nand U46370 (N_46370,N_42517,N_40281);
nor U46371 (N_46371,N_43255,N_43567);
xnor U46372 (N_46372,N_41562,N_42285);
or U46373 (N_46373,N_44019,N_44445);
or U46374 (N_46374,N_43507,N_44159);
and U46375 (N_46375,N_43172,N_42930);
xor U46376 (N_46376,N_42471,N_42707);
nor U46377 (N_46377,N_42329,N_43080);
nor U46378 (N_46378,N_43043,N_44769);
nand U46379 (N_46379,N_42347,N_43133);
nand U46380 (N_46380,N_43665,N_42490);
xor U46381 (N_46381,N_41985,N_43902);
and U46382 (N_46382,N_44574,N_41733);
nand U46383 (N_46383,N_42843,N_41644);
or U46384 (N_46384,N_40367,N_42635);
nor U46385 (N_46385,N_43124,N_41433);
xnor U46386 (N_46386,N_40970,N_44664);
and U46387 (N_46387,N_41076,N_44146);
and U46388 (N_46388,N_40747,N_42156);
nor U46389 (N_46389,N_43390,N_40925);
xor U46390 (N_46390,N_42894,N_41615);
and U46391 (N_46391,N_42426,N_41679);
nand U46392 (N_46392,N_44928,N_42240);
and U46393 (N_46393,N_43425,N_43721);
or U46394 (N_46394,N_41616,N_40356);
or U46395 (N_46395,N_40242,N_44216);
nand U46396 (N_46396,N_43633,N_42673);
or U46397 (N_46397,N_43954,N_43003);
nor U46398 (N_46398,N_43162,N_44910);
xnor U46399 (N_46399,N_40606,N_43828);
xor U46400 (N_46400,N_40536,N_42357);
nand U46401 (N_46401,N_41151,N_43237);
or U46402 (N_46402,N_41500,N_40361);
xor U46403 (N_46403,N_44243,N_42724);
and U46404 (N_46404,N_43015,N_41104);
or U46405 (N_46405,N_41602,N_41135);
nor U46406 (N_46406,N_42772,N_41912);
or U46407 (N_46407,N_42013,N_43104);
nand U46408 (N_46408,N_44965,N_41394);
nand U46409 (N_46409,N_40039,N_42388);
nand U46410 (N_46410,N_44048,N_41893);
or U46411 (N_46411,N_44868,N_41411);
nand U46412 (N_46412,N_44313,N_40174);
nor U46413 (N_46413,N_42436,N_40854);
nand U46414 (N_46414,N_41671,N_41356);
or U46415 (N_46415,N_44017,N_43815);
nor U46416 (N_46416,N_42790,N_43812);
xnor U46417 (N_46417,N_41134,N_42139);
xor U46418 (N_46418,N_44439,N_44941);
and U46419 (N_46419,N_40532,N_42051);
and U46420 (N_46420,N_40739,N_42651);
nor U46421 (N_46421,N_42353,N_41023);
xor U46422 (N_46422,N_41508,N_43147);
or U46423 (N_46423,N_43296,N_42672);
or U46424 (N_46424,N_41966,N_44924);
nor U46425 (N_46425,N_41815,N_44995);
xor U46426 (N_46426,N_40298,N_40664);
and U46427 (N_46427,N_41503,N_43243);
xor U46428 (N_46428,N_41441,N_42925);
or U46429 (N_46429,N_44915,N_41819);
and U46430 (N_46430,N_40637,N_44673);
xor U46431 (N_46431,N_43523,N_42579);
nor U46432 (N_46432,N_40390,N_43171);
nor U46433 (N_46433,N_44040,N_42722);
and U46434 (N_46434,N_42430,N_44783);
nand U46435 (N_46435,N_40135,N_42814);
and U46436 (N_46436,N_42183,N_44286);
or U46437 (N_46437,N_43632,N_44318);
or U46438 (N_46438,N_43552,N_41805);
xnor U46439 (N_46439,N_44175,N_42836);
and U46440 (N_46440,N_41553,N_40232);
nor U46441 (N_46441,N_43423,N_44489);
and U46442 (N_46442,N_44281,N_43520);
and U46443 (N_46443,N_44717,N_41308);
nand U46444 (N_46444,N_43935,N_41286);
or U46445 (N_46445,N_40836,N_41955);
nand U46446 (N_46446,N_44635,N_43699);
nand U46447 (N_46447,N_43493,N_42044);
xnor U46448 (N_46448,N_42235,N_43948);
nor U46449 (N_46449,N_43152,N_44593);
xnor U46450 (N_46450,N_42971,N_44595);
nand U46451 (N_46451,N_43919,N_43248);
nor U46452 (N_46452,N_41498,N_42002);
and U46453 (N_46453,N_40201,N_44182);
and U46454 (N_46454,N_41061,N_42539);
or U46455 (N_46455,N_44822,N_41451);
nand U46456 (N_46456,N_43802,N_42621);
nor U46457 (N_46457,N_42923,N_44084);
xor U46458 (N_46458,N_43700,N_43798);
nor U46459 (N_46459,N_40524,N_42281);
nor U46460 (N_46460,N_43249,N_42167);
nor U46461 (N_46461,N_43189,N_42406);
xnor U46462 (N_46462,N_42486,N_41247);
nand U46463 (N_46463,N_43324,N_42962);
and U46464 (N_46464,N_40340,N_42679);
or U46465 (N_46465,N_44652,N_41318);
xnor U46466 (N_46466,N_40522,N_43271);
nand U46467 (N_46467,N_43900,N_40419);
and U46468 (N_46468,N_42008,N_40884);
nor U46469 (N_46469,N_40624,N_42525);
and U46470 (N_46470,N_40893,N_42927);
xnor U46471 (N_46471,N_42796,N_43365);
or U46472 (N_46472,N_42330,N_40112);
and U46473 (N_46473,N_42259,N_44721);
xor U46474 (N_46474,N_44379,N_43446);
and U46475 (N_46475,N_43166,N_42091);
xnor U46476 (N_46476,N_42714,N_41726);
or U46477 (N_46477,N_41107,N_40722);
nand U46478 (N_46478,N_42855,N_40383);
nand U46479 (N_46479,N_41569,N_41292);
nor U46480 (N_46480,N_43174,N_42902);
xor U46481 (N_46481,N_40220,N_44259);
nor U46482 (N_46482,N_40007,N_44937);
nor U46483 (N_46483,N_43653,N_40831);
nor U46484 (N_46484,N_43380,N_43479);
nor U46485 (N_46485,N_40035,N_44382);
and U46486 (N_46486,N_40771,N_43472);
and U46487 (N_46487,N_44329,N_41011);
nor U46488 (N_46488,N_44520,N_40556);
or U46489 (N_46489,N_44519,N_43749);
nand U46490 (N_46490,N_42571,N_40047);
xor U46491 (N_46491,N_41788,N_41756);
or U46492 (N_46492,N_44598,N_44833);
and U46493 (N_46493,N_44814,N_44580);
nand U46494 (N_46494,N_44647,N_40869);
or U46495 (N_46495,N_43384,N_44068);
nor U46496 (N_46496,N_41153,N_40802);
nand U46497 (N_46497,N_43338,N_42690);
xor U46498 (N_46498,N_43562,N_42318);
or U46499 (N_46499,N_42039,N_43165);
nor U46500 (N_46500,N_40937,N_41768);
nand U46501 (N_46501,N_41141,N_41118);
nor U46502 (N_46502,N_41697,N_42599);
nor U46503 (N_46503,N_44349,N_42989);
nand U46504 (N_46504,N_43054,N_41507);
and U46505 (N_46505,N_41102,N_42641);
xnor U46506 (N_46506,N_40669,N_44016);
or U46507 (N_46507,N_40045,N_44208);
or U46508 (N_46508,N_44828,N_44594);
and U46509 (N_46509,N_42602,N_43216);
xnor U46510 (N_46510,N_41486,N_42225);
and U46511 (N_46511,N_42224,N_40579);
nand U46512 (N_46512,N_43219,N_43364);
xnor U46513 (N_46513,N_42494,N_40284);
and U46514 (N_46514,N_43287,N_42393);
xnor U46515 (N_46515,N_44921,N_41465);
and U46516 (N_46516,N_40950,N_43252);
xor U46517 (N_46517,N_42558,N_44377);
xor U46518 (N_46518,N_41648,N_44812);
or U46519 (N_46519,N_43862,N_41961);
nand U46520 (N_46520,N_40954,N_43754);
and U46521 (N_46521,N_43803,N_44789);
nor U46522 (N_46522,N_44456,N_41589);
or U46523 (N_46523,N_42969,N_42476);
nand U46524 (N_46524,N_42359,N_44562);
nor U46525 (N_46525,N_43487,N_40828);
nor U46526 (N_46526,N_42600,N_43314);
nor U46527 (N_46527,N_41195,N_43304);
nand U46528 (N_46528,N_42509,N_42815);
and U46529 (N_46529,N_40760,N_43458);
nor U46530 (N_46530,N_43993,N_42366);
and U46531 (N_46531,N_41456,N_40529);
nand U46532 (N_46532,N_44688,N_43779);
xor U46533 (N_46533,N_43840,N_41401);
xnor U46534 (N_46534,N_42964,N_44465);
xor U46535 (N_46535,N_41713,N_42063);
and U46536 (N_46536,N_40110,N_43557);
and U46537 (N_46537,N_42671,N_42512);
xnor U46538 (N_46538,N_41550,N_40736);
nand U46539 (N_46539,N_40731,N_43887);
and U46540 (N_46540,N_43148,N_44699);
xor U46541 (N_46541,N_40157,N_40501);
xor U46542 (N_46542,N_42352,N_40018);
or U46543 (N_46543,N_40499,N_42302);
or U46544 (N_46544,N_43573,N_41573);
nor U46545 (N_46545,N_44183,N_42753);
and U46546 (N_46546,N_41455,N_43974);
nand U46547 (N_46547,N_42976,N_41042);
nor U46548 (N_46548,N_43534,N_43012);
and U46549 (N_46549,N_41091,N_40011);
or U46550 (N_46550,N_43836,N_43656);
nor U46551 (N_46551,N_43595,N_42584);
xor U46552 (N_46552,N_44074,N_44207);
and U46553 (N_46553,N_41295,N_40345);
or U46554 (N_46554,N_43269,N_41434);
and U46555 (N_46555,N_43572,N_43256);
and U46556 (N_46556,N_41079,N_41728);
nor U46557 (N_46557,N_41718,N_44516);
xnor U46558 (N_46558,N_44380,N_42822);
and U46559 (N_46559,N_43449,N_42653);
and U46560 (N_46560,N_42108,N_44225);
and U46561 (N_46561,N_44887,N_44649);
or U46562 (N_46562,N_41057,N_43655);
nor U46563 (N_46563,N_42125,N_44620);
and U46564 (N_46564,N_44934,N_42853);
and U46565 (N_46565,N_43885,N_42331);
nand U46566 (N_46566,N_44753,N_40026);
and U46567 (N_46567,N_42174,N_42143);
nor U46568 (N_46568,N_42098,N_40666);
xnor U46569 (N_46569,N_43821,N_44984);
nand U46570 (N_46570,N_41809,N_44241);
xnor U46571 (N_46571,N_42432,N_41766);
and U46572 (N_46572,N_42120,N_44551);
nor U46573 (N_46573,N_43030,N_42913);
and U46574 (N_46574,N_41691,N_44599);
nand U46575 (N_46575,N_41762,N_44498);
xor U46576 (N_46576,N_44085,N_42264);
nand U46577 (N_46577,N_43392,N_43787);
nand U46578 (N_46578,N_42101,N_43879);
nor U46579 (N_46579,N_44373,N_41657);
nor U46580 (N_46580,N_41250,N_44376);
and U46581 (N_46581,N_43355,N_40966);
nor U46582 (N_46582,N_44857,N_44428);
and U46583 (N_46583,N_42859,N_43052);
nor U46584 (N_46584,N_44418,N_43705);
nor U46585 (N_46585,N_42873,N_44679);
xor U46586 (N_46586,N_43087,N_41879);
xnor U46587 (N_46587,N_44410,N_42688);
or U46588 (N_46588,N_41278,N_43868);
nor U46589 (N_46589,N_44169,N_43764);
or U46590 (N_46590,N_43981,N_43769);
and U46591 (N_46591,N_40109,N_43029);
nand U46592 (N_46592,N_40716,N_44691);
xnor U46593 (N_46593,N_41772,N_42195);
and U46594 (N_46594,N_42118,N_43944);
and U46595 (N_46595,N_41899,N_40574);
or U46596 (N_46596,N_40250,N_41002);
or U46597 (N_46597,N_44443,N_40113);
nand U46598 (N_46598,N_40980,N_42941);
xnor U46599 (N_46599,N_41289,N_41911);
and U46600 (N_46600,N_43013,N_41935);
or U46601 (N_46601,N_41640,N_40993);
or U46602 (N_46602,N_40092,N_41632);
and U46603 (N_46603,N_42047,N_44667);
nor U46604 (N_46604,N_44815,N_44658);
xnor U46605 (N_46605,N_43183,N_40265);
xor U46606 (N_46606,N_42454,N_41727);
nand U46607 (N_46607,N_43932,N_41881);
and U46608 (N_46608,N_44902,N_43464);
and U46609 (N_46609,N_44360,N_41843);
and U46610 (N_46610,N_43578,N_44739);
nor U46611 (N_46611,N_43883,N_44861);
nor U46612 (N_46612,N_42728,N_41849);
or U46613 (N_46613,N_40753,N_42627);
or U46614 (N_46614,N_43995,N_42545);
nor U46615 (N_46615,N_43119,N_43864);
or U46616 (N_46616,N_43320,N_42263);
xnor U46617 (N_46617,N_40454,N_41067);
nor U46618 (N_46618,N_42435,N_44448);
or U46619 (N_46619,N_44390,N_43580);
and U46620 (N_46620,N_43362,N_42232);
nor U46621 (N_46621,N_40511,N_43010);
or U46622 (N_46622,N_41581,N_41423);
and U46623 (N_46623,N_43988,N_41544);
and U46624 (N_46624,N_44490,N_43882);
nand U46625 (N_46625,N_40915,N_43429);
nand U46626 (N_46626,N_44438,N_44735);
and U46627 (N_46627,N_41077,N_43786);
and U46628 (N_46628,N_43735,N_44417);
nand U46629 (N_46629,N_41752,N_41618);
xor U46630 (N_46630,N_40456,N_42172);
or U46631 (N_46631,N_44052,N_42217);
and U46632 (N_46632,N_44615,N_44184);
or U46633 (N_46633,N_40483,N_44727);
and U46634 (N_46634,N_42918,N_40322);
and U46635 (N_46635,N_42683,N_41605);
nor U46636 (N_46636,N_42423,N_40078);
nor U46637 (N_46637,N_42608,N_41552);
or U46638 (N_46638,N_43938,N_43826);
xor U46639 (N_46639,N_42102,N_40826);
nor U46640 (N_46640,N_42121,N_40651);
or U46641 (N_46641,N_42391,N_40446);
and U46642 (N_46642,N_40380,N_43931);
xor U46643 (N_46643,N_43389,N_44290);
xnor U46644 (N_46644,N_41086,N_43217);
nand U46645 (N_46645,N_41952,N_41666);
and U46646 (N_46646,N_43278,N_40589);
nor U46647 (N_46647,N_42212,N_43772);
nand U46648 (N_46648,N_40172,N_40750);
nand U46649 (N_46649,N_44278,N_42287);
and U46650 (N_46650,N_44567,N_44545);
nand U46651 (N_46651,N_43397,N_40592);
or U46652 (N_46652,N_43911,N_40516);
nand U46653 (N_46653,N_41653,N_41056);
xnor U46654 (N_46654,N_42117,N_41212);
xor U46655 (N_46655,N_40907,N_40514);
nand U46656 (N_46656,N_42880,N_42113);
nor U46657 (N_46657,N_44588,N_43115);
or U46658 (N_46658,N_44214,N_44473);
nor U46659 (N_46659,N_42296,N_43069);
nor U46660 (N_46660,N_41177,N_41816);
and U46661 (N_46661,N_44962,N_41051);
nor U46662 (N_46662,N_40152,N_40442);
nor U46663 (N_46663,N_42072,N_42324);
nor U46664 (N_46664,N_40353,N_41249);
nand U46665 (N_46665,N_41383,N_41649);
nand U46666 (N_46666,N_41608,N_40208);
nand U46667 (N_46667,N_41958,N_42237);
xnor U46668 (N_46668,N_44842,N_41398);
nor U46669 (N_46669,N_42103,N_42943);
nor U46670 (N_46670,N_40469,N_42110);
xnor U46671 (N_46671,N_40711,N_44319);
or U46672 (N_46672,N_43910,N_42346);
nor U46673 (N_46673,N_41404,N_42879);
nand U46674 (N_46674,N_40488,N_40064);
xor U46675 (N_46675,N_43251,N_41591);
and U46676 (N_46676,N_44303,N_40874);
xor U46677 (N_46677,N_44772,N_44997);
and U46678 (N_46678,N_44385,N_43071);
and U46679 (N_46679,N_40720,N_41038);
or U46680 (N_46680,N_41125,N_41681);
and U46681 (N_46681,N_40478,N_43863);
or U46682 (N_46682,N_42161,N_44432);
and U46683 (N_46683,N_41927,N_41449);
xnor U46684 (N_46684,N_43888,N_44621);
nand U46685 (N_46685,N_40486,N_44761);
nor U46686 (N_46686,N_41298,N_43550);
or U46687 (N_46687,N_44306,N_40545);
nor U46688 (N_46688,N_43452,N_40864);
nand U46689 (N_46689,N_40774,N_43810);
nor U46690 (N_46690,N_44807,N_41267);
or U46691 (N_46691,N_44613,N_42132);
nor U46692 (N_46692,N_42745,N_41918);
xor U46693 (N_46693,N_40158,N_43430);
or U46694 (N_46694,N_42921,N_40248);
xor U46695 (N_46695,N_41324,N_41322);
nor U46696 (N_46696,N_40062,N_43869);
xnor U46697 (N_46697,N_44684,N_43409);
and U46698 (N_46698,N_44927,N_41954);
or U46699 (N_46699,N_43289,N_43939);
or U46700 (N_46700,N_41931,N_43598);
xor U46701 (N_46701,N_41496,N_43759);
nand U46702 (N_46702,N_43434,N_40387);
nor U46703 (N_46703,N_42984,N_40506);
nor U46704 (N_46704,N_41678,N_43943);
xnor U46705 (N_46705,N_40307,N_42887);
xor U46706 (N_46706,N_40466,N_43917);
nor U46707 (N_46707,N_40274,N_41176);
nor U46708 (N_46708,N_40104,N_40639);
nor U46709 (N_46709,N_41168,N_41228);
nand U46710 (N_46710,N_43819,N_43976);
and U46711 (N_46711,N_43695,N_40953);
and U46712 (N_46712,N_40077,N_42776);
or U46713 (N_46713,N_42606,N_44317);
and U46714 (N_46714,N_41306,N_41928);
nand U46715 (N_46715,N_41790,N_40287);
xor U46716 (N_46716,N_44731,N_41328);
nand U46717 (N_46717,N_41533,N_41219);
xor U46718 (N_46718,N_40462,N_40642);
nor U46719 (N_46719,N_41587,N_40625);
nand U46720 (N_46720,N_41235,N_42915);
nand U46721 (N_46721,N_43116,N_41309);
xor U46722 (N_46722,N_40969,N_44130);
nor U46723 (N_46723,N_40277,N_44819);
xnor U46724 (N_46724,N_41490,N_44539);
nor U46725 (N_46725,N_42315,N_43210);
and U46726 (N_46726,N_43433,N_43250);
nand U46727 (N_46727,N_40604,N_40684);
nand U46728 (N_46728,N_43941,N_44512);
or U46729 (N_46729,N_40003,N_42100);
nand U46730 (N_46730,N_43901,N_42601);
and U46731 (N_46731,N_42058,N_40627);
or U46732 (N_46732,N_44996,N_44378);
and U46733 (N_46733,N_42500,N_43348);
or U46734 (N_46734,N_40812,N_42179);
nor U46735 (N_46735,N_42773,N_40346);
and U46736 (N_46736,N_43021,N_42283);
nor U46737 (N_46737,N_44911,N_43401);
xor U46738 (N_46738,N_42888,N_40772);
and U46739 (N_46739,N_40184,N_41342);
or U46740 (N_46740,N_40196,N_43258);
and U46741 (N_46741,N_41696,N_40567);
nor U46742 (N_46742,N_44569,N_41793);
nor U46743 (N_46743,N_40811,N_40100);
nor U46744 (N_46744,N_41282,N_40853);
xnor U46745 (N_46745,N_42271,N_41171);
or U46746 (N_46746,N_42397,N_42095);
nand U46747 (N_46747,N_40851,N_40673);
nand U46748 (N_46748,N_44521,N_42735);
or U46749 (N_46749,N_41659,N_41159);
and U46750 (N_46750,N_41003,N_40829);
nor U46751 (N_46751,N_40871,N_44945);
nor U46752 (N_46752,N_43492,N_44855);
nor U46753 (N_46753,N_43604,N_43712);
nor U46754 (N_46754,N_43610,N_44885);
nor U46755 (N_46755,N_43667,N_40879);
or U46756 (N_46756,N_40523,N_43977);
or U46757 (N_46757,N_41575,N_40742);
xnor U46758 (N_46758,N_40463,N_42811);
nand U46759 (N_46759,N_44852,N_40876);
or U46760 (N_46760,N_42401,N_44045);
and U46761 (N_46761,N_43206,N_41330);
or U46762 (N_46762,N_42693,N_41402);
nor U46763 (N_46763,N_42363,N_40728);
nor U46764 (N_46764,N_42386,N_44900);
or U46765 (N_46765,N_41189,N_41192);
or U46766 (N_46766,N_44991,N_44972);
xor U46767 (N_46767,N_42073,N_43517);
nor U46768 (N_46768,N_44624,N_43242);
and U46769 (N_46769,N_42872,N_42457);
nor U46770 (N_46770,N_43613,N_44137);
or U46771 (N_46771,N_43916,N_42885);
nor U46772 (N_46772,N_43060,N_40743);
xnor U46773 (N_46773,N_41115,N_44354);
nor U46774 (N_46774,N_41227,N_42211);
and U46775 (N_46775,N_43831,N_44578);
or U46776 (N_46776,N_44347,N_40546);
nor U46777 (N_46777,N_43150,N_42459);
nor U46778 (N_46778,N_43535,N_43724);
nand U46779 (N_46779,N_41085,N_41371);
nand U46780 (N_46780,N_44461,N_44558);
nand U46781 (N_46781,N_43045,N_43582);
and U46782 (N_46782,N_41307,N_40660);
nor U46783 (N_46783,N_42433,N_43918);
or U46784 (N_46784,N_41574,N_42439);
nor U46785 (N_46785,N_40703,N_40106);
nand U46786 (N_46786,N_41514,N_44477);
and U46787 (N_46787,N_40900,N_44916);
nor U46788 (N_46788,N_41986,N_44154);
or U46789 (N_46789,N_43224,N_40470);
and U46790 (N_46790,N_42062,N_42995);
nand U46791 (N_46791,N_41531,N_44299);
nand U46792 (N_46792,N_42452,N_42997);
or U46793 (N_46793,N_43463,N_43648);
nor U46794 (N_46794,N_44976,N_44841);
nand U46795 (N_46795,N_42551,N_41207);
and U46796 (N_46796,N_40825,N_40472);
and U46797 (N_46797,N_41349,N_44476);
nor U46798 (N_46798,N_41970,N_42903);
or U46799 (N_46799,N_40230,N_43005);
nand U46800 (N_46800,N_43202,N_43309);
and U46801 (N_46801,N_44745,N_44012);
xnor U46802 (N_46802,N_40566,N_40974);
or U46803 (N_46803,N_43372,N_40149);
nor U46804 (N_46804,N_44994,N_44844);
nand U46805 (N_46805,N_40155,N_44140);
or U46806 (N_46806,N_41479,N_40143);
xnor U46807 (N_46807,N_42088,N_40819);
or U46808 (N_46808,N_41706,N_43200);
nor U46809 (N_46809,N_41337,N_43745);
nor U46810 (N_46810,N_41144,N_43494);
nand U46811 (N_46811,N_44050,N_41901);
or U46812 (N_46812,N_42876,N_43132);
nand U46813 (N_46813,N_41976,N_44108);
or U46814 (N_46814,N_42978,N_43125);
and U46815 (N_46815,N_42170,N_42506);
nand U46816 (N_46816,N_43058,N_43017);
xor U46817 (N_46817,N_40552,N_43641);
xor U46818 (N_46818,N_43574,N_42979);
nand U46819 (N_46819,N_40991,N_40648);
and U46820 (N_46820,N_44064,N_43416);
and U46821 (N_46821,N_40894,N_41190);
and U46822 (N_46822,N_40921,N_40746);
and U46823 (N_46823,N_43489,N_40247);
and U46824 (N_46824,N_44695,N_42216);
nor U46825 (N_46825,N_44028,N_44101);
xnor U46826 (N_46826,N_43669,N_42394);
and U46827 (N_46827,N_41614,N_40983);
nor U46828 (N_46828,N_43110,N_42905);
nand U46829 (N_46829,N_42496,N_42561);
xor U46830 (N_46830,N_43703,N_42104);
xnor U46831 (N_46831,N_42777,N_42169);
or U46832 (N_46832,N_43825,N_44488);
xnor U46833 (N_46833,N_41878,N_44683);
or U46834 (N_46834,N_41010,N_44708);
or U46835 (N_46835,N_41870,N_41944);
nand U46836 (N_46836,N_40978,N_43422);
nand U46837 (N_46837,N_42231,N_40368);
nand U46838 (N_46838,N_43955,N_43684);
xor U46839 (N_46839,N_44510,N_43197);
and U46840 (N_46840,N_44013,N_41715);
and U46841 (N_46841,N_41163,N_41209);
or U46842 (N_46842,N_40404,N_42025);
xor U46843 (N_46843,N_44141,N_41280);
and U46844 (N_46844,N_42554,N_42955);
nand U46845 (N_46845,N_40411,N_42482);
or U46846 (N_46846,N_41432,N_44365);
nand U46847 (N_46847,N_42827,N_43091);
xor U46848 (N_46848,N_40270,N_40916);
nand U46849 (N_46849,N_44240,N_44168);
and U46850 (N_46850,N_41869,N_41095);
and U46851 (N_46851,N_44534,N_41540);
nor U46852 (N_46852,N_43244,N_41784);
nor U46853 (N_46853,N_44375,N_40820);
or U46854 (N_46854,N_41510,N_40200);
or U46855 (N_46855,N_41991,N_44583);
nor U46856 (N_46856,N_44838,N_44131);
nand U46857 (N_46857,N_43731,N_44805);
or U46858 (N_46858,N_42335,N_42870);
and U46859 (N_46859,N_41447,N_42184);
xor U46860 (N_46860,N_40439,N_44042);
and U46861 (N_46861,N_41880,N_41731);
xnor U46862 (N_46862,N_42795,N_44156);
nand U46863 (N_46863,N_44681,N_44366);
xor U46864 (N_46864,N_43025,N_41382);
or U46865 (N_46865,N_43346,N_44515);
and U46866 (N_46866,N_43858,N_40040);
or U46867 (N_46867,N_41064,N_41848);
nor U46868 (N_46868,N_44282,N_43876);
and U46869 (N_46869,N_40889,N_42241);
xor U46870 (N_46870,N_44768,N_43973);
xnor U46871 (N_46871,N_41200,N_44889);
xnor U46872 (N_46872,N_43898,N_40082);
nand U46873 (N_46873,N_41127,N_42067);
xnor U46874 (N_46874,N_44503,N_44362);
nor U46875 (N_46875,N_44668,N_42764);
nand U46876 (N_46876,N_43588,N_43778);
or U46877 (N_46877,N_44142,N_43673);
and U46878 (N_46878,N_44494,N_44774);
nor U46879 (N_46879,N_41112,N_41380);
xnor U46880 (N_46880,N_40898,N_42458);
xor U46881 (N_46881,N_40646,N_44254);
and U46882 (N_46882,N_43650,N_41638);
nand U46883 (N_46883,N_41445,N_43776);
nand U46884 (N_46884,N_42182,N_44869);
xor U46885 (N_46885,N_44680,N_43544);
nor U46886 (N_46886,N_44882,N_41877);
nand U46887 (N_46887,N_42809,N_41557);
xor U46888 (N_46888,N_42470,N_41154);
nor U46889 (N_46889,N_42339,N_43742);
nor U46890 (N_46890,N_43767,N_41988);
nor U46891 (N_46891,N_43266,N_41982);
xnor U46892 (N_46892,N_41186,N_43459);
nand U46893 (N_46893,N_41872,N_42488);
and U46894 (N_46894,N_41582,N_44890);
xnor U46895 (N_46895,N_40801,N_44970);
nor U46896 (N_46896,N_44557,N_42345);
xnor U46897 (N_46897,N_41654,N_41919);
nand U46898 (N_46898,N_40837,N_40093);
xor U46899 (N_46899,N_43813,N_40595);
nor U46900 (N_46900,N_42654,N_42674);
nor U46901 (N_46901,N_40190,N_42911);
nand U46902 (N_46902,N_43297,N_43096);
nor U46903 (N_46903,N_40306,N_40056);
xnor U46904 (N_46904,N_42522,N_41845);
and U46905 (N_46905,N_44230,N_44198);
xor U46906 (N_46906,N_40001,N_43921);
nor U46907 (N_46907,N_42220,N_44765);
or U46908 (N_46908,N_43342,N_41058);
and U46909 (N_46909,N_43007,N_42252);
xnor U46910 (N_46910,N_41987,N_43339);
nand U46911 (N_46911,N_40924,N_40745);
xor U46912 (N_46912,N_42648,N_44528);
xor U46913 (N_46913,N_44409,N_42523);
xnor U46914 (N_46914,N_44353,N_44297);
and U46915 (N_46915,N_44427,N_43755);
and U46916 (N_46916,N_40417,N_44756);
nand U46917 (N_46917,N_44764,N_41274);
or U46918 (N_46918,N_43707,N_44340);
nand U46919 (N_46919,N_44332,N_43597);
nand U46920 (N_46920,N_42274,N_41999);
xnor U46921 (N_46921,N_44371,N_42185);
nor U46922 (N_46922,N_43877,N_41092);
or U46923 (N_46923,N_40057,N_41170);
nand U46924 (N_46924,N_40378,N_42196);
and U46925 (N_46925,N_42810,N_44653);
and U46926 (N_46926,N_42784,N_40594);
or U46927 (N_46927,N_41221,N_41504);
or U46928 (N_46928,N_43528,N_41742);
nor U46929 (N_46929,N_41013,N_42171);
xnor U46930 (N_46930,N_44542,N_42716);
xnor U46931 (N_46931,N_40841,N_44357);
or U46932 (N_46932,N_41842,N_42616);
xnor U46933 (N_46933,N_41027,N_42819);
xor U46934 (N_46934,N_44643,N_40758);
nor U46935 (N_46935,N_41601,N_42668);
xnor U46936 (N_46936,N_41487,N_42029);
and U46937 (N_46937,N_44487,N_40911);
nor U46938 (N_46938,N_42909,N_41494);
and U46939 (N_46939,N_41063,N_42863);
nand U46940 (N_46940,N_41461,N_42221);
and U46941 (N_46941,N_44634,N_44431);
xnor U46942 (N_46942,N_40513,N_43240);
xor U46943 (N_46943,N_43920,N_44549);
or U46944 (N_46944,N_40266,N_42086);
xnor U46945 (N_46945,N_41778,N_44128);
xnor U46946 (N_46946,N_40420,N_42871);
nor U46947 (N_46947,N_42947,N_43100);
xnor U46948 (N_46948,N_41974,N_42854);
or U46949 (N_46949,N_41312,N_44827);
and U46950 (N_46950,N_42074,N_41661);
xor U46951 (N_46951,N_40294,N_42729);
xor U46952 (N_46952,N_42317,N_41121);
nand U46953 (N_46953,N_42840,N_44517);
and U46954 (N_46954,N_42501,N_42824);
and U46955 (N_46955,N_43835,N_42857);
or U46956 (N_46956,N_43211,N_42555);
and U46957 (N_46957,N_40756,N_42499);
xnor U46958 (N_46958,N_40653,N_43402);
nand U46959 (N_46959,N_44676,N_41201);
nand U46960 (N_46960,N_43470,N_42314);
and U46961 (N_46961,N_43584,N_42256);
xnor U46962 (N_46962,N_41588,N_41179);
or U46963 (N_46963,N_40464,N_44939);
nor U46964 (N_46964,N_42192,N_40396);
or U46965 (N_46965,N_40341,N_40959);
or U46966 (N_46966,N_44829,N_42718);
nand U46967 (N_46967,N_43456,N_44185);
or U46968 (N_46968,N_40384,N_44057);
and U46969 (N_46969,N_41505,N_43145);
nor U46970 (N_46970,N_42463,N_42760);
nor U46971 (N_46971,N_41704,N_41631);
nor U46972 (N_46972,N_40012,N_40754);
and U46973 (N_46973,N_44573,N_41329);
nor U46974 (N_46974,N_40455,N_42325);
nor U46975 (N_46975,N_42659,N_40429);
nand U46976 (N_46976,N_42387,N_40229);
nand U46977 (N_46977,N_41370,N_44497);
and U46978 (N_46978,N_40147,N_41543);
nor U46979 (N_46979,N_40452,N_43385);
or U46980 (N_46980,N_42468,N_41530);
xor U46981 (N_46981,N_43870,N_40484);
nor U46982 (N_46982,N_40023,N_44715);
xnor U46983 (N_46983,N_41783,N_43213);
xor U46984 (N_46984,N_44389,N_43592);
nand U46985 (N_46985,N_44138,N_43846);
nand U46986 (N_46986,N_40600,N_42566);
or U46987 (N_46987,N_44401,N_42442);
and U46988 (N_46988,N_40398,N_41083);
or U46989 (N_46989,N_41389,N_41302);
xnor U46990 (N_46990,N_40609,N_42350);
nor U46991 (N_46991,N_41215,N_44960);
nand U46992 (N_46992,N_41687,N_41226);
nor U46993 (N_46993,N_41290,N_43354);
nand U46994 (N_46994,N_40519,N_43568);
nand U46995 (N_46995,N_43635,N_42906);
nand U46996 (N_46996,N_41867,N_42537);
or U46997 (N_46997,N_42000,N_43889);
xor U46998 (N_46998,N_42866,N_43044);
nor U46999 (N_46999,N_40649,N_41333);
or U47000 (N_47000,N_42609,N_41096);
nand U47001 (N_47001,N_40315,N_44248);
or U47002 (N_47002,N_41775,N_41016);
xnor U47003 (N_47003,N_40171,N_40043);
nand U47004 (N_47004,N_42085,N_41773);
or U47005 (N_47005,N_43546,N_41358);
nand U47006 (N_47006,N_41683,N_43405);
xnor U47007 (N_47007,N_44153,N_42059);
or U47008 (N_47008,N_42929,N_41539);
or U47009 (N_47009,N_43323,N_41737);
nor U47010 (N_47010,N_44177,N_44712);
and U47011 (N_47011,N_42552,N_41438);
nand U47012 (N_47012,N_44063,N_41906);
nand U47013 (N_47013,N_41452,N_44339);
and U47014 (N_47014,N_41741,N_41964);
and U47015 (N_47015,N_44750,N_44228);
nor U47016 (N_47016,N_40089,N_40091);
and U47017 (N_47017,N_44009,N_40775);
and U47018 (N_47018,N_41857,N_41365);
or U47019 (N_47019,N_40418,N_44114);
xor U47020 (N_47020,N_44596,N_40908);
nor U47021 (N_47021,N_44462,N_43347);
and U47022 (N_47022,N_44256,N_40272);
xnor U47023 (N_47023,N_42147,N_41116);
nand U47024 (N_47024,N_43924,N_42783);
nor U47025 (N_47025,N_44163,N_42681);
nand U47026 (N_47026,N_42190,N_40170);
xnor U47027 (N_47027,N_43396,N_40882);
nor U47028 (N_47028,N_40402,N_41888);
and U47029 (N_47029,N_44034,N_43768);
or U47030 (N_47030,N_40099,N_43274);
and U47031 (N_47031,N_43762,N_44671);
nor U47032 (N_47032,N_43316,N_40428);
or U47033 (N_47033,N_41641,N_42475);
or U47034 (N_47034,N_41973,N_44020);
nand U47035 (N_47035,N_40435,N_42368);
nor U47036 (N_47036,N_43688,N_41136);
and U47037 (N_47037,N_44352,N_42544);
and U47038 (N_47038,N_42402,N_42258);
xor U47039 (N_47039,N_41323,N_43485);
nand U47040 (N_47040,N_40285,N_41236);
nand U47041 (N_47041,N_42884,N_43959);
nand U47042 (N_47042,N_44274,N_41956);
nand U47043 (N_47043,N_40844,N_43376);
or U47044 (N_47044,N_40800,N_40118);
nand U47045 (N_47045,N_41211,N_44803);
xor U47046 (N_47046,N_40444,N_42736);
nand U47047 (N_47047,N_43602,N_41082);
or U47048 (N_47048,N_40892,N_44786);
or U47049 (N_47049,N_41167,N_41916);
nand U47050 (N_47050,N_40752,N_41084);
nand U47051 (N_47051,N_43426,N_41489);
and U47052 (N_47052,N_40209,N_43551);
or U47053 (N_47053,N_42858,N_41229);
nor U47054 (N_47054,N_43136,N_43842);
xor U47055 (N_47055,N_40582,N_40477);
nor U47056 (N_47056,N_42694,N_44968);
nor U47057 (N_47057,N_40425,N_42413);
and U47058 (N_47058,N_40992,N_41208);
nor U47059 (N_47059,N_41336,N_44197);
xnor U47060 (N_47060,N_44784,N_44726);
nor U47061 (N_47061,N_43689,N_43922);
nand U47062 (N_47062,N_44813,N_44540);
nand U47063 (N_47063,N_44548,N_44157);
and U47064 (N_47064,N_40845,N_44550);
or U47065 (N_47065,N_43505,N_40000);
or U47066 (N_47066,N_40210,N_40533);
nor U47067 (N_47067,N_41814,N_40010);
xor U47068 (N_47068,N_40628,N_43498);
or U47069 (N_47069,N_41395,N_40145);
xnor U47070 (N_47070,N_44061,N_41033);
and U47071 (N_47071,N_40613,N_44088);
and U47072 (N_47072,N_41019,N_40237);
and U47073 (N_47073,N_42680,N_42105);
nor U47074 (N_47074,N_42276,N_43205);
xor U47075 (N_47075,N_40176,N_41132);
nor U47076 (N_47076,N_42816,N_40037);
or U47077 (N_47077,N_44358,N_43615);
and U47078 (N_47078,N_41844,N_40461);
xor U47079 (N_47079,N_43374,N_40139);
and U47080 (N_47080,N_43108,N_44195);
nor U47081 (N_47081,N_44702,N_42465);
nor U47082 (N_47082,N_41635,N_40333);
and U47083 (N_47083,N_43581,N_44233);
or U47084 (N_47084,N_44145,N_43310);
xnor U47085 (N_47085,N_41787,N_41080);
or U47086 (N_47086,N_43880,N_40332);
xnor U47087 (N_47087,N_44092,N_41210);
nor U47088 (N_47088,N_40374,N_43601);
nor U47089 (N_47089,N_44775,N_42878);
nand U47090 (N_47090,N_42381,N_41145);
xor U47091 (N_47091,N_41722,N_40391);
nand U47092 (N_47092,N_41577,N_43751);
nand U47093 (N_47093,N_42805,N_42778);
or U47094 (N_47094,N_44711,N_41293);
nand U47095 (N_47095,N_41198,N_44253);
nand U47096 (N_47096,N_43968,N_42711);
xor U47097 (N_47097,N_41331,N_40494);
nand U47098 (N_47098,N_43496,N_44213);
and U47099 (N_47099,N_43666,N_41458);
nor U47100 (N_47100,N_44656,N_44327);
xor U47101 (N_47101,N_43103,N_42234);
or U47102 (N_47102,N_40098,N_42332);
and U47103 (N_47103,N_42128,N_44817);
nand U47104 (N_47104,N_41188,N_43259);
xor U47105 (N_47105,N_43720,N_44038);
nand U47106 (N_47106,N_40990,N_42922);
or U47107 (N_47107,N_41075,N_43082);
nor U47108 (N_47108,N_44862,N_42576);
nor U47109 (N_47109,N_42803,N_40458);
or U47110 (N_47110,N_43530,N_42992);
nand U47111 (N_47111,N_42447,N_42242);
xnor U47112 (N_47112,N_42483,N_44723);
xor U47113 (N_47113,N_43062,N_41224);
nand U47114 (N_47114,N_42580,N_40212);
nor U47115 (N_47115,N_44285,N_40352);
nor U47116 (N_47116,N_41140,N_40549);
nand U47117 (N_47117,N_40909,N_44865);
nor U47118 (N_47118,N_40050,N_44724);
and U47119 (N_47119,N_43340,N_40260);
nor U47120 (N_47120,N_44526,N_41796);
and U47121 (N_47121,N_44300,N_40636);
and U47122 (N_47122,N_43273,N_42931);
or U47123 (N_47123,N_43820,N_42958);
nor U47124 (N_47124,N_40631,N_42298);
nand U47125 (N_47125,N_44399,N_44514);
nand U47126 (N_47126,N_41744,N_44275);
or U47127 (N_47127,N_43934,N_41181);
xnor U47128 (N_47128,N_44705,N_40183);
and U47129 (N_47129,N_41747,N_42306);
nor U47130 (N_47130,N_43482,N_41996);
nand U47131 (N_47131,N_41825,N_42249);
or U47132 (N_47132,N_41009,N_42340);
xor U47133 (N_47133,N_42438,N_44787);
or U47134 (N_47134,N_40199,N_41419);
nor U47135 (N_47135,N_44777,N_43789);
xnor U47136 (N_47136,N_40297,N_44543);
or U47137 (N_47137,N_43169,N_41818);
and U47138 (N_47138,N_43851,N_44035);
and U47139 (N_47139,N_44637,N_40578);
and U47140 (N_47140,N_44804,N_43328);
nor U47141 (N_47141,N_41757,N_43936);
nor U47142 (N_47142,N_40927,N_44836);
nand U47143 (N_47143,N_43370,N_40465);
xor U47144 (N_47144,N_41859,N_40219);
nor U47145 (N_47145,N_41967,N_42832);
nor U47146 (N_47146,N_44369,N_43118);
or U47147 (N_47147,N_42731,N_41905);
xor U47148 (N_47148,N_40264,N_41702);
and U47149 (N_47149,N_43209,N_42791);
nor U47150 (N_47150,N_43366,N_44136);
or U47151 (N_47151,N_41646,N_41874);
nor U47152 (N_47152,N_44205,N_42443);
and U47153 (N_47153,N_44203,N_43553);
nor U47154 (N_47154,N_44367,N_43006);
nor U47155 (N_47155,N_44642,N_42541);
xor U47156 (N_47156,N_44433,N_41695);
nor U47157 (N_47157,N_40126,N_42577);
or U47158 (N_47158,N_42907,N_40985);
nand U47159 (N_47159,N_40737,N_42570);
xor U47160 (N_47160,N_42320,N_43609);
nor U47161 (N_47161,N_42467,N_43692);
xnor U47162 (N_47162,N_40972,N_44626);
nand U47163 (N_47163,N_44054,N_44840);
nand U47164 (N_47164,N_43188,N_43350);
nor U47165 (N_47165,N_41006,N_42519);
nand U47166 (N_47166,N_41665,N_40569);
and U47167 (N_47167,N_41763,N_42361);
nand U47168 (N_47168,N_40778,N_43035);
nand U47169 (N_47169,N_44215,N_40870);
and U47170 (N_47170,N_43207,N_41776);
nand U47171 (N_47171,N_42280,N_41839);
nor U47172 (N_47172,N_42153,N_42752);
nand U47173 (N_47173,N_40460,N_44998);
xnor U47174 (N_47174,N_40822,N_41939);
nand U47175 (N_47175,N_44337,N_44992);
and U47176 (N_47176,N_42661,N_40555);
nand U47177 (N_47177,N_40422,N_41070);
and U47178 (N_47178,N_43844,N_44026);
nor U47179 (N_47179,N_40038,N_42732);
and U47180 (N_47180,N_41755,N_44071);
nor U47181 (N_47181,N_44973,N_40316);
xor U47182 (N_47182,N_44760,N_44757);
or U47183 (N_47183,N_42748,N_40114);
xnor U47184 (N_47184,N_42831,N_40218);
and U47185 (N_47185,N_40539,N_41579);
nor U47186 (N_47186,N_40835,N_41007);
xor U47187 (N_47187,N_42286,N_43790);
nor U47188 (N_47188,N_41276,N_41943);
or U47189 (N_47189,N_41332,N_41875);
nand U47190 (N_47190,N_42762,N_43774);
nand U47191 (N_47191,N_43621,N_44125);
nand U47192 (N_47192,N_40856,N_42001);
xor U47193 (N_47193,N_41072,N_44586);
or U47194 (N_47194,N_40562,N_40726);
or U47195 (N_47195,N_42749,N_41810);
xor U47196 (N_47196,N_40575,N_44429);
and U47197 (N_47197,N_40645,N_44132);
or U47198 (N_47198,N_42624,N_41239);
xnor U47199 (N_47199,N_40554,N_42823);
xnor U47200 (N_47200,N_41362,N_40414);
or U47201 (N_47201,N_42392,N_43861);
and U47202 (N_47202,N_40591,N_41604);
and U47203 (N_47203,N_42016,N_41353);
or U47204 (N_47204,N_40406,N_40325);
nand U47205 (N_47205,N_43547,N_40348);
xnor U47206 (N_47206,N_41630,N_42593);
or U47207 (N_47207,N_42464,N_41305);
or U47208 (N_47208,N_41868,N_40751);
xnor U47209 (N_47209,N_44894,N_42952);
and U47210 (N_47210,N_42527,N_43480);
nor U47211 (N_47211,N_40655,N_44797);
nor U47212 (N_47212,N_40178,N_41711);
and U47213 (N_47213,N_42379,N_44397);
and U47214 (N_47214,N_42908,N_43512);
or U47215 (N_47215,N_41193,N_41252);
or U47216 (N_47216,N_40006,N_43481);
or U47217 (N_47217,N_44641,N_41253);
xor U47218 (N_47218,N_40963,N_42451);
xor U47219 (N_47219,N_40437,N_40021);
nor U47220 (N_47220,N_40373,N_40761);
or U47221 (N_47221,N_40560,N_42726);
or U47222 (N_47222,N_44555,N_42399);
nand U47223 (N_47223,N_44232,N_44351);
nand U47224 (N_47224,N_43775,N_43837);
and U47225 (N_47225,N_41054,N_41415);
nor U47226 (N_47226,N_43135,N_40282);
or U47227 (N_47227,N_42572,N_44678);
nor U47228 (N_47228,N_41366,N_40166);
or U47229 (N_47229,N_43414,N_40235);
nor U47230 (N_47230,N_41904,N_40392);
nand U47231 (N_47231,N_41682,N_43878);
and U47232 (N_47232,N_42158,N_44044);
or U47233 (N_47233,N_41099,N_40530);
or U47234 (N_47234,N_40749,N_41764);
nor U47235 (N_47235,N_40129,N_40587);
nor U47236 (N_47236,N_41238,N_43740);
nor U47237 (N_47237,N_41528,N_42020);
nor U47238 (N_47238,N_41585,N_40033);
or U47239 (N_47239,N_44795,N_40131);
nor U47240 (N_47240,N_43137,N_43491);
nor U47241 (N_47241,N_40725,N_41443);
nor U47242 (N_47242,N_44265,N_42644);
xnor U47243 (N_47243,N_42846,N_44755);
xor U47244 (N_47244,N_43972,N_40706);
nor U47245 (N_47245,N_43577,N_44322);
and U47246 (N_47246,N_42180,N_42097);
nand U47247 (N_47247,N_40121,N_41138);
or U47248 (N_47248,N_42205,N_41506);
nor U47249 (N_47249,N_41156,N_42407);
or U47250 (N_47250,N_40273,N_44173);
and U47251 (N_47251,N_42358,N_40382);
and U47252 (N_47252,N_43743,N_44147);
and U47253 (N_47253,N_41180,N_44949);
xor U47254 (N_47254,N_40312,N_42588);
and U47255 (N_47255,N_44644,N_44749);
or U47256 (N_47256,N_41364,N_40941);
nor U47257 (N_47257,N_40629,N_43019);
or U47258 (N_47258,N_43872,N_41360);
or U47259 (N_47259,N_40878,N_43685);
xnor U47260 (N_47260,N_43400,N_40241);
nand U47261 (N_47261,N_42697,N_41524);
and U47262 (N_47262,N_42134,N_43441);
xnor U47263 (N_47263,N_43664,N_43387);
xor U47264 (N_47264,N_42026,N_44412);
and U47265 (N_47265,N_40016,N_44674);
and U47266 (N_47266,N_42850,N_41914);
and U47267 (N_47267,N_42019,N_44033);
and U47268 (N_47268,N_40448,N_43522);
and U47269 (N_47269,N_44264,N_44980);
nor U47270 (N_47270,N_42607,N_40288);
and U47271 (N_47271,N_44165,N_42351);
or U47272 (N_47272,N_40897,N_44523);
nor U47273 (N_47273,N_41639,N_40041);
or U47274 (N_47274,N_41537,N_41296);
and U47275 (N_47275,N_43603,N_44370);
nor U47276 (N_47276,N_40997,N_42769);
nand U47277 (N_47277,N_41147,N_43067);
nor U47278 (N_47278,N_41642,N_43780);
nor U47279 (N_47279,N_44288,N_40989);
nand U47280 (N_47280,N_42530,N_43286);
or U47281 (N_47281,N_44956,N_43014);
nand U47282 (N_47282,N_41797,N_42155);
nand U47283 (N_47283,N_44170,N_43325);
or U47284 (N_47284,N_43527,N_43123);
or U47285 (N_47285,N_41436,N_40319);
or U47286 (N_47286,N_42041,N_42024);
or U47287 (N_47287,N_44374,N_42333);
or U47288 (N_47288,N_41287,N_44224);
nand U47289 (N_47289,N_41920,N_40102);
or U47290 (N_47290,N_43059,N_40931);
nand U47291 (N_47291,N_42300,N_44963);
or U47292 (N_47292,N_43377,N_42140);
or U47293 (N_47293,N_41185,N_43403);
and U47294 (N_47294,N_42961,N_43979);
and U47295 (N_47295,N_41428,N_42603);
or U47296 (N_47296,N_40132,N_41892);
xnor U47297 (N_47297,N_41372,N_44974);
nand U47298 (N_47298,N_40547,N_40125);
nand U47299 (N_47299,N_44323,N_42453);
and U47300 (N_47300,N_40564,N_41014);
nor U47301 (N_47301,N_42910,N_40599);
and U47302 (N_47302,N_43616,N_43305);
and U47303 (N_47303,N_44687,N_40335);
and U47304 (N_47304,N_40395,N_42756);
nand U47305 (N_47305,N_40160,N_41834);
or U47306 (N_47306,N_42145,N_42868);
and U47307 (N_47307,N_42597,N_42511);
nand U47308 (N_47308,N_42549,N_43533);
xnor U47309 (N_47309,N_43337,N_41889);
and U47310 (N_47310,N_43203,N_43975);
nand U47311 (N_47311,N_41675,N_44384);
nand U47312 (N_47312,N_43378,N_43903);
nor U47313 (N_47313,N_41178,N_40415);
nand U47314 (N_47314,N_42191,N_43678);
or U47315 (N_47315,N_42344,N_42012);
nand U47316 (N_47316,N_43629,N_44845);
nor U47317 (N_47317,N_43149,N_44920);
nor U47318 (N_47318,N_44426,N_40133);
xor U47319 (N_47319,N_42437,N_42131);
or U47320 (N_47320,N_44663,N_41354);
nor U47321 (N_47321,N_42699,N_41457);
nand U47322 (N_47322,N_42983,N_40194);
nor U47323 (N_47323,N_40534,N_44648);
nor U47324 (N_47324,N_40680,N_42146);
xnor U47325 (N_47325,N_41734,N_44116);
nand U47326 (N_47326,N_40255,N_44729);
nand U47327 (N_47327,N_42946,N_40238);
or U47328 (N_47328,N_42768,N_44266);
and U47329 (N_47329,N_40498,N_40032);
and U47330 (N_47330,N_40490,N_42592);
nor U47331 (N_47331,N_41627,N_43051);
nor U47332 (N_47332,N_44734,N_41921);
xor U47333 (N_47333,N_42604,N_41266);
xor U47334 (N_47334,N_43793,N_44481);
nor U47335 (N_47335,N_43436,N_40095);
or U47336 (N_47336,N_41409,N_43275);
nand U47337 (N_47337,N_44733,N_41182);
and U47338 (N_47338,N_43075,N_43747);
nand U47339 (N_47339,N_44308,N_41275);
nor U47340 (N_47340,N_43785,N_41623);
and U47341 (N_47341,N_43173,N_43018);
nor U47342 (N_47342,N_43351,N_43371);
and U47343 (N_47343,N_44706,N_40067);
nand U47344 (N_47344,N_40863,N_41206);
or U47345 (N_47345,N_44258,N_43852);
xor U47346 (N_47346,N_43620,N_40860);
nand U47347 (N_47347,N_44056,N_42538);
or U47348 (N_47348,N_44150,N_41359);
nor U47349 (N_47349,N_40685,N_41917);
nor U47350 (N_47350,N_40305,N_41406);
nor U47351 (N_47351,N_44513,N_42374);
xnor U47352 (N_47352,N_43718,N_44420);
or U47353 (N_47353,N_42428,N_43246);
nand U47354 (N_47354,N_42480,N_43951);
xor U47355 (N_47355,N_43345,N_44425);
or U47356 (N_47356,N_44849,N_43004);
nor U47357 (N_47357,N_41990,N_40671);
or U47358 (N_47358,N_43049,N_41313);
or U47359 (N_47359,N_44566,N_41497);
xor U47360 (N_47360,N_40430,N_41674);
nand U47361 (N_47361,N_42010,N_40715);
nand U47362 (N_47362,N_42802,N_44024);
xor U47363 (N_47363,N_42477,N_43208);
or U47364 (N_47364,N_43161,N_42450);
nand U47365 (N_47365,N_43156,N_44504);
or U47366 (N_47366,N_41791,N_40818);
nor U47367 (N_47367,N_40689,N_40053);
or U47368 (N_47368,N_40433,N_40182);
xor U47369 (N_47369,N_42064,N_43833);
or U47370 (N_47370,N_43307,N_43419);
nor U47371 (N_47371,N_44422,N_40896);
and U47372 (N_47372,N_42313,N_40707);
xnor U47373 (N_47373,N_41453,N_40858);
nor U47374 (N_47374,N_44211,N_41634);
nand U47375 (N_47375,N_40596,N_44623);
or U47376 (N_47376,N_40123,N_41698);
xnor U47377 (N_47377,N_41066,N_41350);
xor U47378 (N_47378,N_43319,N_41048);
and U47379 (N_47379,N_42526,N_40957);
nor U47380 (N_47380,N_44788,N_41459);
xnor U47381 (N_47381,N_41492,N_42562);
xor U47382 (N_47382,N_41271,N_42737);
or U47383 (N_47383,N_42774,N_44628);
nand U47384 (N_47384,N_40813,N_41405);
nor U47385 (N_47385,N_43532,N_42620);
or U47386 (N_47386,N_40674,N_43038);
nand U47387 (N_47387,N_43654,N_40729);
xnor U47388 (N_47388,N_43282,N_44675);
nand U47389 (N_47389,N_41241,N_42327);
nand U47390 (N_47390,N_40952,N_43040);
nor U47391 (N_47391,N_43856,N_40981);
xor U47392 (N_47392,N_44043,N_43607);
or U47393 (N_47393,N_40162,N_43822);
nand U47394 (N_47394,N_42650,N_44023);
nor U47395 (N_47395,N_40842,N_43733);
or U47396 (N_47396,N_41714,N_40928);
or U47397 (N_47397,N_44364,N_42395);
and U47398 (N_47398,N_40138,N_40688);
and U47399 (N_47399,N_43181,N_43326);
nor U47400 (N_47400,N_41592,N_44989);
and U47401 (N_47401,N_40009,N_41284);
xnor U47402 (N_47402,N_44047,N_41232);
xnor U47403 (N_47403,N_42875,N_40526);
or U47404 (N_47404,N_42763,N_44867);
nand U47405 (N_47405,N_41611,N_44160);
nand U47406 (N_47406,N_43606,N_40204);
xnor U47407 (N_47407,N_42920,N_44078);
and U47408 (N_47408,N_42669,N_40622);
xnor U47409 (N_47409,N_41385,N_43083);
or U47410 (N_47410,N_41840,N_44625);
and U47411 (N_47411,N_41850,N_43726);
nand U47412 (N_47412,N_40700,N_44118);
nor U47413 (N_47413,N_43521,N_41832);
xnor U47414 (N_47414,N_40381,N_41972);
and U47415 (N_47415,N_43639,N_44863);
xor U47416 (N_47416,N_42107,N_41420);
and U47417 (N_47417,N_42825,N_40181);
xnor U47418 (N_47418,N_41556,N_41808);
xnor U47419 (N_47419,N_42751,N_43998);
or U47420 (N_47420,N_42070,N_44099);
xnor U47421 (N_47421,N_43853,N_41580);
nor U47422 (N_47422,N_41598,N_43736);
and U47423 (N_47423,N_44046,N_42684);
xor U47424 (N_47424,N_42877,N_44314);
or U47425 (N_47425,N_41260,N_41450);
and U47426 (N_47426,N_42207,N_40880);
xor U47427 (N_47427,N_41570,N_40068);
xor U47428 (N_47428,N_42111,N_42655);
nand U47429 (N_47429,N_42951,N_44069);
nor U47430 (N_47430,N_43566,N_41558);
and U47431 (N_47431,N_44109,N_40334);
nand U47432 (N_47432,N_40253,N_44161);
xnor U47433 (N_47433,N_42975,N_44499);
or U47434 (N_47434,N_42945,N_40861);
nor U47435 (N_47435,N_42021,N_40833);
or U47436 (N_47436,N_43386,N_43676);
nor U47437 (N_47437,N_43079,N_40061);
nor U47438 (N_47438,N_43418,N_41517);
nand U47439 (N_47439,N_43847,N_42279);
nor U47440 (N_47440,N_44411,N_44475);
nor U47441 (N_47441,N_40705,N_41055);
and U47442 (N_47442,N_42865,N_42424);
or U47443 (N_47443,N_42708,N_44053);
xnor U47444 (N_47444,N_44458,N_41798);
xor U47445 (N_47445,N_42076,N_42489);
nand U47446 (N_47446,N_44728,N_40459);
or U47447 (N_47447,N_44449,N_44419);
nand U47448 (N_47448,N_42446,N_40535);
or U47449 (N_47449,N_40051,N_42498);
and U47450 (N_47450,N_44524,N_41351);
xor U47451 (N_47451,N_42138,N_43230);
nor U47452 (N_47452,N_44988,N_41237);
or U47453 (N_47453,N_44430,N_40712);
and U47454 (N_47454,N_42056,N_43088);
and U47455 (N_47455,N_44767,N_44289);
and U47456 (N_47456,N_44143,N_41217);
nand U47457 (N_47457,N_43704,N_44544);
and U47458 (N_47458,N_44166,N_40940);
nand U47459 (N_47459,N_43306,N_41060);
nand U47460 (N_47460,N_42617,N_43437);
nand U47461 (N_47461,N_40440,N_42938);
nand U47462 (N_47462,N_41139,N_41001);
xor U47463 (N_47463,N_43381,N_41088);
nor U47464 (N_47464,N_40350,N_41636);
and U47465 (N_47465,N_41034,N_40144);
and U47466 (N_47466,N_44059,N_40189);
or U47467 (N_47467,N_44969,N_40824);
and U47468 (N_47468,N_44209,N_44405);
nor U47469 (N_47469,N_41152,N_44600);
nand U47470 (N_47470,N_40947,N_41997);
xnor U47471 (N_47471,N_43649,N_42409);
nor U47472 (N_47472,N_44507,N_43914);
and U47473 (N_47473,N_41538,N_44055);
nand U47474 (N_47474,N_44967,N_42077);
or U47475 (N_47475,N_40355,N_43033);
xnor U47476 (N_47476,N_43291,N_40388);
xnor U47477 (N_47477,N_43694,N_40188);
nor U47478 (N_47478,N_43651,N_44943);
and U47479 (N_47479,N_44348,N_40580);
or U47480 (N_47480,N_44284,N_40323);
or U47481 (N_47481,N_41535,N_42677);
nor U47482 (N_47482,N_41379,N_43946);
xnor U47483 (N_47483,N_40694,N_41162);
or U47484 (N_47484,N_41074,N_40679);
nand U47485 (N_47485,N_43329,N_41563);
nor U47486 (N_47486,N_42284,N_41629);
and U47487 (N_47487,N_40748,N_41750);
xnor U47488 (N_47488,N_40544,N_42595);
nor U47489 (N_47489,N_40806,N_41730);
xnor U47490 (N_47490,N_43055,N_44171);
nand U47491 (N_47491,N_42295,N_42038);
xnor U47492 (N_47492,N_41686,N_43373);
or U47493 (N_47493,N_40476,N_41387);
or U47494 (N_47494,N_43121,N_43983);
nor U47495 (N_47495,N_42427,N_44041);
nor U47496 (N_47496,N_42369,N_40304);
and U47497 (N_47497,N_43526,N_43468);
xor U47498 (N_47498,N_41801,N_44450);
nand U47499 (N_47499,N_43538,N_40245);
and U47500 (N_47500,N_41700,N_40755);
nor U47501 (N_47501,N_41590,N_41925);
xor U47502 (N_47502,N_43773,N_40942);
and U47503 (N_47503,N_41399,N_43598);
nor U47504 (N_47504,N_42326,N_40738);
and U47505 (N_47505,N_43746,N_44816);
or U47506 (N_47506,N_41515,N_44698);
nand U47507 (N_47507,N_43324,N_42041);
nand U47508 (N_47508,N_40179,N_40240);
or U47509 (N_47509,N_42110,N_41553);
nor U47510 (N_47510,N_42846,N_42315);
and U47511 (N_47511,N_40561,N_44801);
nor U47512 (N_47512,N_40590,N_44169);
or U47513 (N_47513,N_40430,N_40292);
and U47514 (N_47514,N_43888,N_40967);
xor U47515 (N_47515,N_41471,N_40134);
xor U47516 (N_47516,N_42226,N_42306);
xor U47517 (N_47517,N_44763,N_44774);
xor U47518 (N_47518,N_40158,N_40971);
or U47519 (N_47519,N_40874,N_41791);
nor U47520 (N_47520,N_41186,N_43297);
xnor U47521 (N_47521,N_42748,N_43470);
xor U47522 (N_47522,N_42596,N_41524);
xnor U47523 (N_47523,N_42052,N_40119);
xnor U47524 (N_47524,N_40711,N_42425);
and U47525 (N_47525,N_42757,N_41635);
or U47526 (N_47526,N_40879,N_42652);
nor U47527 (N_47527,N_40203,N_43044);
nor U47528 (N_47528,N_41997,N_44041);
xnor U47529 (N_47529,N_41403,N_44659);
and U47530 (N_47530,N_41803,N_43474);
or U47531 (N_47531,N_43204,N_41038);
and U47532 (N_47532,N_41545,N_42341);
xnor U47533 (N_47533,N_41312,N_41449);
or U47534 (N_47534,N_44797,N_43589);
or U47535 (N_47535,N_43540,N_44604);
nand U47536 (N_47536,N_41499,N_41688);
or U47537 (N_47537,N_44087,N_42976);
nand U47538 (N_47538,N_44211,N_42040);
or U47539 (N_47539,N_41697,N_40133);
nor U47540 (N_47540,N_40575,N_41401);
xnor U47541 (N_47541,N_40832,N_44772);
and U47542 (N_47542,N_43989,N_40550);
and U47543 (N_47543,N_41177,N_44289);
nand U47544 (N_47544,N_40310,N_40563);
nor U47545 (N_47545,N_42479,N_42684);
or U47546 (N_47546,N_40012,N_42995);
xnor U47547 (N_47547,N_41719,N_42472);
nand U47548 (N_47548,N_44866,N_42184);
xnor U47549 (N_47549,N_43292,N_44870);
xor U47550 (N_47550,N_40106,N_40361);
or U47551 (N_47551,N_41824,N_40503);
and U47552 (N_47552,N_44680,N_42553);
xnor U47553 (N_47553,N_43991,N_40539);
or U47554 (N_47554,N_42967,N_40488);
and U47555 (N_47555,N_42308,N_42175);
or U47556 (N_47556,N_40364,N_42781);
and U47557 (N_47557,N_40936,N_42211);
or U47558 (N_47558,N_44423,N_40038);
and U47559 (N_47559,N_41463,N_41212);
or U47560 (N_47560,N_42155,N_44329);
nor U47561 (N_47561,N_42666,N_41815);
xnor U47562 (N_47562,N_40055,N_43919);
nor U47563 (N_47563,N_44086,N_43194);
and U47564 (N_47564,N_41681,N_42438);
xor U47565 (N_47565,N_42764,N_40957);
nand U47566 (N_47566,N_40522,N_44111);
xor U47567 (N_47567,N_42126,N_44824);
xnor U47568 (N_47568,N_44947,N_44816);
and U47569 (N_47569,N_40981,N_41993);
and U47570 (N_47570,N_40558,N_40365);
and U47571 (N_47571,N_44258,N_43607);
xor U47572 (N_47572,N_40393,N_41603);
nor U47573 (N_47573,N_40671,N_44955);
nand U47574 (N_47574,N_41897,N_44797);
nand U47575 (N_47575,N_42560,N_40655);
nor U47576 (N_47576,N_44941,N_43675);
xor U47577 (N_47577,N_43122,N_44917);
xnor U47578 (N_47578,N_42077,N_40589);
and U47579 (N_47579,N_40515,N_41301);
xor U47580 (N_47580,N_44982,N_42574);
or U47581 (N_47581,N_44561,N_41201);
or U47582 (N_47582,N_40343,N_43793);
xor U47583 (N_47583,N_41417,N_42345);
nor U47584 (N_47584,N_40029,N_42318);
or U47585 (N_47585,N_42240,N_41855);
nor U47586 (N_47586,N_43780,N_40657);
and U47587 (N_47587,N_41135,N_40917);
nor U47588 (N_47588,N_40898,N_44564);
nor U47589 (N_47589,N_41589,N_41921);
nor U47590 (N_47590,N_44819,N_40015);
or U47591 (N_47591,N_41558,N_44413);
nor U47592 (N_47592,N_43460,N_41359);
nor U47593 (N_47593,N_41422,N_41767);
and U47594 (N_47594,N_41661,N_44268);
and U47595 (N_47595,N_42438,N_40494);
and U47596 (N_47596,N_40828,N_44269);
or U47597 (N_47597,N_42651,N_41076);
nand U47598 (N_47598,N_44456,N_41801);
and U47599 (N_47599,N_40308,N_43960);
and U47600 (N_47600,N_40388,N_41819);
xor U47601 (N_47601,N_40257,N_41180);
xnor U47602 (N_47602,N_43355,N_42782);
or U47603 (N_47603,N_42275,N_44595);
and U47604 (N_47604,N_40376,N_41325);
nor U47605 (N_47605,N_43371,N_43524);
or U47606 (N_47606,N_40480,N_43018);
xor U47607 (N_47607,N_43984,N_44965);
or U47608 (N_47608,N_42306,N_43767);
xor U47609 (N_47609,N_42708,N_44638);
nor U47610 (N_47610,N_42982,N_44986);
and U47611 (N_47611,N_41648,N_44295);
nor U47612 (N_47612,N_40049,N_43929);
nor U47613 (N_47613,N_44864,N_43747);
nand U47614 (N_47614,N_42119,N_44262);
and U47615 (N_47615,N_44983,N_43782);
nand U47616 (N_47616,N_43745,N_41883);
xnor U47617 (N_47617,N_44207,N_42890);
xnor U47618 (N_47618,N_42377,N_43936);
nand U47619 (N_47619,N_43403,N_41230);
or U47620 (N_47620,N_42073,N_41163);
nor U47621 (N_47621,N_43882,N_43363);
or U47622 (N_47622,N_41906,N_41330);
xor U47623 (N_47623,N_40359,N_42619);
or U47624 (N_47624,N_42103,N_44344);
nor U47625 (N_47625,N_43849,N_41309);
or U47626 (N_47626,N_41745,N_40228);
nor U47627 (N_47627,N_40136,N_42694);
xor U47628 (N_47628,N_43818,N_41970);
nand U47629 (N_47629,N_42500,N_42205);
nand U47630 (N_47630,N_40555,N_42265);
or U47631 (N_47631,N_40320,N_40719);
and U47632 (N_47632,N_41639,N_43128);
or U47633 (N_47633,N_41166,N_44620);
nand U47634 (N_47634,N_41596,N_42187);
nor U47635 (N_47635,N_44656,N_43025);
nand U47636 (N_47636,N_40000,N_42199);
nor U47637 (N_47637,N_44235,N_40762);
and U47638 (N_47638,N_41943,N_44713);
nor U47639 (N_47639,N_40800,N_40530);
or U47640 (N_47640,N_44789,N_42601);
nor U47641 (N_47641,N_42351,N_41813);
and U47642 (N_47642,N_43957,N_40109);
nor U47643 (N_47643,N_44081,N_42473);
or U47644 (N_47644,N_41025,N_43737);
nor U47645 (N_47645,N_43776,N_42639);
xnor U47646 (N_47646,N_44826,N_40580);
nand U47647 (N_47647,N_42042,N_43092);
xnor U47648 (N_47648,N_44599,N_44046);
xor U47649 (N_47649,N_44276,N_43768);
nand U47650 (N_47650,N_42092,N_44190);
nand U47651 (N_47651,N_41776,N_40675);
xor U47652 (N_47652,N_40939,N_43153);
and U47653 (N_47653,N_43070,N_40631);
nand U47654 (N_47654,N_40578,N_42655);
and U47655 (N_47655,N_44846,N_41291);
or U47656 (N_47656,N_43603,N_40694);
xnor U47657 (N_47657,N_41809,N_42492);
xor U47658 (N_47658,N_41117,N_43851);
nor U47659 (N_47659,N_40493,N_44652);
nand U47660 (N_47660,N_44877,N_42562);
xor U47661 (N_47661,N_41367,N_43017);
xnor U47662 (N_47662,N_43430,N_44543);
nor U47663 (N_47663,N_40219,N_43609);
nor U47664 (N_47664,N_42550,N_40756);
and U47665 (N_47665,N_42466,N_44947);
nor U47666 (N_47666,N_44507,N_44773);
nor U47667 (N_47667,N_40349,N_40613);
nand U47668 (N_47668,N_44532,N_44024);
xnor U47669 (N_47669,N_41977,N_41042);
xnor U47670 (N_47670,N_41997,N_44894);
and U47671 (N_47671,N_43818,N_44681);
nand U47672 (N_47672,N_41200,N_44085);
or U47673 (N_47673,N_43324,N_42994);
nand U47674 (N_47674,N_40520,N_43693);
nand U47675 (N_47675,N_44095,N_43403);
nor U47676 (N_47676,N_44453,N_40840);
nor U47677 (N_47677,N_40318,N_42021);
and U47678 (N_47678,N_42846,N_41350);
xor U47679 (N_47679,N_44190,N_44799);
nor U47680 (N_47680,N_44088,N_43772);
or U47681 (N_47681,N_44625,N_42076);
nand U47682 (N_47682,N_42110,N_41574);
nor U47683 (N_47683,N_44049,N_43421);
nand U47684 (N_47684,N_40315,N_42273);
nand U47685 (N_47685,N_40799,N_44114);
nor U47686 (N_47686,N_40343,N_41417);
xnor U47687 (N_47687,N_43932,N_41547);
or U47688 (N_47688,N_42708,N_41420);
and U47689 (N_47689,N_41388,N_40076);
and U47690 (N_47690,N_43234,N_41129);
xnor U47691 (N_47691,N_44571,N_40436);
or U47692 (N_47692,N_44433,N_44914);
and U47693 (N_47693,N_42914,N_44222);
xnor U47694 (N_47694,N_41799,N_44713);
nor U47695 (N_47695,N_44830,N_41437);
nand U47696 (N_47696,N_44500,N_43034);
nor U47697 (N_47697,N_41861,N_42203);
or U47698 (N_47698,N_42509,N_40543);
nor U47699 (N_47699,N_41586,N_44970);
nand U47700 (N_47700,N_40865,N_44325);
and U47701 (N_47701,N_42461,N_41684);
nand U47702 (N_47702,N_40852,N_41889);
nor U47703 (N_47703,N_43182,N_44422);
and U47704 (N_47704,N_40383,N_43200);
nand U47705 (N_47705,N_42961,N_44938);
xor U47706 (N_47706,N_43412,N_41205);
and U47707 (N_47707,N_41595,N_40451);
nor U47708 (N_47708,N_40165,N_42989);
nand U47709 (N_47709,N_44703,N_41399);
or U47710 (N_47710,N_42987,N_40110);
or U47711 (N_47711,N_42320,N_44198);
or U47712 (N_47712,N_44080,N_42609);
or U47713 (N_47713,N_44949,N_40380);
xor U47714 (N_47714,N_41180,N_41245);
and U47715 (N_47715,N_40281,N_44993);
and U47716 (N_47716,N_42776,N_40871);
nor U47717 (N_47717,N_43257,N_42696);
xnor U47718 (N_47718,N_41725,N_42602);
or U47719 (N_47719,N_42332,N_44265);
nand U47720 (N_47720,N_43626,N_44177);
or U47721 (N_47721,N_41280,N_44896);
xor U47722 (N_47722,N_43526,N_41169);
and U47723 (N_47723,N_41837,N_42448);
nand U47724 (N_47724,N_42842,N_42908);
nand U47725 (N_47725,N_42160,N_44063);
xor U47726 (N_47726,N_40562,N_43184);
or U47727 (N_47727,N_40052,N_44763);
and U47728 (N_47728,N_43240,N_43149);
or U47729 (N_47729,N_44291,N_44024);
nand U47730 (N_47730,N_40394,N_41736);
nor U47731 (N_47731,N_44643,N_42529);
and U47732 (N_47732,N_44033,N_43596);
xor U47733 (N_47733,N_44414,N_41736);
or U47734 (N_47734,N_44737,N_43681);
and U47735 (N_47735,N_42373,N_43526);
nand U47736 (N_47736,N_43466,N_43666);
xor U47737 (N_47737,N_43340,N_41619);
nor U47738 (N_47738,N_41673,N_42330);
xnor U47739 (N_47739,N_44236,N_40235);
nor U47740 (N_47740,N_40275,N_41613);
and U47741 (N_47741,N_42875,N_41273);
or U47742 (N_47742,N_41180,N_41363);
xor U47743 (N_47743,N_41571,N_43860);
nor U47744 (N_47744,N_44398,N_41157);
and U47745 (N_47745,N_42303,N_40097);
or U47746 (N_47746,N_41858,N_44149);
nand U47747 (N_47747,N_41054,N_40096);
nor U47748 (N_47748,N_44108,N_43781);
nor U47749 (N_47749,N_40460,N_41165);
or U47750 (N_47750,N_44046,N_41994);
or U47751 (N_47751,N_40576,N_42503);
or U47752 (N_47752,N_42236,N_40726);
nor U47753 (N_47753,N_42975,N_42704);
or U47754 (N_47754,N_40690,N_44001);
and U47755 (N_47755,N_42230,N_41759);
and U47756 (N_47756,N_43753,N_40832);
and U47757 (N_47757,N_40930,N_41862);
xnor U47758 (N_47758,N_40985,N_41207);
and U47759 (N_47759,N_42098,N_42660);
nor U47760 (N_47760,N_40542,N_40692);
nand U47761 (N_47761,N_40283,N_44657);
xnor U47762 (N_47762,N_44985,N_41810);
xnor U47763 (N_47763,N_40474,N_42569);
and U47764 (N_47764,N_44141,N_42831);
or U47765 (N_47765,N_40813,N_44302);
and U47766 (N_47766,N_44055,N_40618);
and U47767 (N_47767,N_40151,N_44943);
nand U47768 (N_47768,N_44476,N_44212);
xor U47769 (N_47769,N_42921,N_44697);
nand U47770 (N_47770,N_44279,N_41749);
nand U47771 (N_47771,N_44049,N_44593);
xor U47772 (N_47772,N_44603,N_44251);
nand U47773 (N_47773,N_41989,N_40571);
xor U47774 (N_47774,N_44583,N_41408);
and U47775 (N_47775,N_43304,N_40891);
or U47776 (N_47776,N_44925,N_42684);
and U47777 (N_47777,N_42602,N_41660);
or U47778 (N_47778,N_42982,N_40144);
xnor U47779 (N_47779,N_44114,N_43672);
and U47780 (N_47780,N_41098,N_42488);
and U47781 (N_47781,N_43216,N_44729);
nand U47782 (N_47782,N_44030,N_43059);
or U47783 (N_47783,N_43094,N_40383);
and U47784 (N_47784,N_42929,N_44307);
nor U47785 (N_47785,N_41128,N_43143);
nor U47786 (N_47786,N_42690,N_43691);
or U47787 (N_47787,N_41701,N_42606);
nor U47788 (N_47788,N_43962,N_40092);
xnor U47789 (N_47789,N_43581,N_41060);
nor U47790 (N_47790,N_44299,N_42020);
nor U47791 (N_47791,N_41997,N_42435);
and U47792 (N_47792,N_43514,N_41407);
and U47793 (N_47793,N_40992,N_44137);
or U47794 (N_47794,N_44347,N_40990);
nand U47795 (N_47795,N_42711,N_43219);
and U47796 (N_47796,N_42140,N_44480);
xnor U47797 (N_47797,N_42571,N_42155);
nand U47798 (N_47798,N_40708,N_43896);
nor U47799 (N_47799,N_44331,N_44737);
or U47800 (N_47800,N_42669,N_41523);
nor U47801 (N_47801,N_40031,N_44036);
and U47802 (N_47802,N_40461,N_42603);
nor U47803 (N_47803,N_43121,N_42199);
or U47804 (N_47804,N_42755,N_41158);
nor U47805 (N_47805,N_42137,N_44378);
nand U47806 (N_47806,N_41783,N_41247);
nand U47807 (N_47807,N_41572,N_42016);
xnor U47808 (N_47808,N_40296,N_42769);
and U47809 (N_47809,N_44537,N_42121);
and U47810 (N_47810,N_41785,N_42798);
xor U47811 (N_47811,N_41269,N_44856);
or U47812 (N_47812,N_40244,N_40159);
xnor U47813 (N_47813,N_40542,N_41971);
xor U47814 (N_47814,N_42816,N_42041);
or U47815 (N_47815,N_44425,N_41790);
nor U47816 (N_47816,N_44716,N_43584);
or U47817 (N_47817,N_44194,N_40061);
nor U47818 (N_47818,N_41024,N_40837);
nand U47819 (N_47819,N_41986,N_42502);
nor U47820 (N_47820,N_44056,N_44159);
or U47821 (N_47821,N_44963,N_44526);
or U47822 (N_47822,N_41759,N_44391);
and U47823 (N_47823,N_40324,N_44896);
xnor U47824 (N_47824,N_43208,N_44664);
or U47825 (N_47825,N_42737,N_40218);
nor U47826 (N_47826,N_44906,N_40023);
or U47827 (N_47827,N_40826,N_43148);
xor U47828 (N_47828,N_42800,N_41791);
nand U47829 (N_47829,N_43479,N_42232);
and U47830 (N_47830,N_44512,N_40321);
nand U47831 (N_47831,N_41234,N_41776);
and U47832 (N_47832,N_43858,N_41592);
and U47833 (N_47833,N_43202,N_42137);
or U47834 (N_47834,N_42925,N_40414);
or U47835 (N_47835,N_41345,N_40933);
nand U47836 (N_47836,N_42501,N_43371);
or U47837 (N_47837,N_41110,N_44484);
nand U47838 (N_47838,N_41014,N_43690);
or U47839 (N_47839,N_42334,N_42404);
and U47840 (N_47840,N_40619,N_40746);
nand U47841 (N_47841,N_40184,N_41420);
or U47842 (N_47842,N_40984,N_42628);
xor U47843 (N_47843,N_41956,N_42008);
or U47844 (N_47844,N_42985,N_40191);
and U47845 (N_47845,N_44504,N_44363);
or U47846 (N_47846,N_43574,N_43944);
and U47847 (N_47847,N_43072,N_41165);
and U47848 (N_47848,N_44233,N_44200);
and U47849 (N_47849,N_43903,N_44982);
nor U47850 (N_47850,N_42960,N_42267);
nor U47851 (N_47851,N_43349,N_44433);
and U47852 (N_47852,N_43374,N_43843);
or U47853 (N_47853,N_41462,N_42029);
or U47854 (N_47854,N_42131,N_42072);
xnor U47855 (N_47855,N_43463,N_40167);
nor U47856 (N_47856,N_42233,N_44044);
or U47857 (N_47857,N_44731,N_42082);
nor U47858 (N_47858,N_41199,N_43194);
and U47859 (N_47859,N_42292,N_42200);
or U47860 (N_47860,N_41575,N_43090);
and U47861 (N_47861,N_42820,N_43759);
xor U47862 (N_47862,N_42492,N_42414);
nand U47863 (N_47863,N_43402,N_42743);
nand U47864 (N_47864,N_40790,N_40443);
or U47865 (N_47865,N_40376,N_40406);
xnor U47866 (N_47866,N_44523,N_43573);
xnor U47867 (N_47867,N_43539,N_44670);
nor U47868 (N_47868,N_44068,N_40049);
and U47869 (N_47869,N_40670,N_42541);
xor U47870 (N_47870,N_43155,N_41075);
xnor U47871 (N_47871,N_43883,N_43763);
and U47872 (N_47872,N_43581,N_42276);
nor U47873 (N_47873,N_40211,N_43380);
xnor U47874 (N_47874,N_44925,N_44312);
and U47875 (N_47875,N_42097,N_41322);
xor U47876 (N_47876,N_40709,N_43410);
nor U47877 (N_47877,N_41164,N_43065);
or U47878 (N_47878,N_42691,N_43298);
xor U47879 (N_47879,N_44281,N_42777);
nand U47880 (N_47880,N_40365,N_41691);
xor U47881 (N_47881,N_44573,N_42453);
or U47882 (N_47882,N_40760,N_40843);
and U47883 (N_47883,N_44333,N_41494);
or U47884 (N_47884,N_44303,N_40899);
xor U47885 (N_47885,N_40447,N_41883);
or U47886 (N_47886,N_41837,N_42384);
nand U47887 (N_47887,N_40126,N_40412);
or U47888 (N_47888,N_42625,N_43082);
and U47889 (N_47889,N_43250,N_40255);
nand U47890 (N_47890,N_43943,N_40038);
nor U47891 (N_47891,N_40487,N_44954);
nand U47892 (N_47892,N_41666,N_43389);
nand U47893 (N_47893,N_43624,N_42076);
nor U47894 (N_47894,N_40316,N_44971);
xor U47895 (N_47895,N_41989,N_43327);
nand U47896 (N_47896,N_40674,N_44551);
nand U47897 (N_47897,N_43144,N_43158);
nand U47898 (N_47898,N_40331,N_41081);
nor U47899 (N_47899,N_44233,N_42240);
and U47900 (N_47900,N_41919,N_42336);
or U47901 (N_47901,N_41745,N_43815);
nor U47902 (N_47902,N_44636,N_43675);
or U47903 (N_47903,N_41659,N_42053);
nor U47904 (N_47904,N_40491,N_41725);
nor U47905 (N_47905,N_42405,N_44107);
nor U47906 (N_47906,N_41071,N_44534);
and U47907 (N_47907,N_44014,N_42530);
or U47908 (N_47908,N_41526,N_40666);
and U47909 (N_47909,N_42605,N_43785);
or U47910 (N_47910,N_40518,N_41195);
and U47911 (N_47911,N_43501,N_43128);
xor U47912 (N_47912,N_41522,N_42354);
nand U47913 (N_47913,N_40911,N_44374);
or U47914 (N_47914,N_42764,N_41848);
nor U47915 (N_47915,N_44889,N_43420);
nand U47916 (N_47916,N_40819,N_43792);
or U47917 (N_47917,N_42862,N_41978);
nor U47918 (N_47918,N_40670,N_41818);
and U47919 (N_47919,N_44349,N_41880);
or U47920 (N_47920,N_40384,N_43631);
and U47921 (N_47921,N_42124,N_40583);
or U47922 (N_47922,N_42156,N_41564);
xor U47923 (N_47923,N_44211,N_42638);
nor U47924 (N_47924,N_40500,N_42010);
xnor U47925 (N_47925,N_42004,N_44557);
nand U47926 (N_47926,N_44365,N_44354);
and U47927 (N_47927,N_43901,N_43749);
or U47928 (N_47928,N_44146,N_44155);
nor U47929 (N_47929,N_43031,N_43193);
and U47930 (N_47930,N_44953,N_44566);
or U47931 (N_47931,N_43027,N_43170);
and U47932 (N_47932,N_41886,N_41661);
nand U47933 (N_47933,N_43869,N_40704);
nor U47934 (N_47934,N_40990,N_40150);
nand U47935 (N_47935,N_42957,N_44668);
and U47936 (N_47936,N_42508,N_43471);
or U47937 (N_47937,N_41976,N_42433);
nand U47938 (N_47938,N_44623,N_43748);
and U47939 (N_47939,N_42103,N_41098);
or U47940 (N_47940,N_44855,N_44027);
or U47941 (N_47941,N_43332,N_43637);
xnor U47942 (N_47942,N_40353,N_44068);
nor U47943 (N_47943,N_42079,N_40154);
and U47944 (N_47944,N_44642,N_41650);
and U47945 (N_47945,N_42852,N_42105);
and U47946 (N_47946,N_44454,N_40218);
or U47947 (N_47947,N_41524,N_44516);
or U47948 (N_47948,N_42081,N_42939);
and U47949 (N_47949,N_40319,N_42622);
or U47950 (N_47950,N_40235,N_42621);
or U47951 (N_47951,N_41315,N_40689);
or U47952 (N_47952,N_43360,N_43926);
nor U47953 (N_47953,N_44492,N_41956);
or U47954 (N_47954,N_43442,N_40779);
nand U47955 (N_47955,N_41400,N_43320);
nor U47956 (N_47956,N_42694,N_43897);
xnor U47957 (N_47957,N_43730,N_43227);
xor U47958 (N_47958,N_40767,N_40642);
nor U47959 (N_47959,N_44582,N_44246);
nand U47960 (N_47960,N_40892,N_42830);
xor U47961 (N_47961,N_42991,N_43705);
nand U47962 (N_47962,N_42641,N_44265);
and U47963 (N_47963,N_40225,N_41897);
xor U47964 (N_47964,N_42060,N_40859);
nor U47965 (N_47965,N_42304,N_43194);
or U47966 (N_47966,N_40881,N_42635);
xor U47967 (N_47967,N_43850,N_40749);
or U47968 (N_47968,N_41181,N_44630);
and U47969 (N_47969,N_40042,N_42828);
nor U47970 (N_47970,N_42957,N_40792);
xor U47971 (N_47971,N_43995,N_41629);
nand U47972 (N_47972,N_42980,N_42583);
and U47973 (N_47973,N_43436,N_40102);
nand U47974 (N_47974,N_42388,N_41970);
nor U47975 (N_47975,N_42627,N_42184);
nand U47976 (N_47976,N_44378,N_43787);
or U47977 (N_47977,N_40534,N_41450);
xnor U47978 (N_47978,N_41006,N_41983);
nand U47979 (N_47979,N_41133,N_44254);
or U47980 (N_47980,N_41734,N_42428);
and U47981 (N_47981,N_42033,N_43635);
xor U47982 (N_47982,N_42513,N_41661);
nand U47983 (N_47983,N_42217,N_44748);
or U47984 (N_47984,N_42081,N_41100);
nand U47985 (N_47985,N_44965,N_41150);
and U47986 (N_47986,N_41895,N_44322);
nor U47987 (N_47987,N_42232,N_44402);
or U47988 (N_47988,N_42388,N_42679);
nand U47989 (N_47989,N_41958,N_41490);
and U47990 (N_47990,N_41073,N_41862);
nor U47991 (N_47991,N_44451,N_44450);
nor U47992 (N_47992,N_42487,N_44041);
nor U47993 (N_47993,N_40530,N_42526);
xor U47994 (N_47994,N_44040,N_43893);
or U47995 (N_47995,N_40464,N_42103);
xor U47996 (N_47996,N_44077,N_44431);
xor U47997 (N_47997,N_43663,N_44633);
and U47998 (N_47998,N_43822,N_43713);
nand U47999 (N_47999,N_40613,N_44157);
xnor U48000 (N_48000,N_42894,N_44995);
nand U48001 (N_48001,N_44997,N_40990);
and U48002 (N_48002,N_44668,N_43359);
and U48003 (N_48003,N_44729,N_40192);
nor U48004 (N_48004,N_40784,N_41710);
and U48005 (N_48005,N_44413,N_42296);
xnor U48006 (N_48006,N_44793,N_40407);
nor U48007 (N_48007,N_43924,N_44977);
and U48008 (N_48008,N_42657,N_43054);
or U48009 (N_48009,N_43340,N_43545);
nor U48010 (N_48010,N_44408,N_41260);
xor U48011 (N_48011,N_43378,N_44992);
nand U48012 (N_48012,N_43799,N_43211);
or U48013 (N_48013,N_43297,N_43730);
nand U48014 (N_48014,N_41211,N_41790);
or U48015 (N_48015,N_41704,N_44862);
nand U48016 (N_48016,N_41821,N_42104);
nand U48017 (N_48017,N_43543,N_44776);
or U48018 (N_48018,N_43193,N_41216);
nor U48019 (N_48019,N_44113,N_41157);
and U48020 (N_48020,N_40995,N_43608);
xnor U48021 (N_48021,N_42955,N_43232);
nor U48022 (N_48022,N_43471,N_44405);
or U48023 (N_48023,N_42186,N_44318);
nor U48024 (N_48024,N_40914,N_44363);
or U48025 (N_48025,N_44207,N_42779);
and U48026 (N_48026,N_43531,N_42530);
xnor U48027 (N_48027,N_41611,N_40485);
nand U48028 (N_48028,N_44470,N_41266);
or U48029 (N_48029,N_43010,N_40600);
and U48030 (N_48030,N_41822,N_41122);
and U48031 (N_48031,N_43053,N_41225);
xnor U48032 (N_48032,N_44148,N_43611);
and U48033 (N_48033,N_44186,N_44447);
xor U48034 (N_48034,N_42932,N_43837);
xnor U48035 (N_48035,N_44822,N_44953);
or U48036 (N_48036,N_42713,N_40921);
nand U48037 (N_48037,N_40319,N_43439);
nand U48038 (N_48038,N_41790,N_44906);
or U48039 (N_48039,N_42803,N_44773);
and U48040 (N_48040,N_42697,N_42622);
and U48041 (N_48041,N_43491,N_42842);
xnor U48042 (N_48042,N_43418,N_42875);
or U48043 (N_48043,N_43517,N_43678);
or U48044 (N_48044,N_44102,N_44334);
and U48045 (N_48045,N_43502,N_44914);
or U48046 (N_48046,N_44144,N_41570);
nand U48047 (N_48047,N_42465,N_44533);
nand U48048 (N_48048,N_40960,N_41103);
nor U48049 (N_48049,N_43261,N_43857);
and U48050 (N_48050,N_43897,N_41631);
and U48051 (N_48051,N_44272,N_42109);
and U48052 (N_48052,N_44969,N_43949);
or U48053 (N_48053,N_42198,N_42703);
and U48054 (N_48054,N_44746,N_43510);
xnor U48055 (N_48055,N_42970,N_42281);
xnor U48056 (N_48056,N_44663,N_40385);
xor U48057 (N_48057,N_41246,N_43990);
or U48058 (N_48058,N_41926,N_41778);
nand U48059 (N_48059,N_44648,N_44017);
xnor U48060 (N_48060,N_42438,N_42878);
xor U48061 (N_48061,N_44435,N_44975);
nand U48062 (N_48062,N_41022,N_43349);
nand U48063 (N_48063,N_42487,N_40117);
and U48064 (N_48064,N_40012,N_44391);
and U48065 (N_48065,N_40257,N_43256);
nor U48066 (N_48066,N_41485,N_42206);
xnor U48067 (N_48067,N_43962,N_44833);
nor U48068 (N_48068,N_41731,N_40657);
nand U48069 (N_48069,N_44740,N_41362);
xor U48070 (N_48070,N_40123,N_43157);
nand U48071 (N_48071,N_43100,N_42817);
nor U48072 (N_48072,N_44558,N_40046);
or U48073 (N_48073,N_43695,N_43038);
xnor U48074 (N_48074,N_40369,N_44189);
xor U48075 (N_48075,N_42524,N_43367);
or U48076 (N_48076,N_40591,N_44165);
xor U48077 (N_48077,N_42183,N_42280);
nand U48078 (N_48078,N_42098,N_43615);
xnor U48079 (N_48079,N_44117,N_44474);
or U48080 (N_48080,N_40313,N_42939);
nand U48081 (N_48081,N_42360,N_41677);
nor U48082 (N_48082,N_40002,N_43184);
nor U48083 (N_48083,N_42013,N_44460);
and U48084 (N_48084,N_44453,N_43638);
xor U48085 (N_48085,N_43163,N_44735);
or U48086 (N_48086,N_41801,N_44270);
or U48087 (N_48087,N_40175,N_40965);
and U48088 (N_48088,N_41763,N_42820);
nand U48089 (N_48089,N_42098,N_43514);
nand U48090 (N_48090,N_42499,N_44370);
nor U48091 (N_48091,N_43967,N_44548);
and U48092 (N_48092,N_42528,N_44850);
or U48093 (N_48093,N_40533,N_43733);
nor U48094 (N_48094,N_43058,N_43011);
and U48095 (N_48095,N_42023,N_42926);
nor U48096 (N_48096,N_40918,N_44115);
nor U48097 (N_48097,N_41088,N_42313);
or U48098 (N_48098,N_40811,N_41344);
and U48099 (N_48099,N_44844,N_40953);
nand U48100 (N_48100,N_42915,N_41448);
xor U48101 (N_48101,N_43441,N_43999);
xor U48102 (N_48102,N_44044,N_41686);
xnor U48103 (N_48103,N_44204,N_41471);
and U48104 (N_48104,N_42132,N_41616);
nor U48105 (N_48105,N_43963,N_43739);
xor U48106 (N_48106,N_43104,N_40921);
or U48107 (N_48107,N_40026,N_44180);
nand U48108 (N_48108,N_40385,N_44049);
xor U48109 (N_48109,N_41865,N_42969);
or U48110 (N_48110,N_41198,N_44661);
or U48111 (N_48111,N_40622,N_41290);
nand U48112 (N_48112,N_41840,N_40756);
or U48113 (N_48113,N_44182,N_40383);
xor U48114 (N_48114,N_43947,N_44009);
xnor U48115 (N_48115,N_41510,N_40751);
nor U48116 (N_48116,N_42910,N_42808);
nor U48117 (N_48117,N_40460,N_42978);
nor U48118 (N_48118,N_43995,N_41772);
nor U48119 (N_48119,N_43152,N_41520);
and U48120 (N_48120,N_40436,N_41765);
nand U48121 (N_48121,N_41061,N_42981);
xnor U48122 (N_48122,N_40395,N_42740);
nand U48123 (N_48123,N_43064,N_44011);
xor U48124 (N_48124,N_41363,N_41641);
nor U48125 (N_48125,N_41378,N_40681);
nand U48126 (N_48126,N_44615,N_41716);
and U48127 (N_48127,N_40084,N_44225);
nor U48128 (N_48128,N_44197,N_41109);
or U48129 (N_48129,N_40527,N_43811);
nor U48130 (N_48130,N_40459,N_44029);
nor U48131 (N_48131,N_41292,N_40150);
and U48132 (N_48132,N_43679,N_41896);
nand U48133 (N_48133,N_44170,N_42926);
nor U48134 (N_48134,N_42032,N_44474);
xnor U48135 (N_48135,N_44228,N_42531);
nand U48136 (N_48136,N_40242,N_41268);
nor U48137 (N_48137,N_42837,N_44474);
or U48138 (N_48138,N_42584,N_43406);
nor U48139 (N_48139,N_42218,N_43359);
or U48140 (N_48140,N_44856,N_40108);
or U48141 (N_48141,N_40674,N_42138);
nor U48142 (N_48142,N_43271,N_44661);
nor U48143 (N_48143,N_40839,N_40950);
and U48144 (N_48144,N_44681,N_40200);
or U48145 (N_48145,N_44851,N_44008);
or U48146 (N_48146,N_42330,N_44985);
nor U48147 (N_48147,N_44887,N_42982);
or U48148 (N_48148,N_41781,N_44554);
or U48149 (N_48149,N_42753,N_41640);
xnor U48150 (N_48150,N_42330,N_41537);
nand U48151 (N_48151,N_41532,N_44551);
or U48152 (N_48152,N_41460,N_40796);
and U48153 (N_48153,N_40652,N_40251);
and U48154 (N_48154,N_40657,N_43621);
nor U48155 (N_48155,N_43878,N_42708);
nor U48156 (N_48156,N_40879,N_44841);
or U48157 (N_48157,N_42470,N_41439);
nor U48158 (N_48158,N_41552,N_44046);
nand U48159 (N_48159,N_40377,N_43027);
nor U48160 (N_48160,N_42275,N_40578);
and U48161 (N_48161,N_40683,N_40154);
or U48162 (N_48162,N_43327,N_40599);
nor U48163 (N_48163,N_44597,N_41292);
nand U48164 (N_48164,N_40912,N_41713);
xor U48165 (N_48165,N_41116,N_44385);
or U48166 (N_48166,N_41543,N_40511);
nand U48167 (N_48167,N_43680,N_44406);
and U48168 (N_48168,N_41917,N_40481);
xnor U48169 (N_48169,N_40276,N_44315);
or U48170 (N_48170,N_40212,N_44300);
nor U48171 (N_48171,N_41667,N_42354);
xnor U48172 (N_48172,N_40878,N_42609);
or U48173 (N_48173,N_42013,N_42725);
and U48174 (N_48174,N_42589,N_44201);
nand U48175 (N_48175,N_41653,N_43636);
nor U48176 (N_48176,N_44413,N_40764);
nand U48177 (N_48177,N_42556,N_42294);
nor U48178 (N_48178,N_40853,N_43300);
nand U48179 (N_48179,N_41282,N_42281);
and U48180 (N_48180,N_41334,N_41078);
or U48181 (N_48181,N_43406,N_44834);
xor U48182 (N_48182,N_40805,N_44420);
or U48183 (N_48183,N_40827,N_40950);
nand U48184 (N_48184,N_40904,N_44140);
nand U48185 (N_48185,N_44820,N_41350);
nor U48186 (N_48186,N_43687,N_40326);
nand U48187 (N_48187,N_41204,N_43406);
nor U48188 (N_48188,N_42302,N_42391);
or U48189 (N_48189,N_44060,N_43539);
nor U48190 (N_48190,N_44835,N_40716);
and U48191 (N_48191,N_40502,N_42042);
xnor U48192 (N_48192,N_44549,N_44922);
nor U48193 (N_48193,N_44741,N_40973);
or U48194 (N_48194,N_43066,N_41731);
nor U48195 (N_48195,N_41739,N_43069);
xnor U48196 (N_48196,N_44780,N_41634);
nor U48197 (N_48197,N_42774,N_43879);
and U48198 (N_48198,N_42339,N_42993);
xnor U48199 (N_48199,N_44027,N_42007);
or U48200 (N_48200,N_44763,N_40719);
xnor U48201 (N_48201,N_42802,N_43050);
xnor U48202 (N_48202,N_40047,N_43368);
and U48203 (N_48203,N_41541,N_43225);
nand U48204 (N_48204,N_44003,N_40057);
nand U48205 (N_48205,N_41762,N_41986);
xnor U48206 (N_48206,N_41078,N_40568);
or U48207 (N_48207,N_44143,N_43955);
nand U48208 (N_48208,N_40571,N_40140);
nand U48209 (N_48209,N_41803,N_41623);
and U48210 (N_48210,N_40485,N_42560);
and U48211 (N_48211,N_43440,N_43727);
nand U48212 (N_48212,N_42758,N_41499);
nand U48213 (N_48213,N_40462,N_41809);
nand U48214 (N_48214,N_44293,N_44377);
or U48215 (N_48215,N_41582,N_41871);
nor U48216 (N_48216,N_41376,N_43248);
and U48217 (N_48217,N_42708,N_40131);
and U48218 (N_48218,N_42727,N_43263);
nand U48219 (N_48219,N_44964,N_44075);
or U48220 (N_48220,N_43605,N_42249);
nor U48221 (N_48221,N_41025,N_40307);
or U48222 (N_48222,N_42789,N_40893);
nand U48223 (N_48223,N_44298,N_40313);
xnor U48224 (N_48224,N_43378,N_42832);
and U48225 (N_48225,N_41339,N_44090);
nand U48226 (N_48226,N_42180,N_41136);
or U48227 (N_48227,N_43035,N_41754);
and U48228 (N_48228,N_43403,N_41728);
or U48229 (N_48229,N_40738,N_42504);
and U48230 (N_48230,N_40191,N_40473);
and U48231 (N_48231,N_42218,N_40041);
xnor U48232 (N_48232,N_42782,N_42492);
xnor U48233 (N_48233,N_44916,N_43869);
nor U48234 (N_48234,N_43611,N_42802);
xnor U48235 (N_48235,N_40810,N_40108);
xor U48236 (N_48236,N_40708,N_41931);
xor U48237 (N_48237,N_43734,N_40114);
nand U48238 (N_48238,N_44891,N_40564);
and U48239 (N_48239,N_44536,N_44123);
nor U48240 (N_48240,N_44829,N_40908);
nand U48241 (N_48241,N_43649,N_41398);
xnor U48242 (N_48242,N_44273,N_41789);
and U48243 (N_48243,N_43911,N_43219);
or U48244 (N_48244,N_40750,N_40098);
and U48245 (N_48245,N_42007,N_40805);
or U48246 (N_48246,N_41923,N_41783);
nor U48247 (N_48247,N_44829,N_42247);
nand U48248 (N_48248,N_40098,N_40823);
xor U48249 (N_48249,N_44397,N_40756);
and U48250 (N_48250,N_41668,N_42843);
xor U48251 (N_48251,N_43750,N_40728);
nor U48252 (N_48252,N_41666,N_41807);
and U48253 (N_48253,N_41096,N_44959);
or U48254 (N_48254,N_40925,N_43045);
nor U48255 (N_48255,N_42624,N_41997);
and U48256 (N_48256,N_43435,N_42944);
nand U48257 (N_48257,N_41596,N_42616);
nor U48258 (N_48258,N_40760,N_40240);
nand U48259 (N_48259,N_41418,N_44003);
and U48260 (N_48260,N_44826,N_41693);
or U48261 (N_48261,N_40745,N_43107);
or U48262 (N_48262,N_44444,N_41404);
or U48263 (N_48263,N_42741,N_44209);
nor U48264 (N_48264,N_44879,N_43931);
and U48265 (N_48265,N_44018,N_40398);
nor U48266 (N_48266,N_40199,N_41175);
xor U48267 (N_48267,N_41538,N_41512);
nand U48268 (N_48268,N_43561,N_44025);
and U48269 (N_48269,N_43669,N_42489);
or U48270 (N_48270,N_41066,N_41977);
nand U48271 (N_48271,N_41424,N_44118);
nand U48272 (N_48272,N_44680,N_41765);
and U48273 (N_48273,N_40169,N_43060);
xnor U48274 (N_48274,N_40182,N_42146);
or U48275 (N_48275,N_41799,N_41286);
or U48276 (N_48276,N_42087,N_40835);
nand U48277 (N_48277,N_43632,N_40993);
nor U48278 (N_48278,N_40318,N_41012);
nand U48279 (N_48279,N_44258,N_41674);
or U48280 (N_48280,N_43675,N_40583);
nor U48281 (N_48281,N_44258,N_40568);
xnor U48282 (N_48282,N_42515,N_40928);
xor U48283 (N_48283,N_41617,N_44383);
nand U48284 (N_48284,N_41996,N_40805);
and U48285 (N_48285,N_41391,N_42237);
nand U48286 (N_48286,N_43194,N_41900);
or U48287 (N_48287,N_41313,N_40846);
and U48288 (N_48288,N_40802,N_42541);
nand U48289 (N_48289,N_43150,N_41932);
or U48290 (N_48290,N_43769,N_44622);
nor U48291 (N_48291,N_40355,N_40322);
nand U48292 (N_48292,N_40867,N_43740);
or U48293 (N_48293,N_44417,N_43000);
nor U48294 (N_48294,N_42840,N_40926);
xnor U48295 (N_48295,N_43524,N_42689);
nor U48296 (N_48296,N_42602,N_43910);
and U48297 (N_48297,N_43715,N_40434);
and U48298 (N_48298,N_44066,N_42215);
or U48299 (N_48299,N_42899,N_42202);
xor U48300 (N_48300,N_41873,N_40912);
or U48301 (N_48301,N_42102,N_43659);
and U48302 (N_48302,N_44754,N_40248);
or U48303 (N_48303,N_42145,N_40854);
and U48304 (N_48304,N_40638,N_41692);
xor U48305 (N_48305,N_44013,N_43665);
xor U48306 (N_48306,N_42698,N_40715);
or U48307 (N_48307,N_41179,N_42728);
nor U48308 (N_48308,N_43869,N_40433);
nor U48309 (N_48309,N_40799,N_40554);
xnor U48310 (N_48310,N_40267,N_42222);
or U48311 (N_48311,N_40626,N_41949);
and U48312 (N_48312,N_43230,N_43007);
nor U48313 (N_48313,N_44785,N_42864);
nor U48314 (N_48314,N_44552,N_44112);
nand U48315 (N_48315,N_40582,N_44715);
and U48316 (N_48316,N_42879,N_40091);
or U48317 (N_48317,N_44924,N_43521);
nand U48318 (N_48318,N_42119,N_44936);
or U48319 (N_48319,N_41692,N_44389);
nor U48320 (N_48320,N_43368,N_40761);
xor U48321 (N_48321,N_44126,N_42847);
nand U48322 (N_48322,N_40920,N_41492);
nor U48323 (N_48323,N_44442,N_42155);
nor U48324 (N_48324,N_42494,N_40702);
or U48325 (N_48325,N_43571,N_42498);
nand U48326 (N_48326,N_41480,N_41360);
or U48327 (N_48327,N_44451,N_40190);
or U48328 (N_48328,N_41496,N_42228);
xor U48329 (N_48329,N_41979,N_40054);
nor U48330 (N_48330,N_43686,N_42692);
xor U48331 (N_48331,N_42792,N_43295);
and U48332 (N_48332,N_43703,N_42326);
and U48333 (N_48333,N_42805,N_44910);
and U48334 (N_48334,N_40570,N_40615);
and U48335 (N_48335,N_40839,N_41800);
xnor U48336 (N_48336,N_41794,N_44926);
or U48337 (N_48337,N_44564,N_42153);
nand U48338 (N_48338,N_43404,N_43514);
nand U48339 (N_48339,N_42581,N_40635);
and U48340 (N_48340,N_41456,N_43403);
nor U48341 (N_48341,N_41220,N_41908);
and U48342 (N_48342,N_40257,N_42805);
nor U48343 (N_48343,N_44397,N_40384);
nor U48344 (N_48344,N_44282,N_42902);
or U48345 (N_48345,N_41338,N_42780);
nand U48346 (N_48346,N_42451,N_43049);
nand U48347 (N_48347,N_40308,N_44001);
nor U48348 (N_48348,N_44249,N_42248);
nand U48349 (N_48349,N_42913,N_43107);
nor U48350 (N_48350,N_40264,N_42193);
or U48351 (N_48351,N_43609,N_40423);
or U48352 (N_48352,N_42211,N_44566);
and U48353 (N_48353,N_44739,N_43677);
nand U48354 (N_48354,N_40638,N_43419);
nor U48355 (N_48355,N_42561,N_41307);
xnor U48356 (N_48356,N_41176,N_42443);
xor U48357 (N_48357,N_42209,N_43590);
or U48358 (N_48358,N_40214,N_41715);
and U48359 (N_48359,N_44605,N_40464);
or U48360 (N_48360,N_40932,N_41736);
or U48361 (N_48361,N_41524,N_43995);
or U48362 (N_48362,N_42968,N_42282);
and U48363 (N_48363,N_43272,N_43594);
and U48364 (N_48364,N_43763,N_43760);
and U48365 (N_48365,N_42561,N_43525);
nor U48366 (N_48366,N_44612,N_43928);
nor U48367 (N_48367,N_40454,N_43878);
nand U48368 (N_48368,N_41352,N_43034);
or U48369 (N_48369,N_40292,N_42420);
or U48370 (N_48370,N_41025,N_42930);
or U48371 (N_48371,N_43299,N_40151);
xnor U48372 (N_48372,N_42070,N_40032);
nor U48373 (N_48373,N_41596,N_42198);
nand U48374 (N_48374,N_44258,N_41954);
nor U48375 (N_48375,N_40018,N_41182);
xor U48376 (N_48376,N_40777,N_44551);
xnor U48377 (N_48377,N_41221,N_40238);
and U48378 (N_48378,N_41018,N_40295);
xnor U48379 (N_48379,N_40086,N_41052);
or U48380 (N_48380,N_44791,N_41129);
xnor U48381 (N_48381,N_43429,N_43773);
nor U48382 (N_48382,N_40283,N_44630);
nor U48383 (N_48383,N_41282,N_44901);
and U48384 (N_48384,N_43051,N_44208);
nor U48385 (N_48385,N_41942,N_44265);
or U48386 (N_48386,N_40852,N_44796);
or U48387 (N_48387,N_42984,N_42210);
or U48388 (N_48388,N_42988,N_41137);
nand U48389 (N_48389,N_40701,N_43046);
nand U48390 (N_48390,N_44356,N_40957);
xnor U48391 (N_48391,N_42086,N_42630);
or U48392 (N_48392,N_42001,N_43915);
xor U48393 (N_48393,N_42811,N_43963);
nand U48394 (N_48394,N_41849,N_43162);
nand U48395 (N_48395,N_44582,N_40465);
nand U48396 (N_48396,N_44006,N_44976);
or U48397 (N_48397,N_40823,N_42931);
or U48398 (N_48398,N_44010,N_40534);
nor U48399 (N_48399,N_42400,N_43332);
nand U48400 (N_48400,N_40230,N_42284);
and U48401 (N_48401,N_41356,N_41411);
nor U48402 (N_48402,N_42364,N_41296);
and U48403 (N_48403,N_41770,N_42579);
and U48404 (N_48404,N_44015,N_42596);
or U48405 (N_48405,N_44735,N_41712);
and U48406 (N_48406,N_43266,N_40586);
nor U48407 (N_48407,N_43512,N_41378);
or U48408 (N_48408,N_43033,N_41933);
nand U48409 (N_48409,N_42034,N_42161);
or U48410 (N_48410,N_40229,N_42126);
nand U48411 (N_48411,N_40468,N_42351);
and U48412 (N_48412,N_42420,N_44013);
xnor U48413 (N_48413,N_42350,N_44718);
or U48414 (N_48414,N_43282,N_43554);
and U48415 (N_48415,N_42046,N_41275);
and U48416 (N_48416,N_40872,N_41272);
nor U48417 (N_48417,N_40642,N_40778);
or U48418 (N_48418,N_44984,N_43492);
nand U48419 (N_48419,N_42031,N_42836);
nand U48420 (N_48420,N_41427,N_44119);
nand U48421 (N_48421,N_42789,N_41071);
xor U48422 (N_48422,N_43335,N_44234);
nand U48423 (N_48423,N_44222,N_44068);
nor U48424 (N_48424,N_41588,N_41661);
xnor U48425 (N_48425,N_42542,N_40937);
and U48426 (N_48426,N_44102,N_40724);
nor U48427 (N_48427,N_43525,N_42026);
and U48428 (N_48428,N_43650,N_44884);
and U48429 (N_48429,N_42077,N_44024);
nor U48430 (N_48430,N_43702,N_42625);
nor U48431 (N_48431,N_43609,N_40555);
nand U48432 (N_48432,N_41205,N_43381);
or U48433 (N_48433,N_41344,N_42990);
and U48434 (N_48434,N_43365,N_43825);
xnor U48435 (N_48435,N_41549,N_43327);
nand U48436 (N_48436,N_42043,N_44765);
nor U48437 (N_48437,N_44151,N_41106);
nand U48438 (N_48438,N_42044,N_40726);
nor U48439 (N_48439,N_43430,N_40021);
nor U48440 (N_48440,N_44716,N_44316);
nand U48441 (N_48441,N_41816,N_40494);
xnor U48442 (N_48442,N_42988,N_44323);
nor U48443 (N_48443,N_43509,N_44265);
and U48444 (N_48444,N_42700,N_42784);
and U48445 (N_48445,N_40465,N_44530);
or U48446 (N_48446,N_42713,N_40525);
and U48447 (N_48447,N_44876,N_44763);
nor U48448 (N_48448,N_41012,N_44672);
nand U48449 (N_48449,N_42335,N_43044);
xor U48450 (N_48450,N_40101,N_42060);
or U48451 (N_48451,N_41690,N_40348);
nand U48452 (N_48452,N_42972,N_40847);
or U48453 (N_48453,N_43275,N_44500);
xor U48454 (N_48454,N_44268,N_40217);
xor U48455 (N_48455,N_42531,N_43028);
and U48456 (N_48456,N_41246,N_44774);
and U48457 (N_48457,N_42981,N_40128);
nand U48458 (N_48458,N_42293,N_44755);
xor U48459 (N_48459,N_43952,N_40903);
nor U48460 (N_48460,N_42726,N_43072);
nand U48461 (N_48461,N_44111,N_44866);
nand U48462 (N_48462,N_40976,N_42358);
and U48463 (N_48463,N_43566,N_43248);
nand U48464 (N_48464,N_40680,N_40059);
nand U48465 (N_48465,N_40517,N_41978);
xnor U48466 (N_48466,N_42181,N_41643);
nor U48467 (N_48467,N_41061,N_41382);
nand U48468 (N_48468,N_43946,N_43180);
xnor U48469 (N_48469,N_43503,N_40369);
xnor U48470 (N_48470,N_43383,N_40047);
nand U48471 (N_48471,N_42255,N_43194);
or U48472 (N_48472,N_40070,N_44994);
nor U48473 (N_48473,N_43936,N_41195);
nand U48474 (N_48474,N_43699,N_41655);
nand U48475 (N_48475,N_43252,N_43976);
nor U48476 (N_48476,N_43260,N_44735);
and U48477 (N_48477,N_40037,N_43265);
xnor U48478 (N_48478,N_44713,N_43095);
nor U48479 (N_48479,N_42196,N_41413);
xnor U48480 (N_48480,N_40734,N_44731);
xnor U48481 (N_48481,N_41669,N_43728);
and U48482 (N_48482,N_42962,N_40725);
nand U48483 (N_48483,N_40208,N_44336);
nand U48484 (N_48484,N_44526,N_44497);
and U48485 (N_48485,N_44024,N_42609);
or U48486 (N_48486,N_44257,N_44659);
or U48487 (N_48487,N_44287,N_44388);
xnor U48488 (N_48488,N_43536,N_43425);
xnor U48489 (N_48489,N_44138,N_43007);
or U48490 (N_48490,N_43267,N_40041);
and U48491 (N_48491,N_44697,N_42458);
nand U48492 (N_48492,N_41870,N_43936);
or U48493 (N_48493,N_40911,N_40766);
nor U48494 (N_48494,N_44100,N_42041);
nor U48495 (N_48495,N_44168,N_41314);
and U48496 (N_48496,N_43122,N_43521);
nor U48497 (N_48497,N_43570,N_43732);
nor U48498 (N_48498,N_41674,N_41042);
or U48499 (N_48499,N_44463,N_44061);
xor U48500 (N_48500,N_43632,N_43767);
nand U48501 (N_48501,N_43370,N_41294);
nor U48502 (N_48502,N_42419,N_43631);
nor U48503 (N_48503,N_44776,N_44299);
nor U48504 (N_48504,N_40687,N_42552);
xnor U48505 (N_48505,N_42089,N_43721);
nand U48506 (N_48506,N_44237,N_44530);
and U48507 (N_48507,N_43111,N_40325);
nand U48508 (N_48508,N_44161,N_43195);
and U48509 (N_48509,N_42948,N_42262);
nand U48510 (N_48510,N_44669,N_42027);
nand U48511 (N_48511,N_43072,N_41671);
xnor U48512 (N_48512,N_43792,N_44456);
nor U48513 (N_48513,N_42029,N_40716);
nor U48514 (N_48514,N_44052,N_40491);
nand U48515 (N_48515,N_40512,N_43459);
nor U48516 (N_48516,N_42448,N_41701);
xnor U48517 (N_48517,N_43676,N_40099);
nand U48518 (N_48518,N_43044,N_42887);
or U48519 (N_48519,N_42749,N_44327);
nand U48520 (N_48520,N_42563,N_43161);
nor U48521 (N_48521,N_43656,N_41069);
nor U48522 (N_48522,N_44365,N_44084);
xnor U48523 (N_48523,N_40017,N_42797);
xnor U48524 (N_48524,N_44977,N_44986);
xor U48525 (N_48525,N_42696,N_43647);
nand U48526 (N_48526,N_43743,N_44691);
xor U48527 (N_48527,N_41757,N_41520);
nor U48528 (N_48528,N_42990,N_40867);
or U48529 (N_48529,N_42458,N_41028);
xor U48530 (N_48530,N_42875,N_42895);
and U48531 (N_48531,N_41415,N_40135);
or U48532 (N_48532,N_42796,N_40206);
and U48533 (N_48533,N_43736,N_44913);
nor U48534 (N_48534,N_40126,N_42424);
xor U48535 (N_48535,N_43975,N_43065);
and U48536 (N_48536,N_41252,N_41487);
nor U48537 (N_48537,N_43756,N_44248);
nand U48538 (N_48538,N_43182,N_41875);
nand U48539 (N_48539,N_40772,N_40598);
nor U48540 (N_48540,N_40737,N_44887);
nor U48541 (N_48541,N_40339,N_41942);
nor U48542 (N_48542,N_40211,N_42649);
nor U48543 (N_48543,N_42662,N_40824);
xor U48544 (N_48544,N_41125,N_42539);
xor U48545 (N_48545,N_44069,N_44725);
or U48546 (N_48546,N_44459,N_40230);
or U48547 (N_48547,N_44282,N_41815);
nand U48548 (N_48548,N_43963,N_42831);
and U48549 (N_48549,N_44384,N_44734);
xor U48550 (N_48550,N_40381,N_40059);
or U48551 (N_48551,N_43278,N_42699);
and U48552 (N_48552,N_42293,N_44504);
and U48553 (N_48553,N_42294,N_40881);
nand U48554 (N_48554,N_44953,N_42600);
nand U48555 (N_48555,N_43680,N_42099);
or U48556 (N_48556,N_42077,N_42168);
xor U48557 (N_48557,N_44131,N_44114);
and U48558 (N_48558,N_42667,N_43510);
nor U48559 (N_48559,N_43360,N_42016);
or U48560 (N_48560,N_44574,N_42116);
nand U48561 (N_48561,N_41177,N_42528);
nor U48562 (N_48562,N_42079,N_43827);
and U48563 (N_48563,N_44654,N_41179);
and U48564 (N_48564,N_41851,N_41295);
nand U48565 (N_48565,N_42970,N_40734);
nor U48566 (N_48566,N_41953,N_44755);
xor U48567 (N_48567,N_41366,N_42720);
or U48568 (N_48568,N_41290,N_42128);
xor U48569 (N_48569,N_42346,N_43101);
and U48570 (N_48570,N_42286,N_44418);
or U48571 (N_48571,N_40761,N_40832);
xor U48572 (N_48572,N_43311,N_41524);
and U48573 (N_48573,N_42242,N_40537);
and U48574 (N_48574,N_43369,N_41568);
xnor U48575 (N_48575,N_44721,N_41861);
nand U48576 (N_48576,N_41301,N_40085);
or U48577 (N_48577,N_44193,N_44009);
xnor U48578 (N_48578,N_41347,N_42137);
nand U48579 (N_48579,N_42716,N_42544);
xor U48580 (N_48580,N_43986,N_41695);
and U48581 (N_48581,N_41691,N_40898);
or U48582 (N_48582,N_43755,N_40966);
xor U48583 (N_48583,N_42802,N_44365);
nor U48584 (N_48584,N_41980,N_44479);
xnor U48585 (N_48585,N_41342,N_44838);
or U48586 (N_48586,N_44936,N_43617);
nor U48587 (N_48587,N_40592,N_40229);
or U48588 (N_48588,N_42036,N_44435);
or U48589 (N_48589,N_43418,N_42871);
or U48590 (N_48590,N_41626,N_43104);
and U48591 (N_48591,N_40758,N_44633);
and U48592 (N_48592,N_44105,N_44372);
xor U48593 (N_48593,N_42256,N_42304);
xor U48594 (N_48594,N_43071,N_40346);
nor U48595 (N_48595,N_42534,N_43830);
nand U48596 (N_48596,N_44577,N_41280);
and U48597 (N_48597,N_40822,N_43633);
nor U48598 (N_48598,N_41190,N_43486);
and U48599 (N_48599,N_43744,N_41256);
and U48600 (N_48600,N_44171,N_43400);
nor U48601 (N_48601,N_40753,N_41716);
xnor U48602 (N_48602,N_41494,N_40464);
xor U48603 (N_48603,N_42624,N_43689);
or U48604 (N_48604,N_42278,N_42747);
nor U48605 (N_48605,N_43101,N_43369);
or U48606 (N_48606,N_43311,N_42581);
xor U48607 (N_48607,N_44970,N_40670);
xnor U48608 (N_48608,N_43551,N_44871);
or U48609 (N_48609,N_41725,N_44249);
nor U48610 (N_48610,N_41229,N_41712);
and U48611 (N_48611,N_42240,N_43263);
nor U48612 (N_48612,N_41036,N_41955);
nand U48613 (N_48613,N_43126,N_40523);
nor U48614 (N_48614,N_41719,N_44422);
or U48615 (N_48615,N_41106,N_40687);
xor U48616 (N_48616,N_41023,N_43814);
nand U48617 (N_48617,N_44812,N_44069);
nand U48618 (N_48618,N_41743,N_42719);
xor U48619 (N_48619,N_42650,N_40410);
and U48620 (N_48620,N_40555,N_40646);
xnor U48621 (N_48621,N_42213,N_43572);
nand U48622 (N_48622,N_42691,N_41370);
xor U48623 (N_48623,N_40470,N_41970);
and U48624 (N_48624,N_41130,N_44617);
nand U48625 (N_48625,N_40821,N_43350);
nor U48626 (N_48626,N_41180,N_44063);
nand U48627 (N_48627,N_42804,N_42830);
nand U48628 (N_48628,N_41024,N_41310);
xnor U48629 (N_48629,N_40608,N_40026);
or U48630 (N_48630,N_42937,N_43304);
or U48631 (N_48631,N_40371,N_43152);
nor U48632 (N_48632,N_43668,N_41499);
nand U48633 (N_48633,N_43541,N_44300);
xnor U48634 (N_48634,N_42456,N_41959);
or U48635 (N_48635,N_42225,N_40269);
nor U48636 (N_48636,N_41390,N_41235);
nand U48637 (N_48637,N_44718,N_42868);
or U48638 (N_48638,N_42783,N_42342);
xor U48639 (N_48639,N_44579,N_41672);
or U48640 (N_48640,N_40577,N_40558);
nor U48641 (N_48641,N_43339,N_42656);
and U48642 (N_48642,N_42107,N_40022);
or U48643 (N_48643,N_43488,N_41914);
nand U48644 (N_48644,N_44809,N_43211);
xnor U48645 (N_48645,N_42463,N_41716);
xnor U48646 (N_48646,N_42622,N_41697);
xnor U48647 (N_48647,N_42273,N_40601);
and U48648 (N_48648,N_42778,N_41186);
nand U48649 (N_48649,N_41831,N_41424);
nor U48650 (N_48650,N_44930,N_43164);
or U48651 (N_48651,N_40920,N_42427);
nor U48652 (N_48652,N_43731,N_44769);
or U48653 (N_48653,N_44972,N_44770);
xor U48654 (N_48654,N_44859,N_44622);
nand U48655 (N_48655,N_44135,N_42217);
xnor U48656 (N_48656,N_40937,N_41668);
and U48657 (N_48657,N_42285,N_42704);
and U48658 (N_48658,N_43976,N_42439);
nand U48659 (N_48659,N_44152,N_43682);
or U48660 (N_48660,N_40176,N_41102);
or U48661 (N_48661,N_42746,N_44854);
xor U48662 (N_48662,N_43494,N_42655);
nand U48663 (N_48663,N_41820,N_44689);
or U48664 (N_48664,N_41425,N_42167);
and U48665 (N_48665,N_43512,N_42375);
nand U48666 (N_48666,N_41816,N_41743);
nor U48667 (N_48667,N_40319,N_44363);
or U48668 (N_48668,N_41514,N_41382);
xor U48669 (N_48669,N_44605,N_41440);
xor U48670 (N_48670,N_43554,N_44069);
and U48671 (N_48671,N_41938,N_43313);
nand U48672 (N_48672,N_42432,N_44899);
nand U48673 (N_48673,N_41029,N_43954);
or U48674 (N_48674,N_41685,N_43614);
nand U48675 (N_48675,N_42910,N_41522);
or U48676 (N_48676,N_41748,N_42177);
or U48677 (N_48677,N_42362,N_40165);
nor U48678 (N_48678,N_43733,N_42884);
and U48679 (N_48679,N_41048,N_42960);
xnor U48680 (N_48680,N_43754,N_41718);
nand U48681 (N_48681,N_43957,N_43247);
and U48682 (N_48682,N_40145,N_44578);
xnor U48683 (N_48683,N_42629,N_40144);
xnor U48684 (N_48684,N_42369,N_44272);
xnor U48685 (N_48685,N_41427,N_44457);
or U48686 (N_48686,N_42890,N_44355);
and U48687 (N_48687,N_42474,N_42065);
and U48688 (N_48688,N_44799,N_42994);
or U48689 (N_48689,N_40201,N_40147);
and U48690 (N_48690,N_43841,N_40525);
or U48691 (N_48691,N_42239,N_44505);
nor U48692 (N_48692,N_42695,N_41429);
xor U48693 (N_48693,N_44344,N_43375);
or U48694 (N_48694,N_44234,N_40250);
nor U48695 (N_48695,N_42506,N_41156);
xnor U48696 (N_48696,N_41601,N_42285);
nor U48697 (N_48697,N_43554,N_42230);
xor U48698 (N_48698,N_44165,N_44541);
xor U48699 (N_48699,N_41810,N_42311);
or U48700 (N_48700,N_40280,N_40407);
nor U48701 (N_48701,N_40207,N_42132);
and U48702 (N_48702,N_44018,N_41837);
nor U48703 (N_48703,N_43617,N_42643);
or U48704 (N_48704,N_40490,N_41622);
nand U48705 (N_48705,N_43119,N_40845);
xor U48706 (N_48706,N_43184,N_44361);
xnor U48707 (N_48707,N_41505,N_40687);
and U48708 (N_48708,N_43904,N_40392);
or U48709 (N_48709,N_40629,N_44053);
nand U48710 (N_48710,N_44532,N_41159);
and U48711 (N_48711,N_44722,N_42086);
nor U48712 (N_48712,N_40542,N_41030);
and U48713 (N_48713,N_41213,N_40821);
and U48714 (N_48714,N_40417,N_40358);
and U48715 (N_48715,N_44439,N_40946);
and U48716 (N_48716,N_44681,N_41873);
and U48717 (N_48717,N_41066,N_44474);
and U48718 (N_48718,N_44436,N_43731);
xnor U48719 (N_48719,N_42843,N_40363);
or U48720 (N_48720,N_42559,N_42631);
or U48721 (N_48721,N_40165,N_43199);
and U48722 (N_48722,N_41057,N_43879);
or U48723 (N_48723,N_44724,N_42329);
and U48724 (N_48724,N_41552,N_43811);
or U48725 (N_48725,N_41893,N_40822);
and U48726 (N_48726,N_43220,N_40039);
xnor U48727 (N_48727,N_43558,N_43769);
or U48728 (N_48728,N_40419,N_42783);
xnor U48729 (N_48729,N_42425,N_41051);
or U48730 (N_48730,N_42312,N_41518);
and U48731 (N_48731,N_42325,N_43305);
xnor U48732 (N_48732,N_40091,N_44310);
nand U48733 (N_48733,N_42978,N_40503);
or U48734 (N_48734,N_42403,N_42831);
nor U48735 (N_48735,N_43763,N_40907);
xnor U48736 (N_48736,N_40681,N_44933);
or U48737 (N_48737,N_42757,N_44034);
nor U48738 (N_48738,N_43957,N_44456);
nor U48739 (N_48739,N_42886,N_42719);
nand U48740 (N_48740,N_44403,N_42698);
or U48741 (N_48741,N_40679,N_44426);
nor U48742 (N_48742,N_40124,N_41025);
xor U48743 (N_48743,N_42271,N_42048);
and U48744 (N_48744,N_42330,N_41427);
or U48745 (N_48745,N_44802,N_40040);
nand U48746 (N_48746,N_42268,N_44329);
nand U48747 (N_48747,N_41569,N_40165);
nor U48748 (N_48748,N_41580,N_41759);
nor U48749 (N_48749,N_44131,N_44940);
and U48750 (N_48750,N_40934,N_43045);
and U48751 (N_48751,N_41711,N_42571);
xor U48752 (N_48752,N_43339,N_43242);
nand U48753 (N_48753,N_44123,N_41075);
and U48754 (N_48754,N_42351,N_40070);
xnor U48755 (N_48755,N_42080,N_43490);
or U48756 (N_48756,N_43996,N_40439);
or U48757 (N_48757,N_41705,N_42870);
or U48758 (N_48758,N_42667,N_40940);
nand U48759 (N_48759,N_42241,N_41826);
and U48760 (N_48760,N_43723,N_43541);
and U48761 (N_48761,N_41600,N_43445);
or U48762 (N_48762,N_44577,N_41622);
nand U48763 (N_48763,N_40344,N_41788);
and U48764 (N_48764,N_40961,N_42618);
or U48765 (N_48765,N_43732,N_43798);
or U48766 (N_48766,N_40511,N_42324);
and U48767 (N_48767,N_42916,N_40901);
nand U48768 (N_48768,N_42088,N_44071);
nand U48769 (N_48769,N_41591,N_43476);
xor U48770 (N_48770,N_40171,N_42756);
and U48771 (N_48771,N_40567,N_43409);
xnor U48772 (N_48772,N_40914,N_40793);
nand U48773 (N_48773,N_43255,N_43489);
nor U48774 (N_48774,N_40119,N_44673);
xnor U48775 (N_48775,N_40632,N_44300);
nand U48776 (N_48776,N_42037,N_41064);
nand U48777 (N_48777,N_44797,N_41752);
nand U48778 (N_48778,N_43877,N_41980);
nand U48779 (N_48779,N_42465,N_41853);
xnor U48780 (N_48780,N_44571,N_41373);
and U48781 (N_48781,N_43359,N_40847);
or U48782 (N_48782,N_43189,N_43903);
and U48783 (N_48783,N_40718,N_43871);
or U48784 (N_48784,N_41789,N_40107);
or U48785 (N_48785,N_44611,N_40622);
or U48786 (N_48786,N_40421,N_40250);
nand U48787 (N_48787,N_44155,N_43094);
nand U48788 (N_48788,N_44942,N_41126);
xnor U48789 (N_48789,N_41484,N_44734);
or U48790 (N_48790,N_42288,N_42971);
or U48791 (N_48791,N_40696,N_42556);
nand U48792 (N_48792,N_43012,N_40403);
or U48793 (N_48793,N_42784,N_44268);
nor U48794 (N_48794,N_42215,N_44542);
nor U48795 (N_48795,N_44926,N_43254);
nand U48796 (N_48796,N_43617,N_42036);
nand U48797 (N_48797,N_44359,N_43881);
and U48798 (N_48798,N_40144,N_41323);
and U48799 (N_48799,N_40785,N_42828);
and U48800 (N_48800,N_43419,N_41316);
nand U48801 (N_48801,N_44237,N_44388);
nand U48802 (N_48802,N_40122,N_43674);
nand U48803 (N_48803,N_42401,N_40801);
nand U48804 (N_48804,N_43635,N_40874);
or U48805 (N_48805,N_40300,N_41308);
xnor U48806 (N_48806,N_41023,N_43452);
xnor U48807 (N_48807,N_43221,N_40506);
nand U48808 (N_48808,N_42784,N_42251);
and U48809 (N_48809,N_41221,N_42503);
nand U48810 (N_48810,N_41618,N_42467);
nand U48811 (N_48811,N_44544,N_44403);
or U48812 (N_48812,N_43556,N_44801);
nand U48813 (N_48813,N_41066,N_40849);
nand U48814 (N_48814,N_41235,N_42046);
xor U48815 (N_48815,N_43828,N_44661);
nor U48816 (N_48816,N_41385,N_41336);
nor U48817 (N_48817,N_44173,N_42021);
nand U48818 (N_48818,N_41705,N_41249);
and U48819 (N_48819,N_44671,N_42898);
nand U48820 (N_48820,N_40322,N_43766);
xor U48821 (N_48821,N_44232,N_40348);
xnor U48822 (N_48822,N_44493,N_44156);
nand U48823 (N_48823,N_40228,N_41802);
nor U48824 (N_48824,N_42532,N_43556);
nor U48825 (N_48825,N_43222,N_42739);
and U48826 (N_48826,N_43902,N_40111);
or U48827 (N_48827,N_44748,N_44115);
nand U48828 (N_48828,N_41020,N_44459);
nand U48829 (N_48829,N_44149,N_42019);
nor U48830 (N_48830,N_42245,N_44464);
and U48831 (N_48831,N_42206,N_44067);
or U48832 (N_48832,N_41027,N_42597);
nand U48833 (N_48833,N_43111,N_42565);
nor U48834 (N_48834,N_43997,N_42320);
nand U48835 (N_48835,N_40164,N_41806);
nand U48836 (N_48836,N_40293,N_42180);
nor U48837 (N_48837,N_43134,N_40286);
nand U48838 (N_48838,N_41849,N_41907);
nor U48839 (N_48839,N_42532,N_40892);
or U48840 (N_48840,N_40268,N_40346);
nand U48841 (N_48841,N_42746,N_42182);
or U48842 (N_48842,N_42394,N_43202);
or U48843 (N_48843,N_43399,N_40644);
nand U48844 (N_48844,N_44996,N_42525);
or U48845 (N_48845,N_40572,N_44207);
or U48846 (N_48846,N_43644,N_40283);
nor U48847 (N_48847,N_41402,N_42845);
nor U48848 (N_48848,N_40939,N_42811);
and U48849 (N_48849,N_44705,N_42259);
nand U48850 (N_48850,N_42393,N_41565);
nand U48851 (N_48851,N_44575,N_44676);
or U48852 (N_48852,N_40249,N_44419);
nor U48853 (N_48853,N_40771,N_44646);
xnor U48854 (N_48854,N_41868,N_40107);
nor U48855 (N_48855,N_40545,N_42128);
nor U48856 (N_48856,N_40662,N_44262);
nor U48857 (N_48857,N_43894,N_42539);
and U48858 (N_48858,N_43043,N_44062);
nand U48859 (N_48859,N_44499,N_41955);
xnor U48860 (N_48860,N_40741,N_42867);
nand U48861 (N_48861,N_44401,N_44877);
nand U48862 (N_48862,N_41390,N_44905);
nor U48863 (N_48863,N_41757,N_44031);
xnor U48864 (N_48864,N_40933,N_43742);
nand U48865 (N_48865,N_40262,N_43745);
or U48866 (N_48866,N_43813,N_44741);
xnor U48867 (N_48867,N_41234,N_42020);
nand U48868 (N_48868,N_44032,N_44909);
nor U48869 (N_48869,N_40978,N_43447);
nor U48870 (N_48870,N_43899,N_44925);
nor U48871 (N_48871,N_44902,N_41942);
nand U48872 (N_48872,N_42655,N_44775);
nor U48873 (N_48873,N_43965,N_41397);
nor U48874 (N_48874,N_40850,N_41296);
nand U48875 (N_48875,N_44388,N_44365);
nand U48876 (N_48876,N_41093,N_43814);
and U48877 (N_48877,N_44995,N_40936);
or U48878 (N_48878,N_43401,N_44951);
or U48879 (N_48879,N_40296,N_42843);
nand U48880 (N_48880,N_43786,N_43592);
or U48881 (N_48881,N_42889,N_41503);
or U48882 (N_48882,N_42832,N_41104);
xor U48883 (N_48883,N_42908,N_42695);
or U48884 (N_48884,N_42559,N_41117);
xor U48885 (N_48885,N_43919,N_42135);
nor U48886 (N_48886,N_43898,N_42316);
xor U48887 (N_48887,N_41958,N_43459);
nand U48888 (N_48888,N_40016,N_41255);
nor U48889 (N_48889,N_41019,N_41364);
nand U48890 (N_48890,N_41398,N_42069);
xor U48891 (N_48891,N_42933,N_40464);
xor U48892 (N_48892,N_42939,N_41293);
or U48893 (N_48893,N_41389,N_42855);
or U48894 (N_48894,N_44201,N_44624);
xnor U48895 (N_48895,N_41827,N_41657);
and U48896 (N_48896,N_42495,N_44018);
or U48897 (N_48897,N_43720,N_43938);
nand U48898 (N_48898,N_44058,N_42641);
nor U48899 (N_48899,N_42833,N_43840);
xor U48900 (N_48900,N_41976,N_44532);
or U48901 (N_48901,N_43870,N_40261);
and U48902 (N_48902,N_42032,N_43981);
and U48903 (N_48903,N_43723,N_43305);
or U48904 (N_48904,N_40529,N_40445);
xnor U48905 (N_48905,N_43574,N_40074);
and U48906 (N_48906,N_41735,N_41205);
xnor U48907 (N_48907,N_41605,N_44944);
nor U48908 (N_48908,N_41714,N_43708);
nor U48909 (N_48909,N_42544,N_44918);
xor U48910 (N_48910,N_41510,N_40623);
xor U48911 (N_48911,N_40770,N_44529);
xor U48912 (N_48912,N_44863,N_41407);
nor U48913 (N_48913,N_42231,N_41219);
nand U48914 (N_48914,N_43870,N_41864);
nor U48915 (N_48915,N_40122,N_41037);
xnor U48916 (N_48916,N_43291,N_43167);
nor U48917 (N_48917,N_41677,N_40732);
or U48918 (N_48918,N_42054,N_43019);
xnor U48919 (N_48919,N_41127,N_43537);
xor U48920 (N_48920,N_40963,N_44180);
and U48921 (N_48921,N_44110,N_42263);
xnor U48922 (N_48922,N_44367,N_43155);
or U48923 (N_48923,N_41808,N_42241);
xor U48924 (N_48924,N_40729,N_43508);
nand U48925 (N_48925,N_40842,N_43593);
nand U48926 (N_48926,N_43560,N_42995);
xnor U48927 (N_48927,N_41674,N_41433);
and U48928 (N_48928,N_44360,N_42559);
nor U48929 (N_48929,N_40806,N_41260);
nand U48930 (N_48930,N_43684,N_44068);
xnor U48931 (N_48931,N_41742,N_40386);
or U48932 (N_48932,N_40810,N_43145);
nor U48933 (N_48933,N_41431,N_42397);
nand U48934 (N_48934,N_42669,N_43420);
nand U48935 (N_48935,N_43199,N_43126);
and U48936 (N_48936,N_43276,N_42179);
nor U48937 (N_48937,N_43073,N_44243);
and U48938 (N_48938,N_42170,N_42120);
xnor U48939 (N_48939,N_40222,N_40326);
xor U48940 (N_48940,N_41991,N_42327);
nor U48941 (N_48941,N_41287,N_43008);
and U48942 (N_48942,N_42162,N_41167);
or U48943 (N_48943,N_43350,N_40757);
nor U48944 (N_48944,N_41596,N_44156);
nor U48945 (N_48945,N_42202,N_42065);
and U48946 (N_48946,N_44861,N_41613);
and U48947 (N_48947,N_41947,N_42939);
nand U48948 (N_48948,N_44708,N_43186);
nand U48949 (N_48949,N_41252,N_44363);
or U48950 (N_48950,N_42040,N_41021);
or U48951 (N_48951,N_40138,N_42963);
or U48952 (N_48952,N_42143,N_41169);
or U48953 (N_48953,N_41125,N_44040);
or U48954 (N_48954,N_41508,N_40541);
xor U48955 (N_48955,N_43224,N_40439);
xnor U48956 (N_48956,N_40107,N_40752);
or U48957 (N_48957,N_43080,N_44992);
and U48958 (N_48958,N_41950,N_41685);
and U48959 (N_48959,N_44368,N_40565);
nor U48960 (N_48960,N_41953,N_43529);
xnor U48961 (N_48961,N_40168,N_41257);
nor U48962 (N_48962,N_42762,N_40835);
nor U48963 (N_48963,N_44088,N_41374);
nand U48964 (N_48964,N_44648,N_40168);
or U48965 (N_48965,N_42544,N_43122);
and U48966 (N_48966,N_42316,N_42439);
nor U48967 (N_48967,N_44008,N_43274);
nand U48968 (N_48968,N_43739,N_42202);
or U48969 (N_48969,N_41921,N_44116);
xnor U48970 (N_48970,N_41215,N_40743);
or U48971 (N_48971,N_42144,N_41845);
xor U48972 (N_48972,N_40727,N_41827);
xnor U48973 (N_48973,N_44560,N_41766);
and U48974 (N_48974,N_42874,N_43537);
or U48975 (N_48975,N_41870,N_44219);
or U48976 (N_48976,N_42120,N_40778);
nor U48977 (N_48977,N_43443,N_40348);
nand U48978 (N_48978,N_44553,N_44040);
and U48979 (N_48979,N_40370,N_43707);
xor U48980 (N_48980,N_43482,N_41856);
and U48981 (N_48981,N_42515,N_40933);
xor U48982 (N_48982,N_42429,N_40794);
and U48983 (N_48983,N_43829,N_40080);
nor U48984 (N_48984,N_44483,N_42291);
nand U48985 (N_48985,N_42274,N_40581);
xor U48986 (N_48986,N_44758,N_41383);
and U48987 (N_48987,N_41982,N_43411);
nor U48988 (N_48988,N_42899,N_40391);
or U48989 (N_48989,N_44865,N_43100);
and U48990 (N_48990,N_41613,N_43414);
or U48991 (N_48991,N_40819,N_44853);
and U48992 (N_48992,N_41161,N_43303);
xnor U48993 (N_48993,N_40726,N_43815);
and U48994 (N_48994,N_44439,N_43839);
or U48995 (N_48995,N_42060,N_42264);
nand U48996 (N_48996,N_44282,N_43470);
and U48997 (N_48997,N_41012,N_40302);
nor U48998 (N_48998,N_40362,N_40500);
nand U48999 (N_48999,N_42065,N_42660);
xnor U49000 (N_49000,N_44634,N_40524);
nor U49001 (N_49001,N_40159,N_42053);
nand U49002 (N_49002,N_40475,N_43727);
or U49003 (N_49003,N_43508,N_43323);
xor U49004 (N_49004,N_43071,N_42760);
xnor U49005 (N_49005,N_40192,N_43607);
or U49006 (N_49006,N_40702,N_44538);
nor U49007 (N_49007,N_40028,N_44145);
or U49008 (N_49008,N_44637,N_41310);
xor U49009 (N_49009,N_43739,N_44058);
and U49010 (N_49010,N_40550,N_42276);
nand U49011 (N_49011,N_44194,N_44021);
xor U49012 (N_49012,N_42423,N_43216);
nor U49013 (N_49013,N_40908,N_43418);
nand U49014 (N_49014,N_41245,N_40650);
xor U49015 (N_49015,N_41724,N_40374);
or U49016 (N_49016,N_40797,N_42858);
nand U49017 (N_49017,N_40315,N_42687);
nor U49018 (N_49018,N_44946,N_44221);
nand U49019 (N_49019,N_41973,N_40236);
and U49020 (N_49020,N_40528,N_41750);
nor U49021 (N_49021,N_43847,N_41440);
or U49022 (N_49022,N_42764,N_44219);
xor U49023 (N_49023,N_42293,N_43755);
and U49024 (N_49024,N_43543,N_44500);
nand U49025 (N_49025,N_44639,N_42359);
and U49026 (N_49026,N_43689,N_43600);
xnor U49027 (N_49027,N_40162,N_42017);
nand U49028 (N_49028,N_43029,N_40601);
and U49029 (N_49029,N_43762,N_42593);
and U49030 (N_49030,N_44674,N_42093);
xnor U49031 (N_49031,N_41612,N_40706);
nand U49032 (N_49032,N_41146,N_41963);
or U49033 (N_49033,N_41119,N_41423);
nor U49034 (N_49034,N_44239,N_42997);
nand U49035 (N_49035,N_43656,N_40467);
nor U49036 (N_49036,N_40327,N_41509);
and U49037 (N_49037,N_42370,N_42389);
nand U49038 (N_49038,N_43264,N_43082);
and U49039 (N_49039,N_44351,N_43966);
or U49040 (N_49040,N_41837,N_40373);
nor U49041 (N_49041,N_40716,N_40093);
or U49042 (N_49042,N_40191,N_42605);
and U49043 (N_49043,N_44818,N_43139);
nor U49044 (N_49044,N_44570,N_42413);
xnor U49045 (N_49045,N_41735,N_44065);
nand U49046 (N_49046,N_44976,N_44582);
and U49047 (N_49047,N_43596,N_40185);
and U49048 (N_49048,N_41366,N_42637);
nand U49049 (N_49049,N_44466,N_42062);
nand U49050 (N_49050,N_42629,N_42045);
and U49051 (N_49051,N_40670,N_43919);
xnor U49052 (N_49052,N_43678,N_42375);
nand U49053 (N_49053,N_42130,N_40825);
nor U49054 (N_49054,N_41936,N_44035);
or U49055 (N_49055,N_41299,N_44420);
or U49056 (N_49056,N_43640,N_42536);
nor U49057 (N_49057,N_43390,N_41857);
nand U49058 (N_49058,N_42502,N_41170);
xor U49059 (N_49059,N_41637,N_44949);
nand U49060 (N_49060,N_42034,N_42284);
and U49061 (N_49061,N_43712,N_42547);
or U49062 (N_49062,N_44005,N_44750);
nor U49063 (N_49063,N_44184,N_41373);
nand U49064 (N_49064,N_43969,N_42784);
and U49065 (N_49065,N_42748,N_40183);
or U49066 (N_49066,N_44607,N_41034);
and U49067 (N_49067,N_41989,N_43305);
nor U49068 (N_49068,N_44763,N_40128);
nor U49069 (N_49069,N_43291,N_42607);
and U49070 (N_49070,N_41477,N_41352);
xor U49071 (N_49071,N_40135,N_43185);
nand U49072 (N_49072,N_43898,N_41854);
nand U49073 (N_49073,N_43379,N_43688);
and U49074 (N_49074,N_43524,N_43456);
nand U49075 (N_49075,N_40592,N_44013);
and U49076 (N_49076,N_40518,N_41706);
nand U49077 (N_49077,N_41442,N_40835);
or U49078 (N_49078,N_43802,N_43624);
nor U49079 (N_49079,N_41253,N_44507);
xor U49080 (N_49080,N_41811,N_41771);
nand U49081 (N_49081,N_44425,N_43925);
nand U49082 (N_49082,N_40357,N_44693);
nor U49083 (N_49083,N_44804,N_40584);
xnor U49084 (N_49084,N_41988,N_42999);
xor U49085 (N_49085,N_41128,N_44268);
xnor U49086 (N_49086,N_44999,N_41465);
nand U49087 (N_49087,N_44412,N_40251);
nor U49088 (N_49088,N_40645,N_44850);
xnor U49089 (N_49089,N_44105,N_44687);
xnor U49090 (N_49090,N_44640,N_41211);
nand U49091 (N_49091,N_43912,N_42469);
and U49092 (N_49092,N_40173,N_44729);
nand U49093 (N_49093,N_44287,N_42816);
nor U49094 (N_49094,N_43165,N_42302);
xnor U49095 (N_49095,N_43832,N_40353);
nor U49096 (N_49096,N_41552,N_43283);
and U49097 (N_49097,N_42134,N_44815);
nand U49098 (N_49098,N_43638,N_42041);
nand U49099 (N_49099,N_42640,N_44127);
xor U49100 (N_49100,N_42233,N_40656);
or U49101 (N_49101,N_44749,N_43853);
nand U49102 (N_49102,N_40888,N_44557);
or U49103 (N_49103,N_43863,N_40720);
nor U49104 (N_49104,N_44547,N_40428);
or U49105 (N_49105,N_44127,N_41746);
and U49106 (N_49106,N_40374,N_40825);
and U49107 (N_49107,N_43930,N_41588);
and U49108 (N_49108,N_42334,N_40838);
and U49109 (N_49109,N_41431,N_42629);
or U49110 (N_49110,N_44637,N_41990);
and U49111 (N_49111,N_42061,N_44336);
and U49112 (N_49112,N_44554,N_41701);
and U49113 (N_49113,N_44058,N_40401);
or U49114 (N_49114,N_43012,N_43996);
nor U49115 (N_49115,N_43051,N_40205);
nand U49116 (N_49116,N_44048,N_44648);
or U49117 (N_49117,N_44784,N_41509);
nand U49118 (N_49118,N_41816,N_41065);
or U49119 (N_49119,N_41309,N_44826);
xnor U49120 (N_49120,N_43774,N_42040);
xnor U49121 (N_49121,N_43367,N_42503);
or U49122 (N_49122,N_44712,N_40285);
and U49123 (N_49123,N_44552,N_44852);
nand U49124 (N_49124,N_41640,N_41729);
nand U49125 (N_49125,N_40076,N_41563);
and U49126 (N_49126,N_44043,N_40022);
nand U49127 (N_49127,N_42401,N_43829);
and U49128 (N_49128,N_44895,N_41659);
nor U49129 (N_49129,N_44163,N_40202);
xor U49130 (N_49130,N_41355,N_42545);
xor U49131 (N_49131,N_42633,N_43532);
xor U49132 (N_49132,N_44007,N_41307);
or U49133 (N_49133,N_43712,N_40321);
xnor U49134 (N_49134,N_44347,N_42601);
nand U49135 (N_49135,N_43104,N_43171);
nor U49136 (N_49136,N_43951,N_42879);
or U49137 (N_49137,N_43071,N_42731);
or U49138 (N_49138,N_42145,N_44052);
nor U49139 (N_49139,N_42715,N_43314);
or U49140 (N_49140,N_44418,N_40496);
xnor U49141 (N_49141,N_42423,N_41580);
nand U49142 (N_49142,N_41971,N_41557);
nand U49143 (N_49143,N_43741,N_42842);
or U49144 (N_49144,N_43034,N_43455);
and U49145 (N_49145,N_40041,N_43089);
nor U49146 (N_49146,N_41925,N_44697);
nor U49147 (N_49147,N_40485,N_41229);
and U49148 (N_49148,N_41378,N_44726);
or U49149 (N_49149,N_41353,N_41445);
and U49150 (N_49150,N_44407,N_40447);
nor U49151 (N_49151,N_41125,N_40204);
xor U49152 (N_49152,N_43085,N_44270);
nand U49153 (N_49153,N_40281,N_43064);
and U49154 (N_49154,N_41514,N_41571);
or U49155 (N_49155,N_41349,N_43783);
nor U49156 (N_49156,N_44295,N_42058);
nor U49157 (N_49157,N_42695,N_44079);
or U49158 (N_49158,N_43361,N_44829);
nor U49159 (N_49159,N_44768,N_40171);
or U49160 (N_49160,N_41485,N_44061);
and U49161 (N_49161,N_41976,N_42614);
nor U49162 (N_49162,N_41747,N_42932);
nor U49163 (N_49163,N_40058,N_42141);
or U49164 (N_49164,N_42889,N_43929);
nor U49165 (N_49165,N_40896,N_44793);
nor U49166 (N_49166,N_42125,N_41717);
nand U49167 (N_49167,N_42709,N_44619);
or U49168 (N_49168,N_42249,N_42298);
and U49169 (N_49169,N_43791,N_43488);
nand U49170 (N_49170,N_43548,N_44240);
nand U49171 (N_49171,N_44331,N_42969);
or U49172 (N_49172,N_43889,N_43397);
nor U49173 (N_49173,N_42047,N_42890);
xor U49174 (N_49174,N_44572,N_42014);
nand U49175 (N_49175,N_43034,N_44304);
nor U49176 (N_49176,N_42150,N_40476);
nor U49177 (N_49177,N_40912,N_43886);
nor U49178 (N_49178,N_43181,N_41916);
or U49179 (N_49179,N_42050,N_43684);
nor U49180 (N_49180,N_42101,N_44879);
xnor U49181 (N_49181,N_41477,N_43235);
nand U49182 (N_49182,N_42355,N_42332);
nand U49183 (N_49183,N_44798,N_43224);
xnor U49184 (N_49184,N_41135,N_41082);
and U49185 (N_49185,N_42606,N_43850);
and U49186 (N_49186,N_44419,N_43433);
or U49187 (N_49187,N_44213,N_40396);
nor U49188 (N_49188,N_40682,N_40626);
xor U49189 (N_49189,N_44142,N_41389);
nand U49190 (N_49190,N_42883,N_42751);
nand U49191 (N_49191,N_44857,N_43438);
and U49192 (N_49192,N_44767,N_42028);
and U49193 (N_49193,N_40124,N_42298);
and U49194 (N_49194,N_42810,N_43839);
and U49195 (N_49195,N_41820,N_40531);
xnor U49196 (N_49196,N_43745,N_43067);
xnor U49197 (N_49197,N_40246,N_44544);
and U49198 (N_49198,N_43010,N_44193);
nand U49199 (N_49199,N_44207,N_43939);
nor U49200 (N_49200,N_43674,N_42720);
nand U49201 (N_49201,N_43864,N_41220);
or U49202 (N_49202,N_43059,N_43209);
xnor U49203 (N_49203,N_40160,N_41859);
and U49204 (N_49204,N_44340,N_44840);
and U49205 (N_49205,N_43668,N_43972);
nand U49206 (N_49206,N_40503,N_43131);
nand U49207 (N_49207,N_44326,N_41702);
xor U49208 (N_49208,N_43415,N_44185);
nand U49209 (N_49209,N_40150,N_41568);
and U49210 (N_49210,N_41040,N_43452);
or U49211 (N_49211,N_42676,N_41224);
or U49212 (N_49212,N_42675,N_43069);
nand U49213 (N_49213,N_41812,N_41116);
xnor U49214 (N_49214,N_42809,N_42296);
and U49215 (N_49215,N_41467,N_43109);
or U49216 (N_49216,N_43968,N_43314);
nand U49217 (N_49217,N_42028,N_41355);
nand U49218 (N_49218,N_42752,N_43884);
and U49219 (N_49219,N_41835,N_44679);
nand U49220 (N_49220,N_40593,N_42276);
or U49221 (N_49221,N_41049,N_44194);
or U49222 (N_49222,N_40009,N_42389);
or U49223 (N_49223,N_42021,N_40931);
xnor U49224 (N_49224,N_41089,N_43849);
nor U49225 (N_49225,N_41095,N_43759);
nor U49226 (N_49226,N_43207,N_42829);
nand U49227 (N_49227,N_43380,N_43227);
xnor U49228 (N_49228,N_42112,N_43189);
nor U49229 (N_49229,N_40002,N_44118);
and U49230 (N_49230,N_42040,N_42933);
xnor U49231 (N_49231,N_43477,N_40549);
or U49232 (N_49232,N_44559,N_44958);
xnor U49233 (N_49233,N_44300,N_42285);
and U49234 (N_49234,N_42807,N_42623);
or U49235 (N_49235,N_40264,N_42762);
xor U49236 (N_49236,N_40619,N_43906);
nand U49237 (N_49237,N_42749,N_40873);
nand U49238 (N_49238,N_43558,N_43126);
nor U49239 (N_49239,N_42581,N_43490);
and U49240 (N_49240,N_43598,N_40178);
and U49241 (N_49241,N_41945,N_40306);
or U49242 (N_49242,N_44341,N_40561);
or U49243 (N_49243,N_41648,N_43507);
xnor U49244 (N_49244,N_41808,N_40752);
or U49245 (N_49245,N_40459,N_42376);
xor U49246 (N_49246,N_42264,N_44041);
or U49247 (N_49247,N_42765,N_42492);
and U49248 (N_49248,N_41927,N_44130);
xnor U49249 (N_49249,N_44692,N_41044);
nor U49250 (N_49250,N_40681,N_43658);
nor U49251 (N_49251,N_40635,N_43266);
or U49252 (N_49252,N_41009,N_42819);
nor U49253 (N_49253,N_40216,N_42512);
or U49254 (N_49254,N_42357,N_40583);
xnor U49255 (N_49255,N_44301,N_44708);
nand U49256 (N_49256,N_44002,N_41728);
or U49257 (N_49257,N_43803,N_40560);
and U49258 (N_49258,N_43945,N_42845);
and U49259 (N_49259,N_42197,N_40688);
and U49260 (N_49260,N_44401,N_44185);
nand U49261 (N_49261,N_44980,N_42357);
xnor U49262 (N_49262,N_42675,N_40783);
nand U49263 (N_49263,N_43763,N_42194);
or U49264 (N_49264,N_41608,N_40657);
nor U49265 (N_49265,N_41197,N_43975);
or U49266 (N_49266,N_43747,N_41065);
xnor U49267 (N_49267,N_43641,N_43083);
or U49268 (N_49268,N_43094,N_42451);
nor U49269 (N_49269,N_44211,N_41881);
and U49270 (N_49270,N_43812,N_43786);
nor U49271 (N_49271,N_41518,N_44263);
xor U49272 (N_49272,N_41734,N_40885);
or U49273 (N_49273,N_42068,N_40428);
nor U49274 (N_49274,N_40998,N_42274);
nor U49275 (N_49275,N_41550,N_44610);
xor U49276 (N_49276,N_43181,N_43898);
xor U49277 (N_49277,N_43768,N_41769);
and U49278 (N_49278,N_43180,N_41597);
and U49279 (N_49279,N_41235,N_44040);
xor U49280 (N_49280,N_42793,N_41391);
and U49281 (N_49281,N_44174,N_43956);
nand U49282 (N_49282,N_40789,N_40260);
xor U49283 (N_49283,N_40612,N_43500);
nor U49284 (N_49284,N_44497,N_43681);
or U49285 (N_49285,N_43638,N_40713);
xor U49286 (N_49286,N_41465,N_43339);
nand U49287 (N_49287,N_40082,N_44624);
xnor U49288 (N_49288,N_44248,N_42134);
and U49289 (N_49289,N_43576,N_43481);
and U49290 (N_49290,N_43069,N_41877);
or U49291 (N_49291,N_44359,N_43805);
xnor U49292 (N_49292,N_41017,N_43358);
nand U49293 (N_49293,N_42370,N_42899);
or U49294 (N_49294,N_40844,N_42744);
nor U49295 (N_49295,N_44785,N_44570);
or U49296 (N_49296,N_44371,N_40435);
nand U49297 (N_49297,N_43754,N_44336);
xnor U49298 (N_49298,N_44732,N_43138);
and U49299 (N_49299,N_42749,N_44069);
and U49300 (N_49300,N_41803,N_44237);
nand U49301 (N_49301,N_43068,N_42342);
or U49302 (N_49302,N_44867,N_43536);
and U49303 (N_49303,N_41409,N_44245);
nor U49304 (N_49304,N_44016,N_41522);
xor U49305 (N_49305,N_41384,N_44000);
nand U49306 (N_49306,N_41506,N_41959);
or U49307 (N_49307,N_42131,N_41660);
nor U49308 (N_49308,N_42458,N_43357);
and U49309 (N_49309,N_40420,N_43281);
and U49310 (N_49310,N_44248,N_40099);
xor U49311 (N_49311,N_41373,N_42571);
or U49312 (N_49312,N_41323,N_43990);
and U49313 (N_49313,N_41795,N_40992);
and U49314 (N_49314,N_43549,N_44730);
nor U49315 (N_49315,N_40588,N_44871);
nor U49316 (N_49316,N_40699,N_42530);
and U49317 (N_49317,N_42088,N_40614);
or U49318 (N_49318,N_43199,N_43734);
nor U49319 (N_49319,N_43003,N_41467);
and U49320 (N_49320,N_41354,N_40270);
nor U49321 (N_49321,N_42465,N_41485);
xnor U49322 (N_49322,N_43074,N_42742);
and U49323 (N_49323,N_41253,N_40377);
xor U49324 (N_49324,N_43884,N_40408);
or U49325 (N_49325,N_42939,N_40382);
nand U49326 (N_49326,N_43732,N_40114);
xnor U49327 (N_49327,N_41563,N_44714);
and U49328 (N_49328,N_44377,N_41009);
nand U49329 (N_49329,N_44786,N_44626);
xnor U49330 (N_49330,N_41358,N_41149);
or U49331 (N_49331,N_44812,N_44665);
nand U49332 (N_49332,N_41041,N_43643);
xor U49333 (N_49333,N_42293,N_42159);
nand U49334 (N_49334,N_44943,N_43680);
xnor U49335 (N_49335,N_41149,N_40108);
and U49336 (N_49336,N_41824,N_43774);
or U49337 (N_49337,N_44560,N_41824);
nor U49338 (N_49338,N_43125,N_44874);
xnor U49339 (N_49339,N_44178,N_43109);
or U49340 (N_49340,N_44085,N_41897);
nor U49341 (N_49341,N_41259,N_43632);
nand U49342 (N_49342,N_40318,N_42618);
nor U49343 (N_49343,N_42838,N_40181);
nand U49344 (N_49344,N_41278,N_44472);
xnor U49345 (N_49345,N_44441,N_42253);
nand U49346 (N_49346,N_43718,N_42323);
xnor U49347 (N_49347,N_42152,N_42889);
and U49348 (N_49348,N_42259,N_41847);
and U49349 (N_49349,N_43344,N_40235);
nand U49350 (N_49350,N_40382,N_41768);
nor U49351 (N_49351,N_43169,N_43487);
nor U49352 (N_49352,N_42164,N_40473);
nand U49353 (N_49353,N_43909,N_40554);
xnor U49354 (N_49354,N_40738,N_41513);
and U49355 (N_49355,N_44036,N_40789);
nand U49356 (N_49356,N_42773,N_42755);
nor U49357 (N_49357,N_43052,N_40004);
nand U49358 (N_49358,N_41894,N_43466);
nor U49359 (N_49359,N_41366,N_43303);
and U49360 (N_49360,N_42181,N_43353);
and U49361 (N_49361,N_42721,N_41471);
xor U49362 (N_49362,N_41668,N_44776);
and U49363 (N_49363,N_41075,N_40278);
nand U49364 (N_49364,N_42538,N_43580);
nand U49365 (N_49365,N_44262,N_42718);
or U49366 (N_49366,N_40889,N_43516);
or U49367 (N_49367,N_42626,N_43539);
nor U49368 (N_49368,N_44629,N_42594);
nand U49369 (N_49369,N_42295,N_43448);
nand U49370 (N_49370,N_40815,N_43414);
nor U49371 (N_49371,N_44451,N_44050);
xnor U49372 (N_49372,N_44366,N_41452);
nor U49373 (N_49373,N_43004,N_44373);
xnor U49374 (N_49374,N_41094,N_40299);
or U49375 (N_49375,N_42416,N_40545);
nand U49376 (N_49376,N_42617,N_42571);
and U49377 (N_49377,N_42082,N_42622);
or U49378 (N_49378,N_44799,N_42679);
or U49379 (N_49379,N_44100,N_41297);
xor U49380 (N_49380,N_44015,N_44284);
nor U49381 (N_49381,N_42718,N_44707);
or U49382 (N_49382,N_40274,N_44921);
nand U49383 (N_49383,N_40361,N_41305);
nor U49384 (N_49384,N_40644,N_43215);
xnor U49385 (N_49385,N_41732,N_44967);
and U49386 (N_49386,N_44047,N_42260);
xnor U49387 (N_49387,N_40601,N_42565);
and U49388 (N_49388,N_44017,N_42377);
xor U49389 (N_49389,N_42186,N_40037);
or U49390 (N_49390,N_41542,N_42177);
or U49391 (N_49391,N_43001,N_40884);
nand U49392 (N_49392,N_43490,N_43492);
nor U49393 (N_49393,N_42122,N_40702);
and U49394 (N_49394,N_44478,N_43191);
and U49395 (N_49395,N_43699,N_42355);
nand U49396 (N_49396,N_40000,N_43550);
and U49397 (N_49397,N_41954,N_40027);
and U49398 (N_49398,N_41484,N_43860);
xnor U49399 (N_49399,N_44460,N_42214);
xor U49400 (N_49400,N_41683,N_40230);
nand U49401 (N_49401,N_43759,N_43564);
nand U49402 (N_49402,N_44514,N_41295);
nor U49403 (N_49403,N_42975,N_42490);
and U49404 (N_49404,N_42623,N_43408);
nand U49405 (N_49405,N_41581,N_40140);
or U49406 (N_49406,N_40542,N_41968);
nand U49407 (N_49407,N_40764,N_43989);
nor U49408 (N_49408,N_44369,N_40796);
nor U49409 (N_49409,N_42576,N_42246);
nor U49410 (N_49410,N_43081,N_42592);
xnor U49411 (N_49411,N_41940,N_44535);
nor U49412 (N_49412,N_41192,N_41990);
and U49413 (N_49413,N_42195,N_42211);
nor U49414 (N_49414,N_40535,N_44049);
and U49415 (N_49415,N_40150,N_42051);
nor U49416 (N_49416,N_43899,N_41167);
or U49417 (N_49417,N_44076,N_42831);
xor U49418 (N_49418,N_42473,N_43923);
nor U49419 (N_49419,N_41333,N_41983);
or U49420 (N_49420,N_42822,N_42091);
and U49421 (N_49421,N_43623,N_40904);
nor U49422 (N_49422,N_41129,N_42979);
and U49423 (N_49423,N_42885,N_41097);
or U49424 (N_49424,N_43086,N_43958);
nand U49425 (N_49425,N_42864,N_42074);
nor U49426 (N_49426,N_42795,N_41991);
xor U49427 (N_49427,N_43023,N_40834);
nand U49428 (N_49428,N_44678,N_42113);
xnor U49429 (N_49429,N_41056,N_44208);
and U49430 (N_49430,N_40025,N_40283);
and U49431 (N_49431,N_41886,N_43801);
xor U49432 (N_49432,N_43556,N_42074);
or U49433 (N_49433,N_41057,N_43823);
or U49434 (N_49434,N_43461,N_42742);
and U49435 (N_49435,N_44946,N_41600);
xnor U49436 (N_49436,N_40804,N_43989);
nand U49437 (N_49437,N_40721,N_43154);
nand U49438 (N_49438,N_42315,N_40028);
xnor U49439 (N_49439,N_44455,N_42712);
and U49440 (N_49440,N_44467,N_44642);
xnor U49441 (N_49441,N_40608,N_43021);
or U49442 (N_49442,N_43741,N_42937);
nor U49443 (N_49443,N_42086,N_44415);
or U49444 (N_49444,N_43879,N_42962);
and U49445 (N_49445,N_40441,N_44500);
or U49446 (N_49446,N_42915,N_41319);
and U49447 (N_49447,N_43827,N_40602);
xor U49448 (N_49448,N_44441,N_41086);
nand U49449 (N_49449,N_44885,N_43589);
nand U49450 (N_49450,N_43179,N_41798);
nor U49451 (N_49451,N_43004,N_42185);
nor U49452 (N_49452,N_42409,N_44486);
nor U49453 (N_49453,N_40899,N_40577);
nor U49454 (N_49454,N_44989,N_40188);
xor U49455 (N_49455,N_44669,N_40970);
or U49456 (N_49456,N_41401,N_43802);
or U49457 (N_49457,N_42473,N_43642);
nor U49458 (N_49458,N_40726,N_42617);
or U49459 (N_49459,N_44634,N_42389);
nand U49460 (N_49460,N_41069,N_44713);
or U49461 (N_49461,N_43485,N_44698);
nor U49462 (N_49462,N_43652,N_44939);
xor U49463 (N_49463,N_42003,N_42013);
and U49464 (N_49464,N_40777,N_41433);
nor U49465 (N_49465,N_40419,N_40742);
nand U49466 (N_49466,N_43184,N_42807);
and U49467 (N_49467,N_42507,N_44615);
nor U49468 (N_49468,N_43721,N_41285);
or U49469 (N_49469,N_40800,N_41656);
nor U49470 (N_49470,N_42409,N_43797);
xor U49471 (N_49471,N_41581,N_43145);
nor U49472 (N_49472,N_42424,N_44488);
xnor U49473 (N_49473,N_43502,N_43340);
or U49474 (N_49474,N_41538,N_43819);
or U49475 (N_49475,N_44231,N_40167);
or U49476 (N_49476,N_40618,N_44938);
and U49477 (N_49477,N_44288,N_42677);
nor U49478 (N_49478,N_42346,N_42828);
and U49479 (N_49479,N_42688,N_41604);
or U49480 (N_49480,N_44041,N_44508);
or U49481 (N_49481,N_40742,N_42932);
nor U49482 (N_49482,N_40734,N_43947);
and U49483 (N_49483,N_41081,N_40477);
xnor U49484 (N_49484,N_40024,N_40338);
and U49485 (N_49485,N_44137,N_41014);
nand U49486 (N_49486,N_40490,N_41919);
or U49487 (N_49487,N_42807,N_40396);
nand U49488 (N_49488,N_42898,N_41850);
and U49489 (N_49489,N_43508,N_42439);
xnor U49490 (N_49490,N_42666,N_40357);
nand U49491 (N_49491,N_42169,N_41392);
and U49492 (N_49492,N_40715,N_44663);
nor U49493 (N_49493,N_41731,N_41721);
and U49494 (N_49494,N_42306,N_43431);
nand U49495 (N_49495,N_41746,N_41597);
nor U49496 (N_49496,N_42788,N_43407);
nand U49497 (N_49497,N_43926,N_42220);
nand U49498 (N_49498,N_44120,N_43786);
and U49499 (N_49499,N_44108,N_40589);
nor U49500 (N_49500,N_42549,N_42790);
nor U49501 (N_49501,N_40148,N_44011);
and U49502 (N_49502,N_44544,N_44151);
nor U49503 (N_49503,N_43921,N_44851);
nor U49504 (N_49504,N_41025,N_43566);
nand U49505 (N_49505,N_42672,N_44654);
nand U49506 (N_49506,N_41188,N_42688);
nor U49507 (N_49507,N_42514,N_43921);
nor U49508 (N_49508,N_42042,N_40296);
xor U49509 (N_49509,N_42370,N_40900);
or U49510 (N_49510,N_42367,N_44883);
or U49511 (N_49511,N_44104,N_42005);
and U49512 (N_49512,N_43864,N_43351);
nor U49513 (N_49513,N_44903,N_41703);
nor U49514 (N_49514,N_44371,N_42465);
xnor U49515 (N_49515,N_44204,N_42482);
and U49516 (N_49516,N_44428,N_43534);
or U49517 (N_49517,N_42161,N_41887);
or U49518 (N_49518,N_41885,N_41504);
nor U49519 (N_49519,N_44517,N_40999);
and U49520 (N_49520,N_42611,N_43294);
nand U49521 (N_49521,N_41993,N_40040);
nand U49522 (N_49522,N_43971,N_43998);
or U49523 (N_49523,N_43151,N_43426);
and U49524 (N_49524,N_44772,N_44550);
or U49525 (N_49525,N_43618,N_44266);
and U49526 (N_49526,N_43069,N_40878);
nand U49527 (N_49527,N_41187,N_44036);
and U49528 (N_49528,N_41868,N_44976);
nor U49529 (N_49529,N_41536,N_42642);
and U49530 (N_49530,N_44172,N_42356);
xnor U49531 (N_49531,N_41998,N_41065);
or U49532 (N_49532,N_42975,N_44805);
xor U49533 (N_49533,N_41744,N_41651);
or U49534 (N_49534,N_42148,N_40083);
nor U49535 (N_49535,N_43247,N_40661);
and U49536 (N_49536,N_44184,N_44097);
or U49537 (N_49537,N_41116,N_41981);
nand U49538 (N_49538,N_41558,N_43064);
and U49539 (N_49539,N_43047,N_41146);
xnor U49540 (N_49540,N_43177,N_43907);
xor U49541 (N_49541,N_43634,N_43036);
or U49542 (N_49542,N_42065,N_42503);
nand U49543 (N_49543,N_41473,N_43703);
or U49544 (N_49544,N_41902,N_44530);
and U49545 (N_49545,N_40710,N_41824);
and U49546 (N_49546,N_43413,N_40592);
nand U49547 (N_49547,N_44283,N_41151);
nand U49548 (N_49548,N_42124,N_44328);
and U49549 (N_49549,N_41025,N_42067);
nor U49550 (N_49550,N_43046,N_43433);
or U49551 (N_49551,N_40911,N_42422);
xor U49552 (N_49552,N_40044,N_44967);
xor U49553 (N_49553,N_41729,N_42572);
or U49554 (N_49554,N_41986,N_43074);
xor U49555 (N_49555,N_41484,N_44946);
and U49556 (N_49556,N_44111,N_44918);
nor U49557 (N_49557,N_42620,N_41289);
nor U49558 (N_49558,N_43824,N_43441);
nor U49559 (N_49559,N_43941,N_40261);
xor U49560 (N_49560,N_42506,N_41810);
nor U49561 (N_49561,N_40901,N_43824);
nand U49562 (N_49562,N_42725,N_40801);
nor U49563 (N_49563,N_40018,N_40452);
nand U49564 (N_49564,N_44114,N_44387);
or U49565 (N_49565,N_44866,N_41942);
and U49566 (N_49566,N_44266,N_43575);
nor U49567 (N_49567,N_41202,N_43993);
xnor U49568 (N_49568,N_42381,N_43723);
or U49569 (N_49569,N_43768,N_44091);
and U49570 (N_49570,N_43559,N_43863);
nor U49571 (N_49571,N_41906,N_43965);
and U49572 (N_49572,N_41011,N_40605);
xor U49573 (N_49573,N_43153,N_42015);
xnor U49574 (N_49574,N_43373,N_41623);
nor U49575 (N_49575,N_44483,N_40984);
or U49576 (N_49576,N_44982,N_40032);
or U49577 (N_49577,N_40823,N_44695);
or U49578 (N_49578,N_41962,N_40258);
and U49579 (N_49579,N_40115,N_44707);
and U49580 (N_49580,N_40078,N_41720);
or U49581 (N_49581,N_42226,N_42626);
nor U49582 (N_49582,N_44983,N_43023);
xor U49583 (N_49583,N_40618,N_42645);
nand U49584 (N_49584,N_40615,N_41532);
nand U49585 (N_49585,N_41619,N_42570);
nand U49586 (N_49586,N_40186,N_42759);
nand U49587 (N_49587,N_40499,N_43083);
nor U49588 (N_49588,N_43346,N_40966);
and U49589 (N_49589,N_41021,N_41236);
or U49590 (N_49590,N_41107,N_40370);
xor U49591 (N_49591,N_40045,N_41252);
xnor U49592 (N_49592,N_43584,N_43549);
and U49593 (N_49593,N_42300,N_41607);
xor U49594 (N_49594,N_43088,N_41951);
or U49595 (N_49595,N_43470,N_44892);
nand U49596 (N_49596,N_40559,N_44133);
nand U49597 (N_49597,N_40879,N_43484);
nor U49598 (N_49598,N_42949,N_43303);
or U49599 (N_49599,N_40476,N_42806);
xnor U49600 (N_49600,N_44716,N_44458);
or U49601 (N_49601,N_42651,N_44202);
nand U49602 (N_49602,N_40774,N_43368);
nand U49603 (N_49603,N_42597,N_40490);
xnor U49604 (N_49604,N_42063,N_40504);
nand U49605 (N_49605,N_40920,N_44737);
nand U49606 (N_49606,N_43854,N_41467);
xnor U49607 (N_49607,N_40051,N_44956);
and U49608 (N_49608,N_41115,N_43146);
xor U49609 (N_49609,N_43295,N_42403);
xnor U49610 (N_49610,N_41613,N_41540);
nor U49611 (N_49611,N_44686,N_44401);
nor U49612 (N_49612,N_43448,N_44101);
nor U49613 (N_49613,N_44471,N_44995);
or U49614 (N_49614,N_41570,N_40433);
nor U49615 (N_49615,N_42974,N_40718);
nor U49616 (N_49616,N_40355,N_42085);
xnor U49617 (N_49617,N_40646,N_41574);
and U49618 (N_49618,N_41353,N_44043);
xor U49619 (N_49619,N_43374,N_40211);
xnor U49620 (N_49620,N_43489,N_44536);
xnor U49621 (N_49621,N_44704,N_44761);
nor U49622 (N_49622,N_41315,N_44398);
xnor U49623 (N_49623,N_44748,N_42933);
nand U49624 (N_49624,N_40926,N_44099);
xor U49625 (N_49625,N_41372,N_44386);
or U49626 (N_49626,N_41385,N_40368);
xnor U49627 (N_49627,N_41722,N_43255);
or U49628 (N_49628,N_44737,N_44713);
and U49629 (N_49629,N_44180,N_40434);
and U49630 (N_49630,N_40356,N_40830);
or U49631 (N_49631,N_41334,N_42106);
nor U49632 (N_49632,N_41245,N_41185);
and U49633 (N_49633,N_40745,N_41786);
nor U49634 (N_49634,N_42487,N_43968);
xnor U49635 (N_49635,N_41785,N_43665);
nor U49636 (N_49636,N_41284,N_43199);
or U49637 (N_49637,N_42461,N_43004);
and U49638 (N_49638,N_43522,N_43973);
or U49639 (N_49639,N_40245,N_41200);
and U49640 (N_49640,N_42836,N_41394);
nand U49641 (N_49641,N_42787,N_41619);
nand U49642 (N_49642,N_41210,N_43199);
and U49643 (N_49643,N_43253,N_40270);
or U49644 (N_49644,N_42234,N_42119);
and U49645 (N_49645,N_42554,N_41589);
nor U49646 (N_49646,N_43846,N_41969);
nor U49647 (N_49647,N_40704,N_40966);
and U49648 (N_49648,N_42360,N_43602);
and U49649 (N_49649,N_44182,N_44626);
xor U49650 (N_49650,N_41013,N_42677);
nand U49651 (N_49651,N_43839,N_42960);
and U49652 (N_49652,N_42263,N_42871);
xnor U49653 (N_49653,N_41803,N_40461);
xor U49654 (N_49654,N_40387,N_44928);
nand U49655 (N_49655,N_43500,N_40070);
nand U49656 (N_49656,N_44772,N_41183);
xor U49657 (N_49657,N_41762,N_40941);
and U49658 (N_49658,N_44682,N_42588);
xor U49659 (N_49659,N_42673,N_42741);
xnor U49660 (N_49660,N_41446,N_43512);
nor U49661 (N_49661,N_42069,N_43928);
or U49662 (N_49662,N_42267,N_43224);
nand U49663 (N_49663,N_42698,N_40368);
and U49664 (N_49664,N_40830,N_44678);
or U49665 (N_49665,N_42139,N_40961);
and U49666 (N_49666,N_40897,N_44317);
and U49667 (N_49667,N_40480,N_44742);
xnor U49668 (N_49668,N_44048,N_42397);
and U49669 (N_49669,N_44238,N_43404);
or U49670 (N_49670,N_42703,N_42460);
or U49671 (N_49671,N_44037,N_41987);
and U49672 (N_49672,N_44960,N_40701);
and U49673 (N_49673,N_44825,N_44537);
xnor U49674 (N_49674,N_44833,N_40314);
xnor U49675 (N_49675,N_41891,N_44240);
and U49676 (N_49676,N_41250,N_44307);
or U49677 (N_49677,N_43380,N_40135);
xor U49678 (N_49678,N_42955,N_40764);
and U49679 (N_49679,N_44596,N_44235);
xnor U49680 (N_49680,N_40319,N_44133);
xnor U49681 (N_49681,N_43157,N_43607);
or U49682 (N_49682,N_43873,N_44879);
nand U49683 (N_49683,N_43928,N_42378);
nand U49684 (N_49684,N_41471,N_41805);
nor U49685 (N_49685,N_40382,N_43689);
or U49686 (N_49686,N_41878,N_42465);
and U49687 (N_49687,N_40701,N_44182);
nor U49688 (N_49688,N_42131,N_41672);
xnor U49689 (N_49689,N_40882,N_42271);
nor U49690 (N_49690,N_44161,N_43249);
xor U49691 (N_49691,N_41331,N_40884);
and U49692 (N_49692,N_41958,N_44338);
xor U49693 (N_49693,N_44859,N_40005);
xnor U49694 (N_49694,N_41327,N_44960);
xnor U49695 (N_49695,N_41733,N_40981);
or U49696 (N_49696,N_44718,N_41254);
and U49697 (N_49697,N_44896,N_41664);
or U49698 (N_49698,N_41233,N_41264);
nor U49699 (N_49699,N_41850,N_43222);
or U49700 (N_49700,N_44598,N_41564);
nor U49701 (N_49701,N_43892,N_43958);
nor U49702 (N_49702,N_41290,N_40292);
nor U49703 (N_49703,N_44922,N_42463);
or U49704 (N_49704,N_44773,N_40709);
nor U49705 (N_49705,N_41823,N_43694);
xor U49706 (N_49706,N_41064,N_42390);
or U49707 (N_49707,N_42308,N_41564);
or U49708 (N_49708,N_43403,N_43026);
and U49709 (N_49709,N_43486,N_43999);
nor U49710 (N_49710,N_40848,N_41389);
and U49711 (N_49711,N_42890,N_44727);
and U49712 (N_49712,N_44983,N_43677);
nor U49713 (N_49713,N_44110,N_40642);
and U49714 (N_49714,N_43267,N_44078);
or U49715 (N_49715,N_42493,N_40120);
nand U49716 (N_49716,N_42228,N_44703);
nor U49717 (N_49717,N_43560,N_41928);
nand U49718 (N_49718,N_40857,N_42054);
nor U49719 (N_49719,N_40946,N_43761);
nor U49720 (N_49720,N_40036,N_40820);
and U49721 (N_49721,N_42660,N_43643);
and U49722 (N_49722,N_43330,N_43187);
and U49723 (N_49723,N_43805,N_42514);
and U49724 (N_49724,N_40897,N_44180);
nand U49725 (N_49725,N_44337,N_42428);
or U49726 (N_49726,N_44870,N_43864);
and U49727 (N_49727,N_41267,N_43625);
nand U49728 (N_49728,N_44914,N_40870);
and U49729 (N_49729,N_40627,N_44049);
xor U49730 (N_49730,N_40089,N_40288);
or U49731 (N_49731,N_42408,N_44613);
xnor U49732 (N_49732,N_40602,N_40510);
nand U49733 (N_49733,N_42719,N_42880);
xnor U49734 (N_49734,N_43204,N_41938);
nand U49735 (N_49735,N_43830,N_43748);
xnor U49736 (N_49736,N_41531,N_41959);
and U49737 (N_49737,N_41297,N_43258);
nand U49738 (N_49738,N_41691,N_42421);
or U49739 (N_49739,N_43717,N_40483);
and U49740 (N_49740,N_41134,N_41785);
and U49741 (N_49741,N_40050,N_42524);
and U49742 (N_49742,N_40234,N_43775);
xnor U49743 (N_49743,N_42821,N_40479);
xnor U49744 (N_49744,N_41958,N_41358);
and U49745 (N_49745,N_40182,N_41869);
xor U49746 (N_49746,N_41138,N_40970);
or U49747 (N_49747,N_43046,N_44989);
and U49748 (N_49748,N_43886,N_40484);
xnor U49749 (N_49749,N_41705,N_44843);
nand U49750 (N_49750,N_43473,N_43114);
and U49751 (N_49751,N_41680,N_42724);
nand U49752 (N_49752,N_41934,N_44793);
nor U49753 (N_49753,N_44019,N_41513);
nand U49754 (N_49754,N_44867,N_42366);
nor U49755 (N_49755,N_43491,N_40974);
and U49756 (N_49756,N_40844,N_42299);
xnor U49757 (N_49757,N_40566,N_41110);
nor U49758 (N_49758,N_44983,N_41980);
and U49759 (N_49759,N_43596,N_44997);
nor U49760 (N_49760,N_40069,N_41106);
xnor U49761 (N_49761,N_40977,N_43345);
or U49762 (N_49762,N_44253,N_41628);
xnor U49763 (N_49763,N_42572,N_41192);
xnor U49764 (N_49764,N_40884,N_44811);
nor U49765 (N_49765,N_40948,N_40143);
or U49766 (N_49766,N_43977,N_41455);
nor U49767 (N_49767,N_42051,N_43711);
nor U49768 (N_49768,N_44364,N_43890);
nand U49769 (N_49769,N_44983,N_44390);
or U49770 (N_49770,N_42362,N_44908);
and U49771 (N_49771,N_44786,N_41155);
nand U49772 (N_49772,N_43684,N_40196);
and U49773 (N_49773,N_40429,N_41839);
and U49774 (N_49774,N_43720,N_41908);
or U49775 (N_49775,N_43907,N_40160);
nor U49776 (N_49776,N_41138,N_42858);
nor U49777 (N_49777,N_42732,N_43261);
and U49778 (N_49778,N_44028,N_41588);
and U49779 (N_49779,N_41112,N_44031);
nand U49780 (N_49780,N_44455,N_42647);
nand U49781 (N_49781,N_40060,N_40437);
nand U49782 (N_49782,N_40703,N_42466);
nor U49783 (N_49783,N_41366,N_40767);
xnor U49784 (N_49784,N_41078,N_42819);
or U49785 (N_49785,N_41099,N_40774);
nand U49786 (N_49786,N_43290,N_41841);
xnor U49787 (N_49787,N_43588,N_41142);
nor U49788 (N_49788,N_44050,N_40758);
nand U49789 (N_49789,N_40200,N_43059);
xnor U49790 (N_49790,N_40801,N_42352);
xnor U49791 (N_49791,N_41816,N_44472);
nand U49792 (N_49792,N_42770,N_40141);
nand U49793 (N_49793,N_42827,N_41798);
or U49794 (N_49794,N_44955,N_44614);
nand U49795 (N_49795,N_41110,N_44861);
or U49796 (N_49796,N_40229,N_43961);
nor U49797 (N_49797,N_42269,N_41946);
xor U49798 (N_49798,N_44352,N_40404);
nor U49799 (N_49799,N_40831,N_42485);
or U49800 (N_49800,N_40553,N_44181);
nand U49801 (N_49801,N_42324,N_40136);
or U49802 (N_49802,N_43514,N_44341);
nand U49803 (N_49803,N_44868,N_44600);
nor U49804 (N_49804,N_44981,N_42989);
nand U49805 (N_49805,N_43718,N_42626);
xnor U49806 (N_49806,N_41598,N_44644);
and U49807 (N_49807,N_40997,N_44088);
xnor U49808 (N_49808,N_41639,N_42957);
or U49809 (N_49809,N_44536,N_43282);
or U49810 (N_49810,N_42395,N_40504);
nor U49811 (N_49811,N_40310,N_40653);
nand U49812 (N_49812,N_44499,N_41962);
nand U49813 (N_49813,N_41566,N_42978);
or U49814 (N_49814,N_40658,N_41749);
and U49815 (N_49815,N_41674,N_42097);
or U49816 (N_49816,N_44769,N_42136);
nand U49817 (N_49817,N_41232,N_42018);
xor U49818 (N_49818,N_44568,N_44463);
xor U49819 (N_49819,N_41044,N_42430);
nand U49820 (N_49820,N_40550,N_40757);
nand U49821 (N_49821,N_43377,N_42271);
and U49822 (N_49822,N_40781,N_41244);
nand U49823 (N_49823,N_43845,N_41021);
xnor U49824 (N_49824,N_44050,N_41700);
nand U49825 (N_49825,N_44842,N_40189);
xor U49826 (N_49826,N_44586,N_41189);
xor U49827 (N_49827,N_42105,N_41898);
nand U49828 (N_49828,N_44667,N_40909);
nor U49829 (N_49829,N_41228,N_40152);
nor U49830 (N_49830,N_41863,N_43176);
nor U49831 (N_49831,N_40381,N_42756);
nand U49832 (N_49832,N_43267,N_44062);
and U49833 (N_49833,N_43098,N_44828);
nand U49834 (N_49834,N_42285,N_40715);
nand U49835 (N_49835,N_43863,N_41377);
and U49836 (N_49836,N_40224,N_41636);
or U49837 (N_49837,N_40696,N_40875);
or U49838 (N_49838,N_44029,N_43439);
and U49839 (N_49839,N_41895,N_44736);
or U49840 (N_49840,N_41549,N_43097);
or U49841 (N_49841,N_43102,N_42243);
xnor U49842 (N_49842,N_44825,N_43667);
and U49843 (N_49843,N_41069,N_40481);
or U49844 (N_49844,N_44077,N_41677);
and U49845 (N_49845,N_43806,N_40360);
or U49846 (N_49846,N_42300,N_42869);
nor U49847 (N_49847,N_40182,N_43588);
or U49848 (N_49848,N_41663,N_42493);
and U49849 (N_49849,N_41835,N_43442);
xnor U49850 (N_49850,N_42147,N_44068);
xnor U49851 (N_49851,N_41801,N_40427);
nand U49852 (N_49852,N_42411,N_41137);
or U49853 (N_49853,N_44390,N_40569);
xor U49854 (N_49854,N_40009,N_42119);
xnor U49855 (N_49855,N_42963,N_41651);
and U49856 (N_49856,N_42990,N_44372);
nand U49857 (N_49857,N_41605,N_40097);
or U49858 (N_49858,N_43107,N_42346);
and U49859 (N_49859,N_41583,N_41031);
or U49860 (N_49860,N_44863,N_41962);
nand U49861 (N_49861,N_44957,N_42887);
nor U49862 (N_49862,N_41724,N_40432);
nand U49863 (N_49863,N_43040,N_44292);
xnor U49864 (N_49864,N_40215,N_43595);
nand U49865 (N_49865,N_44980,N_42132);
xor U49866 (N_49866,N_42679,N_40097);
nor U49867 (N_49867,N_41369,N_40576);
nor U49868 (N_49868,N_43850,N_40367);
nand U49869 (N_49869,N_40350,N_42775);
and U49870 (N_49870,N_40251,N_41550);
xor U49871 (N_49871,N_43155,N_42235);
nor U49872 (N_49872,N_40359,N_43425);
nand U49873 (N_49873,N_44213,N_41262);
nand U49874 (N_49874,N_40190,N_41420);
xor U49875 (N_49875,N_41886,N_43042);
nand U49876 (N_49876,N_44102,N_40206);
or U49877 (N_49877,N_42624,N_43413);
and U49878 (N_49878,N_43555,N_43862);
or U49879 (N_49879,N_43425,N_44932);
nor U49880 (N_49880,N_43627,N_41135);
nand U49881 (N_49881,N_42781,N_44033);
and U49882 (N_49882,N_41341,N_43218);
or U49883 (N_49883,N_43448,N_44924);
or U49884 (N_49884,N_43961,N_41528);
xnor U49885 (N_49885,N_43084,N_41873);
nor U49886 (N_49886,N_40367,N_43527);
nor U49887 (N_49887,N_43410,N_40845);
and U49888 (N_49888,N_41629,N_44088);
nor U49889 (N_49889,N_41617,N_40841);
xnor U49890 (N_49890,N_41075,N_44513);
nand U49891 (N_49891,N_40007,N_44331);
xor U49892 (N_49892,N_44757,N_43450);
nor U49893 (N_49893,N_42092,N_40917);
xnor U49894 (N_49894,N_42596,N_40918);
nand U49895 (N_49895,N_44654,N_42797);
nor U49896 (N_49896,N_41729,N_42621);
nand U49897 (N_49897,N_44429,N_40075);
and U49898 (N_49898,N_44670,N_40421);
and U49899 (N_49899,N_44598,N_41160);
and U49900 (N_49900,N_40924,N_40867);
nand U49901 (N_49901,N_44092,N_43823);
xor U49902 (N_49902,N_43883,N_41698);
nand U49903 (N_49903,N_41646,N_42494);
and U49904 (N_49904,N_43173,N_42286);
nor U49905 (N_49905,N_44270,N_40549);
xor U49906 (N_49906,N_44906,N_43003);
xnor U49907 (N_49907,N_43736,N_43729);
nor U49908 (N_49908,N_43841,N_41564);
nor U49909 (N_49909,N_43535,N_44126);
or U49910 (N_49910,N_44672,N_44046);
or U49911 (N_49911,N_43292,N_42780);
and U49912 (N_49912,N_42159,N_44863);
xor U49913 (N_49913,N_44276,N_44295);
and U49914 (N_49914,N_42812,N_40894);
xor U49915 (N_49915,N_41660,N_40300);
or U49916 (N_49916,N_43597,N_44232);
xnor U49917 (N_49917,N_44899,N_40765);
and U49918 (N_49918,N_42079,N_44644);
nand U49919 (N_49919,N_44419,N_40926);
xnor U49920 (N_49920,N_41926,N_40211);
xnor U49921 (N_49921,N_43596,N_43084);
xnor U49922 (N_49922,N_44026,N_44301);
and U49923 (N_49923,N_44367,N_44395);
or U49924 (N_49924,N_43179,N_44020);
xnor U49925 (N_49925,N_42735,N_41698);
and U49926 (N_49926,N_42750,N_43377);
nor U49927 (N_49927,N_44500,N_43059);
and U49928 (N_49928,N_41322,N_43279);
and U49929 (N_49929,N_41531,N_41836);
and U49930 (N_49930,N_40888,N_44823);
and U49931 (N_49931,N_41041,N_42317);
or U49932 (N_49932,N_42996,N_43617);
and U49933 (N_49933,N_42106,N_40378);
nor U49934 (N_49934,N_44393,N_43654);
and U49935 (N_49935,N_41375,N_40032);
nand U49936 (N_49936,N_42541,N_43794);
or U49937 (N_49937,N_42390,N_40598);
nor U49938 (N_49938,N_40137,N_42601);
nand U49939 (N_49939,N_44572,N_43393);
or U49940 (N_49940,N_43930,N_42860);
nor U49941 (N_49941,N_42488,N_40922);
xor U49942 (N_49942,N_40075,N_42304);
nand U49943 (N_49943,N_43997,N_44117);
nand U49944 (N_49944,N_40059,N_43144);
nand U49945 (N_49945,N_43963,N_43005);
nor U49946 (N_49946,N_43649,N_42328);
xor U49947 (N_49947,N_41728,N_43388);
nand U49948 (N_49948,N_44787,N_40760);
nand U49949 (N_49949,N_40819,N_41755);
and U49950 (N_49950,N_40005,N_41299);
nand U49951 (N_49951,N_42526,N_42900);
nor U49952 (N_49952,N_43513,N_43813);
nand U49953 (N_49953,N_40066,N_44772);
nand U49954 (N_49954,N_41118,N_44095);
nand U49955 (N_49955,N_41168,N_40859);
nand U49956 (N_49956,N_44670,N_43754);
xor U49957 (N_49957,N_43293,N_44672);
and U49958 (N_49958,N_43760,N_44306);
xor U49959 (N_49959,N_44717,N_44730);
nor U49960 (N_49960,N_40917,N_42291);
and U49961 (N_49961,N_40764,N_42994);
or U49962 (N_49962,N_42253,N_44731);
nand U49963 (N_49963,N_44285,N_41358);
and U49964 (N_49964,N_42786,N_44535);
nor U49965 (N_49965,N_40357,N_42893);
or U49966 (N_49966,N_40378,N_40382);
xnor U49967 (N_49967,N_41567,N_42920);
or U49968 (N_49968,N_40187,N_41138);
nor U49969 (N_49969,N_40791,N_40050);
or U49970 (N_49970,N_43523,N_40174);
xnor U49971 (N_49971,N_42419,N_44155);
nand U49972 (N_49972,N_42283,N_44235);
and U49973 (N_49973,N_43109,N_44144);
nor U49974 (N_49974,N_44027,N_44607);
nand U49975 (N_49975,N_44683,N_41530);
nor U49976 (N_49976,N_43362,N_44268);
and U49977 (N_49977,N_44938,N_40012);
or U49978 (N_49978,N_44587,N_41122);
nand U49979 (N_49979,N_42372,N_42999);
xnor U49980 (N_49980,N_44346,N_41099);
nand U49981 (N_49981,N_43250,N_41333);
nand U49982 (N_49982,N_41208,N_44308);
or U49983 (N_49983,N_43355,N_42065);
xnor U49984 (N_49984,N_40074,N_42041);
nor U49985 (N_49985,N_42708,N_40218);
nand U49986 (N_49986,N_44097,N_43310);
xnor U49987 (N_49987,N_42982,N_44020);
or U49988 (N_49988,N_42426,N_44892);
and U49989 (N_49989,N_41276,N_40447);
nand U49990 (N_49990,N_42909,N_41284);
nor U49991 (N_49991,N_43259,N_40337);
nor U49992 (N_49992,N_43060,N_40122);
nand U49993 (N_49993,N_44656,N_41985);
or U49994 (N_49994,N_43520,N_41351);
nand U49995 (N_49995,N_40322,N_40367);
nor U49996 (N_49996,N_44865,N_42003);
or U49997 (N_49997,N_40573,N_42634);
nor U49998 (N_49998,N_43048,N_44016);
nand U49999 (N_49999,N_40219,N_43588);
nand UO_0 (O_0,N_47855,N_45285);
xor UO_1 (O_1,N_46961,N_47792);
nand UO_2 (O_2,N_45320,N_47427);
xnor UO_3 (O_3,N_48626,N_45158);
or UO_4 (O_4,N_49344,N_45429);
nor UO_5 (O_5,N_45630,N_47941);
xnor UO_6 (O_6,N_49995,N_47768);
xor UO_7 (O_7,N_47955,N_46765);
xnor UO_8 (O_8,N_49613,N_49747);
or UO_9 (O_9,N_45244,N_47045);
xor UO_10 (O_10,N_46785,N_48300);
nor UO_11 (O_11,N_48460,N_47536);
nand UO_12 (O_12,N_48683,N_47908);
or UO_13 (O_13,N_49351,N_49018);
or UO_14 (O_14,N_49542,N_49756);
and UO_15 (O_15,N_48296,N_46536);
and UO_16 (O_16,N_45115,N_48487);
nor UO_17 (O_17,N_45176,N_48452);
and UO_18 (O_18,N_48707,N_46324);
nand UO_19 (O_19,N_46671,N_48503);
or UO_20 (O_20,N_45246,N_49850);
nand UO_21 (O_21,N_45649,N_48987);
and UO_22 (O_22,N_45719,N_46694);
or UO_23 (O_23,N_48163,N_45866);
or UO_24 (O_24,N_49363,N_46243);
nor UO_25 (O_25,N_49380,N_46945);
or UO_26 (O_26,N_48100,N_47502);
xor UO_27 (O_27,N_48011,N_47617);
or UO_28 (O_28,N_47154,N_46731);
and UO_29 (O_29,N_46670,N_46552);
or UO_30 (O_30,N_48245,N_48523);
and UO_31 (O_31,N_47547,N_49111);
or UO_32 (O_32,N_45397,N_46036);
nor UO_33 (O_33,N_46613,N_49818);
xor UO_34 (O_34,N_48637,N_49332);
xnor UO_35 (O_35,N_49639,N_48853);
nand UO_36 (O_36,N_47188,N_49792);
nor UO_37 (O_37,N_46296,N_47211);
nand UO_38 (O_38,N_47107,N_47113);
xnor UO_39 (O_39,N_48224,N_48127);
and UO_40 (O_40,N_45769,N_47311);
or UO_41 (O_41,N_47281,N_45020);
or UO_42 (O_42,N_47487,N_47326);
and UO_43 (O_43,N_47708,N_49952);
xor UO_44 (O_44,N_46002,N_48066);
or UO_45 (O_45,N_47883,N_49274);
nand UO_46 (O_46,N_47544,N_49880);
xor UO_47 (O_47,N_46038,N_46768);
and UO_48 (O_48,N_45153,N_49913);
or UO_49 (O_49,N_47538,N_46096);
xor UO_50 (O_50,N_49116,N_46067);
xor UO_51 (O_51,N_46396,N_47011);
or UO_52 (O_52,N_47589,N_45292);
nand UO_53 (O_53,N_48530,N_45608);
xnor UO_54 (O_54,N_47262,N_48781);
nor UO_55 (O_55,N_48198,N_45822);
or UO_56 (O_56,N_48651,N_49766);
xor UO_57 (O_57,N_48541,N_46283);
nand UO_58 (O_58,N_48383,N_48380);
or UO_59 (O_59,N_45766,N_49686);
or UO_60 (O_60,N_46196,N_45718);
or UO_61 (O_61,N_46594,N_48611);
nor UO_62 (O_62,N_46727,N_49482);
nand UO_63 (O_63,N_46678,N_47638);
or UO_64 (O_64,N_45776,N_48823);
or UO_65 (O_65,N_45642,N_48794);
nor UO_66 (O_66,N_45399,N_49016);
nor UO_67 (O_67,N_45744,N_45934);
xor UO_68 (O_68,N_49675,N_45558);
and UO_69 (O_69,N_46474,N_47972);
nor UO_70 (O_70,N_49439,N_49314);
and UO_71 (O_71,N_49647,N_45536);
or UO_72 (O_72,N_47562,N_49265);
and UO_73 (O_73,N_47237,N_45001);
or UO_74 (O_74,N_49964,N_47714);
xnor UO_75 (O_75,N_48228,N_46397);
and UO_76 (O_76,N_48936,N_49395);
nand UO_77 (O_77,N_45539,N_47897);
nor UO_78 (O_78,N_49712,N_46018);
nor UO_79 (O_79,N_49741,N_46439);
and UO_80 (O_80,N_46776,N_48171);
and UO_81 (O_81,N_46369,N_46920);
or UO_82 (O_82,N_47390,N_45696);
nand UO_83 (O_83,N_45964,N_45820);
xnor UO_84 (O_84,N_49735,N_49803);
or UO_85 (O_85,N_47689,N_47456);
nand UO_86 (O_86,N_45532,N_46786);
nor UO_87 (O_87,N_49057,N_46402);
nand UO_88 (O_88,N_48391,N_47587);
and UO_89 (O_89,N_48483,N_46200);
nand UO_90 (O_90,N_49776,N_49075);
and UO_91 (O_91,N_46887,N_49783);
xnor UO_92 (O_92,N_47543,N_48060);
or UO_93 (O_93,N_45182,N_47610);
nand UO_94 (O_94,N_45212,N_46517);
and UO_95 (O_95,N_46391,N_49628);
nand UO_96 (O_96,N_48803,N_45907);
and UO_97 (O_97,N_49157,N_45356);
or UO_98 (O_98,N_48813,N_49900);
xnor UO_99 (O_99,N_45697,N_45440);
xor UO_100 (O_100,N_48511,N_45217);
and UO_101 (O_101,N_47292,N_45078);
and UO_102 (O_102,N_49863,N_49528);
xnor UO_103 (O_103,N_47927,N_46147);
or UO_104 (O_104,N_45906,N_48795);
nand UO_105 (O_105,N_48415,N_47980);
nor UO_106 (O_106,N_47728,N_49584);
or UO_107 (O_107,N_48569,N_46531);
xnor UO_108 (O_108,N_47119,N_48191);
and UO_109 (O_109,N_48742,N_48165);
nand UO_110 (O_110,N_49607,N_47803);
xor UO_111 (O_111,N_49704,N_48563);
xnor UO_112 (O_112,N_48722,N_48190);
xor UO_113 (O_113,N_46472,N_48879);
and UO_114 (O_114,N_46886,N_48581);
nor UO_115 (O_115,N_49176,N_48967);
nand UO_116 (O_116,N_46263,N_48119);
xnor UO_117 (O_117,N_48605,N_47628);
and UO_118 (O_118,N_47505,N_46921);
xnor UO_119 (O_119,N_49463,N_45493);
nand UO_120 (O_120,N_48176,N_48865);
and UO_121 (O_121,N_47149,N_49240);
or UO_122 (O_122,N_47583,N_49219);
nor UO_123 (O_123,N_49693,N_46749);
or UO_124 (O_124,N_46103,N_49098);
or UO_125 (O_125,N_47381,N_49133);
or UO_126 (O_126,N_45856,N_46646);
nor UO_127 (O_127,N_46815,N_46801);
xnor UO_128 (O_128,N_47644,N_45465);
nand UO_129 (O_129,N_47984,N_46007);
xor UO_130 (O_130,N_45872,N_47013);
and UO_131 (O_131,N_49477,N_46043);
and UO_132 (O_132,N_47240,N_45277);
xnor UO_133 (O_133,N_47258,N_49052);
nand UO_134 (O_134,N_49546,N_47629);
and UO_135 (O_135,N_46923,N_45015);
nand UO_136 (O_136,N_45954,N_47668);
nand UO_137 (O_137,N_45704,N_48345);
nor UO_138 (O_138,N_48792,N_46081);
and UO_139 (O_139,N_49798,N_45681);
nor UO_140 (O_140,N_46253,N_47363);
nor UO_141 (O_141,N_47401,N_45602);
or UO_142 (O_142,N_46453,N_47659);
xor UO_143 (O_143,N_48627,N_45905);
nor UO_144 (O_144,N_48151,N_45275);
nand UO_145 (O_145,N_48752,N_46348);
or UO_146 (O_146,N_46927,N_47546);
and UO_147 (O_147,N_48976,N_47503);
nand UO_148 (O_148,N_47774,N_46130);
or UO_149 (O_149,N_49030,N_48157);
nor UO_150 (O_150,N_46460,N_49605);
xnor UO_151 (O_151,N_47742,N_45668);
nor UO_152 (O_152,N_49327,N_48378);
or UO_153 (O_153,N_46033,N_47540);
or UO_154 (O_154,N_49408,N_46882);
nor UO_155 (O_155,N_46278,N_48618);
nor UO_156 (O_156,N_46559,N_47335);
or UO_157 (O_157,N_48774,N_49040);
nor UO_158 (O_158,N_49451,N_45051);
nand UO_159 (O_159,N_45412,N_48257);
or UO_160 (O_160,N_47901,N_46417);
and UO_161 (O_161,N_46346,N_48331);
and UO_162 (O_162,N_47528,N_49078);
and UO_163 (O_163,N_49370,N_47840);
and UO_164 (O_164,N_49387,N_46644);
and UO_165 (O_165,N_45618,N_48301);
nand UO_166 (O_166,N_49087,N_45407);
nor UO_167 (O_167,N_48540,N_49711);
nor UO_168 (O_168,N_45211,N_46655);
nand UO_169 (O_169,N_48608,N_45162);
or UO_170 (O_170,N_45208,N_46973);
nor UO_171 (O_171,N_48649,N_45846);
xnor UO_172 (O_172,N_49294,N_45816);
xor UO_173 (O_173,N_49550,N_45358);
and UO_174 (O_174,N_45770,N_47454);
xor UO_175 (O_175,N_48821,N_47975);
xor UO_176 (O_176,N_47338,N_45132);
xnor UO_177 (O_177,N_47812,N_47611);
xor UO_178 (O_178,N_48222,N_46438);
or UO_179 (O_179,N_45293,N_45559);
xnor UO_180 (O_180,N_47965,N_49129);
nand UO_181 (O_181,N_49498,N_45875);
nor UO_182 (O_182,N_48588,N_48254);
nand UO_183 (O_183,N_45121,N_49680);
nand UO_184 (O_184,N_48950,N_47506);
nand UO_185 (O_185,N_46011,N_48998);
and UO_186 (O_186,N_47971,N_47523);
and UO_187 (O_187,N_48679,N_48868);
or UO_188 (O_188,N_49088,N_48035);
nor UO_189 (O_189,N_45781,N_48951);
and UO_190 (O_190,N_49886,N_46537);
and UO_191 (O_191,N_47410,N_48286);
nor UO_192 (O_192,N_48969,N_48508);
xor UO_193 (O_193,N_45961,N_45361);
or UO_194 (O_194,N_47344,N_48349);
or UO_195 (O_195,N_47055,N_45930);
and UO_196 (O_196,N_49419,N_47063);
nand UO_197 (O_197,N_49231,N_45013);
nor UO_198 (O_198,N_45918,N_49629);
xor UO_199 (O_199,N_45832,N_49933);
nor UO_200 (O_200,N_49485,N_49271);
xor UO_201 (O_201,N_47167,N_48756);
xor UO_202 (O_202,N_48400,N_46547);
xor UO_203 (O_203,N_47004,N_47664);
or UO_204 (O_204,N_48802,N_45104);
nand UO_205 (O_205,N_47215,N_48136);
nand UO_206 (O_206,N_49927,N_47026);
and UO_207 (O_207,N_49162,N_45924);
and UO_208 (O_208,N_48037,N_46389);
and UO_209 (O_209,N_47478,N_45865);
and UO_210 (O_210,N_45145,N_47632);
nor UO_211 (O_211,N_49764,N_47423);
nor UO_212 (O_212,N_47077,N_47661);
nand UO_213 (O_213,N_47197,N_45159);
xor UO_214 (O_214,N_47655,N_45106);
and UO_215 (O_215,N_46311,N_45108);
or UO_216 (O_216,N_48700,N_49319);
xor UO_217 (O_217,N_45835,N_49807);
or UO_218 (O_218,N_46169,N_48996);
xor UO_219 (O_219,N_45000,N_48582);
nor UO_220 (O_220,N_48462,N_48720);
and UO_221 (O_221,N_49677,N_49665);
xnor UO_222 (O_222,N_49532,N_47067);
xor UO_223 (O_223,N_49867,N_46998);
nand UO_224 (O_224,N_49464,N_49203);
or UO_225 (O_225,N_46798,N_47574);
nand UO_226 (O_226,N_45799,N_49671);
or UO_227 (O_227,N_47373,N_47852);
nor UO_228 (O_228,N_47233,N_49931);
or UO_229 (O_229,N_47571,N_48303);
nor UO_230 (O_230,N_46915,N_45868);
nor UO_231 (O_231,N_49371,N_45887);
nor UO_232 (O_232,N_46667,N_48881);
and UO_233 (O_233,N_47166,N_45323);
xor UO_234 (O_234,N_46643,N_45263);
xor UO_235 (O_235,N_49997,N_45398);
nand UO_236 (O_236,N_47186,N_49590);
nor UO_237 (O_237,N_48428,N_47527);
and UO_238 (O_238,N_45966,N_46160);
nand UO_239 (O_239,N_46704,N_48994);
nand UO_240 (O_240,N_49462,N_46823);
nor UO_241 (O_241,N_45160,N_47616);
or UO_242 (O_242,N_47360,N_45045);
nor UO_243 (O_243,N_45584,N_48762);
xnor UO_244 (O_244,N_47558,N_46037);
xnor UO_245 (O_245,N_48768,N_49309);
or UO_246 (O_246,N_49668,N_47843);
nor UO_247 (O_247,N_45298,N_48084);
or UO_248 (O_248,N_48107,N_48818);
xor UO_249 (O_249,N_49819,N_46116);
nor UO_250 (O_250,N_47860,N_49122);
xor UO_251 (O_251,N_47205,N_45889);
nand UO_252 (O_252,N_45191,N_49942);
nand UO_253 (O_253,N_45152,N_45754);
or UO_254 (O_254,N_45579,N_48687);
nand UO_255 (O_255,N_46529,N_46757);
and UO_256 (O_256,N_47511,N_48528);
or UO_257 (O_257,N_46789,N_45527);
xnor UO_258 (O_258,N_47940,N_45699);
and UO_259 (O_259,N_48447,N_45333);
and UO_260 (O_260,N_49726,N_45128);
and UO_261 (O_261,N_48601,N_46899);
nand UO_262 (O_262,N_46034,N_46608);
or UO_263 (O_263,N_48043,N_49769);
and UO_264 (O_264,N_47873,N_49975);
nor UO_265 (O_265,N_47468,N_46156);
and UO_266 (O_266,N_49367,N_46561);
or UO_267 (O_267,N_49767,N_49476);
or UO_268 (O_268,N_46519,N_47985);
and UO_269 (O_269,N_48032,N_46423);
xnor UO_270 (O_270,N_48816,N_48755);
and UO_271 (O_271,N_47246,N_46216);
nand UO_272 (O_272,N_47919,N_47763);
and UO_273 (O_273,N_46360,N_49833);
nor UO_274 (O_274,N_49345,N_48744);
xor UO_275 (O_275,N_47064,N_45033);
xnor UO_276 (O_276,N_45055,N_47910);
nor UO_277 (O_277,N_46432,N_46732);
and UO_278 (O_278,N_45983,N_49232);
nand UO_279 (O_279,N_46082,N_45800);
and UO_280 (O_280,N_49046,N_46843);
and UO_281 (O_281,N_47966,N_45290);
and UO_282 (O_282,N_47248,N_46467);
nand UO_283 (O_283,N_49812,N_47184);
and UO_284 (O_284,N_49091,N_46351);
or UO_285 (O_285,N_47576,N_46852);
or UO_286 (O_286,N_45252,N_46416);
and UO_287 (O_287,N_48249,N_46215);
nor UO_288 (O_288,N_49457,N_49529);
nor UO_289 (O_289,N_46938,N_49175);
xor UO_290 (O_290,N_46891,N_49159);
nor UO_291 (O_291,N_46113,N_46495);
or UO_292 (O_292,N_45588,N_48164);
and UO_293 (O_293,N_46808,N_49706);
nor UO_294 (O_294,N_45625,N_46967);
xnor UO_295 (O_295,N_45314,N_47802);
xor UO_296 (O_296,N_48199,N_49329);
and UO_297 (O_297,N_46633,N_49672);
or UO_298 (O_298,N_46942,N_45603);
nor UO_299 (O_299,N_47932,N_48516);
and UO_300 (O_300,N_46377,N_47545);
nand UO_301 (O_301,N_47476,N_45388);
nor UO_302 (O_302,N_47025,N_49286);
nor UO_303 (O_303,N_48848,N_49244);
and UO_304 (O_304,N_45953,N_49109);
nor UO_305 (O_305,N_49452,N_46023);
nor UO_306 (O_306,N_46468,N_45083);
nand UO_307 (O_307,N_48510,N_45240);
nand UO_308 (O_308,N_48341,N_48148);
nor UO_309 (O_309,N_45081,N_49843);
or UO_310 (O_310,N_46730,N_47298);
xnor UO_311 (O_311,N_47181,N_47189);
xnor UO_312 (O_312,N_48645,N_49206);
or UO_313 (O_313,N_49701,N_46980);
or UO_314 (O_314,N_46750,N_45210);
nor UO_315 (O_315,N_45111,N_48584);
nand UO_316 (O_316,N_49699,N_46740);
or UO_317 (O_317,N_48898,N_49229);
nor UO_318 (O_318,N_47636,N_49382);
or UO_319 (O_319,N_45386,N_45510);
nand UO_320 (O_320,N_48395,N_46208);
xnor UO_321 (O_321,N_49888,N_46354);
nand UO_322 (O_322,N_45817,N_46479);
xnor UO_323 (O_323,N_45555,N_47660);
nor UO_324 (O_324,N_45620,N_48517);
and UO_325 (O_325,N_48657,N_47073);
nor UO_326 (O_326,N_48680,N_47885);
xor UO_327 (O_327,N_49377,N_49659);
nor UO_328 (O_328,N_49624,N_48172);
xor UO_329 (O_329,N_45171,N_45818);
xor UO_330 (O_330,N_48130,N_48860);
and UO_331 (O_331,N_48883,N_46012);
nor UO_332 (O_332,N_47829,N_47575);
or UO_333 (O_333,N_47471,N_49682);
or UO_334 (O_334,N_46577,N_47332);
or UO_335 (O_335,N_48867,N_48650);
xnor UO_336 (O_336,N_48210,N_46775);
and UO_337 (O_337,N_46609,N_49287);
and UO_338 (O_338,N_46447,N_48385);
xnor UO_339 (O_339,N_45755,N_48693);
and UO_340 (O_340,N_45543,N_47651);
and UO_341 (O_341,N_48068,N_49379);
and UO_342 (O_342,N_47156,N_45309);
and UO_343 (O_343,N_46990,N_49272);
or UO_344 (O_344,N_48390,N_49027);
xor UO_345 (O_345,N_46105,N_45080);
xor UO_346 (O_346,N_47775,N_49369);
nand UO_347 (O_347,N_46855,N_46501);
or UO_348 (O_348,N_49638,N_48009);
xor UO_349 (O_349,N_48134,N_49724);
nor UO_350 (O_350,N_47800,N_45140);
nand UO_351 (O_351,N_46489,N_46247);
nand UO_352 (O_352,N_49144,N_49691);
xor UO_353 (O_353,N_48217,N_48960);
nor UO_354 (O_354,N_47760,N_48067);
or UO_355 (O_355,N_45065,N_49401);
nor UO_356 (O_356,N_49864,N_49011);
and UO_357 (O_357,N_47663,N_49631);
or UO_358 (O_358,N_49822,N_47070);
xor UO_359 (O_359,N_48772,N_46958);
or UO_360 (O_360,N_47424,N_45392);
nand UO_361 (O_361,N_47749,N_48269);
or UO_362 (O_362,N_47261,N_47295);
and UO_363 (O_363,N_48205,N_49178);
xnor UO_364 (O_364,N_48023,N_47875);
nor UO_365 (O_365,N_46231,N_48681);
nand UO_366 (O_366,N_46087,N_46635);
nand UO_367 (O_367,N_46040,N_49879);
nor UO_368 (O_368,N_46875,N_45612);
or UO_369 (O_369,N_48285,N_48292);
nand UO_370 (O_370,N_45583,N_47779);
and UO_371 (O_371,N_48360,N_45423);
or UO_372 (O_372,N_49212,N_47493);
or UO_373 (O_373,N_45272,N_47758);
nor UO_374 (O_374,N_47255,N_46587);
and UO_375 (O_375,N_48850,N_49608);
xor UO_376 (O_376,N_47422,N_46019);
and UO_377 (O_377,N_48320,N_46797);
nand UO_378 (O_378,N_48271,N_47549);
xor UO_379 (O_379,N_48364,N_45726);
or UO_380 (O_380,N_47446,N_46122);
xor UO_381 (O_381,N_46904,N_45258);
and UO_382 (O_382,N_45267,N_49465);
nor UO_383 (O_383,N_45066,N_49891);
xnor UO_384 (O_384,N_45017,N_46123);
nor UO_385 (O_385,N_45435,N_49976);
nor UO_386 (O_386,N_49669,N_47770);
nand UO_387 (O_387,N_45560,N_48577);
and UO_388 (O_388,N_49270,N_45972);
xnor UO_389 (O_389,N_47087,N_45971);
nor UO_390 (O_390,N_47767,N_47526);
or UO_391 (O_391,N_46092,N_47135);
xnor UO_392 (O_392,N_48092,N_49071);
or UO_393 (O_393,N_47507,N_47447);
xnor UO_394 (O_394,N_49578,N_47751);
xnor UO_395 (O_395,N_49224,N_47415);
xnor UO_396 (O_396,N_46390,N_45326);
xor UO_397 (O_397,N_45179,N_49960);
nor UO_398 (O_398,N_49202,N_47286);
or UO_399 (O_399,N_46451,N_49458);
xnor UO_400 (O_400,N_47641,N_46415);
nor UO_401 (O_401,N_48115,N_48726);
xnor UO_402 (O_402,N_48159,N_45879);
or UO_403 (O_403,N_47420,N_48580);
nor UO_404 (O_404,N_46574,N_47701);
xor UO_405 (O_405,N_46992,N_46734);
or UO_406 (O_406,N_47345,N_48658);
or UO_407 (O_407,N_47865,N_49557);
xor UO_408 (O_408,N_48499,N_45069);
nor UO_409 (O_409,N_46521,N_47690);
xor UO_410 (O_410,N_47199,N_45387);
nor UO_411 (O_411,N_46373,N_49311);
xnor UO_412 (O_412,N_46814,N_45752);
nand UO_413 (O_413,N_46159,N_49447);
xor UO_414 (O_414,N_47109,N_49755);
or UO_415 (O_415,N_45890,N_45988);
or UO_416 (O_416,N_47480,N_49749);
or UO_417 (O_417,N_45268,N_47153);
and UO_418 (O_418,N_47715,N_45343);
xnor UO_419 (O_419,N_49047,N_45249);
nand UO_420 (O_420,N_49495,N_46020);
xnor UO_421 (O_421,N_48920,N_46365);
xor UO_422 (O_422,N_49574,N_46166);
nand UO_423 (O_423,N_49932,N_47144);
nor UO_424 (O_424,N_46975,N_45903);
nand UO_425 (O_425,N_46664,N_45531);
xnor UO_426 (O_426,N_45408,N_48990);
and UO_427 (O_427,N_46422,N_49180);
nor UO_428 (O_428,N_47236,N_45825);
or UO_429 (O_429,N_45195,N_46675);
nor UO_430 (O_430,N_47296,N_46319);
or UO_431 (O_431,N_46626,N_46421);
nor UO_432 (O_432,N_46112,N_47577);
or UO_433 (O_433,N_49014,N_49876);
nor UO_434 (O_434,N_46039,N_47250);
and UO_435 (O_435,N_46285,N_48195);
nor UO_436 (O_436,N_46703,N_48997);
nand UO_437 (O_437,N_45498,N_47557);
or UO_438 (O_438,N_49012,N_47483);
or UO_439 (O_439,N_48000,N_49086);
nand UO_440 (O_440,N_45740,N_48007);
or UO_441 (O_441,N_45606,N_45070);
nand UO_442 (O_442,N_46544,N_49784);
and UO_443 (O_443,N_49865,N_47902);
and UO_444 (O_444,N_45050,N_46956);
nor UO_445 (O_445,N_46579,N_49732);
and UO_446 (O_446,N_49762,N_49473);
or UO_447 (O_447,N_48057,N_45652);
nor UO_448 (O_448,N_45554,N_48328);
and UO_449 (O_449,N_45758,N_48667);
or UO_450 (O_450,N_46219,N_46984);
xor UO_451 (O_451,N_46017,N_48698);
xnor UO_452 (O_452,N_47081,N_46403);
nand UO_453 (O_453,N_49245,N_48519);
xnor UO_454 (O_454,N_48955,N_46476);
xor UO_455 (O_455,N_47850,N_45374);
or UO_456 (O_456,N_47169,N_47669);
xor UO_457 (O_457,N_45640,N_45469);
xor UO_458 (O_458,N_49552,N_48836);
nand UO_459 (O_459,N_49899,N_46086);
and UO_460 (O_460,N_46987,N_48216);
nor UO_461 (O_461,N_46430,N_46242);
or UO_462 (O_462,N_49907,N_47846);
and UO_463 (O_463,N_47457,N_49591);
xor UO_464 (O_464,N_47888,N_46518);
xor UO_465 (O_465,N_47137,N_47221);
xnor UO_466 (O_466,N_45657,N_48361);
xor UO_467 (O_467,N_49483,N_49497);
or UO_468 (O_468,N_47569,N_46539);
xor UO_469 (O_469,N_45040,N_47520);
or UO_470 (O_470,N_46210,N_46874);
or UO_471 (O_471,N_48895,N_45393);
or UO_472 (O_472,N_46934,N_46989);
or UO_473 (O_473,N_46362,N_49586);
xor UO_474 (O_474,N_46047,N_45206);
and UO_475 (O_475,N_46142,N_45960);
or UO_476 (O_476,N_48180,N_47445);
and UO_477 (O_477,N_45939,N_47175);
and UO_478 (O_478,N_45748,N_46356);
and UO_479 (O_479,N_45283,N_45250);
xnor UO_480 (O_480,N_47413,N_46716);
and UO_481 (O_481,N_49904,N_47470);
nand UO_482 (O_482,N_45824,N_47256);
nor UO_483 (O_483,N_49950,N_47808);
or UO_484 (O_484,N_47656,N_49655);
and UO_485 (O_485,N_49720,N_49869);
or UO_486 (O_486,N_45097,N_45837);
xnor UO_487 (O_487,N_49107,N_48372);
and UO_488 (O_488,N_47143,N_49601);
nand UO_489 (O_489,N_47716,N_45031);
and UO_490 (O_490,N_46446,N_46572);
nor UO_491 (O_491,N_45129,N_48131);
nor UO_492 (O_492,N_46725,N_46254);
nor UO_493 (O_493,N_48900,N_49005);
nand UO_494 (O_494,N_48471,N_45621);
nor UO_495 (O_495,N_49828,N_45474);
and UO_496 (O_496,N_45230,N_48690);
nor UO_497 (O_497,N_49835,N_49161);
or UO_498 (O_498,N_48399,N_49191);
nor UO_499 (O_499,N_45432,N_45379);
or UO_500 (O_500,N_46014,N_47322);
and UO_501 (O_501,N_48095,N_47667);
nand UO_502 (O_502,N_46056,N_49360);
nor UO_503 (O_503,N_47370,N_48160);
or UO_504 (O_504,N_48518,N_49525);
or UO_505 (O_505,N_46520,N_47497);
nor UO_506 (O_506,N_49799,N_46600);
nand UO_507 (O_507,N_49746,N_49563);
or UO_508 (O_508,N_45226,N_49208);
nor UO_509 (O_509,N_45234,N_49233);
xor UO_510 (O_510,N_47043,N_49028);
or UO_511 (O_511,N_45660,N_45369);
xnor UO_512 (O_512,N_48047,N_48121);
nand UO_513 (O_513,N_47041,N_47872);
nand UO_514 (O_514,N_46638,N_47533);
or UO_515 (O_515,N_47657,N_48593);
and UO_516 (O_516,N_47058,N_48504);
xor UO_517 (O_517,N_49643,N_48579);
or UO_518 (O_518,N_49410,N_48775);
or UO_519 (O_519,N_49708,N_49719);
and UO_520 (O_520,N_49790,N_48948);
nand UO_521 (O_521,N_49507,N_49102);
xor UO_522 (O_522,N_48093,N_48525);
nor UO_523 (O_523,N_47328,N_49895);
nand UO_524 (O_524,N_49909,N_47662);
nand UO_525 (O_525,N_46475,N_49467);
and UO_526 (O_526,N_46174,N_45428);
nand UO_527 (O_527,N_45430,N_46714);
nand UO_528 (O_528,N_46029,N_46293);
and UO_529 (O_529,N_45899,N_49003);
nand UO_530 (O_530,N_47402,N_49970);
nor UO_531 (O_531,N_48875,N_49275);
nor UO_532 (O_532,N_45476,N_47279);
or UO_533 (O_533,N_49069,N_48738);
or UO_534 (O_534,N_49744,N_48218);
and UO_535 (O_535,N_47986,N_47842);
nand UO_536 (O_536,N_47747,N_48851);
and UO_537 (O_537,N_47928,N_47272);
nor UO_538 (O_538,N_49308,N_48805);
xnor UO_539 (O_539,N_49280,N_47780);
or UO_540 (O_540,N_46257,N_46721);
or UO_541 (O_541,N_46756,N_48030);
xor UO_542 (O_542,N_47394,N_49778);
or UO_543 (O_543,N_45395,N_46532);
and UO_544 (O_544,N_46585,N_46106);
xnor UO_545 (O_545,N_45679,N_45994);
and UO_546 (O_546,N_48595,N_47148);
nor UO_547 (O_547,N_46076,N_48348);
xor UO_548 (O_548,N_45844,N_49277);
xor UO_549 (O_549,N_49313,N_47586);
nand UO_550 (O_550,N_47152,N_49676);
or UO_551 (O_551,N_46222,N_49956);
and UO_552 (O_552,N_49988,N_45772);
nand UO_553 (O_553,N_45076,N_46490);
or UO_554 (O_554,N_45406,N_47550);
or UO_555 (O_555,N_48114,N_46862);
nand UO_556 (O_556,N_47572,N_47693);
nand UO_557 (O_557,N_49592,N_46812);
or UO_558 (O_558,N_46653,N_48420);
nor UO_559 (O_559,N_46404,N_45482);
nand UO_560 (O_560,N_47040,N_48090);
nand UO_561 (O_561,N_46688,N_46299);
and UO_562 (O_562,N_47139,N_45542);
nor UO_563 (O_563,N_47640,N_46962);
nand UO_564 (O_564,N_46265,N_45764);
xor UO_565 (O_565,N_45237,N_45405);
or UO_566 (O_566,N_45949,N_45382);
and UO_567 (O_567,N_46760,N_45313);
nor UO_568 (O_568,N_48790,N_48337);
xnor UO_569 (O_569,N_49385,N_49281);
and UO_570 (O_570,N_45282,N_47229);
xnor UO_571 (O_571,N_49815,N_47822);
or UO_572 (O_572,N_49596,N_48660);
xor UO_573 (O_573,N_46845,N_49595);
nand UO_574 (O_574,N_45662,N_49860);
and UO_575 (O_575,N_49508,N_46338);
xor UO_576 (O_576,N_47213,N_48240);
or UO_577 (O_577,N_45470,N_48381);
nor UO_578 (O_578,N_46101,N_47125);
xnor UO_579 (O_579,N_45201,N_46584);
or UO_580 (O_580,N_48064,N_45370);
nand UO_581 (O_581,N_46900,N_48323);
nand UO_582 (O_582,N_46557,N_47930);
nor UO_583 (O_583,N_48437,N_49466);
and UO_584 (O_584,N_45673,N_46692);
xnor UO_585 (O_585,N_49058,N_46911);
or UO_586 (O_586,N_49796,N_47418);
nor UO_587 (O_587,N_48655,N_48904);
nor UO_588 (O_588,N_45485,N_46009);
or UO_589 (O_589,N_46323,N_47563);
nor UO_590 (O_590,N_49481,N_47357);
or UO_591 (O_591,N_46320,N_49236);
or UO_592 (O_592,N_49426,N_45709);
or UO_593 (O_593,N_46192,N_45677);
nor UO_594 (O_594,N_49214,N_48854);
nor UO_595 (O_595,N_45756,N_47553);
nand UO_596 (O_596,N_47383,N_47671);
nor UO_597 (O_597,N_47531,N_47359);
xor UO_598 (O_598,N_48346,N_45582);
nor UO_599 (O_599,N_48138,N_46712);
nand UO_600 (O_600,N_49543,N_45644);
nand UO_601 (O_601,N_48444,N_48873);
nor UO_602 (O_602,N_47091,N_47680);
nor UO_603 (O_603,N_46409,N_48945);
or UO_604 (O_604,N_47581,N_48123);
and UO_605 (O_605,N_48666,N_49140);
or UO_606 (O_606,N_47564,N_48279);
nor UO_607 (O_607,N_47377,N_49670);
and UO_608 (O_608,N_47959,N_47739);
nand UO_609 (O_609,N_49570,N_47477);
xnor UO_610 (O_610,N_49906,N_47356);
or UO_611 (O_611,N_48938,N_46380);
nand UO_612 (O_612,N_45888,N_45224);
or UO_613 (O_613,N_48953,N_48747);
nor UO_614 (O_614,N_47915,N_46541);
nand UO_615 (O_615,N_49025,N_48273);
or UO_616 (O_616,N_49217,N_49339);
and UO_617 (O_617,N_45281,N_49567);
and UO_618 (O_618,N_49681,N_48838);
xnor UO_619 (O_619,N_46689,N_46545);
and UO_620 (O_620,N_48758,N_46059);
or UO_621 (O_621,N_47890,N_45154);
nor UO_622 (O_622,N_48793,N_45340);
nand UO_623 (O_623,N_49442,N_49577);
nand UO_624 (O_624,N_46259,N_48745);
nor UO_625 (O_625,N_46399,N_45882);
nor UO_626 (O_626,N_45401,N_49938);
xor UO_627 (O_627,N_47542,N_47287);
nor UO_628 (O_628,N_48175,N_49667);
nand UO_629 (O_629,N_48470,N_46168);
or UO_630 (O_630,N_48184,N_48226);
nand UO_631 (O_631,N_45347,N_47990);
nand UO_632 (O_632,N_46546,N_47967);
or UO_633 (O_633,N_45658,N_48644);
or UO_634 (O_634,N_46710,N_49320);
xor UO_635 (O_635,N_45384,N_48209);
nor UO_636 (O_636,N_49002,N_45315);
nor UO_637 (O_637,N_48211,N_45355);
xnor UO_638 (O_638,N_49428,N_47886);
and UO_639 (O_639,N_47974,N_49874);
nand UO_640 (O_640,N_47014,N_47052);
xor UO_641 (O_641,N_46940,N_49171);
nand UO_642 (O_642,N_49664,N_47088);
nand UO_643 (O_643,N_46069,N_48734);
xnor UO_644 (O_644,N_47227,N_49612);
nand UO_645 (O_645,N_48677,N_49770);
nor UO_646 (O_646,N_46950,N_49641);
nand UO_647 (O_647,N_48619,N_49186);
and UO_648 (O_648,N_45763,N_47309);
or UO_649 (O_649,N_49760,N_47766);
xor UO_650 (O_650,N_45849,N_47687);
nor UO_651 (O_651,N_47254,N_49696);
nand UO_652 (O_652,N_47953,N_49534);
nand UO_653 (O_653,N_49269,N_45264);
nand UO_654 (O_654,N_47582,N_49658);
or UO_655 (O_655,N_45829,N_48646);
nor UO_656 (O_656,N_48193,N_47686);
xnor UO_657 (O_657,N_47231,N_46287);
nand UO_658 (O_658,N_48607,N_45135);
and UO_659 (O_659,N_46937,N_48459);
nor UO_660 (O_660,N_49929,N_45701);
nand UO_661 (O_661,N_48099,N_48668);
or UO_662 (O_662,N_49341,N_46838);
and UO_663 (O_663,N_49568,N_47201);
nand UO_664 (O_664,N_48636,N_45808);
xnor UO_665 (O_665,N_49153,N_47620);
and UO_666 (O_666,N_49620,N_46129);
nor UO_667 (O_667,N_45523,N_48116);
or UO_668 (O_668,N_49008,N_45847);
xnor UO_669 (O_669,N_47753,N_46488);
xnor UO_670 (O_670,N_45306,N_46121);
and UO_671 (O_671,N_47407,N_49922);
nor UO_672 (O_672,N_45710,N_45500);
nand UO_673 (O_673,N_46702,N_49775);
and UO_674 (O_674,N_46255,N_47913);
nand UO_675 (O_675,N_48600,N_46742);
xor UO_676 (O_676,N_46500,N_45481);
nor UO_677 (O_677,N_47823,N_47978);
xnor UO_678 (O_678,N_49963,N_48319);
or UO_679 (O_679,N_46593,N_45515);
nor UO_680 (O_680,N_49861,N_45591);
or UO_681 (O_681,N_46487,N_45628);
xnor UO_682 (O_682,N_45327,N_48351);
or UO_683 (O_683,N_48526,N_45937);
nand UO_684 (O_684,N_46469,N_48086);
xnor UO_685 (O_685,N_49220,N_47012);
or UO_686 (O_686,N_45341,N_45114);
nand UO_687 (O_687,N_46117,N_47515);
xor UO_688 (O_688,N_49494,N_46084);
and UO_689 (O_689,N_48242,N_48102);
xor UO_690 (O_690,N_49991,N_45149);
or UO_691 (O_691,N_46340,N_48731);
or UO_692 (O_692,N_47994,N_45077);
nand UO_693 (O_693,N_46918,N_47353);
nand UO_694 (O_694,N_46554,N_46819);
nand UO_695 (O_695,N_46223,N_48819);
xnor UO_696 (O_696,N_48880,N_45993);
xnor UO_697 (O_697,N_49593,N_45363);
and UO_698 (O_698,N_49780,N_45936);
xor UO_699 (O_699,N_46393,N_49943);
xor UO_700 (O_700,N_49150,N_48568);
or UO_701 (O_701,N_45675,N_49587);
xor UO_702 (O_702,N_45276,N_45850);
nand UO_703 (O_703,N_45203,N_47720);
or UO_704 (O_704,N_46442,N_46769);
and UO_705 (O_705,N_46758,N_49163);
or UO_706 (O_706,N_45916,N_46914);
nand UO_707 (O_707,N_46787,N_46235);
or UO_708 (O_708,N_45209,N_48350);
xnor UO_709 (O_709,N_47670,N_49980);
and UO_710 (O_710,N_46277,N_45192);
nand UO_711 (O_711,N_47519,N_45062);
xnor UO_712 (O_712,N_45116,N_49703);
and UO_713 (O_713,N_49527,N_45525);
nor UO_714 (O_714,N_49842,N_49189);
nor UO_715 (O_715,N_45426,N_45797);
nor UO_716 (O_716,N_49730,N_46443);
nand UO_717 (O_717,N_46549,N_45042);
or UO_718 (O_718,N_47247,N_46182);
or UO_719 (O_719,N_46063,N_46376);
or UO_720 (O_720,N_45325,N_47449);
nand UO_721 (O_721,N_48080,N_49035);
and UO_722 (O_722,N_48925,N_48808);
nand UO_723 (O_723,N_47997,N_46234);
and UO_724 (O_724,N_45086,N_49136);
xnor UO_725 (O_725,N_49256,N_48622);
xnor UO_726 (O_726,N_49600,N_49615);
and UO_727 (O_727,N_47881,N_45339);
nand UO_728 (O_728,N_49118,N_45198);
nor UO_729 (O_729,N_45505,N_48485);
nand UO_730 (O_730,N_48737,N_48377);
nand UO_731 (O_731,N_49714,N_46031);
nand UO_732 (O_732,N_45848,N_47551);
xnor UO_733 (O_733,N_49413,N_47128);
xor UO_734 (O_734,N_48304,N_46358);
nor UO_735 (O_735,N_49310,N_48307);
nor UO_736 (O_736,N_45010,N_49785);
or UO_737 (O_737,N_46883,N_48652);
or UO_738 (O_738,N_45833,N_49689);
and UO_739 (O_739,N_48829,N_45109);
or UO_740 (O_740,N_49813,N_47441);
xnor UO_741 (O_741,N_45459,N_45036);
xor UO_742 (O_742,N_48458,N_48497);
nor UO_743 (O_743,N_45095,N_48430);
nand UO_744 (O_744,N_49556,N_45992);
nand UO_745 (O_745,N_48703,N_48691);
and UO_746 (O_746,N_45057,N_46669);
or UO_747 (O_747,N_45826,N_47498);
nor UO_748 (O_748,N_49104,N_49374);
nand UO_749 (O_749,N_49353,N_47815);
nand UO_750 (O_750,N_48450,N_45762);
xor UO_751 (O_751,N_49292,N_47727);
or UO_752 (O_752,N_46919,N_47474);
and UO_753 (O_753,N_48861,N_48983);
nand UO_754 (O_754,N_46666,N_49119);
xnor UO_755 (O_755,N_49438,N_49258);
or UO_756 (O_756,N_48486,N_45659);
or UO_757 (O_757,N_49143,N_49375);
xor UO_758 (O_758,N_45626,N_47740);
and UO_759 (O_759,N_45039,N_46912);
or UO_760 (O_760,N_47337,N_48743);
nand UO_761 (O_761,N_45273,N_46289);
nand UO_762 (O_762,N_45118,N_46848);
nand UO_763 (O_763,N_49554,N_45143);
or UO_764 (O_764,N_46970,N_48357);
nor UO_765 (O_765,N_49998,N_46639);
xnor UO_766 (O_766,N_48477,N_49170);
and UO_767 (O_767,N_46602,N_47625);
or UO_768 (O_768,N_48042,N_46425);
xnor UO_769 (O_769,N_47834,N_49616);
or UO_770 (O_770,N_45213,N_45773);
nor UO_771 (O_771,N_47428,N_45750);
and UO_772 (O_772,N_48606,N_46394);
and UO_773 (O_773,N_47379,N_49606);
nor UO_774 (O_774,N_45845,N_46284);
or UO_775 (O_775,N_46748,N_49576);
nor UO_776 (O_776,N_45739,N_45167);
and UO_777 (O_777,N_47757,N_48038);
or UO_778 (O_778,N_47425,N_48529);
nor UO_779 (O_779,N_45862,N_48617);
and UO_780 (O_780,N_48708,N_46582);
xor UO_781 (O_781,N_49694,N_47826);
or UO_782 (O_782,N_49725,N_49300);
nand UO_783 (O_783,N_48203,N_49977);
nand UO_784 (O_784,N_46690,N_45457);
xor UO_785 (O_785,N_45180,N_48126);
or UO_786 (O_786,N_46194,N_48817);
nor UO_787 (O_787,N_48375,N_47317);
and UO_788 (O_788,N_49894,N_48940);
xor UO_789 (O_789,N_45043,N_48952);
nand UO_790 (O_790,N_49722,N_49248);
xor UO_791 (O_791,N_45418,N_46462);
nand UO_792 (O_792,N_45778,N_49034);
xnor UO_793 (O_793,N_46203,N_48110);
or UO_794 (O_794,N_48389,N_46673);
nand UO_795 (O_795,N_47102,N_48986);
nand UO_796 (O_796,N_48327,N_45134);
or UO_797 (O_797,N_45391,N_49283);
nand UO_798 (O_798,N_49290,N_49851);
nor UO_799 (O_799,N_47191,N_49342);
nand UO_800 (O_800,N_49805,N_48501);
nand UO_801 (O_801,N_46830,N_45454);
xor UO_802 (O_802,N_45574,N_49912);
xnor UO_803 (O_803,N_49644,N_48166);
nor UO_804 (O_804,N_48844,N_47643);
xor UO_805 (O_805,N_45239,N_45383);
and UO_806 (O_806,N_49887,N_46661);
nand UO_807 (O_807,N_47340,N_49397);
and UO_808 (O_808,N_46353,N_47608);
or UO_809 (O_809,N_47123,N_49539);
nor UO_810 (O_810,N_47744,N_48778);
or UO_811 (O_811,N_47606,N_49246);
and UO_812 (O_812,N_47274,N_47811);
or UO_813 (O_813,N_49505,N_49145);
or UO_814 (O_814,N_45979,N_49520);
nand UO_815 (O_815,N_48025,N_49128);
xor UO_816 (O_816,N_46176,N_48621);
nor UO_817 (O_817,N_48481,N_48402);
nor UO_818 (O_818,N_48270,N_46836);
nand UO_819 (O_819,N_45068,N_49820);
or UO_820 (O_820,N_47912,N_48724);
nand UO_821 (O_821,N_47906,N_49192);
nor UO_822 (O_822,N_46097,N_45502);
xor UO_823 (O_823,N_47934,N_46445);
nand UO_824 (O_824,N_47729,N_45587);
xor UO_825 (O_825,N_46663,N_45987);
xor UO_826 (O_826,N_47140,N_48368);
xor UO_827 (O_827,N_45099,N_49424);
xnor UO_828 (O_828,N_49019,N_46003);
and UO_829 (O_829,N_49692,N_45223);
xnor UO_830 (O_830,N_48449,N_49503);
nand UO_831 (O_831,N_48957,N_46000);
or UO_832 (O_832,N_45705,N_46152);
nand UO_833 (O_833,N_47522,N_47555);
and UO_834 (O_834,N_47979,N_47399);
xor UO_835 (O_835,N_46601,N_46846);
nor UO_836 (O_836,N_49871,N_48489);
xor UO_837 (O_837,N_48147,N_45260);
nor UO_838 (O_838,N_48834,N_46024);
xnor UO_839 (O_839,N_46636,N_45938);
or UO_840 (O_840,N_48142,N_47388);
and UO_841 (O_841,N_47647,N_47777);
or UO_842 (O_842,N_47570,N_46155);
or UO_843 (O_843,N_47391,N_47068);
nor UO_844 (O_844,N_49197,N_47285);
nand UO_845 (O_845,N_47341,N_48961);
xor UO_846 (O_846,N_48045,N_49121);
nor UO_847 (O_847,N_45442,N_46150);
and UO_848 (O_848,N_49468,N_45419);
and UO_849 (O_849,N_45958,N_48753);
nand UO_850 (O_850,N_49531,N_45170);
nor UO_851 (O_851,N_49023,N_46622);
or UO_852 (O_852,N_47327,N_45049);
xnor UO_853 (O_853,N_45422,N_46183);
and UO_854 (O_854,N_47726,N_47385);
nand UO_855 (O_855,N_49152,N_45274);
xnor UO_856 (O_856,N_45751,N_49551);
xor UO_857 (O_857,N_46719,N_45048);
xor UO_858 (O_858,N_49840,N_46157);
and UO_859 (O_859,N_48974,N_46485);
nand UO_860 (O_860,N_48964,N_45804);
nor UO_861 (O_861,N_46905,N_48293);
nor UO_862 (O_862,N_49808,N_46041);
xor UO_863 (O_863,N_45877,N_47034);
nor UO_864 (O_864,N_46509,N_47639);
xor UO_865 (O_865,N_45692,N_45607);
and UO_866 (O_866,N_49999,N_46534);
nor UO_867 (O_867,N_49969,N_48418);
xor UO_868 (O_868,N_47300,N_46943);
xnor UO_869 (O_869,N_45511,N_48306);
or UO_870 (O_870,N_49130,N_45749);
xnor UO_871 (O_871,N_48822,N_45572);
nand UO_872 (O_872,N_47354,N_46527);
or UO_873 (O_873,N_48312,N_45975);
nor UO_874 (O_874,N_47560,N_49289);
xnor UO_875 (O_875,N_47404,N_49893);
or UO_876 (O_876,N_49801,N_46514);
and UO_877 (O_877,N_47126,N_47121);
xor UO_878 (O_878,N_45445,N_47466);
or UO_879 (O_879,N_49490,N_46779);
xnor UO_880 (O_880,N_48542,N_45881);
xor UO_881 (O_881,N_47330,N_46456);
nor UO_882 (O_882,N_46352,N_46745);
xnor UO_883 (O_883,N_46543,N_46523);
nor UO_884 (O_884,N_45651,N_48576);
and UO_885 (O_885,N_46275,N_47408);
or UO_886 (O_886,N_45544,N_48642);
or UO_887 (O_887,N_49017,N_45464);
xor UO_888 (O_888,N_46162,N_46115);
xnor UO_889 (O_889,N_48069,N_47830);
xnor UO_890 (O_890,N_49181,N_48663);
nand UO_891 (O_891,N_48427,N_49910);
nor UO_892 (O_892,N_47938,N_49123);
and UO_893 (O_893,N_49838,N_47926);
nor UO_894 (O_894,N_45655,N_49340);
and UO_895 (O_895,N_49745,N_48932);
and UO_896 (O_896,N_48049,N_48721);
and UO_897 (O_897,N_48740,N_49182);
and UO_898 (O_898,N_48122,N_45564);
and UO_899 (O_899,N_49890,N_46735);
and UO_900 (O_900,N_48927,N_45110);
nor UO_901 (O_901,N_45506,N_47187);
nor UO_902 (O_902,N_47532,N_48572);
nand UO_903 (O_903,N_47079,N_46681);
nor UO_904 (O_904,N_49433,N_48264);
and UO_905 (O_905,N_48917,N_45366);
or UO_906 (O_906,N_49349,N_49302);
nand UO_907 (O_907,N_48243,N_46371);
nand UO_908 (O_908,N_48761,N_46066);
and UO_909 (O_909,N_49254,N_49402);
nand UO_910 (O_910,N_49789,N_49831);
nor UO_911 (O_911,N_46733,N_47492);
nand UO_912 (O_912,N_49914,N_49583);
nand UO_913 (O_913,N_48376,N_46511);
nand UO_914 (O_914,N_47429,N_47384);
nand UO_915 (O_915,N_47475,N_46890);
xnor UO_916 (O_916,N_49687,N_45927);
and UO_917 (O_917,N_45831,N_47618);
xnor UO_918 (O_918,N_48592,N_47621);
or UO_919 (O_919,N_47214,N_49200);
xnor UO_920 (O_920,N_48214,N_48441);
nand UO_921 (O_921,N_47989,N_45838);
xnor UO_922 (O_922,N_47100,N_47366);
nand UO_923 (O_923,N_47460,N_46310);
nor UO_924 (O_924,N_45472,N_46075);
nand UO_925 (O_925,N_45338,N_49051);
nor UO_926 (O_926,N_49516,N_47485);
and UO_927 (O_927,N_49721,N_48251);
or UO_928 (O_928,N_47697,N_48911);
and UO_929 (O_929,N_48422,N_49449);
nand UO_930 (O_930,N_48678,N_49555);
nand UO_931 (O_931,N_47018,N_49653);
nor UO_932 (O_932,N_45664,N_46676);
and UO_933 (O_933,N_49062,N_47361);
and UO_934 (O_934,N_47369,N_45516);
xor UO_935 (O_935,N_47386,N_46195);
nand UO_936 (O_936,N_47469,N_49544);
nand UO_937 (O_937,N_48594,N_47462);
and UO_938 (O_938,N_49810,N_48559);
or UO_939 (O_939,N_47095,N_49511);
or UO_940 (O_940,N_47922,N_45030);
and UO_941 (O_941,N_45745,N_45700);
nand UO_942 (O_942,N_45551,N_45598);
nor UO_943 (O_943,N_47032,N_49729);
or UO_944 (O_944,N_45627,N_49038);
nor UO_945 (O_945,N_49391,N_46482);
and UO_946 (O_946,N_48914,N_49561);
nand UO_947 (O_947,N_49753,N_49480);
and UO_948 (O_948,N_49120,N_48135);
nand UO_949 (O_949,N_48603,N_45299);
and UO_950 (O_950,N_45873,N_48874);
nor UO_951 (O_951,N_46724,N_46969);
and UO_952 (O_952,N_45530,N_46078);
nor UO_953 (O_953,N_47795,N_45851);
or UO_954 (O_954,N_45577,N_47992);
and UO_955 (O_955,N_45715,N_47183);
and UO_956 (O_956,N_45814,N_45702);
xnor UO_957 (O_957,N_47939,N_47331);
xnor UO_958 (O_958,N_46810,N_48704);
nor UO_959 (O_959,N_49004,N_46272);
or UO_960 (O_960,N_49710,N_45788);
nand UO_961 (O_961,N_45321,N_46806);
and UO_962 (O_962,N_46941,N_48455);
nand UO_963 (O_963,N_45084,N_49418);
xnor UO_964 (O_964,N_48739,N_48767);
and UO_965 (O_965,N_47949,N_49709);
xnor UO_966 (O_966,N_46931,N_48044);
xnor UO_967 (O_967,N_46857,N_46983);
or UO_968 (O_968,N_46098,N_47299);
nand UO_969 (O_969,N_47244,N_48003);
nand UO_970 (O_970,N_46189,N_49947);
or UO_971 (O_971,N_47239,N_47712);
xor UO_972 (O_972,N_45016,N_49662);
xor UO_973 (O_973,N_48864,N_49930);
or UO_974 (O_974,N_49089,N_47268);
or UO_975 (O_975,N_49599,N_48004);
xnor UO_976 (O_976,N_45278,N_48589);
and UO_977 (O_977,N_47482,N_49352);
nor UO_978 (O_978,N_49460,N_47150);
nand UO_979 (O_979,N_48412,N_48682);
and UO_980 (O_980,N_48954,N_46791);
or UO_981 (O_981,N_47008,N_49378);
nand UO_982 (O_982,N_48435,N_46677);
nor UO_983 (O_983,N_47151,N_47916);
nor UO_984 (O_984,N_45279,N_46872);
nand UO_985 (O_985,N_45054,N_48479);
nor UO_986 (O_986,N_46698,N_47734);
nor UO_987 (O_987,N_45189,N_45489);
nand UO_988 (O_988,N_49618,N_46433);
and UO_989 (O_989,N_48672,N_47578);
nand UO_990 (O_990,N_47325,N_46286);
xor UO_991 (O_991,N_46236,N_47884);
and UO_992 (O_992,N_48671,N_49565);
and UO_993 (O_993,N_47987,N_45586);
nand UO_994 (O_994,N_47082,N_47623);
and UO_995 (O_995,N_48661,N_45741);
nand UO_996 (O_996,N_49761,N_47339);
and UO_997 (O_997,N_45215,N_46615);
nor UO_998 (O_998,N_46540,N_45533);
nand UO_999 (O_999,N_46834,N_47275);
nand UO_1000 (O_1000,N_45999,N_49858);
nand UO_1001 (O_1001,N_46065,N_47057);
and UO_1002 (O_1002,N_49082,N_47453);
nor UO_1003 (O_1003,N_46792,N_46367);
nor UO_1004 (O_1004,N_48274,N_48830);
nand UO_1005 (O_1005,N_48062,N_48033);
nor UO_1006 (O_1006,N_47103,N_48723);
xor UO_1007 (O_1007,N_49844,N_47029);
xnor UO_1008 (O_1008,N_46720,N_48553);
and UO_1009 (O_1009,N_47784,N_48615);
nor UO_1010 (O_1010,N_45235,N_46463);
nor UO_1011 (O_1011,N_48206,N_46932);
or UO_1012 (O_1012,N_46308,N_48196);
and UO_1013 (O_1013,N_46385,N_49727);
nand UO_1014 (O_1014,N_48230,N_48426);
and UO_1015 (O_1015,N_49148,N_45410);
or UO_1016 (O_1016,N_48735,N_47573);
and UO_1017 (O_1017,N_46339,N_49368);
nand UO_1018 (O_1018,N_46111,N_48496);
nand UO_1019 (O_1019,N_49614,N_49619);
or UO_1020 (O_1020,N_48669,N_49794);
xor UO_1021 (O_1021,N_46640,N_45959);
nor UO_1022 (O_1022,N_46863,N_45475);
nand UO_1023 (O_1023,N_45220,N_47305);
xor UO_1024 (O_1024,N_49959,N_45075);
or UO_1025 (O_1025,N_49184,N_47847);
and UO_1026 (O_1026,N_45897,N_47134);
or UO_1027 (O_1027,N_47877,N_48109);
and UO_1028 (O_1028,N_49771,N_45375);
or UO_1029 (O_1029,N_49666,N_48783);
and UO_1030 (O_1030,N_47541,N_45287);
nand UO_1031 (O_1031,N_46759,N_48919);
xor UO_1032 (O_1032,N_48310,N_48053);
or UO_1033 (O_1033,N_48771,N_48736);
nor UO_1034 (O_1034,N_48260,N_47465);
or UO_1035 (O_1035,N_48995,N_45981);
nand UO_1036 (O_1036,N_45720,N_48054);
nand UO_1037 (O_1037,N_47867,N_47301);
or UO_1038 (O_1038,N_48842,N_47234);
and UO_1039 (O_1039,N_47798,N_45161);
or UO_1040 (O_1040,N_49255,N_45060);
nand UO_1041 (O_1041,N_49390,N_46127);
xnor UO_1042 (O_1042,N_49954,N_48877);
xnor UO_1043 (O_1043,N_48647,N_46616);
nand UO_1044 (O_1044,N_48469,N_46407);
or UO_1045 (O_1045,N_47718,N_46578);
nand UO_1046 (O_1046,N_46093,N_46091);
and UO_1047 (O_1047,N_47273,N_47849);
nand UO_1048 (O_1048,N_47645,N_45318);
and UO_1049 (O_1049,N_48562,N_46972);
or UO_1050 (O_1050,N_47635,N_47367);
and UO_1051 (O_1051,N_49634,N_47048);
nand UO_1052 (O_1052,N_47521,N_48567);
and UO_1053 (O_1053,N_48336,N_49553);
and UO_1054 (O_1054,N_47136,N_49853);
nor UO_1055 (O_1055,N_46876,N_49399);
xnor UO_1056 (O_1056,N_49384,N_49882);
nand UO_1057 (O_1057,N_45009,N_46273);
and UO_1058 (O_1058,N_47765,N_47098);
xor UO_1059 (O_1059,N_45184,N_46441);
or UO_1060 (O_1060,N_48280,N_45513);
or UO_1061 (O_1061,N_46851,N_49242);
nor UO_1062 (O_1062,N_48773,N_46957);
nand UO_1063 (O_1063,N_48728,N_46207);
and UO_1064 (O_1064,N_46729,N_47595);
and UO_1065 (O_1065,N_47703,N_45216);
or UO_1066 (O_1066,N_45747,N_45920);
or UO_1067 (O_1067,N_48706,N_49781);
or UO_1068 (O_1068,N_46755,N_48169);
nand UO_1069 (O_1069,N_48597,N_49830);
or UO_1070 (O_1070,N_45012,N_45508);
nand UO_1071 (O_1071,N_45779,N_48149);
or UO_1072 (O_1072,N_49821,N_47878);
or UO_1073 (O_1073,N_48776,N_45915);
or UO_1074 (O_1074,N_46457,N_45487);
and UO_1075 (O_1075,N_48174,N_47265);
nor UO_1076 (O_1076,N_45534,N_47138);
nand UO_1077 (O_1077,N_45867,N_46619);
nand UO_1078 (O_1078,N_47209,N_49228);
xor UO_1079 (O_1079,N_47817,N_45046);
and UO_1080 (O_1080,N_48334,N_46313);
nand UO_1081 (O_1081,N_48490,N_46590);
nand UO_1082 (O_1082,N_48639,N_48855);
nand UO_1083 (O_1083,N_48168,N_45221);
or UO_1084 (O_1084,N_49572,N_47937);
xor UO_1085 (O_1085,N_47945,N_47688);
nor UO_1086 (O_1086,N_46553,N_48267);
nor UO_1087 (O_1087,N_46387,N_47731);
nor UO_1088 (O_1088,N_49403,N_46350);
nand UO_1089 (O_1089,N_45218,N_47212);
and UO_1090 (O_1090,N_46592,N_47270);
nand UO_1091 (O_1091,N_45674,N_48362);
nand UO_1092 (O_1092,N_49962,N_45261);
nor UO_1093 (O_1093,N_47190,N_48931);
and UO_1094 (O_1094,N_47622,N_48185);
or UO_1095 (O_1095,N_46172,N_47101);
nor UO_1096 (O_1096,N_46525,N_45717);
or UO_1097 (O_1097,N_48059,N_46778);
nor UO_1098 (O_1098,N_49448,N_48370);
and UO_1099 (O_1099,N_47044,N_46107);
or UO_1100 (O_1100,N_48315,N_46683);
or UO_1101 (O_1101,N_46470,N_49383);
or UO_1102 (O_1102,N_46392,N_47887);
and UO_1103 (O_1103,N_45319,N_45089);
nor UO_1104 (O_1104,N_49646,N_45307);
and UO_1105 (O_1105,N_46408,N_46109);
nand UO_1106 (O_1106,N_46861,N_45127);
xnor UO_1107 (O_1107,N_48814,N_47010);
nor UO_1108 (O_1108,N_45150,N_48662);
and UO_1109 (O_1109,N_48132,N_47450);
nor UO_1110 (O_1110,N_46971,N_47781);
nand UO_1111 (O_1111,N_49636,N_45904);
xor UO_1112 (O_1112,N_46612,N_46839);
and UO_1113 (O_1113,N_49774,N_45694);
or UO_1114 (O_1114,N_46498,N_49488);
and UO_1115 (O_1115,N_48784,N_48125);
or UO_1116 (O_1116,N_49562,N_49836);
and UO_1117 (O_1117,N_45597,N_45289);
xor UO_1118 (O_1118,N_48096,N_47241);
and UO_1119 (O_1119,N_47479,N_46952);
xnor UO_1120 (O_1120,N_48746,N_48150);
and UO_1121 (O_1121,N_46524,N_48548);
or UO_1122 (O_1122,N_49589,N_46149);
and UO_1123 (O_1123,N_46151,N_48807);
nor UO_1124 (O_1124,N_45738,N_49199);
xor UO_1125 (O_1125,N_48417,N_45035);
xnor UO_1126 (O_1126,N_47333,N_47263);
nand UO_1127 (O_1127,N_49972,N_49902);
or UO_1128 (O_1128,N_46916,N_46312);
xor UO_1129 (O_1129,N_47145,N_46821);
or UO_1130 (O_1130,N_45871,N_49700);
and UO_1131 (O_1131,N_48962,N_45478);
and UO_1132 (O_1132,N_49273,N_46492);
and UO_1133 (O_1133,N_45665,N_49039);
or UO_1134 (O_1134,N_47813,N_46700);
nor UO_1135 (O_1135,N_48332,N_46629);
nor UO_1136 (O_1136,N_49847,N_46435);
xor UO_1137 (O_1137,N_46910,N_46064);
nand UO_1138 (O_1138,N_49454,N_45854);
nand UO_1139 (O_1139,N_47440,N_45908);
xor UO_1140 (O_1140,N_46204,N_45310);
nor UO_1141 (O_1141,N_47490,N_46978);
or UO_1142 (O_1142,N_45328,N_47372);
nor UO_1143 (O_1143,N_48513,N_48101);
nand UO_1144 (O_1144,N_47605,N_47921);
or UO_1145 (O_1145,N_46507,N_47117);
and UO_1146 (O_1146,N_46331,N_48295);
xor UO_1147 (O_1147,N_48330,N_46238);
or UO_1148 (O_1148,N_47351,N_48365);
and UO_1149 (O_1149,N_47060,N_45139);
or UO_1150 (O_1150,N_46762,N_49445);
nor UO_1151 (O_1151,N_48146,N_46173);
or UO_1152 (O_1152,N_47962,N_49491);
or UO_1153 (O_1153,N_47192,N_48973);
or UO_1154 (O_1154,N_45795,N_47019);
xnor UO_1155 (O_1155,N_48673,N_47179);
or UO_1156 (O_1156,N_47027,N_48749);
nand UO_1157 (O_1157,N_48788,N_45085);
xor UO_1158 (O_1158,N_46928,N_47304);
and UO_1159 (O_1159,N_45656,N_45518);
and UO_1160 (O_1160,N_49983,N_47868);
xnor UO_1161 (O_1161,N_46877,N_46016);
nor UO_1162 (O_1162,N_49239,N_46229);
and UO_1163 (O_1163,N_46997,N_48113);
or UO_1164 (O_1164,N_47110,N_45957);
or UO_1165 (O_1165,N_46008,N_45807);
xor UO_1166 (O_1166,N_47896,N_47160);
nand UO_1167 (O_1167,N_49955,N_49074);
or UO_1168 (O_1168,N_48558,N_45222);
or UO_1169 (O_1169,N_49101,N_45545);
or UO_1170 (O_1170,N_45593,N_45302);
and UO_1171 (O_1171,N_49226,N_45661);
nor UO_1172 (O_1172,N_49337,N_46542);
nor UO_1173 (O_1173,N_45933,N_48899);
xor UO_1174 (O_1174,N_46771,N_45914);
or UO_1175 (O_1175,N_47282,N_45732);
or UO_1176 (O_1176,N_46906,N_49733);
xnor UO_1177 (O_1177,N_45984,N_47649);
and UO_1178 (O_1178,N_49358,N_48702);
xnor UO_1179 (O_1179,N_49373,N_49325);
or UO_1180 (O_1180,N_46668,N_48034);
or UO_1181 (O_1181,N_48841,N_49407);
nor UO_1182 (O_1182,N_48394,N_48401);
nor UO_1183 (O_1183,N_45725,N_45943);
nand UO_1184 (O_1184,N_46650,N_45156);
xor UO_1185 (O_1185,N_46177,N_49137);
nand UO_1186 (O_1186,N_47588,N_49717);
and UO_1187 (O_1187,N_46767,N_49688);
nand UO_1188 (O_1188,N_49856,N_49317);
nor UO_1189 (O_1189,N_46005,N_46386);
or UO_1190 (O_1190,N_46662,N_45499);
xor UO_1191 (O_1191,N_48476,N_47459);
nor UO_1192 (O_1192,N_47075,N_46213);
xor UO_1193 (O_1193,N_45087,N_45025);
nor UO_1194 (O_1194,N_49404,N_49674);
and UO_1195 (O_1195,N_46693,N_46706);
nand UO_1196 (O_1196,N_49068,N_45497);
nand UO_1197 (O_1197,N_49743,N_46268);
nor UO_1198 (O_1198,N_46685,N_48276);
xor UO_1199 (O_1199,N_49412,N_45452);
or UO_1200 (O_1200,N_47028,N_46747);
nor UO_1201 (O_1201,N_47071,N_47486);
nand UO_1202 (O_1202,N_48313,N_47116);
or UO_1203 (O_1203,N_49207,N_49501);
xnor UO_1204 (O_1204,N_48309,N_45471);
nor UO_1205 (O_1205,N_48889,N_45280);
nor UO_1206 (O_1206,N_49096,N_49021);
nand UO_1207 (O_1207,N_47585,N_46329);
xnor UO_1208 (O_1208,N_49350,N_48088);
nand UO_1209 (O_1209,N_46209,N_45624);
nor UO_1210 (O_1210,N_48970,N_48801);
or UO_1211 (O_1211,N_49305,N_47678);
nor UO_1212 (O_1212,N_45183,N_47097);
nor UO_1213 (O_1213,N_46566,N_47762);
nand UO_1214 (O_1214,N_45501,N_49006);
and UO_1215 (O_1215,N_48815,N_49117);
and UO_1216 (O_1216,N_49857,N_45026);
or UO_1217 (O_1217,N_47909,N_46302);
nor UO_1218 (O_1218,N_47412,N_46614);
and UO_1219 (O_1219,N_47911,N_46370);
or UO_1220 (O_1220,N_48907,N_47580);
nor UO_1221 (O_1221,N_48570,N_46684);
nor UO_1222 (O_1222,N_45852,N_45380);
or UO_1223 (O_1223,N_48234,N_45486);
or UO_1224 (O_1224,N_47257,N_48026);
nand UO_1225 (O_1225,N_48550,N_49492);
nor UO_1226 (O_1226,N_49124,N_48220);
xor UO_1227 (O_1227,N_48186,N_47950);
xnor UO_1228 (O_1228,N_49742,N_45650);
or UO_1229 (O_1229,N_46538,N_48599);
nor UO_1230 (O_1230,N_47232,N_49697);
nor UO_1231 (O_1231,N_48440,N_48464);
nand UO_1232 (O_1232,N_45667,N_48697);
and UO_1233 (O_1233,N_46186,N_48901);
xnor UO_1234 (O_1234,N_45023,N_49768);
xnor UO_1235 (O_1235,N_49429,N_48333);
nor UO_1236 (O_1236,N_49020,N_48947);
and UO_1237 (O_1237,N_47801,N_48717);
and UO_1238 (O_1238,N_49362,N_48013);
and UO_1239 (O_1239,N_48886,N_46015);
nor UO_1240 (O_1240,N_45570,N_47685);
and UO_1241 (O_1241,N_47092,N_49127);
or UO_1242 (O_1242,N_48482,N_48777);
xor UO_1243 (O_1243,N_46624,N_49878);
and UO_1244 (O_1244,N_49718,N_48424);
and UO_1245 (O_1245,N_45635,N_46606);
xnor UO_1246 (O_1246,N_47513,N_49260);
xnor UO_1247 (O_1247,N_49538,N_49472);
xnor UO_1248 (O_1248,N_46180,N_45639);
xnor UO_1249 (O_1249,N_46372,N_49811);
or UO_1250 (O_1250,N_49257,N_48906);
nand UO_1251 (O_1251,N_49673,N_46782);
or UO_1252 (O_1252,N_48942,N_46366);
or UO_1253 (O_1253,N_48277,N_46314);
or UO_1254 (O_1254,N_49487,N_45550);
or UO_1255 (O_1255,N_49037,N_46588);
nand UO_1256 (O_1256,N_45932,N_49267);
or UO_1257 (O_1257,N_49816,N_47841);
or UO_1258 (O_1258,N_46244,N_48048);
and UO_1259 (O_1259,N_45411,N_47007);
nor UO_1260 (O_1260,N_49312,N_46809);
nor UO_1261 (O_1261,N_46261,N_46032);
or UO_1262 (O_1262,N_49475,N_48933);
nor UO_1263 (O_1263,N_45504,N_45576);
or UO_1264 (O_1264,N_49773,N_45801);
or UO_1265 (O_1265,N_49394,N_47637);
xor UO_1266 (O_1266,N_48299,N_46871);
xnor UO_1267 (O_1267,N_49834,N_47368);
and UO_1268 (O_1268,N_45885,N_47220);
nor UO_1269 (O_1269,N_47681,N_46276);
or UO_1270 (O_1270,N_49580,N_47397);
or UO_1271 (O_1271,N_49788,N_45117);
nand UO_1272 (O_1272,N_46770,N_47748);
nand UO_1273 (O_1273,N_45611,N_49450);
nor UO_1274 (O_1274,N_48630,N_46250);
xnor UO_1275 (O_1275,N_48253,N_47864);
nand UO_1276 (O_1276,N_49060,N_46322);
xnor UO_1277 (O_1277,N_46401,N_49739);
nand UO_1278 (O_1278,N_46375,N_46513);
or UO_1279 (O_1279,N_47051,N_48689);
or UO_1280 (O_1280,N_47472,N_45304);
nand UO_1281 (O_1281,N_47021,N_45519);
nor UO_1282 (O_1282,N_47857,N_47552);
nor UO_1283 (O_1283,N_47289,N_45813);
or UO_1284 (O_1284,N_49883,N_48610);
xor UO_1285 (O_1285,N_45103,N_46680);
or UO_1286 (O_1286,N_49982,N_45974);
nand UO_1287 (O_1287,N_47329,N_49173);
xor UO_1288 (O_1288,N_47170,N_48451);
nand UO_1289 (O_1289,N_48543,N_46125);
xnor UO_1290 (O_1290,N_46870,N_49990);
and UO_1291 (O_1291,N_49859,N_48472);
and UO_1292 (O_1292,N_48878,N_48371);
xor UO_1293 (O_1293,N_48354,N_47839);
nand UO_1294 (O_1294,N_47226,N_49896);
and UO_1295 (O_1295,N_45112,N_46596);
nor UO_1296 (O_1296,N_48809,N_46858);
nand UO_1297 (O_1297,N_46741,N_47788);
nand UO_1298 (O_1298,N_45122,N_47677);
or UO_1299 (O_1299,N_48233,N_48887);
or UO_1300 (O_1300,N_47525,N_45451);
or UO_1301 (O_1301,N_47794,N_49814);
or UO_1302 (O_1302,N_49915,N_48227);
or UO_1303 (O_1303,N_49218,N_49331);
nor UO_1304 (O_1304,N_49604,N_47389);
nor UO_1305 (O_1305,N_46802,N_49873);
xnor UO_1306 (O_1306,N_47023,N_45688);
and UO_1307 (O_1307,N_46027,N_46510);
xor UO_1308 (O_1308,N_48965,N_48664);
nor UO_1309 (O_1309,N_46777,N_46589);
nor UO_1310 (O_1310,N_46357,N_48908);
nor UO_1311 (O_1311,N_48514,N_48918);
and UO_1312 (O_1312,N_48991,N_47673);
and UO_1313 (O_1313,N_46294,N_47853);
and UO_1314 (O_1314,N_46922,N_47707);
and UO_1315 (O_1315,N_46496,N_46336);
and UO_1316 (O_1316,N_45594,N_45528);
and UO_1317 (O_1317,N_48640,N_46099);
nand UO_1318 (O_1318,N_45645,N_49131);
or UO_1319 (O_1319,N_48806,N_47024);
nor UO_1320 (O_1320,N_45721,N_46110);
nand UO_1321 (O_1321,N_48760,N_46405);
nand UO_1322 (O_1322,N_47352,N_46641);
nor UO_1323 (O_1323,N_49013,N_48425);
nor UO_1324 (O_1324,N_47743,N_45074);
nor UO_1325 (O_1325,N_45130,N_47514);
xor UO_1326 (O_1326,N_49366,N_49263);
nor UO_1327 (O_1327,N_45458,N_47147);
or UO_1328 (O_1328,N_46108,N_46631);
xor UO_1329 (O_1329,N_48244,N_48494);
xnor UO_1330 (O_1330,N_47430,N_46102);
and UO_1331 (O_1331,N_45680,N_47252);
xnor UO_1332 (O_1332,N_47814,N_45270);
or UO_1333 (O_1333,N_47679,N_45901);
xor UO_1334 (O_1334,N_46560,N_47421);
nand UO_1335 (O_1335,N_45706,N_46061);
xor UO_1336 (O_1336,N_46072,N_47320);
nand UO_1337 (O_1337,N_46986,N_46508);
xor UO_1338 (O_1338,N_48423,N_45970);
nor UO_1339 (O_1339,N_48467,N_45734);
or UO_1340 (O_1340,N_48988,N_45613);
nand UO_1341 (O_1341,N_45599,N_49435);
xnor UO_1342 (O_1342,N_46426,N_46053);
xor UO_1343 (O_1343,N_48006,N_49050);
or UO_1344 (O_1344,N_49581,N_49945);
xor UO_1345 (O_1345,N_49728,N_48493);
nand UO_1346 (O_1346,N_47783,N_45538);
nor UO_1347 (O_1347,N_47963,N_47438);
xor UO_1348 (O_1348,N_49526,N_47579);
xor UO_1349 (O_1349,N_46493,N_49918);
xnor UO_1350 (O_1350,N_48545,N_47310);
or UO_1351 (O_1351,N_48012,N_47031);
nand UO_1352 (O_1352,N_46935,N_46214);
or UO_1353 (O_1353,N_49499,N_48063);
nand UO_1354 (O_1354,N_45768,N_49800);
and UO_1355 (O_1355,N_45473,N_49187);
xor UO_1356 (O_1356,N_48926,N_45623);
and UO_1357 (O_1357,N_47434,N_48120);
xor UO_1358 (O_1358,N_48624,N_48182);
nor UO_1359 (O_1359,N_49201,N_49077);
xor UO_1360 (O_1360,N_48765,N_48999);
xor UO_1361 (O_1361,N_48891,N_46909);
nor UO_1362 (O_1362,N_47516,N_47001);
or UO_1363 (O_1363,N_48856,N_46896);
xor UO_1364 (O_1364,N_49916,N_48769);
and UO_1365 (O_1365,N_45929,N_47495);
nor UO_1366 (O_1366,N_45774,N_46188);
xor UO_1367 (O_1367,N_45869,N_47976);
and UO_1368 (O_1368,N_47510,N_47942);
nor UO_1369 (O_1369,N_45729,N_47676);
xnor UO_1370 (O_1370,N_45571,N_49649);
and UO_1371 (O_1371,N_47832,N_46642);
and UO_1372 (O_1372,N_49110,N_49262);
or UO_1373 (O_1373,N_47172,N_48585);
xor UO_1374 (O_1374,N_45196,N_47463);
and UO_1375 (O_1375,N_45385,N_45242);
nor UO_1376 (O_1376,N_46743,N_47692);
xor UO_1377 (O_1377,N_45707,N_49926);
nand UO_1378 (O_1378,N_46764,N_49957);
or UO_1379 (O_1379,N_46788,N_45349);
nand UO_1380 (O_1380,N_46486,N_48800);
nand UO_1381 (O_1381,N_49365,N_48710);
xor UO_1382 (O_1382,N_46879,N_45503);
and UO_1383 (O_1383,N_48017,N_45592);
and UO_1384 (O_1384,N_46618,N_47319);
and UO_1385 (O_1385,N_48393,N_47761);
xnor UO_1386 (O_1386,N_45641,N_48384);
or UO_1387 (O_1387,N_45251,N_49951);
xnor UO_1388 (O_1388,N_46908,N_46062);
xor UO_1389 (O_1389,N_47118,N_46227);
xnor UO_1390 (O_1390,N_46198,N_45344);
and UO_1391 (O_1391,N_49149,N_47159);
or UO_1392 (O_1392,N_49420,N_45296);
xor UO_1393 (O_1393,N_47863,N_47756);
nor UO_1394 (O_1394,N_45821,N_46888);
and UO_1395 (O_1395,N_48759,N_46930);
xor UO_1396 (O_1396,N_47724,N_49411);
nor UO_1397 (O_1397,N_49103,N_49973);
nand UO_1398 (O_1398,N_45811,N_48915);
nand UO_1399 (O_1399,N_47654,N_45193);
xor UO_1400 (O_1400,N_49359,N_45727);
nor UO_1401 (O_1401,N_48137,N_46088);
or UO_1402 (O_1402,N_46813,N_45352);
or UO_1403 (O_1403,N_49635,N_45919);
and UO_1404 (O_1404,N_49469,N_47033);
nand UO_1405 (O_1405,N_45409,N_48014);
xor UO_1406 (O_1406,N_46090,N_46494);
nor UO_1407 (O_1407,N_49430,N_45840);
nand UO_1408 (O_1408,N_45088,N_45494);
xnor UO_1409 (O_1409,N_46290,N_45479);
nor UO_1410 (O_1410,N_46657,N_49324);
or UO_1411 (O_1411,N_45798,N_47844);
nand UO_1412 (O_1412,N_46028,N_45024);
xnor UO_1413 (O_1413,N_49076,N_47016);
or UO_1414 (O_1414,N_48128,N_48239);
or UO_1415 (O_1415,N_45125,N_48398);
nor UO_1416 (O_1416,N_45098,N_45312);
nor UO_1417 (O_1417,N_46128,N_47193);
or UO_1418 (O_1418,N_45985,N_47894);
nor UO_1419 (O_1419,N_48155,N_47733);
nand UO_1420 (O_1420,N_45297,N_49523);
and UO_1421 (O_1421,N_47918,N_48804);
nand UO_1422 (O_1422,N_48442,N_49530);
and UO_1423 (O_1423,N_45414,N_45730);
and UO_1424 (O_1424,N_45436,N_47626);
xnor UO_1425 (O_1425,N_47501,N_45946);
nand UO_1426 (O_1426,N_48298,N_48178);
and UO_1427 (O_1427,N_48488,N_45759);
nor UO_1428 (O_1428,N_45690,N_49502);
nor UO_1429 (O_1429,N_46966,N_46711);
or UO_1430 (O_1430,N_49989,N_47291);
or UO_1431 (O_1431,N_45269,N_48050);
or UO_1432 (O_1432,N_47249,N_48212);
and UO_1433 (O_1433,N_45056,N_46959);
nand UO_1434 (O_1434,N_46374,N_49967);
nand UO_1435 (O_1435,N_45711,N_47393);
nand UO_1436 (O_1436,N_49048,N_46315);
or UO_1437 (O_1437,N_46892,N_48890);
or UO_1438 (O_1438,N_47173,N_47130);
or UO_1439 (O_1439,N_49158,N_48015);
nand UO_1440 (O_1440,N_46237,N_48979);
nor UO_1441 (O_1441,N_48871,N_45553);
and UO_1442 (O_1442,N_47968,N_49278);
xor UO_1443 (O_1443,N_46158,N_45443);
or UO_1444 (O_1444,N_46225,N_48897);
nor UO_1445 (O_1445,N_48575,N_46562);
nor UO_1446 (O_1446,N_49334,N_49043);
nor UO_1447 (O_1447,N_48432,N_47194);
and UO_1448 (O_1448,N_48466,N_46452);
and UO_1449 (O_1449,N_46021,N_49657);
xor UO_1450 (O_1450,N_46840,N_47072);
xor UO_1451 (O_1451,N_47481,N_49386);
and UO_1452 (O_1452,N_49870,N_47396);
nor UO_1453 (O_1453,N_46865,N_46837);
nand UO_1454 (O_1454,N_45007,N_45682);
xnor UO_1455 (O_1455,N_49825,N_49441);
xnor UO_1456 (O_1456,N_46258,N_45427);
nor UO_1457 (O_1457,N_48261,N_46627);
xor UO_1458 (O_1458,N_49537,N_47185);
or UO_1459 (O_1459,N_46057,N_45708);
nor UO_1460 (O_1460,N_46167,N_49471);
or UO_1461 (O_1461,N_49626,N_48058);
nor UO_1462 (O_1462,N_46827,N_47059);
nor UO_1463 (O_1463,N_45722,N_46154);
nand UO_1464 (O_1464,N_47180,N_48787);
or UO_1465 (O_1465,N_47713,N_49108);
and UO_1466 (O_1466,N_48733,N_48696);
nand UO_1467 (O_1467,N_47861,N_47827);
xor UO_1468 (O_1468,N_48111,N_46994);
nor UO_1469 (O_1469,N_47821,N_47810);
and UO_1470 (O_1470,N_48474,N_47365);
or UO_1471 (O_1471,N_48583,N_45255);
nor UO_1472 (O_1472,N_49364,N_45446);
or UO_1473 (O_1473,N_49141,N_48338);
xnor UO_1474 (O_1474,N_47899,N_46965);
nand UO_1475 (O_1475,N_45236,N_45365);
or UO_1476 (O_1476,N_46071,N_45698);
and UO_1477 (O_1477,N_46739,N_47754);
xnor UO_1478 (O_1478,N_47000,N_47898);
and UO_1479 (O_1479,N_46818,N_45787);
nor UO_1480 (O_1480,N_46466,N_45648);
and UO_1481 (O_1481,N_49303,N_45891);
xnor UO_1482 (O_1482,N_48308,N_46567);
or UO_1483 (O_1483,N_46440,N_47030);
and UO_1484 (O_1484,N_47217,N_49837);
and UO_1485 (O_1485,N_46656,N_45256);
nor UO_1486 (O_1486,N_47178,N_49323);
nand UO_1487 (O_1487,N_45902,N_49326);
and UO_1488 (O_1488,N_48729,N_47035);
xnor UO_1489 (O_1489,N_49630,N_49381);
nand UO_1490 (O_1490,N_48512,N_49737);
or UO_1491 (O_1491,N_49348,N_49772);
xor UO_1492 (O_1492,N_46054,N_49609);
or UO_1493 (O_1493,N_49291,N_49142);
nor UO_1494 (O_1494,N_45253,N_45998);
nand UO_1495 (O_1495,N_45647,N_47467);
nor UO_1496 (O_1496,N_49573,N_46035);
and UO_1497 (O_1497,N_47284,N_48894);
nor UO_1498 (O_1498,N_45733,N_49832);
nor UO_1499 (O_1499,N_49651,N_45034);
nor UO_1500 (O_1500,N_46480,N_45585);
and UO_1501 (O_1501,N_48235,N_48225);
and UO_1502 (O_1502,N_47448,N_46726);
or UO_1503 (O_1503,N_46491,N_46660);
nor UO_1504 (O_1504,N_46880,N_49156);
nor UO_1505 (O_1505,N_48051,N_45164);
nor UO_1506 (O_1506,N_47954,N_45860);
nor UO_1507 (O_1507,N_49678,N_49763);
and UO_1508 (O_1508,N_46530,N_48143);
and UO_1509 (O_1509,N_49661,N_47455);
xnor UO_1510 (O_1510,N_45113,N_48179);
and UO_1511 (O_1511,N_46288,N_45765);
nand UO_1512 (O_1512,N_47529,N_46267);
or UO_1513 (O_1513,N_46179,N_49042);
nor UO_1514 (O_1514,N_47039,N_46458);
nor UO_1515 (O_1515,N_47594,N_48507);
nor UO_1516 (O_1516,N_49564,N_48857);
xor UO_1517 (O_1517,N_46055,N_45695);
or UO_1518 (O_1518,N_47162,N_45204);
xnor UO_1519 (O_1519,N_45857,N_49470);
or UO_1520 (O_1520,N_45354,N_49533);
nand UO_1521 (O_1521,N_45058,N_46783);
or UO_1522 (O_1522,N_47859,N_45562);
nand UO_1523 (O_1523,N_48613,N_45376);
nand UO_1524 (O_1524,N_48779,N_48684);
xnor UO_1525 (O_1525,N_47414,N_45186);
or UO_1526 (O_1526,N_46318,N_49868);
xnor UO_1527 (O_1527,N_47889,N_49400);
nor UO_1528 (O_1528,N_48484,N_49357);
or UO_1529 (O_1529,N_49456,N_48158);
xnor UO_1530 (O_1530,N_45396,N_45126);
nor UO_1531 (O_1531,N_46583,N_49841);
and UO_1532 (O_1532,N_47219,N_45416);
and UO_1533 (O_1533,N_45205,N_47491);
and UO_1534 (O_1534,N_47561,N_45793);
nor UO_1535 (O_1535,N_47882,N_47710);
nor UO_1536 (O_1536,N_49015,N_49548);
and UO_1537 (O_1537,N_46955,N_48537);
and UO_1538 (O_1538,N_47633,N_49295);
nand UO_1539 (O_1539,N_49179,N_49306);
or UO_1540 (O_1540,N_45792,N_49284);
or UO_1541 (O_1541,N_48858,N_45163);
nor UO_1542 (O_1542,N_48105,N_45947);
xor UO_1543 (O_1543,N_48631,N_49919);
nand UO_1544 (O_1544,N_47602,N_45996);
xnor UO_1545 (O_1545,N_48922,N_46869);
xor UO_1546 (O_1546,N_46400,N_49509);
nand UO_1547 (O_1547,N_49504,N_46898);
nor UO_1548 (O_1548,N_49041,N_45806);
xnor UO_1549 (O_1549,N_45786,N_45120);
and UO_1550 (O_1550,N_48173,N_49304);
and UO_1551 (O_1551,N_49652,N_46080);
nand UO_1552 (O_1552,N_45295,N_47038);
xnor UO_1553 (O_1553,N_46576,N_48521);
nand UO_1554 (O_1554,N_49797,N_49237);
nor UO_1555 (O_1555,N_45350,N_45760);
xor UO_1556 (O_1556,N_45791,N_46926);
nand UO_1557 (O_1557,N_48405,N_48406);
or UO_1558 (O_1558,N_48363,N_47378);
or UO_1559 (O_1559,N_48984,N_47315);
nor UO_1560 (O_1560,N_49195,N_47696);
nand UO_1561 (O_1561,N_49924,N_47124);
or UO_1562 (O_1562,N_48571,N_48231);
nor UO_1563 (O_1563,N_48892,N_45450);
nor UO_1564 (O_1564,N_45566,N_49824);
xnor UO_1565 (O_1565,N_48685,N_46535);
xor UO_1566 (O_1566,N_48290,N_46563);
or UO_1567 (O_1567,N_45883,N_46515);
and UO_1568 (O_1568,N_48711,N_49421);
nand UO_1569 (O_1569,N_46085,N_48124);
xnor UO_1570 (O_1570,N_46252,N_48074);
nand UO_1571 (O_1571,N_49908,N_49513);
or UO_1572 (O_1572,N_49946,N_45138);
nor UO_1573 (O_1573,N_49172,N_46044);
nor UO_1574 (O_1574,N_45146,N_48396);
xnor UO_1575 (O_1575,N_49597,N_48262);
and UO_1576 (O_1576,N_47568,N_45913);
and UO_1577 (O_1577,N_48091,N_48913);
xnor UO_1578 (O_1578,N_46042,N_46873);
nand UO_1579 (O_1579,N_48686,N_49061);
xor UO_1580 (O_1580,N_46833,N_45955);
and UO_1581 (O_1581,N_45022,N_48826);
xnor UO_1582 (O_1582,N_46279,N_45329);
or UO_1583 (O_1583,N_45693,N_47607);
xnor UO_1584 (O_1584,N_46533,N_49632);
and UO_1585 (O_1585,N_49750,N_45371);
and UO_1586 (O_1586,N_48985,N_47002);
xnor UO_1587 (O_1587,N_47050,N_46866);
nand UO_1588 (O_1588,N_45895,N_49204);
and UO_1589 (O_1589,N_49984,N_49941);
nor UO_1590 (O_1590,N_47238,N_49793);
xnor UO_1591 (O_1591,N_47948,N_46953);
nand UO_1592 (O_1592,N_45724,N_45228);
or UO_1593 (O_1593,N_49521,N_46805);
xor UO_1594 (O_1594,N_45723,N_45782);
nand UO_1595 (O_1595,N_46503,N_47905);
nor UO_1596 (O_1596,N_48382,N_48078);
nand UO_1597 (O_1597,N_47499,N_47047);
nand UO_1598 (O_1598,N_49642,N_49054);
and UO_1599 (O_1599,N_45468,N_45616);
nor UO_1600 (O_1600,N_47061,N_48001);
xnor UO_1601 (O_1601,N_46193,N_45214);
nand UO_1602 (O_1602,N_45415,N_45402);
and UO_1603 (O_1603,N_47168,N_49132);
nand UO_1604 (O_1604,N_47349,N_45775);
xnor UO_1605 (O_1605,N_46763,N_45173);
or UO_1606 (O_1606,N_46746,N_45336);
nor UO_1607 (O_1607,N_46271,N_47216);
nand UO_1608 (O_1608,N_47235,N_48766);
xnor UO_1609 (O_1609,N_46829,N_47559);
nor UO_1610 (O_1610,N_48468,N_48885);
nand UO_1611 (O_1611,N_46419,N_48665);
xnor UO_1612 (O_1612,N_49259,N_47730);
nor UO_1613 (O_1613,N_45288,N_45094);
nand UO_1614 (O_1614,N_47348,N_45638);
nor UO_1615 (O_1615,N_48495,N_49084);
nor UO_1616 (O_1616,N_45169,N_45390);
xor UO_1617 (O_1617,N_49315,N_48812);
nand UO_1618 (O_1618,N_47769,N_45063);
nand UO_1619 (O_1619,N_46429,N_48421);
or UO_1620 (O_1620,N_48692,N_48546);
nor UO_1621 (O_1621,N_47838,N_47797);
or UO_1622 (O_1622,N_49848,N_46221);
or UO_1623 (O_1623,N_45944,N_49723);
or UO_1624 (O_1624,N_46153,N_45460);
xor UO_1625 (O_1625,N_45492,N_48811);
nor UO_1626 (O_1626,N_48981,N_46708);
xnor UO_1627 (O_1627,N_48089,N_47182);
or UO_1628 (O_1628,N_47371,N_46454);
or UO_1629 (O_1629,N_46143,N_47046);
xnor UO_1630 (O_1630,N_48416,N_48989);
and UO_1631 (O_1631,N_45552,N_46427);
and UO_1632 (O_1632,N_45028,N_49164);
or UO_1633 (O_1633,N_48796,N_45219);
xnor UO_1634 (O_1634,N_48694,N_47406);
nor UO_1635 (O_1635,N_49432,N_47452);
nor UO_1636 (O_1636,N_45663,N_46913);
and UO_1637 (O_1637,N_49423,N_47786);
xor UO_1638 (O_1638,N_45107,N_45830);
nor UO_1639 (O_1639,N_47904,N_45047);
xor UO_1640 (O_1640,N_46256,N_46591);
nor UO_1641 (O_1641,N_47981,N_45188);
nand UO_1642 (O_1642,N_48930,N_47961);
and UO_1643 (O_1643,N_46715,N_45601);
xor UO_1644 (O_1644,N_45950,N_49126);
nor UO_1645 (O_1645,N_49640,N_46414);
nand UO_1646 (O_1646,N_48500,N_45716);
xnor UO_1647 (O_1647,N_48750,N_48839);
xnor UO_1648 (O_1648,N_49715,N_49415);
and UO_1649 (O_1649,N_45968,N_46139);
nand UO_1650 (O_1650,N_46505,N_45334);
nand UO_1651 (O_1651,N_47504,N_45271);
nor UO_1652 (O_1652,N_47141,N_46049);
and UO_1653 (O_1653,N_48625,N_47342);
xor UO_1654 (O_1654,N_48797,N_48265);
nor UO_1655 (O_1655,N_49925,N_49627);
nand UO_1656 (O_1656,N_48616,N_47603);
and UO_1657 (O_1657,N_48538,N_47920);
nor UO_1658 (O_1658,N_49032,N_48118);
nand UO_1659 (O_1659,N_49095,N_48201);
xnor UO_1660 (O_1660,N_47806,N_45495);
nand UO_1661 (O_1661,N_48200,N_46477);
and UO_1662 (O_1662,N_48248,N_46864);
or UO_1663 (O_1663,N_47778,N_45684);
and UO_1664 (O_1664,N_45168,N_49029);
xor UO_1665 (O_1665,N_49569,N_47653);
nand UO_1666 (O_1666,N_48556,N_49392);
nand UO_1667 (O_1667,N_47224,N_47022);
or UO_1668 (O_1668,N_45976,N_45254);
and UO_1669 (O_1669,N_46145,N_49328);
and UO_1670 (O_1670,N_48718,N_46632);
nor UO_1671 (O_1671,N_47277,N_47308);
or UO_1672 (O_1672,N_49804,N_48648);
or UO_1673 (O_1673,N_49205,N_48140);
xor UO_1674 (O_1674,N_46611,N_47017);
nand UO_1675 (O_1675,N_49446,N_48457);
xnor UO_1676 (O_1676,N_48291,N_45580);
nor UO_1677 (O_1677,N_45172,N_48281);
and UO_1678 (O_1678,N_49388,N_45535);
and UO_1679 (O_1679,N_45990,N_47818);
nor UO_1680 (O_1680,N_49623,N_46359);
nor UO_1681 (O_1681,N_49067,N_47020);
and UO_1682 (O_1682,N_45448,N_46444);
and UO_1683 (O_1683,N_47648,N_46761);
nand UO_1684 (O_1684,N_48843,N_47198);
xor UO_1685 (O_1685,N_48972,N_46333);
xor UO_1686 (O_1686,N_45581,N_47358);
nor UO_1687 (O_1687,N_48028,N_45989);
and UO_1688 (O_1688,N_48283,N_49625);
xor UO_1689 (O_1689,N_49826,N_47392);
or UO_1690 (O_1690,N_46674,N_46334);
nor UO_1691 (O_1691,N_48560,N_45563);
xor UO_1692 (O_1692,N_46070,N_49167);
xnor UO_1693 (O_1693,N_47630,N_47015);
xnor UO_1694 (O_1694,N_45187,N_47509);
xor UO_1695 (O_1695,N_46134,N_45761);
and UO_1696 (O_1696,N_49901,N_47741);
xor UO_1697 (O_1697,N_45703,N_45332);
nor UO_1698 (O_1698,N_46342,N_47036);
or UO_1699 (O_1699,N_47601,N_48751);
nor UO_1700 (O_1700,N_47914,N_47161);
or UO_1701 (O_1701,N_49757,N_48461);
nor UO_1702 (O_1702,N_47009,N_48872);
nor UO_1703 (O_1703,N_45286,N_46991);
and UO_1704 (O_1704,N_48505,N_48040);
nand UO_1705 (O_1705,N_45232,N_47554);
nor UO_1706 (O_1706,N_48167,N_46281);
or UO_1707 (O_1707,N_45892,N_45900);
and UO_1708 (O_1708,N_48502,N_46595);
and UO_1709 (O_1709,N_49731,N_49514);
nand UO_1710 (O_1710,N_48419,N_47694);
xor UO_1711 (O_1711,N_45434,N_48549);
nor UO_1712 (O_1712,N_45200,N_46824);
and UO_1713 (O_1713,N_49072,N_47343);
nor UO_1714 (O_1714,N_47804,N_46306);
nand UO_1715 (O_1715,N_46197,N_47375);
nor UO_1716 (O_1716,N_47146,N_46794);
and UO_1717 (O_1717,N_48654,N_49045);
and UO_1718 (O_1718,N_45262,N_46045);
or UO_1719 (O_1719,N_47773,N_49414);
and UO_1720 (O_1720,N_46878,N_47787);
nand UO_1721 (O_1721,N_47518,N_46262);
nor UO_1722 (O_1722,N_47745,N_45575);
and UO_1723 (O_1723,N_49751,N_47970);
nor UO_1724 (O_1724,N_47294,N_48255);
or UO_1725 (O_1725,N_46481,N_45629);
xor UO_1726 (O_1726,N_48145,N_49961);
or UO_1727 (O_1727,N_49376,N_47991);
nand UO_1728 (O_1728,N_46506,N_49734);
nor UO_1729 (O_1729,N_49889,N_48289);
nand UO_1730 (O_1730,N_49210,N_49436);
xnor UO_1731 (O_1731,N_46556,N_46187);
and UO_1732 (O_1732,N_48181,N_47951);
xnor UO_1733 (O_1733,N_47334,N_48551);
xnor UO_1734 (O_1734,N_48321,N_47711);
and UO_1735 (O_1735,N_45884,N_47086);
or UO_1736 (O_1736,N_46298,N_48197);
and UO_1737 (O_1737,N_49261,N_48358);
xnor UO_1738 (O_1738,N_46181,N_47634);
xor UO_1739 (O_1739,N_47796,N_45082);
and UO_1740 (O_1740,N_46335,N_46982);
nor UO_1741 (O_1741,N_46929,N_49296);
and UO_1742 (O_1742,N_46220,N_49026);
and UO_1743 (O_1743,N_46131,N_47132);
nand UO_1744 (O_1744,N_48632,N_47202);
nand UO_1745 (O_1745,N_46148,N_48709);
nand UO_1746 (O_1746,N_47206,N_47435);
or UO_1747 (O_1747,N_46343,N_49911);
xor UO_1748 (O_1748,N_45044,N_48133);
and UO_1749 (O_1749,N_48780,N_47674);
nor UO_1750 (O_1750,N_48097,N_45403);
nor UO_1751 (O_1751,N_46004,N_48578);
and UO_1752 (O_1752,N_47631,N_49897);
xnor UO_1753 (O_1753,N_48566,N_49000);
and UO_1754 (O_1754,N_49405,N_46621);
nand UO_1755 (O_1755,N_49928,N_46686);
nor UO_1756 (O_1756,N_46378,N_45861);
nor UO_1757 (O_1757,N_48036,N_45819);
nand UO_1758 (O_1758,N_45980,N_49252);
and UO_1759 (O_1759,N_45870,N_49055);
nand UO_1760 (O_1760,N_46361,N_45447);
and UO_1761 (O_1761,N_47461,N_45337);
xor UO_1762 (O_1762,N_49266,N_45463);
or UO_1763 (O_1763,N_45301,N_49740);
nor UO_1764 (O_1764,N_49881,N_47093);
or UO_1765 (O_1765,N_49707,N_45147);
xor UO_1766 (O_1766,N_47691,N_45227);
xor UO_1767 (O_1767,N_47078,N_48252);
nand UO_1768 (O_1768,N_47437,N_46630);
xnor UO_1769 (O_1769,N_45002,N_49216);
and UO_1770 (O_1770,N_47500,N_46465);
xor UO_1771 (O_1771,N_47306,N_48832);
nand UO_1772 (O_1772,N_45812,N_47699);
and UO_1773 (O_1773,N_48827,N_49092);
xnor UO_1774 (O_1774,N_46665,N_48534);
nand UO_1775 (O_1775,N_49406,N_46083);
xnor UO_1776 (O_1776,N_45595,N_47382);
or UO_1777 (O_1777,N_49354,N_49940);
nand UO_1778 (O_1778,N_47856,N_49234);
and UO_1779 (O_1779,N_45238,N_47473);
nand UO_1780 (O_1780,N_45248,N_48374);
or UO_1781 (O_1781,N_48129,N_47750);
or UO_1782 (O_1782,N_46449,N_46094);
nand UO_1783 (O_1783,N_45573,N_46604);
nand UO_1784 (O_1784,N_47260,N_45672);
nor UO_1785 (O_1785,N_48106,N_45480);
nor UO_1786 (O_1786,N_48098,N_48443);
nand UO_1787 (O_1787,N_45728,N_48963);
xnor UO_1788 (O_1788,N_46709,N_45093);
nand UO_1789 (O_1789,N_49559,N_48414);
nor UO_1790 (O_1790,N_47062,N_45096);
nor UO_1791 (O_1791,N_48966,N_48413);
or UO_1792 (O_1792,N_46455,N_48928);
and UO_1793 (O_1793,N_45155,N_49484);
nor UO_1794 (O_1794,N_45874,N_45092);
nor UO_1795 (O_1795,N_47210,N_46807);
or UO_1796 (O_1796,N_45689,N_48716);
or UO_1797 (O_1797,N_47746,N_46816);
or UO_1798 (O_1798,N_48314,N_46270);
xor UO_1799 (O_1799,N_46459,N_48977);
nand UO_1800 (O_1800,N_47627,N_47163);
xor UO_1801 (O_1801,N_45381,N_46418);
and UO_1802 (O_1802,N_48112,N_47998);
or UO_1803 (O_1803,N_47417,N_48072);
or UO_1804 (O_1804,N_46104,N_48065);
nor UO_1805 (O_1805,N_48968,N_48294);
nor UO_1806 (O_1806,N_45590,N_48162);
xor UO_1807 (O_1807,N_47933,N_48207);
nor UO_1808 (O_1808,N_49496,N_47791);
nor UO_1809 (O_1809,N_48019,N_45265);
nand UO_1810 (O_1810,N_46598,N_49650);
and UO_1811 (O_1811,N_49777,N_45300);
nand UO_1812 (O_1812,N_45977,N_46902);
xnor UO_1813 (O_1813,N_45567,N_49765);
xor UO_1814 (O_1814,N_48869,N_48356);
nand UO_1815 (O_1815,N_49114,N_48978);
xor UO_1816 (O_1816,N_49227,N_48535);
nand UO_1817 (O_1817,N_49198,N_47042);
and UO_1818 (O_1818,N_48845,N_45614);
nor UO_1819 (O_1819,N_46948,N_46717);
xor UO_1820 (O_1820,N_48463,N_45785);
nor UO_1821 (O_1821,N_47316,N_45880);
or UO_1822 (O_1822,N_45507,N_47364);
nand UO_1823 (O_1823,N_45177,N_46907);
and UO_1824 (O_1824,N_48326,N_47828);
xor UO_1825 (O_1825,N_49316,N_48614);
and UO_1826 (O_1826,N_48232,N_47996);
or UO_1827 (O_1827,N_48202,N_46856);
or UO_1828 (O_1828,N_46341,N_47489);
nor UO_1829 (O_1829,N_47824,N_46687);
nor UO_1830 (O_1830,N_46944,N_46707);
nand UO_1831 (O_1831,N_49758,N_47314);
or UO_1832 (O_1832,N_48903,N_48388);
nand UO_1833 (O_1833,N_49866,N_49500);
xnor UO_1834 (O_1834,N_47400,N_47405);
nor UO_1835 (O_1835,N_47158,N_45926);
nor UO_1836 (O_1836,N_48010,N_45404);
xor UO_1837 (O_1837,N_49099,N_45742);
or UO_1838 (O_1838,N_48949,N_49598);
and UO_1839 (O_1839,N_47809,N_47612);
xnor UO_1840 (O_1840,N_47253,N_45982);
or UO_1841 (O_1841,N_47903,N_49243);
and UO_1842 (O_1842,N_48533,N_46164);
or UO_1843 (O_1843,N_48555,N_46327);
and UO_1844 (O_1844,N_47374,N_47702);
nand UO_1845 (O_1845,N_47218,N_45178);
nand UO_1846 (O_1846,N_49356,N_46718);
xnor UO_1847 (O_1847,N_46228,N_45064);
xor UO_1848 (O_1848,N_47969,N_47923);
nor UO_1849 (O_1849,N_48056,N_48189);
xnor UO_1850 (O_1850,N_47207,N_45090);
and UO_1851 (O_1851,N_49547,N_45637);
and UO_1852 (O_1852,N_47567,N_45790);
and UO_1853 (O_1853,N_45568,N_47658);
nand UO_1854 (O_1854,N_45654,N_47704);
nand UO_1855 (O_1855,N_46894,N_45151);
or UO_1856 (O_1856,N_47738,N_45578);
and UO_1857 (O_1857,N_45921,N_45466);
nor UO_1858 (O_1858,N_45424,N_48373);
nor UO_1859 (O_1859,N_48204,N_48902);
and UO_1860 (O_1860,N_49422,N_49683);
or UO_1861 (O_1861,N_49093,N_46058);
nor UO_1862 (O_1862,N_49230,N_48659);
xnor UO_1863 (O_1863,N_47695,N_47094);
nand UO_1864 (O_1864,N_48318,N_48156);
nor UO_1865 (O_1865,N_45425,N_48317);
nor UO_1866 (O_1866,N_49621,N_47243);
nor UO_1867 (O_1867,N_48714,N_48324);
nand UO_1868 (O_1868,N_47624,N_45842);
nor UO_1869 (O_1869,N_48188,N_47706);
xor UO_1870 (O_1870,N_47650,N_45714);
nand UO_1871 (O_1871,N_45420,N_47323);
or UO_1872 (O_1872,N_46303,N_49221);
nor UO_1873 (O_1873,N_47436,N_46138);
nand UO_1874 (O_1874,N_47833,N_48221);
nor UO_1875 (O_1875,N_46691,N_48386);
nor UO_1876 (O_1876,N_49489,N_46282);
nand UO_1877 (O_1877,N_48039,N_48263);
xor UO_1878 (O_1878,N_46625,N_47439);
xor UO_1879 (O_1879,N_46140,N_49010);
and UO_1880 (O_1880,N_46738,N_49165);
nor UO_1881 (O_1881,N_47157,N_48676);
xnor UO_1882 (O_1882,N_46753,N_48835);
xnor UO_1883 (O_1883,N_46030,N_46939);
nand UO_1884 (O_1884,N_48732,N_48246);
nor UO_1885 (O_1885,N_48081,N_48082);
and UO_1886 (O_1886,N_47419,N_45617);
nor UO_1887 (O_1887,N_48284,N_48935);
or UO_1888 (O_1888,N_49007,N_45928);
xnor UO_1889 (O_1889,N_49416,N_49684);
or UO_1890 (O_1890,N_49022,N_49558);
nor UO_1891 (O_1891,N_48024,N_46344);
nand UO_1892 (O_1892,N_46985,N_48912);
and UO_1893 (O_1893,N_49169,N_46723);
and UO_1894 (O_1894,N_45053,N_47799);
nor UO_1895 (O_1895,N_47195,N_45324);
nand UO_1896 (O_1896,N_47293,N_47484);
xnor UO_1897 (O_1897,N_47764,N_45072);
xnor UO_1898 (O_1898,N_45561,N_47871);
or UO_1899 (O_1899,N_46774,N_46280);
and UO_1900 (O_1900,N_48971,N_45737);
or UO_1901 (O_1901,N_49293,N_47790);
and UO_1902 (O_1902,N_45948,N_49839);
and UO_1903 (O_1903,N_47099,N_49431);
nand UO_1904 (O_1904,N_45952,N_47524);
xor UO_1905 (O_1905,N_46464,N_48825);
and UO_1906 (O_1906,N_46565,N_45967);
nand UO_1907 (O_1907,N_45331,N_49321);
nor UO_1908 (O_1908,N_47869,N_49979);
or UO_1909 (O_1909,N_49934,N_45100);
xor UO_1910 (O_1910,N_48539,N_47858);
or UO_1911 (O_1911,N_47995,N_49787);
or UO_1912 (O_1912,N_45917,N_45367);
or UO_1913 (O_1913,N_48208,N_46804);
or UO_1914 (O_1914,N_48705,N_45997);
nand UO_1915 (O_1915,N_48643,N_46580);
or UO_1916 (O_1916,N_49754,N_45878);
xor UO_1917 (O_1917,N_48609,N_48250);
nand UO_1918 (O_1918,N_48943,N_45619);
and UO_1919 (O_1919,N_48916,N_45810);
and UO_1920 (O_1920,N_49225,N_49066);
xnor UO_1921 (O_1921,N_48027,N_45257);
and UO_1922 (O_1922,N_46917,N_46847);
or UO_1923 (O_1923,N_49506,N_49333);
nand UO_1924 (O_1924,N_48311,N_45137);
nand UO_1925 (O_1925,N_46497,N_46528);
and UO_1926 (O_1926,N_47845,N_48653);
nor UO_1927 (O_1927,N_46233,N_45923);
nor UO_1928 (O_1928,N_48343,N_46013);
nand UO_1929 (O_1929,N_49987,N_48764);
nor UO_1930 (O_1930,N_45565,N_46780);
xor UO_1931 (O_1931,N_45014,N_48061);
or UO_1932 (O_1932,N_45259,N_45653);
and UO_1933 (O_1933,N_46964,N_48719);
nand UO_1934 (O_1934,N_46597,N_46605);
and UO_1935 (O_1935,N_47805,N_48340);
nor UO_1936 (O_1936,N_46502,N_45027);
and UO_1937 (O_1937,N_45541,N_49235);
or UO_1938 (O_1938,N_49877,N_48403);
nor UO_1939 (O_1939,N_47785,N_47535);
and UO_1940 (O_1940,N_47174,N_46672);
nand UO_1941 (O_1941,N_48117,N_46251);
xor UO_1942 (O_1942,N_48366,N_47290);
and UO_1943 (O_1943,N_45029,N_48909);
or UO_1944 (O_1944,N_46933,N_49049);
xnor UO_1945 (O_1945,N_46696,N_46137);
nand UO_1946 (O_1946,N_45940,N_45784);
or UO_1947 (O_1947,N_49965,N_49409);
or UO_1948 (O_1948,N_47614,N_47772);
nor UO_1949 (O_1949,N_47508,N_49849);
or UO_1950 (O_1950,N_48258,N_49053);
nand UO_1951 (O_1951,N_49937,N_45839);
or UO_1952 (O_1952,N_46478,N_48192);
xor UO_1953 (O_1953,N_48236,N_49393);
or UO_1954 (O_1954,N_49298,N_49183);
nor UO_1955 (O_1955,N_46484,N_49398);
nand UO_1956 (O_1956,N_45316,N_46831);
or UO_1957 (O_1957,N_49440,N_47879);
or UO_1958 (O_1958,N_47717,N_46504);
xor UO_1959 (O_1959,N_49036,N_46744);
xor UO_1960 (O_1960,N_46119,N_46558);
xnor UO_1961 (O_1961,N_46300,N_46230);
xor UO_1962 (O_1962,N_46077,N_45520);
or UO_1963 (O_1963,N_47264,N_46412);
nor UO_1964 (O_1964,N_49297,N_48103);
xnor UO_1965 (O_1965,N_45622,N_46901);
nand UO_1966 (O_1966,N_45735,N_48847);
and UO_1967 (O_1967,N_45037,N_48612);
xnor UO_1968 (O_1968,N_45736,N_49461);
xor UO_1969 (O_1969,N_45945,N_48404);
and UO_1970 (O_1970,N_48153,N_46799);
and UO_1971 (O_1971,N_45483,N_49301);
nand UO_1972 (O_1972,N_49855,N_48623);
xnor UO_1973 (O_1973,N_45119,N_48247);
xnor UO_1974 (O_1974,N_46165,N_46963);
nor UO_1975 (O_1975,N_48629,N_47929);
nor UO_1976 (O_1976,N_49080,N_49795);
xor UO_1977 (O_1977,N_48031,N_45041);
xnor UO_1978 (O_1978,N_46095,N_47548);
or UO_1979 (O_1979,N_46555,N_47395);
nand UO_1980 (O_1980,N_45067,N_45631);
xnor UO_1981 (O_1981,N_46301,N_47530);
nand UO_1982 (O_1982,N_45144,N_46304);
nand UO_1983 (O_1983,N_48884,N_47947);
xor UO_1984 (O_1984,N_48982,N_47737);
nor UO_1985 (O_1985,N_47222,N_49138);
nand UO_1986 (O_1986,N_49637,N_46191);
and UO_1987 (O_1987,N_47591,N_47723);
xor UO_1988 (O_1988,N_45894,N_47851);
xor UO_1989 (O_1989,N_48085,N_45713);
or UO_1990 (O_1990,N_46570,N_46974);
or UO_1991 (O_1991,N_48021,N_46199);
or UO_1992 (O_1992,N_47053,N_48046);
or UO_1993 (O_1993,N_45666,N_49921);
nand UO_1994 (O_1994,N_46249,N_46522);
or UO_1995 (O_1995,N_45362,N_46411);
xor UO_1996 (O_1996,N_46790,N_47684);
nand UO_1997 (O_1997,N_47288,N_49097);
nor UO_1998 (O_1998,N_46022,N_47835);
xor UO_1999 (O_1999,N_47880,N_46649);
and UO_2000 (O_2000,N_46795,N_49347);
and UO_2001 (O_2001,N_45142,N_46603);
nor UO_2002 (O_2002,N_46773,N_49993);
xor UO_2003 (O_2003,N_48980,N_49031);
xor UO_2004 (O_2004,N_46473,N_47719);
nand UO_2005 (O_2005,N_46897,N_48587);
nor UO_2006 (O_2006,N_46628,N_46347);
or UO_2007 (O_2007,N_46309,N_47006);
or UO_2008 (O_2008,N_46413,N_49459);
or UO_2009 (O_2009,N_46217,N_47683);
nand UO_2010 (O_2010,N_49125,N_47096);
or UO_2011 (O_2011,N_48602,N_48833);
nor UO_2012 (O_2012,N_46996,N_48882);
or UO_2013 (O_2013,N_47005,N_48018);
and UO_2014 (O_2014,N_48798,N_49090);
and UO_2015 (O_2015,N_46610,N_45059);
nand UO_2016 (O_2016,N_46141,N_49827);
and UO_2017 (O_2017,N_46849,N_47854);
nor UO_2018 (O_2018,N_47204,N_46820);
nor UO_2019 (O_2019,N_46316,N_46995);
and UO_2020 (O_2020,N_46428,N_49588);
and UO_2021 (O_2021,N_46637,N_47646);
xor UO_2022 (O_2022,N_49752,N_47876);
or UO_2023 (O_2023,N_45449,N_46245);
nor UO_2024 (O_2024,N_49986,N_45828);
or UO_2025 (O_2025,N_47433,N_45346);
nor UO_2026 (O_2026,N_48944,N_45038);
or UO_2027 (O_2027,N_45843,N_48975);
nor UO_2028 (O_2028,N_45491,N_49247);
nand UO_2029 (O_2029,N_48302,N_46651);
nand UO_2030 (O_2030,N_49113,N_46548);
nor UO_2031 (O_2031,N_48002,N_49190);
nor UO_2032 (O_2032,N_48367,N_48282);
or UO_2033 (O_2033,N_45011,N_46751);
and UO_2034 (O_2034,N_48586,N_45691);
nand UO_2035 (O_2035,N_45670,N_48741);
or UO_2036 (O_2036,N_49536,N_48073);
nand UO_2037 (O_2037,N_49545,N_46889);
nor UO_2038 (O_2038,N_45963,N_49829);
xor UO_2039 (O_2039,N_47177,N_49139);
xnor UO_2040 (O_2040,N_49453,N_45886);
nor UO_2041 (O_2041,N_46330,N_47380);
and UO_2042 (O_2042,N_48547,N_49185);
xor UO_2043 (O_2043,N_47892,N_45005);
nor UO_2044 (O_2044,N_49307,N_48910);
nand UO_2045 (O_2045,N_47944,N_45294);
or UO_2046 (O_2046,N_46645,N_48958);
xnor UO_2047 (O_2047,N_47203,N_47725);
and UO_2048 (O_2048,N_49389,N_48305);
or UO_2049 (O_2049,N_46448,N_45965);
nand UO_2050 (O_2050,N_46979,N_46853);
and UO_2051 (O_2051,N_49094,N_45438);
xnor UO_2052 (O_2052,N_49994,N_45351);
or UO_2053 (O_2053,N_48799,N_46850);
or UO_2054 (O_2054,N_47891,N_49059);
nand UO_2055 (O_2055,N_49009,N_48862);
nor UO_2056 (O_2056,N_49806,N_48491);
and UO_2057 (O_2057,N_47732,N_46784);
and UO_2058 (O_2058,N_48810,N_45777);
and UO_2059 (O_2059,N_47816,N_45364);
nor UO_2060 (O_2060,N_48020,N_45858);
or UO_2061 (O_2061,N_47165,N_49146);
nand UO_2062 (O_2062,N_45935,N_49716);
or UO_2063 (O_2063,N_49361,N_45225);
or UO_2064 (O_2064,N_47171,N_47496);
nand UO_2065 (O_2065,N_49100,N_45753);
and UO_2066 (O_2066,N_46328,N_47346);
nor UO_2067 (O_2067,N_48641,N_49872);
or UO_2068 (O_2068,N_46884,N_48715);
nand UO_2069 (O_2069,N_49685,N_45439);
nor UO_2070 (O_2070,N_48439,N_49541);
nor UO_2071 (O_2071,N_47956,N_45202);
xnor UO_2072 (O_2072,N_49517,N_47321);
and UO_2073 (O_2073,N_47613,N_46171);
xor UO_2074 (O_2074,N_49540,N_47037);
nor UO_2075 (O_2075,N_45912,N_49575);
nand UO_2076 (O_2076,N_47556,N_45942);
and UO_2077 (O_2077,N_48411,N_45589);
or UO_2078 (O_2078,N_46993,N_48352);
xnor UO_2079 (O_2079,N_45546,N_48223);
or UO_2080 (O_2080,N_48237,N_49443);
or UO_2081 (O_2081,N_47666,N_49663);
and UO_2082 (O_2082,N_48866,N_45389);
xnor UO_2083 (O_2083,N_46264,N_49168);
or UO_2084 (O_2084,N_47793,N_47675);
or UO_2085 (O_2085,N_46800,N_46471);
and UO_2086 (O_2086,N_46178,N_48052);
xor UO_2087 (O_2087,N_45978,N_46483);
nor UO_2088 (O_2088,N_48104,N_47494);
and UO_2089 (O_2089,N_46999,N_47735);
or UO_2090 (O_2090,N_45746,N_45181);
xor UO_2091 (O_2091,N_47752,N_48144);
nor UO_2092 (O_2092,N_49115,N_47917);
xnor UO_2093 (O_2093,N_48934,N_46325);
or UO_2094 (O_2094,N_46946,N_48849);
and UO_2095 (O_2095,N_48859,N_48347);
xor UO_2096 (O_2096,N_48770,N_47426);
or UO_2097 (O_2097,N_45453,N_48108);
and UO_2098 (O_2098,N_49044,N_47105);
nand UO_2099 (O_2099,N_49633,N_49024);
or UO_2100 (O_2100,N_48896,N_47409);
nand UO_2101 (O_2101,N_47983,N_47228);
nand UO_2102 (O_2102,N_46977,N_48993);
and UO_2103 (O_2103,N_45600,N_49522);
nor UO_2104 (O_2104,N_49695,N_47133);
or UO_2105 (O_2105,N_48522,N_49196);
nand UO_2106 (O_2106,N_49705,N_48638);
xor UO_2107 (O_2107,N_49079,N_49679);
nor UO_2108 (O_2108,N_49346,N_46364);
xor UO_2109 (O_2109,N_45101,N_45305);
and UO_2110 (O_2110,N_48071,N_46859);
or UO_2111 (O_2111,N_46010,N_45241);
and UO_2112 (O_2112,N_47112,N_47924);
and UO_2113 (O_2113,N_46383,N_45444);
xor UO_2114 (O_2114,N_45008,N_46766);
or UO_2115 (O_2115,N_46679,N_48392);
nor UO_2116 (O_2116,N_48544,N_46246);
xor UO_2117 (O_2117,N_48022,N_49001);
nor UO_2118 (O_2118,N_49330,N_47848);
nor UO_2119 (O_2119,N_49434,N_46089);
or UO_2120 (O_2120,N_45417,N_48633);
nand UO_2121 (O_2121,N_47084,N_49288);
or UO_2122 (O_2122,N_45073,N_45461);
or UO_2123 (O_2123,N_48215,N_48786);
nor UO_2124 (O_2124,N_48531,N_47517);
nor UO_2125 (O_2125,N_46337,N_48789);
xnor UO_2126 (O_2126,N_48713,N_47709);
and UO_2127 (O_2127,N_49285,N_48387);
and UO_2128 (O_2128,N_49978,N_48083);
xor UO_2129 (O_2129,N_49174,N_46499);
nor UO_2130 (O_2130,N_48727,N_48946);
xor UO_2131 (O_2131,N_49992,N_48075);
and UO_2132 (O_2132,N_48824,N_48359);
and UO_2133 (O_2133,N_48688,N_45610);
xor UO_2134 (O_2134,N_45686,N_48959);
nand UO_2135 (O_2135,N_49905,N_45441);
nand UO_2136 (O_2136,N_48565,N_49936);
xnor UO_2137 (O_2137,N_49809,N_45071);
and UO_2138 (O_2138,N_46599,N_46654);
or UO_2139 (O_2139,N_48278,N_48536);
and UO_2140 (O_2140,N_45910,N_48939);
or UO_2141 (O_2141,N_46046,N_47964);
or UO_2142 (O_2142,N_49594,N_46068);
nand UO_2143 (O_2143,N_47127,N_46345);
xor UO_2144 (O_2144,N_47957,N_49417);
nor UO_2145 (O_2145,N_47403,N_47736);
xor UO_2146 (O_2146,N_45771,N_48863);
or UO_2147 (O_2147,N_47789,N_48077);
and UO_2148 (O_2148,N_49738,N_45456);
nor UO_2149 (O_2149,N_45003,N_46437);
nor UO_2150 (O_2150,N_49194,N_47982);
and UO_2151 (O_2151,N_45517,N_46292);
or UO_2152 (O_2152,N_46381,N_49560);
or UO_2153 (O_2153,N_49188,N_46925);
or UO_2154 (O_2154,N_47593,N_48634);
nor UO_2155 (O_2155,N_47597,N_48929);
or UO_2156 (O_2156,N_46844,N_45421);
nor UO_2157 (O_2157,N_49474,N_49854);
nor UO_2158 (O_2158,N_45105,N_45245);
xnor UO_2159 (O_2159,N_46436,N_48008);
xor UO_2160 (O_2160,N_48410,N_45102);
nand UO_2161 (O_2161,N_47900,N_49211);
nand UO_2162 (O_2162,N_47089,N_48187);
nand UO_2163 (O_2163,N_48635,N_49222);
or UO_2164 (O_2164,N_49845,N_47590);
and UO_2165 (O_2165,N_47297,N_47398);
nand UO_2166 (O_2166,N_45569,N_45091);
xnor UO_2167 (O_2167,N_49085,N_47488);
nor UO_2168 (O_2168,N_48675,N_46248);
xnor UO_2169 (O_2169,N_45431,N_45437);
nor UO_2170 (O_2170,N_48213,N_47512);
or UO_2171 (O_2171,N_48409,N_48628);
or UO_2172 (O_2172,N_47973,N_49033);
nand UO_2173 (O_2173,N_47604,N_46206);
nand UO_2174 (O_2174,N_48465,N_47977);
or UO_2175 (O_2175,N_45308,N_49917);
nand UO_2176 (O_2176,N_49968,N_48238);
or UO_2177 (O_2177,N_45685,N_46398);
xnor UO_2178 (O_2178,N_49372,N_48492);
or UO_2179 (O_2179,N_49166,N_45512);
xnor UO_2180 (O_2180,N_46803,N_47609);
and UO_2181 (O_2181,N_47893,N_48433);
or UO_2182 (O_2182,N_49923,N_49154);
xor UO_2183 (O_2183,N_46951,N_47065);
or UO_2184 (O_2184,N_49656,N_49253);
or UO_2185 (O_2185,N_47347,N_45372);
or UO_2186 (O_2186,N_46722,N_46551);
or UO_2187 (O_2187,N_47302,N_49147);
nand UO_2188 (O_2188,N_49276,N_46120);
nand UO_2189 (O_2189,N_47444,N_48905);
or UO_2190 (O_2190,N_49486,N_48831);
xnor UO_2191 (O_2191,N_46793,N_48876);
nor UO_2192 (O_2192,N_46382,N_45373);
xor UO_2193 (O_2193,N_47907,N_47307);
xor UO_2194 (O_2194,N_48506,N_46658);
nor UO_2195 (O_2195,N_46647,N_48870);
or UO_2196 (O_2196,N_48552,N_45743);
or UO_2197 (O_2197,N_48992,N_46713);
xor UO_2198 (O_2198,N_46212,N_46218);
or UO_2199 (O_2199,N_46114,N_49786);
nand UO_2200 (O_2200,N_47831,N_47054);
or UO_2201 (O_2201,N_45676,N_48288);
or UO_2202 (O_2202,N_45669,N_47652);
xnor UO_2203 (O_2203,N_49846,N_48480);
nand UO_2204 (O_2204,N_45303,N_47122);
and UO_2205 (O_2205,N_49478,N_46586);
and UO_2206 (O_2206,N_45605,N_45853);
or UO_2207 (O_2207,N_45643,N_45311);
nand UO_2208 (O_2208,N_46100,N_48453);
and UO_2209 (O_2209,N_47324,N_48695);
nand UO_2210 (O_2210,N_46132,N_47615);
nor UO_2211 (O_2211,N_47935,N_47245);
and UO_2212 (O_2212,N_49817,N_45836);
nor UO_2213 (O_2213,N_47056,N_49648);
nand UO_2214 (O_2214,N_46326,N_47066);
xnor UO_2215 (O_2215,N_47642,N_45190);
or UO_2216 (O_2216,N_46146,N_48791);
nor UO_2217 (O_2217,N_46947,N_47131);
xnor UO_2218 (O_2218,N_46074,N_48454);
or UO_2219 (O_2219,N_47049,N_47106);
and UO_2220 (O_2220,N_48475,N_49063);
nand UO_2221 (O_2221,N_46581,N_45174);
nor UO_2222 (O_2222,N_47952,N_46564);
nand UO_2223 (O_2223,N_46185,N_48596);
xnor UO_2224 (O_2224,N_45353,N_49238);
xnor UO_2225 (O_2225,N_47432,N_45124);
xnor UO_2226 (O_2226,N_49974,N_45509);
or UO_2227 (O_2227,N_47820,N_49177);
nor UO_2228 (O_2228,N_48229,N_45783);
nor UO_2229 (O_2229,N_48339,N_49791);
nand UO_2230 (O_2230,N_48561,N_46960);
nand UO_2231 (O_2231,N_49106,N_45827);
xnor UO_2232 (O_2232,N_49958,N_46307);
xor UO_2233 (O_2233,N_47771,N_47566);
or UO_2234 (O_2234,N_48434,N_45805);
xor UO_2235 (O_2235,N_49493,N_49535);
or UO_2236 (O_2236,N_48446,N_45973);
nor UO_2237 (O_2237,N_46832,N_45032);
or UO_2238 (O_2238,N_47931,N_48590);
nand UO_2239 (O_2239,N_49971,N_47176);
or UO_2240 (O_2240,N_45893,N_49981);
or UO_2241 (O_2241,N_46893,N_46395);
nand UO_2242 (O_2242,N_46269,N_48275);
nand UO_2243 (O_2243,N_47925,N_47242);
nor UO_2244 (O_2244,N_48154,N_49264);
xnor UO_2245 (O_2245,N_48937,N_45962);
and UO_2246 (O_2246,N_46410,N_49602);
or UO_2247 (O_2247,N_48094,N_45789);
nand UO_2248 (O_2248,N_45876,N_48087);
and UO_2249 (O_2249,N_47431,N_46682);
nor UO_2250 (O_2250,N_49985,N_48941);
nand UO_2251 (O_2251,N_48532,N_48748);
nor UO_2252 (O_2252,N_48287,N_45413);
nand UO_2253 (O_2253,N_47076,N_46239);
nand UO_2254 (O_2254,N_45794,N_46634);
or UO_2255 (O_2255,N_45394,N_45731);
nor UO_2256 (O_2256,N_47350,N_45521);
xor UO_2257 (O_2257,N_48005,N_46550);
or UO_2258 (O_2258,N_45526,N_45345);
nand UO_2259 (O_2259,N_46175,N_47672);
and UO_2260 (O_2260,N_47993,N_47411);
nor UO_2261 (O_2261,N_47271,N_46949);
or UO_2262 (O_2262,N_46936,N_48828);
nor UO_2263 (O_2263,N_45231,N_45951);
xnor UO_2264 (O_2264,N_49282,N_49579);
xor UO_2265 (O_2265,N_49518,N_45969);
or UO_2266 (O_2266,N_46051,N_49713);
xnor UO_2267 (O_2267,N_45922,N_46295);
or UO_2268 (O_2268,N_48344,N_46133);
or UO_2269 (O_2269,N_45557,N_49065);
or UO_2270 (O_2270,N_48956,N_49343);
or UO_2271 (O_2271,N_45634,N_48161);
nand UO_2272 (O_2272,N_46575,N_46052);
xnor UO_2273 (O_2273,N_46006,N_45529);
and UO_2274 (O_2274,N_45061,N_45021);
xor UO_2275 (O_2275,N_48431,N_45455);
or UO_2276 (O_2276,N_47251,N_48152);
nor UO_2277 (O_2277,N_46772,N_46184);
or UO_2278 (O_2278,N_46241,N_49903);
xor UO_2279 (O_2279,N_46828,N_46895);
nand UO_2280 (O_2280,N_47866,N_45609);
nand UO_2281 (O_2281,N_48924,N_48379);
or UO_2282 (O_2282,N_47387,N_48219);
or UO_2283 (O_2283,N_49852,N_47825);
xnor UO_2284 (O_2284,N_49898,N_46205);
xnor UO_2285 (O_2285,N_49268,N_46924);
xnor UO_2286 (O_2286,N_46420,N_45488);
nand UO_2287 (O_2287,N_46450,N_47200);
nand UO_2288 (O_2288,N_49702,N_48782);
and UO_2289 (O_2289,N_47142,N_46623);
xor UO_2290 (O_2290,N_45490,N_48852);
and UO_2291 (O_2291,N_46136,N_46737);
nand UO_2292 (O_2292,N_46026,N_45368);
nand UO_2293 (O_2293,N_46881,N_46867);
or UO_2294 (O_2294,N_45004,N_47230);
or UO_2295 (O_2295,N_45632,N_49479);
nor UO_2296 (O_2296,N_49215,N_45524);
and UO_2297 (O_2297,N_47085,N_48699);
xnor UO_2298 (O_2298,N_47960,N_45911);
nor UO_2299 (O_2299,N_45477,N_45757);
xnor UO_2300 (O_2300,N_46232,N_49948);
xor UO_2301 (O_2301,N_47336,N_46981);
or UO_2302 (O_2302,N_48515,N_47283);
xor UO_2303 (O_2303,N_49427,N_47999);
nand UO_2304 (O_2304,N_46754,N_49585);
and UO_2305 (O_2305,N_47836,N_48141);
nand UO_2306 (O_2306,N_45809,N_45549);
xnor UO_2307 (O_2307,N_49966,N_47895);
xnor UO_2308 (O_2308,N_49884,N_47837);
xor UO_2309 (O_2309,N_49083,N_47946);
and UO_2310 (O_2310,N_48259,N_45462);
nand UO_2311 (O_2311,N_48329,N_45604);
nor UO_2312 (O_2312,N_47312,N_49622);
and UO_2313 (O_2313,N_46516,N_49524);
xnor UO_2314 (O_2314,N_49155,N_49782);
nand UO_2315 (O_2315,N_47721,N_48272);
nand UO_2316 (O_2316,N_48445,N_45767);
and UO_2317 (O_2317,N_47416,N_45342);
and UO_2318 (O_2318,N_46363,N_49515);
and UO_2319 (O_2319,N_48456,N_48429);
xor UO_2320 (O_2320,N_48029,N_48846);
xnor UO_2321 (O_2321,N_48591,N_45131);
and UO_2322 (O_2322,N_45136,N_45712);
and UO_2323 (O_2323,N_46954,N_45377);
nor UO_2324 (O_2324,N_46988,N_45633);
or UO_2325 (O_2325,N_46659,N_48448);
and UO_2326 (O_2326,N_45864,N_45859);
nor UO_2327 (O_2327,N_49802,N_46701);
xnor UO_2328 (O_2328,N_47276,N_46705);
nand UO_2329 (O_2329,N_46384,N_47115);
and UO_2330 (O_2330,N_48730,N_45148);
xor UO_2331 (O_2331,N_45896,N_45596);
and UO_2332 (O_2332,N_48820,N_48670);
and UO_2333 (O_2333,N_48055,N_46842);
and UO_2334 (O_2334,N_45433,N_49566);
and UO_2335 (O_2335,N_49223,N_49437);
and UO_2336 (O_2336,N_46825,N_47208);
xnor UO_2337 (O_2337,N_45141,N_48478);
xor UO_2338 (O_2338,N_45834,N_46379);
and UO_2339 (O_2339,N_48170,N_49603);
and UO_2340 (O_2340,N_45317,N_49736);
xnor UO_2341 (O_2341,N_49582,N_47259);
xnor UO_2342 (O_2342,N_45243,N_47104);
or UO_2343 (O_2343,N_46368,N_48408);
xnor UO_2344 (O_2344,N_45266,N_48325);
or UO_2345 (O_2345,N_48407,N_46903);
xnor UO_2346 (O_2346,N_45678,N_46835);
and UO_2347 (O_2347,N_49611,N_45522);
xnor UO_2348 (O_2348,N_48557,N_48674);
and UO_2349 (O_2349,N_46126,N_49338);
and UO_2350 (O_2350,N_49151,N_48355);
nand UO_2351 (O_2351,N_48266,N_46266);
nand UO_2352 (O_2352,N_49299,N_47362);
nor UO_2353 (O_2353,N_46001,N_48369);
xor UO_2354 (O_2354,N_46461,N_47705);
or UO_2355 (O_2355,N_48436,N_48754);
xor UO_2356 (O_2356,N_48757,N_47870);
or UO_2357 (O_2357,N_45335,N_46736);
and UO_2358 (O_2358,N_46406,N_47819);
and UO_2359 (O_2359,N_47129,N_48921);
and UO_2360 (O_2360,N_48554,N_46697);
and UO_2361 (O_2361,N_46652,N_46226);
or UO_2362 (O_2362,N_48564,N_49944);
or UO_2363 (O_2363,N_46431,N_46424);
nand UO_2364 (O_2364,N_49318,N_46349);
xnor UO_2365 (O_2365,N_46079,N_49885);
and UO_2366 (O_2366,N_45157,N_48473);
nand UO_2367 (O_2367,N_48509,N_49396);
nor UO_2368 (O_2368,N_45615,N_46854);
xnor UO_2369 (O_2369,N_48712,N_45197);
xnor UO_2370 (O_2370,N_48241,N_47223);
xnor UO_2371 (O_2371,N_49056,N_45322);
and UO_2372 (O_2372,N_48070,N_49064);
nor UO_2373 (O_2373,N_49209,N_49571);
nand UO_2374 (O_2374,N_49690,N_49512);
nor UO_2375 (O_2375,N_48139,N_46822);
xnor UO_2376 (O_2376,N_47599,N_49250);
nor UO_2377 (O_2377,N_49249,N_48923);
nor UO_2378 (O_2378,N_45540,N_48177);
xnor UO_2379 (O_2379,N_47090,N_46161);
nor UO_2380 (O_2380,N_45018,N_48016);
and UO_2381 (O_2381,N_45683,N_46699);
xor UO_2382 (O_2382,N_49759,N_47108);
nand UO_2383 (O_2383,N_47442,N_47874);
and UO_2384 (O_2384,N_49425,N_47083);
nand UO_2385 (O_2385,N_45537,N_47759);
and UO_2386 (O_2386,N_45995,N_45898);
or UO_2387 (O_2387,N_48335,N_48183);
or UO_2388 (O_2388,N_46060,N_45671);
xor UO_2389 (O_2389,N_47355,N_47807);
and UO_2390 (O_2390,N_48701,N_45359);
xor UO_2391 (O_2391,N_49996,N_47943);
nand UO_2392 (O_2392,N_45165,N_46135);
or UO_2393 (O_2393,N_49134,N_49322);
or UO_2394 (O_2394,N_47700,N_49610);
or UO_2395 (O_2395,N_49617,N_49748);
and UO_2396 (O_2396,N_48256,N_46695);
nand UO_2397 (O_2397,N_45636,N_47776);
nand UO_2398 (O_2398,N_47376,N_47196);
nor UO_2399 (O_2399,N_46526,N_47596);
xor UO_2400 (O_2400,N_46781,N_45780);
xor UO_2401 (O_2401,N_48527,N_46124);
xor UO_2402 (O_2402,N_45133,N_45348);
or UO_2403 (O_2403,N_47003,N_47313);
or UO_2404 (O_2404,N_47988,N_45019);
nand UO_2405 (O_2405,N_48620,N_46305);
nand UO_2406 (O_2406,N_46512,N_46201);
nor UO_2407 (O_2407,N_46202,N_47600);
nand UO_2408 (O_2408,N_47318,N_46118);
or UO_2409 (O_2409,N_47080,N_47698);
and UO_2410 (O_2410,N_45815,N_45052);
nor UO_2411 (O_2411,N_47682,N_46617);
and UO_2412 (O_2412,N_45166,N_49779);
or UO_2413 (O_2413,N_45229,N_46607);
or UO_2414 (O_2414,N_49698,N_46170);
nor UO_2415 (O_2415,N_45006,N_48785);
nor UO_2416 (O_2416,N_47443,N_46048);
xnor UO_2417 (O_2417,N_45247,N_48656);
and UO_2418 (O_2418,N_47958,N_48763);
xor UO_2419 (O_2419,N_45986,N_49823);
or UO_2420 (O_2420,N_47111,N_46291);
xnor UO_2421 (O_2421,N_47722,N_46144);
and UO_2422 (O_2422,N_48322,N_45841);
xor UO_2423 (O_2423,N_45646,N_45284);
xnor UO_2424 (O_2424,N_47303,N_46728);
xor UO_2425 (O_2425,N_46163,N_45079);
nand UO_2426 (O_2426,N_45330,N_48840);
and UO_2427 (O_2427,N_46817,N_48268);
or UO_2428 (O_2428,N_46571,N_47069);
nor UO_2429 (O_2429,N_45991,N_47619);
nor UO_2430 (O_2430,N_45547,N_49949);
nor UO_2431 (O_2431,N_46224,N_46620);
xor UO_2432 (O_2432,N_47537,N_45855);
xnor UO_2433 (O_2433,N_45357,N_45360);
xnor UO_2434 (O_2434,N_47592,N_46321);
and UO_2435 (O_2435,N_49355,N_46190);
nor UO_2436 (O_2436,N_49510,N_49135);
nor UO_2437 (O_2437,N_46332,N_45194);
nand UO_2438 (O_2438,N_47936,N_45378);
nand UO_2439 (O_2439,N_45496,N_49335);
nand UO_2440 (O_2440,N_49160,N_45863);
nand UO_2441 (O_2441,N_45941,N_47155);
xor UO_2442 (O_2442,N_48604,N_48316);
and UO_2443 (O_2443,N_48438,N_47278);
or UO_2444 (O_2444,N_47269,N_49549);
xor UO_2445 (O_2445,N_45199,N_48725);
nand UO_2446 (O_2446,N_45796,N_46976);
nor UO_2447 (O_2447,N_47565,N_49645);
or UO_2448 (O_2448,N_45400,N_47598);
nand UO_2449 (O_2449,N_46841,N_47267);
nand UO_2450 (O_2450,N_45175,N_49105);
or UO_2451 (O_2451,N_45925,N_45823);
or UO_2452 (O_2452,N_47665,N_47451);
and UO_2453 (O_2453,N_46388,N_47539);
nor UO_2454 (O_2454,N_46885,N_48498);
or UO_2455 (O_2455,N_45548,N_45123);
or UO_2456 (O_2456,N_49070,N_46025);
nand UO_2457 (O_2457,N_47225,N_46297);
nor UO_2458 (O_2458,N_46569,N_46434);
or UO_2459 (O_2459,N_46211,N_47782);
nand UO_2460 (O_2460,N_48520,N_49251);
and UO_2461 (O_2461,N_45956,N_46648);
and UO_2462 (O_2462,N_46317,N_48524);
nor UO_2463 (O_2463,N_46811,N_45233);
nand UO_2464 (O_2464,N_47280,N_49892);
and UO_2465 (O_2465,N_49660,N_49279);
nand UO_2466 (O_2466,N_49862,N_47164);
xnor UO_2467 (O_2467,N_45467,N_47120);
or UO_2468 (O_2468,N_45909,N_45803);
xnor UO_2469 (O_2469,N_48194,N_46260);
nor UO_2470 (O_2470,N_49073,N_49213);
or UO_2471 (O_2471,N_49336,N_48893);
or UO_2472 (O_2472,N_46240,N_45207);
or UO_2473 (O_2473,N_45931,N_45556);
and UO_2474 (O_2474,N_46355,N_47464);
nor UO_2475 (O_2475,N_48353,N_49920);
or UO_2476 (O_2476,N_47534,N_46568);
nor UO_2477 (O_2477,N_48297,N_46860);
nor UO_2478 (O_2478,N_49939,N_48598);
nor UO_2479 (O_2479,N_49444,N_47584);
nor UO_2480 (O_2480,N_48574,N_45514);
nand UO_2481 (O_2481,N_47114,N_49654);
nand UO_2482 (O_2482,N_48888,N_46073);
or UO_2483 (O_2483,N_46868,N_48397);
nand UO_2484 (O_2484,N_45687,N_49112);
xnor UO_2485 (O_2485,N_48573,N_48076);
or UO_2486 (O_2486,N_45484,N_49241);
and UO_2487 (O_2487,N_48041,N_49875);
nand UO_2488 (O_2488,N_49081,N_45185);
and UO_2489 (O_2489,N_47074,N_46796);
or UO_2490 (O_2490,N_47266,N_48079);
and UO_2491 (O_2491,N_47755,N_49935);
or UO_2492 (O_2492,N_47862,N_49953);
or UO_2493 (O_2493,N_45802,N_46752);
or UO_2494 (O_2494,N_46826,N_46968);
or UO_2495 (O_2495,N_45291,N_48837);
and UO_2496 (O_2496,N_49519,N_49193);
nor UO_2497 (O_2497,N_47458,N_46274);
nand UO_2498 (O_2498,N_49455,N_48342);
nor UO_2499 (O_2499,N_46573,N_46050);
xor UO_2500 (O_2500,N_46647,N_45782);
or UO_2501 (O_2501,N_48474,N_45731);
nor UO_2502 (O_2502,N_48872,N_49342);
nor UO_2503 (O_2503,N_48374,N_47994);
xor UO_2504 (O_2504,N_49479,N_48708);
and UO_2505 (O_2505,N_49740,N_48809);
xnor UO_2506 (O_2506,N_49106,N_48398);
xor UO_2507 (O_2507,N_45628,N_46663);
xnor UO_2508 (O_2508,N_45602,N_47920);
nand UO_2509 (O_2509,N_49282,N_47889);
and UO_2510 (O_2510,N_46307,N_45317);
and UO_2511 (O_2511,N_46744,N_48808);
and UO_2512 (O_2512,N_48265,N_49970);
or UO_2513 (O_2513,N_46648,N_48984);
nand UO_2514 (O_2514,N_45333,N_48495);
or UO_2515 (O_2515,N_46219,N_45640);
xnor UO_2516 (O_2516,N_45402,N_45947);
nand UO_2517 (O_2517,N_48839,N_47044);
nor UO_2518 (O_2518,N_46930,N_47779);
nand UO_2519 (O_2519,N_45431,N_49659);
or UO_2520 (O_2520,N_49756,N_48810);
xnor UO_2521 (O_2521,N_47406,N_47999);
xor UO_2522 (O_2522,N_49691,N_48967);
or UO_2523 (O_2523,N_47948,N_46828);
xnor UO_2524 (O_2524,N_48124,N_47037);
and UO_2525 (O_2525,N_47969,N_46573);
or UO_2526 (O_2526,N_47458,N_49713);
xor UO_2527 (O_2527,N_47605,N_46465);
or UO_2528 (O_2528,N_49649,N_46512);
nor UO_2529 (O_2529,N_47373,N_47115);
or UO_2530 (O_2530,N_49228,N_49636);
and UO_2531 (O_2531,N_46275,N_46580);
nand UO_2532 (O_2532,N_49887,N_48731);
nor UO_2533 (O_2533,N_46815,N_46535);
nor UO_2534 (O_2534,N_45574,N_46663);
nor UO_2535 (O_2535,N_48506,N_49072);
or UO_2536 (O_2536,N_49619,N_48736);
or UO_2537 (O_2537,N_48410,N_45010);
xor UO_2538 (O_2538,N_48772,N_46059);
or UO_2539 (O_2539,N_45740,N_49851);
xnor UO_2540 (O_2540,N_49049,N_49261);
xor UO_2541 (O_2541,N_47735,N_48048);
nor UO_2542 (O_2542,N_46701,N_47513);
nand UO_2543 (O_2543,N_45757,N_47670);
nor UO_2544 (O_2544,N_47915,N_45870);
xor UO_2545 (O_2545,N_45250,N_49110);
and UO_2546 (O_2546,N_46548,N_49777);
and UO_2547 (O_2547,N_49969,N_49424);
or UO_2548 (O_2548,N_47570,N_49648);
nand UO_2549 (O_2549,N_48849,N_45866);
or UO_2550 (O_2550,N_49765,N_46770);
and UO_2551 (O_2551,N_49062,N_47507);
nand UO_2552 (O_2552,N_47147,N_47911);
xnor UO_2553 (O_2553,N_49368,N_46776);
nor UO_2554 (O_2554,N_47739,N_46022);
xnor UO_2555 (O_2555,N_48241,N_49144);
nor UO_2556 (O_2556,N_46009,N_46695);
nand UO_2557 (O_2557,N_46080,N_46352);
and UO_2558 (O_2558,N_47028,N_49876);
or UO_2559 (O_2559,N_48572,N_48450);
or UO_2560 (O_2560,N_47262,N_46837);
xnor UO_2561 (O_2561,N_45312,N_48498);
xnor UO_2562 (O_2562,N_45694,N_48462);
xor UO_2563 (O_2563,N_46112,N_48453);
nor UO_2564 (O_2564,N_48179,N_45107);
and UO_2565 (O_2565,N_49046,N_49495);
xnor UO_2566 (O_2566,N_45410,N_46851);
xnor UO_2567 (O_2567,N_46093,N_48168);
nor UO_2568 (O_2568,N_49433,N_46005);
and UO_2569 (O_2569,N_47780,N_49947);
xnor UO_2570 (O_2570,N_46434,N_45888);
nor UO_2571 (O_2571,N_45536,N_49478);
and UO_2572 (O_2572,N_47117,N_45578);
xnor UO_2573 (O_2573,N_45952,N_48084);
xnor UO_2574 (O_2574,N_49475,N_46883);
or UO_2575 (O_2575,N_49143,N_47519);
or UO_2576 (O_2576,N_47443,N_47907);
nor UO_2577 (O_2577,N_46768,N_49475);
nand UO_2578 (O_2578,N_48784,N_49824);
nor UO_2579 (O_2579,N_46986,N_46494);
nand UO_2580 (O_2580,N_49215,N_49865);
and UO_2581 (O_2581,N_49536,N_47063);
xnor UO_2582 (O_2582,N_47620,N_47973);
nor UO_2583 (O_2583,N_49005,N_48059);
and UO_2584 (O_2584,N_49018,N_45048);
nand UO_2585 (O_2585,N_47801,N_49787);
xor UO_2586 (O_2586,N_47653,N_47792);
and UO_2587 (O_2587,N_45550,N_48695);
nor UO_2588 (O_2588,N_48769,N_45229);
nand UO_2589 (O_2589,N_47262,N_45127);
or UO_2590 (O_2590,N_49181,N_49402);
nand UO_2591 (O_2591,N_48186,N_47923);
and UO_2592 (O_2592,N_48332,N_46521);
nand UO_2593 (O_2593,N_45611,N_49900);
and UO_2594 (O_2594,N_48936,N_47363);
or UO_2595 (O_2595,N_47740,N_47710);
nor UO_2596 (O_2596,N_45300,N_45547);
and UO_2597 (O_2597,N_48393,N_47575);
xor UO_2598 (O_2598,N_46811,N_49119);
and UO_2599 (O_2599,N_48687,N_48638);
and UO_2600 (O_2600,N_45881,N_45736);
xnor UO_2601 (O_2601,N_45142,N_49051);
or UO_2602 (O_2602,N_46354,N_49140);
xnor UO_2603 (O_2603,N_48282,N_45104);
xnor UO_2604 (O_2604,N_46144,N_49581);
nor UO_2605 (O_2605,N_48919,N_49013);
and UO_2606 (O_2606,N_47233,N_46130);
xnor UO_2607 (O_2607,N_47900,N_48544);
xnor UO_2608 (O_2608,N_48675,N_46290);
xor UO_2609 (O_2609,N_45209,N_46077);
and UO_2610 (O_2610,N_47119,N_47988);
nand UO_2611 (O_2611,N_48495,N_46916);
nor UO_2612 (O_2612,N_49956,N_45865);
nand UO_2613 (O_2613,N_46685,N_45951);
and UO_2614 (O_2614,N_49795,N_49614);
xor UO_2615 (O_2615,N_49184,N_46481);
nor UO_2616 (O_2616,N_46225,N_47076);
nor UO_2617 (O_2617,N_48483,N_46169);
and UO_2618 (O_2618,N_46928,N_46132);
xnor UO_2619 (O_2619,N_46881,N_45720);
nor UO_2620 (O_2620,N_48489,N_47092);
and UO_2621 (O_2621,N_48911,N_48967);
or UO_2622 (O_2622,N_48829,N_49555);
nand UO_2623 (O_2623,N_48307,N_46155);
nor UO_2624 (O_2624,N_45075,N_47923);
xor UO_2625 (O_2625,N_49126,N_49206);
and UO_2626 (O_2626,N_45787,N_47649);
xor UO_2627 (O_2627,N_49092,N_46755);
nand UO_2628 (O_2628,N_48966,N_48113);
nor UO_2629 (O_2629,N_45435,N_47333);
and UO_2630 (O_2630,N_46381,N_49417);
or UO_2631 (O_2631,N_46699,N_46230);
nor UO_2632 (O_2632,N_45945,N_48096);
nand UO_2633 (O_2633,N_45004,N_49242);
nor UO_2634 (O_2634,N_47116,N_49279);
or UO_2635 (O_2635,N_48457,N_47777);
nand UO_2636 (O_2636,N_48828,N_45279);
and UO_2637 (O_2637,N_45181,N_46367);
nand UO_2638 (O_2638,N_48326,N_48587);
and UO_2639 (O_2639,N_45244,N_45243);
and UO_2640 (O_2640,N_46859,N_49760);
xnor UO_2641 (O_2641,N_47019,N_45763);
or UO_2642 (O_2642,N_47716,N_46197);
or UO_2643 (O_2643,N_46113,N_47801);
and UO_2644 (O_2644,N_48955,N_45165);
nor UO_2645 (O_2645,N_45996,N_47240);
nand UO_2646 (O_2646,N_45687,N_46249);
nor UO_2647 (O_2647,N_47545,N_47966);
nor UO_2648 (O_2648,N_46512,N_46734);
nor UO_2649 (O_2649,N_46440,N_49208);
or UO_2650 (O_2650,N_48367,N_46919);
nand UO_2651 (O_2651,N_46649,N_49055);
nand UO_2652 (O_2652,N_49810,N_45321);
or UO_2653 (O_2653,N_45971,N_47249);
or UO_2654 (O_2654,N_48575,N_48939);
xnor UO_2655 (O_2655,N_48202,N_48677);
nor UO_2656 (O_2656,N_46707,N_48708);
nor UO_2657 (O_2657,N_45803,N_48723);
xor UO_2658 (O_2658,N_45402,N_47891);
nand UO_2659 (O_2659,N_49827,N_47728);
nand UO_2660 (O_2660,N_45316,N_45100);
xnor UO_2661 (O_2661,N_49717,N_49468);
or UO_2662 (O_2662,N_48121,N_45775);
xor UO_2663 (O_2663,N_46486,N_48760);
nand UO_2664 (O_2664,N_48113,N_47985);
or UO_2665 (O_2665,N_47666,N_48834);
and UO_2666 (O_2666,N_47687,N_46664);
nand UO_2667 (O_2667,N_46616,N_49395);
or UO_2668 (O_2668,N_49987,N_48285);
or UO_2669 (O_2669,N_45481,N_47339);
nand UO_2670 (O_2670,N_47702,N_48099);
xnor UO_2671 (O_2671,N_48723,N_46700);
and UO_2672 (O_2672,N_46500,N_47728);
nor UO_2673 (O_2673,N_47831,N_48609);
nand UO_2674 (O_2674,N_45343,N_47095);
xnor UO_2675 (O_2675,N_48096,N_45293);
and UO_2676 (O_2676,N_45738,N_48433);
nor UO_2677 (O_2677,N_47217,N_46470);
nand UO_2678 (O_2678,N_47545,N_46758);
or UO_2679 (O_2679,N_47533,N_47938);
xor UO_2680 (O_2680,N_45251,N_48864);
or UO_2681 (O_2681,N_45283,N_45630);
and UO_2682 (O_2682,N_47287,N_48568);
xnor UO_2683 (O_2683,N_48587,N_46675);
nand UO_2684 (O_2684,N_45555,N_45683);
nor UO_2685 (O_2685,N_47627,N_48090);
xor UO_2686 (O_2686,N_48585,N_49499);
xor UO_2687 (O_2687,N_46383,N_45710);
nor UO_2688 (O_2688,N_45192,N_46686);
xnor UO_2689 (O_2689,N_47134,N_49313);
nand UO_2690 (O_2690,N_45919,N_49649);
nor UO_2691 (O_2691,N_48046,N_49611);
or UO_2692 (O_2692,N_45796,N_48716);
nor UO_2693 (O_2693,N_45324,N_49928);
xor UO_2694 (O_2694,N_47603,N_49346);
nand UO_2695 (O_2695,N_45870,N_49938);
nand UO_2696 (O_2696,N_46808,N_47180);
xor UO_2697 (O_2697,N_47278,N_46979);
xor UO_2698 (O_2698,N_45345,N_47542);
and UO_2699 (O_2699,N_47367,N_46148);
and UO_2700 (O_2700,N_45596,N_45110);
and UO_2701 (O_2701,N_49236,N_47670);
and UO_2702 (O_2702,N_47108,N_46743);
and UO_2703 (O_2703,N_47632,N_47885);
nor UO_2704 (O_2704,N_45018,N_49323);
nand UO_2705 (O_2705,N_49570,N_46576);
or UO_2706 (O_2706,N_47188,N_48529);
or UO_2707 (O_2707,N_47202,N_47979);
and UO_2708 (O_2708,N_45124,N_47350);
nand UO_2709 (O_2709,N_45247,N_49476);
nand UO_2710 (O_2710,N_48345,N_47632);
nand UO_2711 (O_2711,N_48400,N_48596);
or UO_2712 (O_2712,N_48133,N_48393);
and UO_2713 (O_2713,N_46263,N_47217);
and UO_2714 (O_2714,N_49856,N_47402);
xnor UO_2715 (O_2715,N_47640,N_46808);
nor UO_2716 (O_2716,N_49286,N_45976);
nand UO_2717 (O_2717,N_46117,N_47585);
xnor UO_2718 (O_2718,N_46791,N_49726);
nor UO_2719 (O_2719,N_49443,N_47632);
or UO_2720 (O_2720,N_47527,N_49990);
and UO_2721 (O_2721,N_49904,N_49134);
and UO_2722 (O_2722,N_49378,N_47926);
nor UO_2723 (O_2723,N_46679,N_48249);
nor UO_2724 (O_2724,N_49057,N_49641);
and UO_2725 (O_2725,N_45952,N_45833);
nand UO_2726 (O_2726,N_49662,N_48828);
nor UO_2727 (O_2727,N_47230,N_48357);
nand UO_2728 (O_2728,N_46146,N_47009);
nor UO_2729 (O_2729,N_46189,N_46361);
xnor UO_2730 (O_2730,N_45260,N_45139);
and UO_2731 (O_2731,N_48018,N_45233);
and UO_2732 (O_2732,N_46943,N_45069);
and UO_2733 (O_2733,N_47982,N_47328);
nand UO_2734 (O_2734,N_49626,N_48178);
nor UO_2735 (O_2735,N_48037,N_48185);
or UO_2736 (O_2736,N_49065,N_48732);
xor UO_2737 (O_2737,N_49919,N_49204);
xor UO_2738 (O_2738,N_47109,N_49910);
or UO_2739 (O_2739,N_47931,N_49870);
xor UO_2740 (O_2740,N_47230,N_47869);
xnor UO_2741 (O_2741,N_49107,N_45180);
xor UO_2742 (O_2742,N_49205,N_46597);
nand UO_2743 (O_2743,N_46172,N_49607);
xnor UO_2744 (O_2744,N_45927,N_48198);
xnor UO_2745 (O_2745,N_48493,N_46161);
or UO_2746 (O_2746,N_45158,N_48015);
xnor UO_2747 (O_2747,N_49089,N_46773);
xnor UO_2748 (O_2748,N_45802,N_47287);
and UO_2749 (O_2749,N_48426,N_49921);
xor UO_2750 (O_2750,N_48471,N_46904);
xor UO_2751 (O_2751,N_45529,N_48770);
nand UO_2752 (O_2752,N_46377,N_48906);
nor UO_2753 (O_2753,N_47887,N_49114);
and UO_2754 (O_2754,N_47759,N_45330);
nor UO_2755 (O_2755,N_46885,N_48921);
nor UO_2756 (O_2756,N_47366,N_48607);
nand UO_2757 (O_2757,N_49474,N_49081);
nor UO_2758 (O_2758,N_48224,N_49925);
or UO_2759 (O_2759,N_46989,N_45800);
and UO_2760 (O_2760,N_48551,N_45661);
or UO_2761 (O_2761,N_47000,N_48236);
nand UO_2762 (O_2762,N_49386,N_49384);
xnor UO_2763 (O_2763,N_48972,N_49671);
xnor UO_2764 (O_2764,N_46137,N_47781);
and UO_2765 (O_2765,N_45666,N_47421);
or UO_2766 (O_2766,N_48460,N_49341);
nor UO_2767 (O_2767,N_47220,N_46507);
nor UO_2768 (O_2768,N_45171,N_49963);
nor UO_2769 (O_2769,N_47486,N_49471);
nand UO_2770 (O_2770,N_46778,N_48094);
or UO_2771 (O_2771,N_47493,N_45570);
and UO_2772 (O_2772,N_45362,N_47745);
xnor UO_2773 (O_2773,N_49800,N_46792);
or UO_2774 (O_2774,N_47550,N_46628);
nor UO_2775 (O_2775,N_46671,N_45017);
nor UO_2776 (O_2776,N_47032,N_46632);
nand UO_2777 (O_2777,N_47145,N_45071);
xnor UO_2778 (O_2778,N_46190,N_47394);
nor UO_2779 (O_2779,N_47946,N_46885);
nor UO_2780 (O_2780,N_46086,N_47144);
or UO_2781 (O_2781,N_49602,N_47912);
and UO_2782 (O_2782,N_49315,N_47076);
or UO_2783 (O_2783,N_45127,N_46609);
nand UO_2784 (O_2784,N_47813,N_47302);
nand UO_2785 (O_2785,N_49488,N_45343);
nand UO_2786 (O_2786,N_46799,N_48689);
and UO_2787 (O_2787,N_46482,N_47603);
or UO_2788 (O_2788,N_48197,N_46200);
nand UO_2789 (O_2789,N_47796,N_47159);
xor UO_2790 (O_2790,N_48472,N_47532);
nand UO_2791 (O_2791,N_48445,N_49276);
nand UO_2792 (O_2792,N_48834,N_47542);
xor UO_2793 (O_2793,N_48861,N_47913);
and UO_2794 (O_2794,N_45783,N_47504);
nor UO_2795 (O_2795,N_48247,N_49219);
nor UO_2796 (O_2796,N_45119,N_45756);
and UO_2797 (O_2797,N_48497,N_45633);
nand UO_2798 (O_2798,N_46113,N_47057);
xnor UO_2799 (O_2799,N_45646,N_46710);
or UO_2800 (O_2800,N_48034,N_47997);
nand UO_2801 (O_2801,N_49609,N_48998);
and UO_2802 (O_2802,N_46272,N_45362);
nand UO_2803 (O_2803,N_46918,N_48467);
and UO_2804 (O_2804,N_46461,N_49480);
xnor UO_2805 (O_2805,N_46625,N_45894);
and UO_2806 (O_2806,N_49820,N_45249);
nor UO_2807 (O_2807,N_46685,N_47615);
or UO_2808 (O_2808,N_45694,N_48468);
nand UO_2809 (O_2809,N_45616,N_47600);
nand UO_2810 (O_2810,N_48346,N_47521);
and UO_2811 (O_2811,N_45772,N_45495);
or UO_2812 (O_2812,N_46718,N_48933);
nor UO_2813 (O_2813,N_45463,N_47008);
nor UO_2814 (O_2814,N_45895,N_48538);
and UO_2815 (O_2815,N_49547,N_45302);
nor UO_2816 (O_2816,N_46229,N_49130);
nand UO_2817 (O_2817,N_49969,N_48449);
and UO_2818 (O_2818,N_48807,N_47355);
nand UO_2819 (O_2819,N_45008,N_48102);
xnor UO_2820 (O_2820,N_46251,N_45079);
nor UO_2821 (O_2821,N_46830,N_47384);
or UO_2822 (O_2822,N_46757,N_49432);
nor UO_2823 (O_2823,N_49680,N_45809);
or UO_2824 (O_2824,N_49615,N_47784);
and UO_2825 (O_2825,N_46834,N_49268);
xnor UO_2826 (O_2826,N_49965,N_45259);
and UO_2827 (O_2827,N_45001,N_49292);
or UO_2828 (O_2828,N_49026,N_47469);
and UO_2829 (O_2829,N_47681,N_46082);
xor UO_2830 (O_2830,N_49875,N_46711);
or UO_2831 (O_2831,N_49296,N_46416);
xor UO_2832 (O_2832,N_49187,N_49761);
or UO_2833 (O_2833,N_46117,N_46094);
and UO_2834 (O_2834,N_47902,N_49005);
and UO_2835 (O_2835,N_47181,N_46196);
nand UO_2836 (O_2836,N_48676,N_47509);
or UO_2837 (O_2837,N_45951,N_46537);
nor UO_2838 (O_2838,N_45912,N_49485);
and UO_2839 (O_2839,N_48885,N_46267);
nor UO_2840 (O_2840,N_46375,N_45485);
nor UO_2841 (O_2841,N_45974,N_49940);
nand UO_2842 (O_2842,N_47539,N_45663);
nor UO_2843 (O_2843,N_45155,N_45305);
and UO_2844 (O_2844,N_45195,N_45904);
or UO_2845 (O_2845,N_45122,N_45693);
or UO_2846 (O_2846,N_45217,N_49021);
nor UO_2847 (O_2847,N_45424,N_45867);
or UO_2848 (O_2848,N_48693,N_47660);
xnor UO_2849 (O_2849,N_45489,N_49436);
xor UO_2850 (O_2850,N_49678,N_45821);
and UO_2851 (O_2851,N_49006,N_49124);
xor UO_2852 (O_2852,N_49651,N_45946);
and UO_2853 (O_2853,N_48236,N_48397);
or UO_2854 (O_2854,N_45031,N_47986);
or UO_2855 (O_2855,N_45369,N_47931);
xnor UO_2856 (O_2856,N_47384,N_49474);
xor UO_2857 (O_2857,N_49634,N_49016);
and UO_2858 (O_2858,N_48187,N_48962);
or UO_2859 (O_2859,N_46773,N_47742);
and UO_2860 (O_2860,N_48694,N_48047);
nand UO_2861 (O_2861,N_48845,N_47422);
and UO_2862 (O_2862,N_48439,N_45415);
nand UO_2863 (O_2863,N_46060,N_47339);
xnor UO_2864 (O_2864,N_48172,N_49488);
or UO_2865 (O_2865,N_49427,N_48904);
nor UO_2866 (O_2866,N_45007,N_45837);
xor UO_2867 (O_2867,N_48804,N_45396);
or UO_2868 (O_2868,N_47709,N_45783);
xor UO_2869 (O_2869,N_47998,N_47727);
and UO_2870 (O_2870,N_49718,N_47500);
nand UO_2871 (O_2871,N_45604,N_46057);
nor UO_2872 (O_2872,N_49347,N_47315);
or UO_2873 (O_2873,N_46553,N_47266);
xnor UO_2874 (O_2874,N_45237,N_48239);
xnor UO_2875 (O_2875,N_48605,N_49747);
nand UO_2876 (O_2876,N_46718,N_49292);
and UO_2877 (O_2877,N_47059,N_46564);
nor UO_2878 (O_2878,N_47436,N_49676);
or UO_2879 (O_2879,N_49735,N_48532);
and UO_2880 (O_2880,N_45413,N_46808);
xnor UO_2881 (O_2881,N_46519,N_48810);
xnor UO_2882 (O_2882,N_48864,N_48818);
nor UO_2883 (O_2883,N_45952,N_49534);
xor UO_2884 (O_2884,N_47105,N_46098);
nand UO_2885 (O_2885,N_47101,N_46269);
nor UO_2886 (O_2886,N_48538,N_46205);
nand UO_2887 (O_2887,N_47838,N_47871);
and UO_2888 (O_2888,N_48185,N_49039);
nor UO_2889 (O_2889,N_46613,N_47667);
xnor UO_2890 (O_2890,N_45728,N_46834);
or UO_2891 (O_2891,N_49687,N_45641);
nand UO_2892 (O_2892,N_46996,N_48841);
or UO_2893 (O_2893,N_48788,N_45610);
and UO_2894 (O_2894,N_46922,N_46412);
or UO_2895 (O_2895,N_45876,N_45495);
or UO_2896 (O_2896,N_48544,N_46606);
xor UO_2897 (O_2897,N_47985,N_45488);
nand UO_2898 (O_2898,N_48245,N_49171);
nor UO_2899 (O_2899,N_45802,N_46330);
xnor UO_2900 (O_2900,N_47070,N_45771);
xnor UO_2901 (O_2901,N_49817,N_46790);
nand UO_2902 (O_2902,N_48443,N_45612);
nand UO_2903 (O_2903,N_48716,N_45082);
nand UO_2904 (O_2904,N_49987,N_45292);
nor UO_2905 (O_2905,N_48611,N_45948);
nand UO_2906 (O_2906,N_47484,N_46039);
and UO_2907 (O_2907,N_46912,N_48403);
or UO_2908 (O_2908,N_47523,N_49161);
xnor UO_2909 (O_2909,N_48049,N_47539);
nand UO_2910 (O_2910,N_47459,N_49033);
xnor UO_2911 (O_2911,N_49111,N_49722);
nand UO_2912 (O_2912,N_47580,N_48214);
nor UO_2913 (O_2913,N_47760,N_45996);
nor UO_2914 (O_2914,N_48135,N_49213);
nor UO_2915 (O_2915,N_46027,N_46356);
or UO_2916 (O_2916,N_49216,N_46213);
nand UO_2917 (O_2917,N_48287,N_48917);
and UO_2918 (O_2918,N_48519,N_47779);
nand UO_2919 (O_2919,N_48945,N_49041);
xnor UO_2920 (O_2920,N_49072,N_48199);
xor UO_2921 (O_2921,N_48466,N_48558);
or UO_2922 (O_2922,N_49881,N_48949);
or UO_2923 (O_2923,N_45966,N_46055);
nor UO_2924 (O_2924,N_45417,N_49426);
or UO_2925 (O_2925,N_46640,N_46744);
or UO_2926 (O_2926,N_49517,N_45529);
or UO_2927 (O_2927,N_46728,N_46031);
and UO_2928 (O_2928,N_48113,N_47304);
nand UO_2929 (O_2929,N_45075,N_46639);
nand UO_2930 (O_2930,N_45309,N_46749);
nor UO_2931 (O_2931,N_47906,N_45332);
nor UO_2932 (O_2932,N_45179,N_45525);
xor UO_2933 (O_2933,N_49601,N_47285);
or UO_2934 (O_2934,N_47837,N_48251);
xnor UO_2935 (O_2935,N_49031,N_49264);
and UO_2936 (O_2936,N_45595,N_48495);
or UO_2937 (O_2937,N_46798,N_48272);
nor UO_2938 (O_2938,N_49579,N_48173);
nand UO_2939 (O_2939,N_47687,N_47011);
and UO_2940 (O_2940,N_46603,N_49757);
and UO_2941 (O_2941,N_48222,N_45133);
nor UO_2942 (O_2942,N_46308,N_48591);
or UO_2943 (O_2943,N_47932,N_49233);
nor UO_2944 (O_2944,N_46874,N_49618);
or UO_2945 (O_2945,N_46211,N_46710);
and UO_2946 (O_2946,N_45317,N_45886);
nand UO_2947 (O_2947,N_46739,N_45134);
nor UO_2948 (O_2948,N_48036,N_45611);
and UO_2949 (O_2949,N_49210,N_47431);
or UO_2950 (O_2950,N_45657,N_46071);
or UO_2951 (O_2951,N_47881,N_47876);
or UO_2952 (O_2952,N_45306,N_49925);
nor UO_2953 (O_2953,N_45760,N_47024);
nand UO_2954 (O_2954,N_46121,N_48237);
nor UO_2955 (O_2955,N_46362,N_49615);
nor UO_2956 (O_2956,N_47829,N_49362);
nor UO_2957 (O_2957,N_49517,N_47650);
and UO_2958 (O_2958,N_46865,N_47891);
and UO_2959 (O_2959,N_45950,N_47958);
xor UO_2960 (O_2960,N_48691,N_46713);
xnor UO_2961 (O_2961,N_46315,N_47912);
or UO_2962 (O_2962,N_47444,N_49083);
nand UO_2963 (O_2963,N_48782,N_45388);
nand UO_2964 (O_2964,N_48406,N_46917);
and UO_2965 (O_2965,N_47916,N_49233);
and UO_2966 (O_2966,N_49721,N_46901);
or UO_2967 (O_2967,N_48172,N_49661);
and UO_2968 (O_2968,N_48201,N_48272);
nor UO_2969 (O_2969,N_48734,N_46001);
nand UO_2970 (O_2970,N_49158,N_46830);
and UO_2971 (O_2971,N_45513,N_48306);
nor UO_2972 (O_2972,N_45002,N_46525);
nand UO_2973 (O_2973,N_47443,N_45885);
xor UO_2974 (O_2974,N_45615,N_46868);
nand UO_2975 (O_2975,N_45024,N_48372);
and UO_2976 (O_2976,N_47653,N_46404);
nand UO_2977 (O_2977,N_45905,N_46792);
nand UO_2978 (O_2978,N_47149,N_45672);
or UO_2979 (O_2979,N_45370,N_46169);
xnor UO_2980 (O_2980,N_46566,N_46107);
nor UO_2981 (O_2981,N_48459,N_45607);
and UO_2982 (O_2982,N_48893,N_45492);
nand UO_2983 (O_2983,N_46482,N_45836);
nand UO_2984 (O_2984,N_49129,N_47503);
or UO_2985 (O_2985,N_47552,N_46709);
nand UO_2986 (O_2986,N_47133,N_48754);
or UO_2987 (O_2987,N_48274,N_46365);
nand UO_2988 (O_2988,N_47398,N_47388);
xor UO_2989 (O_2989,N_45165,N_48861);
or UO_2990 (O_2990,N_46226,N_49134);
xnor UO_2991 (O_2991,N_46667,N_46497);
xor UO_2992 (O_2992,N_45928,N_48986);
and UO_2993 (O_2993,N_48264,N_45986);
and UO_2994 (O_2994,N_45300,N_46889);
or UO_2995 (O_2995,N_48815,N_46039);
nand UO_2996 (O_2996,N_45142,N_47504);
nor UO_2997 (O_2997,N_49137,N_49983);
nor UO_2998 (O_2998,N_46278,N_49279);
nand UO_2999 (O_2999,N_47444,N_46188);
and UO_3000 (O_3000,N_48639,N_47539);
and UO_3001 (O_3001,N_48174,N_48787);
or UO_3002 (O_3002,N_47531,N_48568);
or UO_3003 (O_3003,N_46403,N_48658);
nor UO_3004 (O_3004,N_48481,N_47322);
and UO_3005 (O_3005,N_48692,N_48491);
nand UO_3006 (O_3006,N_47860,N_45797);
or UO_3007 (O_3007,N_47297,N_45077);
or UO_3008 (O_3008,N_49758,N_46711);
and UO_3009 (O_3009,N_46430,N_47641);
or UO_3010 (O_3010,N_46415,N_47396);
or UO_3011 (O_3011,N_46910,N_48436);
nand UO_3012 (O_3012,N_46701,N_46394);
nor UO_3013 (O_3013,N_46278,N_45802);
or UO_3014 (O_3014,N_48017,N_49571);
nor UO_3015 (O_3015,N_47986,N_49258);
nor UO_3016 (O_3016,N_49468,N_49984);
or UO_3017 (O_3017,N_45455,N_45688);
xnor UO_3018 (O_3018,N_47028,N_46299);
nand UO_3019 (O_3019,N_48707,N_49672);
nand UO_3020 (O_3020,N_49381,N_46559);
nand UO_3021 (O_3021,N_48561,N_46582);
and UO_3022 (O_3022,N_48088,N_46205);
and UO_3023 (O_3023,N_48637,N_47787);
or UO_3024 (O_3024,N_49731,N_49863);
nand UO_3025 (O_3025,N_46511,N_46507);
and UO_3026 (O_3026,N_48100,N_48171);
or UO_3027 (O_3027,N_45502,N_49304);
or UO_3028 (O_3028,N_45046,N_49285);
and UO_3029 (O_3029,N_46081,N_49811);
and UO_3030 (O_3030,N_47074,N_48226);
or UO_3031 (O_3031,N_48634,N_45486);
and UO_3032 (O_3032,N_47994,N_49196);
or UO_3033 (O_3033,N_46824,N_46936);
nor UO_3034 (O_3034,N_47961,N_45503);
or UO_3035 (O_3035,N_49994,N_49043);
and UO_3036 (O_3036,N_49198,N_49814);
or UO_3037 (O_3037,N_49613,N_49344);
xnor UO_3038 (O_3038,N_47217,N_45044);
xnor UO_3039 (O_3039,N_46843,N_49700);
xor UO_3040 (O_3040,N_48844,N_46404);
xor UO_3041 (O_3041,N_47299,N_48042);
xnor UO_3042 (O_3042,N_49856,N_47842);
nand UO_3043 (O_3043,N_45705,N_48162);
xor UO_3044 (O_3044,N_49672,N_46436);
nand UO_3045 (O_3045,N_47514,N_45521);
nand UO_3046 (O_3046,N_46595,N_45999);
xnor UO_3047 (O_3047,N_48939,N_49013);
xnor UO_3048 (O_3048,N_49529,N_49188);
nand UO_3049 (O_3049,N_45617,N_46867);
or UO_3050 (O_3050,N_45895,N_46442);
xnor UO_3051 (O_3051,N_49903,N_46103);
xnor UO_3052 (O_3052,N_45045,N_48409);
xnor UO_3053 (O_3053,N_45996,N_47887);
nor UO_3054 (O_3054,N_49546,N_45561);
nand UO_3055 (O_3055,N_45226,N_47723);
and UO_3056 (O_3056,N_49423,N_45496);
xor UO_3057 (O_3057,N_45123,N_45938);
or UO_3058 (O_3058,N_46126,N_46226);
nand UO_3059 (O_3059,N_48647,N_45429);
and UO_3060 (O_3060,N_47935,N_46341);
nor UO_3061 (O_3061,N_47839,N_48556);
xor UO_3062 (O_3062,N_46969,N_45041);
nor UO_3063 (O_3063,N_48606,N_46021);
nand UO_3064 (O_3064,N_45380,N_48259);
nor UO_3065 (O_3065,N_47978,N_46254);
and UO_3066 (O_3066,N_49069,N_46489);
xnor UO_3067 (O_3067,N_45327,N_48659);
or UO_3068 (O_3068,N_47264,N_47737);
and UO_3069 (O_3069,N_46452,N_49735);
xnor UO_3070 (O_3070,N_49066,N_46450);
xnor UO_3071 (O_3071,N_49320,N_46164);
nand UO_3072 (O_3072,N_46007,N_48403);
nand UO_3073 (O_3073,N_49291,N_45655);
xor UO_3074 (O_3074,N_48722,N_47306);
nand UO_3075 (O_3075,N_46077,N_45785);
nand UO_3076 (O_3076,N_45131,N_49133);
and UO_3077 (O_3077,N_45242,N_45243);
and UO_3078 (O_3078,N_48479,N_45274);
nand UO_3079 (O_3079,N_45555,N_47473);
and UO_3080 (O_3080,N_48225,N_46484);
and UO_3081 (O_3081,N_48847,N_48562);
nor UO_3082 (O_3082,N_48059,N_48531);
and UO_3083 (O_3083,N_48341,N_49649);
or UO_3084 (O_3084,N_48644,N_49145);
or UO_3085 (O_3085,N_48108,N_45300);
or UO_3086 (O_3086,N_46449,N_49431);
xor UO_3087 (O_3087,N_48246,N_49723);
or UO_3088 (O_3088,N_49484,N_45318);
xnor UO_3089 (O_3089,N_48977,N_46853);
or UO_3090 (O_3090,N_48485,N_49686);
nand UO_3091 (O_3091,N_49229,N_49292);
nor UO_3092 (O_3092,N_46720,N_46510);
xor UO_3093 (O_3093,N_47853,N_48593);
nand UO_3094 (O_3094,N_47095,N_47793);
nand UO_3095 (O_3095,N_49912,N_49541);
nor UO_3096 (O_3096,N_46591,N_46599);
nor UO_3097 (O_3097,N_45649,N_49734);
or UO_3098 (O_3098,N_46431,N_49381);
nor UO_3099 (O_3099,N_48417,N_47827);
nor UO_3100 (O_3100,N_45477,N_47987);
and UO_3101 (O_3101,N_48963,N_46237);
nand UO_3102 (O_3102,N_48863,N_47483);
or UO_3103 (O_3103,N_48657,N_49464);
nor UO_3104 (O_3104,N_49495,N_45114);
or UO_3105 (O_3105,N_48898,N_49587);
and UO_3106 (O_3106,N_48366,N_48253);
or UO_3107 (O_3107,N_45077,N_49033);
xnor UO_3108 (O_3108,N_47254,N_45032);
xor UO_3109 (O_3109,N_46127,N_47838);
or UO_3110 (O_3110,N_46649,N_48297);
nand UO_3111 (O_3111,N_45700,N_47878);
and UO_3112 (O_3112,N_47397,N_48691);
nand UO_3113 (O_3113,N_47273,N_47221);
and UO_3114 (O_3114,N_45199,N_46850);
nor UO_3115 (O_3115,N_47967,N_48690);
nand UO_3116 (O_3116,N_49316,N_45016);
xor UO_3117 (O_3117,N_47678,N_49701);
or UO_3118 (O_3118,N_48563,N_49953);
or UO_3119 (O_3119,N_45062,N_46084);
or UO_3120 (O_3120,N_45224,N_45557);
nor UO_3121 (O_3121,N_48928,N_47338);
nor UO_3122 (O_3122,N_45592,N_45423);
or UO_3123 (O_3123,N_46293,N_47195);
and UO_3124 (O_3124,N_49375,N_48092);
or UO_3125 (O_3125,N_49378,N_47842);
and UO_3126 (O_3126,N_48520,N_45349);
nand UO_3127 (O_3127,N_46175,N_46349);
xor UO_3128 (O_3128,N_46622,N_48731);
nor UO_3129 (O_3129,N_47232,N_48523);
or UO_3130 (O_3130,N_49093,N_46342);
and UO_3131 (O_3131,N_49215,N_49474);
nor UO_3132 (O_3132,N_47280,N_48880);
or UO_3133 (O_3133,N_48996,N_49790);
nor UO_3134 (O_3134,N_45008,N_45713);
xor UO_3135 (O_3135,N_46354,N_48124);
nand UO_3136 (O_3136,N_47155,N_45084);
nor UO_3137 (O_3137,N_46040,N_47492);
and UO_3138 (O_3138,N_46817,N_48436);
xor UO_3139 (O_3139,N_48917,N_48332);
nand UO_3140 (O_3140,N_48568,N_46815);
xnor UO_3141 (O_3141,N_47425,N_45953);
nor UO_3142 (O_3142,N_48028,N_47097);
nor UO_3143 (O_3143,N_45987,N_47365);
or UO_3144 (O_3144,N_45117,N_45173);
nand UO_3145 (O_3145,N_47961,N_47641);
nor UO_3146 (O_3146,N_46896,N_48385);
nor UO_3147 (O_3147,N_47611,N_45760);
nor UO_3148 (O_3148,N_45690,N_47869);
or UO_3149 (O_3149,N_47807,N_48644);
nor UO_3150 (O_3150,N_48254,N_46410);
nand UO_3151 (O_3151,N_46401,N_47339);
and UO_3152 (O_3152,N_45165,N_45774);
nor UO_3153 (O_3153,N_49402,N_45261);
nand UO_3154 (O_3154,N_47303,N_47085);
nand UO_3155 (O_3155,N_47904,N_49813);
and UO_3156 (O_3156,N_48859,N_47310);
nor UO_3157 (O_3157,N_49443,N_46384);
nand UO_3158 (O_3158,N_47000,N_46797);
and UO_3159 (O_3159,N_46901,N_45368);
or UO_3160 (O_3160,N_48511,N_49170);
xnor UO_3161 (O_3161,N_45146,N_46920);
nor UO_3162 (O_3162,N_49704,N_48693);
nor UO_3163 (O_3163,N_49469,N_46167);
or UO_3164 (O_3164,N_47213,N_49805);
xnor UO_3165 (O_3165,N_46805,N_49825);
or UO_3166 (O_3166,N_45427,N_49586);
and UO_3167 (O_3167,N_45313,N_47620);
nor UO_3168 (O_3168,N_48331,N_45598);
and UO_3169 (O_3169,N_49666,N_45780);
xnor UO_3170 (O_3170,N_49341,N_48202);
nor UO_3171 (O_3171,N_48609,N_47700);
xnor UO_3172 (O_3172,N_45104,N_45849);
or UO_3173 (O_3173,N_49626,N_48674);
and UO_3174 (O_3174,N_45934,N_45629);
nor UO_3175 (O_3175,N_48297,N_47082);
xor UO_3176 (O_3176,N_49969,N_48011);
xnor UO_3177 (O_3177,N_46626,N_45353);
nand UO_3178 (O_3178,N_48996,N_49603);
nand UO_3179 (O_3179,N_48099,N_48015);
and UO_3180 (O_3180,N_48582,N_45437);
nand UO_3181 (O_3181,N_46159,N_48289);
and UO_3182 (O_3182,N_45755,N_49102);
xor UO_3183 (O_3183,N_48413,N_48105);
xor UO_3184 (O_3184,N_48518,N_48976);
or UO_3185 (O_3185,N_48168,N_45813);
nand UO_3186 (O_3186,N_47679,N_47275);
xor UO_3187 (O_3187,N_47746,N_45938);
xor UO_3188 (O_3188,N_48118,N_46366);
or UO_3189 (O_3189,N_49854,N_46084);
nor UO_3190 (O_3190,N_47573,N_47310);
xnor UO_3191 (O_3191,N_47068,N_46052);
or UO_3192 (O_3192,N_48940,N_49597);
xor UO_3193 (O_3193,N_45882,N_47795);
and UO_3194 (O_3194,N_45940,N_46633);
or UO_3195 (O_3195,N_45732,N_45635);
nand UO_3196 (O_3196,N_45991,N_47664);
xnor UO_3197 (O_3197,N_45106,N_45252);
nand UO_3198 (O_3198,N_47279,N_46123);
or UO_3199 (O_3199,N_45406,N_45794);
xnor UO_3200 (O_3200,N_49059,N_45766);
or UO_3201 (O_3201,N_45794,N_47552);
and UO_3202 (O_3202,N_49468,N_49102);
or UO_3203 (O_3203,N_47642,N_48816);
nand UO_3204 (O_3204,N_49099,N_48215);
nor UO_3205 (O_3205,N_45460,N_46681);
nand UO_3206 (O_3206,N_48082,N_49694);
and UO_3207 (O_3207,N_48691,N_49119);
nand UO_3208 (O_3208,N_46763,N_45124);
nand UO_3209 (O_3209,N_49664,N_45517);
or UO_3210 (O_3210,N_45875,N_45720);
xnor UO_3211 (O_3211,N_48639,N_47583);
or UO_3212 (O_3212,N_49942,N_47054);
or UO_3213 (O_3213,N_45928,N_46944);
or UO_3214 (O_3214,N_46237,N_46394);
nand UO_3215 (O_3215,N_49307,N_47774);
or UO_3216 (O_3216,N_47667,N_49095);
nand UO_3217 (O_3217,N_49812,N_49754);
or UO_3218 (O_3218,N_49146,N_47770);
xor UO_3219 (O_3219,N_45224,N_46296);
xor UO_3220 (O_3220,N_47023,N_48743);
xnor UO_3221 (O_3221,N_48886,N_49149);
or UO_3222 (O_3222,N_46666,N_49744);
and UO_3223 (O_3223,N_49829,N_45024);
or UO_3224 (O_3224,N_46039,N_46967);
xnor UO_3225 (O_3225,N_48964,N_46595);
nor UO_3226 (O_3226,N_46687,N_48231);
xnor UO_3227 (O_3227,N_48095,N_45119);
and UO_3228 (O_3228,N_47224,N_49173);
or UO_3229 (O_3229,N_47074,N_46812);
and UO_3230 (O_3230,N_45095,N_46890);
nor UO_3231 (O_3231,N_47461,N_49628);
or UO_3232 (O_3232,N_47628,N_46672);
or UO_3233 (O_3233,N_46966,N_45064);
nor UO_3234 (O_3234,N_46219,N_46939);
and UO_3235 (O_3235,N_49000,N_46077);
nor UO_3236 (O_3236,N_45661,N_48563);
nand UO_3237 (O_3237,N_46791,N_47653);
and UO_3238 (O_3238,N_46988,N_46504);
and UO_3239 (O_3239,N_45087,N_45990);
xor UO_3240 (O_3240,N_48446,N_49000);
or UO_3241 (O_3241,N_49093,N_45406);
and UO_3242 (O_3242,N_47999,N_47002);
xnor UO_3243 (O_3243,N_47711,N_47166);
nand UO_3244 (O_3244,N_45070,N_47787);
nand UO_3245 (O_3245,N_47677,N_48356);
and UO_3246 (O_3246,N_45203,N_48081);
or UO_3247 (O_3247,N_47802,N_46322);
nor UO_3248 (O_3248,N_47774,N_49439);
nor UO_3249 (O_3249,N_45301,N_48934);
nand UO_3250 (O_3250,N_49803,N_47901);
xor UO_3251 (O_3251,N_47905,N_46354);
nor UO_3252 (O_3252,N_47231,N_46325);
nand UO_3253 (O_3253,N_47787,N_49238);
and UO_3254 (O_3254,N_49318,N_47535);
nand UO_3255 (O_3255,N_49430,N_47870);
or UO_3256 (O_3256,N_45657,N_46898);
nand UO_3257 (O_3257,N_48782,N_49279);
nand UO_3258 (O_3258,N_45137,N_49640);
or UO_3259 (O_3259,N_45361,N_48303);
nand UO_3260 (O_3260,N_48736,N_45416);
and UO_3261 (O_3261,N_45142,N_47086);
or UO_3262 (O_3262,N_49084,N_45011);
xnor UO_3263 (O_3263,N_48309,N_48025);
nor UO_3264 (O_3264,N_48123,N_46326);
nor UO_3265 (O_3265,N_48180,N_45965);
and UO_3266 (O_3266,N_47766,N_49800);
or UO_3267 (O_3267,N_47052,N_47141);
nand UO_3268 (O_3268,N_47102,N_48140);
nand UO_3269 (O_3269,N_46322,N_48145);
nor UO_3270 (O_3270,N_48149,N_48150);
or UO_3271 (O_3271,N_48460,N_47098);
nand UO_3272 (O_3272,N_48123,N_45893);
nor UO_3273 (O_3273,N_45857,N_49365);
nand UO_3274 (O_3274,N_46906,N_45133);
nor UO_3275 (O_3275,N_48913,N_47215);
or UO_3276 (O_3276,N_47095,N_46325);
xnor UO_3277 (O_3277,N_48783,N_46466);
nor UO_3278 (O_3278,N_48349,N_47328);
xor UO_3279 (O_3279,N_48449,N_45173);
or UO_3280 (O_3280,N_45675,N_49862);
nor UO_3281 (O_3281,N_49129,N_48489);
and UO_3282 (O_3282,N_49373,N_47144);
xor UO_3283 (O_3283,N_49109,N_49784);
xor UO_3284 (O_3284,N_46087,N_48876);
nand UO_3285 (O_3285,N_46447,N_46241);
xor UO_3286 (O_3286,N_49149,N_48477);
nand UO_3287 (O_3287,N_48735,N_46921);
nor UO_3288 (O_3288,N_47210,N_47365);
nand UO_3289 (O_3289,N_48855,N_46472);
and UO_3290 (O_3290,N_48994,N_48885);
nor UO_3291 (O_3291,N_47133,N_46625);
nor UO_3292 (O_3292,N_48200,N_47930);
nand UO_3293 (O_3293,N_45747,N_47174);
and UO_3294 (O_3294,N_48918,N_47667);
or UO_3295 (O_3295,N_45030,N_47291);
xnor UO_3296 (O_3296,N_47208,N_45898);
and UO_3297 (O_3297,N_47126,N_48527);
nand UO_3298 (O_3298,N_47665,N_48045);
nor UO_3299 (O_3299,N_47626,N_48888);
or UO_3300 (O_3300,N_45947,N_45348);
nor UO_3301 (O_3301,N_49554,N_49062);
nor UO_3302 (O_3302,N_49004,N_48506);
xor UO_3303 (O_3303,N_46711,N_47458);
xor UO_3304 (O_3304,N_47384,N_45473);
or UO_3305 (O_3305,N_47451,N_46155);
xnor UO_3306 (O_3306,N_45266,N_47474);
nand UO_3307 (O_3307,N_47890,N_48717);
nand UO_3308 (O_3308,N_49774,N_45099);
xnor UO_3309 (O_3309,N_49812,N_46363);
and UO_3310 (O_3310,N_47993,N_47331);
and UO_3311 (O_3311,N_48487,N_49022);
or UO_3312 (O_3312,N_49593,N_45779);
xor UO_3313 (O_3313,N_49258,N_48769);
and UO_3314 (O_3314,N_48749,N_47972);
and UO_3315 (O_3315,N_48898,N_46104);
nor UO_3316 (O_3316,N_45871,N_45421);
nand UO_3317 (O_3317,N_47180,N_45703);
nand UO_3318 (O_3318,N_47343,N_46244);
or UO_3319 (O_3319,N_49809,N_46637);
and UO_3320 (O_3320,N_45507,N_49066);
xor UO_3321 (O_3321,N_46272,N_45085);
nand UO_3322 (O_3322,N_45040,N_46558);
nand UO_3323 (O_3323,N_49944,N_47689);
nor UO_3324 (O_3324,N_48433,N_45916);
nor UO_3325 (O_3325,N_45374,N_46222);
xor UO_3326 (O_3326,N_49614,N_47889);
or UO_3327 (O_3327,N_49578,N_49491);
and UO_3328 (O_3328,N_45949,N_46630);
nand UO_3329 (O_3329,N_46359,N_48287);
and UO_3330 (O_3330,N_46479,N_48948);
and UO_3331 (O_3331,N_46769,N_49734);
xnor UO_3332 (O_3332,N_47613,N_46979);
nor UO_3333 (O_3333,N_46665,N_46420);
xnor UO_3334 (O_3334,N_49447,N_47073);
and UO_3335 (O_3335,N_49791,N_48834);
or UO_3336 (O_3336,N_46729,N_49844);
xor UO_3337 (O_3337,N_45994,N_45462);
nand UO_3338 (O_3338,N_49089,N_46987);
xor UO_3339 (O_3339,N_47914,N_48928);
and UO_3340 (O_3340,N_47774,N_45288);
nor UO_3341 (O_3341,N_48788,N_46502);
or UO_3342 (O_3342,N_49775,N_48916);
or UO_3343 (O_3343,N_46524,N_49460);
and UO_3344 (O_3344,N_45473,N_49826);
or UO_3345 (O_3345,N_48608,N_47070);
and UO_3346 (O_3346,N_48792,N_46097);
xnor UO_3347 (O_3347,N_48911,N_45341);
or UO_3348 (O_3348,N_46907,N_45783);
and UO_3349 (O_3349,N_48120,N_47685);
and UO_3350 (O_3350,N_45184,N_47581);
xor UO_3351 (O_3351,N_47747,N_49881);
nand UO_3352 (O_3352,N_45496,N_45617);
or UO_3353 (O_3353,N_46476,N_49842);
nand UO_3354 (O_3354,N_46148,N_47521);
nand UO_3355 (O_3355,N_49933,N_48639);
nand UO_3356 (O_3356,N_45176,N_48377);
and UO_3357 (O_3357,N_45823,N_48184);
and UO_3358 (O_3358,N_45342,N_48477);
and UO_3359 (O_3359,N_45062,N_46484);
and UO_3360 (O_3360,N_47349,N_45480);
nor UO_3361 (O_3361,N_48618,N_48819);
xor UO_3362 (O_3362,N_48579,N_48104);
or UO_3363 (O_3363,N_47681,N_46952);
xnor UO_3364 (O_3364,N_48644,N_46827);
and UO_3365 (O_3365,N_48281,N_46375);
and UO_3366 (O_3366,N_45867,N_49554);
nand UO_3367 (O_3367,N_49093,N_46851);
and UO_3368 (O_3368,N_46668,N_49939);
and UO_3369 (O_3369,N_45648,N_49184);
nor UO_3370 (O_3370,N_48150,N_47207);
xor UO_3371 (O_3371,N_45514,N_46449);
nor UO_3372 (O_3372,N_48058,N_45933);
or UO_3373 (O_3373,N_46292,N_47727);
nor UO_3374 (O_3374,N_45080,N_49261);
nor UO_3375 (O_3375,N_46091,N_48004);
and UO_3376 (O_3376,N_46856,N_46393);
or UO_3377 (O_3377,N_47152,N_46522);
or UO_3378 (O_3378,N_46311,N_45681);
nor UO_3379 (O_3379,N_45552,N_45221);
nand UO_3380 (O_3380,N_49832,N_45453);
or UO_3381 (O_3381,N_48857,N_46913);
nor UO_3382 (O_3382,N_48641,N_46982);
xor UO_3383 (O_3383,N_46318,N_45548);
and UO_3384 (O_3384,N_49672,N_46040);
nand UO_3385 (O_3385,N_47785,N_45048);
and UO_3386 (O_3386,N_49882,N_49272);
nand UO_3387 (O_3387,N_46373,N_48359);
and UO_3388 (O_3388,N_47123,N_47522);
or UO_3389 (O_3389,N_49021,N_49675);
xor UO_3390 (O_3390,N_47926,N_46326);
xor UO_3391 (O_3391,N_48542,N_47452);
xnor UO_3392 (O_3392,N_47409,N_45838);
nor UO_3393 (O_3393,N_46371,N_45880);
nand UO_3394 (O_3394,N_49966,N_45674);
and UO_3395 (O_3395,N_46973,N_48063);
and UO_3396 (O_3396,N_48377,N_46340);
and UO_3397 (O_3397,N_48071,N_49462);
and UO_3398 (O_3398,N_45432,N_45820);
xnor UO_3399 (O_3399,N_48111,N_48897);
nand UO_3400 (O_3400,N_47617,N_46527);
nor UO_3401 (O_3401,N_47738,N_47487);
or UO_3402 (O_3402,N_48742,N_48095);
or UO_3403 (O_3403,N_47591,N_45758);
and UO_3404 (O_3404,N_45757,N_47857);
nor UO_3405 (O_3405,N_46619,N_47189);
nor UO_3406 (O_3406,N_49457,N_45494);
xor UO_3407 (O_3407,N_48005,N_45063);
nand UO_3408 (O_3408,N_47886,N_49557);
nor UO_3409 (O_3409,N_48307,N_48605);
nor UO_3410 (O_3410,N_49646,N_48484);
xnor UO_3411 (O_3411,N_45582,N_45545);
nand UO_3412 (O_3412,N_46483,N_48523);
or UO_3413 (O_3413,N_49062,N_47732);
xnor UO_3414 (O_3414,N_47252,N_46488);
nand UO_3415 (O_3415,N_48119,N_49050);
nor UO_3416 (O_3416,N_47067,N_47003);
and UO_3417 (O_3417,N_48933,N_45549);
and UO_3418 (O_3418,N_45707,N_46626);
nor UO_3419 (O_3419,N_46126,N_46781);
nor UO_3420 (O_3420,N_48469,N_47831);
and UO_3421 (O_3421,N_45597,N_45657);
nand UO_3422 (O_3422,N_46810,N_47202);
nor UO_3423 (O_3423,N_46225,N_48088);
nor UO_3424 (O_3424,N_45285,N_47831);
or UO_3425 (O_3425,N_49475,N_47887);
nand UO_3426 (O_3426,N_46925,N_48277);
xnor UO_3427 (O_3427,N_47293,N_47259);
nand UO_3428 (O_3428,N_46810,N_48061);
nand UO_3429 (O_3429,N_46817,N_48294);
or UO_3430 (O_3430,N_48721,N_49335);
xnor UO_3431 (O_3431,N_49383,N_49246);
xnor UO_3432 (O_3432,N_48855,N_48048);
or UO_3433 (O_3433,N_46811,N_48642);
and UO_3434 (O_3434,N_48889,N_47406);
xnor UO_3435 (O_3435,N_47835,N_45897);
nand UO_3436 (O_3436,N_46532,N_46443);
nor UO_3437 (O_3437,N_47187,N_46846);
nor UO_3438 (O_3438,N_45301,N_48631);
xnor UO_3439 (O_3439,N_49561,N_49114);
and UO_3440 (O_3440,N_45027,N_48149);
nand UO_3441 (O_3441,N_45097,N_45742);
nand UO_3442 (O_3442,N_45525,N_46690);
nor UO_3443 (O_3443,N_48689,N_48339);
and UO_3444 (O_3444,N_48666,N_48543);
xnor UO_3445 (O_3445,N_46116,N_49404);
xnor UO_3446 (O_3446,N_48891,N_48913);
nand UO_3447 (O_3447,N_46776,N_49383);
and UO_3448 (O_3448,N_46592,N_46051);
xnor UO_3449 (O_3449,N_45366,N_49701);
or UO_3450 (O_3450,N_46683,N_48871);
or UO_3451 (O_3451,N_49894,N_45824);
and UO_3452 (O_3452,N_45140,N_48546);
nor UO_3453 (O_3453,N_49054,N_48894);
nand UO_3454 (O_3454,N_46594,N_46005);
nand UO_3455 (O_3455,N_48059,N_47030);
or UO_3456 (O_3456,N_46630,N_47327);
nand UO_3457 (O_3457,N_49131,N_49796);
nand UO_3458 (O_3458,N_48586,N_49607);
xor UO_3459 (O_3459,N_46275,N_48324);
and UO_3460 (O_3460,N_49855,N_46877);
xor UO_3461 (O_3461,N_48030,N_46660);
nor UO_3462 (O_3462,N_46824,N_49570);
or UO_3463 (O_3463,N_48319,N_48150);
nand UO_3464 (O_3464,N_48334,N_47513);
nor UO_3465 (O_3465,N_49246,N_45141);
and UO_3466 (O_3466,N_45053,N_47823);
xnor UO_3467 (O_3467,N_49959,N_49795);
xor UO_3468 (O_3468,N_46021,N_47631);
nor UO_3469 (O_3469,N_45263,N_46321);
xor UO_3470 (O_3470,N_48449,N_47472);
nor UO_3471 (O_3471,N_45032,N_46045);
and UO_3472 (O_3472,N_45508,N_49239);
nor UO_3473 (O_3473,N_47552,N_45807);
xnor UO_3474 (O_3474,N_45374,N_46282);
xor UO_3475 (O_3475,N_49706,N_48506);
and UO_3476 (O_3476,N_49249,N_45564);
and UO_3477 (O_3477,N_45551,N_47576);
xor UO_3478 (O_3478,N_45072,N_49535);
or UO_3479 (O_3479,N_45150,N_49887);
or UO_3480 (O_3480,N_48561,N_45867);
nor UO_3481 (O_3481,N_46156,N_46612);
nor UO_3482 (O_3482,N_49164,N_49919);
nand UO_3483 (O_3483,N_46820,N_49598);
xnor UO_3484 (O_3484,N_49806,N_47936);
or UO_3485 (O_3485,N_48183,N_47702);
and UO_3486 (O_3486,N_46040,N_48752);
or UO_3487 (O_3487,N_45434,N_48704);
xor UO_3488 (O_3488,N_45809,N_48666);
nand UO_3489 (O_3489,N_47486,N_45273);
nand UO_3490 (O_3490,N_46642,N_48414);
xnor UO_3491 (O_3491,N_47691,N_49093);
and UO_3492 (O_3492,N_46029,N_45574);
xnor UO_3493 (O_3493,N_45371,N_45867);
nor UO_3494 (O_3494,N_49639,N_49147);
nor UO_3495 (O_3495,N_45476,N_48418);
nand UO_3496 (O_3496,N_45161,N_46431);
and UO_3497 (O_3497,N_46135,N_48145);
and UO_3498 (O_3498,N_47083,N_49540);
or UO_3499 (O_3499,N_49250,N_49372);
nand UO_3500 (O_3500,N_45654,N_45537);
xor UO_3501 (O_3501,N_49288,N_47538);
and UO_3502 (O_3502,N_46583,N_46657);
and UO_3503 (O_3503,N_46070,N_46646);
nor UO_3504 (O_3504,N_49423,N_46161);
nor UO_3505 (O_3505,N_49847,N_45920);
nand UO_3506 (O_3506,N_47283,N_48857);
nand UO_3507 (O_3507,N_47677,N_49949);
xnor UO_3508 (O_3508,N_45595,N_45566);
and UO_3509 (O_3509,N_45734,N_47034);
nand UO_3510 (O_3510,N_48390,N_47637);
nor UO_3511 (O_3511,N_45069,N_45453);
nand UO_3512 (O_3512,N_47166,N_47098);
xor UO_3513 (O_3513,N_46759,N_49842);
nor UO_3514 (O_3514,N_49965,N_45934);
nor UO_3515 (O_3515,N_47990,N_47004);
and UO_3516 (O_3516,N_49096,N_45261);
nor UO_3517 (O_3517,N_48741,N_45288);
or UO_3518 (O_3518,N_46222,N_48058);
and UO_3519 (O_3519,N_45618,N_45708);
nand UO_3520 (O_3520,N_49947,N_46865);
nand UO_3521 (O_3521,N_46590,N_45542);
and UO_3522 (O_3522,N_46933,N_46738);
nor UO_3523 (O_3523,N_45029,N_45648);
nand UO_3524 (O_3524,N_49150,N_49806);
nand UO_3525 (O_3525,N_48900,N_48198);
nor UO_3526 (O_3526,N_48595,N_47019);
nand UO_3527 (O_3527,N_45765,N_49667);
xnor UO_3528 (O_3528,N_49249,N_45868);
and UO_3529 (O_3529,N_49800,N_47632);
nand UO_3530 (O_3530,N_49718,N_48920);
nand UO_3531 (O_3531,N_46742,N_48408);
xnor UO_3532 (O_3532,N_49129,N_47250);
nor UO_3533 (O_3533,N_46739,N_48968);
xor UO_3534 (O_3534,N_48163,N_49492);
or UO_3535 (O_3535,N_47191,N_48187);
nor UO_3536 (O_3536,N_46539,N_48571);
or UO_3537 (O_3537,N_48811,N_49885);
xnor UO_3538 (O_3538,N_45577,N_46873);
xor UO_3539 (O_3539,N_48834,N_46004);
nand UO_3540 (O_3540,N_48465,N_47739);
nand UO_3541 (O_3541,N_47939,N_48631);
and UO_3542 (O_3542,N_49828,N_48753);
or UO_3543 (O_3543,N_47390,N_47285);
nand UO_3544 (O_3544,N_48962,N_46652);
xnor UO_3545 (O_3545,N_47722,N_49380);
nand UO_3546 (O_3546,N_47681,N_49977);
or UO_3547 (O_3547,N_49356,N_45595);
xor UO_3548 (O_3548,N_46690,N_45148);
nor UO_3549 (O_3549,N_46941,N_49559);
nand UO_3550 (O_3550,N_48989,N_45793);
xor UO_3551 (O_3551,N_46326,N_47847);
xor UO_3552 (O_3552,N_48757,N_48050);
nand UO_3553 (O_3553,N_47286,N_45167);
or UO_3554 (O_3554,N_49156,N_47557);
nand UO_3555 (O_3555,N_45450,N_48771);
or UO_3556 (O_3556,N_48252,N_46584);
nor UO_3557 (O_3557,N_45996,N_45384);
and UO_3558 (O_3558,N_46613,N_46012);
or UO_3559 (O_3559,N_47987,N_49595);
nor UO_3560 (O_3560,N_48217,N_48215);
nand UO_3561 (O_3561,N_49276,N_45437);
nor UO_3562 (O_3562,N_47640,N_47797);
xor UO_3563 (O_3563,N_46701,N_49362);
xor UO_3564 (O_3564,N_47628,N_47474);
nor UO_3565 (O_3565,N_45638,N_48527);
nor UO_3566 (O_3566,N_45908,N_47919);
nand UO_3567 (O_3567,N_47248,N_49907);
or UO_3568 (O_3568,N_48260,N_47829);
and UO_3569 (O_3569,N_45892,N_49578);
nand UO_3570 (O_3570,N_47710,N_46322);
xor UO_3571 (O_3571,N_48834,N_45005);
or UO_3572 (O_3572,N_47265,N_45477);
nor UO_3573 (O_3573,N_47849,N_48902);
xor UO_3574 (O_3574,N_45575,N_48893);
nor UO_3575 (O_3575,N_47164,N_46757);
nor UO_3576 (O_3576,N_45478,N_47949);
and UO_3577 (O_3577,N_47374,N_46628);
nor UO_3578 (O_3578,N_48731,N_45491);
or UO_3579 (O_3579,N_46911,N_46235);
and UO_3580 (O_3580,N_47630,N_48525);
or UO_3581 (O_3581,N_45636,N_46461);
or UO_3582 (O_3582,N_45640,N_45526);
nand UO_3583 (O_3583,N_48475,N_47632);
and UO_3584 (O_3584,N_45245,N_49103);
and UO_3585 (O_3585,N_47871,N_48754);
and UO_3586 (O_3586,N_47979,N_46294);
or UO_3587 (O_3587,N_45425,N_46622);
and UO_3588 (O_3588,N_46089,N_48619);
nor UO_3589 (O_3589,N_48743,N_49289);
nor UO_3590 (O_3590,N_45305,N_48047);
and UO_3591 (O_3591,N_46977,N_46793);
xnor UO_3592 (O_3592,N_45123,N_49567);
xor UO_3593 (O_3593,N_48443,N_49472);
nand UO_3594 (O_3594,N_48105,N_46015);
nand UO_3595 (O_3595,N_47486,N_47351);
xnor UO_3596 (O_3596,N_47985,N_48471);
and UO_3597 (O_3597,N_48402,N_46715);
xor UO_3598 (O_3598,N_45592,N_46989);
or UO_3599 (O_3599,N_46178,N_48899);
xor UO_3600 (O_3600,N_47065,N_45380);
nand UO_3601 (O_3601,N_47590,N_49893);
and UO_3602 (O_3602,N_47324,N_46210);
nand UO_3603 (O_3603,N_46740,N_49419);
nand UO_3604 (O_3604,N_45130,N_49570);
xor UO_3605 (O_3605,N_45792,N_47066);
or UO_3606 (O_3606,N_47209,N_48874);
nand UO_3607 (O_3607,N_46234,N_47649);
nand UO_3608 (O_3608,N_49788,N_45729);
xor UO_3609 (O_3609,N_48885,N_46870);
xor UO_3610 (O_3610,N_46348,N_45890);
xor UO_3611 (O_3611,N_45964,N_49650);
xnor UO_3612 (O_3612,N_49672,N_46468);
nor UO_3613 (O_3613,N_48678,N_45589);
nand UO_3614 (O_3614,N_45366,N_47998);
nand UO_3615 (O_3615,N_47919,N_46193);
and UO_3616 (O_3616,N_45201,N_48644);
xnor UO_3617 (O_3617,N_47513,N_48065);
xnor UO_3618 (O_3618,N_49604,N_45707);
and UO_3619 (O_3619,N_48465,N_48662);
nand UO_3620 (O_3620,N_49400,N_48090);
and UO_3621 (O_3621,N_49317,N_49907);
or UO_3622 (O_3622,N_47722,N_45917);
and UO_3623 (O_3623,N_47917,N_46520);
nand UO_3624 (O_3624,N_47605,N_49986);
xor UO_3625 (O_3625,N_46959,N_48722);
nand UO_3626 (O_3626,N_45988,N_46135);
xor UO_3627 (O_3627,N_47906,N_45176);
nor UO_3628 (O_3628,N_46629,N_49421);
nor UO_3629 (O_3629,N_47222,N_48647);
and UO_3630 (O_3630,N_47480,N_46588);
nor UO_3631 (O_3631,N_45262,N_45489);
xor UO_3632 (O_3632,N_48038,N_46686);
nor UO_3633 (O_3633,N_45674,N_47690);
or UO_3634 (O_3634,N_45768,N_45549);
nand UO_3635 (O_3635,N_45974,N_49960);
nor UO_3636 (O_3636,N_46241,N_45624);
nor UO_3637 (O_3637,N_46103,N_45224);
nand UO_3638 (O_3638,N_48743,N_45802);
nor UO_3639 (O_3639,N_45114,N_46895);
nor UO_3640 (O_3640,N_46681,N_45843);
nor UO_3641 (O_3641,N_46684,N_48435);
and UO_3642 (O_3642,N_45991,N_48566);
xnor UO_3643 (O_3643,N_46204,N_47430);
xor UO_3644 (O_3644,N_48316,N_46192);
xor UO_3645 (O_3645,N_48426,N_46651);
nor UO_3646 (O_3646,N_46466,N_47820);
nand UO_3647 (O_3647,N_46856,N_48522);
nor UO_3648 (O_3648,N_45507,N_49815);
nand UO_3649 (O_3649,N_49909,N_45954);
and UO_3650 (O_3650,N_46124,N_48137);
nor UO_3651 (O_3651,N_49862,N_48878);
nand UO_3652 (O_3652,N_48746,N_49615);
xor UO_3653 (O_3653,N_45429,N_48957);
nor UO_3654 (O_3654,N_47873,N_46916);
and UO_3655 (O_3655,N_48983,N_49376);
xnor UO_3656 (O_3656,N_46211,N_49982);
and UO_3657 (O_3657,N_47715,N_49777);
xor UO_3658 (O_3658,N_46890,N_48774);
xor UO_3659 (O_3659,N_49371,N_45812);
nand UO_3660 (O_3660,N_47351,N_48286);
nor UO_3661 (O_3661,N_49185,N_47670);
xnor UO_3662 (O_3662,N_49452,N_48474);
nor UO_3663 (O_3663,N_46398,N_45455);
nor UO_3664 (O_3664,N_47444,N_49421);
and UO_3665 (O_3665,N_48478,N_46827);
nand UO_3666 (O_3666,N_48966,N_45013);
and UO_3667 (O_3667,N_49944,N_46769);
nand UO_3668 (O_3668,N_47192,N_48744);
nand UO_3669 (O_3669,N_45628,N_46075);
nor UO_3670 (O_3670,N_45022,N_46709);
nand UO_3671 (O_3671,N_46671,N_46768);
or UO_3672 (O_3672,N_45048,N_46772);
nor UO_3673 (O_3673,N_47577,N_46188);
and UO_3674 (O_3674,N_47955,N_48099);
nand UO_3675 (O_3675,N_47296,N_45875);
nand UO_3676 (O_3676,N_45462,N_46552);
or UO_3677 (O_3677,N_49166,N_47157);
and UO_3678 (O_3678,N_45574,N_46026);
and UO_3679 (O_3679,N_48125,N_45603);
nand UO_3680 (O_3680,N_49955,N_48137);
xnor UO_3681 (O_3681,N_49283,N_49594);
nor UO_3682 (O_3682,N_45196,N_46110);
nor UO_3683 (O_3683,N_46819,N_49055);
nand UO_3684 (O_3684,N_45196,N_45104);
xnor UO_3685 (O_3685,N_48361,N_49643);
nor UO_3686 (O_3686,N_49498,N_47464);
and UO_3687 (O_3687,N_48921,N_46340);
or UO_3688 (O_3688,N_48826,N_48212);
or UO_3689 (O_3689,N_48119,N_47302);
xnor UO_3690 (O_3690,N_45846,N_48041);
nand UO_3691 (O_3691,N_45869,N_46933);
or UO_3692 (O_3692,N_45068,N_46692);
xnor UO_3693 (O_3693,N_49776,N_45416);
nor UO_3694 (O_3694,N_45463,N_47841);
nor UO_3695 (O_3695,N_46880,N_48551);
xor UO_3696 (O_3696,N_47999,N_48898);
xnor UO_3697 (O_3697,N_49569,N_46155);
nor UO_3698 (O_3698,N_49091,N_46500);
nand UO_3699 (O_3699,N_45320,N_49633);
and UO_3700 (O_3700,N_48257,N_46759);
or UO_3701 (O_3701,N_48109,N_48062);
or UO_3702 (O_3702,N_46961,N_45895);
and UO_3703 (O_3703,N_46526,N_46100);
xnor UO_3704 (O_3704,N_45902,N_48120);
nor UO_3705 (O_3705,N_49970,N_47932);
or UO_3706 (O_3706,N_49186,N_48033);
or UO_3707 (O_3707,N_45620,N_47508);
or UO_3708 (O_3708,N_46748,N_46113);
nor UO_3709 (O_3709,N_47364,N_48314);
or UO_3710 (O_3710,N_46367,N_48796);
nand UO_3711 (O_3711,N_47668,N_48048);
xor UO_3712 (O_3712,N_46459,N_46786);
xor UO_3713 (O_3713,N_46143,N_49762);
xnor UO_3714 (O_3714,N_49770,N_49515);
or UO_3715 (O_3715,N_48491,N_45758);
xor UO_3716 (O_3716,N_45870,N_48977);
nand UO_3717 (O_3717,N_48283,N_45593);
nand UO_3718 (O_3718,N_49604,N_47894);
or UO_3719 (O_3719,N_45806,N_46444);
nand UO_3720 (O_3720,N_49210,N_48992);
nand UO_3721 (O_3721,N_47427,N_45089);
xor UO_3722 (O_3722,N_49377,N_45799);
nand UO_3723 (O_3723,N_47850,N_46801);
and UO_3724 (O_3724,N_46933,N_45967);
xor UO_3725 (O_3725,N_49830,N_45579);
nor UO_3726 (O_3726,N_46473,N_49340);
nor UO_3727 (O_3727,N_46526,N_49218);
or UO_3728 (O_3728,N_48600,N_49221);
and UO_3729 (O_3729,N_46473,N_49459);
and UO_3730 (O_3730,N_47145,N_48484);
and UO_3731 (O_3731,N_47239,N_49916);
and UO_3732 (O_3732,N_45271,N_49322);
nor UO_3733 (O_3733,N_46270,N_45280);
and UO_3734 (O_3734,N_46268,N_46463);
nand UO_3735 (O_3735,N_49571,N_49425);
nand UO_3736 (O_3736,N_47660,N_49271);
or UO_3737 (O_3737,N_46672,N_48096);
nand UO_3738 (O_3738,N_48087,N_49888);
and UO_3739 (O_3739,N_45869,N_48140);
nand UO_3740 (O_3740,N_45158,N_49729);
xor UO_3741 (O_3741,N_47657,N_45708);
and UO_3742 (O_3742,N_45244,N_45283);
or UO_3743 (O_3743,N_47122,N_48480);
nand UO_3744 (O_3744,N_48580,N_49508);
nand UO_3745 (O_3745,N_48067,N_48392);
or UO_3746 (O_3746,N_47409,N_48240);
xnor UO_3747 (O_3747,N_46702,N_46078);
and UO_3748 (O_3748,N_49896,N_46888);
xnor UO_3749 (O_3749,N_47738,N_47512);
and UO_3750 (O_3750,N_49585,N_49438);
xor UO_3751 (O_3751,N_45204,N_49582);
and UO_3752 (O_3752,N_48911,N_45561);
or UO_3753 (O_3753,N_49758,N_49735);
nand UO_3754 (O_3754,N_48459,N_47125);
and UO_3755 (O_3755,N_45398,N_45914);
or UO_3756 (O_3756,N_49637,N_46882);
xor UO_3757 (O_3757,N_49133,N_49401);
xnor UO_3758 (O_3758,N_48875,N_47560);
nand UO_3759 (O_3759,N_48213,N_49094);
nand UO_3760 (O_3760,N_49801,N_45731);
or UO_3761 (O_3761,N_49576,N_45524);
xnor UO_3762 (O_3762,N_49116,N_49358);
and UO_3763 (O_3763,N_45319,N_48409);
or UO_3764 (O_3764,N_46293,N_48089);
and UO_3765 (O_3765,N_45578,N_45198);
xor UO_3766 (O_3766,N_48567,N_48169);
nor UO_3767 (O_3767,N_45551,N_47301);
or UO_3768 (O_3768,N_48522,N_49625);
and UO_3769 (O_3769,N_47886,N_49790);
or UO_3770 (O_3770,N_48587,N_45336);
nor UO_3771 (O_3771,N_46728,N_45077);
nor UO_3772 (O_3772,N_49959,N_45356);
and UO_3773 (O_3773,N_48804,N_45727);
xor UO_3774 (O_3774,N_45582,N_45429);
xnor UO_3775 (O_3775,N_47926,N_49475);
nor UO_3776 (O_3776,N_48513,N_47294);
and UO_3777 (O_3777,N_47288,N_48059);
nor UO_3778 (O_3778,N_48640,N_48882);
and UO_3779 (O_3779,N_47857,N_45038);
xor UO_3780 (O_3780,N_48843,N_46618);
or UO_3781 (O_3781,N_46950,N_46765);
nand UO_3782 (O_3782,N_47514,N_49567);
xor UO_3783 (O_3783,N_49498,N_45834);
nand UO_3784 (O_3784,N_48957,N_47149);
nor UO_3785 (O_3785,N_48717,N_48554);
and UO_3786 (O_3786,N_48311,N_48331);
xor UO_3787 (O_3787,N_48960,N_46693);
or UO_3788 (O_3788,N_48749,N_47572);
nand UO_3789 (O_3789,N_45511,N_49419);
or UO_3790 (O_3790,N_47030,N_45672);
nor UO_3791 (O_3791,N_47829,N_45762);
nand UO_3792 (O_3792,N_49117,N_47008);
nor UO_3793 (O_3793,N_48139,N_46168);
or UO_3794 (O_3794,N_47285,N_45274);
or UO_3795 (O_3795,N_45166,N_47230);
nand UO_3796 (O_3796,N_49705,N_48305);
xnor UO_3797 (O_3797,N_46167,N_49654);
and UO_3798 (O_3798,N_46121,N_47217);
and UO_3799 (O_3799,N_48168,N_49525);
or UO_3800 (O_3800,N_49114,N_47155);
nand UO_3801 (O_3801,N_47888,N_48822);
xnor UO_3802 (O_3802,N_46134,N_47334);
and UO_3803 (O_3803,N_48348,N_48381);
and UO_3804 (O_3804,N_47847,N_46851);
nand UO_3805 (O_3805,N_45453,N_46261);
or UO_3806 (O_3806,N_49059,N_45063);
nand UO_3807 (O_3807,N_48916,N_45511);
xor UO_3808 (O_3808,N_47080,N_48781);
nor UO_3809 (O_3809,N_46854,N_48961);
or UO_3810 (O_3810,N_45127,N_48720);
nand UO_3811 (O_3811,N_49486,N_49310);
or UO_3812 (O_3812,N_46945,N_49267);
or UO_3813 (O_3813,N_45691,N_46830);
and UO_3814 (O_3814,N_49096,N_48367);
xor UO_3815 (O_3815,N_49608,N_47552);
and UO_3816 (O_3816,N_49730,N_48703);
or UO_3817 (O_3817,N_49125,N_49406);
nor UO_3818 (O_3818,N_47855,N_48862);
nor UO_3819 (O_3819,N_46984,N_49668);
xor UO_3820 (O_3820,N_45019,N_47871);
or UO_3821 (O_3821,N_49109,N_45240);
or UO_3822 (O_3822,N_47715,N_49916);
xnor UO_3823 (O_3823,N_48963,N_46164);
xnor UO_3824 (O_3824,N_46131,N_48437);
nor UO_3825 (O_3825,N_48728,N_47366);
and UO_3826 (O_3826,N_46133,N_46908);
and UO_3827 (O_3827,N_45130,N_49897);
or UO_3828 (O_3828,N_48241,N_48207);
nand UO_3829 (O_3829,N_47941,N_46637);
or UO_3830 (O_3830,N_45345,N_49176);
xnor UO_3831 (O_3831,N_45844,N_48910);
or UO_3832 (O_3832,N_47790,N_47237);
and UO_3833 (O_3833,N_47918,N_46873);
nand UO_3834 (O_3834,N_49612,N_47272);
nand UO_3835 (O_3835,N_48577,N_47215);
nand UO_3836 (O_3836,N_45270,N_45992);
xnor UO_3837 (O_3837,N_47738,N_49852);
nor UO_3838 (O_3838,N_47393,N_49315);
nand UO_3839 (O_3839,N_49596,N_47714);
nand UO_3840 (O_3840,N_46998,N_48205);
and UO_3841 (O_3841,N_49976,N_49263);
and UO_3842 (O_3842,N_49489,N_48899);
nor UO_3843 (O_3843,N_48530,N_46212);
and UO_3844 (O_3844,N_49534,N_46662);
nor UO_3845 (O_3845,N_47622,N_48688);
xor UO_3846 (O_3846,N_48465,N_45763);
nand UO_3847 (O_3847,N_45430,N_48815);
or UO_3848 (O_3848,N_49867,N_47117);
nand UO_3849 (O_3849,N_48021,N_45967);
nand UO_3850 (O_3850,N_45689,N_47255);
and UO_3851 (O_3851,N_46646,N_49147);
and UO_3852 (O_3852,N_48434,N_48485);
and UO_3853 (O_3853,N_45667,N_46479);
nand UO_3854 (O_3854,N_49899,N_46853);
nor UO_3855 (O_3855,N_47026,N_46914);
or UO_3856 (O_3856,N_45518,N_48993);
xnor UO_3857 (O_3857,N_48921,N_48435);
and UO_3858 (O_3858,N_49369,N_48469);
or UO_3859 (O_3859,N_49835,N_45592);
nor UO_3860 (O_3860,N_48889,N_45471);
and UO_3861 (O_3861,N_48130,N_47076);
nand UO_3862 (O_3862,N_45401,N_49300);
nor UO_3863 (O_3863,N_48481,N_46209);
and UO_3864 (O_3864,N_46147,N_45729);
nand UO_3865 (O_3865,N_46591,N_48221);
or UO_3866 (O_3866,N_48031,N_45965);
and UO_3867 (O_3867,N_48599,N_45210);
or UO_3868 (O_3868,N_49314,N_46993);
or UO_3869 (O_3869,N_46849,N_47486);
and UO_3870 (O_3870,N_49525,N_45657);
nand UO_3871 (O_3871,N_49730,N_46967);
xnor UO_3872 (O_3872,N_48283,N_48006);
xor UO_3873 (O_3873,N_48704,N_46226);
and UO_3874 (O_3874,N_49069,N_48937);
nor UO_3875 (O_3875,N_46408,N_45623);
xnor UO_3876 (O_3876,N_47024,N_46062);
nor UO_3877 (O_3877,N_49023,N_45418);
nor UO_3878 (O_3878,N_46805,N_46643);
or UO_3879 (O_3879,N_45921,N_47706);
or UO_3880 (O_3880,N_47539,N_47562);
nor UO_3881 (O_3881,N_46084,N_47580);
or UO_3882 (O_3882,N_49931,N_45384);
and UO_3883 (O_3883,N_46534,N_46609);
or UO_3884 (O_3884,N_47838,N_49325);
or UO_3885 (O_3885,N_48352,N_47506);
nor UO_3886 (O_3886,N_49529,N_48286);
nor UO_3887 (O_3887,N_47356,N_49300);
nand UO_3888 (O_3888,N_45850,N_45563);
and UO_3889 (O_3889,N_48562,N_49954);
and UO_3890 (O_3890,N_46344,N_47249);
nand UO_3891 (O_3891,N_45824,N_47954);
xnor UO_3892 (O_3892,N_49997,N_45687);
nand UO_3893 (O_3893,N_48746,N_47481);
or UO_3894 (O_3894,N_46162,N_49321);
xor UO_3895 (O_3895,N_45350,N_48810);
xnor UO_3896 (O_3896,N_48959,N_47058);
and UO_3897 (O_3897,N_45071,N_48127);
nor UO_3898 (O_3898,N_48760,N_46224);
or UO_3899 (O_3899,N_49396,N_47682);
nand UO_3900 (O_3900,N_49605,N_45199);
nand UO_3901 (O_3901,N_48583,N_49463);
or UO_3902 (O_3902,N_45641,N_48056);
nand UO_3903 (O_3903,N_46763,N_45732);
xor UO_3904 (O_3904,N_47845,N_45032);
and UO_3905 (O_3905,N_45072,N_47607);
or UO_3906 (O_3906,N_48914,N_49146);
xnor UO_3907 (O_3907,N_48534,N_45056);
or UO_3908 (O_3908,N_47156,N_49965);
nand UO_3909 (O_3909,N_45712,N_46875);
nor UO_3910 (O_3910,N_45537,N_48392);
or UO_3911 (O_3911,N_46726,N_45306);
xnor UO_3912 (O_3912,N_45686,N_45532);
or UO_3913 (O_3913,N_47608,N_48481);
xnor UO_3914 (O_3914,N_47719,N_46549);
xor UO_3915 (O_3915,N_46414,N_47499);
xnor UO_3916 (O_3916,N_49460,N_48231);
xnor UO_3917 (O_3917,N_45945,N_49129);
or UO_3918 (O_3918,N_46278,N_45165);
xnor UO_3919 (O_3919,N_49634,N_49544);
or UO_3920 (O_3920,N_47425,N_49067);
nor UO_3921 (O_3921,N_46145,N_47342);
xor UO_3922 (O_3922,N_49145,N_49457);
nor UO_3923 (O_3923,N_49856,N_48379);
or UO_3924 (O_3924,N_48109,N_49697);
and UO_3925 (O_3925,N_45354,N_49449);
nor UO_3926 (O_3926,N_46399,N_46665);
and UO_3927 (O_3927,N_48256,N_48764);
nand UO_3928 (O_3928,N_47749,N_47987);
nor UO_3929 (O_3929,N_49304,N_49189);
or UO_3930 (O_3930,N_45520,N_47409);
xor UO_3931 (O_3931,N_45066,N_45512);
and UO_3932 (O_3932,N_49387,N_49058);
nand UO_3933 (O_3933,N_46260,N_48802);
xor UO_3934 (O_3934,N_46191,N_49870);
and UO_3935 (O_3935,N_46631,N_47868);
nor UO_3936 (O_3936,N_47705,N_48997);
xnor UO_3937 (O_3937,N_49685,N_49992);
nor UO_3938 (O_3938,N_45886,N_49409);
nor UO_3939 (O_3939,N_45407,N_46700);
nor UO_3940 (O_3940,N_47830,N_47141);
nand UO_3941 (O_3941,N_46822,N_45895);
or UO_3942 (O_3942,N_45166,N_49014);
and UO_3943 (O_3943,N_47226,N_45517);
and UO_3944 (O_3944,N_48438,N_46463);
and UO_3945 (O_3945,N_45292,N_47468);
nand UO_3946 (O_3946,N_49983,N_46741);
xnor UO_3947 (O_3947,N_46041,N_49640);
and UO_3948 (O_3948,N_45146,N_46762);
or UO_3949 (O_3949,N_49719,N_47548);
xnor UO_3950 (O_3950,N_48329,N_47487);
and UO_3951 (O_3951,N_45159,N_48473);
nand UO_3952 (O_3952,N_47215,N_46362);
or UO_3953 (O_3953,N_47582,N_48870);
nor UO_3954 (O_3954,N_46802,N_48963);
xor UO_3955 (O_3955,N_46277,N_49865);
nor UO_3956 (O_3956,N_47116,N_47570);
nor UO_3957 (O_3957,N_46905,N_49057);
nand UO_3958 (O_3958,N_49019,N_49589);
nor UO_3959 (O_3959,N_48268,N_45812);
and UO_3960 (O_3960,N_48617,N_49192);
nor UO_3961 (O_3961,N_46527,N_46477);
and UO_3962 (O_3962,N_48786,N_46184);
xnor UO_3963 (O_3963,N_49199,N_48073);
xor UO_3964 (O_3964,N_46174,N_49487);
xnor UO_3965 (O_3965,N_45786,N_48484);
nand UO_3966 (O_3966,N_48124,N_47185);
nor UO_3967 (O_3967,N_48013,N_46027);
and UO_3968 (O_3968,N_45165,N_45269);
and UO_3969 (O_3969,N_46248,N_47108);
xor UO_3970 (O_3970,N_48966,N_47296);
nand UO_3971 (O_3971,N_48646,N_47363);
nor UO_3972 (O_3972,N_47624,N_47670);
nor UO_3973 (O_3973,N_45642,N_45118);
or UO_3974 (O_3974,N_49468,N_49727);
or UO_3975 (O_3975,N_47568,N_49396);
and UO_3976 (O_3976,N_46470,N_49085);
and UO_3977 (O_3977,N_46811,N_49890);
xor UO_3978 (O_3978,N_49343,N_48345);
nor UO_3979 (O_3979,N_45189,N_47383);
xnor UO_3980 (O_3980,N_48722,N_45601);
and UO_3981 (O_3981,N_49206,N_45693);
xor UO_3982 (O_3982,N_48248,N_49465);
nor UO_3983 (O_3983,N_48564,N_48647);
nor UO_3984 (O_3984,N_46461,N_45962);
nand UO_3985 (O_3985,N_46085,N_45034);
nand UO_3986 (O_3986,N_49277,N_45171);
nor UO_3987 (O_3987,N_47622,N_48534);
nand UO_3988 (O_3988,N_45135,N_48935);
xor UO_3989 (O_3989,N_49818,N_47590);
xor UO_3990 (O_3990,N_47634,N_48918);
and UO_3991 (O_3991,N_49819,N_48373);
nand UO_3992 (O_3992,N_49731,N_49288);
or UO_3993 (O_3993,N_49771,N_46198);
nor UO_3994 (O_3994,N_47452,N_48131);
nand UO_3995 (O_3995,N_47678,N_49638);
nor UO_3996 (O_3996,N_46422,N_48441);
nor UO_3997 (O_3997,N_49398,N_46988);
or UO_3998 (O_3998,N_48404,N_48231);
xnor UO_3999 (O_3999,N_49171,N_47603);
and UO_4000 (O_4000,N_45432,N_46566);
and UO_4001 (O_4001,N_45050,N_45553);
and UO_4002 (O_4002,N_45464,N_49173);
or UO_4003 (O_4003,N_46804,N_49961);
or UO_4004 (O_4004,N_48675,N_45147);
and UO_4005 (O_4005,N_48356,N_49567);
and UO_4006 (O_4006,N_45195,N_47571);
nand UO_4007 (O_4007,N_49688,N_48962);
or UO_4008 (O_4008,N_45017,N_47249);
or UO_4009 (O_4009,N_47985,N_47595);
xnor UO_4010 (O_4010,N_49723,N_47934);
nand UO_4011 (O_4011,N_45341,N_47831);
and UO_4012 (O_4012,N_45595,N_45372);
nor UO_4013 (O_4013,N_47024,N_49557);
and UO_4014 (O_4014,N_49981,N_48215);
or UO_4015 (O_4015,N_47523,N_49392);
xnor UO_4016 (O_4016,N_46184,N_45242);
or UO_4017 (O_4017,N_48905,N_47294);
nor UO_4018 (O_4018,N_46107,N_47001);
xor UO_4019 (O_4019,N_49373,N_49776);
nand UO_4020 (O_4020,N_46164,N_46144);
and UO_4021 (O_4021,N_48080,N_48050);
or UO_4022 (O_4022,N_47342,N_49671);
and UO_4023 (O_4023,N_48942,N_49410);
nor UO_4024 (O_4024,N_47755,N_46102);
xor UO_4025 (O_4025,N_45682,N_45746);
nor UO_4026 (O_4026,N_47271,N_49550);
xor UO_4027 (O_4027,N_48720,N_48218);
xnor UO_4028 (O_4028,N_45779,N_47684);
and UO_4029 (O_4029,N_46771,N_49594);
and UO_4030 (O_4030,N_49966,N_45915);
or UO_4031 (O_4031,N_45724,N_49257);
and UO_4032 (O_4032,N_49652,N_48191);
and UO_4033 (O_4033,N_47555,N_49063);
nor UO_4034 (O_4034,N_49606,N_48435);
xor UO_4035 (O_4035,N_47553,N_48000);
and UO_4036 (O_4036,N_45214,N_45110);
and UO_4037 (O_4037,N_45808,N_46285);
and UO_4038 (O_4038,N_47326,N_46590);
or UO_4039 (O_4039,N_49753,N_47702);
or UO_4040 (O_4040,N_48039,N_47358);
nand UO_4041 (O_4041,N_47874,N_47291);
nand UO_4042 (O_4042,N_48837,N_46321);
and UO_4043 (O_4043,N_45921,N_47814);
and UO_4044 (O_4044,N_46839,N_46501);
and UO_4045 (O_4045,N_45585,N_49209);
nand UO_4046 (O_4046,N_47085,N_46418);
nand UO_4047 (O_4047,N_46474,N_47909);
nor UO_4048 (O_4048,N_49361,N_46306);
nand UO_4049 (O_4049,N_45884,N_48222);
nand UO_4050 (O_4050,N_49886,N_47770);
or UO_4051 (O_4051,N_47459,N_47528);
and UO_4052 (O_4052,N_49768,N_47938);
xnor UO_4053 (O_4053,N_46655,N_48683);
or UO_4054 (O_4054,N_45941,N_45453);
nor UO_4055 (O_4055,N_46492,N_47827);
xnor UO_4056 (O_4056,N_48223,N_49927);
nor UO_4057 (O_4057,N_47064,N_45701);
or UO_4058 (O_4058,N_45128,N_47320);
nand UO_4059 (O_4059,N_47220,N_49625);
nor UO_4060 (O_4060,N_48944,N_46328);
and UO_4061 (O_4061,N_46580,N_48639);
or UO_4062 (O_4062,N_48162,N_46210);
and UO_4063 (O_4063,N_49756,N_47835);
xor UO_4064 (O_4064,N_49651,N_46432);
and UO_4065 (O_4065,N_48545,N_47276);
xor UO_4066 (O_4066,N_47713,N_46677);
xnor UO_4067 (O_4067,N_49743,N_47159);
nor UO_4068 (O_4068,N_46845,N_49532);
xnor UO_4069 (O_4069,N_49590,N_48992);
xor UO_4070 (O_4070,N_46787,N_47635);
or UO_4071 (O_4071,N_46391,N_45599);
and UO_4072 (O_4072,N_49288,N_47476);
or UO_4073 (O_4073,N_49050,N_47317);
nand UO_4074 (O_4074,N_45199,N_48635);
xor UO_4075 (O_4075,N_49224,N_47952);
and UO_4076 (O_4076,N_45074,N_45030);
xnor UO_4077 (O_4077,N_45204,N_46609);
xnor UO_4078 (O_4078,N_49833,N_48195);
or UO_4079 (O_4079,N_49273,N_47444);
xor UO_4080 (O_4080,N_48116,N_48105);
nand UO_4081 (O_4081,N_49268,N_49050);
xnor UO_4082 (O_4082,N_48454,N_48386);
xor UO_4083 (O_4083,N_48007,N_48199);
nor UO_4084 (O_4084,N_46138,N_48191);
nor UO_4085 (O_4085,N_47087,N_49693);
and UO_4086 (O_4086,N_46018,N_45893);
and UO_4087 (O_4087,N_47452,N_47741);
xor UO_4088 (O_4088,N_45263,N_48502);
xnor UO_4089 (O_4089,N_46509,N_48334);
xnor UO_4090 (O_4090,N_48728,N_46529);
nand UO_4091 (O_4091,N_48527,N_49966);
and UO_4092 (O_4092,N_46856,N_46751);
nand UO_4093 (O_4093,N_49353,N_46948);
and UO_4094 (O_4094,N_47974,N_48195);
or UO_4095 (O_4095,N_45371,N_48583);
or UO_4096 (O_4096,N_48647,N_46363);
nor UO_4097 (O_4097,N_48830,N_48365);
nand UO_4098 (O_4098,N_49986,N_46740);
xor UO_4099 (O_4099,N_46738,N_49310);
and UO_4100 (O_4100,N_48273,N_45600);
xor UO_4101 (O_4101,N_47520,N_46370);
or UO_4102 (O_4102,N_45896,N_47754);
xor UO_4103 (O_4103,N_46477,N_49910);
nor UO_4104 (O_4104,N_49201,N_49703);
and UO_4105 (O_4105,N_45503,N_45494);
xor UO_4106 (O_4106,N_47876,N_49404);
and UO_4107 (O_4107,N_48967,N_48239);
nand UO_4108 (O_4108,N_47005,N_45945);
nor UO_4109 (O_4109,N_48812,N_49348);
or UO_4110 (O_4110,N_48106,N_47133);
nor UO_4111 (O_4111,N_46779,N_46943);
nand UO_4112 (O_4112,N_46134,N_47412);
xnor UO_4113 (O_4113,N_49881,N_46017);
xnor UO_4114 (O_4114,N_48201,N_46953);
or UO_4115 (O_4115,N_49060,N_48802);
xor UO_4116 (O_4116,N_47885,N_45311);
nor UO_4117 (O_4117,N_49985,N_47538);
xor UO_4118 (O_4118,N_46507,N_48530);
or UO_4119 (O_4119,N_48936,N_46062);
nand UO_4120 (O_4120,N_46092,N_45347);
xnor UO_4121 (O_4121,N_47795,N_48280);
and UO_4122 (O_4122,N_47808,N_45811);
nor UO_4123 (O_4123,N_48167,N_46379);
nor UO_4124 (O_4124,N_48617,N_48181);
nand UO_4125 (O_4125,N_46284,N_46343);
and UO_4126 (O_4126,N_49451,N_45830);
nor UO_4127 (O_4127,N_46313,N_49475);
and UO_4128 (O_4128,N_49690,N_45408);
xnor UO_4129 (O_4129,N_46783,N_48566);
xor UO_4130 (O_4130,N_48280,N_48663);
nor UO_4131 (O_4131,N_47699,N_49202);
or UO_4132 (O_4132,N_48207,N_48318);
and UO_4133 (O_4133,N_47622,N_46782);
and UO_4134 (O_4134,N_45417,N_46345);
nand UO_4135 (O_4135,N_48663,N_48549);
nor UO_4136 (O_4136,N_49485,N_49840);
or UO_4137 (O_4137,N_45612,N_47897);
nand UO_4138 (O_4138,N_45471,N_47929);
nand UO_4139 (O_4139,N_45659,N_47395);
nor UO_4140 (O_4140,N_49025,N_46166);
nor UO_4141 (O_4141,N_47886,N_46450);
or UO_4142 (O_4142,N_48611,N_46140);
nor UO_4143 (O_4143,N_49869,N_49183);
nor UO_4144 (O_4144,N_46315,N_47717);
and UO_4145 (O_4145,N_46009,N_49660);
or UO_4146 (O_4146,N_45876,N_49778);
and UO_4147 (O_4147,N_46007,N_48523);
or UO_4148 (O_4148,N_46500,N_45678);
and UO_4149 (O_4149,N_49239,N_46807);
nor UO_4150 (O_4150,N_48668,N_45706);
xnor UO_4151 (O_4151,N_48269,N_45279);
and UO_4152 (O_4152,N_45151,N_48603);
and UO_4153 (O_4153,N_48861,N_47907);
xnor UO_4154 (O_4154,N_46450,N_46665);
nand UO_4155 (O_4155,N_46466,N_48637);
and UO_4156 (O_4156,N_47492,N_45244);
nor UO_4157 (O_4157,N_47657,N_45131);
xnor UO_4158 (O_4158,N_49150,N_46562);
and UO_4159 (O_4159,N_48431,N_47768);
and UO_4160 (O_4160,N_46690,N_48604);
xor UO_4161 (O_4161,N_47782,N_46573);
xnor UO_4162 (O_4162,N_48364,N_48120);
and UO_4163 (O_4163,N_45778,N_47838);
xnor UO_4164 (O_4164,N_46269,N_49604);
xnor UO_4165 (O_4165,N_48748,N_47586);
or UO_4166 (O_4166,N_48020,N_45113);
nand UO_4167 (O_4167,N_45643,N_45517);
nor UO_4168 (O_4168,N_47870,N_48027);
xor UO_4169 (O_4169,N_45673,N_47615);
and UO_4170 (O_4170,N_48026,N_46768);
and UO_4171 (O_4171,N_49882,N_45354);
nor UO_4172 (O_4172,N_47339,N_45764);
or UO_4173 (O_4173,N_46982,N_45698);
or UO_4174 (O_4174,N_49970,N_45677);
nor UO_4175 (O_4175,N_46441,N_45588);
nor UO_4176 (O_4176,N_49346,N_47220);
nand UO_4177 (O_4177,N_45522,N_49430);
xnor UO_4178 (O_4178,N_47776,N_46206);
or UO_4179 (O_4179,N_48266,N_47524);
nand UO_4180 (O_4180,N_45221,N_47132);
or UO_4181 (O_4181,N_45734,N_45024);
nor UO_4182 (O_4182,N_48245,N_48102);
xor UO_4183 (O_4183,N_47879,N_46222);
or UO_4184 (O_4184,N_48277,N_45162);
and UO_4185 (O_4185,N_45704,N_45678);
or UO_4186 (O_4186,N_49107,N_45790);
nand UO_4187 (O_4187,N_47059,N_48404);
and UO_4188 (O_4188,N_47582,N_45967);
or UO_4189 (O_4189,N_46274,N_49676);
nor UO_4190 (O_4190,N_47342,N_45119);
xnor UO_4191 (O_4191,N_48359,N_47643);
and UO_4192 (O_4192,N_45268,N_48454);
xor UO_4193 (O_4193,N_47016,N_47405);
xor UO_4194 (O_4194,N_45155,N_48597);
nor UO_4195 (O_4195,N_46994,N_47383);
nor UO_4196 (O_4196,N_45616,N_48013);
xnor UO_4197 (O_4197,N_45205,N_49204);
nor UO_4198 (O_4198,N_47469,N_49806);
and UO_4199 (O_4199,N_47723,N_48126);
and UO_4200 (O_4200,N_47940,N_46898);
nand UO_4201 (O_4201,N_46949,N_46058);
xor UO_4202 (O_4202,N_45770,N_47510);
nand UO_4203 (O_4203,N_48724,N_46041);
nand UO_4204 (O_4204,N_48034,N_45752);
nand UO_4205 (O_4205,N_47845,N_48169);
xnor UO_4206 (O_4206,N_49994,N_45148);
nand UO_4207 (O_4207,N_48196,N_47813);
nor UO_4208 (O_4208,N_48149,N_47089);
xnor UO_4209 (O_4209,N_48959,N_46291);
xor UO_4210 (O_4210,N_48439,N_46481);
or UO_4211 (O_4211,N_49093,N_49667);
xnor UO_4212 (O_4212,N_46025,N_47107);
xnor UO_4213 (O_4213,N_45140,N_45709);
and UO_4214 (O_4214,N_47752,N_45252);
xor UO_4215 (O_4215,N_45954,N_48108);
or UO_4216 (O_4216,N_45234,N_45500);
nor UO_4217 (O_4217,N_49467,N_49454);
and UO_4218 (O_4218,N_49396,N_45330);
nor UO_4219 (O_4219,N_48310,N_49563);
nor UO_4220 (O_4220,N_47041,N_45257);
nor UO_4221 (O_4221,N_47302,N_45966);
and UO_4222 (O_4222,N_48723,N_48444);
nand UO_4223 (O_4223,N_48716,N_49919);
or UO_4224 (O_4224,N_47088,N_48854);
nor UO_4225 (O_4225,N_45393,N_48259);
or UO_4226 (O_4226,N_45241,N_48183);
nor UO_4227 (O_4227,N_47797,N_47153);
nor UO_4228 (O_4228,N_48929,N_47857);
nor UO_4229 (O_4229,N_47947,N_45788);
nand UO_4230 (O_4230,N_45982,N_49273);
or UO_4231 (O_4231,N_48177,N_48484);
and UO_4232 (O_4232,N_49891,N_48990);
nor UO_4233 (O_4233,N_46585,N_45190);
xnor UO_4234 (O_4234,N_49435,N_45146);
xor UO_4235 (O_4235,N_47491,N_47180);
xnor UO_4236 (O_4236,N_49654,N_46309);
xnor UO_4237 (O_4237,N_49356,N_47629);
and UO_4238 (O_4238,N_45246,N_46740);
nand UO_4239 (O_4239,N_48831,N_46095);
xnor UO_4240 (O_4240,N_47134,N_47647);
xor UO_4241 (O_4241,N_48193,N_49991);
or UO_4242 (O_4242,N_46916,N_48803);
nor UO_4243 (O_4243,N_46388,N_49054);
or UO_4244 (O_4244,N_48297,N_48055);
nand UO_4245 (O_4245,N_48307,N_45822);
or UO_4246 (O_4246,N_49540,N_45572);
and UO_4247 (O_4247,N_46715,N_47493);
and UO_4248 (O_4248,N_46047,N_45975);
or UO_4249 (O_4249,N_47822,N_47213);
nand UO_4250 (O_4250,N_48558,N_48147);
nor UO_4251 (O_4251,N_47991,N_46138);
and UO_4252 (O_4252,N_47411,N_47704);
nor UO_4253 (O_4253,N_49017,N_45824);
nand UO_4254 (O_4254,N_48329,N_46553);
nand UO_4255 (O_4255,N_49308,N_49134);
nor UO_4256 (O_4256,N_49530,N_45764);
nand UO_4257 (O_4257,N_49039,N_49292);
or UO_4258 (O_4258,N_46789,N_49395);
or UO_4259 (O_4259,N_49931,N_46991);
xnor UO_4260 (O_4260,N_45311,N_46572);
and UO_4261 (O_4261,N_49051,N_46843);
nand UO_4262 (O_4262,N_48705,N_49891);
and UO_4263 (O_4263,N_47934,N_48697);
nand UO_4264 (O_4264,N_46720,N_47256);
nor UO_4265 (O_4265,N_49610,N_47049);
and UO_4266 (O_4266,N_45186,N_49575);
nand UO_4267 (O_4267,N_49999,N_46697);
or UO_4268 (O_4268,N_49291,N_47960);
nor UO_4269 (O_4269,N_48818,N_46195);
or UO_4270 (O_4270,N_45647,N_47202);
xnor UO_4271 (O_4271,N_46299,N_47448);
or UO_4272 (O_4272,N_49606,N_45880);
nor UO_4273 (O_4273,N_47615,N_46390);
or UO_4274 (O_4274,N_47184,N_46592);
nor UO_4275 (O_4275,N_48815,N_47532);
nand UO_4276 (O_4276,N_45846,N_47593);
xnor UO_4277 (O_4277,N_49155,N_46371);
nor UO_4278 (O_4278,N_49721,N_48129);
nand UO_4279 (O_4279,N_48804,N_46623);
and UO_4280 (O_4280,N_47584,N_49535);
xnor UO_4281 (O_4281,N_45870,N_49607);
nor UO_4282 (O_4282,N_47949,N_46048);
and UO_4283 (O_4283,N_48615,N_45263);
or UO_4284 (O_4284,N_48797,N_48704);
xor UO_4285 (O_4285,N_47128,N_47422);
and UO_4286 (O_4286,N_48088,N_46773);
nand UO_4287 (O_4287,N_47408,N_47103);
nand UO_4288 (O_4288,N_48204,N_46430);
and UO_4289 (O_4289,N_48947,N_45356);
and UO_4290 (O_4290,N_47098,N_48585);
xnor UO_4291 (O_4291,N_48049,N_47733);
or UO_4292 (O_4292,N_49093,N_46838);
nor UO_4293 (O_4293,N_48968,N_49474);
nand UO_4294 (O_4294,N_45625,N_45388);
xor UO_4295 (O_4295,N_47856,N_48720);
xnor UO_4296 (O_4296,N_46298,N_49998);
nand UO_4297 (O_4297,N_46735,N_47723);
nor UO_4298 (O_4298,N_48063,N_49178);
or UO_4299 (O_4299,N_48390,N_45051);
nor UO_4300 (O_4300,N_46129,N_45948);
or UO_4301 (O_4301,N_46121,N_45438);
and UO_4302 (O_4302,N_47585,N_47706);
nor UO_4303 (O_4303,N_45170,N_49208);
and UO_4304 (O_4304,N_46114,N_49568);
or UO_4305 (O_4305,N_48306,N_45903);
nor UO_4306 (O_4306,N_47824,N_48945);
nor UO_4307 (O_4307,N_47593,N_46108);
and UO_4308 (O_4308,N_46640,N_45371);
and UO_4309 (O_4309,N_45770,N_45149);
nor UO_4310 (O_4310,N_47834,N_48369);
nor UO_4311 (O_4311,N_46880,N_47216);
or UO_4312 (O_4312,N_49445,N_46867);
or UO_4313 (O_4313,N_49861,N_48066);
or UO_4314 (O_4314,N_47493,N_45912);
xor UO_4315 (O_4315,N_47229,N_47689);
and UO_4316 (O_4316,N_47833,N_47257);
or UO_4317 (O_4317,N_46482,N_45227);
or UO_4318 (O_4318,N_48070,N_45601);
or UO_4319 (O_4319,N_45482,N_45851);
or UO_4320 (O_4320,N_45403,N_46200);
nand UO_4321 (O_4321,N_48969,N_47238);
nand UO_4322 (O_4322,N_48457,N_45587);
nor UO_4323 (O_4323,N_45523,N_48042);
and UO_4324 (O_4324,N_49593,N_49882);
nand UO_4325 (O_4325,N_49240,N_49301);
xnor UO_4326 (O_4326,N_45214,N_45964);
nor UO_4327 (O_4327,N_49792,N_46772);
or UO_4328 (O_4328,N_49697,N_47190);
nor UO_4329 (O_4329,N_45989,N_47917);
or UO_4330 (O_4330,N_47854,N_45329);
or UO_4331 (O_4331,N_49770,N_46694);
nor UO_4332 (O_4332,N_48890,N_48865);
nor UO_4333 (O_4333,N_45618,N_47566);
and UO_4334 (O_4334,N_48355,N_45954);
nor UO_4335 (O_4335,N_49732,N_47216);
xor UO_4336 (O_4336,N_46299,N_46328);
nand UO_4337 (O_4337,N_46690,N_47860);
and UO_4338 (O_4338,N_45427,N_49309);
or UO_4339 (O_4339,N_49134,N_49582);
xor UO_4340 (O_4340,N_46668,N_48358);
and UO_4341 (O_4341,N_46570,N_48407);
xor UO_4342 (O_4342,N_48720,N_49608);
nor UO_4343 (O_4343,N_46706,N_47426);
nand UO_4344 (O_4344,N_46524,N_49574);
nand UO_4345 (O_4345,N_45607,N_47533);
and UO_4346 (O_4346,N_47430,N_46536);
nor UO_4347 (O_4347,N_47649,N_48452);
or UO_4348 (O_4348,N_48467,N_48379);
and UO_4349 (O_4349,N_46305,N_46673);
or UO_4350 (O_4350,N_48099,N_49160);
nor UO_4351 (O_4351,N_47442,N_48007);
or UO_4352 (O_4352,N_49185,N_45420);
nand UO_4353 (O_4353,N_46728,N_45157);
nor UO_4354 (O_4354,N_47357,N_47813);
nor UO_4355 (O_4355,N_49676,N_47743);
nand UO_4356 (O_4356,N_45658,N_47603);
nor UO_4357 (O_4357,N_47197,N_48333);
nor UO_4358 (O_4358,N_48838,N_48098);
or UO_4359 (O_4359,N_46663,N_48397);
or UO_4360 (O_4360,N_48169,N_46609);
nand UO_4361 (O_4361,N_47195,N_48575);
or UO_4362 (O_4362,N_46590,N_46443);
or UO_4363 (O_4363,N_49600,N_48163);
and UO_4364 (O_4364,N_47130,N_45617);
nor UO_4365 (O_4365,N_49660,N_49227);
xnor UO_4366 (O_4366,N_47441,N_47704);
and UO_4367 (O_4367,N_46273,N_47189);
or UO_4368 (O_4368,N_49454,N_49733);
and UO_4369 (O_4369,N_48095,N_47611);
and UO_4370 (O_4370,N_49506,N_46831);
nor UO_4371 (O_4371,N_48082,N_47961);
and UO_4372 (O_4372,N_49073,N_49366);
nor UO_4373 (O_4373,N_49603,N_46531);
and UO_4374 (O_4374,N_49971,N_48701);
nand UO_4375 (O_4375,N_47299,N_47475);
nand UO_4376 (O_4376,N_46570,N_46104);
nor UO_4377 (O_4377,N_45957,N_47706);
or UO_4378 (O_4378,N_48559,N_48897);
and UO_4379 (O_4379,N_48935,N_48731);
or UO_4380 (O_4380,N_45144,N_47175);
nor UO_4381 (O_4381,N_47675,N_47973);
nand UO_4382 (O_4382,N_45396,N_48619);
and UO_4383 (O_4383,N_46621,N_46978);
and UO_4384 (O_4384,N_47662,N_47934);
nor UO_4385 (O_4385,N_47877,N_46469);
and UO_4386 (O_4386,N_48960,N_45652);
or UO_4387 (O_4387,N_49327,N_45477);
xnor UO_4388 (O_4388,N_47916,N_47509);
nand UO_4389 (O_4389,N_48422,N_46645);
and UO_4390 (O_4390,N_45329,N_49326);
nor UO_4391 (O_4391,N_48135,N_46905);
xor UO_4392 (O_4392,N_49026,N_45046);
or UO_4393 (O_4393,N_48244,N_46621);
nor UO_4394 (O_4394,N_45130,N_45339);
xor UO_4395 (O_4395,N_48287,N_47353);
or UO_4396 (O_4396,N_46142,N_49650);
xnor UO_4397 (O_4397,N_49538,N_46249);
xor UO_4398 (O_4398,N_48290,N_47374);
nor UO_4399 (O_4399,N_45875,N_49339);
or UO_4400 (O_4400,N_47123,N_46913);
and UO_4401 (O_4401,N_48079,N_47799);
xor UO_4402 (O_4402,N_49110,N_46950);
nand UO_4403 (O_4403,N_49068,N_49781);
or UO_4404 (O_4404,N_48635,N_49633);
nor UO_4405 (O_4405,N_49449,N_48832);
nand UO_4406 (O_4406,N_47844,N_47135);
xnor UO_4407 (O_4407,N_46595,N_47361);
xnor UO_4408 (O_4408,N_46791,N_47589);
or UO_4409 (O_4409,N_45920,N_46847);
and UO_4410 (O_4410,N_49666,N_49778);
nor UO_4411 (O_4411,N_47023,N_49122);
and UO_4412 (O_4412,N_49556,N_46212);
or UO_4413 (O_4413,N_45243,N_46494);
nand UO_4414 (O_4414,N_49746,N_48979);
nor UO_4415 (O_4415,N_48903,N_47691);
and UO_4416 (O_4416,N_48087,N_46539);
and UO_4417 (O_4417,N_49919,N_49386);
xnor UO_4418 (O_4418,N_46418,N_47770);
nor UO_4419 (O_4419,N_48136,N_46796);
xor UO_4420 (O_4420,N_47024,N_46748);
nand UO_4421 (O_4421,N_45235,N_47378);
nand UO_4422 (O_4422,N_48808,N_48974);
nor UO_4423 (O_4423,N_48633,N_49976);
nand UO_4424 (O_4424,N_47019,N_46696);
nand UO_4425 (O_4425,N_45656,N_45560);
or UO_4426 (O_4426,N_48153,N_47226);
or UO_4427 (O_4427,N_45630,N_48674);
xor UO_4428 (O_4428,N_48949,N_45843);
nor UO_4429 (O_4429,N_48021,N_45056);
and UO_4430 (O_4430,N_49652,N_49897);
nor UO_4431 (O_4431,N_46130,N_49936);
nand UO_4432 (O_4432,N_48529,N_46244);
nor UO_4433 (O_4433,N_49154,N_46316);
nor UO_4434 (O_4434,N_48465,N_45071);
and UO_4435 (O_4435,N_45394,N_46088);
xnor UO_4436 (O_4436,N_47348,N_46713);
nor UO_4437 (O_4437,N_49110,N_45809);
nor UO_4438 (O_4438,N_46622,N_45074);
nand UO_4439 (O_4439,N_45892,N_46889);
nor UO_4440 (O_4440,N_49967,N_48588);
and UO_4441 (O_4441,N_48390,N_49125);
nor UO_4442 (O_4442,N_48914,N_47716);
and UO_4443 (O_4443,N_45723,N_46741);
nand UO_4444 (O_4444,N_49783,N_47239);
nand UO_4445 (O_4445,N_45449,N_46395);
xor UO_4446 (O_4446,N_47026,N_48213);
nor UO_4447 (O_4447,N_48575,N_45135);
xor UO_4448 (O_4448,N_48866,N_45585);
and UO_4449 (O_4449,N_49014,N_45727);
or UO_4450 (O_4450,N_49517,N_45254);
xnor UO_4451 (O_4451,N_48782,N_48760);
nand UO_4452 (O_4452,N_47205,N_45709);
nor UO_4453 (O_4453,N_46587,N_46474);
nand UO_4454 (O_4454,N_49750,N_46465);
nor UO_4455 (O_4455,N_49461,N_46571);
or UO_4456 (O_4456,N_49284,N_47564);
nor UO_4457 (O_4457,N_48474,N_49785);
or UO_4458 (O_4458,N_47963,N_49238);
nor UO_4459 (O_4459,N_49594,N_47976);
and UO_4460 (O_4460,N_45979,N_47951);
xor UO_4461 (O_4461,N_45692,N_47243);
nor UO_4462 (O_4462,N_48424,N_49781);
or UO_4463 (O_4463,N_47156,N_49267);
or UO_4464 (O_4464,N_46817,N_45103);
or UO_4465 (O_4465,N_49664,N_48647);
nand UO_4466 (O_4466,N_45880,N_47144);
or UO_4467 (O_4467,N_45570,N_47981);
or UO_4468 (O_4468,N_47695,N_47682);
xnor UO_4469 (O_4469,N_46196,N_45026);
xnor UO_4470 (O_4470,N_46402,N_45008);
nor UO_4471 (O_4471,N_49755,N_47728);
nor UO_4472 (O_4472,N_45510,N_46885);
nor UO_4473 (O_4473,N_45305,N_45815);
nand UO_4474 (O_4474,N_45258,N_48541);
nand UO_4475 (O_4475,N_46792,N_49789);
nor UO_4476 (O_4476,N_47482,N_46234);
or UO_4477 (O_4477,N_45368,N_45265);
nand UO_4478 (O_4478,N_46970,N_49571);
and UO_4479 (O_4479,N_49039,N_48302);
xor UO_4480 (O_4480,N_48107,N_47331);
xor UO_4481 (O_4481,N_47034,N_48605);
xnor UO_4482 (O_4482,N_49316,N_47418);
and UO_4483 (O_4483,N_47338,N_47627);
nor UO_4484 (O_4484,N_48882,N_45241);
or UO_4485 (O_4485,N_45795,N_48788);
xnor UO_4486 (O_4486,N_48182,N_46897);
nor UO_4487 (O_4487,N_45629,N_46467);
nor UO_4488 (O_4488,N_47849,N_45692);
xnor UO_4489 (O_4489,N_45105,N_49433);
nand UO_4490 (O_4490,N_46791,N_47351);
and UO_4491 (O_4491,N_46744,N_45789);
and UO_4492 (O_4492,N_48049,N_48766);
nand UO_4493 (O_4493,N_46782,N_48950);
xor UO_4494 (O_4494,N_45569,N_48491);
or UO_4495 (O_4495,N_47715,N_46791);
and UO_4496 (O_4496,N_46959,N_46443);
or UO_4497 (O_4497,N_46138,N_48469);
xor UO_4498 (O_4498,N_47016,N_49832);
nand UO_4499 (O_4499,N_45055,N_48846);
xor UO_4500 (O_4500,N_48660,N_47818);
nor UO_4501 (O_4501,N_45050,N_45973);
xor UO_4502 (O_4502,N_46160,N_48583);
or UO_4503 (O_4503,N_45401,N_45840);
or UO_4504 (O_4504,N_49265,N_47375);
xor UO_4505 (O_4505,N_45959,N_49597);
nor UO_4506 (O_4506,N_49510,N_48484);
xnor UO_4507 (O_4507,N_47572,N_45456);
xnor UO_4508 (O_4508,N_49040,N_49018);
xor UO_4509 (O_4509,N_46259,N_48669);
and UO_4510 (O_4510,N_45926,N_48629);
xor UO_4511 (O_4511,N_48414,N_49804);
xor UO_4512 (O_4512,N_46732,N_45664);
and UO_4513 (O_4513,N_46646,N_49186);
and UO_4514 (O_4514,N_47821,N_47726);
or UO_4515 (O_4515,N_47257,N_46877);
and UO_4516 (O_4516,N_46653,N_46562);
and UO_4517 (O_4517,N_47131,N_49393);
nor UO_4518 (O_4518,N_47106,N_45764);
nor UO_4519 (O_4519,N_46506,N_47255);
nor UO_4520 (O_4520,N_46819,N_46338);
nand UO_4521 (O_4521,N_45348,N_47961);
and UO_4522 (O_4522,N_47729,N_49628);
nor UO_4523 (O_4523,N_49536,N_49303);
nand UO_4524 (O_4524,N_47599,N_49782);
xnor UO_4525 (O_4525,N_49783,N_49635);
nor UO_4526 (O_4526,N_49729,N_49914);
and UO_4527 (O_4527,N_45407,N_45230);
nand UO_4528 (O_4528,N_48100,N_46945);
and UO_4529 (O_4529,N_49888,N_46398);
nor UO_4530 (O_4530,N_48760,N_49114);
and UO_4531 (O_4531,N_46110,N_46736);
xor UO_4532 (O_4532,N_45631,N_45792);
nand UO_4533 (O_4533,N_48141,N_49708);
and UO_4534 (O_4534,N_47191,N_46536);
and UO_4535 (O_4535,N_48407,N_45184);
nand UO_4536 (O_4536,N_46173,N_49326);
or UO_4537 (O_4537,N_48765,N_45777);
and UO_4538 (O_4538,N_47391,N_46471);
and UO_4539 (O_4539,N_46094,N_47796);
or UO_4540 (O_4540,N_45016,N_46263);
or UO_4541 (O_4541,N_46682,N_49353);
or UO_4542 (O_4542,N_47740,N_47504);
nor UO_4543 (O_4543,N_46738,N_45928);
nor UO_4544 (O_4544,N_49408,N_45020);
nor UO_4545 (O_4545,N_48519,N_49769);
nand UO_4546 (O_4546,N_46152,N_46091);
nor UO_4547 (O_4547,N_47953,N_46330);
xor UO_4548 (O_4548,N_49532,N_46855);
and UO_4549 (O_4549,N_45077,N_47934);
nand UO_4550 (O_4550,N_49254,N_47132);
or UO_4551 (O_4551,N_48871,N_46892);
nand UO_4552 (O_4552,N_48193,N_48679);
nor UO_4553 (O_4553,N_49984,N_45369);
xor UO_4554 (O_4554,N_46196,N_47143);
or UO_4555 (O_4555,N_48953,N_46080);
and UO_4556 (O_4556,N_46010,N_45706);
and UO_4557 (O_4557,N_46709,N_45780);
nand UO_4558 (O_4558,N_45003,N_45880);
and UO_4559 (O_4559,N_46262,N_47371);
and UO_4560 (O_4560,N_46541,N_45207);
or UO_4561 (O_4561,N_47730,N_49858);
nor UO_4562 (O_4562,N_47909,N_49182);
nor UO_4563 (O_4563,N_48316,N_49459);
and UO_4564 (O_4564,N_48471,N_47308);
nor UO_4565 (O_4565,N_47341,N_48886);
nor UO_4566 (O_4566,N_49951,N_49677);
nor UO_4567 (O_4567,N_45616,N_46442);
or UO_4568 (O_4568,N_48794,N_48693);
nor UO_4569 (O_4569,N_47010,N_45431);
and UO_4570 (O_4570,N_45045,N_49238);
and UO_4571 (O_4571,N_49815,N_47480);
nor UO_4572 (O_4572,N_48844,N_48242);
nor UO_4573 (O_4573,N_45629,N_45166);
xor UO_4574 (O_4574,N_47495,N_45508);
nand UO_4575 (O_4575,N_45204,N_46276);
and UO_4576 (O_4576,N_48138,N_49444);
nor UO_4577 (O_4577,N_45254,N_48548);
and UO_4578 (O_4578,N_49930,N_46724);
and UO_4579 (O_4579,N_45438,N_45489);
nor UO_4580 (O_4580,N_48040,N_48727);
and UO_4581 (O_4581,N_45634,N_47060);
nand UO_4582 (O_4582,N_49671,N_48882);
nand UO_4583 (O_4583,N_48307,N_48705);
nor UO_4584 (O_4584,N_46217,N_45343);
nor UO_4585 (O_4585,N_45036,N_45936);
and UO_4586 (O_4586,N_46389,N_48057);
nand UO_4587 (O_4587,N_48131,N_45448);
nor UO_4588 (O_4588,N_47260,N_48593);
and UO_4589 (O_4589,N_47380,N_49006);
nor UO_4590 (O_4590,N_46988,N_46945);
nand UO_4591 (O_4591,N_46166,N_48609);
and UO_4592 (O_4592,N_46459,N_49378);
and UO_4593 (O_4593,N_47762,N_45996);
or UO_4594 (O_4594,N_46500,N_45384);
nor UO_4595 (O_4595,N_49196,N_47359);
and UO_4596 (O_4596,N_46480,N_46156);
nor UO_4597 (O_4597,N_47306,N_47529);
or UO_4598 (O_4598,N_49401,N_48190);
or UO_4599 (O_4599,N_49832,N_45802);
and UO_4600 (O_4600,N_45972,N_45484);
or UO_4601 (O_4601,N_47170,N_49651);
nand UO_4602 (O_4602,N_48712,N_48622);
or UO_4603 (O_4603,N_48816,N_46680);
and UO_4604 (O_4604,N_48078,N_48934);
nand UO_4605 (O_4605,N_48847,N_45444);
and UO_4606 (O_4606,N_46201,N_46270);
xnor UO_4607 (O_4607,N_48654,N_47013);
or UO_4608 (O_4608,N_48561,N_45746);
xnor UO_4609 (O_4609,N_46554,N_46912);
or UO_4610 (O_4610,N_45089,N_45842);
or UO_4611 (O_4611,N_46589,N_45501);
and UO_4612 (O_4612,N_47865,N_45899);
nand UO_4613 (O_4613,N_49071,N_45554);
xor UO_4614 (O_4614,N_48027,N_47333);
and UO_4615 (O_4615,N_47059,N_49667);
nand UO_4616 (O_4616,N_46928,N_49374);
nor UO_4617 (O_4617,N_47280,N_45004);
nor UO_4618 (O_4618,N_48771,N_45718);
nor UO_4619 (O_4619,N_45194,N_47511);
xor UO_4620 (O_4620,N_46510,N_46479);
nor UO_4621 (O_4621,N_46765,N_47729);
nand UO_4622 (O_4622,N_46972,N_47651);
nor UO_4623 (O_4623,N_49346,N_47625);
nand UO_4624 (O_4624,N_47483,N_47128);
xnor UO_4625 (O_4625,N_45323,N_49035);
xnor UO_4626 (O_4626,N_48687,N_49208);
nand UO_4627 (O_4627,N_45946,N_46620);
and UO_4628 (O_4628,N_47774,N_47574);
xnor UO_4629 (O_4629,N_47400,N_46832);
or UO_4630 (O_4630,N_45940,N_45287);
nor UO_4631 (O_4631,N_46022,N_48543);
xor UO_4632 (O_4632,N_49760,N_47555);
nor UO_4633 (O_4633,N_49089,N_47589);
nor UO_4634 (O_4634,N_47482,N_49191);
nor UO_4635 (O_4635,N_45909,N_48696);
or UO_4636 (O_4636,N_46303,N_46409);
xnor UO_4637 (O_4637,N_49468,N_46567);
or UO_4638 (O_4638,N_45559,N_46531);
xnor UO_4639 (O_4639,N_46939,N_47836);
nand UO_4640 (O_4640,N_49749,N_49907);
nor UO_4641 (O_4641,N_45089,N_45362);
nand UO_4642 (O_4642,N_46027,N_45817);
or UO_4643 (O_4643,N_47590,N_48135);
nor UO_4644 (O_4644,N_47205,N_45315);
nor UO_4645 (O_4645,N_49621,N_49668);
or UO_4646 (O_4646,N_45623,N_49547);
or UO_4647 (O_4647,N_49681,N_47712);
and UO_4648 (O_4648,N_49422,N_47660);
xnor UO_4649 (O_4649,N_47743,N_49022);
nand UO_4650 (O_4650,N_48640,N_46493);
xor UO_4651 (O_4651,N_45794,N_49650);
nand UO_4652 (O_4652,N_47452,N_46940);
nor UO_4653 (O_4653,N_47690,N_46818);
xnor UO_4654 (O_4654,N_48083,N_45374);
nor UO_4655 (O_4655,N_47382,N_45815);
nor UO_4656 (O_4656,N_49837,N_49031);
or UO_4657 (O_4657,N_45389,N_45843);
nor UO_4658 (O_4658,N_49831,N_45033);
and UO_4659 (O_4659,N_47240,N_46829);
xnor UO_4660 (O_4660,N_49821,N_46126);
and UO_4661 (O_4661,N_47093,N_46759);
nor UO_4662 (O_4662,N_49816,N_49980);
nand UO_4663 (O_4663,N_46002,N_48080);
or UO_4664 (O_4664,N_49151,N_47626);
or UO_4665 (O_4665,N_46584,N_45617);
and UO_4666 (O_4666,N_46767,N_48372);
or UO_4667 (O_4667,N_49219,N_47467);
nor UO_4668 (O_4668,N_47745,N_45380);
nand UO_4669 (O_4669,N_47653,N_47024);
and UO_4670 (O_4670,N_46620,N_49852);
xor UO_4671 (O_4671,N_49037,N_45456);
nor UO_4672 (O_4672,N_47634,N_47136);
xnor UO_4673 (O_4673,N_46353,N_47415);
or UO_4674 (O_4674,N_47638,N_48189);
or UO_4675 (O_4675,N_45291,N_45059);
and UO_4676 (O_4676,N_46998,N_47109);
xnor UO_4677 (O_4677,N_47328,N_49232);
nand UO_4678 (O_4678,N_49603,N_45310);
and UO_4679 (O_4679,N_48752,N_47387);
or UO_4680 (O_4680,N_47393,N_49796);
and UO_4681 (O_4681,N_49389,N_48524);
and UO_4682 (O_4682,N_47283,N_47277);
or UO_4683 (O_4683,N_48281,N_49530);
and UO_4684 (O_4684,N_47196,N_48230);
nor UO_4685 (O_4685,N_45178,N_49229);
nor UO_4686 (O_4686,N_45864,N_47322);
or UO_4687 (O_4687,N_46641,N_48837);
or UO_4688 (O_4688,N_48179,N_49865);
nand UO_4689 (O_4689,N_46916,N_47644);
and UO_4690 (O_4690,N_49397,N_48030);
nand UO_4691 (O_4691,N_48326,N_46118);
nand UO_4692 (O_4692,N_46112,N_48128);
or UO_4693 (O_4693,N_48356,N_48994);
or UO_4694 (O_4694,N_45063,N_46026);
and UO_4695 (O_4695,N_48175,N_45581);
nand UO_4696 (O_4696,N_45255,N_46020);
or UO_4697 (O_4697,N_45792,N_48654);
nor UO_4698 (O_4698,N_47906,N_48290);
nand UO_4699 (O_4699,N_46953,N_48521);
nor UO_4700 (O_4700,N_49175,N_47472);
nand UO_4701 (O_4701,N_46908,N_48631);
nand UO_4702 (O_4702,N_49179,N_48223);
nand UO_4703 (O_4703,N_48225,N_48733);
or UO_4704 (O_4704,N_46622,N_46761);
nand UO_4705 (O_4705,N_45176,N_48235);
nor UO_4706 (O_4706,N_47550,N_48493);
or UO_4707 (O_4707,N_46005,N_48713);
or UO_4708 (O_4708,N_45524,N_46142);
and UO_4709 (O_4709,N_45669,N_46683);
xor UO_4710 (O_4710,N_48970,N_48922);
or UO_4711 (O_4711,N_47460,N_45841);
nand UO_4712 (O_4712,N_46702,N_47212);
nand UO_4713 (O_4713,N_47214,N_49451);
nor UO_4714 (O_4714,N_47799,N_48929);
xnor UO_4715 (O_4715,N_49468,N_45921);
nor UO_4716 (O_4716,N_49530,N_48645);
and UO_4717 (O_4717,N_48494,N_47193);
nor UO_4718 (O_4718,N_49774,N_47647);
or UO_4719 (O_4719,N_48103,N_48173);
or UO_4720 (O_4720,N_48022,N_46693);
nor UO_4721 (O_4721,N_48793,N_46323);
xnor UO_4722 (O_4722,N_47418,N_46165);
and UO_4723 (O_4723,N_49128,N_46660);
xor UO_4724 (O_4724,N_49932,N_48087);
xnor UO_4725 (O_4725,N_45300,N_48092);
xnor UO_4726 (O_4726,N_48636,N_48936);
and UO_4727 (O_4727,N_46406,N_48877);
nand UO_4728 (O_4728,N_47858,N_45718);
or UO_4729 (O_4729,N_45803,N_49455);
or UO_4730 (O_4730,N_48198,N_47706);
nor UO_4731 (O_4731,N_46204,N_47346);
nor UO_4732 (O_4732,N_45141,N_46331);
and UO_4733 (O_4733,N_48762,N_45095);
nor UO_4734 (O_4734,N_45664,N_48056);
xor UO_4735 (O_4735,N_47872,N_45410);
nor UO_4736 (O_4736,N_49495,N_47992);
nor UO_4737 (O_4737,N_49062,N_49748);
nor UO_4738 (O_4738,N_46165,N_47121);
nor UO_4739 (O_4739,N_49129,N_45971);
xnor UO_4740 (O_4740,N_45934,N_48471);
nor UO_4741 (O_4741,N_47671,N_47016);
and UO_4742 (O_4742,N_46262,N_49223);
xor UO_4743 (O_4743,N_48770,N_46147);
and UO_4744 (O_4744,N_47628,N_45498);
and UO_4745 (O_4745,N_47767,N_48531);
or UO_4746 (O_4746,N_48565,N_47184);
or UO_4747 (O_4747,N_47422,N_49071);
and UO_4748 (O_4748,N_48482,N_45236);
xor UO_4749 (O_4749,N_48618,N_45409);
nor UO_4750 (O_4750,N_48633,N_47996);
xor UO_4751 (O_4751,N_48344,N_48079);
or UO_4752 (O_4752,N_49025,N_48553);
and UO_4753 (O_4753,N_49056,N_45693);
nor UO_4754 (O_4754,N_49827,N_49726);
or UO_4755 (O_4755,N_48318,N_45681);
xnor UO_4756 (O_4756,N_49531,N_48663);
nor UO_4757 (O_4757,N_47876,N_46608);
nor UO_4758 (O_4758,N_48955,N_49260);
xor UO_4759 (O_4759,N_46882,N_48810);
nor UO_4760 (O_4760,N_45718,N_47975);
nor UO_4761 (O_4761,N_48359,N_46470);
and UO_4762 (O_4762,N_46985,N_47182);
and UO_4763 (O_4763,N_46468,N_49217);
and UO_4764 (O_4764,N_48800,N_47523);
nor UO_4765 (O_4765,N_46212,N_45787);
nand UO_4766 (O_4766,N_49403,N_49001);
or UO_4767 (O_4767,N_47111,N_47575);
and UO_4768 (O_4768,N_49850,N_49284);
nand UO_4769 (O_4769,N_45854,N_48422);
xor UO_4770 (O_4770,N_45988,N_47707);
xor UO_4771 (O_4771,N_46030,N_47278);
nand UO_4772 (O_4772,N_48781,N_47932);
xnor UO_4773 (O_4773,N_46873,N_46931);
and UO_4774 (O_4774,N_46181,N_47297);
nor UO_4775 (O_4775,N_45986,N_48487);
xnor UO_4776 (O_4776,N_46732,N_46331);
or UO_4777 (O_4777,N_48856,N_47239);
nand UO_4778 (O_4778,N_45863,N_49933);
or UO_4779 (O_4779,N_45654,N_48281);
and UO_4780 (O_4780,N_45566,N_46304);
nor UO_4781 (O_4781,N_48050,N_47244);
nand UO_4782 (O_4782,N_49818,N_49697);
xnor UO_4783 (O_4783,N_49574,N_49737);
or UO_4784 (O_4784,N_49966,N_45158);
nand UO_4785 (O_4785,N_47561,N_45937);
xor UO_4786 (O_4786,N_47757,N_49793);
or UO_4787 (O_4787,N_49597,N_47967);
nand UO_4788 (O_4788,N_49713,N_47507);
or UO_4789 (O_4789,N_45168,N_46813);
or UO_4790 (O_4790,N_49031,N_47965);
xor UO_4791 (O_4791,N_47939,N_47593);
xnor UO_4792 (O_4792,N_45545,N_46349);
or UO_4793 (O_4793,N_46259,N_47785);
or UO_4794 (O_4794,N_46552,N_47582);
and UO_4795 (O_4795,N_49624,N_46108);
xnor UO_4796 (O_4796,N_45932,N_48890);
nand UO_4797 (O_4797,N_48800,N_46832);
and UO_4798 (O_4798,N_45690,N_46832);
xor UO_4799 (O_4799,N_46222,N_47073);
xor UO_4800 (O_4800,N_46408,N_48225);
xor UO_4801 (O_4801,N_48610,N_49699);
nor UO_4802 (O_4802,N_49867,N_45236);
and UO_4803 (O_4803,N_47497,N_45725);
nor UO_4804 (O_4804,N_48282,N_47997);
or UO_4805 (O_4805,N_45710,N_45883);
nand UO_4806 (O_4806,N_48918,N_46529);
and UO_4807 (O_4807,N_45298,N_46151);
and UO_4808 (O_4808,N_47947,N_47101);
xnor UO_4809 (O_4809,N_48978,N_46918);
and UO_4810 (O_4810,N_48427,N_49222);
and UO_4811 (O_4811,N_45909,N_49592);
nor UO_4812 (O_4812,N_45548,N_49171);
xor UO_4813 (O_4813,N_49675,N_49568);
or UO_4814 (O_4814,N_45833,N_46996);
nor UO_4815 (O_4815,N_45027,N_47730);
xnor UO_4816 (O_4816,N_48047,N_49841);
nand UO_4817 (O_4817,N_45105,N_49935);
nor UO_4818 (O_4818,N_48877,N_48684);
nor UO_4819 (O_4819,N_48678,N_46907);
and UO_4820 (O_4820,N_49385,N_47092);
nand UO_4821 (O_4821,N_46379,N_48078);
nand UO_4822 (O_4822,N_47930,N_48299);
or UO_4823 (O_4823,N_45896,N_45983);
and UO_4824 (O_4824,N_46814,N_49293);
nor UO_4825 (O_4825,N_47954,N_48770);
xor UO_4826 (O_4826,N_47222,N_45429);
xnor UO_4827 (O_4827,N_47375,N_47942);
nor UO_4828 (O_4828,N_45178,N_46770);
xor UO_4829 (O_4829,N_46619,N_47431);
nor UO_4830 (O_4830,N_46387,N_47021);
nand UO_4831 (O_4831,N_48995,N_47823);
nor UO_4832 (O_4832,N_47508,N_46649);
nand UO_4833 (O_4833,N_45350,N_45712);
or UO_4834 (O_4834,N_46318,N_45805);
or UO_4835 (O_4835,N_46725,N_48440);
nand UO_4836 (O_4836,N_49235,N_49723);
or UO_4837 (O_4837,N_48733,N_46247);
nand UO_4838 (O_4838,N_46383,N_49145);
or UO_4839 (O_4839,N_49901,N_48499);
xnor UO_4840 (O_4840,N_49962,N_48934);
xor UO_4841 (O_4841,N_47539,N_49886);
nor UO_4842 (O_4842,N_46961,N_46712);
nor UO_4843 (O_4843,N_48617,N_49450);
nand UO_4844 (O_4844,N_45403,N_48912);
and UO_4845 (O_4845,N_48758,N_46378);
xor UO_4846 (O_4846,N_48666,N_46610);
nand UO_4847 (O_4847,N_45870,N_45997);
or UO_4848 (O_4848,N_48378,N_49742);
nor UO_4849 (O_4849,N_48480,N_48886);
and UO_4850 (O_4850,N_45280,N_47131);
and UO_4851 (O_4851,N_48939,N_48403);
nor UO_4852 (O_4852,N_45791,N_48775);
nand UO_4853 (O_4853,N_47802,N_48079);
and UO_4854 (O_4854,N_49056,N_45294);
nor UO_4855 (O_4855,N_45075,N_47311);
xor UO_4856 (O_4856,N_49380,N_48863);
and UO_4857 (O_4857,N_48206,N_47147);
and UO_4858 (O_4858,N_47181,N_49106);
nor UO_4859 (O_4859,N_45572,N_46205);
and UO_4860 (O_4860,N_47723,N_47068);
and UO_4861 (O_4861,N_48672,N_46187);
xnor UO_4862 (O_4862,N_47665,N_46453);
nor UO_4863 (O_4863,N_49522,N_48277);
and UO_4864 (O_4864,N_48524,N_46228);
or UO_4865 (O_4865,N_48163,N_47695);
nor UO_4866 (O_4866,N_47827,N_47198);
and UO_4867 (O_4867,N_46729,N_48665);
and UO_4868 (O_4868,N_47977,N_45586);
xnor UO_4869 (O_4869,N_47752,N_46698);
nand UO_4870 (O_4870,N_46570,N_48680);
and UO_4871 (O_4871,N_48145,N_45324);
and UO_4872 (O_4872,N_49654,N_49777);
nor UO_4873 (O_4873,N_46817,N_48467);
nand UO_4874 (O_4874,N_49421,N_46620);
and UO_4875 (O_4875,N_47197,N_46669);
xnor UO_4876 (O_4876,N_45006,N_45722);
nor UO_4877 (O_4877,N_46452,N_47309);
xor UO_4878 (O_4878,N_49884,N_47462);
xnor UO_4879 (O_4879,N_47455,N_49134);
nor UO_4880 (O_4880,N_46016,N_45116);
or UO_4881 (O_4881,N_45501,N_47352);
nand UO_4882 (O_4882,N_48902,N_46891);
nand UO_4883 (O_4883,N_45833,N_46154);
or UO_4884 (O_4884,N_48286,N_46416);
xor UO_4885 (O_4885,N_48777,N_47140);
and UO_4886 (O_4886,N_47872,N_46525);
nor UO_4887 (O_4887,N_48312,N_45348);
and UO_4888 (O_4888,N_47753,N_48545);
and UO_4889 (O_4889,N_45782,N_45286);
nand UO_4890 (O_4890,N_46231,N_45503);
nor UO_4891 (O_4891,N_47026,N_45294);
and UO_4892 (O_4892,N_49226,N_45101);
and UO_4893 (O_4893,N_46336,N_45437);
nor UO_4894 (O_4894,N_46099,N_49002);
or UO_4895 (O_4895,N_48110,N_45855);
xnor UO_4896 (O_4896,N_47927,N_46689);
nand UO_4897 (O_4897,N_48363,N_47011);
nand UO_4898 (O_4898,N_49938,N_48716);
or UO_4899 (O_4899,N_49173,N_45011);
nand UO_4900 (O_4900,N_47740,N_46740);
or UO_4901 (O_4901,N_46486,N_48669);
or UO_4902 (O_4902,N_45969,N_47340);
xnor UO_4903 (O_4903,N_47144,N_45496);
nand UO_4904 (O_4904,N_45334,N_47666);
and UO_4905 (O_4905,N_49914,N_48501);
or UO_4906 (O_4906,N_46091,N_46086);
or UO_4907 (O_4907,N_45842,N_47091);
and UO_4908 (O_4908,N_48929,N_47812);
xnor UO_4909 (O_4909,N_48629,N_46998);
and UO_4910 (O_4910,N_46259,N_47664);
xor UO_4911 (O_4911,N_45537,N_47344);
or UO_4912 (O_4912,N_45578,N_49934);
xnor UO_4913 (O_4913,N_45492,N_45938);
nand UO_4914 (O_4914,N_49399,N_48156);
and UO_4915 (O_4915,N_47591,N_49587);
nand UO_4916 (O_4916,N_47706,N_47340);
xor UO_4917 (O_4917,N_48804,N_47581);
or UO_4918 (O_4918,N_48584,N_49342);
and UO_4919 (O_4919,N_49188,N_47828);
and UO_4920 (O_4920,N_46526,N_49680);
or UO_4921 (O_4921,N_45254,N_48717);
nand UO_4922 (O_4922,N_49415,N_46626);
or UO_4923 (O_4923,N_45101,N_49530);
and UO_4924 (O_4924,N_48209,N_46729);
nor UO_4925 (O_4925,N_48891,N_48803);
xor UO_4926 (O_4926,N_45183,N_46234);
xor UO_4927 (O_4927,N_48085,N_49124);
nand UO_4928 (O_4928,N_47769,N_46543);
and UO_4929 (O_4929,N_45765,N_48854);
or UO_4930 (O_4930,N_48595,N_48710);
and UO_4931 (O_4931,N_49989,N_47088);
nor UO_4932 (O_4932,N_45451,N_47296);
nand UO_4933 (O_4933,N_49111,N_49998);
or UO_4934 (O_4934,N_45710,N_45558);
nand UO_4935 (O_4935,N_47757,N_49345);
and UO_4936 (O_4936,N_46971,N_48786);
or UO_4937 (O_4937,N_48487,N_47355);
and UO_4938 (O_4938,N_46018,N_48478);
xor UO_4939 (O_4939,N_49514,N_48341);
nand UO_4940 (O_4940,N_46594,N_45654);
nand UO_4941 (O_4941,N_47358,N_48712);
xnor UO_4942 (O_4942,N_46318,N_46302);
and UO_4943 (O_4943,N_48001,N_46168);
nand UO_4944 (O_4944,N_48947,N_45461);
and UO_4945 (O_4945,N_46984,N_47950);
xor UO_4946 (O_4946,N_46512,N_48620);
xor UO_4947 (O_4947,N_47692,N_47552);
or UO_4948 (O_4948,N_47630,N_49418);
and UO_4949 (O_4949,N_47317,N_46628);
xor UO_4950 (O_4950,N_49595,N_46619);
nor UO_4951 (O_4951,N_45873,N_48454);
or UO_4952 (O_4952,N_45763,N_47918);
or UO_4953 (O_4953,N_47347,N_45298);
and UO_4954 (O_4954,N_45113,N_48924);
xor UO_4955 (O_4955,N_47052,N_46678);
or UO_4956 (O_4956,N_46609,N_48355);
nand UO_4957 (O_4957,N_49671,N_46321);
nand UO_4958 (O_4958,N_47656,N_46025);
or UO_4959 (O_4959,N_49200,N_48766);
xor UO_4960 (O_4960,N_49134,N_48415);
xnor UO_4961 (O_4961,N_46446,N_47358);
and UO_4962 (O_4962,N_47417,N_48551);
or UO_4963 (O_4963,N_45489,N_49034);
and UO_4964 (O_4964,N_48772,N_49774);
and UO_4965 (O_4965,N_45036,N_46236);
nand UO_4966 (O_4966,N_45369,N_47150);
and UO_4967 (O_4967,N_45896,N_48799);
nand UO_4968 (O_4968,N_48335,N_46411);
nand UO_4969 (O_4969,N_48818,N_47901);
xor UO_4970 (O_4970,N_46351,N_46788);
and UO_4971 (O_4971,N_45587,N_49167);
and UO_4972 (O_4972,N_45272,N_47528);
or UO_4973 (O_4973,N_48954,N_47679);
or UO_4974 (O_4974,N_49339,N_45897);
nand UO_4975 (O_4975,N_46256,N_48904);
or UO_4976 (O_4976,N_48392,N_48264);
nor UO_4977 (O_4977,N_45217,N_45191);
xnor UO_4978 (O_4978,N_46087,N_48905);
xor UO_4979 (O_4979,N_46112,N_49010);
nand UO_4980 (O_4980,N_46814,N_46070);
xor UO_4981 (O_4981,N_47000,N_49821);
nand UO_4982 (O_4982,N_47649,N_45324);
nand UO_4983 (O_4983,N_49279,N_48735);
nand UO_4984 (O_4984,N_45768,N_48190);
nor UO_4985 (O_4985,N_49537,N_49212);
nor UO_4986 (O_4986,N_48262,N_46609);
nor UO_4987 (O_4987,N_45786,N_47611);
or UO_4988 (O_4988,N_45706,N_45611);
nor UO_4989 (O_4989,N_49828,N_47202);
and UO_4990 (O_4990,N_47695,N_47048);
nor UO_4991 (O_4991,N_47955,N_46242);
or UO_4992 (O_4992,N_49956,N_49086);
or UO_4993 (O_4993,N_45008,N_46143);
xor UO_4994 (O_4994,N_46622,N_49311);
nand UO_4995 (O_4995,N_48384,N_49630);
or UO_4996 (O_4996,N_45868,N_48893);
nand UO_4997 (O_4997,N_48129,N_45059);
nor UO_4998 (O_4998,N_45000,N_48824);
nand UO_4999 (O_4999,N_47640,N_46315);
endmodule