module basic_500_3000_500_60_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_227,In_464);
and U1 (N_1,In_340,In_269);
or U2 (N_2,In_249,In_73);
nand U3 (N_3,In_468,In_476);
xnor U4 (N_4,In_481,In_297);
xnor U5 (N_5,In_32,In_341);
or U6 (N_6,In_343,In_187);
or U7 (N_7,In_172,In_237);
xnor U8 (N_8,In_432,In_117);
nor U9 (N_9,In_107,In_189);
xnor U10 (N_10,In_1,In_61);
nand U11 (N_11,In_7,In_329);
nand U12 (N_12,In_273,In_431);
nand U13 (N_13,In_317,In_39);
nor U14 (N_14,In_424,In_434);
nand U15 (N_15,In_302,In_219);
nand U16 (N_16,In_89,In_496);
nand U17 (N_17,In_473,In_131);
or U18 (N_18,In_147,In_201);
xor U19 (N_19,In_351,In_370);
and U20 (N_20,In_484,In_177);
xor U21 (N_21,In_103,In_488);
nand U22 (N_22,In_45,In_453);
xor U23 (N_23,In_272,In_410);
nor U24 (N_24,In_335,In_72);
nand U25 (N_25,In_190,In_119);
nand U26 (N_26,In_369,In_316);
nand U27 (N_27,In_358,In_67);
or U28 (N_28,In_394,In_19);
nor U29 (N_29,In_135,In_71);
nor U30 (N_30,In_252,In_31);
nand U31 (N_31,In_479,In_170);
and U32 (N_32,In_212,In_356);
nand U33 (N_33,In_198,In_74);
xor U34 (N_34,In_386,In_223);
xnor U35 (N_35,In_346,In_142);
or U36 (N_36,In_195,In_373);
nor U37 (N_37,In_357,In_466);
nor U38 (N_38,In_165,In_287);
nand U39 (N_39,In_129,In_311);
or U40 (N_40,In_152,In_455);
or U41 (N_41,In_469,In_192);
xor U42 (N_42,In_91,In_193);
and U43 (N_43,In_310,In_41);
and U44 (N_44,In_79,In_99);
or U45 (N_45,In_263,In_78);
or U46 (N_46,In_120,In_321);
xnor U47 (N_47,In_282,In_22);
xnor U48 (N_48,In_459,In_150);
nor U49 (N_49,In_445,In_401);
and U50 (N_50,In_236,N_0);
or U51 (N_51,In_8,In_105);
or U52 (N_52,In_332,In_456);
xor U53 (N_53,In_485,In_218);
xor U54 (N_54,N_10,In_243);
xnor U55 (N_55,In_3,N_2);
nor U56 (N_56,In_376,In_256);
and U57 (N_57,In_324,In_377);
nand U58 (N_58,In_204,In_141);
nand U59 (N_59,In_380,In_301);
nand U60 (N_60,In_208,In_126);
nor U61 (N_61,In_76,In_450);
nor U62 (N_62,In_314,In_436);
and U63 (N_63,In_393,In_233);
xnor U64 (N_64,In_54,N_8);
nor U65 (N_65,In_56,In_253);
nand U66 (N_66,In_345,In_104);
and U67 (N_67,In_344,N_11);
xor U68 (N_68,In_100,In_55);
or U69 (N_69,In_77,In_10);
or U70 (N_70,N_7,In_114);
nand U71 (N_71,In_309,In_88);
and U72 (N_72,In_378,N_41);
nand U73 (N_73,In_173,In_110);
or U74 (N_74,In_137,In_251);
nand U75 (N_75,In_97,In_262);
nor U76 (N_76,In_283,In_98);
xnor U77 (N_77,In_144,N_12);
and U78 (N_78,In_199,In_155);
xnor U79 (N_79,In_229,In_48);
nand U80 (N_80,In_388,In_421);
and U81 (N_81,In_15,In_228);
or U82 (N_82,In_460,In_214);
and U83 (N_83,In_402,N_44);
or U84 (N_84,N_35,In_339);
or U85 (N_85,In_37,In_419);
and U86 (N_86,In_348,In_109);
or U87 (N_87,N_31,In_169);
or U88 (N_88,In_175,In_405);
or U89 (N_89,In_379,In_69);
nand U90 (N_90,N_13,In_247);
and U91 (N_91,In_44,In_323);
or U92 (N_92,In_146,In_18);
and U93 (N_93,In_461,In_57);
and U94 (N_94,N_30,In_163);
nor U95 (N_95,In_497,In_66);
and U96 (N_96,In_200,In_25);
and U97 (N_97,In_290,In_420);
and U98 (N_98,In_304,In_327);
xor U99 (N_99,In_52,In_463);
xor U100 (N_100,N_93,In_413);
nand U101 (N_101,N_79,In_211);
or U102 (N_102,N_22,N_34);
or U103 (N_103,In_210,N_32);
and U104 (N_104,N_74,N_46);
xnor U105 (N_105,In_408,N_73);
and U106 (N_106,In_398,In_145);
nand U107 (N_107,In_296,N_82);
xor U108 (N_108,In_470,In_441);
nor U109 (N_109,N_63,In_132);
nand U110 (N_110,In_385,In_375);
nand U111 (N_111,In_58,In_448);
or U112 (N_112,In_166,In_43);
and U113 (N_113,In_221,In_184);
nor U114 (N_114,In_121,In_149);
nor U115 (N_115,In_289,In_34);
nor U116 (N_116,In_112,In_280);
nand U117 (N_117,In_399,In_430);
nand U118 (N_118,In_92,In_384);
nand U119 (N_119,In_482,In_371);
and U120 (N_120,In_276,In_230);
nor U121 (N_121,In_232,In_42);
nor U122 (N_122,In_465,N_16);
xnor U123 (N_123,In_372,N_48);
and U124 (N_124,N_83,In_235);
and U125 (N_125,In_266,In_197);
or U126 (N_126,In_425,In_486);
nor U127 (N_127,N_5,In_106);
nand U128 (N_128,In_29,In_300);
and U129 (N_129,In_354,In_418);
nand U130 (N_130,In_457,N_71);
nand U131 (N_131,In_478,N_4);
or U132 (N_132,In_33,N_9);
and U133 (N_133,In_298,N_94);
nor U134 (N_134,In_40,In_206);
nor U135 (N_135,In_319,In_492);
nand U136 (N_136,N_29,In_254);
or U137 (N_137,In_244,In_387);
or U138 (N_138,In_284,In_6);
or U139 (N_139,In_279,In_242);
or U140 (N_140,In_427,In_390);
xnor U141 (N_141,In_275,N_59);
nand U142 (N_142,In_494,N_40);
or U143 (N_143,In_240,N_49);
nand U144 (N_144,In_239,In_179);
or U145 (N_145,In_412,In_397);
nor U146 (N_146,In_265,In_108);
or U147 (N_147,N_37,N_25);
nor U148 (N_148,In_5,N_70);
nand U149 (N_149,In_21,In_326);
nor U150 (N_150,In_196,In_23);
and U151 (N_151,In_151,In_125);
nand U152 (N_152,In_9,N_137);
xor U153 (N_153,In_264,In_366);
xnor U154 (N_154,In_245,In_382);
or U155 (N_155,N_15,In_30);
or U156 (N_156,N_105,In_130);
or U157 (N_157,In_17,In_451);
or U158 (N_158,In_168,N_50);
and U159 (N_159,In_157,In_27);
nor U160 (N_160,In_20,N_24);
nand U161 (N_161,In_118,In_171);
and U162 (N_162,N_88,N_122);
nand U163 (N_163,In_160,In_320);
or U164 (N_164,N_139,In_299);
and U165 (N_165,In_499,In_83);
nand U166 (N_166,N_19,In_191);
xor U167 (N_167,In_94,In_24);
and U168 (N_168,N_57,N_61);
xnor U169 (N_169,N_127,N_23);
nand U170 (N_170,In_267,In_400);
xnor U171 (N_171,N_101,In_116);
and U172 (N_172,In_225,N_81);
and U173 (N_173,In_102,In_475);
nand U174 (N_174,In_355,In_293);
nor U175 (N_175,N_26,In_101);
nor U176 (N_176,N_146,In_261);
xnor U177 (N_177,N_135,In_277);
or U178 (N_178,N_20,N_130);
xor U179 (N_179,N_132,In_209);
xnor U180 (N_180,N_56,N_142);
nand U181 (N_181,In_14,In_70);
nor U182 (N_182,N_1,In_93);
or U183 (N_183,In_491,In_447);
nand U184 (N_184,In_174,N_77);
xor U185 (N_185,In_95,In_429);
nand U186 (N_186,In_50,N_147);
xor U187 (N_187,N_113,In_161);
and U188 (N_188,N_67,N_18);
nor U189 (N_189,In_85,N_100);
xnor U190 (N_190,In_426,N_104);
xnor U191 (N_191,In_328,In_86);
xor U192 (N_192,In_438,In_474);
nand U193 (N_193,In_493,N_117);
and U194 (N_194,In_442,In_220);
nor U195 (N_195,In_315,N_17);
xor U196 (N_196,In_333,N_68);
and U197 (N_197,N_133,In_477);
and U198 (N_198,In_207,N_90);
nor U199 (N_199,In_128,N_114);
xor U200 (N_200,N_47,In_359);
nand U201 (N_201,In_194,In_483);
and U202 (N_202,In_367,In_183);
nand U203 (N_203,In_417,In_64);
nand U204 (N_204,N_178,In_433);
or U205 (N_205,In_96,N_162);
or U206 (N_206,In_202,N_196);
nor U207 (N_207,N_3,N_165);
nor U208 (N_208,In_188,N_95);
nor U209 (N_209,In_423,In_164);
and U210 (N_210,In_439,In_203);
or U211 (N_211,N_150,In_12);
xor U212 (N_212,In_285,N_144);
and U213 (N_213,In_458,N_38);
nand U214 (N_214,N_155,N_119);
nand U215 (N_215,In_241,N_140);
or U216 (N_216,In_381,In_353);
nand U217 (N_217,N_187,N_42);
and U218 (N_218,In_337,In_480);
and U219 (N_219,N_180,In_305);
nand U220 (N_220,In_124,In_489);
xnor U221 (N_221,N_84,In_122);
and U222 (N_222,N_151,N_103);
nand U223 (N_223,N_163,N_28);
nor U224 (N_224,N_118,In_313);
nor U225 (N_225,N_96,In_374);
nand U226 (N_226,In_139,In_409);
or U227 (N_227,In_404,In_49);
and U228 (N_228,In_234,In_271);
xnor U229 (N_229,In_250,N_183);
nor U230 (N_230,In_389,In_140);
xor U231 (N_231,N_169,N_195);
xnor U232 (N_232,In_338,In_274);
nand U233 (N_233,In_449,In_361);
and U234 (N_234,N_62,In_154);
nor U235 (N_235,In_156,N_154);
xor U236 (N_236,N_106,N_138);
nand U237 (N_237,N_21,N_190);
and U238 (N_238,N_55,In_87);
xor U239 (N_239,In_306,N_168);
and U240 (N_240,In_16,In_454);
nand U241 (N_241,In_281,In_325);
xnor U242 (N_242,In_467,N_161);
nor U243 (N_243,N_173,In_216);
nand U244 (N_244,N_98,N_171);
nor U245 (N_245,N_136,In_428);
nor U246 (N_246,N_92,In_226);
or U247 (N_247,In_115,N_182);
xor U248 (N_248,In_294,In_278);
nor U249 (N_249,In_143,In_472);
or U250 (N_250,N_158,In_176);
nor U251 (N_251,N_87,In_490);
and U252 (N_252,N_160,In_349);
nor U253 (N_253,N_86,In_47);
xnor U254 (N_254,In_403,In_258);
or U255 (N_255,N_231,In_2);
nor U256 (N_256,In_352,In_414);
nor U257 (N_257,N_206,N_244);
nand U258 (N_258,In_416,In_217);
nor U259 (N_259,N_128,N_110);
xor U260 (N_260,N_198,In_334);
nand U261 (N_261,In_336,In_134);
or U262 (N_262,In_80,In_396);
or U263 (N_263,In_260,N_123);
xnor U264 (N_264,In_471,N_134);
nand U265 (N_265,In_362,N_45);
nor U266 (N_266,N_143,N_43);
xor U267 (N_267,In_11,N_184);
xor U268 (N_268,N_202,N_188);
or U269 (N_269,In_65,In_452);
nand U270 (N_270,In_365,N_243);
or U271 (N_271,In_215,In_238);
nand U272 (N_272,N_215,In_178);
nor U273 (N_273,In_368,N_97);
xnor U274 (N_274,In_46,In_81);
or U275 (N_275,In_422,N_217);
or U276 (N_276,In_347,N_52);
and U277 (N_277,N_192,N_66);
nand U278 (N_278,N_248,N_239);
or U279 (N_279,N_39,N_116);
nand U280 (N_280,In_444,In_38);
or U281 (N_281,In_342,In_136);
nand U282 (N_282,In_406,N_112);
nor U283 (N_283,N_60,N_177);
and U284 (N_284,In_392,N_236);
or U285 (N_285,N_69,N_233);
xor U286 (N_286,N_108,N_148);
nand U287 (N_287,In_288,In_123);
nand U288 (N_288,N_27,In_181);
xor U289 (N_289,In_213,In_383);
nand U290 (N_290,In_360,In_322);
and U291 (N_291,In_59,In_53);
nor U292 (N_292,N_65,N_54);
and U293 (N_293,N_102,N_99);
nand U294 (N_294,N_246,N_193);
xnor U295 (N_295,N_53,In_443);
nand U296 (N_296,In_82,In_270);
or U297 (N_297,In_111,N_238);
and U298 (N_298,In_248,N_72);
xnor U299 (N_299,N_172,In_28);
nor U300 (N_300,N_295,N_181);
and U301 (N_301,N_252,In_90);
nand U302 (N_302,In_487,In_63);
nand U303 (N_303,N_175,N_91);
and U304 (N_304,In_159,N_167);
nor U305 (N_305,N_290,In_440);
nor U306 (N_306,N_284,In_498);
nand U307 (N_307,N_152,N_264);
nor U308 (N_308,N_299,In_162);
or U309 (N_309,N_296,N_120);
and U310 (N_310,N_205,N_145);
nand U311 (N_311,In_437,In_231);
and U312 (N_312,N_121,In_167);
nand U313 (N_313,In_312,In_51);
and U314 (N_314,N_224,N_203);
nor U315 (N_315,N_292,In_286);
and U316 (N_316,N_166,N_251);
and U317 (N_317,In_331,N_149);
nand U318 (N_318,N_221,N_269);
nand U319 (N_319,N_237,N_232);
or U320 (N_320,N_170,N_211);
or U321 (N_321,In_158,N_220);
xnor U322 (N_322,In_182,In_257);
nand U323 (N_323,In_318,N_225);
and U324 (N_324,In_36,In_435);
and U325 (N_325,In_133,N_191);
or U326 (N_326,N_254,N_194);
or U327 (N_327,In_268,In_415);
nor U328 (N_328,N_58,N_208);
xnor U329 (N_329,N_261,N_156);
nor U330 (N_330,N_241,N_291);
nand U331 (N_331,N_286,N_275);
nor U332 (N_332,N_107,N_288);
and U333 (N_333,N_285,N_271);
xor U334 (N_334,N_234,N_283);
nand U335 (N_335,In_495,N_210);
nor U336 (N_336,N_214,N_125);
or U337 (N_337,N_204,N_6);
or U338 (N_338,N_247,In_4);
nor U339 (N_339,N_115,In_303);
xor U340 (N_340,N_111,In_60);
and U341 (N_341,N_282,In_259);
xnor U342 (N_342,In_180,In_0);
nand U343 (N_343,N_229,In_407);
and U344 (N_344,N_228,N_64);
xnor U345 (N_345,N_174,N_222);
and U346 (N_346,N_219,N_297);
xnor U347 (N_347,N_131,In_148);
nor U348 (N_348,N_227,In_186);
nor U349 (N_349,N_263,In_138);
and U350 (N_350,N_272,N_319);
and U351 (N_351,N_209,In_84);
xnor U352 (N_352,In_113,N_256);
or U353 (N_353,N_164,N_320);
xnor U354 (N_354,N_250,In_295);
and U355 (N_355,N_331,N_262);
nor U356 (N_356,N_197,N_141);
nand U357 (N_357,N_325,N_347);
and U358 (N_358,N_280,N_344);
or U359 (N_359,N_277,N_345);
nor U360 (N_360,N_268,N_294);
and U361 (N_361,N_333,N_318);
and U362 (N_362,N_329,N_226);
and U363 (N_363,N_157,N_341);
nand U364 (N_364,N_179,N_85);
xor U365 (N_365,In_26,In_222);
and U366 (N_366,N_189,N_335);
nand U367 (N_367,N_300,N_330);
and U368 (N_368,N_304,N_230);
nand U369 (N_369,N_328,N_274);
and U370 (N_370,N_124,N_185);
nand U371 (N_371,In_411,N_259);
and U372 (N_372,In_255,N_337);
xor U373 (N_373,In_75,N_270);
nor U374 (N_374,N_317,In_13);
and U375 (N_375,N_33,N_235);
nand U376 (N_376,N_324,In_35);
xnor U377 (N_377,N_334,N_312);
and U378 (N_378,N_258,N_311);
nor U379 (N_379,In_462,N_308);
and U380 (N_380,N_323,N_159);
nor U381 (N_381,N_200,N_260);
nand U382 (N_382,N_109,N_279);
xor U383 (N_383,N_199,N_276);
xor U384 (N_384,N_293,N_349);
nor U385 (N_385,N_186,N_336);
nand U386 (N_386,N_287,N_242);
and U387 (N_387,N_322,N_89);
and U388 (N_388,N_339,N_313);
xnor U389 (N_389,N_218,N_281);
or U390 (N_390,N_267,N_51);
nor U391 (N_391,N_343,N_255);
and U392 (N_392,In_185,N_305);
or U393 (N_393,In_291,In_62);
xor U394 (N_394,N_36,N_176);
nor U395 (N_395,N_223,In_446);
nor U396 (N_396,N_307,N_212);
or U397 (N_397,N_207,N_273);
or U398 (N_398,N_126,N_80);
xnor U399 (N_399,N_129,N_75);
xnor U400 (N_400,N_321,N_391);
nand U401 (N_401,N_14,In_205);
and U402 (N_402,N_380,N_358);
nor U403 (N_403,In_330,N_378);
xnor U404 (N_404,N_309,N_364);
and U405 (N_405,N_306,N_342);
nor U406 (N_406,N_384,N_377);
nand U407 (N_407,In_153,In_364);
or U408 (N_408,N_370,N_348);
nor U409 (N_409,N_351,N_369);
nor U410 (N_410,N_302,In_292);
nor U411 (N_411,N_346,N_315);
nand U412 (N_412,N_249,N_368);
xor U413 (N_413,N_216,N_392);
nand U414 (N_414,N_356,N_397);
nor U415 (N_415,N_396,In_68);
and U416 (N_416,N_386,N_303);
nand U417 (N_417,N_298,In_395);
or U418 (N_418,N_240,N_265);
nor U419 (N_419,N_393,N_398);
nand U420 (N_420,In_127,N_213);
nand U421 (N_421,N_314,N_301);
xnor U422 (N_422,N_245,N_363);
and U423 (N_423,In_224,N_257);
nor U424 (N_424,N_367,N_371);
and U425 (N_425,N_360,N_373);
and U426 (N_426,N_153,N_350);
xnor U427 (N_427,N_399,N_310);
nor U428 (N_428,N_365,N_394);
or U429 (N_429,N_332,N_78);
nand U430 (N_430,N_266,N_326);
xnor U431 (N_431,N_379,N_382);
nand U432 (N_432,N_362,N_338);
xor U433 (N_433,N_387,N_76);
nand U434 (N_434,In_307,N_327);
nor U435 (N_435,N_385,N_372);
xor U436 (N_436,N_381,In_308);
or U437 (N_437,In_246,N_357);
or U438 (N_438,N_366,N_354);
and U439 (N_439,N_390,N_355);
nor U440 (N_440,N_375,N_253);
or U441 (N_441,N_352,In_391);
nor U442 (N_442,N_376,N_359);
nand U443 (N_443,N_316,N_374);
nor U444 (N_444,N_201,N_383);
nor U445 (N_445,N_361,N_278);
or U446 (N_446,N_289,N_395);
xnor U447 (N_447,N_340,N_388);
and U448 (N_448,N_353,N_389);
nand U449 (N_449,In_363,In_350);
nor U450 (N_450,N_403,N_430);
and U451 (N_451,N_429,N_433);
or U452 (N_452,N_404,N_411);
nand U453 (N_453,N_443,N_440);
and U454 (N_454,N_436,N_410);
nand U455 (N_455,N_423,N_437);
nor U456 (N_456,N_426,N_427);
nand U457 (N_457,N_420,N_405);
or U458 (N_458,N_432,N_449);
nor U459 (N_459,N_418,N_448);
and U460 (N_460,N_442,N_413);
or U461 (N_461,N_445,N_422);
nor U462 (N_462,N_446,N_407);
nand U463 (N_463,N_417,N_447);
nor U464 (N_464,N_425,N_439);
xnor U465 (N_465,N_415,N_406);
or U466 (N_466,N_431,N_400);
or U467 (N_467,N_435,N_412);
nand U468 (N_468,N_409,N_424);
nor U469 (N_469,N_408,N_438);
xor U470 (N_470,N_401,N_444);
and U471 (N_471,N_421,N_419);
and U472 (N_472,N_416,N_414);
xor U473 (N_473,N_428,N_441);
and U474 (N_474,N_402,N_434);
or U475 (N_475,N_443,N_446);
xor U476 (N_476,N_413,N_424);
and U477 (N_477,N_413,N_400);
nand U478 (N_478,N_445,N_411);
or U479 (N_479,N_425,N_409);
xor U480 (N_480,N_443,N_439);
or U481 (N_481,N_415,N_445);
and U482 (N_482,N_427,N_420);
or U483 (N_483,N_440,N_416);
and U484 (N_484,N_443,N_408);
xor U485 (N_485,N_442,N_444);
nand U486 (N_486,N_402,N_436);
nor U487 (N_487,N_418,N_411);
xnor U488 (N_488,N_414,N_431);
or U489 (N_489,N_439,N_414);
and U490 (N_490,N_412,N_431);
and U491 (N_491,N_444,N_405);
xor U492 (N_492,N_446,N_413);
and U493 (N_493,N_420,N_410);
xor U494 (N_494,N_440,N_429);
nor U495 (N_495,N_423,N_421);
xnor U496 (N_496,N_411,N_436);
nor U497 (N_497,N_414,N_405);
nor U498 (N_498,N_409,N_417);
and U499 (N_499,N_412,N_423);
nor U500 (N_500,N_453,N_456);
xnor U501 (N_501,N_459,N_460);
nor U502 (N_502,N_482,N_457);
or U503 (N_503,N_450,N_452);
and U504 (N_504,N_465,N_488);
and U505 (N_505,N_487,N_455);
nand U506 (N_506,N_499,N_492);
and U507 (N_507,N_469,N_498);
or U508 (N_508,N_467,N_473);
xor U509 (N_509,N_496,N_484);
or U510 (N_510,N_494,N_470);
or U511 (N_511,N_451,N_485);
nand U512 (N_512,N_478,N_497);
xor U513 (N_513,N_486,N_491);
xor U514 (N_514,N_468,N_493);
nor U515 (N_515,N_489,N_479);
or U516 (N_516,N_472,N_474);
xor U517 (N_517,N_481,N_475);
and U518 (N_518,N_464,N_458);
and U519 (N_519,N_490,N_471);
xnor U520 (N_520,N_477,N_462);
or U521 (N_521,N_476,N_480);
xor U522 (N_522,N_463,N_466);
xor U523 (N_523,N_495,N_454);
xor U524 (N_524,N_483,N_461);
and U525 (N_525,N_465,N_472);
and U526 (N_526,N_460,N_463);
or U527 (N_527,N_471,N_480);
nor U528 (N_528,N_486,N_482);
nand U529 (N_529,N_498,N_473);
and U530 (N_530,N_455,N_490);
or U531 (N_531,N_456,N_474);
nor U532 (N_532,N_471,N_466);
nand U533 (N_533,N_488,N_476);
or U534 (N_534,N_455,N_476);
nor U535 (N_535,N_472,N_492);
nor U536 (N_536,N_483,N_480);
nand U537 (N_537,N_491,N_496);
xor U538 (N_538,N_467,N_484);
and U539 (N_539,N_493,N_475);
and U540 (N_540,N_452,N_460);
or U541 (N_541,N_453,N_472);
nor U542 (N_542,N_486,N_464);
nand U543 (N_543,N_490,N_485);
nand U544 (N_544,N_488,N_468);
nand U545 (N_545,N_451,N_476);
nand U546 (N_546,N_450,N_492);
nor U547 (N_547,N_480,N_458);
xnor U548 (N_548,N_496,N_475);
nand U549 (N_549,N_488,N_450);
nor U550 (N_550,N_532,N_537);
nor U551 (N_551,N_534,N_515);
nand U552 (N_552,N_542,N_522);
nor U553 (N_553,N_510,N_546);
nand U554 (N_554,N_511,N_526);
xor U555 (N_555,N_548,N_521);
and U556 (N_556,N_536,N_503);
or U557 (N_557,N_508,N_549);
or U558 (N_558,N_518,N_504);
nor U559 (N_559,N_525,N_540);
xnor U560 (N_560,N_516,N_528);
and U561 (N_561,N_543,N_533);
xor U562 (N_562,N_517,N_529);
nand U563 (N_563,N_507,N_547);
nor U564 (N_564,N_524,N_506);
and U565 (N_565,N_513,N_501);
and U566 (N_566,N_530,N_509);
xnor U567 (N_567,N_514,N_512);
xnor U568 (N_568,N_541,N_523);
nor U569 (N_569,N_519,N_505);
or U570 (N_570,N_538,N_531);
and U571 (N_571,N_502,N_535);
xor U572 (N_572,N_539,N_500);
and U573 (N_573,N_520,N_527);
nand U574 (N_574,N_545,N_544);
and U575 (N_575,N_501,N_505);
or U576 (N_576,N_517,N_504);
nor U577 (N_577,N_527,N_504);
nand U578 (N_578,N_548,N_532);
or U579 (N_579,N_523,N_518);
nor U580 (N_580,N_537,N_508);
and U581 (N_581,N_507,N_511);
nor U582 (N_582,N_504,N_515);
nand U583 (N_583,N_537,N_538);
or U584 (N_584,N_535,N_546);
or U585 (N_585,N_510,N_502);
xnor U586 (N_586,N_510,N_548);
nor U587 (N_587,N_523,N_514);
xnor U588 (N_588,N_513,N_528);
and U589 (N_589,N_534,N_519);
and U590 (N_590,N_549,N_546);
and U591 (N_591,N_518,N_529);
and U592 (N_592,N_535,N_505);
xor U593 (N_593,N_528,N_541);
and U594 (N_594,N_508,N_500);
nor U595 (N_595,N_527,N_521);
or U596 (N_596,N_509,N_519);
or U597 (N_597,N_540,N_515);
xnor U598 (N_598,N_549,N_534);
xnor U599 (N_599,N_535,N_510);
nor U600 (N_600,N_551,N_562);
or U601 (N_601,N_560,N_575);
nor U602 (N_602,N_596,N_580);
nor U603 (N_603,N_589,N_559);
nand U604 (N_604,N_568,N_552);
xnor U605 (N_605,N_567,N_592);
and U606 (N_606,N_571,N_555);
nand U607 (N_607,N_565,N_595);
nand U608 (N_608,N_553,N_587);
nand U609 (N_609,N_556,N_597);
or U610 (N_610,N_583,N_572);
nand U611 (N_611,N_585,N_574);
xnor U612 (N_612,N_582,N_576);
or U613 (N_613,N_599,N_593);
or U614 (N_614,N_577,N_570);
or U615 (N_615,N_564,N_579);
xnor U616 (N_616,N_557,N_581);
xor U617 (N_617,N_550,N_591);
nand U618 (N_618,N_594,N_586);
xnor U619 (N_619,N_554,N_563);
and U620 (N_620,N_588,N_561);
xor U621 (N_621,N_566,N_573);
nor U622 (N_622,N_569,N_578);
nand U623 (N_623,N_590,N_598);
and U624 (N_624,N_558,N_584);
nor U625 (N_625,N_596,N_550);
or U626 (N_626,N_562,N_565);
or U627 (N_627,N_566,N_570);
or U628 (N_628,N_576,N_599);
xnor U629 (N_629,N_555,N_553);
xor U630 (N_630,N_579,N_576);
nor U631 (N_631,N_590,N_558);
and U632 (N_632,N_576,N_567);
and U633 (N_633,N_559,N_583);
nand U634 (N_634,N_567,N_587);
or U635 (N_635,N_577,N_596);
nand U636 (N_636,N_559,N_578);
or U637 (N_637,N_571,N_552);
and U638 (N_638,N_583,N_588);
or U639 (N_639,N_593,N_586);
or U640 (N_640,N_565,N_555);
xnor U641 (N_641,N_556,N_566);
and U642 (N_642,N_563,N_598);
nor U643 (N_643,N_567,N_588);
or U644 (N_644,N_556,N_599);
xnor U645 (N_645,N_593,N_563);
nor U646 (N_646,N_554,N_593);
or U647 (N_647,N_556,N_582);
or U648 (N_648,N_590,N_556);
or U649 (N_649,N_581,N_583);
and U650 (N_650,N_613,N_612);
and U651 (N_651,N_629,N_623);
xnor U652 (N_652,N_631,N_639);
or U653 (N_653,N_616,N_647);
xnor U654 (N_654,N_640,N_605);
nand U655 (N_655,N_610,N_648);
or U656 (N_656,N_635,N_630);
or U657 (N_657,N_603,N_606);
nand U658 (N_658,N_607,N_614);
and U659 (N_659,N_644,N_624);
xnor U660 (N_660,N_634,N_646);
or U661 (N_661,N_649,N_611);
and U662 (N_662,N_608,N_621);
nand U663 (N_663,N_632,N_637);
nand U664 (N_664,N_620,N_626);
nor U665 (N_665,N_619,N_645);
xnor U666 (N_666,N_609,N_600);
nor U667 (N_667,N_602,N_627);
nand U668 (N_668,N_642,N_617);
xnor U669 (N_669,N_638,N_601);
or U670 (N_670,N_625,N_615);
nand U671 (N_671,N_633,N_641);
and U672 (N_672,N_604,N_622);
or U673 (N_673,N_628,N_643);
and U674 (N_674,N_618,N_636);
or U675 (N_675,N_619,N_615);
and U676 (N_676,N_642,N_621);
xnor U677 (N_677,N_614,N_635);
nand U678 (N_678,N_614,N_637);
xor U679 (N_679,N_645,N_639);
nor U680 (N_680,N_616,N_629);
nor U681 (N_681,N_648,N_605);
and U682 (N_682,N_618,N_610);
xnor U683 (N_683,N_634,N_610);
xnor U684 (N_684,N_633,N_644);
nor U685 (N_685,N_612,N_609);
xnor U686 (N_686,N_613,N_627);
nor U687 (N_687,N_624,N_612);
xor U688 (N_688,N_600,N_619);
or U689 (N_689,N_617,N_641);
nor U690 (N_690,N_637,N_615);
nor U691 (N_691,N_605,N_646);
nor U692 (N_692,N_634,N_614);
nand U693 (N_693,N_604,N_621);
or U694 (N_694,N_612,N_603);
xnor U695 (N_695,N_608,N_645);
xor U696 (N_696,N_640,N_644);
or U697 (N_697,N_603,N_647);
xnor U698 (N_698,N_611,N_606);
and U699 (N_699,N_621,N_629);
nor U700 (N_700,N_689,N_659);
or U701 (N_701,N_653,N_661);
and U702 (N_702,N_694,N_650);
xor U703 (N_703,N_665,N_696);
nand U704 (N_704,N_697,N_693);
nor U705 (N_705,N_655,N_671);
xor U706 (N_706,N_690,N_674);
nand U707 (N_707,N_652,N_688);
or U708 (N_708,N_666,N_695);
or U709 (N_709,N_685,N_657);
nor U710 (N_710,N_682,N_677);
nor U711 (N_711,N_686,N_678);
or U712 (N_712,N_679,N_663);
nor U713 (N_713,N_656,N_687);
or U714 (N_714,N_664,N_683);
nor U715 (N_715,N_699,N_681);
nand U716 (N_716,N_654,N_691);
xor U717 (N_717,N_662,N_692);
xnor U718 (N_718,N_698,N_673);
nor U719 (N_719,N_667,N_670);
or U720 (N_720,N_672,N_675);
nor U721 (N_721,N_676,N_680);
or U722 (N_722,N_660,N_668);
nand U723 (N_723,N_658,N_669);
or U724 (N_724,N_684,N_651);
xor U725 (N_725,N_681,N_657);
and U726 (N_726,N_676,N_684);
or U727 (N_727,N_652,N_651);
and U728 (N_728,N_698,N_696);
and U729 (N_729,N_685,N_698);
nor U730 (N_730,N_688,N_686);
nor U731 (N_731,N_664,N_654);
or U732 (N_732,N_660,N_692);
xnor U733 (N_733,N_662,N_667);
and U734 (N_734,N_675,N_654);
or U735 (N_735,N_663,N_651);
or U736 (N_736,N_688,N_677);
nor U737 (N_737,N_664,N_659);
xor U738 (N_738,N_684,N_662);
xnor U739 (N_739,N_687,N_683);
and U740 (N_740,N_677,N_673);
nand U741 (N_741,N_676,N_658);
nand U742 (N_742,N_673,N_674);
or U743 (N_743,N_665,N_685);
nand U744 (N_744,N_670,N_699);
nand U745 (N_745,N_672,N_679);
nor U746 (N_746,N_651,N_662);
nand U747 (N_747,N_679,N_657);
and U748 (N_748,N_667,N_652);
nand U749 (N_749,N_690,N_699);
xnor U750 (N_750,N_705,N_706);
and U751 (N_751,N_749,N_703);
nand U752 (N_752,N_700,N_712);
nor U753 (N_753,N_719,N_731);
nand U754 (N_754,N_743,N_735);
xor U755 (N_755,N_707,N_721);
and U756 (N_756,N_715,N_723);
and U757 (N_757,N_720,N_724);
xor U758 (N_758,N_746,N_733);
and U759 (N_759,N_702,N_730);
nand U760 (N_760,N_740,N_734);
and U761 (N_761,N_718,N_741);
nor U762 (N_762,N_710,N_709);
nor U763 (N_763,N_713,N_701);
nor U764 (N_764,N_704,N_716);
nor U765 (N_765,N_717,N_727);
nand U766 (N_766,N_722,N_714);
nand U767 (N_767,N_732,N_747);
xnor U768 (N_768,N_725,N_742);
xnor U769 (N_769,N_737,N_744);
nor U770 (N_770,N_736,N_708);
nand U771 (N_771,N_711,N_739);
nor U772 (N_772,N_729,N_726);
or U773 (N_773,N_748,N_738);
xor U774 (N_774,N_745,N_728);
nor U775 (N_775,N_729,N_721);
xor U776 (N_776,N_726,N_745);
nor U777 (N_777,N_719,N_720);
xor U778 (N_778,N_711,N_701);
and U779 (N_779,N_725,N_700);
nor U780 (N_780,N_708,N_721);
nand U781 (N_781,N_721,N_731);
nor U782 (N_782,N_709,N_720);
xnor U783 (N_783,N_704,N_747);
or U784 (N_784,N_741,N_735);
or U785 (N_785,N_729,N_709);
or U786 (N_786,N_720,N_716);
or U787 (N_787,N_749,N_737);
or U788 (N_788,N_703,N_704);
nor U789 (N_789,N_743,N_717);
nand U790 (N_790,N_731,N_730);
and U791 (N_791,N_719,N_746);
and U792 (N_792,N_701,N_700);
nand U793 (N_793,N_743,N_716);
xnor U794 (N_794,N_737,N_746);
or U795 (N_795,N_744,N_748);
or U796 (N_796,N_742,N_722);
nand U797 (N_797,N_723,N_728);
or U798 (N_798,N_705,N_737);
nor U799 (N_799,N_707,N_739);
nor U800 (N_800,N_799,N_787);
xor U801 (N_801,N_765,N_780);
nand U802 (N_802,N_769,N_773);
and U803 (N_803,N_753,N_772);
nand U804 (N_804,N_792,N_757);
nand U805 (N_805,N_781,N_775);
and U806 (N_806,N_791,N_777);
nand U807 (N_807,N_797,N_782);
nor U808 (N_808,N_752,N_755);
and U809 (N_809,N_766,N_761);
or U810 (N_810,N_798,N_768);
nand U811 (N_811,N_786,N_774);
and U812 (N_812,N_763,N_784);
nor U813 (N_813,N_764,N_793);
xor U814 (N_814,N_779,N_751);
nor U815 (N_815,N_794,N_759);
or U816 (N_816,N_785,N_790);
nand U817 (N_817,N_754,N_758);
or U818 (N_818,N_760,N_783);
nand U819 (N_819,N_796,N_788);
or U820 (N_820,N_756,N_750);
nand U821 (N_821,N_789,N_795);
or U822 (N_822,N_771,N_778);
or U823 (N_823,N_767,N_776);
nand U824 (N_824,N_770,N_762);
nand U825 (N_825,N_768,N_797);
or U826 (N_826,N_782,N_776);
or U827 (N_827,N_755,N_779);
nor U828 (N_828,N_791,N_758);
nor U829 (N_829,N_776,N_792);
nor U830 (N_830,N_775,N_766);
xnor U831 (N_831,N_769,N_796);
and U832 (N_832,N_789,N_778);
nor U833 (N_833,N_779,N_792);
and U834 (N_834,N_790,N_792);
and U835 (N_835,N_751,N_761);
xnor U836 (N_836,N_757,N_766);
xnor U837 (N_837,N_756,N_767);
or U838 (N_838,N_768,N_766);
or U839 (N_839,N_776,N_760);
or U840 (N_840,N_761,N_754);
nand U841 (N_841,N_779,N_776);
and U842 (N_842,N_764,N_762);
nand U843 (N_843,N_788,N_751);
nand U844 (N_844,N_753,N_797);
nor U845 (N_845,N_764,N_792);
or U846 (N_846,N_778,N_773);
nand U847 (N_847,N_769,N_763);
xnor U848 (N_848,N_787,N_774);
and U849 (N_849,N_762,N_754);
nor U850 (N_850,N_803,N_811);
or U851 (N_851,N_808,N_801);
nor U852 (N_852,N_815,N_847);
xnor U853 (N_853,N_816,N_842);
nand U854 (N_854,N_826,N_848);
or U855 (N_855,N_840,N_824);
nand U856 (N_856,N_822,N_839);
or U857 (N_857,N_838,N_844);
or U858 (N_858,N_818,N_841);
nand U859 (N_859,N_807,N_804);
nor U860 (N_860,N_817,N_813);
or U861 (N_861,N_843,N_827);
nor U862 (N_862,N_805,N_831);
xor U863 (N_863,N_812,N_806);
xnor U864 (N_864,N_835,N_836);
or U865 (N_865,N_828,N_821);
and U866 (N_866,N_833,N_820);
nor U867 (N_867,N_800,N_830);
and U868 (N_868,N_845,N_810);
or U869 (N_869,N_846,N_829);
nand U870 (N_870,N_837,N_825);
xnor U871 (N_871,N_814,N_823);
nand U872 (N_872,N_819,N_849);
xnor U873 (N_873,N_832,N_809);
nor U874 (N_874,N_834,N_802);
xor U875 (N_875,N_808,N_816);
nor U876 (N_876,N_802,N_846);
xor U877 (N_877,N_806,N_818);
and U878 (N_878,N_847,N_811);
and U879 (N_879,N_816,N_847);
xnor U880 (N_880,N_827,N_836);
nand U881 (N_881,N_814,N_821);
and U882 (N_882,N_843,N_846);
and U883 (N_883,N_825,N_829);
nand U884 (N_884,N_812,N_808);
nand U885 (N_885,N_814,N_809);
nor U886 (N_886,N_812,N_849);
or U887 (N_887,N_837,N_807);
nor U888 (N_888,N_820,N_843);
xor U889 (N_889,N_801,N_832);
and U890 (N_890,N_848,N_809);
xnor U891 (N_891,N_849,N_809);
nand U892 (N_892,N_818,N_802);
or U893 (N_893,N_847,N_848);
and U894 (N_894,N_848,N_820);
nor U895 (N_895,N_833,N_841);
or U896 (N_896,N_846,N_827);
and U897 (N_897,N_824,N_837);
or U898 (N_898,N_807,N_831);
xor U899 (N_899,N_842,N_843);
and U900 (N_900,N_861,N_887);
and U901 (N_901,N_851,N_894);
nand U902 (N_902,N_854,N_868);
nor U903 (N_903,N_875,N_895);
nor U904 (N_904,N_899,N_857);
nor U905 (N_905,N_871,N_859);
nand U906 (N_906,N_879,N_850);
nor U907 (N_907,N_860,N_858);
xnor U908 (N_908,N_891,N_866);
nor U909 (N_909,N_878,N_872);
nand U910 (N_910,N_889,N_873);
nor U911 (N_911,N_897,N_863);
nand U912 (N_912,N_883,N_862);
nand U913 (N_913,N_892,N_890);
and U914 (N_914,N_864,N_870);
nor U915 (N_915,N_896,N_869);
or U916 (N_916,N_884,N_855);
xnor U917 (N_917,N_865,N_874);
nand U918 (N_918,N_885,N_888);
xor U919 (N_919,N_880,N_886);
nor U920 (N_920,N_881,N_898);
or U921 (N_921,N_852,N_893);
nand U922 (N_922,N_876,N_853);
and U923 (N_923,N_882,N_856);
xor U924 (N_924,N_877,N_867);
and U925 (N_925,N_885,N_898);
nand U926 (N_926,N_885,N_876);
and U927 (N_927,N_861,N_889);
nand U928 (N_928,N_898,N_882);
or U929 (N_929,N_853,N_863);
xor U930 (N_930,N_897,N_884);
nor U931 (N_931,N_851,N_881);
and U932 (N_932,N_854,N_888);
nor U933 (N_933,N_866,N_852);
and U934 (N_934,N_853,N_879);
nand U935 (N_935,N_871,N_874);
nand U936 (N_936,N_899,N_896);
or U937 (N_937,N_888,N_878);
or U938 (N_938,N_877,N_875);
and U939 (N_939,N_866,N_864);
nor U940 (N_940,N_855,N_851);
xor U941 (N_941,N_891,N_850);
xor U942 (N_942,N_855,N_882);
and U943 (N_943,N_881,N_877);
xnor U944 (N_944,N_861,N_898);
and U945 (N_945,N_864,N_881);
nor U946 (N_946,N_871,N_851);
nand U947 (N_947,N_894,N_890);
or U948 (N_948,N_892,N_881);
nand U949 (N_949,N_882,N_878);
nand U950 (N_950,N_902,N_904);
nand U951 (N_951,N_947,N_911);
or U952 (N_952,N_906,N_915);
and U953 (N_953,N_922,N_941);
nor U954 (N_954,N_920,N_908);
nand U955 (N_955,N_921,N_929);
nor U956 (N_956,N_945,N_917);
and U957 (N_957,N_946,N_932);
and U958 (N_958,N_927,N_928);
nand U959 (N_959,N_931,N_903);
or U960 (N_960,N_942,N_940);
or U961 (N_961,N_907,N_937);
or U962 (N_962,N_918,N_930);
or U963 (N_963,N_938,N_905);
nand U964 (N_964,N_919,N_910);
or U965 (N_965,N_913,N_935);
nand U966 (N_966,N_934,N_924);
nor U967 (N_967,N_912,N_901);
and U968 (N_968,N_925,N_948);
xnor U969 (N_969,N_939,N_944);
or U970 (N_970,N_916,N_949);
nand U971 (N_971,N_926,N_900);
nor U972 (N_972,N_943,N_909);
nor U973 (N_973,N_914,N_936);
xnor U974 (N_974,N_933,N_923);
nand U975 (N_975,N_901,N_933);
and U976 (N_976,N_915,N_937);
nand U977 (N_977,N_928,N_917);
xor U978 (N_978,N_928,N_937);
xnor U979 (N_979,N_916,N_913);
xnor U980 (N_980,N_925,N_934);
and U981 (N_981,N_944,N_917);
nor U982 (N_982,N_931,N_913);
or U983 (N_983,N_936,N_932);
and U984 (N_984,N_915,N_934);
nand U985 (N_985,N_932,N_903);
nand U986 (N_986,N_907,N_920);
or U987 (N_987,N_937,N_900);
nor U988 (N_988,N_944,N_924);
nand U989 (N_989,N_919,N_900);
xnor U990 (N_990,N_908,N_919);
and U991 (N_991,N_945,N_929);
and U992 (N_992,N_933,N_939);
nand U993 (N_993,N_940,N_914);
nand U994 (N_994,N_913,N_932);
xnor U995 (N_995,N_937,N_949);
or U996 (N_996,N_932,N_911);
xor U997 (N_997,N_914,N_928);
or U998 (N_998,N_912,N_932);
nand U999 (N_999,N_906,N_949);
or U1000 (N_1000,N_996,N_986);
nor U1001 (N_1001,N_995,N_982);
and U1002 (N_1002,N_987,N_990);
or U1003 (N_1003,N_969,N_971);
and U1004 (N_1004,N_950,N_999);
and U1005 (N_1005,N_967,N_977);
xor U1006 (N_1006,N_973,N_983);
or U1007 (N_1007,N_972,N_981);
nor U1008 (N_1008,N_985,N_993);
xor U1009 (N_1009,N_984,N_953);
nor U1010 (N_1010,N_965,N_976);
or U1011 (N_1011,N_952,N_968);
and U1012 (N_1012,N_998,N_956);
nor U1013 (N_1013,N_975,N_954);
or U1014 (N_1014,N_997,N_970);
or U1015 (N_1015,N_979,N_980);
nand U1016 (N_1016,N_964,N_963);
nor U1017 (N_1017,N_959,N_994);
nand U1018 (N_1018,N_955,N_974);
and U1019 (N_1019,N_961,N_989);
and U1020 (N_1020,N_957,N_951);
or U1021 (N_1021,N_962,N_978);
or U1022 (N_1022,N_966,N_992);
and U1023 (N_1023,N_960,N_958);
nand U1024 (N_1024,N_988,N_991);
nand U1025 (N_1025,N_990,N_956);
or U1026 (N_1026,N_970,N_988);
xor U1027 (N_1027,N_956,N_976);
xor U1028 (N_1028,N_972,N_964);
xor U1029 (N_1029,N_951,N_998);
nor U1030 (N_1030,N_958,N_975);
xnor U1031 (N_1031,N_962,N_986);
nand U1032 (N_1032,N_968,N_998);
or U1033 (N_1033,N_957,N_998);
and U1034 (N_1034,N_962,N_969);
and U1035 (N_1035,N_967,N_954);
or U1036 (N_1036,N_981,N_988);
nor U1037 (N_1037,N_999,N_990);
nor U1038 (N_1038,N_955,N_990);
nand U1039 (N_1039,N_972,N_956);
nand U1040 (N_1040,N_987,N_955);
nand U1041 (N_1041,N_954,N_989);
xnor U1042 (N_1042,N_989,N_964);
or U1043 (N_1043,N_955,N_952);
and U1044 (N_1044,N_984,N_968);
nand U1045 (N_1045,N_992,N_970);
nand U1046 (N_1046,N_984,N_975);
nor U1047 (N_1047,N_959,N_970);
nor U1048 (N_1048,N_950,N_998);
nand U1049 (N_1049,N_961,N_962);
nor U1050 (N_1050,N_1026,N_1033);
nor U1051 (N_1051,N_1042,N_1046);
or U1052 (N_1052,N_1030,N_1018);
and U1053 (N_1053,N_1040,N_1003);
nor U1054 (N_1054,N_1004,N_1021);
nor U1055 (N_1055,N_1005,N_1000);
nor U1056 (N_1056,N_1017,N_1027);
xnor U1057 (N_1057,N_1020,N_1045);
xnor U1058 (N_1058,N_1006,N_1016);
nand U1059 (N_1059,N_1048,N_1011);
and U1060 (N_1060,N_1007,N_1029);
nand U1061 (N_1061,N_1043,N_1025);
nor U1062 (N_1062,N_1014,N_1022);
nand U1063 (N_1063,N_1002,N_1023);
nand U1064 (N_1064,N_1009,N_1034);
nor U1065 (N_1065,N_1032,N_1039);
or U1066 (N_1066,N_1013,N_1036);
and U1067 (N_1067,N_1041,N_1024);
xor U1068 (N_1068,N_1008,N_1037);
xor U1069 (N_1069,N_1035,N_1044);
nand U1070 (N_1070,N_1001,N_1010);
nor U1071 (N_1071,N_1019,N_1049);
and U1072 (N_1072,N_1012,N_1028);
nand U1073 (N_1073,N_1038,N_1031);
nor U1074 (N_1074,N_1015,N_1047);
or U1075 (N_1075,N_1044,N_1000);
nor U1076 (N_1076,N_1007,N_1022);
or U1077 (N_1077,N_1031,N_1015);
or U1078 (N_1078,N_1002,N_1046);
or U1079 (N_1079,N_1020,N_1015);
or U1080 (N_1080,N_1047,N_1022);
xnor U1081 (N_1081,N_1020,N_1001);
xnor U1082 (N_1082,N_1029,N_1015);
and U1083 (N_1083,N_1021,N_1040);
and U1084 (N_1084,N_1018,N_1003);
nand U1085 (N_1085,N_1030,N_1021);
xor U1086 (N_1086,N_1010,N_1022);
xor U1087 (N_1087,N_1031,N_1026);
nand U1088 (N_1088,N_1029,N_1025);
or U1089 (N_1089,N_1030,N_1034);
or U1090 (N_1090,N_1034,N_1037);
or U1091 (N_1091,N_1012,N_1006);
xor U1092 (N_1092,N_1009,N_1047);
nor U1093 (N_1093,N_1015,N_1025);
nand U1094 (N_1094,N_1001,N_1036);
and U1095 (N_1095,N_1044,N_1006);
nor U1096 (N_1096,N_1045,N_1024);
xnor U1097 (N_1097,N_1031,N_1040);
nor U1098 (N_1098,N_1039,N_1000);
nor U1099 (N_1099,N_1013,N_1006);
and U1100 (N_1100,N_1098,N_1091);
xnor U1101 (N_1101,N_1069,N_1060);
nand U1102 (N_1102,N_1080,N_1094);
nand U1103 (N_1103,N_1054,N_1076);
nor U1104 (N_1104,N_1066,N_1096);
nand U1105 (N_1105,N_1084,N_1061);
and U1106 (N_1106,N_1070,N_1079);
and U1107 (N_1107,N_1067,N_1071);
nand U1108 (N_1108,N_1062,N_1057);
or U1109 (N_1109,N_1063,N_1072);
xor U1110 (N_1110,N_1093,N_1082);
xor U1111 (N_1111,N_1059,N_1058);
nor U1112 (N_1112,N_1085,N_1050);
or U1113 (N_1113,N_1089,N_1081);
and U1114 (N_1114,N_1088,N_1053);
xnor U1115 (N_1115,N_1073,N_1092);
and U1116 (N_1116,N_1068,N_1065);
nand U1117 (N_1117,N_1078,N_1087);
xnor U1118 (N_1118,N_1074,N_1075);
nor U1119 (N_1119,N_1056,N_1086);
nor U1120 (N_1120,N_1052,N_1099);
and U1121 (N_1121,N_1077,N_1051);
nand U1122 (N_1122,N_1055,N_1083);
and U1123 (N_1123,N_1095,N_1097);
and U1124 (N_1124,N_1090,N_1064);
nor U1125 (N_1125,N_1053,N_1080);
nor U1126 (N_1126,N_1064,N_1096);
or U1127 (N_1127,N_1073,N_1075);
or U1128 (N_1128,N_1068,N_1077);
xor U1129 (N_1129,N_1065,N_1054);
and U1130 (N_1130,N_1091,N_1096);
nor U1131 (N_1131,N_1096,N_1092);
nand U1132 (N_1132,N_1070,N_1076);
xor U1133 (N_1133,N_1050,N_1056);
xnor U1134 (N_1134,N_1055,N_1063);
and U1135 (N_1135,N_1058,N_1065);
xor U1136 (N_1136,N_1068,N_1088);
and U1137 (N_1137,N_1066,N_1063);
nor U1138 (N_1138,N_1086,N_1085);
nand U1139 (N_1139,N_1061,N_1053);
and U1140 (N_1140,N_1090,N_1076);
and U1141 (N_1141,N_1059,N_1066);
nand U1142 (N_1142,N_1080,N_1067);
or U1143 (N_1143,N_1091,N_1085);
nand U1144 (N_1144,N_1095,N_1080);
or U1145 (N_1145,N_1070,N_1052);
xor U1146 (N_1146,N_1060,N_1062);
xnor U1147 (N_1147,N_1082,N_1051);
nand U1148 (N_1148,N_1073,N_1074);
and U1149 (N_1149,N_1075,N_1069);
or U1150 (N_1150,N_1146,N_1141);
or U1151 (N_1151,N_1103,N_1121);
nand U1152 (N_1152,N_1104,N_1123);
xor U1153 (N_1153,N_1139,N_1120);
and U1154 (N_1154,N_1135,N_1129);
nand U1155 (N_1155,N_1108,N_1136);
nand U1156 (N_1156,N_1114,N_1130);
nand U1157 (N_1157,N_1144,N_1109);
and U1158 (N_1158,N_1125,N_1119);
nand U1159 (N_1159,N_1133,N_1116);
nand U1160 (N_1160,N_1102,N_1107);
xor U1161 (N_1161,N_1145,N_1124);
nand U1162 (N_1162,N_1122,N_1111);
xnor U1163 (N_1163,N_1128,N_1117);
and U1164 (N_1164,N_1115,N_1105);
and U1165 (N_1165,N_1149,N_1127);
and U1166 (N_1166,N_1113,N_1100);
nand U1167 (N_1167,N_1134,N_1106);
and U1168 (N_1168,N_1126,N_1131);
xor U1169 (N_1169,N_1138,N_1112);
nand U1170 (N_1170,N_1143,N_1101);
nor U1171 (N_1171,N_1148,N_1110);
nand U1172 (N_1172,N_1118,N_1137);
xnor U1173 (N_1173,N_1142,N_1147);
and U1174 (N_1174,N_1132,N_1140);
and U1175 (N_1175,N_1146,N_1119);
nand U1176 (N_1176,N_1123,N_1112);
or U1177 (N_1177,N_1136,N_1140);
or U1178 (N_1178,N_1114,N_1121);
nand U1179 (N_1179,N_1116,N_1111);
xor U1180 (N_1180,N_1100,N_1112);
and U1181 (N_1181,N_1138,N_1120);
xnor U1182 (N_1182,N_1143,N_1126);
nand U1183 (N_1183,N_1147,N_1127);
and U1184 (N_1184,N_1104,N_1113);
nor U1185 (N_1185,N_1145,N_1141);
nand U1186 (N_1186,N_1148,N_1136);
and U1187 (N_1187,N_1124,N_1147);
or U1188 (N_1188,N_1109,N_1147);
or U1189 (N_1189,N_1111,N_1117);
xnor U1190 (N_1190,N_1124,N_1107);
xnor U1191 (N_1191,N_1100,N_1140);
xnor U1192 (N_1192,N_1137,N_1148);
and U1193 (N_1193,N_1131,N_1132);
xor U1194 (N_1194,N_1148,N_1124);
nand U1195 (N_1195,N_1119,N_1118);
nor U1196 (N_1196,N_1138,N_1119);
nor U1197 (N_1197,N_1129,N_1120);
nand U1198 (N_1198,N_1103,N_1146);
or U1199 (N_1199,N_1147,N_1115);
and U1200 (N_1200,N_1190,N_1173);
and U1201 (N_1201,N_1196,N_1164);
nor U1202 (N_1202,N_1169,N_1181);
or U1203 (N_1203,N_1161,N_1195);
nor U1204 (N_1204,N_1189,N_1160);
xnor U1205 (N_1205,N_1194,N_1178);
nor U1206 (N_1206,N_1159,N_1192);
xnor U1207 (N_1207,N_1180,N_1158);
nor U1208 (N_1208,N_1170,N_1188);
nand U1209 (N_1209,N_1151,N_1197);
xor U1210 (N_1210,N_1154,N_1171);
xnor U1211 (N_1211,N_1185,N_1182);
and U1212 (N_1212,N_1198,N_1177);
or U1213 (N_1213,N_1153,N_1152);
nand U1214 (N_1214,N_1199,N_1163);
and U1215 (N_1215,N_1175,N_1166);
xor U1216 (N_1216,N_1165,N_1157);
or U1217 (N_1217,N_1184,N_1162);
or U1218 (N_1218,N_1186,N_1183);
xor U1219 (N_1219,N_1156,N_1193);
or U1220 (N_1220,N_1176,N_1167);
nand U1221 (N_1221,N_1174,N_1150);
nand U1222 (N_1222,N_1172,N_1187);
and U1223 (N_1223,N_1191,N_1168);
nor U1224 (N_1224,N_1155,N_1179);
nor U1225 (N_1225,N_1198,N_1193);
nor U1226 (N_1226,N_1164,N_1189);
or U1227 (N_1227,N_1152,N_1191);
or U1228 (N_1228,N_1166,N_1167);
and U1229 (N_1229,N_1172,N_1173);
or U1230 (N_1230,N_1150,N_1168);
xor U1231 (N_1231,N_1159,N_1183);
or U1232 (N_1232,N_1158,N_1165);
or U1233 (N_1233,N_1199,N_1190);
and U1234 (N_1234,N_1176,N_1152);
and U1235 (N_1235,N_1161,N_1171);
and U1236 (N_1236,N_1157,N_1182);
nand U1237 (N_1237,N_1158,N_1152);
xnor U1238 (N_1238,N_1162,N_1193);
and U1239 (N_1239,N_1150,N_1154);
nor U1240 (N_1240,N_1176,N_1191);
or U1241 (N_1241,N_1172,N_1191);
or U1242 (N_1242,N_1162,N_1198);
or U1243 (N_1243,N_1183,N_1154);
nor U1244 (N_1244,N_1164,N_1159);
nand U1245 (N_1245,N_1187,N_1184);
and U1246 (N_1246,N_1192,N_1193);
nor U1247 (N_1247,N_1160,N_1159);
nor U1248 (N_1248,N_1180,N_1177);
or U1249 (N_1249,N_1192,N_1166);
nor U1250 (N_1250,N_1240,N_1220);
nand U1251 (N_1251,N_1215,N_1245);
xnor U1252 (N_1252,N_1206,N_1236);
nand U1253 (N_1253,N_1231,N_1230);
and U1254 (N_1254,N_1201,N_1209);
nor U1255 (N_1255,N_1211,N_1229);
nor U1256 (N_1256,N_1203,N_1243);
nand U1257 (N_1257,N_1249,N_1246);
nand U1258 (N_1258,N_1233,N_1225);
and U1259 (N_1259,N_1219,N_1235);
nor U1260 (N_1260,N_1228,N_1210);
nand U1261 (N_1261,N_1237,N_1213);
xnor U1262 (N_1262,N_1208,N_1204);
and U1263 (N_1263,N_1242,N_1248);
nor U1264 (N_1264,N_1202,N_1218);
or U1265 (N_1265,N_1224,N_1239);
nor U1266 (N_1266,N_1216,N_1241);
nor U1267 (N_1267,N_1234,N_1222);
and U1268 (N_1268,N_1217,N_1214);
nor U1269 (N_1269,N_1212,N_1223);
nor U1270 (N_1270,N_1232,N_1244);
nand U1271 (N_1271,N_1205,N_1247);
nor U1272 (N_1272,N_1200,N_1238);
nand U1273 (N_1273,N_1221,N_1207);
and U1274 (N_1274,N_1226,N_1227);
or U1275 (N_1275,N_1247,N_1235);
nand U1276 (N_1276,N_1206,N_1229);
and U1277 (N_1277,N_1238,N_1230);
and U1278 (N_1278,N_1210,N_1218);
or U1279 (N_1279,N_1225,N_1249);
nand U1280 (N_1280,N_1246,N_1224);
or U1281 (N_1281,N_1215,N_1212);
nand U1282 (N_1282,N_1245,N_1203);
xor U1283 (N_1283,N_1211,N_1245);
or U1284 (N_1284,N_1228,N_1240);
or U1285 (N_1285,N_1235,N_1221);
and U1286 (N_1286,N_1210,N_1223);
xor U1287 (N_1287,N_1221,N_1237);
and U1288 (N_1288,N_1241,N_1224);
or U1289 (N_1289,N_1225,N_1234);
or U1290 (N_1290,N_1245,N_1218);
nor U1291 (N_1291,N_1247,N_1229);
and U1292 (N_1292,N_1245,N_1217);
nand U1293 (N_1293,N_1200,N_1228);
nor U1294 (N_1294,N_1232,N_1200);
nand U1295 (N_1295,N_1206,N_1205);
or U1296 (N_1296,N_1221,N_1201);
xor U1297 (N_1297,N_1200,N_1206);
xor U1298 (N_1298,N_1212,N_1210);
nand U1299 (N_1299,N_1223,N_1230);
nand U1300 (N_1300,N_1297,N_1290);
and U1301 (N_1301,N_1252,N_1268);
or U1302 (N_1302,N_1294,N_1266);
nor U1303 (N_1303,N_1288,N_1280);
nor U1304 (N_1304,N_1255,N_1293);
or U1305 (N_1305,N_1251,N_1258);
and U1306 (N_1306,N_1286,N_1262);
or U1307 (N_1307,N_1281,N_1295);
nor U1308 (N_1308,N_1257,N_1298);
or U1309 (N_1309,N_1250,N_1275);
nor U1310 (N_1310,N_1277,N_1269);
or U1311 (N_1311,N_1285,N_1292);
nand U1312 (N_1312,N_1263,N_1296);
nand U1313 (N_1313,N_1267,N_1278);
xor U1314 (N_1314,N_1276,N_1272);
xnor U1315 (N_1315,N_1261,N_1287);
xor U1316 (N_1316,N_1270,N_1260);
and U1317 (N_1317,N_1289,N_1274);
or U1318 (N_1318,N_1299,N_1282);
nor U1319 (N_1319,N_1284,N_1279);
nand U1320 (N_1320,N_1254,N_1264);
and U1321 (N_1321,N_1265,N_1256);
nand U1322 (N_1322,N_1259,N_1283);
nand U1323 (N_1323,N_1273,N_1271);
or U1324 (N_1324,N_1291,N_1253);
xnor U1325 (N_1325,N_1261,N_1289);
nand U1326 (N_1326,N_1288,N_1257);
nor U1327 (N_1327,N_1254,N_1293);
and U1328 (N_1328,N_1275,N_1282);
or U1329 (N_1329,N_1266,N_1296);
and U1330 (N_1330,N_1280,N_1278);
or U1331 (N_1331,N_1291,N_1286);
or U1332 (N_1332,N_1277,N_1265);
nor U1333 (N_1333,N_1294,N_1256);
and U1334 (N_1334,N_1287,N_1279);
and U1335 (N_1335,N_1268,N_1283);
xnor U1336 (N_1336,N_1267,N_1280);
and U1337 (N_1337,N_1285,N_1286);
nor U1338 (N_1338,N_1295,N_1290);
nand U1339 (N_1339,N_1256,N_1286);
nand U1340 (N_1340,N_1289,N_1257);
and U1341 (N_1341,N_1274,N_1277);
xnor U1342 (N_1342,N_1251,N_1290);
xor U1343 (N_1343,N_1281,N_1272);
and U1344 (N_1344,N_1250,N_1263);
or U1345 (N_1345,N_1287,N_1282);
nor U1346 (N_1346,N_1283,N_1255);
nor U1347 (N_1347,N_1258,N_1257);
or U1348 (N_1348,N_1266,N_1264);
nor U1349 (N_1349,N_1267,N_1292);
and U1350 (N_1350,N_1317,N_1335);
and U1351 (N_1351,N_1336,N_1334);
or U1352 (N_1352,N_1311,N_1315);
nand U1353 (N_1353,N_1326,N_1306);
nand U1354 (N_1354,N_1321,N_1332);
and U1355 (N_1355,N_1302,N_1347);
and U1356 (N_1356,N_1341,N_1340);
and U1357 (N_1357,N_1324,N_1305);
xnor U1358 (N_1358,N_1314,N_1320);
nand U1359 (N_1359,N_1301,N_1346);
and U1360 (N_1360,N_1330,N_1325);
xor U1361 (N_1361,N_1331,N_1323);
and U1362 (N_1362,N_1312,N_1338);
and U1363 (N_1363,N_1318,N_1344);
xor U1364 (N_1364,N_1307,N_1342);
and U1365 (N_1365,N_1345,N_1310);
and U1366 (N_1366,N_1319,N_1339);
or U1367 (N_1367,N_1303,N_1349);
or U1368 (N_1368,N_1322,N_1300);
and U1369 (N_1369,N_1313,N_1329);
or U1370 (N_1370,N_1333,N_1348);
and U1371 (N_1371,N_1327,N_1343);
nor U1372 (N_1372,N_1328,N_1309);
and U1373 (N_1373,N_1308,N_1316);
and U1374 (N_1374,N_1304,N_1337);
and U1375 (N_1375,N_1310,N_1338);
and U1376 (N_1376,N_1310,N_1328);
xor U1377 (N_1377,N_1339,N_1325);
nand U1378 (N_1378,N_1301,N_1338);
nor U1379 (N_1379,N_1343,N_1302);
xnor U1380 (N_1380,N_1338,N_1328);
nor U1381 (N_1381,N_1349,N_1315);
and U1382 (N_1382,N_1341,N_1301);
nand U1383 (N_1383,N_1336,N_1313);
nor U1384 (N_1384,N_1306,N_1313);
or U1385 (N_1385,N_1303,N_1304);
nor U1386 (N_1386,N_1336,N_1346);
nand U1387 (N_1387,N_1314,N_1317);
and U1388 (N_1388,N_1319,N_1320);
and U1389 (N_1389,N_1309,N_1342);
xnor U1390 (N_1390,N_1322,N_1301);
or U1391 (N_1391,N_1334,N_1316);
xnor U1392 (N_1392,N_1308,N_1343);
nand U1393 (N_1393,N_1317,N_1303);
xnor U1394 (N_1394,N_1329,N_1331);
or U1395 (N_1395,N_1316,N_1331);
nor U1396 (N_1396,N_1303,N_1302);
or U1397 (N_1397,N_1334,N_1319);
xnor U1398 (N_1398,N_1331,N_1344);
nand U1399 (N_1399,N_1316,N_1348);
and U1400 (N_1400,N_1383,N_1399);
nand U1401 (N_1401,N_1372,N_1389);
or U1402 (N_1402,N_1355,N_1379);
or U1403 (N_1403,N_1398,N_1378);
or U1404 (N_1404,N_1363,N_1370);
or U1405 (N_1405,N_1350,N_1396);
or U1406 (N_1406,N_1387,N_1368);
nand U1407 (N_1407,N_1382,N_1358);
nor U1408 (N_1408,N_1377,N_1397);
or U1409 (N_1409,N_1360,N_1352);
nor U1410 (N_1410,N_1354,N_1357);
or U1411 (N_1411,N_1353,N_1384);
and U1412 (N_1412,N_1366,N_1391);
nor U1413 (N_1413,N_1365,N_1394);
nor U1414 (N_1414,N_1374,N_1393);
and U1415 (N_1415,N_1359,N_1371);
and U1416 (N_1416,N_1361,N_1395);
or U1417 (N_1417,N_1381,N_1373);
nor U1418 (N_1418,N_1369,N_1364);
and U1419 (N_1419,N_1388,N_1375);
or U1420 (N_1420,N_1351,N_1356);
or U1421 (N_1421,N_1376,N_1385);
xnor U1422 (N_1422,N_1386,N_1392);
or U1423 (N_1423,N_1367,N_1362);
nand U1424 (N_1424,N_1390,N_1380);
nor U1425 (N_1425,N_1392,N_1398);
or U1426 (N_1426,N_1368,N_1377);
and U1427 (N_1427,N_1398,N_1369);
nand U1428 (N_1428,N_1362,N_1359);
nor U1429 (N_1429,N_1380,N_1388);
or U1430 (N_1430,N_1386,N_1363);
nand U1431 (N_1431,N_1353,N_1389);
nand U1432 (N_1432,N_1360,N_1390);
xor U1433 (N_1433,N_1385,N_1353);
or U1434 (N_1434,N_1353,N_1375);
xnor U1435 (N_1435,N_1384,N_1374);
or U1436 (N_1436,N_1387,N_1372);
or U1437 (N_1437,N_1362,N_1379);
nand U1438 (N_1438,N_1355,N_1397);
and U1439 (N_1439,N_1352,N_1398);
nor U1440 (N_1440,N_1359,N_1351);
and U1441 (N_1441,N_1370,N_1367);
or U1442 (N_1442,N_1398,N_1373);
and U1443 (N_1443,N_1397,N_1350);
or U1444 (N_1444,N_1392,N_1383);
xnor U1445 (N_1445,N_1352,N_1399);
and U1446 (N_1446,N_1389,N_1352);
nor U1447 (N_1447,N_1357,N_1366);
nand U1448 (N_1448,N_1383,N_1350);
nor U1449 (N_1449,N_1391,N_1398);
nor U1450 (N_1450,N_1440,N_1402);
or U1451 (N_1451,N_1426,N_1412);
xor U1452 (N_1452,N_1418,N_1401);
and U1453 (N_1453,N_1407,N_1404);
nand U1454 (N_1454,N_1417,N_1427);
and U1455 (N_1455,N_1415,N_1431);
nand U1456 (N_1456,N_1448,N_1442);
or U1457 (N_1457,N_1433,N_1414);
and U1458 (N_1458,N_1410,N_1406);
xnor U1459 (N_1459,N_1443,N_1423);
or U1460 (N_1460,N_1408,N_1446);
or U1461 (N_1461,N_1437,N_1444);
nor U1462 (N_1462,N_1416,N_1428);
or U1463 (N_1463,N_1432,N_1435);
nand U1464 (N_1464,N_1441,N_1400);
and U1465 (N_1465,N_1436,N_1419);
nand U1466 (N_1466,N_1411,N_1422);
nand U1467 (N_1467,N_1439,N_1434);
and U1468 (N_1468,N_1413,N_1424);
and U1469 (N_1469,N_1420,N_1438);
or U1470 (N_1470,N_1449,N_1421);
or U1471 (N_1471,N_1403,N_1447);
or U1472 (N_1472,N_1445,N_1425);
and U1473 (N_1473,N_1405,N_1430);
xnor U1474 (N_1474,N_1429,N_1409);
or U1475 (N_1475,N_1440,N_1415);
xor U1476 (N_1476,N_1435,N_1421);
nand U1477 (N_1477,N_1438,N_1408);
or U1478 (N_1478,N_1411,N_1420);
nor U1479 (N_1479,N_1404,N_1414);
or U1480 (N_1480,N_1445,N_1419);
nand U1481 (N_1481,N_1448,N_1410);
xor U1482 (N_1482,N_1406,N_1431);
xor U1483 (N_1483,N_1434,N_1432);
xnor U1484 (N_1484,N_1443,N_1422);
xor U1485 (N_1485,N_1407,N_1417);
nand U1486 (N_1486,N_1411,N_1417);
nand U1487 (N_1487,N_1432,N_1433);
nand U1488 (N_1488,N_1431,N_1430);
nand U1489 (N_1489,N_1408,N_1403);
xnor U1490 (N_1490,N_1447,N_1426);
and U1491 (N_1491,N_1400,N_1405);
nor U1492 (N_1492,N_1427,N_1413);
nor U1493 (N_1493,N_1426,N_1439);
xnor U1494 (N_1494,N_1443,N_1419);
nor U1495 (N_1495,N_1431,N_1421);
xor U1496 (N_1496,N_1403,N_1448);
and U1497 (N_1497,N_1427,N_1414);
nand U1498 (N_1498,N_1416,N_1448);
nand U1499 (N_1499,N_1441,N_1427);
nand U1500 (N_1500,N_1498,N_1477);
and U1501 (N_1501,N_1467,N_1478);
and U1502 (N_1502,N_1482,N_1458);
and U1503 (N_1503,N_1466,N_1452);
nand U1504 (N_1504,N_1484,N_1453);
xnor U1505 (N_1505,N_1456,N_1462);
xnor U1506 (N_1506,N_1460,N_1480);
nor U1507 (N_1507,N_1457,N_1455);
and U1508 (N_1508,N_1494,N_1468);
nor U1509 (N_1509,N_1454,N_1472);
nand U1510 (N_1510,N_1471,N_1487);
xor U1511 (N_1511,N_1474,N_1486);
nand U1512 (N_1512,N_1451,N_1461);
nand U1513 (N_1513,N_1464,N_1459);
or U1514 (N_1514,N_1499,N_1476);
or U1515 (N_1515,N_1470,N_1465);
xor U1516 (N_1516,N_1450,N_1475);
or U1517 (N_1517,N_1493,N_1463);
nor U1518 (N_1518,N_1483,N_1490);
or U1519 (N_1519,N_1491,N_1497);
and U1520 (N_1520,N_1488,N_1479);
or U1521 (N_1521,N_1485,N_1492);
nor U1522 (N_1522,N_1495,N_1473);
and U1523 (N_1523,N_1496,N_1481);
and U1524 (N_1524,N_1469,N_1489);
and U1525 (N_1525,N_1471,N_1457);
nand U1526 (N_1526,N_1479,N_1499);
nor U1527 (N_1527,N_1455,N_1462);
nor U1528 (N_1528,N_1454,N_1487);
xnor U1529 (N_1529,N_1459,N_1494);
nor U1530 (N_1530,N_1492,N_1487);
nand U1531 (N_1531,N_1469,N_1471);
nor U1532 (N_1532,N_1464,N_1451);
and U1533 (N_1533,N_1454,N_1450);
nand U1534 (N_1534,N_1480,N_1491);
nor U1535 (N_1535,N_1468,N_1489);
and U1536 (N_1536,N_1490,N_1498);
nand U1537 (N_1537,N_1483,N_1491);
nor U1538 (N_1538,N_1495,N_1486);
and U1539 (N_1539,N_1454,N_1482);
nand U1540 (N_1540,N_1479,N_1453);
or U1541 (N_1541,N_1475,N_1471);
and U1542 (N_1542,N_1459,N_1478);
and U1543 (N_1543,N_1481,N_1491);
xnor U1544 (N_1544,N_1490,N_1453);
nor U1545 (N_1545,N_1450,N_1465);
nor U1546 (N_1546,N_1486,N_1482);
or U1547 (N_1547,N_1484,N_1473);
or U1548 (N_1548,N_1450,N_1489);
nor U1549 (N_1549,N_1456,N_1473);
and U1550 (N_1550,N_1507,N_1512);
and U1551 (N_1551,N_1524,N_1500);
xnor U1552 (N_1552,N_1529,N_1502);
nand U1553 (N_1553,N_1541,N_1516);
and U1554 (N_1554,N_1525,N_1539);
or U1555 (N_1555,N_1514,N_1517);
and U1556 (N_1556,N_1522,N_1543);
or U1557 (N_1557,N_1508,N_1532);
and U1558 (N_1558,N_1518,N_1546);
nor U1559 (N_1559,N_1548,N_1549);
or U1560 (N_1560,N_1515,N_1511);
nand U1561 (N_1561,N_1531,N_1501);
or U1562 (N_1562,N_1526,N_1528);
nor U1563 (N_1563,N_1519,N_1538);
or U1564 (N_1564,N_1504,N_1503);
nand U1565 (N_1565,N_1523,N_1540);
nand U1566 (N_1566,N_1521,N_1536);
xnor U1567 (N_1567,N_1506,N_1513);
xnor U1568 (N_1568,N_1547,N_1542);
or U1569 (N_1569,N_1537,N_1535);
nand U1570 (N_1570,N_1510,N_1520);
and U1571 (N_1571,N_1533,N_1534);
xnor U1572 (N_1572,N_1545,N_1527);
and U1573 (N_1573,N_1505,N_1509);
xor U1574 (N_1574,N_1544,N_1530);
nor U1575 (N_1575,N_1545,N_1514);
and U1576 (N_1576,N_1547,N_1548);
nor U1577 (N_1577,N_1549,N_1510);
nand U1578 (N_1578,N_1503,N_1515);
nor U1579 (N_1579,N_1542,N_1539);
or U1580 (N_1580,N_1518,N_1521);
xnor U1581 (N_1581,N_1521,N_1507);
xnor U1582 (N_1582,N_1542,N_1521);
and U1583 (N_1583,N_1527,N_1534);
nand U1584 (N_1584,N_1502,N_1510);
nand U1585 (N_1585,N_1509,N_1503);
nor U1586 (N_1586,N_1508,N_1544);
nand U1587 (N_1587,N_1532,N_1526);
xor U1588 (N_1588,N_1531,N_1528);
nand U1589 (N_1589,N_1514,N_1542);
xnor U1590 (N_1590,N_1510,N_1529);
nor U1591 (N_1591,N_1517,N_1535);
and U1592 (N_1592,N_1533,N_1500);
nand U1593 (N_1593,N_1527,N_1508);
nand U1594 (N_1594,N_1545,N_1533);
nand U1595 (N_1595,N_1508,N_1528);
nor U1596 (N_1596,N_1514,N_1527);
nor U1597 (N_1597,N_1542,N_1518);
xnor U1598 (N_1598,N_1508,N_1530);
nor U1599 (N_1599,N_1539,N_1518);
and U1600 (N_1600,N_1551,N_1561);
nor U1601 (N_1601,N_1567,N_1589);
or U1602 (N_1602,N_1584,N_1569);
xnor U1603 (N_1603,N_1588,N_1598);
xor U1604 (N_1604,N_1585,N_1596);
or U1605 (N_1605,N_1577,N_1571);
or U1606 (N_1606,N_1581,N_1568);
nand U1607 (N_1607,N_1566,N_1565);
xor U1608 (N_1608,N_1560,N_1578);
nand U1609 (N_1609,N_1559,N_1557);
nand U1610 (N_1610,N_1594,N_1591);
xnor U1611 (N_1611,N_1572,N_1554);
and U1612 (N_1612,N_1576,N_1597);
or U1613 (N_1613,N_1563,N_1555);
and U1614 (N_1614,N_1595,N_1579);
or U1615 (N_1615,N_1556,N_1553);
nand U1616 (N_1616,N_1590,N_1575);
or U1617 (N_1617,N_1562,N_1587);
or U1618 (N_1618,N_1599,N_1593);
and U1619 (N_1619,N_1580,N_1592);
nor U1620 (N_1620,N_1550,N_1586);
xor U1621 (N_1621,N_1570,N_1583);
and U1622 (N_1622,N_1552,N_1564);
or U1623 (N_1623,N_1574,N_1573);
xor U1624 (N_1624,N_1582,N_1558);
xor U1625 (N_1625,N_1578,N_1550);
or U1626 (N_1626,N_1557,N_1594);
nor U1627 (N_1627,N_1599,N_1597);
nor U1628 (N_1628,N_1588,N_1592);
nand U1629 (N_1629,N_1557,N_1590);
and U1630 (N_1630,N_1589,N_1565);
xor U1631 (N_1631,N_1567,N_1562);
nand U1632 (N_1632,N_1550,N_1582);
xnor U1633 (N_1633,N_1562,N_1574);
nor U1634 (N_1634,N_1556,N_1596);
xnor U1635 (N_1635,N_1554,N_1578);
or U1636 (N_1636,N_1574,N_1595);
nand U1637 (N_1637,N_1579,N_1581);
xnor U1638 (N_1638,N_1550,N_1587);
xor U1639 (N_1639,N_1574,N_1556);
xnor U1640 (N_1640,N_1577,N_1552);
nand U1641 (N_1641,N_1552,N_1578);
nor U1642 (N_1642,N_1570,N_1584);
nand U1643 (N_1643,N_1564,N_1591);
or U1644 (N_1644,N_1565,N_1580);
xnor U1645 (N_1645,N_1559,N_1583);
or U1646 (N_1646,N_1589,N_1553);
nor U1647 (N_1647,N_1590,N_1589);
and U1648 (N_1648,N_1580,N_1585);
or U1649 (N_1649,N_1586,N_1554);
xor U1650 (N_1650,N_1648,N_1607);
nand U1651 (N_1651,N_1639,N_1602);
nand U1652 (N_1652,N_1622,N_1640);
and U1653 (N_1653,N_1633,N_1600);
nor U1654 (N_1654,N_1634,N_1631);
nor U1655 (N_1655,N_1635,N_1620);
or U1656 (N_1656,N_1646,N_1643);
nor U1657 (N_1657,N_1629,N_1644);
nand U1658 (N_1658,N_1604,N_1612);
xnor U1659 (N_1659,N_1606,N_1625);
xnor U1660 (N_1660,N_1645,N_1611);
nor U1661 (N_1661,N_1609,N_1613);
nor U1662 (N_1662,N_1649,N_1610);
or U1663 (N_1663,N_1605,N_1608);
xor U1664 (N_1664,N_1623,N_1616);
nor U1665 (N_1665,N_1619,N_1637);
and U1666 (N_1666,N_1628,N_1632);
or U1667 (N_1667,N_1618,N_1614);
xnor U1668 (N_1668,N_1601,N_1641);
or U1669 (N_1669,N_1627,N_1621);
nand U1670 (N_1670,N_1636,N_1638);
nand U1671 (N_1671,N_1630,N_1647);
xnor U1672 (N_1672,N_1603,N_1624);
and U1673 (N_1673,N_1642,N_1626);
xor U1674 (N_1674,N_1617,N_1615);
nor U1675 (N_1675,N_1622,N_1646);
nor U1676 (N_1676,N_1635,N_1629);
nand U1677 (N_1677,N_1621,N_1626);
nor U1678 (N_1678,N_1644,N_1631);
and U1679 (N_1679,N_1631,N_1636);
nor U1680 (N_1680,N_1647,N_1612);
and U1681 (N_1681,N_1634,N_1628);
nand U1682 (N_1682,N_1632,N_1609);
xor U1683 (N_1683,N_1618,N_1627);
nor U1684 (N_1684,N_1622,N_1615);
nor U1685 (N_1685,N_1609,N_1637);
and U1686 (N_1686,N_1621,N_1602);
nor U1687 (N_1687,N_1605,N_1628);
xor U1688 (N_1688,N_1620,N_1610);
nor U1689 (N_1689,N_1641,N_1605);
nand U1690 (N_1690,N_1607,N_1606);
xor U1691 (N_1691,N_1630,N_1614);
or U1692 (N_1692,N_1638,N_1609);
xnor U1693 (N_1693,N_1627,N_1648);
nand U1694 (N_1694,N_1617,N_1627);
nand U1695 (N_1695,N_1613,N_1634);
nand U1696 (N_1696,N_1610,N_1626);
nor U1697 (N_1697,N_1612,N_1600);
or U1698 (N_1698,N_1634,N_1609);
nor U1699 (N_1699,N_1601,N_1616);
xnor U1700 (N_1700,N_1660,N_1673);
nand U1701 (N_1701,N_1671,N_1664);
nor U1702 (N_1702,N_1668,N_1678);
nor U1703 (N_1703,N_1652,N_1685);
nand U1704 (N_1704,N_1674,N_1667);
nor U1705 (N_1705,N_1654,N_1699);
and U1706 (N_1706,N_1669,N_1680);
xnor U1707 (N_1707,N_1683,N_1679);
or U1708 (N_1708,N_1657,N_1684);
xnor U1709 (N_1709,N_1670,N_1686);
and U1710 (N_1710,N_1697,N_1690);
nor U1711 (N_1711,N_1691,N_1687);
nor U1712 (N_1712,N_1672,N_1677);
nand U1713 (N_1713,N_1675,N_1651);
and U1714 (N_1714,N_1682,N_1658);
nand U1715 (N_1715,N_1666,N_1681);
or U1716 (N_1716,N_1661,N_1698);
nor U1717 (N_1717,N_1655,N_1650);
nor U1718 (N_1718,N_1663,N_1696);
nor U1719 (N_1719,N_1662,N_1688);
or U1720 (N_1720,N_1695,N_1694);
xor U1721 (N_1721,N_1693,N_1692);
or U1722 (N_1722,N_1659,N_1653);
xor U1723 (N_1723,N_1656,N_1689);
nand U1724 (N_1724,N_1665,N_1676);
nor U1725 (N_1725,N_1654,N_1666);
and U1726 (N_1726,N_1685,N_1689);
nor U1727 (N_1727,N_1678,N_1675);
nand U1728 (N_1728,N_1697,N_1656);
nor U1729 (N_1729,N_1660,N_1679);
nand U1730 (N_1730,N_1668,N_1651);
xor U1731 (N_1731,N_1696,N_1651);
and U1732 (N_1732,N_1668,N_1664);
xor U1733 (N_1733,N_1688,N_1660);
or U1734 (N_1734,N_1668,N_1696);
and U1735 (N_1735,N_1662,N_1676);
nand U1736 (N_1736,N_1669,N_1653);
or U1737 (N_1737,N_1673,N_1675);
and U1738 (N_1738,N_1655,N_1652);
nand U1739 (N_1739,N_1667,N_1678);
or U1740 (N_1740,N_1669,N_1662);
xor U1741 (N_1741,N_1689,N_1673);
and U1742 (N_1742,N_1690,N_1665);
xor U1743 (N_1743,N_1680,N_1653);
or U1744 (N_1744,N_1672,N_1697);
nor U1745 (N_1745,N_1679,N_1677);
xnor U1746 (N_1746,N_1669,N_1684);
nand U1747 (N_1747,N_1688,N_1652);
and U1748 (N_1748,N_1680,N_1698);
or U1749 (N_1749,N_1660,N_1681);
nand U1750 (N_1750,N_1740,N_1719);
xor U1751 (N_1751,N_1706,N_1700);
nand U1752 (N_1752,N_1729,N_1711);
or U1753 (N_1753,N_1702,N_1748);
and U1754 (N_1754,N_1744,N_1749);
and U1755 (N_1755,N_1709,N_1745);
nand U1756 (N_1756,N_1732,N_1707);
nor U1757 (N_1757,N_1731,N_1721);
or U1758 (N_1758,N_1722,N_1701);
and U1759 (N_1759,N_1736,N_1746);
nor U1760 (N_1760,N_1718,N_1715);
xor U1761 (N_1761,N_1723,N_1733);
nor U1762 (N_1762,N_1728,N_1743);
nand U1763 (N_1763,N_1704,N_1720);
nor U1764 (N_1764,N_1703,N_1737);
xor U1765 (N_1765,N_1710,N_1717);
xor U1766 (N_1766,N_1742,N_1712);
nor U1767 (N_1767,N_1708,N_1713);
and U1768 (N_1768,N_1730,N_1735);
or U1769 (N_1769,N_1734,N_1738);
xor U1770 (N_1770,N_1741,N_1726);
nand U1771 (N_1771,N_1716,N_1714);
xor U1772 (N_1772,N_1724,N_1725);
xor U1773 (N_1773,N_1747,N_1739);
nand U1774 (N_1774,N_1727,N_1705);
or U1775 (N_1775,N_1721,N_1739);
xnor U1776 (N_1776,N_1723,N_1714);
or U1777 (N_1777,N_1730,N_1703);
and U1778 (N_1778,N_1702,N_1712);
nand U1779 (N_1779,N_1738,N_1746);
nand U1780 (N_1780,N_1726,N_1706);
nor U1781 (N_1781,N_1704,N_1736);
and U1782 (N_1782,N_1732,N_1729);
or U1783 (N_1783,N_1701,N_1719);
nand U1784 (N_1784,N_1704,N_1742);
xor U1785 (N_1785,N_1724,N_1738);
xor U1786 (N_1786,N_1734,N_1726);
and U1787 (N_1787,N_1733,N_1741);
and U1788 (N_1788,N_1717,N_1734);
nor U1789 (N_1789,N_1743,N_1727);
xor U1790 (N_1790,N_1745,N_1726);
nand U1791 (N_1791,N_1748,N_1720);
xor U1792 (N_1792,N_1709,N_1730);
and U1793 (N_1793,N_1745,N_1737);
nand U1794 (N_1794,N_1700,N_1744);
nor U1795 (N_1795,N_1705,N_1729);
or U1796 (N_1796,N_1722,N_1742);
nor U1797 (N_1797,N_1745,N_1732);
or U1798 (N_1798,N_1730,N_1741);
xor U1799 (N_1799,N_1710,N_1728);
or U1800 (N_1800,N_1787,N_1753);
and U1801 (N_1801,N_1776,N_1790);
xor U1802 (N_1802,N_1799,N_1781);
xnor U1803 (N_1803,N_1794,N_1779);
xor U1804 (N_1804,N_1752,N_1784);
xnor U1805 (N_1805,N_1756,N_1778);
xnor U1806 (N_1806,N_1797,N_1755);
nor U1807 (N_1807,N_1767,N_1773);
or U1808 (N_1808,N_1754,N_1777);
and U1809 (N_1809,N_1786,N_1789);
or U1810 (N_1810,N_1795,N_1760);
xnor U1811 (N_1811,N_1780,N_1798);
and U1812 (N_1812,N_1768,N_1775);
and U1813 (N_1813,N_1793,N_1757);
and U1814 (N_1814,N_1766,N_1761);
or U1815 (N_1815,N_1770,N_1764);
xnor U1816 (N_1816,N_1785,N_1791);
or U1817 (N_1817,N_1774,N_1788);
and U1818 (N_1818,N_1782,N_1762);
and U1819 (N_1819,N_1771,N_1769);
xnor U1820 (N_1820,N_1758,N_1759);
xor U1821 (N_1821,N_1751,N_1796);
nand U1822 (N_1822,N_1765,N_1772);
nor U1823 (N_1823,N_1750,N_1763);
xnor U1824 (N_1824,N_1783,N_1792);
nand U1825 (N_1825,N_1785,N_1781);
or U1826 (N_1826,N_1764,N_1755);
and U1827 (N_1827,N_1756,N_1754);
nor U1828 (N_1828,N_1798,N_1784);
nand U1829 (N_1829,N_1798,N_1795);
and U1830 (N_1830,N_1758,N_1767);
xor U1831 (N_1831,N_1783,N_1785);
and U1832 (N_1832,N_1768,N_1777);
xor U1833 (N_1833,N_1768,N_1763);
or U1834 (N_1834,N_1761,N_1765);
or U1835 (N_1835,N_1752,N_1779);
or U1836 (N_1836,N_1765,N_1757);
xnor U1837 (N_1837,N_1784,N_1766);
xor U1838 (N_1838,N_1797,N_1765);
xor U1839 (N_1839,N_1751,N_1790);
or U1840 (N_1840,N_1788,N_1781);
and U1841 (N_1841,N_1763,N_1775);
or U1842 (N_1842,N_1761,N_1769);
xor U1843 (N_1843,N_1796,N_1755);
nand U1844 (N_1844,N_1758,N_1790);
or U1845 (N_1845,N_1780,N_1783);
nor U1846 (N_1846,N_1760,N_1781);
xnor U1847 (N_1847,N_1756,N_1786);
or U1848 (N_1848,N_1754,N_1764);
and U1849 (N_1849,N_1789,N_1793);
or U1850 (N_1850,N_1803,N_1841);
xnor U1851 (N_1851,N_1831,N_1810);
or U1852 (N_1852,N_1827,N_1835);
nor U1853 (N_1853,N_1840,N_1845);
and U1854 (N_1854,N_1817,N_1839);
nand U1855 (N_1855,N_1838,N_1815);
xor U1856 (N_1856,N_1807,N_1836);
xor U1857 (N_1857,N_1809,N_1805);
or U1858 (N_1858,N_1837,N_1808);
and U1859 (N_1859,N_1832,N_1823);
and U1860 (N_1860,N_1818,N_1802);
nor U1861 (N_1861,N_1829,N_1820);
xnor U1862 (N_1862,N_1846,N_1821);
nand U1863 (N_1863,N_1819,N_1804);
or U1864 (N_1864,N_1814,N_1822);
or U1865 (N_1865,N_1800,N_1828);
or U1866 (N_1866,N_1849,N_1843);
nand U1867 (N_1867,N_1825,N_1842);
nor U1868 (N_1868,N_1833,N_1813);
nand U1869 (N_1869,N_1830,N_1847);
or U1870 (N_1870,N_1812,N_1816);
and U1871 (N_1871,N_1801,N_1824);
nor U1872 (N_1872,N_1834,N_1844);
nand U1873 (N_1873,N_1848,N_1826);
and U1874 (N_1874,N_1806,N_1811);
or U1875 (N_1875,N_1839,N_1815);
nand U1876 (N_1876,N_1803,N_1815);
nand U1877 (N_1877,N_1835,N_1810);
xor U1878 (N_1878,N_1840,N_1841);
nor U1879 (N_1879,N_1848,N_1840);
or U1880 (N_1880,N_1816,N_1831);
nand U1881 (N_1881,N_1801,N_1806);
and U1882 (N_1882,N_1834,N_1842);
nand U1883 (N_1883,N_1814,N_1815);
nor U1884 (N_1884,N_1841,N_1848);
or U1885 (N_1885,N_1809,N_1849);
or U1886 (N_1886,N_1832,N_1802);
xnor U1887 (N_1887,N_1849,N_1837);
or U1888 (N_1888,N_1826,N_1840);
nand U1889 (N_1889,N_1812,N_1847);
or U1890 (N_1890,N_1808,N_1806);
or U1891 (N_1891,N_1836,N_1827);
and U1892 (N_1892,N_1804,N_1812);
nor U1893 (N_1893,N_1833,N_1800);
nor U1894 (N_1894,N_1808,N_1843);
or U1895 (N_1895,N_1813,N_1808);
nor U1896 (N_1896,N_1827,N_1822);
and U1897 (N_1897,N_1807,N_1820);
or U1898 (N_1898,N_1812,N_1831);
nand U1899 (N_1899,N_1800,N_1802);
nand U1900 (N_1900,N_1864,N_1889);
and U1901 (N_1901,N_1891,N_1862);
nand U1902 (N_1902,N_1898,N_1887);
and U1903 (N_1903,N_1871,N_1878);
xor U1904 (N_1904,N_1880,N_1875);
xnor U1905 (N_1905,N_1888,N_1857);
xnor U1906 (N_1906,N_1860,N_1856);
nor U1907 (N_1907,N_1884,N_1882);
and U1908 (N_1908,N_1850,N_1852);
xnor U1909 (N_1909,N_1876,N_1853);
xnor U1910 (N_1910,N_1851,N_1883);
nand U1911 (N_1911,N_1865,N_1870);
or U1912 (N_1912,N_1894,N_1861);
xnor U1913 (N_1913,N_1885,N_1879);
xnor U1914 (N_1914,N_1854,N_1881);
xnor U1915 (N_1915,N_1868,N_1866);
nor U1916 (N_1916,N_1874,N_1869);
or U1917 (N_1917,N_1872,N_1892);
nor U1918 (N_1918,N_1896,N_1897);
xnor U1919 (N_1919,N_1858,N_1893);
or U1920 (N_1920,N_1895,N_1867);
nand U1921 (N_1921,N_1877,N_1859);
xnor U1922 (N_1922,N_1873,N_1899);
and U1923 (N_1923,N_1855,N_1890);
xor U1924 (N_1924,N_1886,N_1863);
nand U1925 (N_1925,N_1888,N_1858);
xor U1926 (N_1926,N_1858,N_1866);
nor U1927 (N_1927,N_1875,N_1859);
and U1928 (N_1928,N_1878,N_1886);
or U1929 (N_1929,N_1878,N_1895);
nand U1930 (N_1930,N_1869,N_1853);
xnor U1931 (N_1931,N_1877,N_1875);
nor U1932 (N_1932,N_1887,N_1867);
xor U1933 (N_1933,N_1866,N_1876);
or U1934 (N_1934,N_1895,N_1881);
and U1935 (N_1935,N_1854,N_1885);
and U1936 (N_1936,N_1863,N_1872);
nor U1937 (N_1937,N_1876,N_1889);
nand U1938 (N_1938,N_1879,N_1899);
nor U1939 (N_1939,N_1894,N_1891);
and U1940 (N_1940,N_1885,N_1868);
xor U1941 (N_1941,N_1867,N_1850);
or U1942 (N_1942,N_1851,N_1863);
and U1943 (N_1943,N_1887,N_1878);
nor U1944 (N_1944,N_1868,N_1862);
or U1945 (N_1945,N_1860,N_1859);
nor U1946 (N_1946,N_1889,N_1887);
xnor U1947 (N_1947,N_1850,N_1898);
nor U1948 (N_1948,N_1869,N_1859);
and U1949 (N_1949,N_1885,N_1860);
nor U1950 (N_1950,N_1908,N_1918);
nor U1951 (N_1951,N_1905,N_1941);
or U1952 (N_1952,N_1922,N_1901);
and U1953 (N_1953,N_1930,N_1915);
nand U1954 (N_1954,N_1902,N_1940);
and U1955 (N_1955,N_1900,N_1936);
or U1956 (N_1956,N_1911,N_1927);
nand U1957 (N_1957,N_1933,N_1921);
nand U1958 (N_1958,N_1925,N_1924);
nand U1959 (N_1959,N_1906,N_1907);
nand U1960 (N_1960,N_1935,N_1947);
nand U1961 (N_1961,N_1926,N_1945);
or U1962 (N_1962,N_1928,N_1914);
and U1963 (N_1963,N_1944,N_1917);
and U1964 (N_1964,N_1934,N_1946);
and U1965 (N_1965,N_1904,N_1903);
nor U1966 (N_1966,N_1942,N_1910);
or U1967 (N_1967,N_1923,N_1916);
xor U1968 (N_1968,N_1949,N_1937);
and U1969 (N_1969,N_1932,N_1948);
xnor U1970 (N_1970,N_1919,N_1939);
and U1971 (N_1971,N_1920,N_1909);
nor U1972 (N_1972,N_1938,N_1913);
or U1973 (N_1973,N_1929,N_1931);
nand U1974 (N_1974,N_1912,N_1943);
and U1975 (N_1975,N_1945,N_1928);
and U1976 (N_1976,N_1947,N_1902);
nor U1977 (N_1977,N_1900,N_1931);
xor U1978 (N_1978,N_1925,N_1901);
xor U1979 (N_1979,N_1943,N_1918);
nor U1980 (N_1980,N_1939,N_1935);
and U1981 (N_1981,N_1904,N_1940);
nand U1982 (N_1982,N_1922,N_1905);
xor U1983 (N_1983,N_1929,N_1932);
or U1984 (N_1984,N_1935,N_1933);
nand U1985 (N_1985,N_1905,N_1920);
xor U1986 (N_1986,N_1919,N_1943);
or U1987 (N_1987,N_1936,N_1928);
xor U1988 (N_1988,N_1926,N_1942);
or U1989 (N_1989,N_1924,N_1910);
nand U1990 (N_1990,N_1937,N_1902);
nor U1991 (N_1991,N_1900,N_1943);
or U1992 (N_1992,N_1928,N_1913);
and U1993 (N_1993,N_1914,N_1905);
nand U1994 (N_1994,N_1900,N_1902);
nand U1995 (N_1995,N_1911,N_1918);
xor U1996 (N_1996,N_1902,N_1914);
nand U1997 (N_1997,N_1943,N_1910);
and U1998 (N_1998,N_1919,N_1921);
nor U1999 (N_1999,N_1913,N_1904);
or U2000 (N_2000,N_1956,N_1964);
nor U2001 (N_2001,N_1959,N_1986);
or U2002 (N_2002,N_1996,N_1953);
and U2003 (N_2003,N_1955,N_1991);
and U2004 (N_2004,N_1952,N_1998);
or U2005 (N_2005,N_1975,N_1983);
or U2006 (N_2006,N_1985,N_1988);
or U2007 (N_2007,N_1974,N_1966);
and U2008 (N_2008,N_1982,N_1987);
nand U2009 (N_2009,N_1958,N_1984);
or U2010 (N_2010,N_1970,N_1960);
nand U2011 (N_2011,N_1957,N_1997);
nand U2012 (N_2012,N_1969,N_1981);
nor U2013 (N_2013,N_1951,N_1980);
and U2014 (N_2014,N_1954,N_1999);
nand U2015 (N_2015,N_1963,N_1971);
or U2016 (N_2016,N_1968,N_1979);
and U2017 (N_2017,N_1994,N_1973);
xnor U2018 (N_2018,N_1967,N_1950);
nor U2019 (N_2019,N_1989,N_1992);
xnor U2020 (N_2020,N_1995,N_1972);
or U2021 (N_2021,N_1976,N_1965);
and U2022 (N_2022,N_1978,N_1961);
and U2023 (N_2023,N_1993,N_1977);
or U2024 (N_2024,N_1990,N_1962);
nor U2025 (N_2025,N_1999,N_1958);
and U2026 (N_2026,N_1975,N_1960);
xnor U2027 (N_2027,N_1971,N_1965);
and U2028 (N_2028,N_1952,N_1972);
nand U2029 (N_2029,N_1954,N_1953);
nor U2030 (N_2030,N_1994,N_1962);
and U2031 (N_2031,N_1982,N_1964);
or U2032 (N_2032,N_1993,N_1996);
and U2033 (N_2033,N_1973,N_1953);
xor U2034 (N_2034,N_1961,N_1995);
nor U2035 (N_2035,N_1985,N_1999);
nor U2036 (N_2036,N_1978,N_1977);
and U2037 (N_2037,N_1992,N_1959);
xnor U2038 (N_2038,N_1964,N_1999);
and U2039 (N_2039,N_1964,N_1963);
or U2040 (N_2040,N_1978,N_1968);
nor U2041 (N_2041,N_1951,N_1975);
or U2042 (N_2042,N_1998,N_1973);
nor U2043 (N_2043,N_1963,N_1953);
nor U2044 (N_2044,N_1978,N_1970);
nand U2045 (N_2045,N_1969,N_1961);
nand U2046 (N_2046,N_1977,N_1980);
or U2047 (N_2047,N_1981,N_1973);
and U2048 (N_2048,N_1970,N_1953);
xor U2049 (N_2049,N_1965,N_1960);
or U2050 (N_2050,N_2005,N_2048);
and U2051 (N_2051,N_2036,N_2012);
and U2052 (N_2052,N_2024,N_2003);
nand U2053 (N_2053,N_2023,N_2032);
or U2054 (N_2054,N_2026,N_2037);
and U2055 (N_2055,N_2034,N_2013);
and U2056 (N_2056,N_2014,N_2004);
and U2057 (N_2057,N_2001,N_2010);
nand U2058 (N_2058,N_2018,N_2021);
and U2059 (N_2059,N_2035,N_2002);
and U2060 (N_2060,N_2025,N_2039);
and U2061 (N_2061,N_2047,N_2043);
and U2062 (N_2062,N_2031,N_2015);
nand U2063 (N_2063,N_2016,N_2045);
and U2064 (N_2064,N_2046,N_2022);
or U2065 (N_2065,N_2019,N_2041);
nor U2066 (N_2066,N_2009,N_2017);
xnor U2067 (N_2067,N_2007,N_2049);
nor U2068 (N_2068,N_2040,N_2008);
and U2069 (N_2069,N_2011,N_2038);
nand U2070 (N_2070,N_2020,N_2027);
xor U2071 (N_2071,N_2029,N_2006);
nor U2072 (N_2072,N_2030,N_2000);
and U2073 (N_2073,N_2042,N_2033);
or U2074 (N_2074,N_2028,N_2044);
xnor U2075 (N_2075,N_2025,N_2032);
or U2076 (N_2076,N_2009,N_2047);
and U2077 (N_2077,N_2036,N_2001);
nor U2078 (N_2078,N_2049,N_2027);
nand U2079 (N_2079,N_2039,N_2017);
nand U2080 (N_2080,N_2029,N_2043);
nor U2081 (N_2081,N_2012,N_2042);
nand U2082 (N_2082,N_2001,N_2023);
or U2083 (N_2083,N_2047,N_2028);
nand U2084 (N_2084,N_2002,N_2018);
and U2085 (N_2085,N_2029,N_2038);
and U2086 (N_2086,N_2007,N_2023);
or U2087 (N_2087,N_2026,N_2001);
or U2088 (N_2088,N_2017,N_2027);
and U2089 (N_2089,N_2044,N_2019);
nor U2090 (N_2090,N_2031,N_2048);
nor U2091 (N_2091,N_2030,N_2041);
or U2092 (N_2092,N_2047,N_2013);
xnor U2093 (N_2093,N_2018,N_2030);
nand U2094 (N_2094,N_2004,N_2022);
nand U2095 (N_2095,N_2029,N_2013);
or U2096 (N_2096,N_2003,N_2004);
nand U2097 (N_2097,N_2001,N_2003);
nor U2098 (N_2098,N_2036,N_2019);
nor U2099 (N_2099,N_2022,N_2031);
nand U2100 (N_2100,N_2082,N_2055);
nor U2101 (N_2101,N_2086,N_2057);
or U2102 (N_2102,N_2063,N_2085);
nand U2103 (N_2103,N_2054,N_2098);
xnor U2104 (N_2104,N_2072,N_2095);
or U2105 (N_2105,N_2099,N_2092);
xor U2106 (N_2106,N_2050,N_2076);
or U2107 (N_2107,N_2056,N_2090);
nor U2108 (N_2108,N_2051,N_2087);
nor U2109 (N_2109,N_2073,N_2091);
nand U2110 (N_2110,N_2088,N_2078);
nand U2111 (N_2111,N_2096,N_2080);
xnor U2112 (N_2112,N_2068,N_2061);
xnor U2113 (N_2113,N_2062,N_2067);
nor U2114 (N_2114,N_2066,N_2071);
nor U2115 (N_2115,N_2089,N_2053);
xor U2116 (N_2116,N_2060,N_2081);
and U2117 (N_2117,N_2058,N_2070);
and U2118 (N_2118,N_2059,N_2094);
nand U2119 (N_2119,N_2077,N_2079);
nand U2120 (N_2120,N_2065,N_2052);
nor U2121 (N_2121,N_2084,N_2097);
nand U2122 (N_2122,N_2075,N_2069);
xor U2123 (N_2123,N_2074,N_2093);
nand U2124 (N_2124,N_2083,N_2064);
and U2125 (N_2125,N_2088,N_2093);
xnor U2126 (N_2126,N_2078,N_2074);
nand U2127 (N_2127,N_2053,N_2088);
and U2128 (N_2128,N_2063,N_2090);
or U2129 (N_2129,N_2097,N_2098);
and U2130 (N_2130,N_2079,N_2091);
nor U2131 (N_2131,N_2070,N_2085);
and U2132 (N_2132,N_2060,N_2053);
and U2133 (N_2133,N_2090,N_2086);
xor U2134 (N_2134,N_2063,N_2058);
or U2135 (N_2135,N_2070,N_2081);
nor U2136 (N_2136,N_2099,N_2069);
nand U2137 (N_2137,N_2059,N_2083);
nor U2138 (N_2138,N_2058,N_2098);
xor U2139 (N_2139,N_2095,N_2050);
xnor U2140 (N_2140,N_2083,N_2072);
or U2141 (N_2141,N_2082,N_2073);
nand U2142 (N_2142,N_2057,N_2099);
nand U2143 (N_2143,N_2081,N_2097);
xor U2144 (N_2144,N_2060,N_2080);
and U2145 (N_2145,N_2099,N_2070);
xnor U2146 (N_2146,N_2086,N_2061);
or U2147 (N_2147,N_2080,N_2087);
nand U2148 (N_2148,N_2077,N_2075);
nand U2149 (N_2149,N_2098,N_2084);
xor U2150 (N_2150,N_2110,N_2132);
nand U2151 (N_2151,N_2130,N_2133);
and U2152 (N_2152,N_2129,N_2140);
nor U2153 (N_2153,N_2141,N_2126);
nand U2154 (N_2154,N_2148,N_2121);
or U2155 (N_2155,N_2134,N_2147);
xnor U2156 (N_2156,N_2128,N_2124);
nand U2157 (N_2157,N_2114,N_2109);
or U2158 (N_2158,N_2115,N_2131);
nor U2159 (N_2159,N_2145,N_2100);
nand U2160 (N_2160,N_2106,N_2102);
xnor U2161 (N_2161,N_2127,N_2111);
nor U2162 (N_2162,N_2118,N_2139);
or U2163 (N_2163,N_2122,N_2104);
and U2164 (N_2164,N_2137,N_2149);
nand U2165 (N_2165,N_2123,N_2113);
nand U2166 (N_2166,N_2101,N_2146);
or U2167 (N_2167,N_2144,N_2143);
nor U2168 (N_2168,N_2107,N_2120);
and U2169 (N_2169,N_2116,N_2136);
nand U2170 (N_2170,N_2142,N_2119);
nor U2171 (N_2171,N_2135,N_2103);
and U2172 (N_2172,N_2112,N_2125);
nor U2173 (N_2173,N_2108,N_2105);
or U2174 (N_2174,N_2117,N_2138);
nand U2175 (N_2175,N_2122,N_2124);
or U2176 (N_2176,N_2131,N_2130);
xor U2177 (N_2177,N_2142,N_2146);
or U2178 (N_2178,N_2118,N_2147);
or U2179 (N_2179,N_2104,N_2111);
xor U2180 (N_2180,N_2123,N_2146);
nand U2181 (N_2181,N_2111,N_2102);
and U2182 (N_2182,N_2101,N_2135);
or U2183 (N_2183,N_2113,N_2131);
and U2184 (N_2184,N_2113,N_2132);
or U2185 (N_2185,N_2120,N_2133);
nand U2186 (N_2186,N_2130,N_2116);
and U2187 (N_2187,N_2126,N_2129);
nor U2188 (N_2188,N_2119,N_2103);
and U2189 (N_2189,N_2135,N_2123);
or U2190 (N_2190,N_2146,N_2118);
nand U2191 (N_2191,N_2132,N_2117);
and U2192 (N_2192,N_2121,N_2103);
nor U2193 (N_2193,N_2129,N_2144);
or U2194 (N_2194,N_2122,N_2133);
and U2195 (N_2195,N_2137,N_2100);
and U2196 (N_2196,N_2119,N_2133);
or U2197 (N_2197,N_2118,N_2140);
and U2198 (N_2198,N_2119,N_2116);
nand U2199 (N_2199,N_2132,N_2109);
nor U2200 (N_2200,N_2159,N_2184);
nor U2201 (N_2201,N_2194,N_2152);
nand U2202 (N_2202,N_2186,N_2198);
or U2203 (N_2203,N_2150,N_2189);
nor U2204 (N_2204,N_2182,N_2153);
nor U2205 (N_2205,N_2178,N_2176);
or U2206 (N_2206,N_2174,N_2164);
and U2207 (N_2207,N_2196,N_2165);
and U2208 (N_2208,N_2170,N_2155);
nand U2209 (N_2209,N_2191,N_2181);
nand U2210 (N_2210,N_2163,N_2166);
xnor U2211 (N_2211,N_2160,N_2156);
and U2212 (N_2212,N_2193,N_2188);
xnor U2213 (N_2213,N_2187,N_2179);
or U2214 (N_2214,N_2173,N_2180);
or U2215 (N_2215,N_2151,N_2190);
or U2216 (N_2216,N_2162,N_2172);
or U2217 (N_2217,N_2175,N_2167);
xnor U2218 (N_2218,N_2161,N_2171);
nand U2219 (N_2219,N_2169,N_2185);
or U2220 (N_2220,N_2183,N_2197);
xor U2221 (N_2221,N_2168,N_2195);
or U2222 (N_2222,N_2192,N_2154);
nand U2223 (N_2223,N_2158,N_2199);
nor U2224 (N_2224,N_2157,N_2177);
nand U2225 (N_2225,N_2186,N_2199);
xnor U2226 (N_2226,N_2157,N_2152);
or U2227 (N_2227,N_2193,N_2192);
nor U2228 (N_2228,N_2151,N_2178);
or U2229 (N_2229,N_2167,N_2168);
and U2230 (N_2230,N_2178,N_2181);
or U2231 (N_2231,N_2180,N_2186);
nor U2232 (N_2232,N_2184,N_2154);
xnor U2233 (N_2233,N_2179,N_2165);
xnor U2234 (N_2234,N_2151,N_2162);
and U2235 (N_2235,N_2188,N_2160);
or U2236 (N_2236,N_2182,N_2171);
or U2237 (N_2237,N_2191,N_2174);
nor U2238 (N_2238,N_2190,N_2176);
or U2239 (N_2239,N_2169,N_2162);
or U2240 (N_2240,N_2154,N_2195);
and U2241 (N_2241,N_2167,N_2161);
nand U2242 (N_2242,N_2187,N_2160);
or U2243 (N_2243,N_2151,N_2186);
nor U2244 (N_2244,N_2177,N_2196);
xor U2245 (N_2245,N_2176,N_2195);
and U2246 (N_2246,N_2180,N_2187);
xor U2247 (N_2247,N_2195,N_2190);
and U2248 (N_2248,N_2159,N_2181);
nor U2249 (N_2249,N_2191,N_2189);
nand U2250 (N_2250,N_2223,N_2242);
xor U2251 (N_2251,N_2211,N_2209);
nand U2252 (N_2252,N_2232,N_2220);
nand U2253 (N_2253,N_2218,N_2243);
and U2254 (N_2254,N_2230,N_2226);
nor U2255 (N_2255,N_2241,N_2236);
xnor U2256 (N_2256,N_2216,N_2219);
nor U2257 (N_2257,N_2217,N_2207);
nand U2258 (N_2258,N_2202,N_2231);
nand U2259 (N_2259,N_2245,N_2206);
or U2260 (N_2260,N_2248,N_2214);
or U2261 (N_2261,N_2208,N_2237);
nand U2262 (N_2262,N_2249,N_2224);
nand U2263 (N_2263,N_2239,N_2221);
nand U2264 (N_2264,N_2212,N_2228);
nand U2265 (N_2265,N_2215,N_2229);
and U2266 (N_2266,N_2204,N_2205);
nor U2267 (N_2267,N_2238,N_2201);
nand U2268 (N_2268,N_2233,N_2200);
or U2269 (N_2269,N_2203,N_2227);
or U2270 (N_2270,N_2225,N_2234);
nand U2271 (N_2271,N_2222,N_2210);
or U2272 (N_2272,N_2235,N_2246);
or U2273 (N_2273,N_2240,N_2213);
nand U2274 (N_2274,N_2244,N_2247);
nand U2275 (N_2275,N_2244,N_2234);
xnor U2276 (N_2276,N_2236,N_2219);
xnor U2277 (N_2277,N_2225,N_2210);
nand U2278 (N_2278,N_2214,N_2241);
nor U2279 (N_2279,N_2233,N_2208);
and U2280 (N_2280,N_2234,N_2246);
xor U2281 (N_2281,N_2200,N_2249);
xor U2282 (N_2282,N_2229,N_2238);
xnor U2283 (N_2283,N_2225,N_2244);
nor U2284 (N_2284,N_2207,N_2212);
xnor U2285 (N_2285,N_2238,N_2218);
or U2286 (N_2286,N_2238,N_2233);
and U2287 (N_2287,N_2203,N_2200);
xor U2288 (N_2288,N_2203,N_2243);
and U2289 (N_2289,N_2247,N_2211);
nand U2290 (N_2290,N_2201,N_2214);
and U2291 (N_2291,N_2245,N_2200);
xor U2292 (N_2292,N_2240,N_2202);
nor U2293 (N_2293,N_2203,N_2207);
nor U2294 (N_2294,N_2238,N_2223);
or U2295 (N_2295,N_2238,N_2216);
and U2296 (N_2296,N_2226,N_2212);
nor U2297 (N_2297,N_2204,N_2237);
nor U2298 (N_2298,N_2244,N_2215);
and U2299 (N_2299,N_2219,N_2221);
xor U2300 (N_2300,N_2263,N_2259);
and U2301 (N_2301,N_2255,N_2287);
or U2302 (N_2302,N_2277,N_2256);
nor U2303 (N_2303,N_2260,N_2262);
or U2304 (N_2304,N_2295,N_2288);
and U2305 (N_2305,N_2285,N_2286);
or U2306 (N_2306,N_2281,N_2250);
xor U2307 (N_2307,N_2269,N_2273);
and U2308 (N_2308,N_2294,N_2278);
or U2309 (N_2309,N_2275,N_2251);
xnor U2310 (N_2310,N_2290,N_2258);
nand U2311 (N_2311,N_2267,N_2266);
nand U2312 (N_2312,N_2265,N_2270);
nand U2313 (N_2313,N_2283,N_2271);
and U2314 (N_2314,N_2293,N_2284);
nor U2315 (N_2315,N_2298,N_2252);
xor U2316 (N_2316,N_2274,N_2292);
or U2317 (N_2317,N_2264,N_2261);
and U2318 (N_2318,N_2280,N_2276);
nor U2319 (N_2319,N_2299,N_2289);
nor U2320 (N_2320,N_2257,N_2268);
or U2321 (N_2321,N_2254,N_2272);
nand U2322 (N_2322,N_2297,N_2291);
xnor U2323 (N_2323,N_2296,N_2279);
xor U2324 (N_2324,N_2282,N_2253);
xor U2325 (N_2325,N_2266,N_2275);
or U2326 (N_2326,N_2273,N_2290);
or U2327 (N_2327,N_2272,N_2260);
nand U2328 (N_2328,N_2257,N_2270);
and U2329 (N_2329,N_2277,N_2267);
xnor U2330 (N_2330,N_2264,N_2263);
nand U2331 (N_2331,N_2292,N_2283);
xor U2332 (N_2332,N_2292,N_2285);
nand U2333 (N_2333,N_2293,N_2274);
and U2334 (N_2334,N_2298,N_2291);
nor U2335 (N_2335,N_2263,N_2279);
and U2336 (N_2336,N_2270,N_2287);
nor U2337 (N_2337,N_2254,N_2266);
nor U2338 (N_2338,N_2271,N_2274);
or U2339 (N_2339,N_2299,N_2261);
xor U2340 (N_2340,N_2270,N_2289);
or U2341 (N_2341,N_2275,N_2281);
and U2342 (N_2342,N_2254,N_2268);
xor U2343 (N_2343,N_2269,N_2284);
or U2344 (N_2344,N_2282,N_2264);
or U2345 (N_2345,N_2257,N_2287);
xnor U2346 (N_2346,N_2250,N_2288);
or U2347 (N_2347,N_2293,N_2258);
nor U2348 (N_2348,N_2250,N_2283);
nor U2349 (N_2349,N_2265,N_2290);
nor U2350 (N_2350,N_2306,N_2314);
nor U2351 (N_2351,N_2325,N_2332);
nand U2352 (N_2352,N_2313,N_2345);
nor U2353 (N_2353,N_2315,N_2304);
nand U2354 (N_2354,N_2303,N_2309);
and U2355 (N_2355,N_2347,N_2318);
xnor U2356 (N_2356,N_2317,N_2312);
xor U2357 (N_2357,N_2348,N_2327);
nor U2358 (N_2358,N_2336,N_2322);
nor U2359 (N_2359,N_2335,N_2320);
nand U2360 (N_2360,N_2324,N_2339);
or U2361 (N_2361,N_2307,N_2334);
nand U2362 (N_2362,N_2337,N_2300);
xor U2363 (N_2363,N_2344,N_2338);
xor U2364 (N_2364,N_2305,N_2328);
and U2365 (N_2365,N_2342,N_2329);
or U2366 (N_2366,N_2323,N_2321);
xor U2367 (N_2367,N_2331,N_2341);
and U2368 (N_2368,N_2316,N_2308);
nand U2369 (N_2369,N_2333,N_2319);
or U2370 (N_2370,N_2330,N_2310);
xor U2371 (N_2371,N_2340,N_2302);
xor U2372 (N_2372,N_2311,N_2343);
nor U2373 (N_2373,N_2301,N_2349);
or U2374 (N_2374,N_2346,N_2326);
xnor U2375 (N_2375,N_2332,N_2342);
or U2376 (N_2376,N_2306,N_2308);
and U2377 (N_2377,N_2338,N_2347);
nand U2378 (N_2378,N_2311,N_2322);
nand U2379 (N_2379,N_2344,N_2320);
and U2380 (N_2380,N_2315,N_2309);
or U2381 (N_2381,N_2331,N_2330);
or U2382 (N_2382,N_2300,N_2317);
or U2383 (N_2383,N_2310,N_2322);
nand U2384 (N_2384,N_2320,N_2300);
xnor U2385 (N_2385,N_2338,N_2305);
xnor U2386 (N_2386,N_2321,N_2335);
nor U2387 (N_2387,N_2316,N_2344);
and U2388 (N_2388,N_2349,N_2333);
nor U2389 (N_2389,N_2304,N_2335);
nand U2390 (N_2390,N_2321,N_2340);
xnor U2391 (N_2391,N_2339,N_2347);
xnor U2392 (N_2392,N_2305,N_2341);
and U2393 (N_2393,N_2326,N_2300);
and U2394 (N_2394,N_2330,N_2314);
xor U2395 (N_2395,N_2325,N_2339);
xor U2396 (N_2396,N_2305,N_2345);
nor U2397 (N_2397,N_2341,N_2313);
or U2398 (N_2398,N_2326,N_2335);
nor U2399 (N_2399,N_2334,N_2333);
or U2400 (N_2400,N_2372,N_2395);
nand U2401 (N_2401,N_2358,N_2354);
and U2402 (N_2402,N_2382,N_2397);
and U2403 (N_2403,N_2384,N_2385);
nor U2404 (N_2404,N_2377,N_2398);
xnor U2405 (N_2405,N_2374,N_2391);
or U2406 (N_2406,N_2350,N_2386);
nand U2407 (N_2407,N_2383,N_2376);
nand U2408 (N_2408,N_2380,N_2363);
and U2409 (N_2409,N_2373,N_2378);
nor U2410 (N_2410,N_2392,N_2366);
nor U2411 (N_2411,N_2356,N_2361);
nand U2412 (N_2412,N_2351,N_2362);
and U2413 (N_2413,N_2371,N_2352);
nand U2414 (N_2414,N_2393,N_2394);
and U2415 (N_2415,N_2387,N_2390);
and U2416 (N_2416,N_2379,N_2396);
or U2417 (N_2417,N_2367,N_2375);
or U2418 (N_2418,N_2357,N_2389);
xnor U2419 (N_2419,N_2369,N_2381);
xor U2420 (N_2420,N_2353,N_2368);
nand U2421 (N_2421,N_2364,N_2399);
or U2422 (N_2422,N_2355,N_2359);
nor U2423 (N_2423,N_2370,N_2360);
xnor U2424 (N_2424,N_2388,N_2365);
and U2425 (N_2425,N_2351,N_2395);
or U2426 (N_2426,N_2370,N_2380);
nand U2427 (N_2427,N_2368,N_2360);
nor U2428 (N_2428,N_2352,N_2373);
and U2429 (N_2429,N_2394,N_2385);
xor U2430 (N_2430,N_2376,N_2398);
nand U2431 (N_2431,N_2376,N_2393);
nor U2432 (N_2432,N_2371,N_2364);
nand U2433 (N_2433,N_2353,N_2352);
nand U2434 (N_2434,N_2350,N_2365);
nand U2435 (N_2435,N_2356,N_2396);
or U2436 (N_2436,N_2353,N_2398);
and U2437 (N_2437,N_2351,N_2357);
nand U2438 (N_2438,N_2387,N_2350);
nor U2439 (N_2439,N_2363,N_2361);
and U2440 (N_2440,N_2385,N_2351);
and U2441 (N_2441,N_2384,N_2356);
xnor U2442 (N_2442,N_2359,N_2374);
xnor U2443 (N_2443,N_2381,N_2372);
and U2444 (N_2444,N_2392,N_2351);
nor U2445 (N_2445,N_2368,N_2396);
and U2446 (N_2446,N_2387,N_2396);
or U2447 (N_2447,N_2350,N_2362);
and U2448 (N_2448,N_2369,N_2356);
and U2449 (N_2449,N_2377,N_2389);
nand U2450 (N_2450,N_2404,N_2431);
nand U2451 (N_2451,N_2425,N_2408);
and U2452 (N_2452,N_2407,N_2416);
xor U2453 (N_2453,N_2436,N_2441);
and U2454 (N_2454,N_2420,N_2443);
and U2455 (N_2455,N_2422,N_2402);
xnor U2456 (N_2456,N_2411,N_2435);
nand U2457 (N_2457,N_2406,N_2446);
nand U2458 (N_2458,N_2413,N_2414);
and U2459 (N_2459,N_2403,N_2417);
nor U2460 (N_2460,N_2427,N_2419);
xnor U2461 (N_2461,N_2426,N_2440);
xor U2462 (N_2462,N_2409,N_2432);
and U2463 (N_2463,N_2405,N_2434);
xnor U2464 (N_2464,N_2438,N_2448);
xor U2465 (N_2465,N_2421,N_2444);
nand U2466 (N_2466,N_2415,N_2449);
or U2467 (N_2467,N_2428,N_2401);
xor U2468 (N_2468,N_2412,N_2410);
or U2469 (N_2469,N_2433,N_2400);
xor U2470 (N_2470,N_2429,N_2445);
and U2471 (N_2471,N_2442,N_2418);
nand U2472 (N_2472,N_2430,N_2424);
nand U2473 (N_2473,N_2447,N_2439);
xor U2474 (N_2474,N_2437,N_2423);
nor U2475 (N_2475,N_2430,N_2407);
nor U2476 (N_2476,N_2402,N_2430);
xnor U2477 (N_2477,N_2419,N_2412);
nor U2478 (N_2478,N_2412,N_2406);
xnor U2479 (N_2479,N_2441,N_2438);
or U2480 (N_2480,N_2444,N_2443);
xnor U2481 (N_2481,N_2413,N_2412);
or U2482 (N_2482,N_2417,N_2401);
and U2483 (N_2483,N_2439,N_2410);
nand U2484 (N_2484,N_2440,N_2400);
nand U2485 (N_2485,N_2403,N_2439);
nor U2486 (N_2486,N_2409,N_2404);
nand U2487 (N_2487,N_2403,N_2424);
or U2488 (N_2488,N_2422,N_2434);
or U2489 (N_2489,N_2407,N_2449);
nand U2490 (N_2490,N_2420,N_2409);
nand U2491 (N_2491,N_2443,N_2431);
and U2492 (N_2492,N_2431,N_2438);
or U2493 (N_2493,N_2428,N_2425);
or U2494 (N_2494,N_2427,N_2433);
xnor U2495 (N_2495,N_2449,N_2446);
and U2496 (N_2496,N_2407,N_2433);
xor U2497 (N_2497,N_2407,N_2440);
nor U2498 (N_2498,N_2446,N_2444);
xnor U2499 (N_2499,N_2433,N_2447);
xor U2500 (N_2500,N_2492,N_2475);
and U2501 (N_2501,N_2483,N_2462);
nor U2502 (N_2502,N_2456,N_2460);
or U2503 (N_2503,N_2489,N_2454);
and U2504 (N_2504,N_2490,N_2472);
and U2505 (N_2505,N_2477,N_2493);
xor U2506 (N_2506,N_2453,N_2468);
nand U2507 (N_2507,N_2496,N_2458);
nor U2508 (N_2508,N_2457,N_2473);
xor U2509 (N_2509,N_2476,N_2495);
nand U2510 (N_2510,N_2471,N_2499);
nand U2511 (N_2511,N_2469,N_2479);
nand U2512 (N_2512,N_2467,N_2474);
nor U2513 (N_2513,N_2452,N_2481);
or U2514 (N_2514,N_2494,N_2498);
and U2515 (N_2515,N_2480,N_2466);
and U2516 (N_2516,N_2488,N_2486);
nand U2517 (N_2517,N_2455,N_2484);
or U2518 (N_2518,N_2470,N_2450);
nand U2519 (N_2519,N_2465,N_2451);
nand U2520 (N_2520,N_2497,N_2482);
nor U2521 (N_2521,N_2464,N_2485);
or U2522 (N_2522,N_2491,N_2478);
and U2523 (N_2523,N_2459,N_2461);
nor U2524 (N_2524,N_2487,N_2463);
nand U2525 (N_2525,N_2497,N_2473);
xor U2526 (N_2526,N_2451,N_2491);
or U2527 (N_2527,N_2493,N_2452);
or U2528 (N_2528,N_2476,N_2497);
or U2529 (N_2529,N_2465,N_2461);
nand U2530 (N_2530,N_2464,N_2483);
nor U2531 (N_2531,N_2498,N_2458);
nand U2532 (N_2532,N_2472,N_2484);
and U2533 (N_2533,N_2472,N_2488);
or U2534 (N_2534,N_2491,N_2498);
xor U2535 (N_2535,N_2465,N_2470);
nand U2536 (N_2536,N_2481,N_2461);
nand U2537 (N_2537,N_2493,N_2475);
nand U2538 (N_2538,N_2466,N_2457);
xnor U2539 (N_2539,N_2456,N_2499);
nand U2540 (N_2540,N_2491,N_2485);
nand U2541 (N_2541,N_2453,N_2470);
or U2542 (N_2542,N_2484,N_2494);
nor U2543 (N_2543,N_2454,N_2460);
and U2544 (N_2544,N_2452,N_2494);
nor U2545 (N_2545,N_2470,N_2472);
or U2546 (N_2546,N_2453,N_2496);
nor U2547 (N_2547,N_2498,N_2481);
nor U2548 (N_2548,N_2492,N_2464);
nor U2549 (N_2549,N_2465,N_2482);
or U2550 (N_2550,N_2511,N_2505);
or U2551 (N_2551,N_2523,N_2517);
nand U2552 (N_2552,N_2503,N_2512);
or U2553 (N_2553,N_2518,N_2526);
and U2554 (N_2554,N_2538,N_2540);
and U2555 (N_2555,N_2546,N_2501);
xnor U2556 (N_2556,N_2529,N_2530);
nor U2557 (N_2557,N_2504,N_2537);
nor U2558 (N_2558,N_2535,N_2507);
nor U2559 (N_2559,N_2539,N_2532);
or U2560 (N_2560,N_2508,N_2548);
nor U2561 (N_2561,N_2534,N_2544);
nand U2562 (N_2562,N_2513,N_2510);
nand U2563 (N_2563,N_2545,N_2500);
xor U2564 (N_2564,N_2520,N_2533);
nand U2565 (N_2565,N_2543,N_2527);
or U2566 (N_2566,N_2515,N_2542);
nor U2567 (N_2567,N_2506,N_2519);
and U2568 (N_2568,N_2502,N_2509);
nor U2569 (N_2569,N_2536,N_2541);
xor U2570 (N_2570,N_2524,N_2516);
nand U2571 (N_2571,N_2521,N_2549);
or U2572 (N_2572,N_2522,N_2531);
nand U2573 (N_2573,N_2528,N_2514);
and U2574 (N_2574,N_2547,N_2525);
nand U2575 (N_2575,N_2516,N_2510);
xnor U2576 (N_2576,N_2531,N_2534);
nand U2577 (N_2577,N_2506,N_2527);
or U2578 (N_2578,N_2518,N_2547);
and U2579 (N_2579,N_2530,N_2528);
xnor U2580 (N_2580,N_2511,N_2548);
nor U2581 (N_2581,N_2514,N_2541);
nand U2582 (N_2582,N_2532,N_2525);
and U2583 (N_2583,N_2528,N_2548);
nor U2584 (N_2584,N_2518,N_2500);
xor U2585 (N_2585,N_2528,N_2532);
and U2586 (N_2586,N_2538,N_2524);
or U2587 (N_2587,N_2502,N_2528);
or U2588 (N_2588,N_2549,N_2505);
nor U2589 (N_2589,N_2547,N_2515);
nor U2590 (N_2590,N_2501,N_2529);
or U2591 (N_2591,N_2535,N_2521);
xnor U2592 (N_2592,N_2505,N_2529);
or U2593 (N_2593,N_2512,N_2509);
nor U2594 (N_2594,N_2535,N_2538);
or U2595 (N_2595,N_2517,N_2511);
nor U2596 (N_2596,N_2516,N_2500);
and U2597 (N_2597,N_2523,N_2525);
nor U2598 (N_2598,N_2542,N_2502);
nand U2599 (N_2599,N_2502,N_2507);
and U2600 (N_2600,N_2587,N_2559);
nor U2601 (N_2601,N_2562,N_2588);
and U2602 (N_2602,N_2554,N_2590);
nand U2603 (N_2603,N_2566,N_2592);
nor U2604 (N_2604,N_2599,N_2581);
or U2605 (N_2605,N_2596,N_2574);
nand U2606 (N_2606,N_2573,N_2576);
and U2607 (N_2607,N_2580,N_2572);
nor U2608 (N_2608,N_2567,N_2575);
or U2609 (N_2609,N_2594,N_2593);
nand U2610 (N_2610,N_2579,N_2595);
xor U2611 (N_2611,N_2564,N_2582);
or U2612 (N_2612,N_2583,N_2569);
xnor U2613 (N_2613,N_2585,N_2584);
nand U2614 (N_2614,N_2560,N_2558);
nand U2615 (N_2615,N_2597,N_2550);
or U2616 (N_2616,N_2577,N_2563);
nand U2617 (N_2617,N_2570,N_2557);
xor U2618 (N_2618,N_2565,N_2561);
or U2619 (N_2619,N_2589,N_2551);
xor U2620 (N_2620,N_2556,N_2568);
or U2621 (N_2621,N_2555,N_2578);
nand U2622 (N_2622,N_2586,N_2598);
xor U2623 (N_2623,N_2591,N_2571);
xnor U2624 (N_2624,N_2552,N_2553);
or U2625 (N_2625,N_2564,N_2598);
nand U2626 (N_2626,N_2596,N_2599);
nor U2627 (N_2627,N_2552,N_2569);
nor U2628 (N_2628,N_2595,N_2568);
xor U2629 (N_2629,N_2582,N_2588);
nand U2630 (N_2630,N_2588,N_2555);
xor U2631 (N_2631,N_2560,N_2567);
nand U2632 (N_2632,N_2560,N_2571);
or U2633 (N_2633,N_2588,N_2596);
xnor U2634 (N_2634,N_2570,N_2593);
nor U2635 (N_2635,N_2563,N_2564);
or U2636 (N_2636,N_2551,N_2584);
nor U2637 (N_2637,N_2588,N_2583);
xor U2638 (N_2638,N_2588,N_2593);
nand U2639 (N_2639,N_2551,N_2575);
and U2640 (N_2640,N_2564,N_2556);
xnor U2641 (N_2641,N_2577,N_2559);
nor U2642 (N_2642,N_2555,N_2574);
nand U2643 (N_2643,N_2568,N_2583);
nand U2644 (N_2644,N_2571,N_2557);
xor U2645 (N_2645,N_2567,N_2591);
or U2646 (N_2646,N_2558,N_2583);
and U2647 (N_2647,N_2561,N_2574);
nor U2648 (N_2648,N_2580,N_2557);
or U2649 (N_2649,N_2571,N_2587);
nand U2650 (N_2650,N_2610,N_2646);
and U2651 (N_2651,N_2608,N_2631);
nand U2652 (N_2652,N_2603,N_2606);
and U2653 (N_2653,N_2627,N_2607);
and U2654 (N_2654,N_2619,N_2625);
nor U2655 (N_2655,N_2616,N_2602);
nor U2656 (N_2656,N_2613,N_2600);
nand U2657 (N_2657,N_2649,N_2624);
xnor U2658 (N_2658,N_2609,N_2637);
nand U2659 (N_2659,N_2642,N_2643);
nor U2660 (N_2660,N_2621,N_2611);
nand U2661 (N_2661,N_2622,N_2620);
or U2662 (N_2662,N_2617,N_2618);
nor U2663 (N_2663,N_2629,N_2615);
nand U2664 (N_2664,N_2630,N_2628);
nand U2665 (N_2665,N_2647,N_2604);
or U2666 (N_2666,N_2614,N_2626);
and U2667 (N_2667,N_2623,N_2605);
and U2668 (N_2668,N_2633,N_2640);
and U2669 (N_2669,N_2612,N_2636);
or U2670 (N_2670,N_2632,N_2635);
nor U2671 (N_2671,N_2645,N_2601);
or U2672 (N_2672,N_2634,N_2644);
nor U2673 (N_2673,N_2641,N_2638);
or U2674 (N_2674,N_2648,N_2639);
nand U2675 (N_2675,N_2624,N_2645);
nor U2676 (N_2676,N_2619,N_2607);
nor U2677 (N_2677,N_2606,N_2621);
nor U2678 (N_2678,N_2616,N_2631);
or U2679 (N_2679,N_2622,N_2639);
nand U2680 (N_2680,N_2642,N_2601);
or U2681 (N_2681,N_2621,N_2639);
xor U2682 (N_2682,N_2648,N_2640);
xnor U2683 (N_2683,N_2612,N_2610);
nand U2684 (N_2684,N_2643,N_2618);
and U2685 (N_2685,N_2617,N_2641);
and U2686 (N_2686,N_2646,N_2611);
and U2687 (N_2687,N_2610,N_2637);
or U2688 (N_2688,N_2618,N_2634);
xnor U2689 (N_2689,N_2643,N_2626);
nor U2690 (N_2690,N_2638,N_2625);
or U2691 (N_2691,N_2624,N_2600);
or U2692 (N_2692,N_2602,N_2644);
nand U2693 (N_2693,N_2619,N_2635);
and U2694 (N_2694,N_2601,N_2644);
xnor U2695 (N_2695,N_2608,N_2606);
nor U2696 (N_2696,N_2623,N_2620);
nor U2697 (N_2697,N_2634,N_2611);
and U2698 (N_2698,N_2624,N_2623);
nor U2699 (N_2699,N_2638,N_2607);
or U2700 (N_2700,N_2658,N_2651);
or U2701 (N_2701,N_2668,N_2671);
nor U2702 (N_2702,N_2690,N_2663);
nor U2703 (N_2703,N_2659,N_2664);
or U2704 (N_2704,N_2652,N_2669);
nor U2705 (N_2705,N_2660,N_2654);
nor U2706 (N_2706,N_2695,N_2675);
xor U2707 (N_2707,N_2650,N_2678);
and U2708 (N_2708,N_2662,N_2673);
nand U2709 (N_2709,N_2665,N_2666);
nor U2710 (N_2710,N_2676,N_2653);
xnor U2711 (N_2711,N_2657,N_2688);
xor U2712 (N_2712,N_2681,N_2670);
and U2713 (N_2713,N_2697,N_2686);
or U2714 (N_2714,N_2674,N_2687);
or U2715 (N_2715,N_2667,N_2682);
xor U2716 (N_2716,N_2698,N_2679);
nand U2717 (N_2717,N_2685,N_2689);
nand U2718 (N_2718,N_2656,N_2677);
xnor U2719 (N_2719,N_2684,N_2680);
nor U2720 (N_2720,N_2693,N_2694);
or U2721 (N_2721,N_2699,N_2683);
nand U2722 (N_2722,N_2661,N_2692);
nor U2723 (N_2723,N_2696,N_2672);
or U2724 (N_2724,N_2691,N_2655);
xnor U2725 (N_2725,N_2655,N_2677);
and U2726 (N_2726,N_2650,N_2676);
xnor U2727 (N_2727,N_2683,N_2654);
xnor U2728 (N_2728,N_2667,N_2693);
nand U2729 (N_2729,N_2675,N_2666);
nand U2730 (N_2730,N_2657,N_2673);
or U2731 (N_2731,N_2697,N_2696);
nand U2732 (N_2732,N_2696,N_2677);
xor U2733 (N_2733,N_2688,N_2653);
nor U2734 (N_2734,N_2662,N_2656);
or U2735 (N_2735,N_2651,N_2650);
nor U2736 (N_2736,N_2668,N_2655);
and U2737 (N_2737,N_2687,N_2665);
or U2738 (N_2738,N_2683,N_2659);
nand U2739 (N_2739,N_2686,N_2696);
nand U2740 (N_2740,N_2673,N_2695);
xor U2741 (N_2741,N_2672,N_2671);
or U2742 (N_2742,N_2661,N_2656);
nand U2743 (N_2743,N_2696,N_2692);
xnor U2744 (N_2744,N_2662,N_2660);
and U2745 (N_2745,N_2689,N_2661);
xnor U2746 (N_2746,N_2688,N_2669);
and U2747 (N_2747,N_2684,N_2698);
xor U2748 (N_2748,N_2688,N_2650);
and U2749 (N_2749,N_2665,N_2698);
xor U2750 (N_2750,N_2737,N_2709);
and U2751 (N_2751,N_2700,N_2718);
xnor U2752 (N_2752,N_2726,N_2706);
nor U2753 (N_2753,N_2704,N_2707);
or U2754 (N_2754,N_2749,N_2730);
xor U2755 (N_2755,N_2733,N_2705);
or U2756 (N_2756,N_2715,N_2717);
or U2757 (N_2757,N_2713,N_2746);
or U2758 (N_2758,N_2745,N_2719);
nor U2759 (N_2759,N_2723,N_2724);
or U2760 (N_2760,N_2741,N_2734);
nand U2761 (N_2761,N_2729,N_2736);
and U2762 (N_2762,N_2728,N_2727);
nand U2763 (N_2763,N_2735,N_2711);
nor U2764 (N_2764,N_2716,N_2702);
or U2765 (N_2765,N_2738,N_2731);
or U2766 (N_2766,N_2701,N_2744);
nor U2767 (N_2767,N_2703,N_2742);
or U2768 (N_2768,N_2725,N_2743);
nand U2769 (N_2769,N_2720,N_2712);
xnor U2770 (N_2770,N_2710,N_2739);
nor U2771 (N_2771,N_2732,N_2708);
or U2772 (N_2772,N_2721,N_2747);
nor U2773 (N_2773,N_2740,N_2722);
xor U2774 (N_2774,N_2748,N_2714);
nand U2775 (N_2775,N_2716,N_2707);
nand U2776 (N_2776,N_2742,N_2745);
xor U2777 (N_2777,N_2735,N_2742);
and U2778 (N_2778,N_2736,N_2748);
xnor U2779 (N_2779,N_2704,N_2705);
nand U2780 (N_2780,N_2741,N_2731);
or U2781 (N_2781,N_2718,N_2736);
xnor U2782 (N_2782,N_2744,N_2733);
nand U2783 (N_2783,N_2700,N_2724);
xnor U2784 (N_2784,N_2749,N_2729);
xnor U2785 (N_2785,N_2731,N_2748);
and U2786 (N_2786,N_2734,N_2713);
nor U2787 (N_2787,N_2711,N_2709);
nand U2788 (N_2788,N_2737,N_2740);
nand U2789 (N_2789,N_2728,N_2706);
nand U2790 (N_2790,N_2724,N_2729);
or U2791 (N_2791,N_2708,N_2702);
nand U2792 (N_2792,N_2738,N_2717);
xor U2793 (N_2793,N_2728,N_2715);
xor U2794 (N_2794,N_2718,N_2748);
nor U2795 (N_2795,N_2721,N_2742);
and U2796 (N_2796,N_2720,N_2711);
nor U2797 (N_2797,N_2728,N_2711);
or U2798 (N_2798,N_2709,N_2730);
or U2799 (N_2799,N_2736,N_2743);
or U2800 (N_2800,N_2792,N_2750);
and U2801 (N_2801,N_2760,N_2795);
xnor U2802 (N_2802,N_2784,N_2791);
or U2803 (N_2803,N_2753,N_2769);
nand U2804 (N_2804,N_2752,N_2794);
nor U2805 (N_2805,N_2770,N_2767);
xnor U2806 (N_2806,N_2786,N_2758);
or U2807 (N_2807,N_2763,N_2765);
nand U2808 (N_2808,N_2782,N_2790);
and U2809 (N_2809,N_2772,N_2796);
and U2810 (N_2810,N_2779,N_2777);
and U2811 (N_2811,N_2799,N_2762);
or U2812 (N_2812,N_2771,N_2783);
and U2813 (N_2813,N_2781,N_2793);
nand U2814 (N_2814,N_2776,N_2788);
xnor U2815 (N_2815,N_2798,N_2773);
nor U2816 (N_2816,N_2751,N_2774);
nand U2817 (N_2817,N_2755,N_2756);
nor U2818 (N_2818,N_2754,N_2768);
nand U2819 (N_2819,N_2766,N_2775);
nor U2820 (N_2820,N_2757,N_2797);
or U2821 (N_2821,N_2780,N_2759);
xnor U2822 (N_2822,N_2764,N_2787);
nand U2823 (N_2823,N_2778,N_2789);
nand U2824 (N_2824,N_2785,N_2761);
xor U2825 (N_2825,N_2750,N_2783);
nor U2826 (N_2826,N_2799,N_2773);
nand U2827 (N_2827,N_2754,N_2762);
nand U2828 (N_2828,N_2776,N_2761);
or U2829 (N_2829,N_2795,N_2790);
nand U2830 (N_2830,N_2786,N_2763);
nand U2831 (N_2831,N_2783,N_2793);
xor U2832 (N_2832,N_2771,N_2777);
nor U2833 (N_2833,N_2764,N_2763);
and U2834 (N_2834,N_2777,N_2757);
or U2835 (N_2835,N_2795,N_2778);
or U2836 (N_2836,N_2792,N_2782);
nor U2837 (N_2837,N_2764,N_2794);
nor U2838 (N_2838,N_2792,N_2775);
or U2839 (N_2839,N_2782,N_2775);
xor U2840 (N_2840,N_2763,N_2778);
and U2841 (N_2841,N_2761,N_2791);
or U2842 (N_2842,N_2791,N_2771);
and U2843 (N_2843,N_2751,N_2768);
nor U2844 (N_2844,N_2769,N_2788);
or U2845 (N_2845,N_2781,N_2792);
xor U2846 (N_2846,N_2799,N_2775);
xnor U2847 (N_2847,N_2788,N_2755);
xnor U2848 (N_2848,N_2783,N_2797);
nor U2849 (N_2849,N_2754,N_2785);
and U2850 (N_2850,N_2803,N_2838);
xnor U2851 (N_2851,N_2828,N_2801);
xnor U2852 (N_2852,N_2844,N_2819);
nor U2853 (N_2853,N_2847,N_2826);
xnor U2854 (N_2854,N_2811,N_2815);
and U2855 (N_2855,N_2800,N_2813);
or U2856 (N_2856,N_2802,N_2806);
nor U2857 (N_2857,N_2824,N_2830);
xor U2858 (N_2858,N_2841,N_2842);
or U2859 (N_2859,N_2845,N_2817);
nand U2860 (N_2860,N_2833,N_2807);
and U2861 (N_2861,N_2810,N_2829);
xor U2862 (N_2862,N_2834,N_2814);
nand U2863 (N_2863,N_2809,N_2827);
nor U2864 (N_2864,N_2846,N_2818);
nand U2865 (N_2865,N_2804,N_2825);
and U2866 (N_2866,N_2823,N_2816);
nor U2867 (N_2867,N_2835,N_2839);
and U2868 (N_2868,N_2808,N_2812);
nand U2869 (N_2869,N_2821,N_2805);
nor U2870 (N_2870,N_2848,N_2849);
nor U2871 (N_2871,N_2820,N_2840);
or U2872 (N_2872,N_2832,N_2836);
xnor U2873 (N_2873,N_2822,N_2843);
xor U2874 (N_2874,N_2831,N_2837);
nor U2875 (N_2875,N_2843,N_2812);
or U2876 (N_2876,N_2817,N_2808);
nand U2877 (N_2877,N_2839,N_2806);
xnor U2878 (N_2878,N_2802,N_2803);
or U2879 (N_2879,N_2824,N_2846);
and U2880 (N_2880,N_2821,N_2825);
xnor U2881 (N_2881,N_2800,N_2809);
nand U2882 (N_2882,N_2835,N_2826);
nand U2883 (N_2883,N_2821,N_2801);
or U2884 (N_2884,N_2818,N_2815);
or U2885 (N_2885,N_2807,N_2824);
nand U2886 (N_2886,N_2830,N_2821);
xor U2887 (N_2887,N_2842,N_2843);
and U2888 (N_2888,N_2803,N_2844);
or U2889 (N_2889,N_2842,N_2800);
or U2890 (N_2890,N_2805,N_2842);
nor U2891 (N_2891,N_2823,N_2802);
xor U2892 (N_2892,N_2834,N_2837);
nor U2893 (N_2893,N_2815,N_2804);
xnor U2894 (N_2894,N_2826,N_2815);
nor U2895 (N_2895,N_2847,N_2849);
nand U2896 (N_2896,N_2834,N_2848);
or U2897 (N_2897,N_2811,N_2834);
and U2898 (N_2898,N_2847,N_2821);
xor U2899 (N_2899,N_2835,N_2810);
nor U2900 (N_2900,N_2886,N_2885);
or U2901 (N_2901,N_2887,N_2899);
nor U2902 (N_2902,N_2850,N_2874);
and U2903 (N_2903,N_2868,N_2857);
or U2904 (N_2904,N_2881,N_2864);
and U2905 (N_2905,N_2876,N_2862);
xnor U2906 (N_2906,N_2873,N_2895);
or U2907 (N_2907,N_2871,N_2880);
or U2908 (N_2908,N_2882,N_2851);
nand U2909 (N_2909,N_2860,N_2890);
and U2910 (N_2910,N_2866,N_2869);
xor U2911 (N_2911,N_2877,N_2891);
nor U2912 (N_2912,N_2884,N_2888);
nor U2913 (N_2913,N_2896,N_2879);
nor U2914 (N_2914,N_2897,N_2852);
nand U2915 (N_2915,N_2861,N_2893);
and U2916 (N_2916,N_2898,N_2863);
and U2917 (N_2917,N_2872,N_2894);
xnor U2918 (N_2918,N_2883,N_2858);
nor U2919 (N_2919,N_2855,N_2870);
xnor U2920 (N_2920,N_2875,N_2867);
xor U2921 (N_2921,N_2853,N_2892);
and U2922 (N_2922,N_2878,N_2889);
xor U2923 (N_2923,N_2854,N_2865);
nor U2924 (N_2924,N_2856,N_2859);
nor U2925 (N_2925,N_2865,N_2895);
nor U2926 (N_2926,N_2860,N_2889);
nor U2927 (N_2927,N_2874,N_2896);
or U2928 (N_2928,N_2872,N_2880);
xor U2929 (N_2929,N_2869,N_2890);
nand U2930 (N_2930,N_2878,N_2852);
or U2931 (N_2931,N_2888,N_2870);
nand U2932 (N_2932,N_2867,N_2850);
or U2933 (N_2933,N_2854,N_2893);
and U2934 (N_2934,N_2871,N_2850);
or U2935 (N_2935,N_2860,N_2875);
and U2936 (N_2936,N_2851,N_2863);
or U2937 (N_2937,N_2889,N_2850);
and U2938 (N_2938,N_2850,N_2890);
nand U2939 (N_2939,N_2885,N_2899);
or U2940 (N_2940,N_2857,N_2853);
nor U2941 (N_2941,N_2875,N_2877);
or U2942 (N_2942,N_2857,N_2874);
xnor U2943 (N_2943,N_2888,N_2868);
and U2944 (N_2944,N_2865,N_2875);
nand U2945 (N_2945,N_2863,N_2856);
and U2946 (N_2946,N_2877,N_2871);
and U2947 (N_2947,N_2881,N_2883);
xor U2948 (N_2948,N_2852,N_2856);
nor U2949 (N_2949,N_2865,N_2891);
and U2950 (N_2950,N_2944,N_2927);
and U2951 (N_2951,N_2902,N_2919);
xnor U2952 (N_2952,N_2947,N_2935);
nor U2953 (N_2953,N_2941,N_2912);
nor U2954 (N_2954,N_2913,N_2946);
nand U2955 (N_2955,N_2948,N_2939);
or U2956 (N_2956,N_2907,N_2925);
and U2957 (N_2957,N_2940,N_2932);
or U2958 (N_2958,N_2900,N_2906);
and U2959 (N_2959,N_2911,N_2915);
or U2960 (N_2960,N_2917,N_2924);
or U2961 (N_2961,N_2904,N_2909);
nand U2962 (N_2962,N_2922,N_2936);
and U2963 (N_2963,N_2949,N_2908);
or U2964 (N_2964,N_2929,N_2905);
or U2965 (N_2965,N_2938,N_2920);
xor U2966 (N_2966,N_2933,N_2930);
xnor U2967 (N_2967,N_2921,N_2910);
nor U2968 (N_2968,N_2916,N_2934);
nor U2969 (N_2969,N_2918,N_2926);
nand U2970 (N_2970,N_2945,N_2943);
xor U2971 (N_2971,N_2901,N_2928);
xnor U2972 (N_2972,N_2942,N_2923);
and U2973 (N_2973,N_2914,N_2931);
nor U2974 (N_2974,N_2903,N_2937);
nor U2975 (N_2975,N_2910,N_2920);
nand U2976 (N_2976,N_2939,N_2928);
and U2977 (N_2977,N_2933,N_2912);
or U2978 (N_2978,N_2929,N_2904);
or U2979 (N_2979,N_2909,N_2947);
nor U2980 (N_2980,N_2912,N_2900);
or U2981 (N_2981,N_2941,N_2909);
or U2982 (N_2982,N_2920,N_2924);
nand U2983 (N_2983,N_2940,N_2939);
xnor U2984 (N_2984,N_2936,N_2912);
nor U2985 (N_2985,N_2901,N_2922);
xor U2986 (N_2986,N_2905,N_2908);
nor U2987 (N_2987,N_2910,N_2940);
nor U2988 (N_2988,N_2922,N_2943);
xor U2989 (N_2989,N_2940,N_2925);
xor U2990 (N_2990,N_2940,N_2924);
nand U2991 (N_2991,N_2918,N_2904);
nor U2992 (N_2992,N_2945,N_2908);
nand U2993 (N_2993,N_2908,N_2904);
or U2994 (N_2994,N_2949,N_2922);
nand U2995 (N_2995,N_2902,N_2941);
and U2996 (N_2996,N_2916,N_2936);
xor U2997 (N_2997,N_2945,N_2924);
nor U2998 (N_2998,N_2929,N_2919);
nor U2999 (N_2999,N_2917,N_2948);
nor UO_0 (O_0,N_2958,N_2970);
xnor UO_1 (O_1,N_2973,N_2954);
and UO_2 (O_2,N_2984,N_2994);
nor UO_3 (O_3,N_2950,N_2961);
and UO_4 (O_4,N_2988,N_2999);
or UO_5 (O_5,N_2996,N_2965);
nor UO_6 (O_6,N_2963,N_2977);
nand UO_7 (O_7,N_2966,N_2985);
or UO_8 (O_8,N_2952,N_2976);
or UO_9 (O_9,N_2971,N_2987);
xnor UO_10 (O_10,N_2991,N_2980);
xor UO_11 (O_11,N_2962,N_2995);
nor UO_12 (O_12,N_2986,N_2959);
or UO_13 (O_13,N_2957,N_2979);
nor UO_14 (O_14,N_2960,N_2951);
and UO_15 (O_15,N_2953,N_2997);
nand UO_16 (O_16,N_2982,N_2981);
xor UO_17 (O_17,N_2983,N_2964);
nor UO_18 (O_18,N_2978,N_2975);
xor UO_19 (O_19,N_2992,N_2955);
nor UO_20 (O_20,N_2969,N_2967);
and UO_21 (O_21,N_2989,N_2998);
xnor UO_22 (O_22,N_2956,N_2968);
or UO_23 (O_23,N_2990,N_2993);
nor UO_24 (O_24,N_2974,N_2972);
or UO_25 (O_25,N_2990,N_2956);
nor UO_26 (O_26,N_2956,N_2969);
or UO_27 (O_27,N_2957,N_2970);
nand UO_28 (O_28,N_2989,N_2983);
or UO_29 (O_29,N_2968,N_2986);
nand UO_30 (O_30,N_2979,N_2970);
or UO_31 (O_31,N_2952,N_2997);
nand UO_32 (O_32,N_2957,N_2988);
xnor UO_33 (O_33,N_2989,N_2992);
and UO_34 (O_34,N_2990,N_2957);
or UO_35 (O_35,N_2982,N_2960);
nand UO_36 (O_36,N_2987,N_2967);
or UO_37 (O_37,N_2951,N_2998);
and UO_38 (O_38,N_2987,N_2965);
xor UO_39 (O_39,N_2959,N_2973);
nor UO_40 (O_40,N_2951,N_2975);
and UO_41 (O_41,N_2996,N_2985);
xnor UO_42 (O_42,N_2983,N_2971);
nor UO_43 (O_43,N_2973,N_2956);
and UO_44 (O_44,N_2996,N_2972);
or UO_45 (O_45,N_2986,N_2955);
and UO_46 (O_46,N_2996,N_2950);
nor UO_47 (O_47,N_2953,N_2959);
nand UO_48 (O_48,N_2986,N_2966);
and UO_49 (O_49,N_2989,N_2952);
nor UO_50 (O_50,N_2962,N_2954);
xor UO_51 (O_51,N_2986,N_2963);
nor UO_52 (O_52,N_2960,N_2952);
and UO_53 (O_53,N_2975,N_2966);
or UO_54 (O_54,N_2960,N_2957);
nor UO_55 (O_55,N_2977,N_2998);
and UO_56 (O_56,N_2980,N_2988);
or UO_57 (O_57,N_2978,N_2980);
nand UO_58 (O_58,N_2992,N_2987);
nand UO_59 (O_59,N_2962,N_2951);
nand UO_60 (O_60,N_2974,N_2990);
nor UO_61 (O_61,N_2968,N_2962);
or UO_62 (O_62,N_2991,N_2967);
nand UO_63 (O_63,N_2985,N_2971);
or UO_64 (O_64,N_2985,N_2963);
and UO_65 (O_65,N_2993,N_2998);
xor UO_66 (O_66,N_2995,N_2981);
nor UO_67 (O_67,N_2982,N_2967);
nor UO_68 (O_68,N_2969,N_2986);
or UO_69 (O_69,N_2983,N_2991);
xor UO_70 (O_70,N_2983,N_2965);
or UO_71 (O_71,N_2997,N_2996);
xnor UO_72 (O_72,N_2979,N_2981);
and UO_73 (O_73,N_2952,N_2955);
nand UO_74 (O_74,N_2979,N_2983);
xor UO_75 (O_75,N_2989,N_2967);
and UO_76 (O_76,N_2974,N_2975);
nand UO_77 (O_77,N_2970,N_2984);
and UO_78 (O_78,N_2994,N_2958);
and UO_79 (O_79,N_2970,N_2972);
and UO_80 (O_80,N_2993,N_2969);
nor UO_81 (O_81,N_2971,N_2962);
or UO_82 (O_82,N_2962,N_2987);
xnor UO_83 (O_83,N_2981,N_2989);
nand UO_84 (O_84,N_2956,N_2963);
xnor UO_85 (O_85,N_2956,N_2999);
and UO_86 (O_86,N_2962,N_2950);
or UO_87 (O_87,N_2979,N_2987);
nand UO_88 (O_88,N_2957,N_2973);
nand UO_89 (O_89,N_2957,N_2994);
xor UO_90 (O_90,N_2952,N_2982);
and UO_91 (O_91,N_2991,N_2952);
or UO_92 (O_92,N_2969,N_2975);
and UO_93 (O_93,N_2978,N_2996);
or UO_94 (O_94,N_2950,N_2979);
or UO_95 (O_95,N_2961,N_2951);
xnor UO_96 (O_96,N_2978,N_2990);
nand UO_97 (O_97,N_2974,N_2983);
and UO_98 (O_98,N_2994,N_2961);
xnor UO_99 (O_99,N_2998,N_2983);
nor UO_100 (O_100,N_2988,N_2956);
and UO_101 (O_101,N_2958,N_2963);
or UO_102 (O_102,N_2955,N_2995);
nand UO_103 (O_103,N_2993,N_2972);
and UO_104 (O_104,N_2964,N_2982);
and UO_105 (O_105,N_2968,N_2982);
nor UO_106 (O_106,N_2986,N_2978);
and UO_107 (O_107,N_2962,N_2958);
and UO_108 (O_108,N_2967,N_2981);
and UO_109 (O_109,N_2997,N_2960);
nor UO_110 (O_110,N_2963,N_2980);
nand UO_111 (O_111,N_2963,N_2983);
nand UO_112 (O_112,N_2959,N_2971);
or UO_113 (O_113,N_2983,N_2969);
and UO_114 (O_114,N_2985,N_2979);
and UO_115 (O_115,N_2961,N_2980);
and UO_116 (O_116,N_2966,N_2967);
nor UO_117 (O_117,N_2961,N_2989);
or UO_118 (O_118,N_2961,N_2974);
nor UO_119 (O_119,N_2966,N_2964);
nor UO_120 (O_120,N_2974,N_2969);
or UO_121 (O_121,N_2980,N_2985);
or UO_122 (O_122,N_2999,N_2958);
or UO_123 (O_123,N_2961,N_2993);
xnor UO_124 (O_124,N_2994,N_2951);
and UO_125 (O_125,N_2965,N_2955);
nand UO_126 (O_126,N_2998,N_2972);
xnor UO_127 (O_127,N_2965,N_2984);
and UO_128 (O_128,N_2954,N_2957);
xnor UO_129 (O_129,N_2951,N_2992);
xnor UO_130 (O_130,N_2975,N_2982);
nand UO_131 (O_131,N_2986,N_2957);
xor UO_132 (O_132,N_2988,N_2952);
and UO_133 (O_133,N_2952,N_2972);
and UO_134 (O_134,N_2968,N_2958);
and UO_135 (O_135,N_2954,N_2952);
and UO_136 (O_136,N_2990,N_2994);
or UO_137 (O_137,N_2984,N_2997);
or UO_138 (O_138,N_2979,N_2973);
nand UO_139 (O_139,N_2997,N_2970);
and UO_140 (O_140,N_2971,N_2980);
nand UO_141 (O_141,N_2971,N_2979);
xor UO_142 (O_142,N_2982,N_2970);
xor UO_143 (O_143,N_2986,N_2958);
nor UO_144 (O_144,N_2954,N_2990);
nor UO_145 (O_145,N_2980,N_2957);
nor UO_146 (O_146,N_2961,N_2995);
nand UO_147 (O_147,N_2973,N_2970);
xor UO_148 (O_148,N_2965,N_2993);
and UO_149 (O_149,N_2959,N_2964);
and UO_150 (O_150,N_2969,N_2992);
xnor UO_151 (O_151,N_2955,N_2950);
and UO_152 (O_152,N_2968,N_2963);
and UO_153 (O_153,N_2976,N_2980);
nand UO_154 (O_154,N_2957,N_2989);
and UO_155 (O_155,N_2957,N_2978);
xnor UO_156 (O_156,N_2982,N_2987);
xnor UO_157 (O_157,N_2968,N_2960);
nor UO_158 (O_158,N_2965,N_2981);
nor UO_159 (O_159,N_2991,N_2953);
nor UO_160 (O_160,N_2969,N_2951);
and UO_161 (O_161,N_2996,N_2961);
xor UO_162 (O_162,N_2958,N_2971);
nand UO_163 (O_163,N_2958,N_2966);
or UO_164 (O_164,N_2973,N_2988);
xnor UO_165 (O_165,N_2971,N_2996);
and UO_166 (O_166,N_2959,N_2985);
or UO_167 (O_167,N_2997,N_2977);
and UO_168 (O_168,N_2978,N_2951);
nand UO_169 (O_169,N_2982,N_2983);
or UO_170 (O_170,N_2963,N_2979);
and UO_171 (O_171,N_2958,N_2952);
xnor UO_172 (O_172,N_2974,N_2998);
nand UO_173 (O_173,N_2987,N_2980);
nor UO_174 (O_174,N_2996,N_2967);
and UO_175 (O_175,N_2969,N_2977);
or UO_176 (O_176,N_2953,N_2967);
and UO_177 (O_177,N_2965,N_2986);
nor UO_178 (O_178,N_2968,N_2983);
nand UO_179 (O_179,N_2965,N_2969);
nand UO_180 (O_180,N_2976,N_2994);
or UO_181 (O_181,N_2972,N_2967);
nand UO_182 (O_182,N_2979,N_2994);
or UO_183 (O_183,N_2958,N_2956);
nand UO_184 (O_184,N_2979,N_2977);
nor UO_185 (O_185,N_2963,N_2967);
and UO_186 (O_186,N_2967,N_2973);
xor UO_187 (O_187,N_2995,N_2960);
xnor UO_188 (O_188,N_2984,N_2950);
nand UO_189 (O_189,N_2981,N_2987);
nor UO_190 (O_190,N_2997,N_2971);
or UO_191 (O_191,N_2977,N_2988);
or UO_192 (O_192,N_2988,N_2984);
nand UO_193 (O_193,N_2990,N_2981);
or UO_194 (O_194,N_2999,N_2980);
xnor UO_195 (O_195,N_2983,N_2955);
xnor UO_196 (O_196,N_2959,N_2989);
and UO_197 (O_197,N_2964,N_2977);
and UO_198 (O_198,N_2977,N_2986);
nand UO_199 (O_199,N_2953,N_2990);
nand UO_200 (O_200,N_2959,N_2962);
or UO_201 (O_201,N_2950,N_2997);
nand UO_202 (O_202,N_2997,N_2962);
nand UO_203 (O_203,N_2952,N_2957);
or UO_204 (O_204,N_2980,N_2997);
xnor UO_205 (O_205,N_2962,N_2952);
and UO_206 (O_206,N_2955,N_2976);
nor UO_207 (O_207,N_2982,N_2980);
and UO_208 (O_208,N_2960,N_2986);
and UO_209 (O_209,N_2990,N_2965);
xnor UO_210 (O_210,N_2997,N_2978);
nor UO_211 (O_211,N_2954,N_2996);
or UO_212 (O_212,N_2997,N_2999);
nand UO_213 (O_213,N_2977,N_2980);
nand UO_214 (O_214,N_2981,N_2988);
and UO_215 (O_215,N_2976,N_2990);
xnor UO_216 (O_216,N_2983,N_2994);
nand UO_217 (O_217,N_2973,N_2999);
nand UO_218 (O_218,N_2969,N_2990);
nor UO_219 (O_219,N_2996,N_2963);
nand UO_220 (O_220,N_2991,N_2989);
nand UO_221 (O_221,N_2958,N_2995);
and UO_222 (O_222,N_2972,N_2963);
nand UO_223 (O_223,N_2978,N_2962);
nor UO_224 (O_224,N_2976,N_2999);
nor UO_225 (O_225,N_2974,N_2997);
and UO_226 (O_226,N_2953,N_2979);
or UO_227 (O_227,N_2992,N_2976);
xor UO_228 (O_228,N_2964,N_2967);
xor UO_229 (O_229,N_2982,N_2963);
nor UO_230 (O_230,N_2953,N_2955);
or UO_231 (O_231,N_2986,N_2992);
xnor UO_232 (O_232,N_2975,N_2990);
nor UO_233 (O_233,N_2962,N_2994);
and UO_234 (O_234,N_2961,N_2998);
nor UO_235 (O_235,N_2979,N_2972);
and UO_236 (O_236,N_2973,N_2955);
nor UO_237 (O_237,N_2969,N_2979);
or UO_238 (O_238,N_2960,N_2955);
nor UO_239 (O_239,N_2965,N_2963);
and UO_240 (O_240,N_2960,N_2991);
nor UO_241 (O_241,N_2999,N_2964);
and UO_242 (O_242,N_2981,N_2955);
or UO_243 (O_243,N_2993,N_2959);
xnor UO_244 (O_244,N_2991,N_2999);
xor UO_245 (O_245,N_2984,N_2951);
or UO_246 (O_246,N_2958,N_2954);
xnor UO_247 (O_247,N_2989,N_2973);
or UO_248 (O_248,N_2970,N_2980);
and UO_249 (O_249,N_2981,N_2968);
or UO_250 (O_250,N_2962,N_2965);
or UO_251 (O_251,N_2964,N_2972);
and UO_252 (O_252,N_2973,N_2963);
and UO_253 (O_253,N_2985,N_2997);
xnor UO_254 (O_254,N_2988,N_2979);
nand UO_255 (O_255,N_2954,N_2950);
nand UO_256 (O_256,N_2962,N_2956);
nand UO_257 (O_257,N_2989,N_2994);
and UO_258 (O_258,N_2971,N_2969);
nor UO_259 (O_259,N_2967,N_2992);
or UO_260 (O_260,N_2995,N_2985);
nor UO_261 (O_261,N_2983,N_2962);
or UO_262 (O_262,N_2987,N_2964);
and UO_263 (O_263,N_2973,N_2987);
and UO_264 (O_264,N_2957,N_2961);
nor UO_265 (O_265,N_2986,N_2961);
or UO_266 (O_266,N_2994,N_2972);
and UO_267 (O_267,N_2998,N_2992);
xor UO_268 (O_268,N_2974,N_2953);
nor UO_269 (O_269,N_2954,N_2970);
xor UO_270 (O_270,N_2993,N_2996);
nand UO_271 (O_271,N_2984,N_2990);
nand UO_272 (O_272,N_2966,N_2996);
or UO_273 (O_273,N_2961,N_2966);
nand UO_274 (O_274,N_2964,N_2995);
and UO_275 (O_275,N_2962,N_2961);
nand UO_276 (O_276,N_2994,N_2995);
nand UO_277 (O_277,N_2966,N_2972);
nor UO_278 (O_278,N_2993,N_2999);
and UO_279 (O_279,N_2956,N_2964);
nand UO_280 (O_280,N_2979,N_2984);
and UO_281 (O_281,N_2990,N_2958);
and UO_282 (O_282,N_2950,N_2969);
or UO_283 (O_283,N_2995,N_2988);
or UO_284 (O_284,N_2967,N_2965);
nand UO_285 (O_285,N_2971,N_2999);
and UO_286 (O_286,N_2968,N_2976);
nor UO_287 (O_287,N_2958,N_2975);
xor UO_288 (O_288,N_2951,N_2957);
nor UO_289 (O_289,N_2976,N_2998);
and UO_290 (O_290,N_2950,N_2991);
xor UO_291 (O_291,N_2952,N_2978);
nor UO_292 (O_292,N_2989,N_2951);
nor UO_293 (O_293,N_2987,N_2954);
or UO_294 (O_294,N_2982,N_2985);
or UO_295 (O_295,N_2977,N_2987);
or UO_296 (O_296,N_2982,N_2976);
and UO_297 (O_297,N_2988,N_2965);
and UO_298 (O_298,N_2969,N_2954);
nand UO_299 (O_299,N_2958,N_2951);
and UO_300 (O_300,N_2952,N_2969);
xnor UO_301 (O_301,N_2995,N_2952);
and UO_302 (O_302,N_2960,N_2963);
and UO_303 (O_303,N_2972,N_2983);
and UO_304 (O_304,N_2956,N_2993);
nor UO_305 (O_305,N_2966,N_2987);
and UO_306 (O_306,N_2998,N_2984);
and UO_307 (O_307,N_2958,N_2984);
or UO_308 (O_308,N_2979,N_2951);
and UO_309 (O_309,N_2968,N_2994);
xor UO_310 (O_310,N_2992,N_2991);
and UO_311 (O_311,N_2987,N_2972);
or UO_312 (O_312,N_2980,N_2965);
xor UO_313 (O_313,N_2954,N_2971);
xnor UO_314 (O_314,N_2953,N_2976);
nor UO_315 (O_315,N_2978,N_2992);
xor UO_316 (O_316,N_2970,N_2966);
xnor UO_317 (O_317,N_2986,N_2991);
nand UO_318 (O_318,N_2977,N_2985);
or UO_319 (O_319,N_2957,N_2991);
nor UO_320 (O_320,N_2985,N_2972);
or UO_321 (O_321,N_2978,N_2956);
xnor UO_322 (O_322,N_2968,N_2952);
or UO_323 (O_323,N_2969,N_2991);
nand UO_324 (O_324,N_2956,N_2977);
and UO_325 (O_325,N_2981,N_2977);
xnor UO_326 (O_326,N_2987,N_2961);
nor UO_327 (O_327,N_2987,N_2958);
xnor UO_328 (O_328,N_2975,N_2953);
nand UO_329 (O_329,N_2977,N_2958);
or UO_330 (O_330,N_2975,N_2962);
nand UO_331 (O_331,N_2998,N_2954);
or UO_332 (O_332,N_2976,N_2978);
nand UO_333 (O_333,N_2984,N_2999);
xnor UO_334 (O_334,N_2978,N_2963);
or UO_335 (O_335,N_2976,N_2979);
xnor UO_336 (O_336,N_2989,N_2995);
and UO_337 (O_337,N_2997,N_2993);
and UO_338 (O_338,N_2998,N_2994);
nor UO_339 (O_339,N_2960,N_2998);
xor UO_340 (O_340,N_2995,N_2991);
and UO_341 (O_341,N_2954,N_2966);
nand UO_342 (O_342,N_2976,N_2981);
nor UO_343 (O_343,N_2993,N_2966);
or UO_344 (O_344,N_2955,N_2963);
or UO_345 (O_345,N_2957,N_2962);
xor UO_346 (O_346,N_2995,N_2987);
and UO_347 (O_347,N_2968,N_2971);
nand UO_348 (O_348,N_2956,N_2971);
xnor UO_349 (O_349,N_2992,N_2995);
and UO_350 (O_350,N_2964,N_2984);
nor UO_351 (O_351,N_2993,N_2955);
nand UO_352 (O_352,N_2969,N_2953);
or UO_353 (O_353,N_2958,N_2978);
nand UO_354 (O_354,N_2958,N_2976);
and UO_355 (O_355,N_2978,N_2989);
xor UO_356 (O_356,N_2993,N_2989);
xor UO_357 (O_357,N_2959,N_2955);
nand UO_358 (O_358,N_2998,N_2971);
or UO_359 (O_359,N_2972,N_2982);
and UO_360 (O_360,N_2951,N_2974);
nand UO_361 (O_361,N_2959,N_2976);
xor UO_362 (O_362,N_2990,N_2955);
or UO_363 (O_363,N_2970,N_2999);
and UO_364 (O_364,N_2960,N_2996);
or UO_365 (O_365,N_2965,N_2972);
and UO_366 (O_366,N_2960,N_2989);
xor UO_367 (O_367,N_2966,N_2963);
or UO_368 (O_368,N_2980,N_2995);
and UO_369 (O_369,N_2975,N_2993);
nand UO_370 (O_370,N_2969,N_2961);
xor UO_371 (O_371,N_2951,N_2952);
and UO_372 (O_372,N_2992,N_2952);
nand UO_373 (O_373,N_2955,N_2967);
xnor UO_374 (O_374,N_2963,N_2988);
and UO_375 (O_375,N_2976,N_2961);
xnor UO_376 (O_376,N_2999,N_2985);
xnor UO_377 (O_377,N_2978,N_2966);
xor UO_378 (O_378,N_2987,N_2998);
nand UO_379 (O_379,N_2978,N_2988);
xnor UO_380 (O_380,N_2981,N_2963);
xor UO_381 (O_381,N_2994,N_2980);
xor UO_382 (O_382,N_2963,N_2951);
and UO_383 (O_383,N_2980,N_2967);
xor UO_384 (O_384,N_2993,N_2995);
and UO_385 (O_385,N_2987,N_2993);
nor UO_386 (O_386,N_2950,N_2983);
nand UO_387 (O_387,N_2972,N_2999);
nand UO_388 (O_388,N_2950,N_2968);
xnor UO_389 (O_389,N_2989,N_2953);
nand UO_390 (O_390,N_2964,N_2978);
and UO_391 (O_391,N_2983,N_2997);
and UO_392 (O_392,N_2961,N_2960);
xnor UO_393 (O_393,N_2968,N_2954);
xor UO_394 (O_394,N_2991,N_2990);
and UO_395 (O_395,N_2972,N_2950);
nand UO_396 (O_396,N_2999,N_2963);
xor UO_397 (O_397,N_2964,N_2994);
nand UO_398 (O_398,N_2959,N_2961);
or UO_399 (O_399,N_2958,N_2972);
and UO_400 (O_400,N_2960,N_2976);
nand UO_401 (O_401,N_2981,N_2986);
and UO_402 (O_402,N_2980,N_2964);
xor UO_403 (O_403,N_2997,N_2951);
or UO_404 (O_404,N_2951,N_2988);
xor UO_405 (O_405,N_2977,N_2955);
or UO_406 (O_406,N_2981,N_2992);
nand UO_407 (O_407,N_2965,N_2956);
or UO_408 (O_408,N_2987,N_2960);
or UO_409 (O_409,N_2988,N_2986);
nor UO_410 (O_410,N_2996,N_2989);
or UO_411 (O_411,N_2967,N_2976);
nand UO_412 (O_412,N_2993,N_2963);
xnor UO_413 (O_413,N_2977,N_2990);
or UO_414 (O_414,N_2979,N_2990);
nand UO_415 (O_415,N_2988,N_2950);
or UO_416 (O_416,N_2982,N_2988);
xnor UO_417 (O_417,N_2997,N_2966);
xnor UO_418 (O_418,N_2960,N_2971);
xor UO_419 (O_419,N_2970,N_2991);
and UO_420 (O_420,N_2959,N_2968);
nand UO_421 (O_421,N_2955,N_2970);
and UO_422 (O_422,N_2959,N_2984);
nor UO_423 (O_423,N_2955,N_2991);
and UO_424 (O_424,N_2953,N_2965);
nand UO_425 (O_425,N_2984,N_2974);
and UO_426 (O_426,N_2990,N_2980);
xor UO_427 (O_427,N_2997,N_2958);
nand UO_428 (O_428,N_2987,N_2994);
or UO_429 (O_429,N_2977,N_2982);
nor UO_430 (O_430,N_2972,N_2973);
nor UO_431 (O_431,N_2959,N_2969);
xnor UO_432 (O_432,N_2974,N_2970);
or UO_433 (O_433,N_2950,N_2974);
xnor UO_434 (O_434,N_2973,N_2998);
or UO_435 (O_435,N_2976,N_2972);
or UO_436 (O_436,N_2987,N_2976);
and UO_437 (O_437,N_2978,N_2983);
and UO_438 (O_438,N_2953,N_2999);
nand UO_439 (O_439,N_2951,N_2967);
or UO_440 (O_440,N_2992,N_2963);
and UO_441 (O_441,N_2971,N_2963);
and UO_442 (O_442,N_2989,N_2958);
and UO_443 (O_443,N_2965,N_2968);
or UO_444 (O_444,N_2953,N_2985);
nor UO_445 (O_445,N_2954,N_2984);
nand UO_446 (O_446,N_2965,N_2952);
and UO_447 (O_447,N_2958,N_2973);
or UO_448 (O_448,N_2956,N_2975);
nand UO_449 (O_449,N_2961,N_2973);
and UO_450 (O_450,N_2970,N_2962);
or UO_451 (O_451,N_2987,N_2983);
and UO_452 (O_452,N_2991,N_2963);
nor UO_453 (O_453,N_2952,N_2981);
nor UO_454 (O_454,N_2966,N_2999);
nand UO_455 (O_455,N_2990,N_2983);
and UO_456 (O_456,N_2966,N_2952);
nand UO_457 (O_457,N_2990,N_2951);
nand UO_458 (O_458,N_2953,N_2962);
nor UO_459 (O_459,N_2997,N_2954);
and UO_460 (O_460,N_2963,N_2970);
xor UO_461 (O_461,N_2957,N_2975);
nand UO_462 (O_462,N_2988,N_2970);
xnor UO_463 (O_463,N_2951,N_2970);
and UO_464 (O_464,N_2974,N_2980);
xor UO_465 (O_465,N_2979,N_2986);
and UO_466 (O_466,N_2970,N_2953);
nand UO_467 (O_467,N_2956,N_2992);
nand UO_468 (O_468,N_2983,N_2977);
or UO_469 (O_469,N_2975,N_2983);
nor UO_470 (O_470,N_2999,N_2994);
or UO_471 (O_471,N_2999,N_2954);
and UO_472 (O_472,N_2957,N_2959);
xor UO_473 (O_473,N_2999,N_2998);
or UO_474 (O_474,N_2981,N_2956);
nand UO_475 (O_475,N_2968,N_2989);
and UO_476 (O_476,N_2969,N_2973);
xnor UO_477 (O_477,N_2993,N_2982);
nor UO_478 (O_478,N_2951,N_2973);
or UO_479 (O_479,N_2959,N_2960);
xor UO_480 (O_480,N_2985,N_2986);
and UO_481 (O_481,N_2976,N_2962);
xnor UO_482 (O_482,N_2969,N_2972);
or UO_483 (O_483,N_2993,N_2983);
and UO_484 (O_484,N_2976,N_2984);
or UO_485 (O_485,N_2990,N_2971);
nor UO_486 (O_486,N_2969,N_2994);
or UO_487 (O_487,N_2955,N_2957);
xnor UO_488 (O_488,N_2997,N_2998);
nor UO_489 (O_489,N_2962,N_2992);
xnor UO_490 (O_490,N_2986,N_2984);
nor UO_491 (O_491,N_2954,N_2985);
nor UO_492 (O_492,N_2995,N_2971);
nor UO_493 (O_493,N_2971,N_2957);
xor UO_494 (O_494,N_2988,N_2991);
nor UO_495 (O_495,N_2974,N_2954);
and UO_496 (O_496,N_2951,N_2985);
and UO_497 (O_497,N_2972,N_2954);
nand UO_498 (O_498,N_2985,N_2981);
and UO_499 (O_499,N_2981,N_2984);
endmodule